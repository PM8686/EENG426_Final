magic
tech sky130l
timestamp 1731220585
<< m1 >>
rect 3008 3599 3012 3635
rect 1176 3495 1180 3531
rect 1304 3439 1308 3471
rect 2408 3435 2412 3475
rect 976 3331 980 3367
rect 352 3175 356 3211
rect 848 3119 852 3171
rect 2984 2919 2988 2975
rect 240 2623 244 2655
rect 736 2623 740 2655
rect 2096 2651 2100 2687
rect 2904 2651 2908 2687
rect 2672 2595 2676 2627
rect 2880 2483 2884 2527
rect 3128 2435 3132 2467
rect 2312 2327 2316 2363
rect 2424 2327 2428 2363
rect 2776 2311 2780 2355
rect 1168 2187 1172 2223
rect 2928 2171 2932 2207
rect 2864 1847 2868 1883
rect 2168 1783 2172 1815
rect 328 1671 332 1723
rect 2888 1623 2892 1655
rect 1616 1319 1620 1351
rect 1288 1135 1292 1207
rect 3088 1131 3092 1163
rect 792 927 796 1031
rect 2632 971 2636 1003
rect 536 715 540 751
rect 208 315 212 347
<< m2c >>
rect 3008 3635 3012 3639
rect 264 3631 268 3635
rect 392 3631 396 3635
rect 528 3631 532 3635
rect 664 3631 668 3635
rect 800 3631 804 3635
rect 936 3631 940 3635
rect 1080 3631 1084 3635
rect 1224 3631 1228 3635
rect 2184 3595 2188 3599
rect 2472 3595 2476 3599
rect 2760 3595 2764 3599
rect 3008 3595 3012 3599
rect 3048 3595 3052 3599
rect 1928 3583 1932 3587
rect 2008 3583 2012 3587
rect 2096 3583 2100 3587
rect 2200 3583 2204 3587
rect 2320 3583 2324 3587
rect 2448 3583 2452 3587
rect 2584 3583 2588 3587
rect 2720 3583 2724 3587
rect 2856 3583 2860 3587
rect 3000 3583 3004 3587
rect 3144 3583 3148 3587
rect 3288 3583 3292 3587
rect 648 3567 652 3571
rect 1208 3567 1212 3571
rect 1176 3531 1180 3535
rect 2568 3519 2572 3523
rect 2984 3519 2988 3523
rect 216 3491 220 3495
rect 336 3491 340 3495
rect 448 3491 452 3495
rect 560 3491 564 3495
rect 664 3491 668 3495
rect 768 3491 772 3495
rect 864 3491 868 3495
rect 952 3491 956 3495
rect 1040 3491 1044 3495
rect 1128 3491 1132 3495
rect 1176 3491 1180 3495
rect 1216 3491 1220 3495
rect 1304 3491 1308 3495
rect 1392 3491 1396 3495
rect 1480 3491 1484 3495
rect 2408 3475 2412 3479
rect 256 3471 260 3475
rect 392 3471 396 3475
rect 528 3471 532 3475
rect 648 3471 652 3475
rect 760 3471 764 3475
rect 864 3471 868 3475
rect 968 3471 972 3475
rect 1064 3471 1068 3475
rect 1160 3471 1164 3475
rect 1256 3471 1260 3475
rect 1304 3471 1308 3475
rect 1352 3471 1356 3475
rect 2000 3443 2004 3447
rect 2184 3443 2188 3447
rect 2368 3443 2372 3447
rect 1304 3435 1308 3439
rect 2544 3443 2548 3447
rect 2704 3443 2708 3447
rect 2856 3443 2860 3447
rect 2992 3443 2996 3447
rect 3112 3443 3116 3447
rect 3224 3443 3228 3447
rect 3336 3443 3340 3447
rect 3448 3443 3452 3447
rect 3536 3443 3540 3447
rect 2032 3431 2036 3435
rect 2152 3431 2156 3435
rect 2280 3431 2284 3435
rect 2408 3431 2412 3435
rect 2416 3431 2420 3435
rect 2560 3431 2564 3435
rect 2704 3431 2708 3435
rect 2856 3431 2860 3435
rect 3024 3431 3028 3435
rect 3192 3431 3196 3435
rect 3368 3431 3372 3435
rect 3536 3431 3540 3435
rect 240 3407 244 3411
rect 1336 3407 1340 3411
rect 976 3367 980 3371
rect 2688 3367 2692 3371
rect 248 3327 252 3331
rect 400 3327 404 3331
rect 544 3327 548 3331
rect 680 3327 684 3331
rect 808 3327 812 3331
rect 928 3327 932 3331
rect 976 3327 980 3331
rect 1048 3327 1052 3331
rect 1160 3327 1164 3331
rect 1272 3327 1276 3331
rect 1384 3327 1388 3331
rect 232 3311 236 3315
rect 392 3311 396 3315
rect 544 3311 548 3315
rect 696 3311 700 3315
rect 840 3311 844 3315
rect 976 3311 980 3315
rect 1112 3311 1116 3315
rect 1240 3311 1244 3315
rect 1368 3311 1372 3315
rect 1496 3311 1500 3315
rect 2048 3291 2052 3295
rect 2184 3291 2188 3295
rect 2328 3291 2332 3295
rect 2472 3291 2476 3295
rect 2616 3291 2620 3295
rect 2760 3291 2764 3295
rect 2904 3291 2908 3295
rect 3056 3291 3060 3295
rect 3216 3291 3220 3295
rect 3384 3291 3388 3295
rect 3536 3291 3540 3295
rect 1952 3279 1956 3283
rect 2088 3279 2092 3283
rect 2216 3279 2220 3283
rect 2344 3279 2348 3283
rect 2472 3279 2476 3283
rect 2616 3279 2620 3283
rect 2768 3279 2772 3283
rect 2944 3279 2948 3283
rect 3136 3279 3140 3283
rect 3336 3279 3340 3283
rect 3536 3279 3540 3283
rect 1480 3247 1484 3251
rect 2328 3215 2332 3219
rect 352 3211 356 3215
rect 168 3171 172 3175
rect 304 3171 308 3175
rect 352 3171 356 3175
rect 448 3171 452 3175
rect 608 3171 612 3175
rect 768 3171 772 3175
rect 848 3171 852 3175
rect 928 3171 932 3175
rect 1080 3171 1084 3175
rect 1224 3171 1228 3175
rect 1360 3171 1364 3175
rect 1496 3171 1500 3175
rect 1640 3171 1644 3175
rect 200 3151 204 3155
rect 344 3151 348 3155
rect 488 3151 492 3155
rect 632 3151 636 3155
rect 768 3151 772 3155
rect 896 3151 900 3155
rect 1016 3151 1020 3155
rect 1128 3151 1132 3155
rect 1232 3151 1236 3155
rect 1336 3151 1340 3155
rect 1432 3151 1436 3155
rect 1520 3151 1524 3155
rect 1608 3151 1612 3155
rect 1696 3151 1700 3155
rect 1776 3151 1780 3155
rect 1928 3139 1932 3143
rect 2040 3139 2044 3143
rect 2176 3139 2180 3143
rect 2328 3139 2332 3143
rect 2488 3139 2492 3143
rect 2656 3139 2660 3143
rect 2832 3139 2836 3143
rect 3008 3139 3012 3143
rect 3184 3139 3188 3143
rect 3360 3139 3364 3143
rect 3536 3139 3540 3143
rect 1928 3127 1932 3131
rect 2096 3127 2100 3131
rect 2288 3127 2292 3131
rect 2480 3127 2484 3131
rect 2672 3127 2676 3131
rect 2856 3127 2860 3131
rect 3040 3127 3044 3131
rect 3224 3127 3228 3131
rect 3416 3127 3420 3131
rect 848 3115 852 3119
rect 2464 3063 2468 3067
rect 3400 3063 3404 3067
rect 168 2999 172 3003
rect 256 2999 260 3003
rect 360 2999 364 3003
rect 472 2999 476 3003
rect 584 2999 588 3003
rect 696 2999 700 3003
rect 184 2975 188 2979
rect 344 2975 348 2979
rect 512 2975 516 2979
rect 672 2975 676 2979
rect 824 2975 828 2979
rect 968 2975 972 2979
rect 1104 2975 1108 2979
rect 1224 2975 1228 2979
rect 1336 2975 1340 2979
rect 1448 2975 1452 2979
rect 1560 2975 1564 2979
rect 1672 2975 1676 2979
rect 2232 2975 2236 2979
rect 2368 2975 2372 2979
rect 2512 2975 2516 2979
rect 2656 2975 2660 2979
rect 2800 2975 2804 2979
rect 2936 2975 2940 2979
rect 2984 2975 2988 2979
rect 3072 2975 3076 2979
rect 3216 2975 3220 2979
rect 3360 2975 3364 2979
rect 2152 2951 2156 2955
rect 2232 2951 2236 2955
rect 2312 2951 2316 2955
rect 2392 2951 2396 2955
rect 2472 2951 2476 2955
rect 2552 2951 2556 2955
rect 2632 2951 2636 2955
rect 2720 2951 2724 2955
rect 2816 2951 2820 2955
rect 2936 2951 2940 2955
rect 3064 2951 3068 2955
rect 3208 2951 3212 2955
rect 3360 2951 3364 2955
rect 3520 2951 3524 2955
rect 2984 2915 2988 2919
rect 1656 2911 1660 2915
rect 2136 2887 2140 2891
rect 2800 2887 2804 2891
rect 3344 2887 3348 2891
rect 184 2835 188 2839
rect 344 2835 348 2839
rect 504 2835 508 2839
rect 664 2835 668 2839
rect 816 2835 820 2839
rect 960 2835 964 2839
rect 1088 2835 1092 2839
rect 1208 2835 1212 2839
rect 1320 2835 1324 2839
rect 1424 2835 1428 2839
rect 1520 2835 1524 2839
rect 1624 2835 1628 2839
rect 1728 2835 1732 2839
rect 168 2819 172 2823
rect 272 2819 276 2823
rect 408 2819 412 2823
rect 560 2819 564 2823
rect 712 2819 716 2823
rect 872 2819 876 2823
rect 1024 2819 1028 2823
rect 1168 2819 1172 2823
rect 1304 2819 1308 2823
rect 1432 2819 1436 2823
rect 1552 2819 1556 2823
rect 1672 2819 1676 2823
rect 1776 2819 1780 2823
rect 2080 2811 2084 2815
rect 2168 2811 2172 2815
rect 2272 2811 2276 2815
rect 2376 2811 2380 2815
rect 2496 2811 2500 2815
rect 2624 2811 2628 2815
rect 2760 2811 2764 2815
rect 2912 2811 2916 2815
rect 3064 2811 3068 2815
rect 3224 2811 3228 2815
rect 3392 2811 3396 2815
rect 3536 2811 3540 2815
rect 1928 2787 1932 2791
rect 2040 2787 2044 2791
rect 2192 2787 2196 2791
rect 2352 2787 2356 2791
rect 2512 2787 2516 2791
rect 2664 2787 2668 2791
rect 2816 2787 2820 2791
rect 2968 2787 2972 2791
rect 3112 2787 3116 2791
rect 3256 2787 3260 2791
rect 3408 2787 3412 2791
rect 3536 2787 3540 2791
rect 392 2755 396 2759
rect 1760 2755 1764 2759
rect 3240 2723 3244 2727
rect 2096 2687 2100 2691
rect 168 2675 172 2679
rect 264 2675 268 2679
rect 400 2675 404 2679
rect 544 2675 548 2679
rect 696 2675 700 2679
rect 848 2675 852 2679
rect 1008 2675 1012 2679
rect 1168 2675 1172 2679
rect 1320 2675 1324 2679
rect 1480 2675 1484 2679
rect 1640 2675 1644 2679
rect 1776 2675 1780 2679
rect 168 2655 172 2659
rect 240 2655 244 2659
rect 304 2655 308 2659
rect 472 2655 476 2659
rect 648 2655 652 2659
rect 736 2655 740 2659
rect 816 2655 820 2659
rect 976 2655 980 2659
rect 1128 2655 1132 2659
rect 1272 2655 1276 2659
rect 1424 2655 1428 2659
rect 1576 2655 1580 2659
rect 240 2619 244 2623
rect 2904 2687 2908 2691
rect 1928 2647 1932 2651
rect 2096 2647 2100 2651
rect 2136 2647 2140 2651
rect 2360 2647 2364 2651
rect 2568 2647 2572 2651
rect 2768 2647 2772 2651
rect 2904 2647 2908 2651
rect 2944 2647 2948 2651
rect 3104 2647 3108 2651
rect 3256 2647 3260 2651
rect 3408 2647 3412 2651
rect 3536 2647 3540 2651
rect 1928 2627 1932 2631
rect 2080 2627 2084 2631
rect 2288 2627 2292 2631
rect 2520 2627 2524 2631
rect 2672 2627 2676 2631
rect 2776 2627 2780 2631
rect 3040 2627 3044 2631
rect 3312 2627 3316 2631
rect 736 2619 740 2623
rect 456 2591 460 2595
rect 2672 2591 2676 2595
rect 2760 2563 2764 2567
rect 2880 2527 2884 2531
rect 168 2511 172 2515
rect 256 2511 260 2515
rect 400 2511 404 2515
rect 560 2511 564 2515
rect 736 2511 740 2515
rect 912 2511 916 2515
rect 1080 2511 1084 2515
rect 1240 2511 1244 2515
rect 1392 2511 1396 2515
rect 1544 2511 1548 2515
rect 1704 2511 1708 2515
rect 168 2495 172 2499
rect 248 2495 252 2499
rect 328 2495 332 2499
rect 416 2495 420 2499
rect 536 2495 540 2499
rect 672 2495 676 2499
rect 808 2495 812 2499
rect 952 2495 956 2499
rect 1088 2495 1092 2499
rect 1216 2495 1220 2499
rect 1336 2495 1340 2499
rect 1456 2495 1460 2499
rect 1576 2495 1580 2499
rect 1696 2495 1700 2499
rect 1928 2487 1932 2491
rect 2040 2487 2044 2491
rect 2192 2487 2196 2491
rect 2352 2487 2356 2491
rect 2504 2487 2508 2491
rect 2656 2487 2660 2491
rect 2792 2487 2796 2491
rect 2920 2487 2924 2491
rect 3040 2487 3044 2491
rect 3152 2487 3156 2491
rect 3256 2487 3260 2491
rect 3352 2487 3356 2491
rect 3456 2487 3460 2491
rect 3536 2487 3540 2491
rect 2880 2479 2884 2483
rect 2024 2467 2028 2471
rect 2152 2467 2156 2471
rect 2288 2467 2292 2471
rect 2432 2467 2436 2471
rect 2576 2467 2580 2471
rect 2728 2467 2732 2471
rect 2888 2467 2892 2471
rect 3048 2467 3052 2471
rect 3128 2467 3132 2471
rect 3216 2467 3220 2471
rect 3384 2467 3388 2471
rect 3536 2467 3540 2471
rect 3128 2431 3132 2435
rect 2560 2403 2564 2407
rect 2312 2363 2316 2367
rect 1096 2343 1100 2347
rect 1176 2343 1180 2347
rect 1256 2343 1260 2347
rect 1336 2343 1340 2347
rect 1416 2343 1420 2347
rect 1496 2343 1500 2347
rect 2424 2363 2428 2367
rect 2776 2355 2780 2359
rect 384 2323 388 2327
rect 464 2323 468 2327
rect 544 2323 548 2327
rect 624 2323 628 2327
rect 704 2323 708 2327
rect 784 2323 788 2327
rect 864 2323 868 2327
rect 944 2323 948 2327
rect 1024 2323 1028 2327
rect 1104 2323 1108 2327
rect 1184 2323 1188 2327
rect 1264 2323 1268 2327
rect 1344 2323 1348 2327
rect 2176 2323 2180 2327
rect 2272 2323 2276 2327
rect 2312 2323 2316 2327
rect 2376 2323 2380 2327
rect 2424 2323 2428 2327
rect 2488 2323 2492 2327
rect 2608 2323 2612 2327
rect 2736 2323 2740 2327
rect 2880 2323 2884 2327
rect 3040 2323 3044 2327
rect 3208 2323 3212 2327
rect 3384 2323 3388 2327
rect 3536 2323 3540 2327
rect 2304 2307 2308 2311
rect 2384 2307 2388 2311
rect 2464 2307 2468 2311
rect 2544 2307 2548 2311
rect 2624 2307 2628 2311
rect 2704 2307 2708 2311
rect 2776 2307 2780 2311
rect 2784 2307 2788 2311
rect 2872 2307 2876 2311
rect 2960 2307 2964 2311
rect 2528 2243 2532 2247
rect 1168 2223 1172 2227
rect 2928 2207 2932 2211
rect 408 2183 412 2187
rect 488 2183 492 2187
rect 568 2183 572 2187
rect 648 2183 652 2187
rect 728 2183 732 2187
rect 808 2183 812 2187
rect 888 2183 892 2187
rect 968 2183 972 2187
rect 1048 2183 1052 2187
rect 1128 2183 1132 2187
rect 1168 2183 1172 2187
rect 1208 2183 1212 2187
rect 1288 2183 1292 2187
rect 2344 2167 2348 2171
rect 2432 2167 2436 2171
rect 2528 2167 2532 2171
rect 2632 2167 2636 2171
rect 2752 2167 2756 2171
rect 2888 2167 2892 2171
rect 2928 2167 2932 2171
rect 3040 2167 3044 2171
rect 3208 2167 3212 2171
rect 3384 2167 3388 2171
rect 3536 2167 3540 2171
rect 336 2159 340 2163
rect 432 2159 436 2163
rect 528 2159 532 2163
rect 624 2159 628 2163
rect 712 2159 716 2163
rect 800 2159 804 2163
rect 888 2159 892 2163
rect 976 2159 980 2163
rect 1064 2159 1068 2163
rect 1152 2159 1156 2163
rect 1248 2159 1252 2163
rect 1928 2151 1932 2155
rect 2008 2151 2012 2155
rect 2136 2151 2140 2155
rect 2272 2151 2276 2155
rect 2416 2151 2420 2155
rect 2568 2151 2572 2155
rect 2720 2151 2724 2155
rect 2872 2151 2876 2155
rect 3032 2151 3036 2155
rect 3200 2151 3204 2155
rect 3376 2151 3380 2155
rect 3536 2151 3540 2155
rect 320 2095 324 2099
rect 1912 2087 1916 2091
rect 2552 2087 2556 2091
rect 3360 2087 3364 2091
rect 240 2007 244 2011
rect 360 2007 364 2011
rect 480 2007 484 2011
rect 608 2007 612 2011
rect 736 2007 740 2011
rect 856 2007 860 2011
rect 976 2007 980 2011
rect 1096 2007 1100 2011
rect 1208 2007 1212 2011
rect 1312 2007 1316 2011
rect 1408 2007 1412 2011
rect 1504 2007 1508 2011
rect 1600 2007 1604 2011
rect 1696 2007 1700 2011
rect 1776 2007 1780 2011
rect 2000 2003 2004 2007
rect 2248 2003 2252 2007
rect 2480 2003 2484 2007
rect 2688 2003 2692 2007
rect 2872 2003 2876 2007
rect 3032 2003 3036 2007
rect 3176 2003 3180 2007
rect 3304 2003 3308 2007
rect 3432 2003 3436 2007
rect 3536 2003 3540 2007
rect 216 1991 220 1995
rect 376 1991 380 1995
rect 544 1991 548 1995
rect 712 1991 716 1995
rect 880 1991 884 1995
rect 1040 1991 1044 1995
rect 1192 1991 1196 1995
rect 1336 1991 1340 1995
rect 1472 1991 1476 1995
rect 1608 1991 1612 1995
rect 1744 1991 1748 1995
rect 1984 1991 1988 1995
rect 2104 1991 2108 1995
rect 2224 1991 2228 1995
rect 2344 1991 2348 1995
rect 2472 1991 2476 1995
rect 2608 1991 2612 1995
rect 2768 1991 2772 1995
rect 2944 1991 2948 1995
rect 3144 1991 3148 1995
rect 3352 1991 3356 1995
rect 3536 1991 3540 1995
rect 200 1927 204 1931
rect 1728 1927 1732 1931
rect 2328 1927 2332 1931
rect 2456 1927 2460 1931
rect 2864 1883 2868 1887
rect 168 1847 172 1851
rect 272 1847 276 1851
rect 408 1847 412 1851
rect 560 1847 564 1851
rect 720 1847 724 1851
rect 880 1847 884 1851
rect 1040 1847 1044 1851
rect 1192 1847 1196 1851
rect 1336 1847 1340 1851
rect 1488 1847 1492 1851
rect 1640 1847 1644 1851
rect 2096 1843 2100 1847
rect 2184 1843 2188 1847
rect 2272 1843 2276 1847
rect 2352 1843 2356 1847
rect 2432 1843 2436 1847
rect 2520 1843 2524 1847
rect 2608 1843 2612 1847
rect 2696 1843 2700 1847
rect 2792 1843 2796 1847
rect 2864 1843 2868 1847
rect 2904 1843 2908 1847
rect 3024 1843 3028 1847
rect 3152 1843 3156 1847
rect 3280 1843 3284 1847
rect 3416 1843 3420 1847
rect 3536 1843 3540 1847
rect 168 1831 172 1835
rect 312 1831 316 1835
rect 496 1831 500 1835
rect 688 1831 692 1835
rect 872 1831 876 1835
rect 1048 1831 1052 1835
rect 1216 1831 1220 1835
rect 1376 1831 1380 1835
rect 1536 1831 1540 1835
rect 1704 1831 1708 1835
rect 2120 1815 2124 1819
rect 2168 1815 2172 1819
rect 2264 1815 2268 1819
rect 2424 1815 2428 1819
rect 2584 1815 2588 1819
rect 2744 1815 2748 1819
rect 2904 1815 2908 1819
rect 3056 1815 3060 1819
rect 3200 1815 3204 1819
rect 3344 1815 3348 1819
rect 3496 1815 3500 1819
rect 2168 1779 2172 1783
rect 1688 1767 1692 1771
rect 2728 1751 2732 1755
rect 2888 1751 2892 1755
rect 3480 1751 3484 1755
rect 328 1723 332 1727
rect 168 1683 172 1687
rect 248 1683 252 1687
rect 376 1683 380 1687
rect 528 1683 532 1687
rect 696 1683 700 1687
rect 872 1683 876 1687
rect 1040 1683 1044 1687
rect 1200 1683 1204 1687
rect 1352 1683 1356 1687
rect 1496 1683 1500 1687
rect 1640 1683 1644 1687
rect 1776 1683 1780 1687
rect 2136 1671 2140 1675
rect 2272 1671 2276 1675
rect 2416 1671 2420 1675
rect 2560 1671 2564 1675
rect 2696 1671 2700 1675
rect 2832 1671 2836 1675
rect 2960 1671 2964 1675
rect 3080 1671 3084 1675
rect 3192 1671 3196 1675
rect 3304 1671 3308 1675
rect 3424 1671 3428 1675
rect 3536 1671 3540 1675
rect 168 1667 172 1671
rect 320 1667 324 1671
rect 328 1667 332 1671
rect 504 1667 508 1671
rect 696 1667 700 1671
rect 880 1667 884 1671
rect 1056 1667 1060 1671
rect 1224 1667 1228 1671
rect 1384 1667 1388 1671
rect 1544 1667 1548 1671
rect 1704 1667 1708 1671
rect 1992 1655 1996 1659
rect 2112 1655 2116 1659
rect 2240 1655 2244 1659
rect 2376 1655 2380 1659
rect 2520 1655 2524 1659
rect 2664 1655 2668 1659
rect 2808 1655 2812 1659
rect 2888 1655 2892 1659
rect 2952 1655 2956 1659
rect 3096 1655 3100 1659
rect 3248 1655 3252 1659
rect 3400 1655 3404 1659
rect 3536 1655 3540 1659
rect 2888 1619 2892 1623
rect 2792 1591 2796 1595
rect 192 1527 196 1531
rect 320 1527 324 1531
rect 456 1527 460 1531
rect 600 1527 604 1531
rect 744 1527 748 1531
rect 880 1527 884 1531
rect 1016 1527 1020 1531
rect 1152 1527 1156 1531
rect 1280 1527 1284 1531
rect 1408 1527 1412 1531
rect 1544 1527 1548 1531
rect 256 1511 260 1515
rect 400 1511 404 1515
rect 544 1511 548 1515
rect 680 1511 684 1515
rect 808 1511 812 1515
rect 928 1511 932 1515
rect 1040 1511 1044 1515
rect 1144 1511 1148 1515
rect 1240 1511 1244 1515
rect 1344 1511 1348 1515
rect 1448 1511 1452 1515
rect 1928 1507 1932 1511
rect 2080 1507 2084 1511
rect 2240 1507 2244 1511
rect 2400 1507 2404 1511
rect 2560 1507 2564 1511
rect 2720 1507 2724 1511
rect 2872 1507 2876 1511
rect 3016 1507 3020 1511
rect 3152 1507 3156 1511
rect 3288 1507 3292 1511
rect 3424 1507 3428 1511
rect 3536 1507 3540 1511
rect 1928 1487 1932 1491
rect 2032 1487 2036 1491
rect 2160 1487 2164 1491
rect 2296 1487 2300 1491
rect 2440 1487 2444 1491
rect 2592 1487 2596 1491
rect 2744 1487 2748 1491
rect 2904 1487 2908 1491
rect 3064 1487 3068 1491
rect 3224 1487 3228 1491
rect 3392 1487 3396 1491
rect 3536 1487 3540 1491
rect 2280 1423 2284 1427
rect 2576 1423 2580 1427
rect 288 1363 292 1367
rect 384 1363 388 1367
rect 480 1363 484 1367
rect 576 1363 580 1367
rect 664 1363 668 1367
rect 752 1363 756 1367
rect 840 1363 844 1367
rect 952 1363 956 1367
rect 1080 1363 1084 1367
rect 1240 1363 1244 1367
rect 1416 1363 1420 1367
rect 1608 1363 1612 1367
rect 1776 1363 1780 1367
rect 384 1351 388 1355
rect 496 1351 500 1355
rect 616 1351 620 1355
rect 752 1351 756 1355
rect 888 1351 892 1355
rect 1032 1351 1036 1355
rect 1168 1351 1172 1355
rect 1304 1351 1308 1355
rect 1432 1351 1436 1355
rect 1552 1351 1556 1355
rect 1616 1351 1620 1355
rect 1672 1351 1676 1355
rect 1776 1351 1780 1355
rect 1928 1347 1932 1351
rect 2056 1347 2060 1351
rect 2200 1347 2204 1351
rect 2336 1347 2340 1351
rect 2464 1347 2468 1351
rect 2584 1347 2588 1351
rect 2704 1347 2708 1351
rect 2824 1347 2828 1351
rect 2944 1347 2948 1351
rect 1952 1327 1956 1331
rect 2072 1327 2076 1331
rect 2208 1327 2212 1331
rect 2344 1327 2348 1331
rect 2480 1327 2484 1331
rect 2616 1327 2620 1331
rect 2744 1327 2748 1331
rect 2864 1327 2868 1331
rect 2976 1327 2980 1331
rect 3088 1327 3092 1331
rect 3208 1327 3212 1331
rect 1616 1315 1620 1319
rect 736 1287 740 1291
rect 3192 1263 3196 1267
rect 344 1207 348 1211
rect 448 1207 452 1211
rect 568 1207 572 1211
rect 704 1207 708 1211
rect 848 1207 852 1211
rect 992 1207 996 1211
rect 1136 1207 1140 1211
rect 1272 1207 1276 1211
rect 1288 1207 1292 1211
rect 1408 1207 1412 1211
rect 1536 1207 1540 1211
rect 1664 1207 1668 1211
rect 1776 1207 1780 1211
rect 264 1195 268 1199
rect 440 1195 444 1199
rect 616 1195 620 1199
rect 784 1195 788 1199
rect 952 1195 956 1199
rect 1104 1195 1108 1199
rect 1248 1195 1252 1199
rect 1392 1195 1396 1199
rect 1528 1195 1532 1199
rect 1664 1195 1668 1199
rect 1776 1195 1780 1199
rect 1928 1179 1932 1183
rect 2104 1179 2108 1183
rect 2304 1179 2308 1183
rect 2504 1179 2508 1183
rect 2696 1179 2700 1183
rect 2880 1179 2884 1183
rect 3056 1179 3060 1183
rect 3224 1179 3228 1183
rect 3392 1179 3396 1183
rect 3536 1179 3540 1183
rect 1928 1163 1932 1167
rect 2008 1163 2012 1167
rect 2112 1163 2116 1167
rect 2240 1163 2244 1167
rect 2392 1163 2396 1167
rect 2552 1163 2556 1167
rect 2712 1163 2716 1167
rect 2864 1163 2868 1167
rect 3008 1163 3012 1167
rect 3088 1163 3092 1167
rect 3152 1163 3156 1167
rect 3288 1163 3292 1167
rect 3424 1163 3428 1167
rect 3536 1163 3540 1167
rect 600 1131 604 1135
rect 1288 1131 1292 1135
rect 1648 1131 1652 1135
rect 3088 1127 3092 1131
rect 2536 1099 2540 1103
rect 176 1051 180 1055
rect 312 1051 316 1055
rect 456 1051 460 1055
rect 600 1051 604 1055
rect 744 1051 748 1055
rect 880 1051 884 1055
rect 1008 1051 1012 1055
rect 1136 1051 1140 1055
rect 1256 1051 1260 1055
rect 1376 1051 1380 1055
rect 1504 1051 1508 1055
rect 168 1031 172 1035
rect 288 1031 292 1035
rect 432 1031 436 1035
rect 576 1031 580 1035
rect 712 1031 716 1035
rect 792 1031 796 1035
rect 832 1031 836 1035
rect 952 1031 956 1035
rect 1064 1031 1068 1035
rect 1168 1031 1172 1035
rect 1272 1031 1276 1035
rect 1384 1031 1388 1035
rect 2200 1015 2204 1019
rect 2288 1015 2292 1019
rect 2392 1015 2396 1019
rect 2512 1015 2516 1019
rect 2640 1015 2644 1019
rect 2784 1015 2788 1019
rect 2928 1015 2932 1019
rect 3080 1015 3084 1019
rect 3240 1015 3244 1019
rect 3400 1015 3404 1019
rect 3536 1015 3540 1019
rect 2328 1003 2332 1007
rect 2408 1003 2412 1007
rect 2496 1003 2500 1007
rect 2592 1003 2596 1007
rect 2632 1003 2636 1007
rect 2696 1003 2700 1007
rect 2808 1003 2812 1007
rect 2936 1003 2940 1007
rect 3080 1003 3084 1007
rect 3232 1003 3236 1007
rect 3392 1003 3396 1007
rect 3536 1003 3540 1007
rect 2632 967 2636 971
rect 2920 939 2924 943
rect 792 923 796 927
rect 168 883 172 887
rect 248 883 252 887
rect 360 883 364 887
rect 480 883 484 887
rect 600 883 604 887
rect 720 883 724 887
rect 832 883 836 887
rect 944 883 948 887
rect 1048 883 1052 887
rect 1152 883 1156 887
rect 1256 883 1260 887
rect 1360 883 1364 887
rect 168 863 172 867
rect 280 863 284 867
rect 424 863 428 867
rect 584 863 588 867
rect 744 863 748 867
rect 896 863 900 867
rect 1040 863 1044 867
rect 1176 863 1180 867
rect 1304 863 1308 867
rect 1424 863 1428 867
rect 1544 863 1548 867
rect 1672 863 1676 867
rect 2312 855 2316 859
rect 2392 855 2396 859
rect 2472 855 2476 859
rect 2552 855 2556 859
rect 2640 855 2644 859
rect 2736 855 2740 859
rect 2840 855 2844 859
rect 2944 855 2948 859
rect 3048 855 3052 859
rect 3144 855 3148 859
rect 3248 855 3252 859
rect 3352 855 3356 859
rect 3456 855 3460 859
rect 3536 855 3540 859
rect 2192 831 2196 835
rect 2272 831 2276 835
rect 2352 831 2356 835
rect 2448 831 2452 835
rect 2560 831 2564 835
rect 2680 831 2684 835
rect 2808 831 2812 835
rect 2936 831 2940 835
rect 3064 831 3068 835
rect 3184 831 3188 835
rect 3304 831 3308 835
rect 3432 831 3436 835
rect 3536 831 3540 835
rect 536 751 540 755
rect 168 711 172 715
rect 296 711 300 715
rect 464 711 468 715
rect 536 711 540 715
rect 640 711 644 715
rect 816 711 820 715
rect 984 711 988 715
rect 1136 711 1140 715
rect 1280 711 1284 715
rect 1416 711 1420 715
rect 1544 711 1548 715
rect 1672 711 1676 715
rect 1776 711 1780 715
rect 320 687 324 691
rect 432 687 436 691
rect 552 687 556 691
rect 680 687 684 691
rect 808 687 812 691
rect 928 687 932 691
rect 1048 687 1052 691
rect 1160 687 1164 691
rect 1272 687 1276 691
rect 1376 687 1380 691
rect 1480 687 1484 691
rect 1584 687 1588 691
rect 1688 687 1692 691
rect 1776 687 1780 691
rect 1928 683 1932 687
rect 2008 683 2012 687
rect 2104 683 2108 687
rect 2216 683 2220 687
rect 2344 683 2348 687
rect 2480 683 2484 687
rect 2624 683 2628 687
rect 2776 683 2780 687
rect 2928 683 2932 687
rect 3080 683 3084 687
rect 3232 683 3236 687
rect 3392 683 3396 687
rect 3536 683 3540 687
rect 1928 667 1932 671
rect 2120 667 2124 671
rect 2320 667 2324 671
rect 2504 667 2508 671
rect 2680 667 2684 671
rect 2856 667 2860 671
rect 3032 667 3036 671
rect 3208 667 3212 671
rect 3384 667 3388 671
rect 3536 667 3540 671
rect 344 543 348 547
rect 424 543 428 547
rect 504 543 508 547
rect 592 543 596 547
rect 680 543 684 547
rect 768 543 772 547
rect 856 543 860 547
rect 944 543 948 547
rect 1032 543 1036 547
rect 1120 543 1124 547
rect 1208 543 1212 547
rect 1296 543 1300 547
rect 1928 523 1932 527
rect 2008 523 2012 527
rect 2120 523 2124 527
rect 2248 523 2252 527
rect 2384 523 2388 527
rect 2528 523 2532 527
rect 2680 523 2684 527
rect 2840 523 2844 527
rect 3008 523 3012 527
rect 3184 523 3188 527
rect 3368 523 3372 527
rect 3536 523 3540 527
rect 264 519 268 523
rect 368 519 372 523
rect 464 519 468 523
rect 560 519 564 523
rect 656 519 660 523
rect 744 519 748 523
rect 832 519 836 523
rect 920 519 924 523
rect 1008 519 1012 523
rect 1096 519 1100 523
rect 1184 519 1188 523
rect 1272 519 1276 523
rect 2176 511 2180 515
rect 2256 511 2260 515
rect 2352 511 2356 515
rect 2456 511 2460 515
rect 2576 511 2580 515
rect 2712 511 2716 515
rect 2864 511 2868 515
rect 3024 511 3028 515
rect 3200 511 3204 515
rect 3376 511 3380 515
rect 3536 511 3540 515
rect 168 371 172 375
rect 280 371 284 375
rect 408 371 412 375
rect 528 371 532 375
rect 640 371 644 375
rect 752 371 756 375
rect 856 371 860 375
rect 952 371 956 375
rect 1040 371 1044 375
rect 1136 371 1140 375
rect 1232 371 1236 375
rect 1328 371 1332 375
rect 2368 367 2372 371
rect 2448 367 2452 371
rect 2528 367 2532 371
rect 2616 367 2620 371
rect 2720 367 2724 371
rect 2832 367 2836 371
rect 2960 367 2964 371
rect 3104 367 3108 371
rect 3248 367 3252 371
rect 3400 367 3404 371
rect 3536 367 3540 371
rect 168 347 172 351
rect 208 347 212 351
rect 272 347 276 351
rect 400 347 404 351
rect 536 347 540 351
rect 672 347 676 351
rect 800 347 804 351
rect 920 347 924 351
rect 1032 347 1036 351
rect 1144 347 1148 351
rect 1248 347 1252 351
rect 1352 347 1356 351
rect 1464 347 1468 351
rect 2104 347 2108 351
rect 2192 347 2196 351
rect 2288 347 2292 351
rect 2400 347 2404 351
rect 2528 347 2532 351
rect 2664 347 2668 351
rect 2800 347 2804 351
rect 2936 347 2940 351
rect 3064 347 3068 351
rect 3192 347 3196 351
rect 3312 347 3316 351
rect 3432 347 3436 351
rect 3536 347 3540 351
rect 208 311 212 315
rect 520 283 524 287
rect 256 199 260 203
rect 368 199 372 203
rect 496 199 500 203
rect 632 199 636 203
rect 768 199 772 203
rect 904 199 908 203
rect 1040 199 1044 203
rect 1168 199 1172 203
rect 1288 199 1292 203
rect 1400 199 1404 203
rect 1512 199 1516 203
rect 1632 199 1636 203
rect 1928 199 1932 203
rect 2016 199 2020 203
rect 2128 199 2132 203
rect 2256 199 2260 203
rect 2392 199 2396 203
rect 2536 199 2540 203
rect 2680 199 2684 203
rect 2824 199 2828 203
rect 2968 199 2972 203
rect 3112 199 3116 203
rect 3256 199 3260 203
rect 3408 199 3412 203
rect 3536 199 3540 203
rect 1928 175 1932 179
rect 2008 175 2012 179
rect 2112 175 2116 179
rect 2232 175 2236 179
rect 2360 175 2364 179
rect 2488 175 2492 179
rect 2608 175 2612 179
rect 2728 175 2732 179
rect 2840 175 2844 179
rect 2944 175 2948 179
rect 3040 175 3044 179
rect 3136 175 3140 179
rect 3232 175 3236 179
rect 3328 175 3332 179
rect 3424 175 3428 179
rect 184 155 188 159
rect 264 155 268 159
rect 344 155 348 159
rect 424 155 428 159
rect 504 155 508 159
rect 584 155 588 159
rect 672 155 676 159
rect 760 155 764 159
rect 848 155 852 159
rect 936 155 940 159
rect 1024 155 1028 159
rect 1112 155 1116 159
rect 1192 155 1196 159
rect 1272 155 1276 159
rect 1360 155 1364 159
rect 1448 155 1452 159
rect 1536 155 1540 159
rect 1616 155 1620 159
rect 1696 155 1700 159
rect 1776 155 1780 159
<< m2 >>
rect 2150 3648 2156 3649
rect 1870 3645 1876 3646
rect 1870 3641 1871 3645
rect 1875 3641 1876 3645
rect 2150 3644 2151 3648
rect 2155 3644 2156 3648
rect 2150 3643 2156 3644
rect 2438 3648 2444 3649
rect 2438 3644 2439 3648
rect 2443 3644 2444 3648
rect 2438 3643 2444 3644
rect 2726 3648 2732 3649
rect 2726 3644 2727 3648
rect 2731 3644 2732 3648
rect 2726 3643 2732 3644
rect 3014 3648 3020 3649
rect 3014 3644 3015 3648
rect 3019 3644 3020 3648
rect 3014 3643 3020 3644
rect 3590 3645 3596 3646
rect 1870 3640 1876 3641
rect 3590 3641 3591 3645
rect 3595 3641 3596 3645
rect 3590 3640 3596 3641
rect 2242 3639 2248 3640
rect 2242 3638 2243 3639
rect 2213 3636 2243 3638
rect 194 3635 200 3636
rect 194 3631 195 3635
rect 199 3634 200 3635
rect 263 3635 269 3636
rect 263 3634 264 3635
rect 199 3632 264 3634
rect 199 3631 200 3632
rect 194 3630 200 3631
rect 263 3631 264 3632
rect 268 3631 269 3635
rect 263 3630 269 3631
rect 290 3635 296 3636
rect 290 3631 291 3635
rect 295 3634 296 3635
rect 391 3635 397 3636
rect 391 3634 392 3635
rect 295 3632 392 3634
rect 295 3631 296 3632
rect 290 3630 296 3631
rect 391 3631 392 3632
rect 396 3631 397 3635
rect 391 3630 397 3631
rect 418 3635 424 3636
rect 418 3631 419 3635
rect 423 3634 424 3635
rect 527 3635 533 3636
rect 527 3634 528 3635
rect 423 3632 528 3634
rect 423 3631 424 3632
rect 418 3630 424 3631
rect 527 3631 528 3632
rect 532 3631 533 3635
rect 527 3630 533 3631
rect 554 3635 560 3636
rect 554 3631 555 3635
rect 559 3634 560 3635
rect 663 3635 669 3636
rect 663 3634 664 3635
rect 559 3632 664 3634
rect 559 3631 560 3632
rect 554 3630 560 3631
rect 663 3631 664 3632
rect 668 3631 669 3635
rect 663 3630 669 3631
rect 799 3635 808 3636
rect 799 3631 800 3635
rect 807 3631 808 3635
rect 799 3630 808 3631
rect 826 3635 832 3636
rect 826 3631 827 3635
rect 831 3634 832 3635
rect 935 3635 941 3636
rect 935 3634 936 3635
rect 831 3632 936 3634
rect 831 3631 832 3632
rect 826 3630 832 3631
rect 935 3631 936 3632
rect 940 3631 941 3635
rect 935 3630 941 3631
rect 962 3635 968 3636
rect 962 3631 963 3635
rect 967 3634 968 3635
rect 1079 3635 1085 3636
rect 1079 3634 1080 3635
rect 967 3632 1080 3634
rect 967 3631 968 3632
rect 962 3630 968 3631
rect 1079 3631 1080 3632
rect 1084 3631 1085 3635
rect 1079 3630 1085 3631
rect 1106 3635 1112 3636
rect 1106 3631 1107 3635
rect 1111 3634 1112 3635
rect 1223 3635 1229 3636
rect 1223 3634 1224 3635
rect 1111 3632 1224 3634
rect 1111 3631 1112 3632
rect 1106 3630 1112 3631
rect 1223 3631 1224 3632
rect 1228 3631 1229 3635
rect 2242 3635 2243 3636
rect 2247 3635 2248 3639
rect 2510 3639 2516 3640
rect 2510 3638 2511 3639
rect 2501 3636 2511 3638
rect 2242 3634 2248 3635
rect 2510 3635 2511 3636
rect 2515 3635 2516 3639
rect 3007 3639 3013 3640
rect 3007 3638 3008 3639
rect 2789 3636 3008 3638
rect 2510 3634 2516 3635
rect 3007 3635 3008 3636
rect 3012 3635 3013 3639
rect 3086 3639 3092 3640
rect 3086 3638 3087 3639
rect 3077 3636 3087 3638
rect 3007 3634 3013 3635
rect 3086 3635 3087 3636
rect 3091 3635 3092 3639
rect 3086 3634 3092 3635
rect 1223 3630 1229 3631
rect 1870 3628 1876 3629
rect 142 3626 148 3627
rect 142 3622 143 3626
rect 147 3622 148 3626
rect 142 3621 148 3622
rect 238 3626 244 3627
rect 238 3622 239 3626
rect 243 3622 244 3626
rect 238 3621 244 3622
rect 366 3626 372 3627
rect 366 3622 367 3626
rect 371 3622 372 3626
rect 366 3621 372 3622
rect 502 3626 508 3627
rect 502 3622 503 3626
rect 507 3622 508 3626
rect 502 3621 508 3622
rect 638 3626 644 3627
rect 638 3622 639 3626
rect 643 3622 644 3626
rect 638 3621 644 3622
rect 774 3626 780 3627
rect 774 3622 775 3626
rect 779 3622 780 3626
rect 774 3621 780 3622
rect 910 3626 916 3627
rect 910 3622 911 3626
rect 915 3622 916 3626
rect 910 3621 916 3622
rect 1054 3626 1060 3627
rect 1054 3622 1055 3626
rect 1059 3622 1060 3626
rect 1054 3621 1060 3622
rect 1198 3626 1204 3627
rect 1198 3622 1199 3626
rect 1203 3622 1204 3626
rect 1870 3624 1871 3628
rect 1875 3624 1876 3628
rect 1870 3623 1876 3624
rect 3590 3628 3596 3629
rect 3590 3624 3591 3628
rect 3595 3624 3596 3628
rect 3590 3623 3596 3624
rect 1198 3621 1204 3622
rect 2158 3610 2164 3611
rect 110 3608 116 3609
rect 110 3604 111 3608
rect 115 3604 116 3608
rect 110 3603 116 3604
rect 1830 3608 1836 3609
rect 1830 3604 1831 3608
rect 1835 3604 1836 3608
rect 2158 3606 2159 3610
rect 2163 3606 2164 3610
rect 2158 3605 2164 3606
rect 2446 3610 2452 3611
rect 2446 3606 2447 3610
rect 2451 3606 2452 3610
rect 2446 3605 2452 3606
rect 2734 3610 2740 3611
rect 2734 3606 2735 3610
rect 2739 3606 2740 3610
rect 2734 3605 2740 3606
rect 3022 3610 3028 3611
rect 3022 3606 3023 3610
rect 3027 3606 3028 3610
rect 3022 3605 3028 3606
rect 1830 3603 1836 3604
rect 194 3599 200 3600
rect 194 3595 195 3599
rect 199 3595 200 3599
rect 194 3594 200 3595
rect 290 3599 296 3600
rect 290 3595 291 3599
rect 295 3595 296 3599
rect 290 3594 296 3595
rect 418 3599 424 3600
rect 418 3595 419 3599
rect 423 3595 424 3599
rect 418 3594 424 3595
rect 554 3599 560 3600
rect 554 3595 555 3599
rect 559 3595 560 3599
rect 554 3594 560 3595
rect 826 3599 832 3600
rect 826 3595 827 3599
rect 831 3595 832 3599
rect 826 3594 832 3595
rect 962 3599 968 3600
rect 962 3595 963 3599
rect 967 3595 968 3599
rect 962 3594 968 3595
rect 1106 3599 1112 3600
rect 1106 3595 1107 3599
rect 1111 3595 1112 3599
rect 1106 3594 1112 3595
rect 2182 3599 2189 3600
rect 2182 3595 2183 3599
rect 2188 3595 2189 3599
rect 2182 3594 2189 3595
rect 2471 3599 2477 3600
rect 2471 3595 2472 3599
rect 2476 3598 2477 3599
rect 2502 3599 2508 3600
rect 2502 3598 2503 3599
rect 2476 3596 2503 3598
rect 2476 3595 2477 3596
rect 2471 3594 2477 3595
rect 2502 3595 2503 3596
rect 2507 3595 2508 3599
rect 2502 3594 2508 3595
rect 2510 3599 2516 3600
rect 2510 3595 2511 3599
rect 2515 3598 2516 3599
rect 2759 3599 2765 3600
rect 2759 3598 2760 3599
rect 2515 3596 2760 3598
rect 2515 3595 2516 3596
rect 2510 3594 2516 3595
rect 2759 3595 2760 3596
rect 2764 3595 2765 3599
rect 2759 3594 2765 3595
rect 3007 3599 3013 3600
rect 3007 3595 3008 3599
rect 3012 3598 3013 3599
rect 3047 3599 3053 3600
rect 3047 3598 3048 3599
rect 3012 3596 3048 3598
rect 3012 3595 3013 3596
rect 3007 3594 3013 3595
rect 3047 3595 3048 3596
rect 3052 3595 3053 3599
rect 3047 3594 3053 3595
rect 3270 3595 3276 3596
rect 3270 3594 3271 3595
rect 3080 3592 3271 3594
rect 110 3591 116 3592
rect 110 3587 111 3591
rect 115 3587 116 3591
rect 1830 3591 1836 3592
rect 110 3586 116 3587
rect 134 3588 140 3589
rect 134 3584 135 3588
rect 139 3584 140 3588
rect 134 3583 140 3584
rect 230 3588 236 3589
rect 230 3584 231 3588
rect 235 3584 236 3588
rect 230 3583 236 3584
rect 358 3588 364 3589
rect 358 3584 359 3588
rect 363 3584 364 3588
rect 358 3583 364 3584
rect 494 3588 500 3589
rect 494 3584 495 3588
rect 499 3584 500 3588
rect 494 3583 500 3584
rect 630 3588 636 3589
rect 630 3584 631 3588
rect 635 3584 636 3588
rect 630 3583 636 3584
rect 766 3588 772 3589
rect 766 3584 767 3588
rect 771 3584 772 3588
rect 766 3583 772 3584
rect 902 3588 908 3589
rect 902 3584 903 3588
rect 907 3584 908 3588
rect 902 3583 908 3584
rect 1046 3588 1052 3589
rect 1046 3584 1047 3588
rect 1051 3584 1052 3588
rect 1046 3583 1052 3584
rect 1190 3588 1196 3589
rect 1190 3584 1191 3588
rect 1195 3584 1196 3588
rect 1830 3587 1831 3591
rect 1835 3587 1836 3591
rect 1830 3586 1836 3587
rect 1927 3587 1936 3588
rect 1190 3583 1196 3584
rect 1927 3583 1928 3587
rect 1935 3583 1936 3587
rect 1927 3582 1936 3583
rect 1954 3587 1960 3588
rect 1954 3583 1955 3587
rect 1959 3586 1960 3587
rect 2007 3587 2013 3588
rect 2007 3586 2008 3587
rect 1959 3584 2008 3586
rect 1959 3583 1960 3584
rect 1954 3582 1960 3583
rect 2007 3583 2008 3584
rect 2012 3583 2013 3587
rect 2007 3582 2013 3583
rect 2034 3587 2040 3588
rect 2034 3583 2035 3587
rect 2039 3586 2040 3587
rect 2095 3587 2101 3588
rect 2095 3586 2096 3587
rect 2039 3584 2096 3586
rect 2039 3583 2040 3584
rect 2034 3582 2040 3583
rect 2095 3583 2096 3584
rect 2100 3583 2101 3587
rect 2095 3582 2101 3583
rect 2122 3587 2128 3588
rect 2122 3583 2123 3587
rect 2127 3586 2128 3587
rect 2199 3587 2205 3588
rect 2199 3586 2200 3587
rect 2127 3584 2200 3586
rect 2127 3583 2128 3584
rect 2122 3582 2128 3583
rect 2199 3583 2200 3584
rect 2204 3583 2205 3587
rect 2199 3582 2205 3583
rect 2242 3587 2248 3588
rect 2242 3583 2243 3587
rect 2247 3586 2248 3587
rect 2319 3587 2325 3588
rect 2319 3586 2320 3587
rect 2247 3584 2320 3586
rect 2247 3583 2248 3584
rect 2242 3582 2248 3583
rect 2319 3583 2320 3584
rect 2324 3583 2325 3587
rect 2319 3582 2325 3583
rect 2346 3587 2352 3588
rect 2346 3583 2347 3587
rect 2351 3586 2352 3587
rect 2447 3587 2453 3588
rect 2447 3586 2448 3587
rect 2351 3584 2448 3586
rect 2351 3583 2352 3584
rect 2346 3582 2352 3583
rect 2447 3583 2448 3584
rect 2452 3583 2453 3587
rect 2447 3582 2453 3583
rect 2474 3587 2480 3588
rect 2474 3583 2475 3587
rect 2479 3586 2480 3587
rect 2583 3587 2589 3588
rect 2583 3586 2584 3587
rect 2479 3584 2584 3586
rect 2479 3583 2480 3584
rect 2474 3582 2480 3583
rect 2583 3583 2584 3584
rect 2588 3583 2589 3587
rect 2583 3582 2589 3583
rect 2719 3587 2725 3588
rect 2719 3583 2720 3587
rect 2724 3586 2725 3587
rect 2746 3587 2752 3588
rect 2724 3584 2734 3586
rect 2724 3583 2725 3584
rect 2719 3582 2725 3583
rect 2730 3583 2736 3584
rect 2730 3579 2731 3583
rect 2735 3579 2736 3583
rect 2746 3583 2747 3587
rect 2751 3586 2752 3587
rect 2855 3587 2861 3588
rect 2855 3586 2856 3587
rect 2751 3584 2856 3586
rect 2751 3583 2752 3584
rect 2746 3582 2752 3583
rect 2855 3583 2856 3584
rect 2860 3583 2861 3587
rect 2855 3582 2861 3583
rect 2999 3587 3005 3588
rect 2999 3583 3000 3587
rect 3004 3586 3005 3587
rect 3080 3586 3082 3592
rect 3270 3591 3271 3592
rect 3275 3591 3276 3595
rect 3270 3590 3276 3591
rect 3004 3584 3082 3586
rect 3086 3587 3092 3588
rect 3004 3583 3005 3584
rect 2999 3582 3005 3583
rect 3086 3583 3087 3587
rect 3091 3586 3092 3587
rect 3143 3587 3149 3588
rect 3143 3586 3144 3587
rect 3091 3584 3144 3586
rect 3091 3583 3092 3584
rect 3086 3582 3092 3583
rect 3143 3583 3144 3584
rect 3148 3583 3149 3587
rect 3143 3582 3149 3583
rect 3170 3587 3176 3588
rect 3170 3583 3171 3587
rect 3175 3586 3176 3587
rect 3287 3587 3293 3588
rect 3287 3586 3288 3587
rect 3175 3584 3288 3586
rect 3175 3583 3176 3584
rect 3170 3582 3176 3583
rect 3287 3583 3288 3584
rect 3292 3583 3293 3587
rect 3287 3582 3293 3583
rect 1902 3578 1908 3579
rect 1902 3574 1903 3578
rect 1907 3574 1908 3578
rect 1902 3573 1908 3574
rect 1982 3578 1988 3579
rect 1982 3574 1983 3578
rect 1987 3574 1988 3578
rect 1982 3573 1988 3574
rect 2070 3578 2076 3579
rect 2070 3574 2071 3578
rect 2075 3574 2076 3578
rect 2070 3573 2076 3574
rect 2174 3578 2180 3579
rect 2174 3574 2175 3578
rect 2179 3574 2180 3578
rect 2174 3573 2180 3574
rect 2294 3578 2300 3579
rect 2294 3574 2295 3578
rect 2299 3574 2300 3578
rect 2294 3573 2300 3574
rect 2422 3578 2428 3579
rect 2422 3574 2423 3578
rect 2427 3574 2428 3578
rect 2422 3573 2428 3574
rect 2558 3578 2564 3579
rect 2558 3574 2559 3578
rect 2563 3574 2564 3578
rect 2558 3573 2564 3574
rect 2694 3578 2700 3579
rect 2730 3578 2736 3579
rect 2830 3578 2836 3579
rect 2694 3574 2695 3578
rect 2699 3574 2700 3578
rect 2694 3573 2700 3574
rect 2830 3574 2831 3578
rect 2835 3574 2836 3578
rect 2830 3573 2836 3574
rect 2974 3578 2980 3579
rect 2974 3574 2975 3578
rect 2979 3574 2980 3578
rect 2974 3573 2980 3574
rect 3118 3578 3124 3579
rect 3118 3574 3119 3578
rect 3123 3574 3124 3578
rect 3118 3573 3124 3574
rect 3262 3578 3268 3579
rect 3262 3574 3263 3578
rect 3267 3574 3268 3578
rect 3262 3573 3268 3574
rect 450 3571 456 3572
rect 450 3567 451 3571
rect 455 3570 456 3571
rect 647 3571 653 3572
rect 647 3570 648 3571
rect 455 3568 648 3570
rect 455 3567 456 3568
rect 450 3566 456 3567
rect 647 3567 648 3568
rect 652 3567 653 3571
rect 647 3566 653 3567
rect 802 3571 808 3572
rect 802 3567 803 3571
rect 807 3570 808 3571
rect 910 3571 916 3572
rect 910 3570 911 3571
rect 807 3568 911 3570
rect 807 3567 808 3568
rect 802 3566 808 3567
rect 910 3567 911 3568
rect 915 3567 916 3571
rect 910 3566 916 3567
rect 1054 3571 1060 3572
rect 1054 3567 1055 3571
rect 1059 3570 1060 3571
rect 1207 3571 1213 3572
rect 1207 3570 1208 3571
rect 1059 3568 1208 3570
rect 1059 3567 1060 3568
rect 1054 3566 1060 3567
rect 1207 3567 1208 3568
rect 1212 3567 1213 3571
rect 1207 3566 1213 3567
rect 1870 3560 1876 3561
rect 1870 3556 1871 3560
rect 1875 3556 1876 3560
rect 1870 3555 1876 3556
rect 3590 3560 3596 3561
rect 3590 3556 3591 3560
rect 3595 3556 3596 3560
rect 3590 3555 3596 3556
rect 1954 3551 1960 3552
rect 1954 3547 1955 3551
rect 1959 3547 1960 3551
rect 1954 3546 1960 3547
rect 2034 3551 2040 3552
rect 2034 3547 2035 3551
rect 2039 3547 2040 3551
rect 2034 3546 2040 3547
rect 2122 3551 2128 3552
rect 2122 3547 2123 3551
rect 2127 3547 2128 3551
rect 2122 3546 2128 3547
rect 2182 3551 2188 3552
rect 2182 3547 2183 3551
rect 2187 3547 2188 3551
rect 2182 3546 2188 3547
rect 2346 3551 2352 3552
rect 2346 3547 2347 3551
rect 2351 3547 2352 3551
rect 2346 3546 2352 3547
rect 2474 3551 2480 3552
rect 2474 3547 2475 3551
rect 2479 3547 2480 3551
rect 2474 3546 2480 3547
rect 2746 3551 2752 3552
rect 2746 3547 2747 3551
rect 2751 3547 2752 3551
rect 2746 3546 2752 3547
rect 2838 3551 2844 3552
rect 2838 3547 2839 3551
rect 2843 3547 2844 3551
rect 2838 3546 2844 3547
rect 3170 3551 3176 3552
rect 3170 3547 3171 3551
rect 3175 3547 3176 3551
rect 3170 3546 3176 3547
rect 3270 3551 3276 3552
rect 3270 3547 3271 3551
rect 3275 3547 3276 3551
rect 3270 3546 3276 3547
rect 182 3544 188 3545
rect 110 3541 116 3542
rect 110 3537 111 3541
rect 115 3537 116 3541
rect 182 3540 183 3544
rect 187 3540 188 3544
rect 182 3539 188 3540
rect 302 3544 308 3545
rect 302 3540 303 3544
rect 307 3540 308 3544
rect 302 3539 308 3540
rect 414 3544 420 3545
rect 414 3540 415 3544
rect 419 3540 420 3544
rect 414 3539 420 3540
rect 526 3544 532 3545
rect 526 3540 527 3544
rect 531 3540 532 3544
rect 526 3539 532 3540
rect 630 3544 636 3545
rect 630 3540 631 3544
rect 635 3540 636 3544
rect 630 3539 636 3540
rect 734 3544 740 3545
rect 734 3540 735 3544
rect 739 3540 740 3544
rect 734 3539 740 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 918 3544 924 3545
rect 918 3540 919 3544
rect 923 3540 924 3544
rect 918 3539 924 3540
rect 1006 3544 1012 3545
rect 1006 3540 1007 3544
rect 1011 3540 1012 3544
rect 1006 3539 1012 3540
rect 1094 3544 1100 3545
rect 1094 3540 1095 3544
rect 1099 3540 1100 3544
rect 1094 3539 1100 3540
rect 1182 3544 1188 3545
rect 1182 3540 1183 3544
rect 1187 3540 1188 3544
rect 1182 3539 1188 3540
rect 1270 3544 1276 3545
rect 1270 3540 1271 3544
rect 1275 3540 1276 3544
rect 1270 3539 1276 3540
rect 1358 3544 1364 3545
rect 1358 3540 1359 3544
rect 1363 3540 1364 3544
rect 1358 3539 1364 3540
rect 1446 3544 1452 3545
rect 1446 3540 1447 3544
rect 1451 3540 1452 3544
rect 1870 3543 1876 3544
rect 1446 3539 1452 3540
rect 1830 3541 1836 3542
rect 110 3536 116 3537
rect 1830 3537 1831 3541
rect 1835 3537 1836 3541
rect 1870 3539 1871 3543
rect 1875 3539 1876 3543
rect 3590 3543 3596 3544
rect 1870 3538 1876 3539
rect 1894 3540 1900 3541
rect 1830 3536 1836 3537
rect 1894 3536 1895 3540
rect 1899 3536 1900 3540
rect 258 3535 264 3536
rect 258 3534 259 3535
rect 245 3532 259 3534
rect 258 3531 259 3532
rect 263 3531 264 3535
rect 382 3535 388 3536
rect 382 3534 383 3535
rect 365 3532 383 3534
rect 258 3530 264 3531
rect 382 3531 383 3532
rect 387 3531 388 3535
rect 602 3535 608 3536
rect 602 3534 603 3535
rect 382 3530 388 3531
rect 242 3527 248 3528
rect 110 3524 116 3525
rect 110 3520 111 3524
rect 115 3520 116 3524
rect 242 3523 243 3527
rect 247 3526 248 3527
rect 432 3526 434 3533
rect 589 3532 603 3534
rect 602 3531 603 3532
rect 607 3531 608 3535
rect 706 3535 712 3536
rect 706 3534 707 3535
rect 693 3532 707 3534
rect 602 3530 608 3531
rect 706 3531 707 3532
rect 711 3531 712 3535
rect 806 3535 812 3536
rect 806 3534 807 3535
rect 797 3532 807 3534
rect 706 3530 712 3531
rect 806 3531 807 3532
rect 811 3531 812 3535
rect 898 3535 904 3536
rect 898 3534 899 3535
rect 893 3532 899 3534
rect 806 3530 812 3531
rect 898 3531 899 3532
rect 903 3531 904 3535
rect 898 3530 904 3531
rect 910 3535 916 3536
rect 910 3531 911 3535
rect 915 3534 916 3535
rect 1074 3535 1080 3536
rect 1074 3534 1075 3535
rect 915 3532 937 3534
rect 1069 3532 1075 3534
rect 915 3531 916 3532
rect 910 3530 916 3531
rect 1074 3531 1075 3532
rect 1079 3531 1080 3535
rect 1175 3535 1181 3536
rect 1175 3534 1176 3535
rect 1157 3532 1176 3534
rect 1074 3530 1080 3531
rect 1175 3531 1176 3532
rect 1180 3531 1181 3535
rect 1250 3535 1256 3536
rect 1250 3534 1251 3535
rect 1245 3532 1251 3534
rect 1175 3530 1181 3531
rect 1250 3531 1251 3532
rect 1255 3531 1256 3535
rect 1338 3535 1344 3536
rect 1338 3534 1339 3535
rect 1333 3532 1339 3534
rect 1250 3530 1256 3531
rect 1338 3531 1339 3532
rect 1343 3531 1344 3535
rect 1426 3535 1432 3536
rect 1426 3534 1427 3535
rect 1421 3532 1427 3534
rect 1338 3530 1344 3531
rect 1426 3531 1427 3532
rect 1431 3531 1432 3535
rect 1426 3530 1432 3531
rect 1434 3535 1440 3536
rect 1894 3535 1900 3536
rect 1974 3540 1980 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 2062 3540 2068 3541
rect 2062 3536 2063 3540
rect 2067 3536 2068 3540
rect 2062 3535 2068 3536
rect 2166 3540 2172 3541
rect 2166 3536 2167 3540
rect 2171 3536 2172 3540
rect 2166 3535 2172 3536
rect 2286 3540 2292 3541
rect 2286 3536 2287 3540
rect 2291 3536 2292 3540
rect 2286 3535 2292 3536
rect 2414 3540 2420 3541
rect 2414 3536 2415 3540
rect 2419 3536 2420 3540
rect 2414 3535 2420 3536
rect 2550 3540 2556 3541
rect 2550 3536 2551 3540
rect 2555 3536 2556 3540
rect 2550 3535 2556 3536
rect 2686 3540 2692 3541
rect 2686 3536 2687 3540
rect 2691 3536 2692 3540
rect 2686 3535 2692 3536
rect 2822 3540 2828 3541
rect 2822 3536 2823 3540
rect 2827 3536 2828 3540
rect 2822 3535 2828 3536
rect 2966 3540 2972 3541
rect 2966 3536 2967 3540
rect 2971 3536 2972 3540
rect 2966 3535 2972 3536
rect 3110 3540 3116 3541
rect 3110 3536 3111 3540
rect 3115 3536 3116 3540
rect 3110 3535 3116 3536
rect 3254 3540 3260 3541
rect 3254 3536 3255 3540
rect 3259 3536 3260 3540
rect 3590 3539 3591 3543
rect 3595 3539 3596 3543
rect 3590 3538 3596 3539
rect 3254 3535 3260 3536
rect 1434 3531 1435 3535
rect 1439 3534 1440 3535
rect 1439 3532 1465 3534
rect 1439 3531 1440 3532
rect 1434 3530 1440 3531
rect 247 3524 434 3526
rect 1830 3524 1836 3525
rect 247 3523 248 3524
rect 242 3522 248 3523
rect 110 3519 116 3520
rect 1830 3520 1831 3524
rect 1835 3520 1836 3524
rect 1830 3519 1836 3520
rect 2558 3523 2564 3524
rect 2558 3519 2559 3523
rect 2563 3522 2564 3523
rect 2567 3523 2573 3524
rect 2567 3522 2568 3523
rect 2563 3520 2568 3522
rect 2563 3519 2564 3520
rect 2558 3518 2564 3519
rect 2567 3519 2568 3520
rect 2572 3519 2573 3523
rect 2567 3518 2573 3519
rect 2983 3523 2992 3524
rect 2983 3519 2984 3523
rect 2991 3519 2992 3523
rect 2983 3518 2992 3519
rect 190 3506 196 3507
rect 190 3502 191 3506
rect 195 3502 196 3506
rect 190 3501 196 3502
rect 310 3506 316 3507
rect 310 3502 311 3506
rect 315 3502 316 3506
rect 310 3501 316 3502
rect 422 3506 428 3507
rect 422 3502 423 3506
rect 427 3502 428 3506
rect 422 3501 428 3502
rect 534 3506 540 3507
rect 534 3502 535 3506
rect 539 3502 540 3506
rect 534 3501 540 3502
rect 638 3506 644 3507
rect 638 3502 639 3506
rect 643 3502 644 3506
rect 638 3501 644 3502
rect 742 3506 748 3507
rect 742 3502 743 3506
rect 747 3502 748 3506
rect 742 3501 748 3502
rect 838 3506 844 3507
rect 838 3502 839 3506
rect 843 3502 844 3506
rect 838 3501 844 3502
rect 926 3506 932 3507
rect 926 3502 927 3506
rect 931 3502 932 3506
rect 926 3501 932 3502
rect 1014 3506 1020 3507
rect 1014 3502 1015 3506
rect 1019 3502 1020 3506
rect 1014 3501 1020 3502
rect 1102 3506 1108 3507
rect 1102 3502 1103 3506
rect 1107 3502 1108 3506
rect 1102 3501 1108 3502
rect 1190 3506 1196 3507
rect 1190 3502 1191 3506
rect 1195 3502 1196 3506
rect 1190 3501 1196 3502
rect 1278 3506 1284 3507
rect 1278 3502 1279 3506
rect 1283 3502 1284 3506
rect 1278 3501 1284 3502
rect 1366 3506 1372 3507
rect 1366 3502 1367 3506
rect 1371 3502 1372 3506
rect 1366 3501 1372 3502
rect 1454 3506 1460 3507
rect 1454 3502 1455 3506
rect 1459 3502 1460 3506
rect 1454 3501 1460 3502
rect 1966 3496 1972 3497
rect 215 3495 221 3496
rect 215 3491 216 3495
rect 220 3494 221 3495
rect 242 3495 248 3496
rect 242 3494 243 3495
rect 220 3492 243 3494
rect 220 3491 221 3492
rect 215 3490 221 3491
rect 242 3491 243 3492
rect 247 3491 248 3495
rect 242 3490 248 3491
rect 258 3495 264 3496
rect 258 3491 259 3495
rect 263 3494 264 3495
rect 335 3495 341 3496
rect 335 3494 336 3495
rect 263 3492 336 3494
rect 263 3491 264 3492
rect 258 3490 264 3491
rect 335 3491 336 3492
rect 340 3491 341 3495
rect 335 3490 341 3491
rect 447 3495 456 3496
rect 447 3491 448 3495
rect 455 3491 456 3495
rect 447 3490 456 3491
rect 559 3495 565 3496
rect 559 3491 560 3495
rect 564 3494 565 3495
rect 602 3495 608 3496
rect 564 3492 598 3494
rect 564 3491 565 3492
rect 559 3490 565 3491
rect 596 3486 598 3492
rect 602 3491 603 3495
rect 607 3494 608 3495
rect 663 3495 669 3496
rect 663 3494 664 3495
rect 607 3492 664 3494
rect 607 3491 608 3492
rect 602 3490 608 3491
rect 663 3491 664 3492
rect 668 3491 669 3495
rect 663 3490 669 3491
rect 706 3495 712 3496
rect 706 3491 707 3495
rect 711 3494 712 3495
rect 767 3495 773 3496
rect 767 3494 768 3495
rect 711 3492 768 3494
rect 711 3491 712 3492
rect 706 3490 712 3491
rect 767 3491 768 3492
rect 772 3491 773 3495
rect 767 3490 773 3491
rect 806 3495 812 3496
rect 806 3491 807 3495
rect 811 3494 812 3495
rect 863 3495 869 3496
rect 863 3494 864 3495
rect 811 3492 864 3494
rect 811 3491 812 3492
rect 806 3490 812 3491
rect 863 3491 864 3492
rect 868 3491 869 3495
rect 863 3490 869 3491
rect 898 3495 904 3496
rect 898 3491 899 3495
rect 903 3494 904 3495
rect 951 3495 957 3496
rect 951 3494 952 3495
rect 903 3492 952 3494
rect 903 3491 904 3492
rect 898 3490 904 3491
rect 951 3491 952 3492
rect 956 3491 957 3495
rect 951 3490 957 3491
rect 1039 3495 1045 3496
rect 1039 3491 1040 3495
rect 1044 3494 1045 3495
rect 1054 3495 1060 3496
rect 1054 3494 1055 3495
rect 1044 3492 1055 3494
rect 1044 3491 1045 3492
rect 1039 3490 1045 3491
rect 1054 3491 1055 3492
rect 1059 3491 1060 3495
rect 1054 3490 1060 3491
rect 1074 3495 1080 3496
rect 1074 3491 1075 3495
rect 1079 3494 1080 3495
rect 1127 3495 1133 3496
rect 1127 3494 1128 3495
rect 1079 3492 1128 3494
rect 1079 3491 1080 3492
rect 1074 3490 1080 3491
rect 1127 3491 1128 3492
rect 1132 3491 1133 3495
rect 1127 3490 1133 3491
rect 1175 3495 1181 3496
rect 1175 3491 1176 3495
rect 1180 3494 1181 3495
rect 1215 3495 1221 3496
rect 1215 3494 1216 3495
rect 1180 3492 1216 3494
rect 1180 3491 1181 3492
rect 1175 3490 1181 3491
rect 1215 3491 1216 3492
rect 1220 3491 1221 3495
rect 1215 3490 1221 3491
rect 1250 3495 1256 3496
rect 1250 3491 1251 3495
rect 1255 3494 1256 3495
rect 1303 3495 1309 3496
rect 1303 3494 1304 3495
rect 1255 3492 1304 3494
rect 1255 3491 1256 3492
rect 1250 3490 1256 3491
rect 1303 3491 1304 3492
rect 1308 3491 1309 3495
rect 1303 3490 1309 3491
rect 1338 3495 1344 3496
rect 1338 3491 1339 3495
rect 1343 3494 1344 3495
rect 1391 3495 1397 3496
rect 1391 3494 1392 3495
rect 1343 3492 1392 3494
rect 1343 3491 1344 3492
rect 1338 3490 1344 3491
rect 1391 3491 1392 3492
rect 1396 3491 1397 3495
rect 1391 3490 1397 3491
rect 1426 3495 1432 3496
rect 1426 3491 1427 3495
rect 1431 3494 1432 3495
rect 1479 3495 1485 3496
rect 1479 3494 1480 3495
rect 1431 3492 1480 3494
rect 1431 3491 1432 3492
rect 1426 3490 1432 3491
rect 1479 3491 1480 3492
rect 1484 3491 1485 3495
rect 1479 3490 1485 3491
rect 1870 3493 1876 3494
rect 1870 3489 1871 3493
rect 1875 3489 1876 3493
rect 1966 3492 1967 3496
rect 1971 3492 1972 3496
rect 1966 3491 1972 3492
rect 2150 3496 2156 3497
rect 2150 3492 2151 3496
rect 2155 3492 2156 3496
rect 2150 3491 2156 3492
rect 2334 3496 2340 3497
rect 2334 3492 2335 3496
rect 2339 3492 2340 3496
rect 2334 3491 2340 3492
rect 2510 3496 2516 3497
rect 2510 3492 2511 3496
rect 2515 3492 2516 3496
rect 2510 3491 2516 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2822 3496 2828 3497
rect 2822 3492 2823 3496
rect 2827 3492 2828 3496
rect 2822 3491 2828 3492
rect 2958 3496 2964 3497
rect 2958 3492 2959 3496
rect 2963 3492 2964 3496
rect 2958 3491 2964 3492
rect 3078 3496 3084 3497
rect 3078 3492 3079 3496
rect 3083 3492 3084 3496
rect 3078 3491 3084 3492
rect 3190 3496 3196 3497
rect 3190 3492 3191 3496
rect 3195 3492 3196 3496
rect 3190 3491 3196 3492
rect 3302 3496 3308 3497
rect 3302 3492 3303 3496
rect 3307 3492 3308 3496
rect 3302 3491 3308 3492
rect 3414 3496 3420 3497
rect 3414 3492 3415 3496
rect 3419 3492 3420 3496
rect 3414 3491 3420 3492
rect 3502 3496 3508 3497
rect 3502 3492 3503 3496
rect 3507 3492 3508 3496
rect 3502 3491 3508 3492
rect 3590 3493 3596 3494
rect 1870 3488 1876 3489
rect 3590 3489 3591 3493
rect 3595 3489 3596 3493
rect 3590 3488 3596 3489
rect 846 3487 852 3488
rect 846 3486 847 3487
rect 596 3484 847 3486
rect 846 3483 847 3484
rect 851 3483 852 3487
rect 846 3482 852 3483
rect 1930 3487 1936 3488
rect 1930 3483 1931 3487
rect 1935 3486 1936 3487
rect 2034 3487 2040 3488
rect 1935 3484 1985 3486
rect 1935 3483 1936 3484
rect 1930 3482 1936 3483
rect 2034 3483 2035 3487
rect 2039 3486 2040 3487
rect 2402 3487 2408 3488
rect 2039 3484 2169 3486
rect 2039 3483 2040 3484
rect 2034 3482 2040 3483
rect 2396 3478 2398 3485
rect 2402 3483 2403 3487
rect 2407 3486 2408 3487
rect 2738 3487 2744 3488
rect 2407 3484 2529 3486
rect 2407 3483 2408 3484
rect 2402 3482 2408 3483
rect 2732 3480 2734 3485
rect 2738 3483 2739 3487
rect 2743 3486 2744 3487
rect 3042 3487 3048 3488
rect 3042 3486 3043 3487
rect 2743 3484 2841 3486
rect 3021 3484 3043 3486
rect 2743 3483 2744 3484
rect 2738 3482 2744 3483
rect 3042 3483 3043 3484
rect 3047 3483 3048 3487
rect 3158 3487 3164 3488
rect 3158 3486 3159 3487
rect 3141 3484 3159 3486
rect 3042 3482 3048 3483
rect 3158 3483 3159 3484
rect 3163 3483 3164 3487
rect 3270 3487 3276 3488
rect 3270 3486 3271 3487
rect 3253 3484 3271 3486
rect 3158 3482 3164 3483
rect 3270 3483 3271 3484
rect 3275 3483 3276 3487
rect 3382 3487 3388 3488
rect 3382 3486 3383 3487
rect 3365 3484 3383 3486
rect 3270 3482 3276 3483
rect 3382 3483 3383 3484
rect 3387 3483 3388 3487
rect 3482 3487 3488 3488
rect 3482 3486 3483 3487
rect 3477 3484 3483 3486
rect 3382 3482 3388 3483
rect 3482 3483 3483 3484
rect 3487 3483 3488 3487
rect 3482 3482 3488 3483
rect 3564 3480 3566 3485
rect 2407 3479 2413 3480
rect 2407 3478 2408 3479
rect 1870 3476 1876 3477
rect 2396 3476 2408 3478
rect 255 3475 261 3476
rect 255 3471 256 3475
rect 260 3474 261 3475
rect 374 3475 380 3476
rect 374 3474 375 3475
rect 260 3472 375 3474
rect 260 3471 261 3472
rect 255 3470 261 3471
rect 374 3471 375 3472
rect 379 3471 380 3475
rect 374 3470 380 3471
rect 382 3475 388 3476
rect 382 3471 383 3475
rect 387 3474 388 3475
rect 391 3475 397 3476
rect 391 3474 392 3475
rect 387 3472 392 3474
rect 387 3471 388 3472
rect 382 3470 388 3471
rect 391 3471 392 3472
rect 396 3471 397 3475
rect 391 3470 397 3471
rect 518 3475 524 3476
rect 518 3471 519 3475
rect 523 3474 524 3475
rect 527 3475 533 3476
rect 527 3474 528 3475
rect 523 3472 528 3474
rect 523 3471 524 3472
rect 518 3470 524 3471
rect 527 3471 528 3472
rect 532 3471 533 3475
rect 527 3470 533 3471
rect 554 3475 560 3476
rect 554 3471 555 3475
rect 559 3474 560 3475
rect 647 3475 653 3476
rect 647 3474 648 3475
rect 559 3472 648 3474
rect 559 3471 560 3472
rect 554 3470 560 3471
rect 647 3471 648 3472
rect 652 3471 653 3475
rect 647 3470 653 3471
rect 674 3475 680 3476
rect 674 3471 675 3475
rect 679 3474 680 3475
rect 759 3475 765 3476
rect 759 3474 760 3475
rect 679 3472 760 3474
rect 679 3471 680 3472
rect 674 3470 680 3471
rect 759 3471 760 3472
rect 764 3471 765 3475
rect 759 3470 765 3471
rect 786 3475 792 3476
rect 786 3471 787 3475
rect 791 3474 792 3475
rect 863 3475 869 3476
rect 863 3474 864 3475
rect 791 3472 864 3474
rect 791 3471 792 3472
rect 786 3470 792 3471
rect 863 3471 864 3472
rect 868 3471 869 3475
rect 863 3470 869 3471
rect 967 3475 973 3476
rect 967 3471 968 3475
rect 972 3474 973 3475
rect 986 3475 992 3476
rect 986 3474 987 3475
rect 972 3472 987 3474
rect 972 3471 973 3472
rect 967 3470 973 3471
rect 986 3471 987 3472
rect 991 3471 992 3475
rect 986 3470 992 3471
rect 994 3475 1000 3476
rect 994 3471 995 3475
rect 999 3474 1000 3475
rect 1063 3475 1069 3476
rect 1063 3474 1064 3475
rect 999 3472 1064 3474
rect 999 3471 1000 3472
rect 994 3470 1000 3471
rect 1063 3471 1064 3472
rect 1068 3471 1069 3475
rect 1063 3470 1069 3471
rect 1090 3475 1096 3476
rect 1090 3471 1091 3475
rect 1095 3474 1096 3475
rect 1159 3475 1165 3476
rect 1159 3474 1160 3475
rect 1095 3472 1160 3474
rect 1095 3471 1096 3472
rect 1090 3470 1096 3471
rect 1159 3471 1160 3472
rect 1164 3471 1165 3475
rect 1159 3470 1165 3471
rect 1206 3475 1212 3476
rect 1206 3471 1207 3475
rect 1211 3474 1212 3475
rect 1255 3475 1261 3476
rect 1255 3474 1256 3475
rect 1211 3472 1256 3474
rect 1211 3471 1212 3472
rect 1206 3470 1212 3471
rect 1255 3471 1256 3472
rect 1260 3471 1261 3475
rect 1255 3470 1261 3471
rect 1303 3475 1309 3476
rect 1303 3471 1304 3475
rect 1308 3474 1309 3475
rect 1351 3475 1357 3476
rect 1351 3474 1352 3475
rect 1308 3472 1352 3474
rect 1308 3471 1309 3472
rect 1303 3470 1309 3471
rect 1351 3471 1352 3472
rect 1356 3471 1357 3475
rect 1870 3472 1871 3476
rect 1875 3472 1876 3476
rect 2407 3475 2408 3476
rect 2412 3475 2413 3479
rect 2407 3474 2413 3475
rect 2730 3479 2736 3480
rect 2730 3475 2731 3479
rect 2735 3475 2736 3479
rect 2730 3474 2736 3475
rect 3562 3479 3568 3480
rect 3562 3475 3563 3479
rect 3567 3475 3568 3479
rect 3562 3474 3568 3475
rect 3590 3476 3596 3477
rect 1870 3471 1876 3472
rect 3590 3472 3591 3476
rect 3595 3472 3596 3476
rect 3590 3471 3596 3472
rect 1351 3470 1357 3471
rect 230 3466 236 3467
rect 230 3462 231 3466
rect 235 3462 236 3466
rect 230 3461 236 3462
rect 366 3466 372 3467
rect 366 3462 367 3466
rect 371 3462 372 3466
rect 366 3461 372 3462
rect 502 3466 508 3467
rect 502 3462 503 3466
rect 507 3462 508 3466
rect 502 3461 508 3462
rect 622 3466 628 3467
rect 622 3462 623 3466
rect 627 3462 628 3466
rect 622 3461 628 3462
rect 734 3466 740 3467
rect 734 3462 735 3466
rect 739 3462 740 3466
rect 734 3461 740 3462
rect 838 3466 844 3467
rect 838 3462 839 3466
rect 843 3462 844 3466
rect 838 3461 844 3462
rect 942 3466 948 3467
rect 942 3462 943 3466
rect 947 3462 948 3466
rect 942 3461 948 3462
rect 1038 3466 1044 3467
rect 1038 3462 1039 3466
rect 1043 3462 1044 3466
rect 1038 3461 1044 3462
rect 1134 3466 1140 3467
rect 1134 3462 1135 3466
rect 1139 3462 1140 3466
rect 1134 3461 1140 3462
rect 1230 3466 1236 3467
rect 1230 3462 1231 3466
rect 1235 3462 1236 3466
rect 1230 3461 1236 3462
rect 1326 3466 1332 3467
rect 1326 3462 1327 3466
rect 1331 3462 1332 3466
rect 1326 3461 1332 3462
rect 1974 3458 1980 3459
rect 1974 3454 1975 3458
rect 1979 3454 1980 3458
rect 1974 3453 1980 3454
rect 2158 3458 2164 3459
rect 2158 3454 2159 3458
rect 2163 3454 2164 3458
rect 2158 3453 2164 3454
rect 2342 3458 2348 3459
rect 2342 3454 2343 3458
rect 2347 3454 2348 3458
rect 2342 3453 2348 3454
rect 2518 3458 2524 3459
rect 2518 3454 2519 3458
rect 2523 3454 2524 3458
rect 2518 3453 2524 3454
rect 2678 3458 2684 3459
rect 2678 3454 2679 3458
rect 2683 3454 2684 3458
rect 2678 3453 2684 3454
rect 2830 3458 2836 3459
rect 2830 3454 2831 3458
rect 2835 3454 2836 3458
rect 2830 3453 2836 3454
rect 2966 3458 2972 3459
rect 2966 3454 2967 3458
rect 2971 3454 2972 3458
rect 2966 3453 2972 3454
rect 3086 3458 3092 3459
rect 3086 3454 3087 3458
rect 3091 3454 3092 3458
rect 3086 3453 3092 3454
rect 3198 3458 3204 3459
rect 3198 3454 3199 3458
rect 3203 3454 3204 3458
rect 3198 3453 3204 3454
rect 3310 3458 3316 3459
rect 3310 3454 3311 3458
rect 3315 3454 3316 3458
rect 3310 3453 3316 3454
rect 3422 3458 3428 3459
rect 3422 3454 3423 3458
rect 3427 3454 3428 3458
rect 3422 3453 3428 3454
rect 3510 3458 3516 3459
rect 3510 3454 3511 3458
rect 3515 3454 3516 3458
rect 3510 3453 3516 3454
rect 110 3448 116 3449
rect 110 3444 111 3448
rect 115 3444 116 3448
rect 110 3443 116 3444
rect 1830 3448 1836 3449
rect 1830 3444 1831 3448
rect 1835 3444 1836 3448
rect 1830 3443 1836 3444
rect 1999 3447 2005 3448
rect 1999 3443 2000 3447
rect 2004 3446 2005 3447
rect 2034 3447 2040 3448
rect 2034 3446 2035 3447
rect 2004 3444 2035 3446
rect 2004 3443 2005 3444
rect 1999 3442 2005 3443
rect 2034 3443 2035 3444
rect 2039 3443 2040 3447
rect 2034 3442 2040 3443
rect 2178 3447 2189 3448
rect 2178 3443 2179 3447
rect 2183 3443 2184 3447
rect 2188 3443 2189 3447
rect 2178 3442 2189 3443
rect 2367 3447 2373 3448
rect 2367 3443 2368 3447
rect 2372 3446 2373 3447
rect 2402 3447 2408 3448
rect 2402 3446 2403 3447
rect 2372 3444 2403 3446
rect 2372 3443 2373 3444
rect 2367 3442 2373 3443
rect 2402 3443 2403 3444
rect 2407 3443 2408 3447
rect 2402 3442 2408 3443
rect 2543 3447 2549 3448
rect 2543 3443 2544 3447
rect 2548 3446 2549 3447
rect 2558 3447 2564 3448
rect 2558 3446 2559 3447
rect 2548 3444 2559 3446
rect 2548 3443 2549 3444
rect 2543 3442 2549 3443
rect 2558 3443 2559 3444
rect 2563 3443 2564 3447
rect 2558 3442 2564 3443
rect 2703 3447 2709 3448
rect 2703 3443 2704 3447
rect 2708 3446 2709 3447
rect 2738 3447 2744 3448
rect 2738 3446 2739 3447
rect 2708 3444 2739 3446
rect 2708 3443 2709 3444
rect 2703 3442 2709 3443
rect 2738 3443 2739 3444
rect 2743 3443 2744 3447
rect 2738 3442 2744 3443
rect 2854 3447 2861 3448
rect 2854 3443 2855 3447
rect 2860 3443 2861 3447
rect 2854 3442 2861 3443
rect 2986 3447 2997 3448
rect 2986 3443 2987 3447
rect 2991 3443 2992 3447
rect 2996 3443 2997 3447
rect 2986 3442 2997 3443
rect 3042 3447 3048 3448
rect 3042 3443 3043 3447
rect 3047 3446 3048 3447
rect 3111 3447 3117 3448
rect 3111 3446 3112 3447
rect 3047 3444 3112 3446
rect 3047 3443 3048 3444
rect 3042 3442 3048 3443
rect 3111 3443 3112 3444
rect 3116 3443 3117 3447
rect 3111 3442 3117 3443
rect 3158 3447 3164 3448
rect 3158 3443 3159 3447
rect 3163 3446 3164 3447
rect 3223 3447 3229 3448
rect 3223 3446 3224 3447
rect 3163 3444 3224 3446
rect 3163 3443 3164 3444
rect 3158 3442 3164 3443
rect 3223 3443 3224 3444
rect 3228 3443 3229 3447
rect 3223 3442 3229 3443
rect 3270 3447 3276 3448
rect 3270 3443 3271 3447
rect 3275 3446 3276 3447
rect 3335 3447 3341 3448
rect 3335 3446 3336 3447
rect 3275 3444 3336 3446
rect 3275 3443 3276 3444
rect 3270 3442 3276 3443
rect 3335 3443 3336 3444
rect 3340 3443 3341 3447
rect 3335 3442 3341 3443
rect 3382 3447 3388 3448
rect 3382 3443 3383 3447
rect 3387 3446 3388 3447
rect 3447 3447 3453 3448
rect 3447 3446 3448 3447
rect 3387 3444 3448 3446
rect 3387 3443 3388 3444
rect 3382 3442 3388 3443
rect 3447 3443 3448 3444
rect 3452 3443 3453 3447
rect 3447 3442 3453 3443
rect 3482 3447 3488 3448
rect 3482 3443 3483 3447
rect 3487 3446 3488 3447
rect 3535 3447 3541 3448
rect 3535 3446 3536 3447
rect 3487 3444 3536 3446
rect 3487 3443 3488 3444
rect 3482 3442 3488 3443
rect 3535 3443 3536 3444
rect 3540 3443 3541 3447
rect 3535 3442 3541 3443
rect 2052 3440 2162 3442
rect 374 3439 380 3440
rect 374 3435 375 3439
rect 379 3435 380 3439
rect 374 3434 380 3435
rect 554 3439 560 3440
rect 554 3435 555 3439
rect 559 3435 560 3439
rect 554 3434 560 3435
rect 674 3439 680 3440
rect 674 3435 675 3439
rect 679 3435 680 3439
rect 674 3434 680 3435
rect 786 3439 792 3440
rect 786 3435 787 3439
rect 791 3435 792 3439
rect 786 3434 792 3435
rect 846 3439 852 3440
rect 846 3435 847 3439
rect 851 3435 852 3439
rect 846 3434 852 3435
rect 994 3439 1000 3440
rect 994 3435 995 3439
rect 999 3435 1000 3439
rect 994 3434 1000 3435
rect 1090 3439 1096 3440
rect 1090 3435 1091 3439
rect 1095 3435 1096 3439
rect 1206 3439 1212 3440
rect 1206 3438 1207 3439
rect 1189 3436 1207 3438
rect 1090 3434 1096 3435
rect 1206 3435 1207 3436
rect 1211 3435 1212 3439
rect 1303 3439 1309 3440
rect 1303 3438 1304 3439
rect 1285 3436 1304 3438
rect 1206 3434 1212 3435
rect 1303 3435 1304 3436
rect 1308 3435 1309 3439
rect 1303 3434 1309 3435
rect 2031 3435 2037 3436
rect 110 3431 116 3432
rect 110 3427 111 3431
rect 115 3427 116 3431
rect 1830 3431 1836 3432
rect 110 3426 116 3427
rect 222 3428 228 3429
rect 222 3424 223 3428
rect 227 3424 228 3428
rect 222 3423 228 3424
rect 358 3428 364 3429
rect 358 3424 359 3428
rect 363 3424 364 3428
rect 358 3423 364 3424
rect 494 3428 500 3429
rect 494 3424 495 3428
rect 499 3424 500 3428
rect 494 3423 500 3424
rect 614 3428 620 3429
rect 614 3424 615 3428
rect 619 3424 620 3428
rect 614 3423 620 3424
rect 726 3428 732 3429
rect 726 3424 727 3428
rect 731 3424 732 3428
rect 726 3423 732 3424
rect 830 3428 836 3429
rect 830 3424 831 3428
rect 835 3424 836 3428
rect 830 3423 836 3424
rect 934 3428 940 3429
rect 934 3424 935 3428
rect 939 3424 940 3428
rect 934 3423 940 3424
rect 1030 3428 1036 3429
rect 1030 3424 1031 3428
rect 1035 3424 1036 3428
rect 1030 3423 1036 3424
rect 1126 3428 1132 3429
rect 1126 3424 1127 3428
rect 1131 3424 1132 3428
rect 1126 3423 1132 3424
rect 1222 3428 1228 3429
rect 1222 3424 1223 3428
rect 1227 3424 1228 3428
rect 1222 3423 1228 3424
rect 1318 3428 1324 3429
rect 1318 3424 1319 3428
rect 1323 3424 1324 3428
rect 1830 3427 1831 3431
rect 1835 3427 1836 3431
rect 2031 3431 2032 3435
rect 2036 3434 2037 3435
rect 2052 3434 2054 3440
rect 2160 3438 2162 3440
rect 2262 3439 2268 3440
rect 2262 3438 2263 3439
rect 2160 3436 2263 3438
rect 2036 3432 2054 3434
rect 2058 3435 2064 3436
rect 2036 3431 2037 3432
rect 2031 3430 2037 3431
rect 2058 3431 2059 3435
rect 2063 3434 2064 3435
rect 2151 3435 2157 3436
rect 2151 3434 2152 3435
rect 2063 3432 2152 3434
rect 2063 3431 2064 3432
rect 2058 3430 2064 3431
rect 2151 3431 2152 3432
rect 2156 3431 2157 3435
rect 2262 3435 2263 3436
rect 2267 3435 2268 3439
rect 2262 3434 2268 3435
rect 2279 3435 2288 3436
rect 2151 3430 2157 3431
rect 2279 3431 2280 3435
rect 2287 3431 2288 3435
rect 2279 3430 2288 3431
rect 2407 3435 2413 3436
rect 2407 3431 2408 3435
rect 2412 3434 2413 3435
rect 2415 3435 2421 3436
rect 2415 3434 2416 3435
rect 2412 3432 2416 3434
rect 2412 3431 2413 3432
rect 2407 3430 2413 3431
rect 2415 3431 2416 3432
rect 2420 3431 2421 3435
rect 2415 3430 2421 3431
rect 2442 3435 2448 3436
rect 2442 3431 2443 3435
rect 2447 3434 2448 3435
rect 2559 3435 2565 3436
rect 2559 3434 2560 3435
rect 2447 3432 2560 3434
rect 2447 3431 2448 3432
rect 2442 3430 2448 3431
rect 2559 3431 2560 3432
rect 2564 3431 2565 3435
rect 2559 3430 2565 3431
rect 2586 3435 2592 3436
rect 2586 3431 2587 3435
rect 2591 3434 2592 3435
rect 2703 3435 2709 3436
rect 2703 3434 2704 3435
rect 2591 3432 2704 3434
rect 2591 3431 2592 3432
rect 2586 3430 2592 3431
rect 2703 3431 2704 3432
rect 2708 3431 2709 3435
rect 2703 3430 2709 3431
rect 2855 3435 2861 3436
rect 2855 3431 2856 3435
rect 2860 3434 2861 3435
rect 3006 3435 3012 3436
rect 3006 3434 3007 3435
rect 2860 3432 3007 3434
rect 2860 3431 2861 3432
rect 2855 3430 2861 3431
rect 3006 3431 3007 3432
rect 3011 3431 3012 3435
rect 3006 3430 3012 3431
rect 3023 3435 3029 3436
rect 3023 3431 3024 3435
rect 3028 3434 3029 3435
rect 3174 3435 3180 3436
rect 3174 3434 3175 3435
rect 3028 3432 3175 3434
rect 3028 3431 3029 3432
rect 3023 3430 3029 3431
rect 3174 3431 3175 3432
rect 3179 3431 3180 3435
rect 3174 3430 3180 3431
rect 3191 3435 3197 3436
rect 3191 3431 3192 3435
rect 3196 3434 3197 3435
rect 3350 3435 3356 3436
rect 3350 3434 3351 3435
rect 3196 3432 3351 3434
rect 3196 3431 3197 3432
rect 3191 3430 3197 3431
rect 3350 3431 3351 3432
rect 3355 3431 3356 3435
rect 3350 3430 3356 3431
rect 3358 3435 3364 3436
rect 3358 3431 3359 3435
rect 3363 3434 3364 3435
rect 3367 3435 3373 3436
rect 3367 3434 3368 3435
rect 3363 3432 3368 3434
rect 3363 3431 3364 3432
rect 3358 3430 3364 3431
rect 3367 3431 3368 3432
rect 3372 3431 3373 3435
rect 3367 3430 3373 3431
rect 3535 3435 3541 3436
rect 3535 3431 3536 3435
rect 3540 3434 3541 3435
rect 3562 3435 3568 3436
rect 3562 3434 3563 3435
rect 3540 3432 3563 3434
rect 3540 3431 3541 3432
rect 3535 3430 3541 3431
rect 3562 3431 3563 3432
rect 3567 3431 3568 3435
rect 3562 3430 3568 3431
rect 1830 3426 1836 3427
rect 2006 3426 2012 3427
rect 1318 3423 1324 3424
rect 2006 3422 2007 3426
rect 2011 3422 2012 3426
rect 2006 3421 2012 3422
rect 2126 3426 2132 3427
rect 2126 3422 2127 3426
rect 2131 3422 2132 3426
rect 2126 3421 2132 3422
rect 2254 3426 2260 3427
rect 2254 3422 2255 3426
rect 2259 3422 2260 3426
rect 2254 3421 2260 3422
rect 2390 3426 2396 3427
rect 2390 3422 2391 3426
rect 2395 3422 2396 3426
rect 2390 3421 2396 3422
rect 2534 3426 2540 3427
rect 2534 3422 2535 3426
rect 2539 3422 2540 3426
rect 2534 3421 2540 3422
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2830 3426 2836 3427
rect 2830 3422 2831 3426
rect 2835 3422 2836 3426
rect 2830 3421 2836 3422
rect 2998 3426 3004 3427
rect 2998 3422 2999 3426
rect 3003 3422 3004 3426
rect 2998 3421 3004 3422
rect 3166 3426 3172 3427
rect 3166 3422 3167 3426
rect 3171 3422 3172 3426
rect 3166 3421 3172 3422
rect 3342 3426 3348 3427
rect 3342 3422 3343 3426
rect 3347 3422 3348 3426
rect 3342 3421 3348 3422
rect 3510 3426 3516 3427
rect 3510 3422 3511 3426
rect 3515 3422 3516 3426
rect 3510 3421 3516 3422
rect 239 3411 248 3412
rect 239 3407 240 3411
rect 247 3407 248 3411
rect 239 3406 248 3407
rect 1246 3411 1252 3412
rect 1246 3407 1247 3411
rect 1251 3410 1252 3411
rect 1335 3411 1341 3412
rect 1335 3410 1336 3411
rect 1251 3408 1336 3410
rect 1251 3407 1252 3408
rect 1246 3406 1252 3407
rect 1335 3407 1336 3408
rect 1340 3407 1341 3411
rect 1335 3406 1341 3407
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 2058 3399 2064 3400
rect 2058 3395 2059 3399
rect 2063 3395 2064 3399
rect 2058 3394 2064 3395
rect 2178 3399 2184 3400
rect 2178 3395 2179 3399
rect 2183 3395 2184 3399
rect 2178 3394 2184 3395
rect 2262 3399 2268 3400
rect 2262 3395 2263 3399
rect 2267 3395 2268 3399
rect 2262 3394 2268 3395
rect 2442 3399 2448 3400
rect 2442 3395 2443 3399
rect 2447 3395 2448 3399
rect 2442 3394 2448 3395
rect 2586 3399 2592 3400
rect 2586 3395 2587 3399
rect 2591 3395 2592 3399
rect 2586 3394 2592 3395
rect 2854 3399 2860 3400
rect 2854 3395 2855 3399
rect 2859 3395 2860 3399
rect 2854 3394 2860 3395
rect 3006 3399 3012 3400
rect 3006 3395 3007 3399
rect 3011 3395 3012 3399
rect 3006 3394 3012 3395
rect 3174 3399 3180 3400
rect 3174 3395 3175 3399
rect 3179 3395 3180 3399
rect 3174 3394 3180 3395
rect 3350 3399 3356 3400
rect 3350 3395 3351 3399
rect 3355 3395 3356 3399
rect 3350 3394 3356 3395
rect 3534 3399 3540 3400
rect 3534 3395 3535 3399
rect 3539 3395 3540 3399
rect 3534 3394 3540 3395
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 3590 3391 3596 3392
rect 1870 3386 1876 3387
rect 1998 3388 2004 3389
rect 1998 3384 1999 3388
rect 2003 3384 2004 3388
rect 1998 3383 2004 3384
rect 2118 3388 2124 3389
rect 2118 3384 2119 3388
rect 2123 3384 2124 3388
rect 2118 3383 2124 3384
rect 2246 3388 2252 3389
rect 2246 3384 2247 3388
rect 2251 3384 2252 3388
rect 2246 3383 2252 3384
rect 2382 3388 2388 3389
rect 2382 3384 2383 3388
rect 2387 3384 2388 3388
rect 2382 3383 2388 3384
rect 2526 3388 2532 3389
rect 2526 3384 2527 3388
rect 2531 3384 2532 3388
rect 2526 3383 2532 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2822 3388 2828 3389
rect 2822 3384 2823 3388
rect 2827 3384 2828 3388
rect 2822 3383 2828 3384
rect 2990 3388 2996 3389
rect 2990 3384 2991 3388
rect 2995 3384 2996 3388
rect 2990 3383 2996 3384
rect 3158 3388 3164 3389
rect 3158 3384 3159 3388
rect 3163 3384 3164 3388
rect 3158 3383 3164 3384
rect 3334 3388 3340 3389
rect 3334 3384 3335 3388
rect 3339 3384 3340 3388
rect 3334 3383 3340 3384
rect 3502 3388 3508 3389
rect 3502 3384 3503 3388
rect 3507 3384 3508 3388
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3502 3383 3508 3384
rect 214 3380 220 3381
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 214 3376 215 3380
rect 219 3376 220 3380
rect 214 3375 220 3376
rect 366 3380 372 3381
rect 366 3376 367 3380
rect 371 3376 372 3380
rect 366 3375 372 3376
rect 510 3380 516 3381
rect 510 3376 511 3380
rect 515 3376 516 3380
rect 510 3375 516 3376
rect 646 3380 652 3381
rect 646 3376 647 3380
rect 651 3376 652 3380
rect 646 3375 652 3376
rect 774 3380 780 3381
rect 774 3376 775 3380
rect 779 3376 780 3380
rect 774 3375 780 3376
rect 894 3380 900 3381
rect 894 3376 895 3380
rect 899 3376 900 3380
rect 894 3375 900 3376
rect 1014 3380 1020 3381
rect 1014 3376 1015 3380
rect 1019 3376 1020 3380
rect 1014 3375 1020 3376
rect 1126 3380 1132 3381
rect 1126 3376 1127 3380
rect 1131 3376 1132 3380
rect 1126 3375 1132 3376
rect 1238 3380 1244 3381
rect 1238 3376 1239 3380
rect 1243 3376 1244 3380
rect 1238 3375 1244 3376
rect 1350 3380 1356 3381
rect 1350 3376 1351 3380
rect 1355 3376 1356 3380
rect 1350 3375 1356 3376
rect 1830 3377 1836 3378
rect 110 3372 116 3373
rect 1830 3373 1831 3377
rect 1835 3373 1836 3377
rect 1830 3372 1836 3373
rect 282 3371 288 3372
rect 282 3370 283 3371
rect 277 3368 283 3370
rect 282 3367 283 3368
rect 287 3367 288 3371
rect 578 3371 584 3372
rect 376 3368 385 3370
rect 282 3366 288 3367
rect 374 3367 380 3368
rect 374 3363 375 3367
rect 379 3363 380 3367
rect 374 3362 380 3363
rect 518 3367 524 3368
rect 518 3363 519 3367
rect 523 3366 524 3367
rect 528 3366 530 3369
rect 578 3367 579 3371
rect 583 3370 584 3371
rect 714 3371 720 3372
rect 583 3368 665 3370
rect 583 3367 584 3368
rect 578 3366 584 3367
rect 714 3367 715 3371
rect 719 3370 720 3371
rect 975 3371 981 3372
rect 975 3370 976 3371
rect 719 3368 793 3370
rect 957 3368 976 3370
rect 719 3367 720 3368
rect 714 3366 720 3367
rect 975 3367 976 3368
rect 980 3367 981 3371
rect 1094 3371 1100 3372
rect 1094 3370 1095 3371
rect 1077 3368 1095 3370
rect 975 3366 981 3367
rect 1094 3367 1095 3368
rect 1099 3367 1100 3371
rect 1206 3371 1212 3372
rect 1206 3370 1207 3371
rect 1189 3368 1207 3370
rect 1094 3366 1100 3367
rect 1206 3367 1207 3368
rect 1211 3367 1212 3371
rect 1318 3371 1324 3372
rect 1318 3370 1319 3371
rect 1301 3368 1319 3370
rect 1206 3366 1212 3367
rect 1318 3367 1319 3368
rect 1323 3367 1324 3371
rect 1318 3366 1324 3367
rect 1326 3371 1332 3372
rect 1326 3367 1327 3371
rect 1331 3370 1332 3371
rect 2618 3371 2624 3372
rect 1331 3368 1369 3370
rect 1331 3367 1332 3368
rect 1326 3366 1332 3367
rect 2618 3367 2619 3371
rect 2623 3370 2624 3371
rect 2687 3371 2693 3372
rect 2687 3370 2688 3371
rect 2623 3368 2688 3370
rect 2623 3367 2624 3368
rect 2618 3366 2624 3367
rect 2687 3367 2688 3368
rect 2692 3367 2693 3371
rect 2687 3366 2693 3367
rect 523 3364 530 3366
rect 523 3363 524 3364
rect 518 3362 524 3363
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 1830 3360 1836 3361
rect 1830 3356 1831 3360
rect 1835 3356 1836 3360
rect 1830 3355 1836 3356
rect 2014 3344 2020 3345
rect 222 3342 228 3343
rect 222 3338 223 3342
rect 227 3338 228 3342
rect 222 3337 228 3338
rect 374 3342 380 3343
rect 374 3338 375 3342
rect 379 3338 380 3342
rect 374 3337 380 3338
rect 518 3342 524 3343
rect 518 3338 519 3342
rect 523 3338 524 3342
rect 518 3337 524 3338
rect 654 3342 660 3343
rect 654 3338 655 3342
rect 659 3338 660 3342
rect 654 3337 660 3338
rect 782 3342 788 3343
rect 782 3338 783 3342
rect 787 3338 788 3342
rect 782 3337 788 3338
rect 902 3342 908 3343
rect 902 3338 903 3342
rect 907 3338 908 3342
rect 902 3337 908 3338
rect 1022 3342 1028 3343
rect 1022 3338 1023 3342
rect 1027 3338 1028 3342
rect 1022 3337 1028 3338
rect 1134 3342 1140 3343
rect 1134 3338 1135 3342
rect 1139 3338 1140 3342
rect 1134 3337 1140 3338
rect 1246 3342 1252 3343
rect 1246 3338 1247 3342
rect 1251 3338 1252 3342
rect 1246 3337 1252 3338
rect 1358 3342 1364 3343
rect 1358 3338 1359 3342
rect 1363 3338 1364 3342
rect 1358 3337 1364 3338
rect 1870 3341 1876 3342
rect 1870 3337 1871 3341
rect 1875 3337 1876 3341
rect 2014 3340 2015 3344
rect 2019 3340 2020 3344
rect 2014 3339 2020 3340
rect 2150 3344 2156 3345
rect 2150 3340 2151 3344
rect 2155 3340 2156 3344
rect 2150 3339 2156 3340
rect 2294 3344 2300 3345
rect 2294 3340 2295 3344
rect 2299 3340 2300 3344
rect 2294 3339 2300 3340
rect 2438 3344 2444 3345
rect 2438 3340 2439 3344
rect 2443 3340 2444 3344
rect 2438 3339 2444 3340
rect 2582 3344 2588 3345
rect 2582 3340 2583 3344
rect 2587 3340 2588 3344
rect 2582 3339 2588 3340
rect 2726 3344 2732 3345
rect 2726 3340 2727 3344
rect 2731 3340 2732 3344
rect 2726 3339 2732 3340
rect 2870 3344 2876 3345
rect 2870 3340 2871 3344
rect 2875 3340 2876 3344
rect 2870 3339 2876 3340
rect 3022 3344 3028 3345
rect 3022 3340 3023 3344
rect 3027 3340 3028 3344
rect 3022 3339 3028 3340
rect 3182 3344 3188 3345
rect 3182 3340 3183 3344
rect 3187 3340 3188 3344
rect 3182 3339 3188 3340
rect 3350 3344 3356 3345
rect 3350 3340 3351 3344
rect 3355 3340 3356 3344
rect 3350 3339 3356 3340
rect 3502 3344 3508 3345
rect 3502 3340 3503 3344
rect 3507 3340 3508 3344
rect 3502 3339 3508 3340
rect 3590 3341 3596 3342
rect 1870 3336 1876 3337
rect 3590 3337 3591 3341
rect 3595 3337 3596 3341
rect 3590 3336 3596 3337
rect 2106 3335 2112 3336
rect 2106 3334 2107 3335
rect 2077 3332 2107 3334
rect 242 3331 253 3332
rect 242 3327 243 3331
rect 247 3327 248 3331
rect 252 3327 253 3331
rect 242 3326 253 3327
rect 282 3331 288 3332
rect 282 3327 283 3331
rect 287 3330 288 3331
rect 399 3331 405 3332
rect 399 3330 400 3331
rect 287 3328 400 3330
rect 287 3327 288 3328
rect 282 3326 288 3327
rect 399 3327 400 3328
rect 404 3327 405 3331
rect 399 3326 405 3327
rect 543 3331 549 3332
rect 543 3327 544 3331
rect 548 3330 549 3331
rect 578 3331 584 3332
rect 578 3330 579 3331
rect 548 3328 579 3330
rect 548 3327 549 3328
rect 543 3326 549 3327
rect 578 3327 579 3328
rect 583 3327 584 3331
rect 578 3326 584 3327
rect 679 3331 685 3332
rect 679 3327 680 3331
rect 684 3330 685 3331
rect 714 3331 720 3332
rect 714 3330 715 3331
rect 684 3328 715 3330
rect 684 3327 685 3328
rect 679 3326 685 3327
rect 714 3327 715 3328
rect 719 3327 720 3331
rect 714 3326 720 3327
rect 807 3331 813 3332
rect 807 3327 808 3331
rect 812 3330 813 3331
rect 822 3331 828 3332
rect 822 3330 823 3331
rect 812 3328 823 3330
rect 812 3327 813 3328
rect 807 3326 813 3327
rect 822 3327 823 3328
rect 827 3327 828 3331
rect 822 3326 828 3327
rect 926 3331 933 3332
rect 926 3327 927 3331
rect 932 3327 933 3331
rect 926 3326 933 3327
rect 975 3331 981 3332
rect 975 3327 976 3331
rect 980 3330 981 3331
rect 1047 3331 1053 3332
rect 1047 3330 1048 3331
rect 980 3328 1048 3330
rect 980 3327 981 3328
rect 975 3326 981 3327
rect 1047 3327 1048 3328
rect 1052 3327 1053 3331
rect 1047 3326 1053 3327
rect 1094 3331 1100 3332
rect 1094 3327 1095 3331
rect 1099 3330 1100 3331
rect 1159 3331 1165 3332
rect 1159 3330 1160 3331
rect 1099 3328 1160 3330
rect 1099 3327 1100 3328
rect 1094 3326 1100 3327
rect 1159 3327 1160 3328
rect 1164 3327 1165 3331
rect 1159 3326 1165 3327
rect 1206 3331 1212 3332
rect 1206 3327 1207 3331
rect 1211 3330 1212 3331
rect 1271 3331 1277 3332
rect 1271 3330 1272 3331
rect 1211 3328 1272 3330
rect 1211 3327 1212 3328
rect 1206 3326 1212 3327
rect 1271 3327 1272 3328
rect 1276 3327 1277 3331
rect 1271 3326 1277 3327
rect 1318 3331 1324 3332
rect 1318 3327 1319 3331
rect 1323 3330 1324 3331
rect 1383 3331 1389 3332
rect 1383 3330 1384 3331
rect 1323 3328 1384 3330
rect 1323 3327 1324 3328
rect 1318 3326 1324 3327
rect 1383 3327 1384 3328
rect 1388 3327 1389 3331
rect 2106 3331 2107 3332
rect 2111 3331 2112 3335
rect 2246 3335 2252 3336
rect 2246 3334 2247 3335
rect 2213 3332 2247 3334
rect 2106 3330 2112 3331
rect 2246 3331 2247 3332
rect 2251 3331 2252 3335
rect 2246 3330 2252 3331
rect 2282 3335 2288 3336
rect 2282 3331 2283 3335
rect 2287 3334 2288 3335
rect 2506 3335 2512 3336
rect 2287 3332 2313 3334
rect 2287 3331 2288 3332
rect 2282 3330 2288 3331
rect 2500 3328 2502 3333
rect 2506 3331 2507 3335
rect 2511 3334 2512 3335
rect 2794 3335 2800 3336
rect 2794 3334 2795 3335
rect 2511 3332 2601 3334
rect 2789 3332 2795 3334
rect 2511 3331 2512 3332
rect 2506 3330 2512 3331
rect 2794 3331 2795 3332
rect 2799 3331 2800 3335
rect 2970 3335 2976 3336
rect 2970 3334 2971 3335
rect 2933 3332 2971 3334
rect 2794 3330 2800 3331
rect 2970 3331 2971 3332
rect 2975 3331 2976 3335
rect 3126 3335 3132 3336
rect 3126 3334 3127 3335
rect 3085 3332 3127 3334
rect 2970 3330 2976 3331
rect 3126 3331 3127 3332
rect 3131 3331 3132 3335
rect 3290 3335 3296 3336
rect 3290 3334 3291 3335
rect 3245 3332 3291 3334
rect 3126 3330 3132 3331
rect 3290 3331 3291 3332
rect 3295 3331 3296 3335
rect 3290 3330 3296 3331
rect 3358 3331 3364 3332
rect 1383 3326 1389 3327
rect 2498 3327 2504 3328
rect 1870 3324 1876 3325
rect 1870 3320 1871 3324
rect 1875 3320 1876 3324
rect 2498 3323 2499 3327
rect 2503 3323 2504 3327
rect 3358 3327 3359 3331
rect 3363 3330 3364 3331
rect 3368 3330 3370 3333
rect 3363 3328 3370 3330
rect 3564 3328 3566 3333
rect 3363 3327 3364 3328
rect 3358 3326 3364 3327
rect 3562 3327 3568 3328
rect 2498 3322 2504 3323
rect 3562 3323 3563 3327
rect 3567 3323 3568 3327
rect 3562 3322 3568 3323
rect 3590 3324 3596 3325
rect 1870 3319 1876 3320
rect 3590 3320 3591 3324
rect 3595 3320 3596 3324
rect 3590 3319 3596 3320
rect 231 3315 237 3316
rect 231 3311 232 3315
rect 236 3314 237 3315
rect 298 3315 304 3316
rect 298 3314 299 3315
rect 236 3312 299 3314
rect 236 3311 237 3312
rect 231 3310 237 3311
rect 298 3311 299 3312
rect 303 3311 304 3315
rect 298 3310 304 3311
rect 382 3315 388 3316
rect 382 3311 383 3315
rect 387 3314 388 3315
rect 391 3315 397 3316
rect 391 3314 392 3315
rect 387 3312 392 3314
rect 387 3311 388 3312
rect 382 3310 388 3311
rect 391 3311 392 3312
rect 396 3311 397 3315
rect 391 3310 397 3311
rect 543 3315 552 3316
rect 543 3311 544 3315
rect 551 3311 552 3315
rect 543 3310 552 3311
rect 570 3315 576 3316
rect 570 3311 571 3315
rect 575 3314 576 3315
rect 695 3315 701 3316
rect 695 3314 696 3315
rect 575 3312 696 3314
rect 575 3311 576 3312
rect 570 3310 576 3311
rect 695 3311 696 3312
rect 700 3311 701 3315
rect 695 3310 701 3311
rect 722 3315 728 3316
rect 722 3311 723 3315
rect 727 3314 728 3315
rect 839 3315 845 3316
rect 839 3314 840 3315
rect 727 3312 840 3314
rect 727 3311 728 3312
rect 722 3310 728 3311
rect 839 3311 840 3312
rect 844 3311 845 3315
rect 839 3310 845 3311
rect 975 3315 984 3316
rect 975 3311 976 3315
rect 983 3311 984 3315
rect 975 3310 984 3311
rect 1002 3315 1008 3316
rect 1002 3311 1003 3315
rect 1007 3314 1008 3315
rect 1111 3315 1117 3316
rect 1111 3314 1112 3315
rect 1007 3312 1112 3314
rect 1007 3311 1008 3312
rect 1002 3310 1008 3311
rect 1111 3311 1112 3312
rect 1116 3311 1117 3315
rect 1111 3310 1117 3311
rect 1166 3315 1172 3316
rect 1166 3311 1167 3315
rect 1171 3314 1172 3315
rect 1239 3315 1245 3316
rect 1239 3314 1240 3315
rect 1171 3312 1240 3314
rect 1171 3311 1172 3312
rect 1166 3310 1172 3311
rect 1239 3311 1240 3312
rect 1244 3311 1245 3315
rect 1239 3310 1245 3311
rect 1266 3315 1272 3316
rect 1266 3311 1267 3315
rect 1271 3314 1272 3315
rect 1367 3315 1373 3316
rect 1367 3314 1368 3315
rect 1271 3312 1368 3314
rect 1271 3311 1272 3312
rect 1266 3310 1272 3311
rect 1367 3311 1368 3312
rect 1372 3311 1373 3315
rect 1367 3310 1373 3311
rect 1394 3315 1400 3316
rect 1394 3311 1395 3315
rect 1399 3314 1400 3315
rect 1495 3315 1501 3316
rect 1495 3314 1496 3315
rect 1399 3312 1496 3314
rect 1399 3311 1400 3312
rect 1394 3310 1400 3311
rect 1495 3311 1496 3312
rect 1500 3311 1501 3315
rect 1495 3310 1501 3311
rect 206 3306 212 3307
rect 206 3302 207 3306
rect 211 3302 212 3306
rect 206 3301 212 3302
rect 366 3306 372 3307
rect 366 3302 367 3306
rect 371 3302 372 3306
rect 366 3301 372 3302
rect 518 3306 524 3307
rect 518 3302 519 3306
rect 523 3302 524 3306
rect 518 3301 524 3302
rect 670 3306 676 3307
rect 670 3302 671 3306
rect 675 3302 676 3306
rect 670 3301 676 3302
rect 814 3306 820 3307
rect 814 3302 815 3306
rect 819 3302 820 3306
rect 814 3301 820 3302
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1086 3306 1092 3307
rect 1086 3302 1087 3306
rect 1091 3302 1092 3306
rect 1086 3301 1092 3302
rect 1214 3306 1220 3307
rect 1214 3302 1215 3306
rect 1219 3302 1220 3306
rect 1214 3301 1220 3302
rect 1342 3306 1348 3307
rect 1342 3302 1343 3306
rect 1347 3302 1348 3306
rect 1342 3301 1348 3302
rect 1470 3306 1476 3307
rect 1470 3302 1471 3306
rect 1475 3302 1476 3306
rect 1470 3301 1476 3302
rect 2022 3306 2028 3307
rect 2022 3302 2023 3306
rect 2027 3302 2028 3306
rect 2022 3301 2028 3302
rect 2158 3306 2164 3307
rect 2158 3302 2159 3306
rect 2163 3302 2164 3306
rect 2158 3301 2164 3302
rect 2302 3306 2308 3307
rect 2302 3302 2303 3306
rect 2307 3302 2308 3306
rect 2302 3301 2308 3302
rect 2446 3306 2452 3307
rect 2446 3302 2447 3306
rect 2451 3302 2452 3306
rect 2446 3301 2452 3302
rect 2590 3306 2596 3307
rect 2590 3302 2591 3306
rect 2595 3302 2596 3306
rect 2590 3301 2596 3302
rect 2734 3306 2740 3307
rect 2734 3302 2735 3306
rect 2739 3302 2740 3306
rect 2734 3301 2740 3302
rect 2878 3306 2884 3307
rect 2878 3302 2879 3306
rect 2883 3302 2884 3306
rect 2878 3301 2884 3302
rect 3030 3306 3036 3307
rect 3030 3302 3031 3306
rect 3035 3302 3036 3306
rect 3030 3301 3036 3302
rect 3190 3306 3196 3307
rect 3190 3302 3191 3306
rect 3195 3302 3196 3306
rect 3190 3301 3196 3302
rect 3358 3306 3364 3307
rect 3358 3302 3359 3306
rect 3363 3302 3364 3306
rect 3358 3301 3364 3302
rect 3510 3306 3516 3307
rect 3510 3302 3511 3306
rect 3515 3302 3516 3306
rect 3510 3301 3516 3302
rect 1978 3295 1984 3296
rect 1978 3291 1979 3295
rect 1983 3294 1984 3295
rect 2047 3295 2053 3296
rect 2047 3294 2048 3295
rect 1983 3292 2048 3294
rect 1983 3291 1984 3292
rect 1978 3290 1984 3291
rect 2047 3291 2048 3292
rect 2052 3291 2053 3295
rect 2047 3290 2053 3291
rect 2106 3295 2112 3296
rect 2106 3291 2107 3295
rect 2111 3294 2112 3295
rect 2183 3295 2189 3296
rect 2183 3294 2184 3295
rect 2111 3292 2184 3294
rect 2111 3291 2112 3292
rect 2106 3290 2112 3291
rect 2183 3291 2184 3292
rect 2188 3291 2189 3295
rect 2183 3290 2189 3291
rect 2246 3295 2252 3296
rect 2246 3291 2247 3295
rect 2251 3294 2252 3295
rect 2327 3295 2333 3296
rect 2327 3294 2328 3295
rect 2251 3292 2328 3294
rect 2251 3291 2252 3292
rect 2246 3290 2252 3291
rect 2327 3291 2328 3292
rect 2332 3291 2333 3295
rect 2327 3290 2333 3291
rect 2471 3295 2477 3296
rect 2471 3291 2472 3295
rect 2476 3294 2477 3295
rect 2506 3295 2512 3296
rect 2506 3294 2507 3295
rect 2476 3292 2507 3294
rect 2476 3291 2477 3292
rect 2471 3290 2477 3291
rect 2506 3291 2507 3292
rect 2511 3291 2512 3295
rect 2506 3290 2512 3291
rect 2615 3295 2624 3296
rect 2615 3291 2616 3295
rect 2623 3291 2624 3295
rect 2615 3290 2624 3291
rect 2759 3295 2765 3296
rect 2759 3291 2760 3295
rect 2764 3294 2765 3295
rect 2786 3295 2792 3296
rect 2786 3294 2787 3295
rect 2764 3292 2787 3294
rect 2764 3291 2765 3292
rect 2759 3290 2765 3291
rect 2786 3291 2787 3292
rect 2791 3291 2792 3295
rect 2786 3290 2792 3291
rect 2794 3295 2800 3296
rect 2794 3291 2795 3295
rect 2799 3294 2800 3295
rect 2903 3295 2909 3296
rect 2903 3294 2904 3295
rect 2799 3292 2904 3294
rect 2799 3291 2800 3292
rect 2794 3290 2800 3291
rect 2903 3291 2904 3292
rect 2908 3291 2909 3295
rect 2903 3290 2909 3291
rect 2970 3295 2976 3296
rect 2970 3291 2971 3295
rect 2975 3294 2976 3295
rect 3055 3295 3061 3296
rect 3055 3294 3056 3295
rect 2975 3292 3056 3294
rect 2975 3291 2976 3292
rect 2970 3290 2976 3291
rect 3055 3291 3056 3292
rect 3060 3291 3061 3295
rect 3055 3290 3061 3291
rect 3126 3295 3132 3296
rect 3126 3291 3127 3295
rect 3131 3294 3132 3295
rect 3215 3295 3221 3296
rect 3215 3294 3216 3295
rect 3131 3292 3216 3294
rect 3131 3291 3132 3292
rect 3126 3290 3132 3291
rect 3215 3291 3216 3292
rect 3220 3291 3221 3295
rect 3215 3290 3221 3291
rect 3290 3295 3296 3296
rect 3290 3291 3291 3295
rect 3295 3294 3296 3295
rect 3383 3295 3389 3296
rect 3383 3294 3384 3295
rect 3295 3292 3384 3294
rect 3295 3291 3296 3292
rect 3290 3290 3296 3291
rect 3383 3291 3384 3292
rect 3388 3291 3389 3295
rect 3383 3290 3389 3291
rect 3534 3295 3541 3296
rect 3534 3291 3535 3295
rect 3540 3291 3541 3295
rect 3534 3290 3541 3291
rect 110 3288 116 3289
rect 110 3284 111 3288
rect 115 3284 116 3288
rect 110 3283 116 3284
rect 1830 3288 1836 3289
rect 1830 3284 1831 3288
rect 1835 3284 1836 3288
rect 1830 3283 1836 3284
rect 1951 3283 1957 3284
rect 258 3279 264 3280
rect 258 3275 259 3279
rect 263 3275 264 3279
rect 258 3274 264 3275
rect 298 3279 304 3280
rect 298 3275 299 3279
rect 303 3278 304 3279
rect 570 3279 576 3280
rect 303 3276 377 3278
rect 303 3275 304 3276
rect 298 3274 304 3275
rect 570 3275 571 3279
rect 575 3275 576 3279
rect 570 3274 576 3275
rect 722 3279 728 3280
rect 722 3275 723 3279
rect 727 3275 728 3279
rect 722 3274 728 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 1002 3279 1008 3280
rect 1002 3275 1003 3279
rect 1007 3275 1008 3279
rect 1166 3279 1172 3280
rect 1166 3278 1167 3279
rect 1141 3276 1167 3278
rect 1002 3274 1008 3275
rect 1166 3275 1167 3276
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1266 3279 1272 3280
rect 1266 3275 1267 3279
rect 1271 3275 1272 3279
rect 1266 3274 1272 3275
rect 1394 3279 1400 3280
rect 1394 3275 1395 3279
rect 1399 3275 1400 3279
rect 1951 3279 1952 3283
rect 1956 3282 1957 3283
rect 2070 3283 2076 3284
rect 2070 3282 2071 3283
rect 1956 3280 2071 3282
rect 1956 3279 1957 3280
rect 1951 3278 1957 3279
rect 2070 3279 2071 3280
rect 2075 3279 2076 3283
rect 2070 3278 2076 3279
rect 2087 3283 2093 3284
rect 2087 3279 2088 3283
rect 2092 3282 2093 3283
rect 2198 3283 2204 3284
rect 2198 3282 2199 3283
rect 2092 3280 2199 3282
rect 2092 3279 2093 3280
rect 2087 3278 2093 3279
rect 2198 3279 2199 3280
rect 2203 3279 2204 3283
rect 2198 3278 2204 3279
rect 2210 3283 2221 3284
rect 2210 3279 2211 3283
rect 2215 3279 2216 3283
rect 2220 3279 2221 3283
rect 2210 3278 2221 3279
rect 2343 3283 2349 3284
rect 2343 3279 2344 3283
rect 2348 3282 2349 3283
rect 2454 3283 2460 3284
rect 2454 3282 2455 3283
rect 2348 3280 2455 3282
rect 2348 3279 2349 3280
rect 2343 3278 2349 3279
rect 2454 3279 2455 3280
rect 2459 3279 2460 3283
rect 2454 3278 2460 3279
rect 2471 3283 2477 3284
rect 2471 3279 2472 3283
rect 2476 3282 2477 3283
rect 2498 3283 2504 3284
rect 2498 3282 2499 3283
rect 2476 3280 2499 3282
rect 2476 3279 2477 3280
rect 2471 3278 2477 3279
rect 2498 3279 2499 3280
rect 2503 3279 2504 3283
rect 2498 3278 2504 3279
rect 2614 3283 2621 3284
rect 2614 3279 2615 3283
rect 2620 3279 2621 3283
rect 2614 3278 2621 3279
rect 2642 3283 2648 3284
rect 2642 3279 2643 3283
rect 2647 3282 2648 3283
rect 2767 3283 2773 3284
rect 2767 3282 2768 3283
rect 2647 3280 2768 3282
rect 2647 3279 2648 3280
rect 2642 3278 2648 3279
rect 2767 3279 2768 3280
rect 2772 3279 2773 3283
rect 2767 3278 2773 3279
rect 2794 3283 2800 3284
rect 2794 3279 2795 3283
rect 2799 3282 2800 3283
rect 2943 3283 2949 3284
rect 2943 3282 2944 3283
rect 2799 3280 2944 3282
rect 2799 3279 2800 3280
rect 2794 3278 2800 3279
rect 2943 3279 2944 3280
rect 2948 3279 2949 3283
rect 2943 3278 2949 3279
rect 2970 3283 2976 3284
rect 2970 3279 2971 3283
rect 2975 3282 2976 3283
rect 3135 3283 3141 3284
rect 3135 3282 3136 3283
rect 2975 3280 3136 3282
rect 2975 3279 2976 3280
rect 2970 3278 2976 3279
rect 3135 3279 3136 3280
rect 3140 3279 3141 3283
rect 3135 3278 3141 3279
rect 3162 3283 3168 3284
rect 3162 3279 3163 3283
rect 3167 3282 3168 3283
rect 3335 3283 3341 3284
rect 3335 3282 3336 3283
rect 3167 3280 3336 3282
rect 3167 3279 3168 3280
rect 3162 3278 3168 3279
rect 3335 3279 3336 3280
rect 3340 3279 3341 3283
rect 3335 3278 3341 3279
rect 3535 3283 3541 3284
rect 3535 3279 3536 3283
rect 3540 3282 3541 3283
rect 3562 3283 3568 3284
rect 3562 3282 3563 3283
rect 3540 3280 3563 3282
rect 3540 3279 3541 3280
rect 3535 3278 3541 3279
rect 3562 3279 3563 3280
rect 3567 3279 3568 3283
rect 3562 3278 3568 3279
rect 1394 3274 1400 3275
rect 1926 3274 1932 3275
rect 110 3271 116 3272
rect 110 3267 111 3271
rect 115 3267 116 3271
rect 1830 3271 1836 3272
rect 110 3266 116 3267
rect 198 3268 204 3269
rect 198 3264 199 3268
rect 203 3264 204 3268
rect 198 3263 204 3264
rect 358 3268 364 3269
rect 358 3264 359 3268
rect 363 3264 364 3268
rect 358 3263 364 3264
rect 510 3268 516 3269
rect 510 3264 511 3268
rect 515 3264 516 3268
rect 510 3263 516 3264
rect 662 3268 668 3269
rect 662 3264 663 3268
rect 667 3264 668 3268
rect 662 3263 668 3264
rect 806 3268 812 3269
rect 806 3264 807 3268
rect 811 3264 812 3268
rect 806 3263 812 3264
rect 942 3268 948 3269
rect 942 3264 943 3268
rect 947 3264 948 3268
rect 942 3263 948 3264
rect 1078 3268 1084 3269
rect 1078 3264 1079 3268
rect 1083 3264 1084 3268
rect 1078 3263 1084 3264
rect 1206 3268 1212 3269
rect 1206 3264 1207 3268
rect 1211 3264 1212 3268
rect 1206 3263 1212 3264
rect 1334 3268 1340 3269
rect 1334 3264 1335 3268
rect 1339 3264 1340 3268
rect 1334 3263 1340 3264
rect 1462 3268 1468 3269
rect 1462 3264 1463 3268
rect 1467 3264 1468 3268
rect 1830 3267 1831 3271
rect 1835 3267 1836 3271
rect 1926 3270 1927 3274
rect 1931 3270 1932 3274
rect 1926 3269 1932 3270
rect 2062 3274 2068 3275
rect 2062 3270 2063 3274
rect 2067 3270 2068 3274
rect 2062 3269 2068 3270
rect 2190 3274 2196 3275
rect 2190 3270 2191 3274
rect 2195 3270 2196 3274
rect 2190 3269 2196 3270
rect 2318 3274 2324 3275
rect 2318 3270 2319 3274
rect 2323 3270 2324 3274
rect 2318 3269 2324 3270
rect 2446 3274 2452 3275
rect 2446 3270 2447 3274
rect 2451 3270 2452 3274
rect 2446 3269 2452 3270
rect 2590 3274 2596 3275
rect 2590 3270 2591 3274
rect 2595 3270 2596 3274
rect 2590 3269 2596 3270
rect 2742 3274 2748 3275
rect 2742 3270 2743 3274
rect 2747 3270 2748 3274
rect 2742 3269 2748 3270
rect 2918 3274 2924 3275
rect 2918 3270 2919 3274
rect 2923 3270 2924 3274
rect 2918 3269 2924 3270
rect 3110 3274 3116 3275
rect 3110 3270 3111 3274
rect 3115 3270 3116 3274
rect 3110 3269 3116 3270
rect 3310 3274 3316 3275
rect 3310 3270 3311 3274
rect 3315 3270 3316 3274
rect 3310 3269 3316 3270
rect 3510 3274 3516 3275
rect 3510 3270 3511 3274
rect 3515 3270 3516 3274
rect 3510 3269 3516 3270
rect 1830 3266 1836 3267
rect 1462 3263 1468 3264
rect 1870 3256 1876 3257
rect 1870 3252 1871 3256
rect 1875 3252 1876 3256
rect 1398 3251 1404 3252
rect 1398 3247 1399 3251
rect 1403 3250 1404 3251
rect 1479 3251 1485 3252
rect 1870 3251 1876 3252
rect 3590 3256 3596 3257
rect 3590 3252 3591 3256
rect 3595 3252 3596 3256
rect 3590 3251 3596 3252
rect 1479 3250 1480 3251
rect 1403 3248 1480 3250
rect 1403 3247 1404 3248
rect 1398 3246 1404 3247
rect 1479 3247 1480 3248
rect 1484 3247 1485 3251
rect 1479 3246 1485 3247
rect 1978 3247 1984 3248
rect 1978 3243 1979 3247
rect 1983 3243 1984 3247
rect 1978 3242 1984 3243
rect 2070 3247 2076 3248
rect 2070 3243 2071 3247
rect 2075 3243 2076 3247
rect 2070 3242 2076 3243
rect 2198 3247 2204 3248
rect 2198 3243 2199 3247
rect 2203 3243 2204 3247
rect 2198 3242 2204 3243
rect 2454 3247 2460 3248
rect 2454 3243 2455 3247
rect 2459 3243 2460 3247
rect 2454 3242 2460 3243
rect 2642 3247 2648 3248
rect 2642 3243 2643 3247
rect 2647 3243 2648 3247
rect 2642 3242 2648 3243
rect 2794 3247 2800 3248
rect 2794 3243 2795 3247
rect 2799 3243 2800 3247
rect 2794 3242 2800 3243
rect 2970 3247 2976 3248
rect 2970 3243 2971 3247
rect 2975 3243 2976 3247
rect 2970 3242 2976 3243
rect 3162 3247 3168 3248
rect 3162 3243 3163 3247
rect 3167 3243 3168 3247
rect 3162 3242 3168 3243
rect 3318 3247 3324 3248
rect 3318 3243 3319 3247
rect 3323 3243 3324 3247
rect 3318 3242 3324 3243
rect 3534 3247 3540 3248
rect 3534 3243 3535 3247
rect 3539 3243 3540 3247
rect 3534 3242 3540 3243
rect 1870 3239 1876 3240
rect 1870 3235 1871 3239
rect 1875 3235 1876 3239
rect 3590 3239 3596 3240
rect 1870 3234 1876 3235
rect 1918 3236 1924 3237
rect 1918 3232 1919 3236
rect 1923 3232 1924 3236
rect 1918 3231 1924 3232
rect 2054 3236 2060 3237
rect 2054 3232 2055 3236
rect 2059 3232 2060 3236
rect 2054 3231 2060 3232
rect 2182 3236 2188 3237
rect 2182 3232 2183 3236
rect 2187 3232 2188 3236
rect 2182 3231 2188 3232
rect 2310 3236 2316 3237
rect 2310 3232 2311 3236
rect 2315 3232 2316 3236
rect 2310 3231 2316 3232
rect 2438 3236 2444 3237
rect 2438 3232 2439 3236
rect 2443 3232 2444 3236
rect 2438 3231 2444 3232
rect 2582 3236 2588 3237
rect 2582 3232 2583 3236
rect 2587 3232 2588 3236
rect 2582 3231 2588 3232
rect 2734 3236 2740 3237
rect 2734 3232 2735 3236
rect 2739 3232 2740 3236
rect 2734 3231 2740 3232
rect 2910 3236 2916 3237
rect 2910 3232 2911 3236
rect 2915 3232 2916 3236
rect 2910 3231 2916 3232
rect 3102 3236 3108 3237
rect 3102 3232 3103 3236
rect 3107 3232 3108 3236
rect 3102 3231 3108 3232
rect 3302 3236 3308 3237
rect 3302 3232 3303 3236
rect 3307 3232 3308 3236
rect 3302 3231 3308 3232
rect 3502 3236 3508 3237
rect 3502 3232 3503 3236
rect 3507 3232 3508 3236
rect 3590 3235 3591 3239
rect 3595 3235 3596 3239
rect 3590 3234 3596 3235
rect 3502 3231 3508 3232
rect 134 3224 140 3225
rect 110 3221 116 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 134 3220 135 3224
rect 139 3220 140 3224
rect 134 3219 140 3220
rect 270 3224 276 3225
rect 270 3220 271 3224
rect 275 3220 276 3224
rect 270 3219 276 3220
rect 414 3224 420 3225
rect 414 3220 415 3224
rect 419 3220 420 3224
rect 414 3219 420 3220
rect 574 3224 580 3225
rect 574 3220 575 3224
rect 579 3220 580 3224
rect 574 3219 580 3220
rect 734 3224 740 3225
rect 734 3220 735 3224
rect 739 3220 740 3224
rect 734 3219 740 3220
rect 894 3224 900 3225
rect 894 3220 895 3224
rect 899 3220 900 3224
rect 894 3219 900 3220
rect 1046 3224 1052 3225
rect 1046 3220 1047 3224
rect 1051 3220 1052 3224
rect 1046 3219 1052 3220
rect 1190 3224 1196 3225
rect 1190 3220 1191 3224
rect 1195 3220 1196 3224
rect 1190 3219 1196 3220
rect 1326 3224 1332 3225
rect 1326 3220 1327 3224
rect 1331 3220 1332 3224
rect 1326 3219 1332 3220
rect 1462 3224 1468 3225
rect 1462 3220 1463 3224
rect 1467 3220 1468 3224
rect 1462 3219 1468 3220
rect 1606 3224 1612 3225
rect 1606 3220 1607 3224
rect 1611 3220 1612 3224
rect 1606 3219 1612 3220
rect 1830 3221 1836 3222
rect 110 3216 116 3217
rect 1830 3217 1831 3221
rect 1835 3217 1836 3221
rect 1830 3216 1836 3217
rect 2326 3219 2333 3220
rect 202 3215 208 3216
rect 202 3214 203 3215
rect 197 3212 203 3214
rect 202 3211 203 3212
rect 207 3211 208 3215
rect 351 3215 357 3216
rect 351 3214 352 3215
rect 333 3212 352 3214
rect 202 3210 208 3211
rect 351 3211 352 3212
rect 356 3211 357 3215
rect 546 3215 552 3216
rect 351 3210 357 3211
rect 194 3207 200 3208
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 194 3203 195 3207
rect 199 3206 200 3207
rect 432 3206 434 3213
rect 546 3211 547 3215
rect 551 3214 552 3215
rect 642 3215 648 3216
rect 551 3212 593 3214
rect 551 3211 552 3212
rect 546 3210 552 3211
rect 642 3211 643 3215
rect 647 3214 648 3215
rect 802 3215 808 3216
rect 647 3212 753 3214
rect 647 3211 648 3212
rect 642 3210 648 3211
rect 802 3211 803 3215
rect 807 3214 808 3215
rect 1114 3215 1120 3216
rect 1114 3214 1115 3215
rect 807 3212 913 3214
rect 1109 3212 1115 3214
rect 807 3211 808 3212
rect 802 3210 808 3211
rect 1114 3211 1115 3212
rect 1119 3211 1120 3215
rect 1282 3215 1288 3216
rect 1282 3214 1283 3215
rect 1253 3212 1283 3214
rect 1114 3210 1120 3211
rect 1282 3211 1283 3212
rect 1287 3211 1288 3215
rect 1418 3215 1424 3216
rect 1418 3214 1419 3215
rect 1389 3212 1419 3214
rect 1282 3210 1288 3211
rect 1418 3211 1419 3212
rect 1423 3211 1424 3215
rect 1558 3215 1564 3216
rect 1558 3214 1559 3215
rect 1525 3212 1559 3214
rect 1418 3210 1424 3211
rect 1558 3211 1559 3212
rect 1563 3211 1564 3215
rect 1558 3210 1564 3211
rect 1586 3215 1592 3216
rect 1586 3211 1587 3215
rect 1591 3214 1592 3215
rect 2326 3215 2327 3219
rect 2332 3215 2333 3219
rect 2326 3214 2333 3215
rect 1591 3212 1625 3214
rect 1591 3211 1592 3212
rect 1586 3210 1592 3211
rect 199 3204 434 3206
rect 1830 3204 1836 3205
rect 199 3203 200 3204
rect 194 3202 200 3203
rect 110 3199 116 3200
rect 1830 3200 1831 3204
rect 1835 3200 1836 3204
rect 1830 3199 1836 3200
rect 1894 3192 1900 3193
rect 1870 3189 1876 3190
rect 142 3186 148 3187
rect 142 3182 143 3186
rect 147 3182 148 3186
rect 142 3181 148 3182
rect 278 3186 284 3187
rect 278 3182 279 3186
rect 283 3182 284 3186
rect 278 3181 284 3182
rect 422 3186 428 3187
rect 422 3182 423 3186
rect 427 3182 428 3186
rect 422 3181 428 3182
rect 582 3186 588 3187
rect 582 3182 583 3186
rect 587 3182 588 3186
rect 582 3181 588 3182
rect 742 3186 748 3187
rect 742 3182 743 3186
rect 747 3182 748 3186
rect 742 3181 748 3182
rect 902 3186 908 3187
rect 902 3182 903 3186
rect 907 3182 908 3186
rect 902 3181 908 3182
rect 1054 3186 1060 3187
rect 1054 3182 1055 3186
rect 1059 3182 1060 3186
rect 1054 3181 1060 3182
rect 1198 3186 1204 3187
rect 1198 3182 1199 3186
rect 1203 3182 1204 3186
rect 1198 3181 1204 3182
rect 1334 3186 1340 3187
rect 1334 3182 1335 3186
rect 1339 3182 1340 3186
rect 1334 3181 1340 3182
rect 1470 3186 1476 3187
rect 1470 3182 1471 3186
rect 1475 3182 1476 3186
rect 1470 3181 1476 3182
rect 1614 3186 1620 3187
rect 1614 3182 1615 3186
rect 1619 3182 1620 3186
rect 1870 3185 1871 3189
rect 1875 3185 1876 3189
rect 1894 3188 1895 3192
rect 1899 3188 1900 3192
rect 1894 3187 1900 3188
rect 2006 3192 2012 3193
rect 2006 3188 2007 3192
rect 2011 3188 2012 3192
rect 2006 3187 2012 3188
rect 2142 3192 2148 3193
rect 2142 3188 2143 3192
rect 2147 3188 2148 3192
rect 2142 3187 2148 3188
rect 2294 3192 2300 3193
rect 2294 3188 2295 3192
rect 2299 3188 2300 3192
rect 2294 3187 2300 3188
rect 2454 3192 2460 3193
rect 2454 3188 2455 3192
rect 2459 3188 2460 3192
rect 2454 3187 2460 3188
rect 2622 3192 2628 3193
rect 2622 3188 2623 3192
rect 2627 3188 2628 3192
rect 2622 3187 2628 3188
rect 2798 3192 2804 3193
rect 2798 3188 2799 3192
rect 2803 3188 2804 3192
rect 2798 3187 2804 3188
rect 2974 3192 2980 3193
rect 2974 3188 2975 3192
rect 2979 3188 2980 3192
rect 2974 3187 2980 3188
rect 3150 3192 3156 3193
rect 3150 3188 3151 3192
rect 3155 3188 3156 3192
rect 3150 3187 3156 3188
rect 3326 3192 3332 3193
rect 3326 3188 3327 3192
rect 3331 3188 3332 3192
rect 3326 3187 3332 3188
rect 3502 3192 3508 3193
rect 3502 3188 3503 3192
rect 3507 3188 3508 3192
rect 3502 3187 3508 3188
rect 3590 3189 3596 3190
rect 1870 3184 1876 3185
rect 3590 3185 3591 3189
rect 3595 3185 3596 3189
rect 3590 3184 3596 3185
rect 1962 3183 1968 3184
rect 1962 3182 1963 3183
rect 1614 3181 1620 3182
rect 1957 3180 1963 3182
rect 1962 3179 1963 3180
rect 1967 3179 1968 3183
rect 2090 3183 2096 3184
rect 2090 3182 2091 3183
rect 2069 3180 2091 3182
rect 1962 3178 1968 3179
rect 2090 3179 2091 3180
rect 2095 3179 2096 3183
rect 2210 3183 2216 3184
rect 2210 3182 2211 3183
rect 2205 3180 2211 3182
rect 2090 3178 2096 3179
rect 2210 3179 2211 3180
rect 2215 3179 2216 3183
rect 2370 3183 2376 3184
rect 2370 3182 2371 3183
rect 2357 3180 2371 3182
rect 2210 3178 2216 3179
rect 2370 3179 2371 3180
rect 2375 3179 2376 3183
rect 2614 3183 2620 3184
rect 2464 3180 2473 3182
rect 2370 3178 2376 3179
rect 2462 3179 2468 3180
rect 167 3175 173 3176
rect 167 3171 168 3175
rect 172 3174 173 3175
rect 194 3175 200 3176
rect 194 3174 195 3175
rect 172 3172 195 3174
rect 172 3171 173 3172
rect 167 3170 173 3171
rect 194 3171 195 3172
rect 199 3171 200 3175
rect 194 3170 200 3171
rect 258 3175 264 3176
rect 258 3171 259 3175
rect 263 3174 264 3175
rect 303 3175 309 3176
rect 303 3174 304 3175
rect 263 3172 304 3174
rect 263 3171 264 3172
rect 258 3170 264 3171
rect 303 3171 304 3172
rect 308 3171 309 3175
rect 303 3170 309 3171
rect 351 3175 357 3176
rect 351 3171 352 3175
rect 356 3174 357 3175
rect 447 3175 453 3176
rect 447 3174 448 3175
rect 356 3172 448 3174
rect 356 3171 357 3172
rect 351 3170 357 3171
rect 447 3171 448 3172
rect 452 3171 453 3175
rect 447 3170 453 3171
rect 607 3175 613 3176
rect 607 3171 608 3175
rect 612 3174 613 3175
rect 642 3175 648 3176
rect 642 3174 643 3175
rect 612 3172 643 3174
rect 612 3171 613 3172
rect 607 3170 613 3171
rect 642 3171 643 3172
rect 647 3171 648 3175
rect 642 3170 648 3171
rect 767 3175 773 3176
rect 767 3171 768 3175
rect 772 3174 773 3175
rect 802 3175 808 3176
rect 802 3174 803 3175
rect 772 3172 803 3174
rect 772 3171 773 3172
rect 767 3170 773 3171
rect 802 3171 803 3172
rect 807 3171 808 3175
rect 802 3170 808 3171
rect 847 3175 853 3176
rect 847 3171 848 3175
rect 852 3174 853 3175
rect 927 3175 933 3176
rect 927 3174 928 3175
rect 852 3172 928 3174
rect 852 3171 853 3172
rect 847 3170 853 3171
rect 927 3171 928 3172
rect 932 3171 933 3175
rect 927 3170 933 3171
rect 1078 3175 1085 3176
rect 1078 3171 1079 3175
rect 1084 3171 1085 3175
rect 1078 3170 1085 3171
rect 1114 3175 1120 3176
rect 1114 3171 1115 3175
rect 1119 3174 1120 3175
rect 1223 3175 1229 3176
rect 1223 3174 1224 3175
rect 1119 3172 1224 3174
rect 1119 3171 1120 3172
rect 1114 3170 1120 3171
rect 1223 3171 1224 3172
rect 1228 3171 1229 3175
rect 1223 3170 1229 3171
rect 1282 3175 1288 3176
rect 1282 3171 1283 3175
rect 1287 3174 1288 3175
rect 1359 3175 1365 3176
rect 1359 3174 1360 3175
rect 1287 3172 1360 3174
rect 1287 3171 1288 3172
rect 1282 3170 1288 3171
rect 1359 3171 1360 3172
rect 1364 3171 1365 3175
rect 1359 3170 1365 3171
rect 1418 3175 1424 3176
rect 1418 3171 1419 3175
rect 1423 3174 1424 3175
rect 1495 3175 1501 3176
rect 1495 3174 1496 3175
rect 1423 3172 1496 3174
rect 1423 3171 1424 3172
rect 1418 3170 1424 3171
rect 1495 3171 1496 3172
rect 1500 3171 1501 3175
rect 1495 3170 1501 3171
rect 1558 3175 1564 3176
rect 1558 3171 1559 3175
rect 1563 3174 1564 3175
rect 1639 3175 1645 3176
rect 1639 3174 1640 3175
rect 1563 3172 1640 3174
rect 1563 3171 1564 3172
rect 1558 3170 1564 3171
rect 1639 3171 1640 3172
rect 1644 3171 1645 3175
rect 2462 3175 2463 3179
rect 2467 3175 2468 3179
rect 2614 3179 2615 3183
rect 2619 3182 2620 3183
rect 2690 3183 2696 3184
rect 2619 3180 2641 3182
rect 2619 3179 2620 3180
rect 2614 3178 2620 3179
rect 2690 3179 2691 3183
rect 2695 3182 2696 3183
rect 2914 3183 2920 3184
rect 2695 3180 2817 3182
rect 2695 3179 2696 3180
rect 2690 3178 2696 3179
rect 2914 3179 2915 3183
rect 2919 3182 2920 3183
rect 3262 3183 3268 3184
rect 3262 3182 3263 3183
rect 2919 3180 2993 3182
rect 3213 3180 3263 3182
rect 2919 3179 2920 3180
rect 2914 3178 2920 3179
rect 3262 3179 3263 3180
rect 3267 3179 3268 3183
rect 3398 3183 3404 3184
rect 3398 3182 3399 3183
rect 3389 3180 3399 3182
rect 3262 3178 3268 3179
rect 3398 3179 3399 3180
rect 3403 3179 3404 3183
rect 3398 3178 3404 3179
rect 2462 3174 2468 3175
rect 3210 3175 3216 3176
rect 1639 3170 1645 3171
rect 1870 3172 1876 3173
rect 1870 3168 1871 3172
rect 1875 3168 1876 3172
rect 3210 3171 3211 3175
rect 3215 3174 3216 3175
rect 3520 3174 3522 3181
rect 3215 3172 3522 3174
rect 3590 3172 3596 3173
rect 3215 3171 3216 3172
rect 3210 3170 3216 3171
rect 1870 3167 1876 3168
rect 3590 3168 3591 3172
rect 3595 3168 3596 3172
rect 3590 3167 3596 3168
rect 199 3155 208 3156
rect 199 3151 200 3155
rect 207 3151 208 3155
rect 199 3150 208 3151
rect 226 3155 232 3156
rect 226 3151 227 3155
rect 231 3154 232 3155
rect 343 3155 349 3156
rect 343 3154 344 3155
rect 231 3152 344 3154
rect 231 3151 232 3152
rect 226 3150 232 3151
rect 343 3151 344 3152
rect 348 3151 349 3155
rect 343 3150 349 3151
rect 487 3155 493 3156
rect 487 3151 488 3155
rect 492 3154 493 3155
rect 498 3155 504 3156
rect 498 3154 499 3155
rect 492 3152 499 3154
rect 492 3151 493 3152
rect 487 3150 493 3151
rect 498 3151 499 3152
rect 503 3151 504 3155
rect 498 3150 504 3151
rect 514 3155 520 3156
rect 514 3151 515 3155
rect 519 3154 520 3155
rect 631 3155 637 3156
rect 631 3154 632 3155
rect 519 3152 632 3154
rect 519 3151 520 3152
rect 514 3150 520 3151
rect 631 3151 632 3152
rect 636 3151 637 3155
rect 631 3150 637 3151
rect 658 3155 664 3156
rect 658 3151 659 3155
rect 663 3154 664 3155
rect 767 3155 773 3156
rect 767 3154 768 3155
rect 663 3152 768 3154
rect 663 3151 664 3152
rect 658 3150 664 3151
rect 767 3151 768 3152
rect 772 3151 773 3155
rect 767 3150 773 3151
rect 895 3155 901 3156
rect 895 3151 896 3155
rect 900 3154 901 3155
rect 910 3155 916 3156
rect 910 3154 911 3155
rect 900 3152 911 3154
rect 900 3151 901 3152
rect 895 3150 901 3151
rect 910 3151 911 3152
rect 915 3151 916 3155
rect 910 3150 916 3151
rect 922 3155 928 3156
rect 922 3151 923 3155
rect 927 3154 928 3155
rect 1015 3155 1021 3156
rect 1015 3154 1016 3155
rect 927 3152 1016 3154
rect 927 3151 928 3152
rect 922 3150 928 3151
rect 1015 3151 1016 3152
rect 1020 3151 1021 3155
rect 1015 3150 1021 3151
rect 1042 3155 1048 3156
rect 1042 3151 1043 3155
rect 1047 3154 1048 3155
rect 1127 3155 1133 3156
rect 1127 3154 1128 3155
rect 1047 3152 1128 3154
rect 1047 3151 1048 3152
rect 1042 3150 1048 3151
rect 1127 3151 1128 3152
rect 1132 3151 1133 3155
rect 1127 3150 1133 3151
rect 1154 3155 1160 3156
rect 1154 3151 1155 3155
rect 1159 3154 1160 3155
rect 1231 3155 1237 3156
rect 1231 3154 1232 3155
rect 1159 3152 1232 3154
rect 1159 3151 1160 3152
rect 1154 3150 1160 3151
rect 1231 3151 1232 3152
rect 1236 3151 1237 3155
rect 1231 3150 1237 3151
rect 1258 3155 1264 3156
rect 1258 3151 1259 3155
rect 1263 3154 1264 3155
rect 1335 3155 1341 3156
rect 1335 3154 1336 3155
rect 1263 3152 1336 3154
rect 1263 3151 1264 3152
rect 1258 3150 1264 3151
rect 1335 3151 1336 3152
rect 1340 3151 1341 3155
rect 1335 3150 1341 3151
rect 1362 3155 1368 3156
rect 1362 3151 1363 3155
rect 1367 3154 1368 3155
rect 1431 3155 1437 3156
rect 1431 3154 1432 3155
rect 1367 3152 1432 3154
rect 1367 3151 1368 3152
rect 1362 3150 1368 3151
rect 1431 3151 1432 3152
rect 1436 3151 1437 3155
rect 1431 3150 1437 3151
rect 1458 3155 1464 3156
rect 1458 3151 1459 3155
rect 1463 3154 1464 3155
rect 1519 3155 1525 3156
rect 1519 3154 1520 3155
rect 1463 3152 1520 3154
rect 1463 3151 1464 3152
rect 1458 3150 1464 3151
rect 1519 3151 1520 3152
rect 1524 3151 1525 3155
rect 1519 3150 1525 3151
rect 1546 3155 1552 3156
rect 1546 3151 1547 3155
rect 1551 3154 1552 3155
rect 1607 3155 1613 3156
rect 1607 3154 1608 3155
rect 1551 3152 1608 3154
rect 1551 3151 1552 3152
rect 1546 3150 1552 3151
rect 1607 3151 1608 3152
rect 1612 3151 1613 3155
rect 1607 3150 1613 3151
rect 1634 3155 1640 3156
rect 1634 3151 1635 3155
rect 1639 3154 1640 3155
rect 1695 3155 1701 3156
rect 1695 3154 1696 3155
rect 1639 3152 1696 3154
rect 1639 3151 1640 3152
rect 1634 3150 1640 3151
rect 1695 3151 1696 3152
rect 1700 3151 1701 3155
rect 1695 3150 1701 3151
rect 1722 3155 1728 3156
rect 1722 3151 1723 3155
rect 1727 3154 1728 3155
rect 1775 3155 1781 3156
rect 1775 3154 1776 3155
rect 1727 3152 1776 3154
rect 1727 3151 1728 3152
rect 1722 3150 1728 3151
rect 1775 3151 1776 3152
rect 1780 3151 1781 3155
rect 1775 3150 1781 3151
rect 1902 3154 1908 3155
rect 1902 3150 1903 3154
rect 1907 3150 1908 3154
rect 1902 3149 1908 3150
rect 2014 3154 2020 3155
rect 2014 3150 2015 3154
rect 2019 3150 2020 3154
rect 2014 3149 2020 3150
rect 2150 3154 2156 3155
rect 2150 3150 2151 3154
rect 2155 3150 2156 3154
rect 2150 3149 2156 3150
rect 2302 3154 2308 3155
rect 2302 3150 2303 3154
rect 2307 3150 2308 3154
rect 2302 3149 2308 3150
rect 2462 3154 2468 3155
rect 2462 3150 2463 3154
rect 2467 3150 2468 3154
rect 2462 3149 2468 3150
rect 2630 3154 2636 3155
rect 2630 3150 2631 3154
rect 2635 3150 2636 3154
rect 2630 3149 2636 3150
rect 2806 3154 2812 3155
rect 2806 3150 2807 3154
rect 2811 3150 2812 3154
rect 2806 3149 2812 3150
rect 2982 3154 2988 3155
rect 2982 3150 2983 3154
rect 2987 3150 2988 3154
rect 2982 3149 2988 3150
rect 3158 3154 3164 3155
rect 3158 3150 3159 3154
rect 3163 3150 3164 3154
rect 3158 3149 3164 3150
rect 3334 3154 3340 3155
rect 3334 3150 3335 3154
rect 3339 3150 3340 3154
rect 3334 3149 3340 3150
rect 3510 3154 3516 3155
rect 3510 3150 3511 3154
rect 3515 3150 3516 3154
rect 3510 3149 3516 3150
rect 174 3146 180 3147
rect 174 3142 175 3146
rect 179 3142 180 3146
rect 174 3141 180 3142
rect 318 3146 324 3147
rect 318 3142 319 3146
rect 323 3142 324 3146
rect 318 3141 324 3142
rect 462 3146 468 3147
rect 462 3142 463 3146
rect 467 3142 468 3146
rect 462 3141 468 3142
rect 606 3146 612 3147
rect 606 3142 607 3146
rect 611 3142 612 3146
rect 606 3141 612 3142
rect 742 3146 748 3147
rect 742 3142 743 3146
rect 747 3142 748 3146
rect 742 3141 748 3142
rect 870 3146 876 3147
rect 870 3142 871 3146
rect 875 3142 876 3146
rect 870 3141 876 3142
rect 990 3146 996 3147
rect 990 3142 991 3146
rect 995 3142 996 3146
rect 990 3141 996 3142
rect 1102 3146 1108 3147
rect 1102 3142 1103 3146
rect 1107 3142 1108 3146
rect 1102 3141 1108 3142
rect 1206 3146 1212 3147
rect 1206 3142 1207 3146
rect 1211 3142 1212 3146
rect 1206 3141 1212 3142
rect 1310 3146 1316 3147
rect 1310 3142 1311 3146
rect 1315 3142 1316 3146
rect 1310 3141 1316 3142
rect 1406 3146 1412 3147
rect 1406 3142 1407 3146
rect 1411 3142 1412 3146
rect 1406 3141 1412 3142
rect 1494 3146 1500 3147
rect 1494 3142 1495 3146
rect 1499 3142 1500 3146
rect 1494 3141 1500 3142
rect 1582 3146 1588 3147
rect 1582 3142 1583 3146
rect 1587 3142 1588 3146
rect 1582 3141 1588 3142
rect 1670 3146 1676 3147
rect 1670 3142 1671 3146
rect 1675 3142 1676 3146
rect 1670 3141 1676 3142
rect 1750 3146 1756 3147
rect 1750 3142 1751 3146
rect 1755 3142 1756 3146
rect 1750 3141 1756 3142
rect 1926 3143 1933 3144
rect 1926 3139 1927 3143
rect 1932 3139 1933 3143
rect 1926 3138 1933 3139
rect 1962 3143 1968 3144
rect 1962 3139 1963 3143
rect 1967 3142 1968 3143
rect 2039 3143 2045 3144
rect 2039 3142 2040 3143
rect 1967 3140 2040 3142
rect 1967 3139 1968 3140
rect 1962 3138 1968 3139
rect 2039 3139 2040 3140
rect 2044 3139 2045 3143
rect 2039 3138 2045 3139
rect 2090 3143 2096 3144
rect 2090 3139 2091 3143
rect 2095 3142 2096 3143
rect 2175 3143 2181 3144
rect 2175 3142 2176 3143
rect 2095 3140 2176 3142
rect 2095 3139 2096 3140
rect 2090 3138 2096 3139
rect 2175 3139 2176 3140
rect 2180 3139 2181 3143
rect 2175 3138 2181 3139
rect 2326 3143 2333 3144
rect 2326 3139 2327 3143
rect 2332 3139 2333 3143
rect 2326 3138 2333 3139
rect 2370 3143 2376 3144
rect 2370 3139 2371 3143
rect 2375 3142 2376 3143
rect 2487 3143 2493 3144
rect 2487 3142 2488 3143
rect 2375 3140 2488 3142
rect 2375 3139 2376 3140
rect 2370 3138 2376 3139
rect 2487 3139 2488 3140
rect 2492 3139 2493 3143
rect 2487 3138 2493 3139
rect 2655 3143 2661 3144
rect 2655 3139 2656 3143
rect 2660 3142 2661 3143
rect 2690 3143 2696 3144
rect 2690 3142 2691 3143
rect 2660 3140 2691 3142
rect 2660 3139 2661 3140
rect 2655 3138 2661 3139
rect 2690 3139 2691 3140
rect 2695 3139 2696 3143
rect 2690 3138 2696 3139
rect 2831 3143 2837 3144
rect 2831 3139 2832 3143
rect 2836 3142 2837 3143
rect 2914 3143 2920 3144
rect 2914 3142 2915 3143
rect 2836 3140 2915 3142
rect 2836 3139 2837 3140
rect 2831 3138 2837 3139
rect 2914 3139 2915 3140
rect 2919 3139 2920 3143
rect 2914 3138 2920 3139
rect 3006 3143 3013 3144
rect 3006 3139 3007 3143
rect 3012 3139 3013 3143
rect 3006 3138 3013 3139
rect 3183 3143 3189 3144
rect 3183 3139 3184 3143
rect 3188 3142 3189 3143
rect 3210 3143 3216 3144
rect 3210 3142 3211 3143
rect 3188 3140 3211 3142
rect 3188 3139 3189 3140
rect 3183 3138 3189 3139
rect 3210 3139 3211 3140
rect 3215 3139 3216 3143
rect 3210 3138 3216 3139
rect 3262 3143 3268 3144
rect 3262 3139 3263 3143
rect 3267 3142 3268 3143
rect 3359 3143 3365 3144
rect 3359 3142 3360 3143
rect 3267 3140 3360 3142
rect 3267 3139 3268 3140
rect 3262 3138 3268 3139
rect 3359 3139 3360 3140
rect 3364 3139 3365 3143
rect 3359 3138 3365 3139
rect 3534 3143 3541 3144
rect 3534 3139 3535 3143
rect 3540 3139 3541 3143
rect 3534 3138 3541 3139
rect 1927 3131 1933 3132
rect 1927 3130 1928 3131
rect 110 3128 116 3129
rect 110 3124 111 3128
rect 115 3124 116 3128
rect 110 3123 116 3124
rect 1830 3128 1836 3129
rect 1830 3124 1831 3128
rect 1835 3124 1836 3128
rect 1830 3123 1836 3124
rect 1844 3128 1928 3130
rect 226 3119 232 3120
rect 226 3115 227 3119
rect 231 3115 232 3119
rect 226 3114 232 3115
rect 358 3119 364 3120
rect 358 3115 359 3119
rect 363 3115 364 3119
rect 358 3114 364 3115
rect 514 3119 520 3120
rect 514 3115 515 3119
rect 519 3115 520 3119
rect 514 3114 520 3115
rect 658 3119 664 3120
rect 658 3115 659 3119
rect 663 3115 664 3119
rect 847 3119 853 3120
rect 847 3118 848 3119
rect 797 3116 848 3118
rect 658 3114 664 3115
rect 847 3115 848 3116
rect 852 3115 853 3119
rect 847 3114 853 3115
rect 922 3119 928 3120
rect 922 3115 923 3119
rect 927 3115 928 3119
rect 922 3114 928 3115
rect 1042 3119 1048 3120
rect 1042 3115 1043 3119
rect 1047 3115 1048 3119
rect 1042 3114 1048 3115
rect 1154 3119 1160 3120
rect 1154 3115 1155 3119
rect 1159 3115 1160 3119
rect 1154 3114 1160 3115
rect 1258 3119 1264 3120
rect 1258 3115 1259 3119
rect 1263 3115 1264 3119
rect 1258 3114 1264 3115
rect 1362 3119 1368 3120
rect 1362 3115 1363 3119
rect 1367 3115 1368 3119
rect 1362 3114 1368 3115
rect 1458 3119 1464 3120
rect 1458 3115 1459 3119
rect 1463 3115 1464 3119
rect 1458 3114 1464 3115
rect 1546 3119 1552 3120
rect 1546 3115 1547 3119
rect 1551 3115 1552 3119
rect 1546 3114 1552 3115
rect 1634 3119 1640 3120
rect 1634 3115 1635 3119
rect 1639 3115 1640 3119
rect 1634 3114 1640 3115
rect 1722 3119 1728 3120
rect 1722 3115 1723 3119
rect 1727 3115 1728 3119
rect 1844 3118 1846 3128
rect 1927 3127 1928 3128
rect 1932 3127 1933 3131
rect 1927 3126 1933 3127
rect 2095 3131 2101 3132
rect 2095 3127 2096 3131
rect 2100 3130 2101 3131
rect 2114 3131 2120 3132
rect 2114 3130 2115 3131
rect 2100 3128 2115 3130
rect 2100 3127 2101 3128
rect 2095 3126 2101 3127
rect 2114 3127 2115 3128
rect 2119 3127 2120 3131
rect 2114 3126 2120 3127
rect 2122 3131 2128 3132
rect 2122 3127 2123 3131
rect 2127 3130 2128 3131
rect 2287 3131 2293 3132
rect 2287 3130 2288 3131
rect 2127 3128 2288 3130
rect 2127 3127 2128 3128
rect 2122 3126 2128 3127
rect 2287 3127 2288 3128
rect 2292 3127 2293 3131
rect 2287 3126 2293 3127
rect 2470 3131 2476 3132
rect 2470 3127 2471 3131
rect 2475 3130 2476 3131
rect 2479 3131 2485 3132
rect 2479 3130 2480 3131
rect 2475 3128 2480 3130
rect 2475 3127 2476 3128
rect 2470 3126 2476 3127
rect 2479 3127 2480 3128
rect 2484 3127 2485 3131
rect 2479 3126 2485 3127
rect 2671 3131 2677 3132
rect 2671 3127 2672 3131
rect 2676 3130 2677 3131
rect 2682 3131 2688 3132
rect 2682 3130 2683 3131
rect 2676 3128 2683 3130
rect 2676 3127 2677 3128
rect 2671 3126 2677 3127
rect 2682 3127 2683 3128
rect 2687 3127 2688 3131
rect 2682 3126 2688 3127
rect 2698 3131 2704 3132
rect 2698 3127 2699 3131
rect 2703 3130 2704 3131
rect 2855 3131 2861 3132
rect 2855 3130 2856 3131
rect 2703 3128 2856 3130
rect 2703 3127 2704 3128
rect 2698 3126 2704 3127
rect 2855 3127 2856 3128
rect 2860 3127 2861 3131
rect 2855 3126 2861 3127
rect 3039 3131 3048 3132
rect 3039 3127 3040 3131
rect 3047 3127 3048 3131
rect 3039 3126 3048 3127
rect 3066 3131 3072 3132
rect 3066 3127 3067 3131
rect 3071 3130 3072 3131
rect 3223 3131 3229 3132
rect 3223 3130 3224 3131
rect 3071 3128 3224 3130
rect 3071 3127 3072 3128
rect 3066 3126 3072 3127
rect 3223 3127 3224 3128
rect 3228 3127 3229 3131
rect 3223 3126 3229 3127
rect 3398 3131 3404 3132
rect 3398 3127 3399 3131
rect 3403 3130 3404 3131
rect 3415 3131 3421 3132
rect 3415 3130 3416 3131
rect 3403 3128 3416 3130
rect 3403 3127 3404 3128
rect 3398 3126 3404 3127
rect 3415 3127 3416 3128
rect 3420 3127 3421 3131
rect 3415 3126 3421 3127
rect 1805 3116 1846 3118
rect 1902 3122 1908 3123
rect 1902 3118 1903 3122
rect 1907 3118 1908 3122
rect 1902 3117 1908 3118
rect 2070 3122 2076 3123
rect 2070 3118 2071 3122
rect 2075 3118 2076 3122
rect 2070 3117 2076 3118
rect 2262 3122 2268 3123
rect 2262 3118 2263 3122
rect 2267 3118 2268 3122
rect 2262 3117 2268 3118
rect 2454 3122 2460 3123
rect 2454 3118 2455 3122
rect 2459 3118 2460 3122
rect 2454 3117 2460 3118
rect 2646 3122 2652 3123
rect 2646 3118 2647 3122
rect 2651 3118 2652 3122
rect 2646 3117 2652 3118
rect 2830 3122 2836 3123
rect 2830 3118 2831 3122
rect 2835 3118 2836 3122
rect 2830 3117 2836 3118
rect 3014 3122 3020 3123
rect 3014 3118 3015 3122
rect 3019 3118 3020 3122
rect 3014 3117 3020 3118
rect 3198 3122 3204 3123
rect 3198 3118 3199 3122
rect 3203 3118 3204 3122
rect 3198 3117 3204 3118
rect 3390 3122 3396 3123
rect 3390 3118 3391 3122
rect 3395 3118 3396 3122
rect 3390 3117 3396 3118
rect 1722 3114 1728 3115
rect 110 3111 116 3112
rect 110 3107 111 3111
rect 115 3107 116 3111
rect 1830 3111 1836 3112
rect 110 3106 116 3107
rect 166 3108 172 3109
rect 166 3104 167 3108
rect 171 3104 172 3108
rect 166 3103 172 3104
rect 310 3108 316 3109
rect 310 3104 311 3108
rect 315 3104 316 3108
rect 310 3103 316 3104
rect 454 3108 460 3109
rect 454 3104 455 3108
rect 459 3104 460 3108
rect 454 3103 460 3104
rect 598 3108 604 3109
rect 598 3104 599 3108
rect 603 3104 604 3108
rect 598 3103 604 3104
rect 734 3108 740 3109
rect 734 3104 735 3108
rect 739 3104 740 3108
rect 734 3103 740 3104
rect 862 3108 868 3109
rect 862 3104 863 3108
rect 867 3104 868 3108
rect 862 3103 868 3104
rect 982 3108 988 3109
rect 982 3104 983 3108
rect 987 3104 988 3108
rect 982 3103 988 3104
rect 1094 3108 1100 3109
rect 1094 3104 1095 3108
rect 1099 3104 1100 3108
rect 1094 3103 1100 3104
rect 1198 3108 1204 3109
rect 1198 3104 1199 3108
rect 1203 3104 1204 3108
rect 1198 3103 1204 3104
rect 1302 3108 1308 3109
rect 1302 3104 1303 3108
rect 1307 3104 1308 3108
rect 1302 3103 1308 3104
rect 1398 3108 1404 3109
rect 1398 3104 1399 3108
rect 1403 3104 1404 3108
rect 1398 3103 1404 3104
rect 1486 3108 1492 3109
rect 1486 3104 1487 3108
rect 1491 3104 1492 3108
rect 1486 3103 1492 3104
rect 1574 3108 1580 3109
rect 1574 3104 1575 3108
rect 1579 3104 1580 3108
rect 1574 3103 1580 3104
rect 1662 3108 1668 3109
rect 1662 3104 1663 3108
rect 1667 3104 1668 3108
rect 1662 3103 1668 3104
rect 1742 3108 1748 3109
rect 1742 3104 1743 3108
rect 1747 3104 1748 3108
rect 1830 3107 1831 3111
rect 1835 3107 1836 3111
rect 1830 3106 1836 3107
rect 1742 3103 1748 3104
rect 1870 3104 1876 3105
rect 1870 3100 1871 3104
rect 1875 3100 1876 3104
rect 1870 3099 1876 3100
rect 3590 3104 3596 3105
rect 3590 3100 3591 3104
rect 3595 3100 3596 3104
rect 3590 3099 3596 3100
rect 1926 3095 1932 3096
rect 1926 3091 1927 3095
rect 1931 3091 1932 3095
rect 1926 3090 1932 3091
rect 2122 3095 2128 3096
rect 2122 3091 2123 3095
rect 2127 3091 2128 3095
rect 2122 3090 2128 3091
rect 2314 3095 2320 3096
rect 2314 3091 2315 3095
rect 2319 3091 2320 3095
rect 2314 3090 2320 3091
rect 2698 3095 2704 3096
rect 2698 3091 2699 3095
rect 2703 3091 2704 3095
rect 3006 3095 3012 3096
rect 3006 3094 3007 3095
rect 2885 3092 3007 3094
rect 2698 3090 2704 3091
rect 3006 3091 3007 3092
rect 3011 3091 3012 3095
rect 3006 3090 3012 3091
rect 3066 3095 3072 3096
rect 3066 3091 3067 3095
rect 3071 3091 3072 3095
rect 3282 3095 3288 3096
rect 3282 3094 3283 3095
rect 3253 3092 3283 3094
rect 3066 3090 3072 3091
rect 3282 3091 3283 3092
rect 3287 3091 3288 3095
rect 3282 3090 3288 3091
rect 1870 3087 1876 3088
rect 1870 3083 1871 3087
rect 1875 3083 1876 3087
rect 3590 3087 3596 3088
rect 1870 3082 1876 3083
rect 1894 3084 1900 3085
rect 1894 3080 1895 3084
rect 1899 3080 1900 3084
rect 1894 3079 1900 3080
rect 2062 3084 2068 3085
rect 2062 3080 2063 3084
rect 2067 3080 2068 3084
rect 2062 3079 2068 3080
rect 2254 3084 2260 3085
rect 2254 3080 2255 3084
rect 2259 3080 2260 3084
rect 2254 3079 2260 3080
rect 2446 3084 2452 3085
rect 2446 3080 2447 3084
rect 2451 3080 2452 3084
rect 2446 3079 2452 3080
rect 2638 3084 2644 3085
rect 2638 3080 2639 3084
rect 2643 3080 2644 3084
rect 2638 3079 2644 3080
rect 2822 3084 2828 3085
rect 2822 3080 2823 3084
rect 2827 3080 2828 3084
rect 2822 3079 2828 3080
rect 3006 3084 3012 3085
rect 3006 3080 3007 3084
rect 3011 3080 3012 3084
rect 3006 3079 3012 3080
rect 3190 3084 3196 3085
rect 3190 3080 3191 3084
rect 3195 3080 3196 3084
rect 3190 3079 3196 3080
rect 3382 3084 3388 3085
rect 3382 3080 3383 3084
rect 3387 3080 3388 3084
rect 3590 3083 3591 3087
rect 3595 3083 3596 3087
rect 3590 3082 3596 3083
rect 3382 3079 3388 3080
rect 2114 3067 2120 3068
rect 2114 3063 2115 3067
rect 2119 3066 2120 3067
rect 2463 3067 2469 3068
rect 2463 3066 2464 3067
rect 2119 3064 2464 3066
rect 2119 3063 2120 3064
rect 2114 3062 2120 3063
rect 2463 3063 2464 3064
rect 2468 3063 2469 3067
rect 2463 3062 2469 3063
rect 3042 3067 3048 3068
rect 3042 3063 3043 3067
rect 3047 3066 3048 3067
rect 3399 3067 3405 3068
rect 3399 3066 3400 3067
rect 3047 3064 3400 3066
rect 3047 3063 3048 3064
rect 3042 3062 3048 3063
rect 3399 3063 3400 3064
rect 3404 3063 3405 3067
rect 3399 3062 3405 3063
rect 134 3052 140 3053
rect 110 3049 116 3050
rect 110 3045 111 3049
rect 115 3045 116 3049
rect 134 3048 135 3052
rect 139 3048 140 3052
rect 134 3047 140 3048
rect 222 3052 228 3053
rect 222 3048 223 3052
rect 227 3048 228 3052
rect 222 3047 228 3048
rect 326 3052 332 3053
rect 326 3048 327 3052
rect 331 3048 332 3052
rect 326 3047 332 3048
rect 438 3052 444 3053
rect 438 3048 439 3052
rect 443 3048 444 3052
rect 438 3047 444 3048
rect 550 3052 556 3053
rect 550 3048 551 3052
rect 555 3048 556 3052
rect 550 3047 556 3048
rect 662 3052 668 3053
rect 662 3048 663 3052
rect 667 3048 668 3052
rect 662 3047 668 3048
rect 1830 3049 1836 3050
rect 110 3044 116 3045
rect 1830 3045 1831 3049
rect 1835 3045 1836 3049
rect 1830 3044 1836 3045
rect 202 3043 208 3044
rect 196 3036 198 3041
rect 202 3039 203 3043
rect 207 3042 208 3043
rect 290 3043 296 3044
rect 207 3040 241 3042
rect 207 3039 208 3040
rect 202 3038 208 3039
rect 290 3039 291 3043
rect 295 3042 296 3043
rect 506 3043 512 3044
rect 295 3040 345 3042
rect 295 3039 296 3040
rect 290 3038 296 3039
rect 500 3036 502 3041
rect 506 3039 507 3043
rect 511 3042 512 3043
rect 618 3043 624 3044
rect 511 3040 569 3042
rect 511 3039 512 3040
rect 506 3038 512 3039
rect 618 3039 619 3043
rect 623 3042 624 3043
rect 623 3040 681 3042
rect 623 3039 624 3040
rect 618 3038 624 3039
rect 194 3035 200 3036
rect 110 3032 116 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 194 3031 195 3035
rect 199 3031 200 3035
rect 194 3030 200 3031
rect 498 3035 504 3036
rect 498 3031 499 3035
rect 503 3031 504 3035
rect 498 3030 504 3031
rect 1830 3032 1836 3033
rect 110 3027 116 3028
rect 1830 3028 1831 3032
rect 1835 3028 1836 3032
rect 1830 3027 1836 3028
rect 2198 3028 2204 3029
rect 1870 3025 1876 3026
rect 1870 3021 1871 3025
rect 1875 3021 1876 3025
rect 2198 3024 2199 3028
rect 2203 3024 2204 3028
rect 2198 3023 2204 3024
rect 2334 3028 2340 3029
rect 2334 3024 2335 3028
rect 2339 3024 2340 3028
rect 2334 3023 2340 3024
rect 2478 3028 2484 3029
rect 2478 3024 2479 3028
rect 2483 3024 2484 3028
rect 2478 3023 2484 3024
rect 2622 3028 2628 3029
rect 2622 3024 2623 3028
rect 2627 3024 2628 3028
rect 2622 3023 2628 3024
rect 2766 3028 2772 3029
rect 2766 3024 2767 3028
rect 2771 3024 2772 3028
rect 2766 3023 2772 3024
rect 2902 3028 2908 3029
rect 2902 3024 2903 3028
rect 2907 3024 2908 3028
rect 2902 3023 2908 3024
rect 3038 3028 3044 3029
rect 3038 3024 3039 3028
rect 3043 3024 3044 3028
rect 3038 3023 3044 3024
rect 3182 3028 3188 3029
rect 3182 3024 3183 3028
rect 3187 3024 3188 3028
rect 3182 3023 3188 3024
rect 3326 3028 3332 3029
rect 3326 3024 3327 3028
rect 3331 3024 3332 3028
rect 3326 3023 3332 3024
rect 3590 3025 3596 3026
rect 1870 3020 1876 3021
rect 3590 3021 3591 3025
rect 3595 3021 3596 3025
rect 3590 3020 3596 3021
rect 2426 3019 2432 3020
rect 2426 3018 2427 3019
rect 142 3014 148 3015
rect 142 3010 143 3014
rect 147 3010 148 3014
rect 142 3009 148 3010
rect 230 3014 236 3015
rect 230 3010 231 3014
rect 235 3010 236 3014
rect 230 3009 236 3010
rect 334 3014 340 3015
rect 334 3010 335 3014
rect 339 3010 340 3014
rect 334 3009 340 3010
rect 446 3014 452 3015
rect 446 3010 447 3014
rect 451 3010 452 3014
rect 446 3009 452 3010
rect 558 3014 564 3015
rect 558 3010 559 3014
rect 563 3010 564 3014
rect 558 3009 564 3010
rect 670 3014 676 3015
rect 670 3010 671 3014
rect 675 3010 676 3014
rect 2260 3012 2262 3017
rect 2397 3016 2427 3018
rect 2426 3015 2427 3016
rect 2431 3015 2432 3019
rect 2690 3019 2696 3020
rect 2426 3014 2432 3015
rect 670 3009 676 3010
rect 2258 3011 2264 3012
rect 1870 3008 1876 3009
rect 1870 3004 1871 3008
rect 1875 3004 1876 3008
rect 2258 3007 2259 3011
rect 2263 3007 2264 3011
rect 2258 3006 2264 3007
rect 2266 3011 2272 3012
rect 2266 3007 2267 3011
rect 2271 3010 2272 3011
rect 2496 3010 2498 3017
rect 2684 3012 2686 3017
rect 2690 3015 2691 3019
rect 2695 3018 2696 3019
rect 2834 3019 2840 3020
rect 2695 3016 2785 3018
rect 2695 3015 2696 3016
rect 2690 3014 2696 3015
rect 2834 3015 2835 3019
rect 2839 3018 2840 3019
rect 3106 3019 3112 3020
rect 2839 3016 2921 3018
rect 2839 3015 2840 3016
rect 2834 3014 2840 3015
rect 3100 3012 3102 3017
rect 3106 3015 3107 3019
rect 3111 3018 3112 3019
rect 3250 3019 3256 3020
rect 3111 3016 3201 3018
rect 3111 3015 3112 3016
rect 3106 3014 3112 3015
rect 3250 3015 3251 3019
rect 3255 3018 3256 3019
rect 3255 3016 3345 3018
rect 3255 3015 3256 3016
rect 3250 3014 3256 3015
rect 2271 3008 2498 3010
rect 2682 3011 2688 3012
rect 2271 3007 2272 3008
rect 2266 3006 2272 3007
rect 2682 3007 2683 3011
rect 2687 3007 2688 3011
rect 2682 3006 2688 3007
rect 3098 3011 3104 3012
rect 3098 3007 3099 3011
rect 3103 3007 3104 3011
rect 3098 3006 3104 3007
rect 3590 3008 3596 3009
rect 167 3003 173 3004
rect 167 2999 168 3003
rect 172 3002 173 3003
rect 202 3003 208 3004
rect 202 3002 203 3003
rect 172 3000 203 3002
rect 172 2999 173 3000
rect 167 2998 173 2999
rect 202 2999 203 3000
rect 207 2999 208 3003
rect 202 2998 208 2999
rect 255 3003 261 3004
rect 255 2999 256 3003
rect 260 3002 261 3003
rect 290 3003 296 3004
rect 290 3002 291 3003
rect 260 3000 291 3002
rect 260 2999 261 3000
rect 255 2998 261 2999
rect 290 2999 291 3000
rect 295 2999 296 3003
rect 290 2998 296 2999
rect 358 3003 365 3004
rect 358 2999 359 3003
rect 364 2999 365 3003
rect 358 2998 365 2999
rect 471 3003 477 3004
rect 471 2999 472 3003
rect 476 3002 477 3003
rect 506 3003 512 3004
rect 506 3002 507 3003
rect 476 3000 507 3002
rect 476 2999 477 3000
rect 471 2998 477 2999
rect 506 2999 507 3000
rect 511 2999 512 3003
rect 506 2998 512 2999
rect 583 3003 589 3004
rect 583 2999 584 3003
rect 588 3002 589 3003
rect 618 3003 624 3004
rect 618 3002 619 3003
rect 588 3000 619 3002
rect 588 2999 589 3000
rect 583 2998 589 2999
rect 618 2999 619 3000
rect 623 2999 624 3003
rect 618 2998 624 2999
rect 695 3003 701 3004
rect 695 2999 696 3003
rect 700 3002 701 3003
rect 806 3003 812 3004
rect 1870 3003 1876 3004
rect 3590 3004 3591 3008
rect 3595 3004 3596 3008
rect 3590 3003 3596 3004
rect 806 3002 807 3003
rect 700 3000 807 3002
rect 700 2999 701 3000
rect 695 2998 701 2999
rect 806 2999 807 3000
rect 811 2999 812 3003
rect 806 2998 812 2999
rect 2206 2990 2212 2991
rect 1262 2987 1268 2988
rect 1262 2986 1263 2987
rect 1064 2984 1263 2986
rect 183 2979 189 2980
rect 183 2975 184 2979
rect 188 2978 189 2979
rect 194 2979 200 2980
rect 194 2978 195 2979
rect 188 2976 195 2978
rect 188 2975 189 2976
rect 183 2974 189 2975
rect 194 2975 195 2976
rect 199 2975 200 2979
rect 194 2974 200 2975
rect 210 2979 216 2980
rect 210 2975 211 2979
rect 215 2978 216 2979
rect 343 2979 349 2980
rect 343 2978 344 2979
rect 215 2976 344 2978
rect 215 2975 216 2976
rect 210 2974 216 2975
rect 343 2975 344 2976
rect 348 2975 349 2979
rect 343 2974 349 2975
rect 511 2979 517 2980
rect 511 2975 512 2979
rect 516 2978 517 2979
rect 530 2979 536 2980
rect 530 2978 531 2979
rect 516 2976 531 2978
rect 516 2975 517 2976
rect 511 2974 517 2975
rect 530 2975 531 2976
rect 535 2975 536 2979
rect 530 2974 536 2975
rect 538 2979 544 2980
rect 538 2975 539 2979
rect 543 2978 544 2979
rect 671 2979 677 2980
rect 671 2978 672 2979
rect 543 2976 672 2978
rect 543 2975 544 2976
rect 538 2974 544 2975
rect 671 2975 672 2976
rect 676 2975 677 2979
rect 671 2974 677 2975
rect 698 2979 704 2980
rect 698 2975 699 2979
rect 703 2978 704 2979
rect 823 2979 829 2980
rect 823 2978 824 2979
rect 703 2976 824 2978
rect 703 2975 704 2976
rect 698 2974 704 2975
rect 823 2975 824 2976
rect 828 2975 829 2979
rect 823 2974 829 2975
rect 967 2979 973 2980
rect 967 2975 968 2979
rect 972 2978 973 2979
rect 1064 2978 1066 2984
rect 1262 2983 1263 2984
rect 1267 2983 1268 2987
rect 2206 2986 2207 2990
rect 2211 2986 2212 2990
rect 2206 2985 2212 2986
rect 2342 2990 2348 2991
rect 2342 2986 2343 2990
rect 2347 2986 2348 2990
rect 2342 2985 2348 2986
rect 2486 2990 2492 2991
rect 2486 2986 2487 2990
rect 2491 2986 2492 2990
rect 2486 2985 2492 2986
rect 2630 2990 2636 2991
rect 2630 2986 2631 2990
rect 2635 2986 2636 2990
rect 2630 2985 2636 2986
rect 2774 2990 2780 2991
rect 2774 2986 2775 2990
rect 2779 2986 2780 2990
rect 2774 2985 2780 2986
rect 2910 2990 2916 2991
rect 2910 2986 2911 2990
rect 2915 2986 2916 2990
rect 2910 2985 2916 2986
rect 3046 2990 3052 2991
rect 3046 2986 3047 2990
rect 3051 2986 3052 2990
rect 3046 2985 3052 2986
rect 3190 2990 3196 2991
rect 3190 2986 3191 2990
rect 3195 2986 3196 2990
rect 3190 2985 3196 2986
rect 3334 2990 3340 2991
rect 3334 2986 3335 2990
rect 3339 2986 3340 2990
rect 3334 2985 3340 2986
rect 1262 2982 1268 2983
rect 972 2976 1066 2978
rect 1070 2979 1076 2980
rect 972 2975 973 2976
rect 967 2974 973 2975
rect 1070 2975 1071 2979
rect 1075 2978 1076 2979
rect 1103 2979 1109 2980
rect 1103 2978 1104 2979
rect 1075 2976 1104 2978
rect 1075 2975 1076 2976
rect 1070 2974 1076 2975
rect 1103 2975 1104 2976
rect 1108 2975 1109 2979
rect 1103 2974 1109 2975
rect 1130 2979 1136 2980
rect 1130 2975 1131 2979
rect 1135 2978 1136 2979
rect 1223 2979 1229 2980
rect 1223 2978 1224 2979
rect 1135 2976 1224 2978
rect 1135 2975 1136 2976
rect 1130 2974 1136 2975
rect 1223 2975 1224 2976
rect 1228 2975 1229 2979
rect 1223 2974 1229 2975
rect 1250 2979 1256 2980
rect 1250 2975 1251 2979
rect 1255 2978 1256 2979
rect 1335 2979 1341 2980
rect 1335 2978 1336 2979
rect 1255 2976 1336 2978
rect 1255 2975 1256 2976
rect 1250 2974 1256 2975
rect 1335 2975 1336 2976
rect 1340 2975 1341 2979
rect 1335 2974 1341 2975
rect 1362 2979 1368 2980
rect 1362 2975 1363 2979
rect 1367 2978 1368 2979
rect 1447 2979 1453 2980
rect 1447 2978 1448 2979
rect 1367 2976 1448 2978
rect 1367 2975 1368 2976
rect 1362 2974 1368 2975
rect 1447 2975 1448 2976
rect 1452 2975 1453 2979
rect 1447 2974 1453 2975
rect 1474 2979 1480 2980
rect 1474 2975 1475 2979
rect 1479 2978 1480 2979
rect 1559 2979 1565 2980
rect 1559 2978 1560 2979
rect 1479 2976 1560 2978
rect 1479 2975 1480 2976
rect 1474 2974 1480 2975
rect 1559 2975 1560 2976
rect 1564 2975 1565 2979
rect 1559 2974 1565 2975
rect 1586 2979 1592 2980
rect 1586 2975 1587 2979
rect 1591 2978 1592 2979
rect 1671 2979 1677 2980
rect 1671 2978 1672 2979
rect 1591 2976 1672 2978
rect 1591 2975 1592 2976
rect 1586 2974 1592 2975
rect 1671 2975 1672 2976
rect 1676 2975 1677 2979
rect 1671 2974 1677 2975
rect 2231 2979 2237 2980
rect 2231 2975 2232 2979
rect 2236 2978 2237 2979
rect 2266 2979 2272 2980
rect 2266 2978 2267 2979
rect 2236 2976 2267 2978
rect 2236 2975 2237 2976
rect 2231 2974 2237 2975
rect 2266 2975 2267 2976
rect 2271 2975 2272 2979
rect 2266 2974 2272 2975
rect 2314 2979 2320 2980
rect 2314 2975 2315 2979
rect 2319 2978 2320 2979
rect 2367 2979 2373 2980
rect 2367 2978 2368 2979
rect 2319 2976 2368 2978
rect 2319 2975 2320 2976
rect 2314 2974 2320 2975
rect 2367 2975 2368 2976
rect 2372 2975 2373 2979
rect 2367 2974 2373 2975
rect 2426 2979 2432 2980
rect 2426 2975 2427 2979
rect 2431 2978 2432 2979
rect 2511 2979 2517 2980
rect 2511 2978 2512 2979
rect 2431 2976 2512 2978
rect 2431 2975 2432 2976
rect 2426 2974 2432 2975
rect 2511 2975 2512 2976
rect 2516 2975 2517 2979
rect 2511 2974 2517 2975
rect 2655 2979 2661 2980
rect 2655 2975 2656 2979
rect 2660 2978 2661 2979
rect 2690 2979 2696 2980
rect 2690 2978 2691 2979
rect 2660 2976 2691 2978
rect 2660 2975 2661 2976
rect 2655 2974 2661 2975
rect 2690 2975 2691 2976
rect 2695 2975 2696 2979
rect 2690 2974 2696 2975
rect 2799 2979 2805 2980
rect 2799 2975 2800 2979
rect 2804 2978 2805 2979
rect 2834 2979 2840 2980
rect 2834 2978 2835 2979
rect 2804 2976 2835 2978
rect 2804 2975 2805 2976
rect 2799 2974 2805 2975
rect 2834 2975 2835 2976
rect 2839 2975 2840 2979
rect 2834 2974 2840 2975
rect 2935 2979 2941 2980
rect 2935 2975 2936 2979
rect 2940 2978 2941 2979
rect 2983 2979 2989 2980
rect 2983 2978 2984 2979
rect 2940 2976 2984 2978
rect 2940 2975 2941 2976
rect 2935 2974 2941 2975
rect 2983 2975 2984 2976
rect 2988 2975 2989 2979
rect 2983 2974 2989 2975
rect 3071 2979 3077 2980
rect 3071 2975 3072 2979
rect 3076 2978 3077 2979
rect 3106 2979 3112 2980
rect 3106 2978 3107 2979
rect 3076 2976 3107 2978
rect 3076 2975 3077 2976
rect 3071 2974 3077 2975
rect 3106 2975 3107 2976
rect 3111 2975 3112 2979
rect 3106 2974 3112 2975
rect 3215 2979 3221 2980
rect 3215 2975 3216 2979
rect 3220 2978 3221 2979
rect 3250 2979 3256 2980
rect 3250 2978 3251 2979
rect 3220 2976 3251 2978
rect 3220 2975 3221 2976
rect 3215 2974 3221 2975
rect 3250 2975 3251 2976
rect 3255 2975 3256 2979
rect 3250 2974 3256 2975
rect 3282 2979 3288 2980
rect 3282 2975 3283 2979
rect 3287 2978 3288 2979
rect 3359 2979 3365 2980
rect 3359 2978 3360 2979
rect 3287 2976 3360 2978
rect 3287 2975 3288 2976
rect 3282 2974 3288 2975
rect 3359 2975 3360 2976
rect 3364 2975 3365 2979
rect 3359 2974 3365 2975
rect 158 2970 164 2971
rect 158 2966 159 2970
rect 163 2966 164 2970
rect 158 2965 164 2966
rect 318 2970 324 2971
rect 318 2966 319 2970
rect 323 2966 324 2970
rect 318 2965 324 2966
rect 486 2970 492 2971
rect 486 2966 487 2970
rect 491 2966 492 2970
rect 486 2965 492 2966
rect 646 2970 652 2971
rect 646 2966 647 2970
rect 651 2966 652 2970
rect 646 2965 652 2966
rect 798 2970 804 2971
rect 798 2966 799 2970
rect 803 2966 804 2970
rect 798 2965 804 2966
rect 942 2970 948 2971
rect 942 2966 943 2970
rect 947 2966 948 2970
rect 942 2965 948 2966
rect 1078 2970 1084 2971
rect 1078 2966 1079 2970
rect 1083 2966 1084 2970
rect 1078 2965 1084 2966
rect 1198 2970 1204 2971
rect 1198 2966 1199 2970
rect 1203 2966 1204 2970
rect 1198 2965 1204 2966
rect 1310 2970 1316 2971
rect 1310 2966 1311 2970
rect 1315 2966 1316 2970
rect 1310 2965 1316 2966
rect 1422 2970 1428 2971
rect 1422 2966 1423 2970
rect 1427 2966 1428 2970
rect 1422 2965 1428 2966
rect 1534 2970 1540 2971
rect 1534 2966 1535 2970
rect 1539 2966 1540 2970
rect 1534 2965 1540 2966
rect 1646 2970 1652 2971
rect 1646 2966 1647 2970
rect 1651 2966 1652 2970
rect 1646 2965 1652 2966
rect 2151 2955 2157 2956
rect 110 2952 116 2953
rect 110 2948 111 2952
rect 115 2948 116 2952
rect 110 2947 116 2948
rect 1830 2952 1836 2953
rect 1830 2948 1831 2952
rect 1835 2948 1836 2952
rect 2151 2951 2152 2955
rect 2156 2954 2157 2955
rect 2214 2955 2220 2956
rect 2214 2954 2215 2955
rect 2156 2952 2215 2954
rect 2156 2951 2157 2952
rect 2151 2950 2157 2951
rect 2214 2951 2215 2952
rect 2219 2951 2220 2955
rect 2214 2950 2220 2951
rect 2231 2955 2237 2956
rect 2231 2951 2232 2955
rect 2236 2954 2237 2955
rect 2258 2955 2264 2956
rect 2258 2954 2259 2955
rect 2236 2952 2259 2954
rect 2236 2951 2237 2952
rect 2231 2950 2237 2951
rect 2258 2951 2259 2952
rect 2263 2951 2264 2955
rect 2258 2950 2264 2951
rect 2311 2955 2320 2956
rect 2311 2951 2312 2955
rect 2319 2951 2320 2955
rect 2311 2950 2320 2951
rect 2350 2955 2356 2956
rect 2350 2951 2351 2955
rect 2355 2954 2356 2955
rect 2391 2955 2397 2956
rect 2391 2954 2392 2955
rect 2355 2952 2392 2954
rect 2355 2951 2356 2952
rect 2350 2950 2356 2951
rect 2391 2951 2392 2952
rect 2396 2951 2397 2955
rect 2391 2950 2397 2951
rect 2418 2955 2424 2956
rect 2418 2951 2419 2955
rect 2423 2954 2424 2955
rect 2471 2955 2477 2956
rect 2471 2954 2472 2955
rect 2423 2952 2472 2954
rect 2423 2951 2424 2952
rect 2418 2950 2424 2951
rect 2471 2951 2472 2952
rect 2476 2951 2477 2955
rect 2471 2950 2477 2951
rect 2498 2955 2504 2956
rect 2498 2951 2499 2955
rect 2503 2954 2504 2955
rect 2551 2955 2557 2956
rect 2551 2954 2552 2955
rect 2503 2952 2552 2954
rect 2503 2951 2504 2952
rect 2498 2950 2504 2951
rect 2551 2951 2552 2952
rect 2556 2951 2557 2955
rect 2551 2950 2557 2951
rect 2578 2955 2584 2956
rect 2578 2951 2579 2955
rect 2583 2954 2584 2955
rect 2631 2955 2637 2956
rect 2631 2954 2632 2955
rect 2583 2952 2632 2954
rect 2583 2951 2584 2952
rect 2578 2950 2584 2951
rect 2631 2951 2632 2952
rect 2636 2951 2637 2955
rect 2631 2950 2637 2951
rect 2658 2955 2664 2956
rect 2658 2951 2659 2955
rect 2663 2954 2664 2955
rect 2719 2955 2725 2956
rect 2719 2954 2720 2955
rect 2663 2952 2720 2954
rect 2663 2951 2664 2952
rect 2658 2950 2664 2951
rect 2719 2951 2720 2952
rect 2724 2951 2725 2955
rect 2719 2950 2725 2951
rect 2746 2955 2752 2956
rect 2746 2951 2747 2955
rect 2751 2954 2752 2955
rect 2815 2955 2821 2956
rect 2815 2954 2816 2955
rect 2751 2952 2816 2954
rect 2751 2951 2752 2952
rect 2746 2950 2752 2951
rect 2815 2951 2816 2952
rect 2820 2951 2821 2955
rect 2815 2950 2821 2951
rect 2935 2955 2941 2956
rect 2935 2951 2936 2955
rect 2940 2954 2941 2955
rect 2946 2955 2952 2956
rect 2946 2954 2947 2955
rect 2940 2952 2947 2954
rect 2940 2951 2941 2952
rect 2935 2950 2941 2951
rect 2946 2951 2947 2952
rect 2951 2951 2952 2955
rect 2946 2950 2952 2951
rect 2962 2955 2968 2956
rect 2962 2951 2963 2955
rect 2967 2954 2968 2955
rect 3063 2955 3069 2956
rect 3063 2954 3064 2955
rect 2967 2952 3064 2954
rect 2967 2951 2968 2952
rect 2962 2950 2968 2951
rect 3063 2951 3064 2952
rect 3068 2951 3069 2955
rect 3063 2950 3069 2951
rect 3098 2955 3104 2956
rect 3098 2951 3099 2955
rect 3103 2954 3104 2955
rect 3207 2955 3213 2956
rect 3207 2954 3208 2955
rect 3103 2952 3208 2954
rect 3103 2951 3104 2952
rect 3098 2950 3104 2951
rect 3207 2951 3208 2952
rect 3212 2951 3213 2955
rect 3207 2950 3213 2951
rect 3234 2955 3240 2956
rect 3234 2951 3235 2955
rect 3239 2954 3240 2955
rect 3359 2955 3365 2956
rect 3359 2954 3360 2955
rect 3239 2952 3360 2954
rect 3239 2951 3240 2952
rect 3234 2950 3240 2951
rect 3359 2951 3360 2952
rect 3364 2951 3365 2955
rect 3359 2950 3365 2951
rect 3438 2955 3444 2956
rect 3438 2951 3439 2955
rect 3443 2954 3444 2955
rect 3519 2955 3525 2956
rect 3519 2954 3520 2955
rect 3443 2952 3520 2954
rect 3443 2951 3444 2952
rect 3438 2950 3444 2951
rect 3519 2951 3520 2952
rect 3524 2951 3525 2955
rect 3519 2950 3525 2951
rect 1830 2947 1836 2948
rect 2126 2946 2132 2947
rect 210 2943 216 2944
rect 210 2939 211 2943
rect 215 2939 216 2943
rect 210 2938 216 2939
rect 342 2943 348 2944
rect 342 2939 343 2943
rect 347 2939 348 2943
rect 342 2938 348 2939
rect 538 2943 544 2944
rect 538 2939 539 2943
rect 543 2939 544 2943
rect 538 2938 544 2939
rect 698 2943 704 2944
rect 698 2939 699 2943
rect 703 2939 704 2943
rect 698 2938 704 2939
rect 806 2943 812 2944
rect 806 2939 807 2943
rect 811 2939 812 2943
rect 1070 2943 1076 2944
rect 1070 2942 1071 2943
rect 997 2940 1071 2942
rect 806 2938 812 2939
rect 1070 2939 1071 2940
rect 1075 2939 1076 2943
rect 1070 2938 1076 2939
rect 1130 2943 1136 2944
rect 1130 2939 1131 2943
rect 1135 2939 1136 2943
rect 1130 2938 1136 2939
rect 1250 2943 1256 2944
rect 1250 2939 1251 2943
rect 1255 2939 1256 2943
rect 1250 2938 1256 2939
rect 1362 2943 1368 2944
rect 1362 2939 1363 2943
rect 1367 2939 1368 2943
rect 1362 2938 1368 2939
rect 1474 2943 1480 2944
rect 1474 2939 1475 2943
rect 1479 2939 1480 2943
rect 1474 2938 1480 2939
rect 1586 2943 1592 2944
rect 1586 2939 1587 2943
rect 1591 2939 1592 2943
rect 2126 2942 2127 2946
rect 2131 2942 2132 2946
rect 2126 2941 2132 2942
rect 2206 2946 2212 2947
rect 2206 2942 2207 2946
rect 2211 2942 2212 2946
rect 2206 2941 2212 2942
rect 2286 2946 2292 2947
rect 2286 2942 2287 2946
rect 2291 2942 2292 2946
rect 2286 2941 2292 2942
rect 2366 2946 2372 2947
rect 2366 2942 2367 2946
rect 2371 2942 2372 2946
rect 2366 2941 2372 2942
rect 2446 2946 2452 2947
rect 2446 2942 2447 2946
rect 2451 2942 2452 2946
rect 2446 2941 2452 2942
rect 2526 2946 2532 2947
rect 2526 2942 2527 2946
rect 2531 2942 2532 2946
rect 2526 2941 2532 2942
rect 2606 2946 2612 2947
rect 2606 2942 2607 2946
rect 2611 2942 2612 2946
rect 2606 2941 2612 2942
rect 2694 2946 2700 2947
rect 2694 2942 2695 2946
rect 2699 2942 2700 2946
rect 2694 2941 2700 2942
rect 2790 2946 2796 2947
rect 2790 2942 2791 2946
rect 2795 2942 2796 2946
rect 2790 2941 2796 2942
rect 2910 2946 2916 2947
rect 2910 2942 2911 2946
rect 2915 2942 2916 2946
rect 2910 2941 2916 2942
rect 3038 2946 3044 2947
rect 3038 2942 3039 2946
rect 3043 2942 3044 2946
rect 3038 2941 3044 2942
rect 3182 2946 3188 2947
rect 3182 2942 3183 2946
rect 3187 2942 3188 2946
rect 3182 2941 3188 2942
rect 3334 2946 3340 2947
rect 3334 2942 3335 2946
rect 3339 2942 3340 2946
rect 3334 2941 3340 2942
rect 3494 2946 3500 2947
rect 3494 2942 3495 2946
rect 3499 2942 3500 2946
rect 3494 2941 3500 2942
rect 1586 2938 1592 2939
rect 110 2935 116 2936
rect 110 2931 111 2935
rect 115 2931 116 2935
rect 1830 2935 1836 2936
rect 110 2930 116 2931
rect 150 2932 156 2933
rect 150 2928 151 2932
rect 155 2928 156 2932
rect 150 2927 156 2928
rect 310 2932 316 2933
rect 310 2928 311 2932
rect 315 2928 316 2932
rect 310 2927 316 2928
rect 478 2932 484 2933
rect 478 2928 479 2932
rect 483 2928 484 2932
rect 478 2927 484 2928
rect 638 2932 644 2933
rect 638 2928 639 2932
rect 643 2928 644 2932
rect 638 2927 644 2928
rect 790 2932 796 2933
rect 790 2928 791 2932
rect 795 2928 796 2932
rect 790 2927 796 2928
rect 934 2932 940 2933
rect 934 2928 935 2932
rect 939 2928 940 2932
rect 934 2927 940 2928
rect 1070 2932 1076 2933
rect 1070 2928 1071 2932
rect 1075 2928 1076 2932
rect 1070 2927 1076 2928
rect 1190 2932 1196 2933
rect 1190 2928 1191 2932
rect 1195 2928 1196 2932
rect 1190 2927 1196 2928
rect 1302 2932 1308 2933
rect 1302 2928 1303 2932
rect 1307 2928 1308 2932
rect 1302 2927 1308 2928
rect 1414 2932 1420 2933
rect 1414 2928 1415 2932
rect 1419 2928 1420 2932
rect 1414 2927 1420 2928
rect 1526 2932 1532 2933
rect 1526 2928 1527 2932
rect 1531 2928 1532 2932
rect 1526 2927 1532 2928
rect 1638 2932 1644 2933
rect 1638 2928 1639 2932
rect 1643 2928 1644 2932
rect 1830 2931 1831 2935
rect 1835 2931 1836 2935
rect 1830 2930 1836 2931
rect 1638 2927 1644 2928
rect 1870 2928 1876 2929
rect 1870 2924 1871 2928
rect 1875 2924 1876 2928
rect 1870 2923 1876 2924
rect 3590 2928 3596 2929
rect 3590 2924 3591 2928
rect 3595 2924 3596 2928
rect 3590 2923 3596 2924
rect 2214 2919 2220 2920
rect 1426 2915 1432 2916
rect 1426 2911 1427 2915
rect 1431 2914 1432 2915
rect 1655 2915 1661 2916
rect 1655 2914 1656 2915
rect 1431 2912 1656 2914
rect 1431 2911 1432 2912
rect 1426 2910 1432 2911
rect 1655 2911 1656 2912
rect 1660 2911 1661 2915
rect 2214 2915 2215 2919
rect 2219 2915 2220 2919
rect 2350 2919 2356 2920
rect 2350 2918 2351 2919
rect 2341 2916 2351 2918
rect 2214 2914 2220 2915
rect 2350 2915 2351 2916
rect 2355 2915 2356 2919
rect 2350 2914 2356 2915
rect 2418 2919 2424 2920
rect 2418 2915 2419 2919
rect 2423 2915 2424 2919
rect 2418 2914 2424 2915
rect 2498 2919 2504 2920
rect 2498 2915 2499 2919
rect 2503 2915 2504 2919
rect 2498 2914 2504 2915
rect 2578 2919 2584 2920
rect 2578 2915 2579 2919
rect 2583 2915 2584 2919
rect 2578 2914 2584 2915
rect 2658 2919 2664 2920
rect 2658 2915 2659 2919
rect 2663 2915 2664 2919
rect 2658 2914 2664 2915
rect 2746 2919 2752 2920
rect 2746 2915 2747 2919
rect 2751 2915 2752 2919
rect 2746 2914 2752 2915
rect 2962 2919 2968 2920
rect 2962 2915 2963 2919
rect 2967 2915 2968 2919
rect 2962 2914 2968 2915
rect 2983 2919 2989 2920
rect 2983 2915 2984 2919
rect 2988 2918 2989 2919
rect 3234 2919 3240 2920
rect 2988 2916 3049 2918
rect 2988 2915 2989 2916
rect 2983 2914 2989 2915
rect 3234 2915 3235 2919
rect 3239 2915 3240 2919
rect 3234 2914 3240 2915
rect 3534 2919 3540 2920
rect 3534 2915 3535 2919
rect 3539 2915 3540 2919
rect 3534 2914 3540 2915
rect 1655 2910 1661 2911
rect 1870 2911 1876 2912
rect 1870 2907 1871 2911
rect 1875 2907 1876 2911
rect 3590 2911 3596 2912
rect 1870 2906 1876 2907
rect 2118 2908 2124 2909
rect 2118 2904 2119 2908
rect 2123 2904 2124 2908
rect 2118 2903 2124 2904
rect 2198 2908 2204 2909
rect 2198 2904 2199 2908
rect 2203 2904 2204 2908
rect 2198 2903 2204 2904
rect 2278 2908 2284 2909
rect 2278 2904 2279 2908
rect 2283 2904 2284 2908
rect 2278 2903 2284 2904
rect 2358 2908 2364 2909
rect 2358 2904 2359 2908
rect 2363 2904 2364 2908
rect 2358 2903 2364 2904
rect 2438 2908 2444 2909
rect 2438 2904 2439 2908
rect 2443 2904 2444 2908
rect 2438 2903 2444 2904
rect 2518 2908 2524 2909
rect 2518 2904 2519 2908
rect 2523 2904 2524 2908
rect 2518 2903 2524 2904
rect 2598 2908 2604 2909
rect 2598 2904 2599 2908
rect 2603 2904 2604 2908
rect 2598 2903 2604 2904
rect 2686 2908 2692 2909
rect 2686 2904 2687 2908
rect 2691 2904 2692 2908
rect 2686 2903 2692 2904
rect 2782 2908 2788 2909
rect 2782 2904 2783 2908
rect 2787 2904 2788 2908
rect 2782 2903 2788 2904
rect 2902 2908 2908 2909
rect 2902 2904 2903 2908
rect 2907 2904 2908 2908
rect 2902 2903 2908 2904
rect 3030 2908 3036 2909
rect 3030 2904 3031 2908
rect 3035 2904 3036 2908
rect 3030 2903 3036 2904
rect 3174 2908 3180 2909
rect 3174 2904 3175 2908
rect 3179 2904 3180 2908
rect 3174 2903 3180 2904
rect 3326 2908 3332 2909
rect 3326 2904 3327 2908
rect 3331 2904 3332 2908
rect 3326 2903 3332 2904
rect 3486 2908 3492 2909
rect 3486 2904 3487 2908
rect 3491 2904 3492 2908
rect 3590 2907 3591 2911
rect 3595 2907 3596 2911
rect 3590 2906 3596 2907
rect 3486 2903 3492 2904
rect 2082 2891 2088 2892
rect 150 2888 156 2889
rect 110 2885 116 2886
rect 110 2881 111 2885
rect 115 2881 116 2885
rect 150 2884 151 2888
rect 155 2884 156 2888
rect 150 2883 156 2884
rect 310 2888 316 2889
rect 310 2884 311 2888
rect 315 2884 316 2888
rect 310 2883 316 2884
rect 470 2888 476 2889
rect 470 2884 471 2888
rect 475 2884 476 2888
rect 470 2883 476 2884
rect 630 2888 636 2889
rect 630 2884 631 2888
rect 635 2884 636 2888
rect 630 2883 636 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 926 2888 932 2889
rect 926 2884 927 2888
rect 931 2884 932 2888
rect 926 2883 932 2884
rect 1054 2888 1060 2889
rect 1054 2884 1055 2888
rect 1059 2884 1060 2888
rect 1054 2883 1060 2884
rect 1174 2888 1180 2889
rect 1174 2884 1175 2888
rect 1179 2884 1180 2888
rect 1174 2883 1180 2884
rect 1286 2888 1292 2889
rect 1286 2884 1287 2888
rect 1291 2884 1292 2888
rect 1286 2883 1292 2884
rect 1390 2888 1396 2889
rect 1390 2884 1391 2888
rect 1395 2884 1396 2888
rect 1390 2883 1396 2884
rect 1486 2888 1492 2889
rect 1486 2884 1487 2888
rect 1491 2884 1492 2888
rect 1486 2883 1492 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1590 2883 1596 2884
rect 1694 2888 1700 2889
rect 1694 2884 1695 2888
rect 1699 2884 1700 2888
rect 2082 2887 2083 2891
rect 2087 2890 2088 2891
rect 2135 2891 2141 2892
rect 2135 2890 2136 2891
rect 2087 2888 2136 2890
rect 2087 2887 2088 2888
rect 2082 2886 2088 2887
rect 2135 2887 2136 2888
rect 2140 2887 2141 2891
rect 2135 2886 2141 2887
rect 2626 2891 2632 2892
rect 2626 2887 2627 2891
rect 2631 2890 2632 2891
rect 2799 2891 2805 2892
rect 2799 2890 2800 2891
rect 2631 2888 2800 2890
rect 2631 2887 2632 2888
rect 2626 2886 2632 2887
rect 2799 2887 2800 2888
rect 2804 2887 2805 2891
rect 2799 2886 2805 2887
rect 3226 2891 3232 2892
rect 3226 2887 3227 2891
rect 3231 2890 3232 2891
rect 3343 2891 3349 2892
rect 3343 2890 3344 2891
rect 3231 2888 3344 2890
rect 3231 2887 3232 2888
rect 3226 2886 3232 2887
rect 3343 2887 3344 2888
rect 3348 2887 3349 2891
rect 3343 2886 3349 2887
rect 1694 2883 1700 2884
rect 1830 2885 1836 2886
rect 110 2880 116 2881
rect 1830 2881 1831 2885
rect 1835 2881 1836 2885
rect 1830 2880 1836 2881
rect 218 2879 224 2880
rect 152 2876 169 2878
rect 150 2875 156 2876
rect 150 2871 151 2875
rect 155 2871 156 2875
rect 218 2875 219 2879
rect 223 2878 224 2879
rect 538 2879 544 2880
rect 223 2876 329 2878
rect 223 2875 224 2876
rect 218 2874 224 2875
rect 532 2872 534 2877
rect 538 2875 539 2879
rect 543 2878 544 2879
rect 698 2879 704 2880
rect 543 2876 649 2878
rect 543 2875 544 2876
rect 538 2874 544 2875
rect 698 2875 699 2879
rect 703 2878 704 2879
rect 1014 2879 1020 2880
rect 1014 2878 1015 2879
rect 703 2876 801 2878
rect 989 2876 1015 2878
rect 703 2875 704 2876
rect 698 2874 704 2875
rect 1014 2875 1015 2876
rect 1019 2875 1020 2879
rect 1122 2879 1128 2880
rect 1122 2878 1123 2879
rect 1117 2876 1123 2878
rect 1014 2874 1020 2875
rect 1122 2875 1123 2876
rect 1127 2875 1128 2879
rect 1254 2879 1260 2880
rect 1254 2878 1255 2879
rect 1237 2876 1255 2878
rect 1122 2874 1128 2875
rect 1254 2875 1255 2876
rect 1259 2875 1260 2879
rect 1254 2874 1260 2875
rect 1262 2879 1268 2880
rect 1262 2875 1263 2879
rect 1267 2878 1268 2879
rect 1462 2879 1468 2880
rect 1462 2878 1463 2879
rect 1267 2876 1305 2878
rect 1453 2876 1463 2878
rect 1267 2875 1268 2876
rect 1262 2874 1268 2875
rect 1462 2875 1463 2876
rect 1467 2875 1468 2879
rect 1562 2879 1568 2880
rect 1562 2878 1563 2879
rect 1549 2876 1563 2878
rect 1462 2874 1468 2875
rect 1562 2875 1563 2876
rect 1567 2875 1568 2879
rect 1666 2879 1672 2880
rect 1666 2878 1667 2879
rect 1653 2876 1667 2878
rect 1562 2874 1568 2875
rect 1666 2875 1667 2876
rect 1671 2875 1672 2879
rect 1666 2874 1672 2875
rect 1674 2879 1680 2880
rect 1674 2875 1675 2879
rect 1679 2878 1680 2879
rect 1679 2876 1713 2878
rect 1679 2875 1680 2876
rect 1674 2874 1680 2875
rect 150 2870 156 2871
rect 530 2871 536 2872
rect 110 2868 116 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 530 2867 531 2871
rect 535 2867 536 2871
rect 530 2866 536 2867
rect 1830 2868 1836 2869
rect 110 2863 116 2864
rect 1830 2864 1831 2868
rect 1835 2864 1836 2868
rect 1830 2863 1836 2864
rect 2046 2864 2052 2865
rect 1870 2861 1876 2862
rect 1870 2857 1871 2861
rect 1875 2857 1876 2861
rect 2046 2860 2047 2864
rect 2051 2860 2052 2864
rect 2046 2859 2052 2860
rect 2134 2864 2140 2865
rect 2134 2860 2135 2864
rect 2139 2860 2140 2864
rect 2134 2859 2140 2860
rect 2238 2864 2244 2865
rect 2238 2860 2239 2864
rect 2243 2860 2244 2864
rect 2238 2859 2244 2860
rect 2342 2864 2348 2865
rect 2342 2860 2343 2864
rect 2347 2860 2348 2864
rect 2342 2859 2348 2860
rect 2462 2864 2468 2865
rect 2462 2860 2463 2864
rect 2467 2860 2468 2864
rect 2462 2859 2468 2860
rect 2590 2864 2596 2865
rect 2590 2860 2591 2864
rect 2595 2860 2596 2864
rect 2590 2859 2596 2860
rect 2726 2864 2732 2865
rect 2726 2860 2727 2864
rect 2731 2860 2732 2864
rect 2726 2859 2732 2860
rect 2878 2864 2884 2865
rect 2878 2860 2879 2864
rect 2883 2860 2884 2864
rect 2878 2859 2884 2860
rect 3030 2864 3036 2865
rect 3030 2860 3031 2864
rect 3035 2860 3036 2864
rect 3030 2859 3036 2860
rect 3190 2864 3196 2865
rect 3190 2860 3191 2864
rect 3195 2860 3196 2864
rect 3190 2859 3196 2860
rect 3358 2864 3364 2865
rect 3358 2860 3359 2864
rect 3363 2860 3364 2864
rect 3358 2859 3364 2860
rect 3502 2864 3508 2865
rect 3502 2860 3503 2864
rect 3507 2860 3508 2864
rect 3502 2859 3508 2860
rect 3590 2861 3596 2862
rect 1870 2856 1876 2857
rect 3590 2857 3591 2861
rect 3595 2857 3596 2861
rect 3590 2856 3596 2857
rect 2114 2855 2120 2856
rect 2114 2854 2115 2855
rect 2109 2852 2115 2854
rect 2114 2851 2115 2852
rect 2119 2851 2120 2855
rect 2306 2855 2312 2856
rect 158 2850 164 2851
rect 158 2846 159 2850
rect 163 2846 164 2850
rect 158 2845 164 2846
rect 318 2850 324 2851
rect 318 2846 319 2850
rect 323 2846 324 2850
rect 318 2845 324 2846
rect 478 2850 484 2851
rect 478 2846 479 2850
rect 483 2846 484 2850
rect 478 2845 484 2846
rect 638 2850 644 2851
rect 638 2846 639 2850
rect 643 2846 644 2850
rect 638 2845 644 2846
rect 790 2850 796 2851
rect 790 2846 791 2850
rect 795 2846 796 2850
rect 790 2845 796 2846
rect 934 2850 940 2851
rect 934 2846 935 2850
rect 939 2846 940 2850
rect 934 2845 940 2846
rect 1062 2850 1068 2851
rect 1062 2846 1063 2850
rect 1067 2846 1068 2850
rect 1062 2845 1068 2846
rect 1182 2850 1188 2851
rect 1182 2846 1183 2850
rect 1187 2846 1188 2850
rect 1182 2845 1188 2846
rect 1294 2850 1300 2851
rect 1294 2846 1295 2850
rect 1299 2846 1300 2850
rect 1294 2845 1300 2846
rect 1398 2850 1404 2851
rect 1398 2846 1399 2850
rect 1403 2846 1404 2850
rect 1398 2845 1404 2846
rect 1494 2850 1500 2851
rect 1494 2846 1495 2850
rect 1499 2846 1500 2850
rect 1494 2845 1500 2846
rect 1598 2850 1604 2851
rect 1598 2846 1599 2850
rect 1603 2846 1604 2850
rect 1598 2845 1604 2846
rect 1702 2850 1708 2851
rect 2114 2850 2120 2851
rect 1702 2846 1703 2850
rect 1707 2846 1708 2850
rect 2196 2848 2198 2853
rect 1702 2845 1708 2846
rect 2194 2847 2200 2848
rect 1870 2844 1876 2845
rect 1870 2840 1871 2844
rect 1875 2840 1876 2844
rect 2194 2843 2195 2847
rect 2199 2843 2200 2847
rect 2300 2846 2302 2853
rect 2306 2851 2307 2855
rect 2311 2854 2312 2855
rect 2410 2855 2416 2856
rect 2311 2852 2361 2854
rect 2311 2851 2312 2852
rect 2306 2850 2312 2851
rect 2410 2851 2411 2855
rect 2415 2854 2416 2855
rect 2682 2855 2688 2856
rect 2682 2854 2683 2855
rect 2415 2852 2481 2854
rect 2653 2852 2683 2854
rect 2415 2851 2416 2852
rect 2410 2850 2416 2851
rect 2682 2851 2683 2852
rect 2687 2851 2688 2855
rect 2794 2855 2800 2856
rect 2794 2854 2795 2855
rect 2789 2852 2795 2854
rect 2682 2850 2688 2851
rect 2794 2851 2795 2852
rect 2799 2851 2800 2855
rect 2946 2855 2952 2856
rect 2946 2854 2947 2855
rect 2941 2852 2947 2854
rect 2794 2850 2800 2851
rect 2946 2851 2947 2852
rect 2951 2851 2952 2855
rect 2946 2850 2952 2851
rect 2958 2855 2964 2856
rect 2958 2851 2959 2855
rect 2963 2854 2964 2855
rect 3098 2855 3104 2856
rect 2963 2852 3049 2854
rect 2963 2851 2964 2852
rect 2958 2850 2964 2851
rect 3098 2851 3099 2855
rect 3103 2854 3104 2855
rect 3438 2855 3444 2856
rect 3438 2854 3439 2855
rect 3103 2852 3209 2854
rect 3421 2852 3439 2854
rect 3103 2851 3104 2852
rect 3098 2850 3104 2851
rect 3438 2851 3439 2852
rect 3443 2851 3444 2855
rect 3438 2850 3444 2851
rect 3564 2848 3566 2853
rect 2314 2847 2320 2848
rect 2314 2846 2315 2847
rect 2300 2844 2315 2846
rect 2194 2842 2200 2843
rect 2314 2843 2315 2844
rect 2319 2843 2320 2847
rect 2314 2842 2320 2843
rect 3562 2847 3568 2848
rect 3562 2843 3563 2847
rect 3567 2843 3568 2847
rect 3562 2842 3568 2843
rect 3590 2844 3596 2845
rect 183 2839 189 2840
rect 183 2835 184 2839
rect 188 2838 189 2839
rect 218 2839 224 2840
rect 218 2838 219 2839
rect 188 2836 219 2838
rect 188 2835 189 2836
rect 183 2834 189 2835
rect 218 2835 219 2836
rect 223 2835 224 2839
rect 218 2834 224 2835
rect 342 2839 349 2840
rect 342 2835 343 2839
rect 348 2835 349 2839
rect 342 2834 349 2835
rect 503 2839 509 2840
rect 503 2835 504 2839
rect 508 2838 509 2839
rect 538 2839 544 2840
rect 538 2838 539 2839
rect 508 2836 539 2838
rect 508 2835 509 2836
rect 503 2834 509 2835
rect 538 2835 539 2836
rect 543 2835 544 2839
rect 538 2834 544 2835
rect 663 2839 669 2840
rect 663 2835 664 2839
rect 668 2838 669 2839
rect 698 2839 704 2840
rect 698 2838 699 2839
rect 668 2836 699 2838
rect 668 2835 669 2836
rect 663 2834 669 2835
rect 698 2835 699 2836
rect 703 2835 704 2839
rect 698 2834 704 2835
rect 815 2839 821 2840
rect 815 2835 816 2839
rect 820 2838 821 2839
rect 854 2839 860 2840
rect 854 2838 855 2839
rect 820 2836 855 2838
rect 820 2835 821 2836
rect 815 2834 821 2835
rect 854 2835 855 2836
rect 859 2835 860 2839
rect 854 2834 860 2835
rect 959 2839 965 2840
rect 959 2835 960 2839
rect 964 2838 965 2839
rect 1006 2839 1012 2840
rect 1006 2838 1007 2839
rect 964 2836 1007 2838
rect 964 2835 965 2836
rect 959 2834 965 2835
rect 1006 2835 1007 2836
rect 1011 2835 1012 2839
rect 1006 2834 1012 2835
rect 1014 2839 1020 2840
rect 1014 2835 1015 2839
rect 1019 2838 1020 2839
rect 1087 2839 1093 2840
rect 1087 2838 1088 2839
rect 1019 2836 1088 2838
rect 1019 2835 1020 2836
rect 1014 2834 1020 2835
rect 1087 2835 1088 2836
rect 1092 2835 1093 2839
rect 1087 2834 1093 2835
rect 1122 2839 1128 2840
rect 1122 2835 1123 2839
rect 1127 2838 1128 2839
rect 1207 2839 1213 2840
rect 1207 2838 1208 2839
rect 1127 2836 1208 2838
rect 1127 2835 1128 2836
rect 1122 2834 1128 2835
rect 1207 2835 1208 2836
rect 1212 2835 1213 2839
rect 1207 2834 1213 2835
rect 1254 2839 1260 2840
rect 1254 2835 1255 2839
rect 1259 2838 1260 2839
rect 1319 2839 1325 2840
rect 1319 2838 1320 2839
rect 1259 2836 1320 2838
rect 1259 2835 1260 2836
rect 1254 2834 1260 2835
rect 1319 2835 1320 2836
rect 1324 2835 1325 2839
rect 1319 2834 1325 2835
rect 1423 2839 1432 2840
rect 1423 2835 1424 2839
rect 1431 2835 1432 2839
rect 1423 2834 1432 2835
rect 1462 2839 1468 2840
rect 1462 2835 1463 2839
rect 1467 2838 1468 2839
rect 1519 2839 1525 2840
rect 1519 2838 1520 2839
rect 1467 2836 1520 2838
rect 1467 2835 1468 2836
rect 1462 2834 1468 2835
rect 1519 2835 1520 2836
rect 1524 2835 1525 2839
rect 1519 2834 1525 2835
rect 1562 2839 1568 2840
rect 1562 2835 1563 2839
rect 1567 2838 1568 2839
rect 1623 2839 1629 2840
rect 1623 2838 1624 2839
rect 1567 2836 1624 2838
rect 1567 2835 1568 2836
rect 1562 2834 1568 2835
rect 1623 2835 1624 2836
rect 1628 2835 1629 2839
rect 1623 2834 1629 2835
rect 1666 2839 1672 2840
rect 1666 2835 1667 2839
rect 1671 2838 1672 2839
rect 1727 2839 1733 2840
rect 1870 2839 1876 2840
rect 3590 2840 3591 2844
rect 3595 2840 3596 2844
rect 3590 2839 3596 2840
rect 1727 2838 1728 2839
rect 1671 2836 1728 2838
rect 1671 2835 1672 2836
rect 1666 2834 1672 2835
rect 1727 2835 1728 2836
rect 1732 2835 1733 2839
rect 1727 2834 1733 2835
rect 1286 2831 1292 2832
rect 1286 2830 1287 2831
rect 1159 2828 1287 2830
rect 150 2823 156 2824
rect 150 2819 151 2823
rect 155 2822 156 2823
rect 167 2823 173 2824
rect 167 2822 168 2823
rect 155 2820 168 2822
rect 155 2819 156 2820
rect 150 2818 156 2819
rect 167 2819 168 2820
rect 172 2819 173 2823
rect 167 2818 173 2819
rect 194 2823 200 2824
rect 194 2819 195 2823
rect 199 2822 200 2823
rect 271 2823 277 2824
rect 271 2822 272 2823
rect 199 2820 272 2822
rect 199 2819 200 2820
rect 194 2818 200 2819
rect 271 2819 272 2820
rect 276 2819 277 2823
rect 271 2818 277 2819
rect 298 2823 304 2824
rect 298 2819 299 2823
rect 303 2822 304 2823
rect 407 2823 413 2824
rect 407 2822 408 2823
rect 303 2820 408 2822
rect 303 2819 304 2820
rect 298 2818 304 2819
rect 407 2819 408 2820
rect 412 2819 413 2823
rect 407 2818 413 2819
rect 559 2823 565 2824
rect 559 2819 560 2823
rect 564 2822 565 2823
rect 570 2823 576 2824
rect 570 2822 571 2823
rect 564 2820 571 2822
rect 564 2819 565 2820
rect 559 2818 565 2819
rect 570 2819 571 2820
rect 575 2819 576 2823
rect 570 2818 576 2819
rect 586 2823 592 2824
rect 586 2819 587 2823
rect 591 2822 592 2823
rect 711 2823 717 2824
rect 711 2822 712 2823
rect 591 2820 712 2822
rect 591 2819 592 2820
rect 586 2818 592 2819
rect 711 2819 712 2820
rect 716 2819 717 2823
rect 711 2818 717 2819
rect 738 2823 744 2824
rect 738 2819 739 2823
rect 743 2822 744 2823
rect 871 2823 877 2824
rect 871 2822 872 2823
rect 743 2820 872 2822
rect 743 2819 744 2820
rect 738 2818 744 2819
rect 871 2819 872 2820
rect 876 2819 877 2823
rect 871 2818 877 2819
rect 1023 2823 1029 2824
rect 1023 2819 1024 2823
rect 1028 2822 1029 2823
rect 1159 2822 1161 2828
rect 1286 2827 1287 2828
rect 1291 2827 1292 2831
rect 1286 2826 1292 2827
rect 2054 2826 2060 2827
rect 1028 2820 1161 2822
rect 1167 2823 1173 2824
rect 1028 2819 1029 2820
rect 1023 2818 1029 2819
rect 1167 2819 1168 2823
rect 1172 2822 1173 2823
rect 1202 2823 1208 2824
rect 1202 2822 1203 2823
rect 1172 2820 1203 2822
rect 1172 2819 1173 2820
rect 1167 2818 1173 2819
rect 1202 2819 1203 2820
rect 1207 2819 1208 2823
rect 1202 2818 1208 2819
rect 1230 2823 1236 2824
rect 1230 2819 1231 2823
rect 1235 2822 1236 2823
rect 1303 2823 1309 2824
rect 1303 2822 1304 2823
rect 1235 2820 1304 2822
rect 1235 2819 1236 2820
rect 1230 2818 1236 2819
rect 1303 2819 1304 2820
rect 1308 2819 1309 2823
rect 1303 2818 1309 2819
rect 1431 2823 1440 2824
rect 1431 2819 1432 2823
rect 1439 2819 1440 2823
rect 1431 2818 1440 2819
rect 1458 2823 1464 2824
rect 1458 2819 1459 2823
rect 1463 2822 1464 2823
rect 1551 2823 1557 2824
rect 1551 2822 1552 2823
rect 1463 2820 1552 2822
rect 1463 2819 1464 2820
rect 1458 2818 1464 2819
rect 1551 2819 1552 2820
rect 1556 2819 1557 2823
rect 1551 2818 1557 2819
rect 1578 2823 1584 2824
rect 1578 2819 1579 2823
rect 1583 2822 1584 2823
rect 1671 2823 1677 2824
rect 1671 2822 1672 2823
rect 1583 2820 1672 2822
rect 1583 2819 1584 2820
rect 1578 2818 1584 2819
rect 1671 2819 1672 2820
rect 1676 2819 1677 2823
rect 1671 2818 1677 2819
rect 1714 2823 1720 2824
rect 1714 2819 1715 2823
rect 1719 2822 1720 2823
rect 1775 2823 1781 2824
rect 1775 2822 1776 2823
rect 1719 2820 1776 2822
rect 1719 2819 1720 2820
rect 1714 2818 1720 2819
rect 1775 2819 1776 2820
rect 1780 2819 1781 2823
rect 2054 2822 2055 2826
rect 2059 2822 2060 2826
rect 2054 2821 2060 2822
rect 2142 2826 2148 2827
rect 2142 2822 2143 2826
rect 2147 2822 2148 2826
rect 2142 2821 2148 2822
rect 2246 2826 2252 2827
rect 2246 2822 2247 2826
rect 2251 2822 2252 2826
rect 2246 2821 2252 2822
rect 2350 2826 2356 2827
rect 2350 2822 2351 2826
rect 2355 2822 2356 2826
rect 2350 2821 2356 2822
rect 2470 2826 2476 2827
rect 2470 2822 2471 2826
rect 2475 2822 2476 2826
rect 2470 2821 2476 2822
rect 2598 2826 2604 2827
rect 2598 2822 2599 2826
rect 2603 2822 2604 2826
rect 2598 2821 2604 2822
rect 2734 2826 2740 2827
rect 2734 2822 2735 2826
rect 2739 2822 2740 2826
rect 2734 2821 2740 2822
rect 2886 2826 2892 2827
rect 2886 2822 2887 2826
rect 2891 2822 2892 2826
rect 2886 2821 2892 2822
rect 3038 2826 3044 2827
rect 3038 2822 3039 2826
rect 3043 2822 3044 2826
rect 3038 2821 3044 2822
rect 3198 2826 3204 2827
rect 3198 2822 3199 2826
rect 3203 2822 3204 2826
rect 3198 2821 3204 2822
rect 3366 2826 3372 2827
rect 3366 2822 3367 2826
rect 3371 2822 3372 2826
rect 3366 2821 3372 2822
rect 3510 2826 3516 2827
rect 3510 2822 3511 2826
rect 3515 2822 3516 2826
rect 3510 2821 3516 2822
rect 1775 2818 1781 2819
rect 2079 2815 2088 2816
rect 142 2814 148 2815
rect 142 2810 143 2814
rect 147 2810 148 2814
rect 142 2809 148 2810
rect 246 2814 252 2815
rect 246 2810 247 2814
rect 251 2810 252 2814
rect 246 2809 252 2810
rect 382 2814 388 2815
rect 382 2810 383 2814
rect 387 2810 388 2814
rect 382 2809 388 2810
rect 534 2814 540 2815
rect 534 2810 535 2814
rect 539 2810 540 2814
rect 534 2809 540 2810
rect 686 2814 692 2815
rect 686 2810 687 2814
rect 691 2810 692 2814
rect 686 2809 692 2810
rect 846 2814 852 2815
rect 846 2810 847 2814
rect 851 2810 852 2814
rect 846 2809 852 2810
rect 998 2814 1004 2815
rect 998 2810 999 2814
rect 1003 2810 1004 2814
rect 998 2809 1004 2810
rect 1142 2814 1148 2815
rect 1142 2810 1143 2814
rect 1147 2810 1148 2814
rect 1142 2809 1148 2810
rect 1278 2814 1284 2815
rect 1278 2810 1279 2814
rect 1283 2810 1284 2814
rect 1278 2809 1284 2810
rect 1406 2814 1412 2815
rect 1406 2810 1407 2814
rect 1411 2810 1412 2814
rect 1406 2809 1412 2810
rect 1526 2814 1532 2815
rect 1526 2810 1527 2814
rect 1531 2810 1532 2814
rect 1526 2809 1532 2810
rect 1646 2814 1652 2815
rect 1646 2810 1647 2814
rect 1651 2810 1652 2814
rect 1646 2809 1652 2810
rect 1750 2814 1756 2815
rect 1750 2810 1751 2814
rect 1755 2810 1756 2814
rect 2079 2811 2080 2815
rect 2087 2811 2088 2815
rect 2079 2810 2088 2811
rect 2114 2815 2120 2816
rect 2114 2811 2115 2815
rect 2119 2814 2120 2815
rect 2167 2815 2173 2816
rect 2167 2814 2168 2815
rect 2119 2812 2168 2814
rect 2119 2811 2120 2812
rect 2114 2810 2120 2811
rect 2167 2811 2168 2812
rect 2172 2811 2173 2815
rect 2167 2810 2173 2811
rect 2271 2815 2277 2816
rect 2271 2811 2272 2815
rect 2276 2814 2277 2815
rect 2306 2815 2312 2816
rect 2306 2814 2307 2815
rect 2276 2812 2307 2814
rect 2276 2811 2277 2812
rect 2271 2810 2277 2811
rect 2306 2811 2307 2812
rect 2311 2811 2312 2815
rect 2306 2810 2312 2811
rect 2375 2815 2381 2816
rect 2375 2811 2376 2815
rect 2380 2814 2381 2815
rect 2410 2815 2416 2816
rect 2410 2814 2411 2815
rect 2380 2812 2411 2814
rect 2380 2811 2381 2812
rect 2375 2810 2381 2811
rect 2410 2811 2411 2812
rect 2415 2811 2416 2815
rect 2410 2810 2416 2811
rect 2494 2815 2501 2816
rect 2494 2811 2495 2815
rect 2500 2811 2501 2815
rect 2494 2810 2501 2811
rect 2623 2815 2632 2816
rect 2623 2811 2624 2815
rect 2631 2811 2632 2815
rect 2623 2810 2632 2811
rect 2682 2815 2688 2816
rect 2682 2811 2683 2815
rect 2687 2814 2688 2815
rect 2759 2815 2765 2816
rect 2759 2814 2760 2815
rect 2687 2812 2760 2814
rect 2687 2811 2688 2812
rect 2682 2810 2688 2811
rect 2759 2811 2760 2812
rect 2764 2811 2765 2815
rect 2759 2810 2765 2811
rect 2794 2815 2800 2816
rect 2794 2811 2795 2815
rect 2799 2814 2800 2815
rect 2911 2815 2917 2816
rect 2911 2814 2912 2815
rect 2799 2812 2912 2814
rect 2799 2811 2800 2812
rect 2794 2810 2800 2811
rect 2911 2811 2912 2812
rect 2916 2811 2917 2815
rect 2911 2810 2917 2811
rect 3063 2815 3069 2816
rect 3063 2811 3064 2815
rect 3068 2814 3069 2815
rect 3098 2815 3104 2816
rect 3098 2814 3099 2815
rect 3068 2812 3099 2814
rect 3068 2811 3069 2812
rect 3063 2810 3069 2811
rect 3098 2811 3099 2812
rect 3103 2811 3104 2815
rect 3098 2810 3104 2811
rect 3223 2815 3232 2816
rect 3223 2811 3224 2815
rect 3231 2811 3232 2815
rect 3223 2810 3232 2811
rect 3390 2815 3397 2816
rect 3390 2811 3391 2815
rect 3396 2811 3397 2815
rect 3390 2810 3397 2811
rect 3534 2815 3541 2816
rect 3534 2811 3535 2815
rect 3540 2811 3541 2815
rect 3534 2810 3541 2811
rect 1750 2809 1756 2810
rect 2022 2799 2028 2800
rect 2022 2798 2023 2799
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 1830 2796 1836 2797
rect 1830 2792 1831 2796
rect 1835 2792 1836 2796
rect 1948 2796 2023 2798
rect 1830 2791 1836 2792
rect 1927 2791 1933 2792
rect 194 2787 200 2788
rect 194 2783 195 2787
rect 199 2783 200 2787
rect 194 2782 200 2783
rect 298 2787 304 2788
rect 298 2783 299 2787
rect 303 2783 304 2787
rect 298 2782 304 2783
rect 586 2787 592 2788
rect 586 2783 587 2787
rect 591 2783 592 2787
rect 586 2782 592 2783
rect 738 2787 744 2788
rect 738 2783 739 2787
rect 743 2783 744 2787
rect 738 2782 744 2783
rect 854 2787 860 2788
rect 854 2783 855 2787
rect 859 2783 860 2787
rect 854 2782 860 2783
rect 1006 2787 1012 2788
rect 1006 2783 1007 2787
rect 1011 2783 1012 2787
rect 1230 2787 1236 2788
rect 1230 2786 1231 2787
rect 1197 2784 1231 2786
rect 1006 2782 1012 2783
rect 1230 2783 1231 2784
rect 1235 2783 1236 2787
rect 1230 2782 1236 2783
rect 1286 2787 1292 2788
rect 1286 2783 1287 2787
rect 1291 2783 1292 2787
rect 1286 2782 1292 2783
rect 1458 2787 1464 2788
rect 1458 2783 1459 2787
rect 1463 2783 1464 2787
rect 1458 2782 1464 2783
rect 1578 2787 1584 2788
rect 1578 2783 1579 2787
rect 1583 2783 1584 2787
rect 1714 2787 1720 2788
rect 1714 2786 1715 2787
rect 1701 2784 1715 2786
rect 1578 2782 1584 2783
rect 1714 2783 1715 2784
rect 1719 2783 1720 2787
rect 1927 2787 1928 2791
rect 1932 2790 1933 2791
rect 1948 2790 1950 2796
rect 2022 2795 2023 2796
rect 2027 2795 2028 2799
rect 2022 2794 2028 2795
rect 1932 2788 1950 2790
rect 1954 2791 1960 2792
rect 1932 2787 1933 2788
rect 1927 2786 1933 2787
rect 1954 2787 1955 2791
rect 1959 2790 1960 2791
rect 2039 2791 2045 2792
rect 2039 2790 2040 2791
rect 1959 2788 2040 2790
rect 1959 2787 1960 2788
rect 1954 2786 1960 2787
rect 2039 2787 2040 2788
rect 2044 2787 2045 2791
rect 2039 2786 2045 2787
rect 2191 2791 2200 2792
rect 2191 2787 2192 2791
rect 2199 2787 2200 2791
rect 2191 2786 2200 2787
rect 2218 2791 2224 2792
rect 2218 2787 2219 2791
rect 2223 2790 2224 2791
rect 2351 2791 2357 2792
rect 2351 2790 2352 2791
rect 2223 2788 2352 2790
rect 2223 2787 2224 2788
rect 2218 2786 2224 2787
rect 2351 2787 2352 2788
rect 2356 2787 2357 2791
rect 2351 2786 2357 2787
rect 2418 2791 2424 2792
rect 2418 2787 2419 2791
rect 2423 2790 2424 2791
rect 2511 2791 2517 2792
rect 2511 2790 2512 2791
rect 2423 2788 2512 2790
rect 2423 2787 2424 2788
rect 2418 2786 2424 2787
rect 2511 2787 2512 2788
rect 2516 2787 2517 2791
rect 2511 2786 2517 2787
rect 2663 2791 2672 2792
rect 2663 2787 2664 2791
rect 2671 2787 2672 2791
rect 2663 2786 2672 2787
rect 2690 2791 2696 2792
rect 2690 2787 2691 2791
rect 2695 2790 2696 2791
rect 2815 2791 2821 2792
rect 2815 2790 2816 2791
rect 2695 2788 2816 2790
rect 2695 2787 2696 2788
rect 2690 2786 2696 2787
rect 2815 2787 2816 2788
rect 2820 2787 2821 2791
rect 2815 2786 2821 2787
rect 2842 2791 2848 2792
rect 2842 2787 2843 2791
rect 2847 2790 2848 2791
rect 2967 2791 2973 2792
rect 2967 2790 2968 2791
rect 2847 2788 2968 2790
rect 2847 2787 2848 2788
rect 2842 2786 2848 2787
rect 2967 2787 2968 2788
rect 2972 2787 2973 2791
rect 2967 2786 2973 2787
rect 2994 2791 3000 2792
rect 2994 2787 2995 2791
rect 2999 2790 3000 2791
rect 3111 2791 3117 2792
rect 3111 2790 3112 2791
rect 2999 2788 3112 2790
rect 2999 2787 3000 2788
rect 2994 2786 3000 2787
rect 3111 2787 3112 2788
rect 3116 2787 3117 2791
rect 3111 2786 3117 2787
rect 3138 2791 3144 2792
rect 3138 2787 3139 2791
rect 3143 2790 3144 2791
rect 3255 2791 3261 2792
rect 3255 2790 3256 2791
rect 3143 2788 3256 2790
rect 3143 2787 3144 2788
rect 3138 2786 3144 2787
rect 3255 2787 3256 2788
rect 3260 2787 3261 2791
rect 3255 2786 3261 2787
rect 3407 2791 3413 2792
rect 3407 2787 3408 2791
rect 3412 2790 3413 2791
rect 3442 2791 3448 2792
rect 3442 2790 3443 2791
rect 3412 2788 3443 2790
rect 3412 2787 3413 2788
rect 3407 2786 3413 2787
rect 3442 2787 3443 2788
rect 3447 2787 3448 2791
rect 3442 2786 3448 2787
rect 3535 2791 3541 2792
rect 3535 2787 3536 2791
rect 3540 2790 3541 2791
rect 3562 2791 3568 2792
rect 3562 2790 3563 2791
rect 3540 2788 3563 2790
rect 3540 2787 3541 2788
rect 3535 2786 3541 2787
rect 3562 2787 3563 2788
rect 3567 2787 3568 2791
rect 3562 2786 3568 2787
rect 1714 2782 1720 2783
rect 1902 2782 1908 2783
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 1830 2779 1836 2780
rect 110 2774 116 2775
rect 134 2776 140 2777
rect 134 2772 135 2776
rect 139 2772 140 2776
rect 134 2771 140 2772
rect 238 2776 244 2777
rect 238 2772 239 2776
rect 243 2772 244 2776
rect 238 2771 244 2772
rect 374 2776 380 2777
rect 374 2772 375 2776
rect 379 2772 380 2776
rect 374 2771 380 2772
rect 526 2776 532 2777
rect 526 2772 527 2776
rect 531 2772 532 2776
rect 526 2771 532 2772
rect 678 2776 684 2777
rect 678 2772 679 2776
rect 683 2772 684 2776
rect 678 2771 684 2772
rect 838 2776 844 2777
rect 838 2772 839 2776
rect 843 2772 844 2776
rect 838 2771 844 2772
rect 990 2776 996 2777
rect 990 2772 991 2776
rect 995 2772 996 2776
rect 990 2771 996 2772
rect 1134 2776 1140 2777
rect 1134 2772 1135 2776
rect 1139 2772 1140 2776
rect 1134 2771 1140 2772
rect 1270 2776 1276 2777
rect 1270 2772 1271 2776
rect 1275 2772 1276 2776
rect 1270 2771 1276 2772
rect 1398 2776 1404 2777
rect 1398 2772 1399 2776
rect 1403 2772 1404 2776
rect 1398 2771 1404 2772
rect 1518 2776 1524 2777
rect 1518 2772 1519 2776
rect 1523 2772 1524 2776
rect 1518 2771 1524 2772
rect 1638 2776 1644 2777
rect 1638 2772 1639 2776
rect 1643 2772 1644 2776
rect 1638 2771 1644 2772
rect 1742 2776 1748 2777
rect 1742 2772 1743 2776
rect 1747 2772 1748 2776
rect 1830 2775 1831 2779
rect 1835 2775 1836 2779
rect 1902 2778 1903 2782
rect 1907 2778 1908 2782
rect 1902 2777 1908 2778
rect 2014 2782 2020 2783
rect 2014 2778 2015 2782
rect 2019 2778 2020 2782
rect 2014 2777 2020 2778
rect 2166 2782 2172 2783
rect 2166 2778 2167 2782
rect 2171 2778 2172 2782
rect 2166 2777 2172 2778
rect 2326 2782 2332 2783
rect 2326 2778 2327 2782
rect 2331 2778 2332 2782
rect 2326 2777 2332 2778
rect 2486 2782 2492 2783
rect 2486 2778 2487 2782
rect 2491 2778 2492 2782
rect 2486 2777 2492 2778
rect 2638 2782 2644 2783
rect 2638 2778 2639 2782
rect 2643 2778 2644 2782
rect 2638 2777 2644 2778
rect 2790 2782 2796 2783
rect 2790 2778 2791 2782
rect 2795 2778 2796 2782
rect 2790 2777 2796 2778
rect 2942 2782 2948 2783
rect 2942 2778 2943 2782
rect 2947 2778 2948 2782
rect 2942 2777 2948 2778
rect 3086 2782 3092 2783
rect 3086 2778 3087 2782
rect 3091 2778 3092 2782
rect 3086 2777 3092 2778
rect 3230 2782 3236 2783
rect 3230 2778 3231 2782
rect 3235 2778 3236 2782
rect 3230 2777 3236 2778
rect 3382 2782 3388 2783
rect 3382 2778 3383 2782
rect 3387 2778 3388 2782
rect 3382 2777 3388 2778
rect 3510 2782 3516 2783
rect 3510 2778 3511 2782
rect 3515 2778 3516 2782
rect 3510 2777 3516 2778
rect 1830 2774 1836 2775
rect 1742 2771 1748 2772
rect 1870 2764 1876 2765
rect 1870 2760 1871 2764
rect 1875 2760 1876 2764
rect 391 2759 400 2760
rect 391 2755 392 2759
rect 399 2755 400 2759
rect 391 2754 400 2755
rect 1730 2759 1736 2760
rect 1730 2755 1731 2759
rect 1735 2758 1736 2759
rect 1759 2759 1765 2760
rect 1870 2759 1876 2760
rect 3590 2764 3596 2765
rect 3590 2760 3591 2764
rect 3595 2760 3596 2764
rect 3590 2759 3596 2760
rect 1759 2758 1760 2759
rect 1735 2756 1760 2758
rect 1735 2755 1736 2756
rect 1730 2754 1736 2755
rect 1759 2755 1760 2756
rect 1764 2755 1765 2759
rect 1759 2754 1765 2755
rect 1954 2755 1960 2756
rect 1954 2751 1955 2755
rect 1959 2751 1960 2755
rect 1954 2750 1960 2751
rect 2066 2755 2072 2756
rect 2066 2751 2067 2755
rect 2071 2751 2072 2755
rect 2066 2750 2072 2751
rect 2218 2755 2224 2756
rect 2218 2751 2219 2755
rect 2223 2751 2224 2755
rect 2218 2750 2224 2751
rect 2358 2755 2364 2756
rect 2358 2751 2359 2755
rect 2363 2751 2364 2755
rect 2358 2750 2364 2751
rect 2494 2755 2500 2756
rect 2494 2751 2495 2755
rect 2499 2751 2500 2755
rect 2494 2750 2500 2751
rect 2690 2755 2696 2756
rect 2690 2751 2691 2755
rect 2695 2751 2696 2755
rect 2690 2750 2696 2751
rect 2842 2755 2848 2756
rect 2842 2751 2843 2755
rect 2847 2751 2848 2755
rect 2842 2750 2848 2751
rect 2994 2755 3000 2756
rect 2994 2751 2995 2755
rect 2999 2751 3000 2755
rect 2994 2750 3000 2751
rect 3138 2755 3144 2756
rect 3138 2751 3139 2755
rect 3143 2751 3144 2755
rect 3138 2750 3144 2751
rect 3390 2755 3396 2756
rect 3390 2751 3391 2755
rect 3395 2751 3396 2755
rect 3390 2750 3396 2751
rect 3534 2755 3540 2756
rect 3534 2751 3535 2755
rect 3539 2751 3540 2755
rect 3534 2750 3540 2751
rect 1870 2747 1876 2748
rect 1870 2743 1871 2747
rect 1875 2743 1876 2747
rect 3590 2747 3596 2748
rect 1870 2742 1876 2743
rect 1894 2744 1900 2745
rect 1894 2740 1895 2744
rect 1899 2740 1900 2744
rect 1894 2739 1900 2740
rect 2006 2744 2012 2745
rect 2006 2740 2007 2744
rect 2011 2740 2012 2744
rect 2006 2739 2012 2740
rect 2158 2744 2164 2745
rect 2158 2740 2159 2744
rect 2163 2740 2164 2744
rect 2158 2739 2164 2740
rect 2318 2744 2324 2745
rect 2318 2740 2319 2744
rect 2323 2740 2324 2744
rect 2318 2739 2324 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2630 2744 2636 2745
rect 2630 2740 2631 2744
rect 2635 2740 2636 2744
rect 2630 2739 2636 2740
rect 2782 2744 2788 2745
rect 2782 2740 2783 2744
rect 2787 2740 2788 2744
rect 2782 2739 2788 2740
rect 2934 2744 2940 2745
rect 2934 2740 2935 2744
rect 2939 2740 2940 2744
rect 2934 2739 2940 2740
rect 3078 2744 3084 2745
rect 3078 2740 3079 2744
rect 3083 2740 3084 2744
rect 3078 2739 3084 2740
rect 3222 2744 3228 2745
rect 3222 2740 3223 2744
rect 3227 2740 3228 2744
rect 3222 2739 3228 2740
rect 3374 2744 3380 2745
rect 3374 2740 3375 2744
rect 3379 2740 3380 2744
rect 3374 2739 3380 2740
rect 3502 2744 3508 2745
rect 3502 2740 3503 2744
rect 3507 2740 3508 2744
rect 3590 2743 3591 2747
rect 3595 2743 3596 2747
rect 3590 2742 3596 2743
rect 3502 2739 3508 2740
rect 134 2728 140 2729
rect 110 2725 116 2726
rect 110 2721 111 2725
rect 115 2721 116 2725
rect 134 2724 135 2728
rect 139 2724 140 2728
rect 134 2723 140 2724
rect 230 2728 236 2729
rect 230 2724 231 2728
rect 235 2724 236 2728
rect 230 2723 236 2724
rect 366 2728 372 2729
rect 366 2724 367 2728
rect 371 2724 372 2728
rect 366 2723 372 2724
rect 510 2728 516 2729
rect 510 2724 511 2728
rect 515 2724 516 2728
rect 510 2723 516 2724
rect 662 2728 668 2729
rect 662 2724 663 2728
rect 667 2724 668 2728
rect 662 2723 668 2724
rect 814 2728 820 2729
rect 814 2724 815 2728
rect 819 2724 820 2728
rect 814 2723 820 2724
rect 974 2728 980 2729
rect 974 2724 975 2728
rect 979 2724 980 2728
rect 974 2723 980 2724
rect 1134 2728 1140 2729
rect 1134 2724 1135 2728
rect 1139 2724 1140 2728
rect 1134 2723 1140 2724
rect 1286 2728 1292 2729
rect 1286 2724 1287 2728
rect 1291 2724 1292 2728
rect 1286 2723 1292 2724
rect 1446 2728 1452 2729
rect 1446 2724 1447 2728
rect 1451 2724 1452 2728
rect 1446 2723 1452 2724
rect 1606 2728 1612 2729
rect 1606 2724 1607 2728
rect 1611 2724 1612 2728
rect 1606 2723 1612 2724
rect 1742 2728 1748 2729
rect 1742 2724 1743 2728
rect 1747 2724 1748 2728
rect 3138 2727 3144 2728
rect 1742 2723 1748 2724
rect 1830 2725 1836 2726
rect 110 2720 116 2721
rect 1830 2721 1831 2725
rect 1835 2721 1836 2725
rect 3138 2723 3139 2727
rect 3143 2726 3144 2727
rect 3239 2727 3245 2728
rect 3239 2726 3240 2727
rect 3143 2724 3240 2726
rect 3143 2723 3144 2724
rect 3138 2722 3144 2723
rect 3239 2723 3240 2724
rect 3244 2723 3245 2727
rect 3239 2722 3245 2723
rect 1830 2720 1836 2721
rect 202 2719 208 2720
rect 196 2712 198 2717
rect 202 2715 203 2719
rect 207 2718 208 2719
rect 298 2719 304 2720
rect 207 2716 249 2718
rect 207 2715 208 2716
rect 202 2714 208 2715
rect 298 2715 299 2719
rect 303 2718 304 2719
rect 578 2719 584 2720
rect 303 2716 385 2718
rect 303 2715 304 2716
rect 298 2714 304 2715
rect 572 2712 574 2717
rect 578 2715 579 2719
rect 583 2718 584 2719
rect 730 2719 736 2720
rect 583 2716 681 2718
rect 583 2715 584 2716
rect 578 2714 584 2715
rect 730 2715 731 2719
rect 735 2718 736 2719
rect 1070 2719 1076 2720
rect 1070 2718 1071 2719
rect 735 2716 833 2718
rect 1037 2716 1071 2718
rect 735 2715 736 2716
rect 730 2714 736 2715
rect 1070 2715 1071 2716
rect 1075 2715 1076 2719
rect 1202 2719 1208 2720
rect 1202 2718 1203 2719
rect 1197 2716 1203 2718
rect 1070 2714 1076 2715
rect 1202 2715 1203 2716
rect 1207 2715 1208 2719
rect 1202 2714 1208 2715
rect 1222 2719 1228 2720
rect 1222 2715 1223 2719
rect 1227 2718 1228 2719
rect 1354 2719 1360 2720
rect 1227 2716 1305 2718
rect 1227 2715 1228 2716
rect 1222 2714 1228 2715
rect 1354 2715 1355 2719
rect 1359 2718 1360 2719
rect 1842 2719 1848 2720
rect 1842 2718 1843 2719
rect 1359 2716 1465 2718
rect 1359 2715 1360 2716
rect 1354 2714 1360 2715
rect 1668 2714 1670 2717
rect 1805 2716 1843 2718
rect 1738 2715 1744 2716
rect 1738 2714 1739 2715
rect 1668 2712 1739 2714
rect 194 2711 200 2712
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 194 2707 195 2711
rect 199 2707 200 2711
rect 194 2706 200 2707
rect 570 2711 576 2712
rect 570 2707 571 2711
rect 575 2707 576 2711
rect 1738 2711 1739 2712
rect 1743 2711 1744 2715
rect 1842 2715 1843 2716
rect 1847 2715 1848 2719
rect 1842 2714 1848 2715
rect 1738 2710 1744 2711
rect 570 2706 576 2707
rect 1830 2708 1836 2709
rect 110 2703 116 2704
rect 1830 2704 1831 2708
rect 1835 2704 1836 2708
rect 1830 2703 1836 2704
rect 1894 2700 1900 2701
rect 1870 2697 1876 2698
rect 1870 2693 1871 2697
rect 1875 2693 1876 2697
rect 1894 2696 1895 2700
rect 1899 2696 1900 2700
rect 1894 2695 1900 2696
rect 2102 2700 2108 2701
rect 2102 2696 2103 2700
rect 2107 2696 2108 2700
rect 2102 2695 2108 2696
rect 2326 2700 2332 2701
rect 2326 2696 2327 2700
rect 2331 2696 2332 2700
rect 2326 2695 2332 2696
rect 2534 2700 2540 2701
rect 2534 2696 2535 2700
rect 2539 2696 2540 2700
rect 2534 2695 2540 2696
rect 2734 2700 2740 2701
rect 2734 2696 2735 2700
rect 2739 2696 2740 2700
rect 2734 2695 2740 2696
rect 2910 2700 2916 2701
rect 2910 2696 2911 2700
rect 2915 2696 2916 2700
rect 2910 2695 2916 2696
rect 3070 2700 3076 2701
rect 3070 2696 3071 2700
rect 3075 2696 3076 2700
rect 3070 2695 3076 2696
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3374 2700 3380 2701
rect 3374 2696 3375 2700
rect 3379 2696 3380 2700
rect 3374 2695 3380 2696
rect 3502 2700 3508 2701
rect 3502 2696 3503 2700
rect 3507 2696 3508 2700
rect 3502 2695 3508 2696
rect 3590 2697 3596 2698
rect 1870 2692 1876 2693
rect 3590 2693 3591 2697
rect 3595 2693 3596 2697
rect 3590 2692 3596 2693
rect 2095 2691 2101 2692
rect 142 2690 148 2691
rect 142 2686 143 2690
rect 147 2686 148 2690
rect 142 2685 148 2686
rect 238 2690 244 2691
rect 238 2686 239 2690
rect 243 2686 244 2690
rect 238 2685 244 2686
rect 374 2690 380 2691
rect 374 2686 375 2690
rect 379 2686 380 2690
rect 374 2685 380 2686
rect 518 2690 524 2691
rect 518 2686 519 2690
rect 523 2686 524 2690
rect 518 2685 524 2686
rect 670 2690 676 2691
rect 670 2686 671 2690
rect 675 2686 676 2690
rect 670 2685 676 2686
rect 822 2690 828 2691
rect 822 2686 823 2690
rect 827 2686 828 2690
rect 822 2685 828 2686
rect 982 2690 988 2691
rect 982 2686 983 2690
rect 987 2686 988 2690
rect 982 2685 988 2686
rect 1142 2690 1148 2691
rect 1142 2686 1143 2690
rect 1147 2686 1148 2690
rect 1142 2685 1148 2686
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1454 2690 1460 2691
rect 1454 2686 1455 2690
rect 1459 2686 1460 2690
rect 1454 2685 1460 2686
rect 1614 2690 1620 2691
rect 1614 2686 1615 2690
rect 1619 2686 1620 2690
rect 1614 2685 1620 2686
rect 1750 2690 1756 2691
rect 2095 2690 2096 2691
rect 1750 2686 1751 2690
rect 1755 2686 1756 2690
rect 1957 2688 2096 2690
rect 2095 2687 2096 2688
rect 2100 2687 2101 2691
rect 2454 2691 2460 2692
rect 2454 2690 2455 2691
rect 2095 2686 2101 2687
rect 1750 2685 1756 2686
rect 2022 2683 2028 2684
rect 1870 2680 1876 2681
rect 167 2679 173 2680
rect 167 2675 168 2679
rect 172 2678 173 2679
rect 202 2679 208 2680
rect 202 2678 203 2679
rect 172 2676 203 2678
rect 172 2675 173 2676
rect 167 2674 173 2675
rect 202 2675 203 2676
rect 207 2675 208 2679
rect 202 2674 208 2675
rect 263 2679 269 2680
rect 263 2675 264 2679
rect 268 2678 269 2679
rect 298 2679 304 2680
rect 298 2678 299 2679
rect 268 2676 299 2678
rect 268 2675 269 2676
rect 263 2674 269 2675
rect 298 2675 299 2676
rect 303 2675 304 2679
rect 298 2674 304 2675
rect 394 2679 405 2680
rect 394 2675 395 2679
rect 399 2675 400 2679
rect 404 2675 405 2679
rect 394 2674 405 2675
rect 543 2679 549 2680
rect 543 2675 544 2679
rect 548 2678 549 2679
rect 578 2679 584 2680
rect 578 2678 579 2679
rect 548 2676 579 2678
rect 548 2675 549 2676
rect 543 2674 549 2675
rect 578 2675 579 2676
rect 583 2675 584 2679
rect 578 2674 584 2675
rect 695 2679 701 2680
rect 695 2675 696 2679
rect 700 2678 701 2679
rect 730 2679 736 2680
rect 730 2678 731 2679
rect 700 2676 731 2678
rect 700 2675 701 2676
rect 695 2674 701 2675
rect 730 2675 731 2676
rect 735 2675 736 2679
rect 730 2674 736 2675
rect 842 2679 853 2680
rect 842 2675 843 2679
rect 847 2675 848 2679
rect 852 2675 853 2679
rect 842 2674 853 2675
rect 1006 2679 1013 2680
rect 1006 2675 1007 2679
rect 1012 2675 1013 2679
rect 1006 2674 1013 2675
rect 1070 2679 1076 2680
rect 1070 2675 1071 2679
rect 1075 2678 1076 2679
rect 1167 2679 1173 2680
rect 1167 2678 1168 2679
rect 1075 2676 1168 2678
rect 1075 2675 1076 2676
rect 1070 2674 1076 2675
rect 1167 2675 1168 2676
rect 1172 2675 1173 2679
rect 1167 2674 1173 2675
rect 1319 2679 1325 2680
rect 1319 2675 1320 2679
rect 1324 2678 1325 2679
rect 1354 2679 1360 2680
rect 1354 2678 1355 2679
rect 1324 2676 1355 2678
rect 1324 2675 1325 2676
rect 1319 2674 1325 2675
rect 1354 2675 1355 2676
rect 1359 2675 1360 2679
rect 1354 2674 1360 2675
rect 1479 2679 1485 2680
rect 1479 2675 1480 2679
rect 1484 2678 1485 2679
rect 1558 2679 1564 2680
rect 1558 2678 1559 2679
rect 1484 2676 1559 2678
rect 1484 2675 1485 2676
rect 1479 2674 1485 2675
rect 1558 2675 1559 2676
rect 1563 2675 1564 2679
rect 1558 2674 1564 2675
rect 1639 2679 1645 2680
rect 1639 2675 1640 2679
rect 1644 2678 1645 2679
rect 1730 2679 1736 2680
rect 1730 2678 1731 2679
rect 1644 2676 1731 2678
rect 1644 2675 1645 2676
rect 1639 2674 1645 2675
rect 1730 2675 1731 2676
rect 1735 2675 1736 2679
rect 1730 2674 1736 2675
rect 1738 2679 1744 2680
rect 1738 2675 1739 2679
rect 1743 2678 1744 2679
rect 1775 2679 1781 2680
rect 1775 2678 1776 2679
rect 1743 2676 1776 2678
rect 1743 2675 1744 2676
rect 1738 2674 1744 2675
rect 1775 2675 1776 2676
rect 1780 2675 1781 2679
rect 1870 2676 1871 2680
rect 1875 2676 1876 2680
rect 2022 2679 2023 2683
rect 2027 2682 2028 2683
rect 2120 2682 2122 2689
rect 2389 2688 2455 2690
rect 2454 2687 2455 2688
rect 2459 2687 2460 2691
rect 2454 2686 2460 2687
rect 2478 2691 2484 2692
rect 2478 2687 2479 2691
rect 2483 2690 2484 2691
rect 2903 2691 2909 2692
rect 2903 2690 2904 2691
rect 2483 2688 2553 2690
rect 2797 2688 2904 2690
rect 2483 2687 2484 2688
rect 2478 2686 2484 2687
rect 2903 2687 2904 2688
rect 2908 2687 2909 2691
rect 3014 2691 3020 2692
rect 3014 2690 3015 2691
rect 2973 2688 3015 2690
rect 2903 2686 2909 2687
rect 3014 2687 3015 2688
rect 3019 2687 3020 2691
rect 3170 2691 3176 2692
rect 3170 2690 3171 2691
rect 3133 2688 3171 2690
rect 3014 2686 3020 2687
rect 3170 2687 3171 2688
rect 3175 2687 3176 2691
rect 3322 2691 3328 2692
rect 3322 2690 3323 2691
rect 3285 2688 3323 2690
rect 3170 2686 3176 2687
rect 3322 2687 3323 2688
rect 3327 2687 3328 2691
rect 3442 2691 3448 2692
rect 3442 2690 3443 2691
rect 3437 2688 3443 2690
rect 3322 2686 3328 2687
rect 3442 2687 3443 2688
rect 3447 2687 3448 2691
rect 3570 2691 3576 2692
rect 3570 2690 3571 2691
rect 3565 2688 3571 2690
rect 3442 2686 3448 2687
rect 3570 2687 3571 2688
rect 3575 2687 3576 2691
rect 3570 2686 3576 2687
rect 2027 2680 2122 2682
rect 3590 2680 3596 2681
rect 2027 2679 2028 2680
rect 2022 2678 2028 2679
rect 1870 2675 1876 2676
rect 3590 2676 3591 2680
rect 3595 2676 3596 2680
rect 3590 2675 3596 2676
rect 1775 2674 1781 2675
rect 1902 2662 1908 2663
rect 167 2659 173 2660
rect 167 2655 168 2659
rect 172 2658 173 2659
rect 194 2659 200 2660
rect 194 2658 195 2659
rect 172 2656 195 2658
rect 172 2655 173 2656
rect 167 2654 173 2655
rect 194 2655 195 2656
rect 199 2655 200 2659
rect 194 2654 200 2655
rect 239 2659 245 2660
rect 239 2655 240 2659
rect 244 2658 245 2659
rect 303 2659 309 2660
rect 303 2658 304 2659
rect 244 2656 304 2658
rect 244 2655 245 2656
rect 239 2654 245 2655
rect 303 2655 304 2656
rect 308 2655 309 2659
rect 303 2654 309 2655
rect 330 2659 336 2660
rect 330 2655 331 2659
rect 335 2658 336 2659
rect 471 2659 477 2660
rect 471 2658 472 2659
rect 335 2656 472 2658
rect 335 2655 336 2656
rect 330 2654 336 2655
rect 471 2655 472 2656
rect 476 2655 477 2659
rect 471 2654 477 2655
rect 586 2659 592 2660
rect 586 2655 587 2659
rect 591 2658 592 2659
rect 647 2659 653 2660
rect 647 2658 648 2659
rect 591 2656 648 2658
rect 591 2655 592 2656
rect 586 2654 592 2655
rect 647 2655 648 2656
rect 652 2655 653 2659
rect 647 2654 653 2655
rect 735 2659 741 2660
rect 735 2655 736 2659
rect 740 2658 741 2659
rect 815 2659 821 2660
rect 815 2658 816 2659
rect 740 2656 816 2658
rect 740 2655 741 2656
rect 735 2654 741 2655
rect 815 2655 816 2656
rect 820 2655 821 2659
rect 815 2654 821 2655
rect 975 2659 981 2660
rect 975 2655 976 2659
rect 980 2658 981 2659
rect 990 2659 996 2660
rect 990 2658 991 2659
rect 980 2656 991 2658
rect 980 2655 981 2656
rect 975 2654 981 2655
rect 990 2655 991 2656
rect 995 2655 996 2659
rect 990 2654 996 2655
rect 1002 2659 1008 2660
rect 1002 2655 1003 2659
rect 1007 2658 1008 2659
rect 1127 2659 1133 2660
rect 1127 2658 1128 2659
rect 1007 2656 1128 2658
rect 1007 2655 1008 2656
rect 1002 2654 1008 2655
rect 1127 2655 1128 2656
rect 1132 2655 1133 2659
rect 1127 2654 1133 2655
rect 1154 2659 1160 2660
rect 1154 2655 1155 2659
rect 1159 2658 1160 2659
rect 1271 2659 1277 2660
rect 1271 2658 1272 2659
rect 1159 2656 1272 2658
rect 1159 2655 1160 2656
rect 1154 2654 1160 2655
rect 1271 2655 1272 2656
rect 1276 2655 1277 2659
rect 1271 2654 1277 2655
rect 1390 2659 1396 2660
rect 1390 2655 1391 2659
rect 1395 2658 1396 2659
rect 1423 2659 1429 2660
rect 1423 2658 1424 2659
rect 1395 2656 1424 2658
rect 1395 2655 1396 2656
rect 1390 2654 1396 2655
rect 1423 2655 1424 2656
rect 1428 2655 1429 2659
rect 1423 2654 1429 2655
rect 1542 2659 1548 2660
rect 1542 2655 1543 2659
rect 1547 2658 1548 2659
rect 1575 2659 1581 2660
rect 1575 2658 1576 2659
rect 1547 2656 1576 2658
rect 1547 2655 1548 2656
rect 1542 2654 1548 2655
rect 1575 2655 1576 2656
rect 1580 2655 1581 2659
rect 1902 2658 1903 2662
rect 1907 2658 1908 2662
rect 1902 2657 1908 2658
rect 2110 2662 2116 2663
rect 2110 2658 2111 2662
rect 2115 2658 2116 2662
rect 2110 2657 2116 2658
rect 2334 2662 2340 2663
rect 2334 2658 2335 2662
rect 2339 2658 2340 2662
rect 2334 2657 2340 2658
rect 2542 2662 2548 2663
rect 2542 2658 2543 2662
rect 2547 2658 2548 2662
rect 2542 2657 2548 2658
rect 2742 2662 2748 2663
rect 2742 2658 2743 2662
rect 2747 2658 2748 2662
rect 2742 2657 2748 2658
rect 2918 2662 2924 2663
rect 2918 2658 2919 2662
rect 2923 2658 2924 2662
rect 2918 2657 2924 2658
rect 3078 2662 3084 2663
rect 3078 2658 3079 2662
rect 3083 2658 3084 2662
rect 3078 2657 3084 2658
rect 3230 2662 3236 2663
rect 3230 2658 3231 2662
rect 3235 2658 3236 2662
rect 3230 2657 3236 2658
rect 3382 2662 3388 2663
rect 3382 2658 3383 2662
rect 3387 2658 3388 2662
rect 3382 2657 3388 2658
rect 3510 2662 3516 2663
rect 3510 2658 3511 2662
rect 3515 2658 3516 2662
rect 3510 2657 3516 2658
rect 1575 2654 1581 2655
rect 1842 2651 1848 2652
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 278 2650 284 2651
rect 278 2646 279 2650
rect 283 2646 284 2650
rect 278 2645 284 2646
rect 446 2650 452 2651
rect 446 2646 447 2650
rect 451 2646 452 2650
rect 446 2645 452 2646
rect 622 2650 628 2651
rect 622 2646 623 2650
rect 627 2646 628 2650
rect 622 2645 628 2646
rect 790 2650 796 2651
rect 790 2646 791 2650
rect 795 2646 796 2650
rect 790 2645 796 2646
rect 950 2650 956 2651
rect 950 2646 951 2650
rect 955 2646 956 2650
rect 950 2645 956 2646
rect 1102 2650 1108 2651
rect 1102 2646 1103 2650
rect 1107 2646 1108 2650
rect 1102 2645 1108 2646
rect 1246 2650 1252 2651
rect 1246 2646 1247 2650
rect 1251 2646 1252 2650
rect 1246 2645 1252 2646
rect 1398 2650 1404 2651
rect 1398 2646 1399 2650
rect 1403 2646 1404 2650
rect 1398 2645 1404 2646
rect 1550 2650 1556 2651
rect 1550 2646 1551 2650
rect 1555 2646 1556 2650
rect 1842 2647 1843 2651
rect 1847 2650 1848 2651
rect 1927 2651 1933 2652
rect 1927 2650 1928 2651
rect 1847 2648 1928 2650
rect 1847 2647 1848 2648
rect 1842 2646 1848 2647
rect 1927 2647 1928 2648
rect 1932 2647 1933 2651
rect 1927 2646 1933 2647
rect 2095 2651 2101 2652
rect 2095 2647 2096 2651
rect 2100 2650 2101 2651
rect 2135 2651 2141 2652
rect 2135 2650 2136 2651
rect 2100 2648 2136 2650
rect 2100 2647 2101 2648
rect 2095 2646 2101 2647
rect 2135 2647 2136 2648
rect 2140 2647 2141 2651
rect 2135 2646 2141 2647
rect 2358 2651 2365 2652
rect 2358 2647 2359 2651
rect 2364 2647 2365 2651
rect 2358 2646 2365 2647
rect 2454 2651 2460 2652
rect 2454 2647 2455 2651
rect 2459 2650 2460 2651
rect 2567 2651 2573 2652
rect 2567 2650 2568 2651
rect 2459 2648 2568 2650
rect 2459 2647 2460 2648
rect 2454 2646 2460 2647
rect 2567 2647 2568 2648
rect 2572 2647 2573 2651
rect 2567 2646 2573 2647
rect 2767 2651 2776 2652
rect 2767 2647 2768 2651
rect 2775 2647 2776 2651
rect 2767 2646 2776 2647
rect 2903 2651 2909 2652
rect 2903 2647 2904 2651
rect 2908 2650 2909 2651
rect 2943 2651 2949 2652
rect 2943 2650 2944 2651
rect 2908 2648 2944 2650
rect 2908 2647 2909 2648
rect 2903 2646 2909 2647
rect 2943 2647 2944 2648
rect 2948 2647 2949 2651
rect 2943 2646 2949 2647
rect 3014 2651 3020 2652
rect 3014 2647 3015 2651
rect 3019 2650 3020 2651
rect 3103 2651 3109 2652
rect 3103 2650 3104 2651
rect 3019 2648 3104 2650
rect 3019 2647 3020 2648
rect 3014 2646 3020 2647
rect 3103 2647 3104 2648
rect 3108 2647 3109 2651
rect 3103 2646 3109 2647
rect 3170 2651 3176 2652
rect 3170 2647 3171 2651
rect 3175 2650 3176 2651
rect 3255 2651 3261 2652
rect 3255 2650 3256 2651
rect 3175 2648 3256 2650
rect 3175 2647 3176 2648
rect 3170 2646 3176 2647
rect 3255 2647 3256 2648
rect 3260 2647 3261 2651
rect 3255 2646 3261 2647
rect 3322 2651 3328 2652
rect 3322 2647 3323 2651
rect 3327 2650 3328 2651
rect 3407 2651 3413 2652
rect 3407 2650 3408 2651
rect 3327 2648 3408 2650
rect 3327 2647 3328 2648
rect 3322 2646 3328 2647
rect 3407 2647 3408 2648
rect 3412 2647 3413 2651
rect 3407 2646 3413 2647
rect 3534 2651 3541 2652
rect 3534 2647 3535 2651
rect 3540 2647 3541 2651
rect 3534 2646 3541 2647
rect 1550 2645 1556 2646
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 1927 2631 1936 2632
rect 1927 2627 1928 2631
rect 1935 2627 1936 2631
rect 1927 2626 1936 2627
rect 1954 2631 1960 2632
rect 1954 2627 1955 2631
rect 1959 2630 1960 2631
rect 2079 2631 2085 2632
rect 2079 2630 2080 2631
rect 1959 2628 2080 2630
rect 1959 2627 1960 2628
rect 1954 2626 1960 2627
rect 2079 2627 2080 2628
rect 2084 2627 2085 2631
rect 2079 2626 2085 2627
rect 2254 2631 2260 2632
rect 2254 2627 2255 2631
rect 2259 2630 2260 2631
rect 2287 2631 2293 2632
rect 2287 2630 2288 2631
rect 2259 2628 2288 2630
rect 2259 2627 2260 2628
rect 2254 2626 2260 2627
rect 2287 2627 2288 2628
rect 2292 2627 2293 2631
rect 2287 2626 2293 2627
rect 2314 2631 2320 2632
rect 2314 2627 2315 2631
rect 2319 2630 2320 2631
rect 2519 2631 2525 2632
rect 2519 2630 2520 2631
rect 2319 2628 2520 2630
rect 2319 2627 2320 2628
rect 2314 2626 2320 2627
rect 2519 2627 2520 2628
rect 2524 2627 2525 2631
rect 2519 2626 2525 2627
rect 2671 2631 2677 2632
rect 2671 2627 2672 2631
rect 2676 2630 2677 2631
rect 2775 2631 2781 2632
rect 2775 2630 2776 2631
rect 2676 2628 2776 2630
rect 2676 2627 2677 2628
rect 2671 2626 2677 2627
rect 2775 2627 2776 2628
rect 2780 2627 2781 2631
rect 2775 2626 2781 2627
rect 3039 2631 3045 2632
rect 3039 2627 3040 2631
rect 3044 2630 3045 2631
rect 3294 2631 3300 2632
rect 3294 2630 3295 2631
rect 3044 2628 3295 2630
rect 3044 2627 3045 2628
rect 3039 2626 3045 2627
rect 3294 2627 3295 2628
rect 3299 2627 3300 2631
rect 3294 2626 3300 2627
rect 3302 2631 3308 2632
rect 3302 2627 3303 2631
rect 3307 2630 3308 2631
rect 3311 2631 3317 2632
rect 3311 2630 3312 2631
rect 3307 2628 3312 2630
rect 3307 2627 3308 2628
rect 3302 2626 3308 2627
rect 3311 2627 3312 2628
rect 3316 2627 3317 2631
rect 3311 2626 3317 2627
rect 239 2623 245 2624
rect 239 2622 240 2623
rect 197 2620 240 2622
rect 239 2619 240 2620
rect 244 2619 245 2623
rect 239 2618 245 2619
rect 330 2623 336 2624
rect 330 2619 331 2623
rect 335 2619 336 2623
rect 735 2623 741 2624
rect 735 2622 736 2623
rect 677 2620 736 2622
rect 330 2618 336 2619
rect 735 2619 736 2620
rect 740 2619 741 2623
rect 735 2618 741 2619
rect 842 2623 848 2624
rect 842 2619 843 2623
rect 847 2619 848 2623
rect 842 2618 848 2619
rect 1002 2623 1008 2624
rect 1002 2619 1003 2623
rect 1007 2619 1008 2623
rect 1002 2618 1008 2619
rect 1154 2623 1160 2624
rect 1154 2619 1155 2623
rect 1159 2619 1160 2623
rect 1390 2623 1396 2624
rect 1390 2622 1391 2623
rect 1301 2620 1391 2622
rect 1154 2618 1160 2619
rect 1390 2619 1391 2620
rect 1395 2619 1396 2623
rect 1542 2623 1548 2624
rect 1542 2622 1543 2623
rect 1453 2620 1543 2622
rect 1390 2618 1396 2619
rect 1542 2619 1543 2620
rect 1547 2619 1548 2623
rect 1542 2618 1548 2619
rect 1558 2623 1564 2624
rect 1558 2619 1559 2623
rect 1563 2619 1564 2623
rect 1558 2618 1564 2619
rect 1902 2622 1908 2623
rect 1902 2618 1903 2622
rect 1907 2618 1908 2622
rect 1902 2617 1908 2618
rect 2054 2622 2060 2623
rect 2054 2618 2055 2622
rect 2059 2618 2060 2622
rect 2054 2617 2060 2618
rect 2262 2622 2268 2623
rect 2262 2618 2263 2622
rect 2267 2618 2268 2622
rect 2262 2617 2268 2618
rect 2494 2622 2500 2623
rect 2494 2618 2495 2622
rect 2499 2618 2500 2622
rect 2494 2617 2500 2618
rect 2750 2622 2756 2623
rect 2750 2618 2751 2622
rect 2755 2618 2756 2622
rect 2750 2617 2756 2618
rect 3014 2622 3020 2623
rect 3014 2618 3015 2622
rect 3019 2618 3020 2622
rect 3014 2617 3020 2618
rect 3286 2622 3292 2623
rect 3286 2618 3287 2622
rect 3291 2618 3292 2622
rect 3286 2617 3292 2618
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 1830 2615 1836 2616
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 270 2612 276 2613
rect 270 2608 271 2612
rect 275 2608 276 2612
rect 270 2607 276 2608
rect 438 2612 444 2613
rect 438 2608 439 2612
rect 443 2608 444 2612
rect 438 2607 444 2608
rect 614 2612 620 2613
rect 614 2608 615 2612
rect 619 2608 620 2612
rect 614 2607 620 2608
rect 782 2612 788 2613
rect 782 2608 783 2612
rect 787 2608 788 2612
rect 782 2607 788 2608
rect 942 2612 948 2613
rect 942 2608 943 2612
rect 947 2608 948 2612
rect 942 2607 948 2608
rect 1094 2612 1100 2613
rect 1094 2608 1095 2612
rect 1099 2608 1100 2612
rect 1094 2607 1100 2608
rect 1238 2612 1244 2613
rect 1238 2608 1239 2612
rect 1243 2608 1244 2612
rect 1238 2607 1244 2608
rect 1390 2612 1396 2613
rect 1390 2608 1391 2612
rect 1395 2608 1396 2612
rect 1390 2607 1396 2608
rect 1542 2612 1548 2613
rect 1542 2608 1543 2612
rect 1547 2608 1548 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1542 2607 1548 2608
rect 1870 2604 1876 2605
rect 1870 2600 1871 2604
rect 1875 2600 1876 2604
rect 1870 2599 1876 2600
rect 3590 2604 3596 2605
rect 3590 2600 3591 2604
rect 3595 2600 3596 2604
rect 3590 2599 3596 2600
rect 402 2595 408 2596
rect 402 2591 403 2595
rect 407 2594 408 2595
rect 455 2595 461 2596
rect 455 2594 456 2595
rect 407 2592 456 2594
rect 407 2591 408 2592
rect 402 2590 408 2591
rect 455 2591 456 2592
rect 460 2591 461 2595
rect 455 2590 461 2591
rect 1954 2595 1960 2596
rect 1954 2591 1955 2595
rect 1959 2591 1960 2595
rect 2254 2595 2260 2596
rect 2254 2594 2255 2595
rect 2109 2592 2255 2594
rect 1954 2590 1960 2591
rect 2254 2591 2255 2592
rect 2259 2591 2260 2595
rect 2254 2590 2260 2591
rect 2314 2595 2320 2596
rect 2314 2591 2315 2595
rect 2319 2591 2320 2595
rect 2671 2595 2677 2596
rect 2671 2594 2672 2595
rect 2549 2592 2672 2594
rect 2314 2590 2320 2591
rect 2671 2591 2672 2592
rect 2676 2591 2677 2595
rect 2671 2590 2677 2591
rect 3038 2595 3044 2596
rect 3038 2591 3039 2595
rect 3043 2591 3044 2595
rect 3038 2590 3044 2591
rect 3294 2595 3300 2596
rect 3294 2591 3295 2595
rect 3299 2591 3300 2595
rect 3294 2590 3300 2591
rect 1870 2587 1876 2588
rect 1870 2583 1871 2587
rect 1875 2583 1876 2587
rect 3590 2587 3596 2588
rect 1870 2582 1876 2583
rect 1894 2584 1900 2585
rect 1894 2580 1895 2584
rect 1899 2580 1900 2584
rect 1894 2579 1900 2580
rect 2046 2584 2052 2585
rect 2046 2580 2047 2584
rect 2051 2580 2052 2584
rect 2046 2579 2052 2580
rect 2254 2584 2260 2585
rect 2254 2580 2255 2584
rect 2259 2580 2260 2584
rect 2254 2579 2260 2580
rect 2486 2584 2492 2585
rect 2486 2580 2487 2584
rect 2491 2580 2492 2584
rect 2486 2579 2492 2580
rect 2742 2584 2748 2585
rect 2742 2580 2743 2584
rect 2747 2580 2748 2584
rect 2742 2579 2748 2580
rect 3006 2584 3012 2585
rect 3006 2580 3007 2584
rect 3011 2580 3012 2584
rect 3006 2579 3012 2580
rect 3278 2584 3284 2585
rect 3278 2580 3279 2584
rect 3283 2580 3284 2584
rect 3590 2583 3591 2587
rect 3595 2583 3596 2587
rect 3590 2582 3596 2583
rect 3278 2579 3284 2580
rect 2658 2567 2664 2568
rect 134 2564 140 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 134 2560 135 2564
rect 139 2560 140 2564
rect 134 2559 140 2560
rect 222 2564 228 2565
rect 222 2560 223 2564
rect 227 2560 228 2564
rect 222 2559 228 2560
rect 366 2564 372 2565
rect 366 2560 367 2564
rect 371 2560 372 2564
rect 366 2559 372 2560
rect 526 2564 532 2565
rect 526 2560 527 2564
rect 531 2560 532 2564
rect 526 2559 532 2560
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 878 2564 884 2565
rect 878 2560 879 2564
rect 883 2560 884 2564
rect 878 2559 884 2560
rect 1046 2564 1052 2565
rect 1046 2560 1047 2564
rect 1051 2560 1052 2564
rect 1046 2559 1052 2560
rect 1206 2564 1212 2565
rect 1206 2560 1207 2564
rect 1211 2560 1212 2564
rect 1206 2559 1212 2560
rect 1358 2564 1364 2565
rect 1358 2560 1359 2564
rect 1363 2560 1364 2564
rect 1358 2559 1364 2560
rect 1510 2564 1516 2565
rect 1510 2560 1511 2564
rect 1515 2560 1516 2564
rect 1510 2559 1516 2560
rect 1670 2564 1676 2565
rect 1670 2560 1671 2564
rect 1675 2560 1676 2564
rect 2658 2563 2659 2567
rect 2663 2566 2664 2567
rect 2759 2567 2765 2568
rect 2759 2566 2760 2567
rect 2663 2564 2760 2566
rect 2663 2563 2664 2564
rect 2658 2562 2664 2563
rect 2759 2563 2760 2564
rect 2764 2563 2765 2567
rect 2759 2562 2765 2563
rect 1670 2559 1676 2560
rect 1830 2561 1836 2562
rect 110 2556 116 2557
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1830 2556 1836 2557
rect 202 2555 208 2556
rect 196 2548 198 2553
rect 202 2551 203 2555
rect 207 2554 208 2555
rect 290 2555 296 2556
rect 207 2552 241 2554
rect 207 2551 208 2552
rect 202 2550 208 2551
rect 290 2551 291 2555
rect 295 2554 296 2555
rect 594 2555 600 2556
rect 295 2552 385 2554
rect 295 2551 296 2552
rect 290 2550 296 2551
rect 588 2548 590 2553
rect 594 2551 595 2555
rect 599 2554 600 2555
rect 770 2555 776 2556
rect 599 2552 721 2554
rect 599 2551 600 2552
rect 594 2550 600 2551
rect 770 2551 771 2555
rect 775 2554 776 2555
rect 990 2555 996 2556
rect 775 2552 897 2554
rect 775 2551 776 2552
rect 770 2550 776 2551
rect 990 2551 991 2555
rect 995 2554 996 2555
rect 1114 2555 1120 2556
rect 995 2552 1065 2554
rect 995 2551 996 2552
rect 990 2550 996 2551
rect 1114 2551 1115 2555
rect 1119 2554 1120 2555
rect 1274 2555 1280 2556
rect 1119 2552 1225 2554
rect 1119 2551 1120 2552
rect 1114 2550 1120 2551
rect 1274 2551 1275 2555
rect 1279 2554 1280 2555
rect 1426 2555 1432 2556
rect 1279 2552 1377 2554
rect 1279 2551 1280 2552
rect 1274 2550 1280 2551
rect 1426 2551 1427 2555
rect 1431 2554 1432 2555
rect 1578 2555 1584 2556
rect 1431 2552 1529 2554
rect 1431 2551 1432 2552
rect 1426 2550 1432 2551
rect 1578 2551 1579 2555
rect 1583 2554 1584 2555
rect 1583 2552 1689 2554
rect 1583 2551 1584 2552
rect 1578 2550 1584 2551
rect 194 2547 200 2548
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 194 2543 195 2547
rect 199 2543 200 2547
rect 194 2542 200 2543
rect 586 2547 592 2548
rect 586 2543 587 2547
rect 591 2543 592 2547
rect 586 2542 592 2543
rect 1830 2544 1836 2545
rect 110 2539 116 2540
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 1894 2540 1900 2541
rect 1870 2537 1876 2538
rect 1870 2533 1871 2537
rect 1875 2533 1876 2537
rect 1894 2536 1895 2540
rect 1899 2536 1900 2540
rect 1894 2535 1900 2536
rect 2006 2540 2012 2541
rect 2006 2536 2007 2540
rect 2011 2536 2012 2540
rect 2006 2535 2012 2536
rect 2158 2540 2164 2541
rect 2158 2536 2159 2540
rect 2163 2536 2164 2540
rect 2158 2535 2164 2536
rect 2318 2540 2324 2541
rect 2318 2536 2319 2540
rect 2323 2536 2324 2540
rect 2318 2535 2324 2536
rect 2470 2540 2476 2541
rect 2470 2536 2471 2540
rect 2475 2536 2476 2540
rect 2470 2535 2476 2536
rect 2622 2540 2628 2541
rect 2622 2536 2623 2540
rect 2627 2536 2628 2540
rect 2622 2535 2628 2536
rect 2758 2540 2764 2541
rect 2758 2536 2759 2540
rect 2763 2536 2764 2540
rect 2758 2535 2764 2536
rect 2886 2540 2892 2541
rect 2886 2536 2887 2540
rect 2891 2536 2892 2540
rect 2886 2535 2892 2536
rect 3006 2540 3012 2541
rect 3006 2536 3007 2540
rect 3011 2536 3012 2540
rect 3006 2535 3012 2536
rect 3118 2540 3124 2541
rect 3118 2536 3119 2540
rect 3123 2536 3124 2540
rect 3118 2535 3124 2536
rect 3222 2540 3228 2541
rect 3222 2536 3223 2540
rect 3227 2536 3228 2540
rect 3222 2535 3228 2536
rect 3318 2540 3324 2541
rect 3318 2536 3319 2540
rect 3323 2536 3324 2540
rect 3318 2535 3324 2536
rect 3422 2540 3428 2541
rect 3422 2536 3423 2540
rect 3427 2536 3428 2540
rect 3422 2535 3428 2536
rect 3502 2540 3508 2541
rect 3502 2536 3503 2540
rect 3507 2536 3508 2540
rect 3502 2535 3508 2536
rect 3590 2537 3596 2538
rect 1870 2532 1876 2533
rect 3590 2533 3591 2537
rect 3595 2533 3596 2537
rect 3590 2532 3596 2533
rect 1962 2531 1968 2532
rect 1962 2530 1963 2531
rect 1957 2528 1963 2530
rect 1962 2527 1963 2528
rect 1967 2527 1968 2531
rect 2106 2531 2112 2532
rect 2106 2530 2107 2531
rect 2069 2528 2107 2530
rect 142 2526 148 2527
rect 142 2522 143 2526
rect 147 2522 148 2526
rect 142 2521 148 2522
rect 230 2526 236 2527
rect 230 2522 231 2526
rect 235 2522 236 2526
rect 230 2521 236 2522
rect 374 2526 380 2527
rect 374 2522 375 2526
rect 379 2522 380 2526
rect 374 2521 380 2522
rect 534 2526 540 2527
rect 534 2522 535 2526
rect 539 2522 540 2526
rect 534 2521 540 2522
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 886 2526 892 2527
rect 886 2522 887 2526
rect 891 2522 892 2526
rect 886 2521 892 2522
rect 1054 2526 1060 2527
rect 1054 2522 1055 2526
rect 1059 2522 1060 2526
rect 1054 2521 1060 2522
rect 1214 2526 1220 2527
rect 1214 2522 1215 2526
rect 1219 2522 1220 2526
rect 1214 2521 1220 2522
rect 1366 2526 1372 2527
rect 1366 2522 1367 2526
rect 1371 2522 1372 2526
rect 1366 2521 1372 2522
rect 1518 2526 1524 2527
rect 1518 2522 1519 2526
rect 1523 2522 1524 2526
rect 1518 2521 1524 2522
rect 1678 2526 1684 2527
rect 1962 2526 1968 2527
rect 2106 2527 2107 2528
rect 2111 2527 2112 2531
rect 2262 2531 2268 2532
rect 2262 2530 2263 2531
rect 2221 2528 2263 2530
rect 2106 2526 2112 2527
rect 2262 2527 2263 2528
rect 2267 2527 2268 2531
rect 2418 2531 2424 2532
rect 2418 2530 2419 2531
rect 2381 2528 2419 2530
rect 2262 2526 2268 2527
rect 2418 2527 2419 2528
rect 2423 2527 2424 2531
rect 2418 2526 2424 2527
rect 2426 2531 2432 2532
rect 2426 2527 2427 2531
rect 2431 2530 2432 2531
rect 2714 2531 2720 2532
rect 2714 2530 2715 2531
rect 2431 2528 2489 2530
rect 2685 2528 2715 2530
rect 2431 2527 2432 2528
rect 2426 2526 2432 2527
rect 2714 2527 2715 2528
rect 2719 2527 2720 2531
rect 2879 2531 2885 2532
rect 2879 2530 2880 2531
rect 2821 2528 2880 2530
rect 2714 2526 2720 2527
rect 2879 2527 2880 2528
rect 2884 2527 2885 2531
rect 2954 2531 2960 2532
rect 2879 2526 2885 2527
rect 1678 2522 1679 2526
rect 1683 2522 1684 2526
rect 1678 2521 1684 2522
rect 2682 2523 2688 2524
rect 1870 2520 1876 2521
rect 1870 2516 1871 2520
rect 1875 2516 1876 2520
rect 2682 2519 2683 2523
rect 2687 2522 2688 2523
rect 2904 2522 2906 2529
rect 2954 2527 2955 2531
rect 2959 2530 2960 2531
rect 3074 2531 3080 2532
rect 2959 2528 3025 2530
rect 2959 2527 2960 2528
rect 2954 2526 2960 2527
rect 3074 2527 3075 2531
rect 3079 2530 3080 2531
rect 3290 2531 3296 2532
rect 3079 2528 3137 2530
rect 3079 2527 3080 2528
rect 3074 2526 3080 2527
rect 2687 2520 2906 2522
rect 3284 2522 3286 2529
rect 3290 2527 3291 2531
rect 3295 2530 3296 2531
rect 3386 2531 3392 2532
rect 3295 2528 3337 2530
rect 3295 2527 3296 2528
rect 3290 2526 3296 2527
rect 3386 2527 3387 2531
rect 3391 2530 3392 2531
rect 3391 2528 3441 2530
rect 3391 2527 3392 2528
rect 3386 2526 3392 2527
rect 3564 2524 3566 2529
rect 3302 2523 3308 2524
rect 3302 2522 3303 2523
rect 3284 2520 3303 2522
rect 2687 2519 2688 2520
rect 2682 2518 2688 2519
rect 3302 2519 3303 2520
rect 3307 2519 3308 2523
rect 3302 2518 3308 2519
rect 3562 2523 3568 2524
rect 3562 2519 3563 2523
rect 3567 2519 3568 2523
rect 3562 2518 3568 2519
rect 3590 2520 3596 2521
rect 167 2515 173 2516
rect 167 2511 168 2515
rect 172 2514 173 2515
rect 202 2515 208 2516
rect 202 2514 203 2515
rect 172 2512 203 2514
rect 172 2511 173 2512
rect 167 2510 173 2511
rect 202 2511 203 2512
rect 207 2511 208 2515
rect 202 2510 208 2511
rect 255 2515 261 2516
rect 255 2511 256 2515
rect 260 2514 261 2515
rect 290 2515 296 2516
rect 290 2514 291 2515
rect 260 2512 291 2514
rect 260 2511 261 2512
rect 255 2510 261 2511
rect 290 2511 291 2512
rect 295 2511 296 2515
rect 290 2510 296 2511
rect 399 2515 408 2516
rect 399 2511 400 2515
rect 407 2511 408 2515
rect 399 2510 408 2511
rect 559 2515 565 2516
rect 559 2511 560 2515
rect 564 2514 565 2515
rect 594 2515 600 2516
rect 594 2514 595 2515
rect 564 2512 595 2514
rect 564 2511 565 2512
rect 559 2510 565 2511
rect 594 2511 595 2512
rect 599 2511 600 2515
rect 594 2510 600 2511
rect 735 2515 741 2516
rect 735 2511 736 2515
rect 740 2514 741 2515
rect 770 2515 776 2516
rect 770 2514 771 2515
rect 740 2512 771 2514
rect 740 2511 741 2512
rect 735 2510 741 2511
rect 770 2511 771 2512
rect 775 2511 776 2515
rect 770 2510 776 2511
rect 911 2515 917 2516
rect 911 2511 912 2515
rect 916 2514 917 2515
rect 934 2515 940 2516
rect 934 2514 935 2515
rect 916 2512 935 2514
rect 916 2511 917 2512
rect 911 2510 917 2511
rect 934 2511 935 2512
rect 939 2511 940 2515
rect 934 2510 940 2511
rect 1079 2515 1085 2516
rect 1079 2511 1080 2515
rect 1084 2514 1085 2515
rect 1114 2515 1120 2516
rect 1114 2514 1115 2515
rect 1084 2512 1115 2514
rect 1084 2511 1085 2512
rect 1079 2510 1085 2511
rect 1114 2511 1115 2512
rect 1119 2511 1120 2515
rect 1114 2510 1120 2511
rect 1239 2515 1245 2516
rect 1239 2511 1240 2515
rect 1244 2514 1245 2515
rect 1274 2515 1280 2516
rect 1274 2514 1275 2515
rect 1244 2512 1275 2514
rect 1244 2511 1245 2512
rect 1239 2510 1245 2511
rect 1274 2511 1275 2512
rect 1279 2511 1280 2515
rect 1274 2510 1280 2511
rect 1391 2515 1397 2516
rect 1391 2511 1392 2515
rect 1396 2514 1397 2515
rect 1426 2515 1432 2516
rect 1426 2514 1427 2515
rect 1396 2512 1427 2514
rect 1396 2511 1397 2512
rect 1391 2510 1397 2511
rect 1426 2511 1427 2512
rect 1431 2511 1432 2515
rect 1426 2510 1432 2511
rect 1543 2515 1549 2516
rect 1543 2511 1544 2515
rect 1548 2514 1549 2515
rect 1578 2515 1584 2516
rect 1578 2514 1579 2515
rect 1548 2512 1579 2514
rect 1548 2511 1549 2512
rect 1543 2510 1549 2511
rect 1578 2511 1579 2512
rect 1583 2511 1584 2515
rect 1578 2510 1584 2511
rect 1702 2515 1709 2516
rect 1870 2515 1876 2516
rect 3590 2516 3591 2520
rect 3595 2516 3596 2520
rect 3590 2515 3596 2516
rect 1702 2511 1703 2515
rect 1708 2511 1709 2515
rect 1702 2510 1709 2511
rect 1902 2502 1908 2503
rect 167 2499 173 2500
rect 167 2495 168 2499
rect 172 2498 173 2499
rect 194 2499 200 2500
rect 194 2498 195 2499
rect 172 2496 195 2498
rect 172 2495 173 2496
rect 167 2494 173 2495
rect 194 2495 195 2496
rect 199 2495 200 2499
rect 194 2494 200 2495
rect 214 2499 220 2500
rect 214 2495 215 2499
rect 219 2498 220 2499
rect 247 2499 253 2500
rect 247 2498 248 2499
rect 219 2496 248 2498
rect 219 2495 220 2496
rect 214 2494 220 2495
rect 247 2495 248 2496
rect 252 2495 253 2499
rect 247 2494 253 2495
rect 274 2499 280 2500
rect 274 2495 275 2499
rect 279 2498 280 2499
rect 327 2499 333 2500
rect 327 2498 328 2499
rect 279 2496 328 2498
rect 279 2495 280 2496
rect 274 2494 280 2495
rect 327 2495 328 2496
rect 332 2495 333 2499
rect 327 2494 333 2495
rect 354 2499 360 2500
rect 354 2495 355 2499
rect 359 2498 360 2499
rect 415 2499 421 2500
rect 415 2498 416 2499
rect 359 2496 416 2498
rect 359 2495 360 2496
rect 354 2494 360 2495
rect 415 2495 416 2496
rect 420 2495 421 2499
rect 415 2494 421 2495
rect 442 2499 448 2500
rect 442 2495 443 2499
rect 447 2498 448 2499
rect 535 2499 541 2500
rect 535 2498 536 2499
rect 447 2496 536 2498
rect 447 2495 448 2496
rect 442 2494 448 2495
rect 535 2495 536 2496
rect 540 2495 541 2499
rect 535 2494 541 2495
rect 562 2499 568 2500
rect 562 2495 563 2499
rect 567 2498 568 2499
rect 671 2499 677 2500
rect 671 2498 672 2499
rect 567 2496 672 2498
rect 567 2495 568 2496
rect 562 2494 568 2495
rect 671 2495 672 2496
rect 676 2495 677 2499
rect 671 2494 677 2495
rect 698 2499 704 2500
rect 698 2495 699 2499
rect 703 2498 704 2499
rect 807 2499 813 2500
rect 807 2498 808 2499
rect 703 2496 808 2498
rect 703 2495 704 2496
rect 698 2494 704 2495
rect 807 2495 808 2496
rect 812 2495 813 2499
rect 807 2494 813 2495
rect 834 2499 840 2500
rect 834 2495 835 2499
rect 839 2498 840 2499
rect 951 2499 957 2500
rect 951 2498 952 2499
rect 839 2496 952 2498
rect 839 2495 840 2496
rect 834 2494 840 2495
rect 951 2495 952 2496
rect 956 2495 957 2499
rect 951 2494 957 2495
rect 1087 2499 1093 2500
rect 1087 2495 1088 2499
rect 1092 2498 1093 2499
rect 1134 2499 1140 2500
rect 1134 2498 1135 2499
rect 1092 2496 1135 2498
rect 1092 2495 1093 2496
rect 1087 2494 1093 2495
rect 1134 2495 1135 2496
rect 1139 2495 1140 2499
rect 1134 2494 1140 2495
rect 1142 2499 1148 2500
rect 1142 2495 1143 2499
rect 1147 2498 1148 2499
rect 1215 2499 1221 2500
rect 1215 2498 1216 2499
rect 1147 2496 1216 2498
rect 1147 2495 1148 2496
rect 1142 2494 1148 2495
rect 1215 2495 1216 2496
rect 1220 2495 1221 2499
rect 1215 2494 1221 2495
rect 1242 2499 1248 2500
rect 1242 2495 1243 2499
rect 1247 2498 1248 2499
rect 1335 2499 1341 2500
rect 1335 2498 1336 2499
rect 1247 2496 1336 2498
rect 1247 2495 1248 2496
rect 1242 2494 1248 2495
rect 1335 2495 1336 2496
rect 1340 2495 1341 2499
rect 1335 2494 1341 2495
rect 1422 2499 1428 2500
rect 1422 2495 1423 2499
rect 1427 2498 1428 2499
rect 1455 2499 1461 2500
rect 1455 2498 1456 2499
rect 1427 2496 1456 2498
rect 1427 2495 1428 2496
rect 1422 2494 1428 2495
rect 1455 2495 1456 2496
rect 1460 2495 1461 2499
rect 1455 2494 1461 2495
rect 1482 2499 1488 2500
rect 1482 2495 1483 2499
rect 1487 2498 1488 2499
rect 1575 2499 1581 2500
rect 1575 2498 1576 2499
rect 1487 2496 1576 2498
rect 1487 2495 1488 2496
rect 1482 2494 1488 2495
rect 1575 2495 1576 2496
rect 1580 2495 1581 2499
rect 1575 2494 1581 2495
rect 1602 2499 1608 2500
rect 1602 2495 1603 2499
rect 1607 2498 1608 2499
rect 1695 2499 1701 2500
rect 1695 2498 1696 2499
rect 1607 2496 1696 2498
rect 1607 2495 1608 2496
rect 1602 2494 1608 2495
rect 1695 2495 1696 2496
rect 1700 2495 1701 2499
rect 1902 2498 1903 2502
rect 1907 2498 1908 2502
rect 1902 2497 1908 2498
rect 2014 2502 2020 2503
rect 2014 2498 2015 2502
rect 2019 2498 2020 2502
rect 2014 2497 2020 2498
rect 2166 2502 2172 2503
rect 2166 2498 2167 2502
rect 2171 2498 2172 2502
rect 2166 2497 2172 2498
rect 2326 2502 2332 2503
rect 2326 2498 2327 2502
rect 2331 2498 2332 2502
rect 2326 2497 2332 2498
rect 2478 2502 2484 2503
rect 2478 2498 2479 2502
rect 2483 2498 2484 2502
rect 2478 2497 2484 2498
rect 2630 2502 2636 2503
rect 2630 2498 2631 2502
rect 2635 2498 2636 2502
rect 2630 2497 2636 2498
rect 2766 2502 2772 2503
rect 2766 2498 2767 2502
rect 2771 2498 2772 2502
rect 2766 2497 2772 2498
rect 2894 2502 2900 2503
rect 2894 2498 2895 2502
rect 2899 2498 2900 2502
rect 2894 2497 2900 2498
rect 3014 2502 3020 2503
rect 3014 2498 3015 2502
rect 3019 2498 3020 2502
rect 3014 2497 3020 2498
rect 3126 2502 3132 2503
rect 3126 2498 3127 2502
rect 3131 2498 3132 2502
rect 3126 2497 3132 2498
rect 3230 2502 3236 2503
rect 3230 2498 3231 2502
rect 3235 2498 3236 2502
rect 3230 2497 3236 2498
rect 3326 2502 3332 2503
rect 3326 2498 3327 2502
rect 3331 2498 3332 2502
rect 3326 2497 3332 2498
rect 3430 2502 3436 2503
rect 3430 2498 3431 2502
rect 3435 2498 3436 2502
rect 3430 2497 3436 2498
rect 3510 2502 3516 2503
rect 3510 2498 3511 2502
rect 3515 2498 3516 2502
rect 3510 2497 3516 2498
rect 1695 2494 1701 2495
rect 1927 2491 1936 2492
rect 142 2490 148 2491
rect 142 2486 143 2490
rect 147 2486 148 2490
rect 142 2485 148 2486
rect 222 2490 228 2491
rect 222 2486 223 2490
rect 227 2486 228 2490
rect 222 2485 228 2486
rect 302 2490 308 2491
rect 302 2486 303 2490
rect 307 2486 308 2490
rect 302 2485 308 2486
rect 390 2490 396 2491
rect 390 2486 391 2490
rect 395 2486 396 2490
rect 390 2485 396 2486
rect 510 2490 516 2491
rect 510 2486 511 2490
rect 515 2486 516 2490
rect 510 2485 516 2486
rect 646 2490 652 2491
rect 646 2486 647 2490
rect 651 2486 652 2490
rect 646 2485 652 2486
rect 782 2490 788 2491
rect 782 2486 783 2490
rect 787 2486 788 2490
rect 782 2485 788 2486
rect 926 2490 932 2491
rect 926 2486 927 2490
rect 931 2486 932 2490
rect 926 2485 932 2486
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1310 2490 1316 2491
rect 1310 2486 1311 2490
rect 1315 2486 1316 2490
rect 1310 2485 1316 2486
rect 1430 2490 1436 2491
rect 1430 2486 1431 2490
rect 1435 2486 1436 2490
rect 1430 2485 1436 2486
rect 1550 2490 1556 2491
rect 1550 2486 1551 2490
rect 1555 2486 1556 2490
rect 1550 2485 1556 2486
rect 1670 2490 1676 2491
rect 1670 2486 1671 2490
rect 1675 2486 1676 2490
rect 1927 2487 1928 2491
rect 1935 2487 1936 2491
rect 1927 2486 1936 2487
rect 1962 2491 1968 2492
rect 1962 2487 1963 2491
rect 1967 2490 1968 2491
rect 2039 2491 2045 2492
rect 2039 2490 2040 2491
rect 1967 2488 2040 2490
rect 1967 2487 1968 2488
rect 1962 2486 1968 2487
rect 2039 2487 2040 2488
rect 2044 2487 2045 2491
rect 2039 2486 2045 2487
rect 2106 2491 2112 2492
rect 2106 2487 2107 2491
rect 2111 2490 2112 2491
rect 2191 2491 2197 2492
rect 2191 2490 2192 2491
rect 2111 2488 2192 2490
rect 2111 2487 2112 2488
rect 2106 2486 2112 2487
rect 2191 2487 2192 2488
rect 2196 2487 2197 2491
rect 2191 2486 2197 2487
rect 2262 2491 2268 2492
rect 2262 2487 2263 2491
rect 2267 2490 2268 2491
rect 2351 2491 2357 2492
rect 2351 2490 2352 2491
rect 2267 2488 2352 2490
rect 2267 2487 2268 2488
rect 2262 2486 2268 2487
rect 2351 2487 2352 2488
rect 2356 2487 2357 2491
rect 2351 2486 2357 2487
rect 2418 2491 2424 2492
rect 2418 2487 2419 2491
rect 2423 2490 2424 2491
rect 2503 2491 2509 2492
rect 2503 2490 2504 2491
rect 2423 2488 2504 2490
rect 2423 2487 2424 2488
rect 2418 2486 2424 2487
rect 2503 2487 2504 2488
rect 2508 2487 2509 2491
rect 2503 2486 2509 2487
rect 2655 2491 2661 2492
rect 2655 2487 2656 2491
rect 2660 2490 2661 2491
rect 2682 2491 2688 2492
rect 2682 2490 2683 2491
rect 2660 2488 2683 2490
rect 2660 2487 2661 2488
rect 2655 2486 2661 2487
rect 2682 2487 2683 2488
rect 2687 2487 2688 2491
rect 2682 2486 2688 2487
rect 2714 2491 2720 2492
rect 2714 2487 2715 2491
rect 2719 2490 2720 2491
rect 2791 2491 2797 2492
rect 2791 2490 2792 2491
rect 2719 2488 2792 2490
rect 2719 2487 2720 2488
rect 2714 2486 2720 2487
rect 2791 2487 2792 2488
rect 2796 2487 2797 2491
rect 2791 2486 2797 2487
rect 2919 2491 2925 2492
rect 2919 2487 2920 2491
rect 2924 2490 2925 2491
rect 2954 2491 2960 2492
rect 2954 2490 2955 2491
rect 2924 2488 2955 2490
rect 2924 2487 2925 2488
rect 2919 2486 2925 2487
rect 2954 2487 2955 2488
rect 2959 2487 2960 2491
rect 2954 2486 2960 2487
rect 3038 2491 3045 2492
rect 3038 2487 3039 2491
rect 3044 2487 3045 2491
rect 3151 2491 3157 2492
rect 3151 2490 3152 2491
rect 3038 2486 3045 2487
rect 3048 2488 3152 2490
rect 1670 2485 1676 2486
rect 2879 2483 2885 2484
rect 2426 2479 2432 2480
rect 2426 2478 2427 2479
rect 2044 2476 2427 2478
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 2023 2471 2029 2472
rect 2023 2467 2024 2471
rect 2028 2470 2029 2471
rect 2044 2470 2046 2476
rect 2426 2475 2427 2476
rect 2431 2475 2432 2479
rect 2879 2479 2880 2483
rect 2884 2482 2885 2483
rect 3048 2482 3050 2488
rect 3151 2487 3152 2488
rect 3156 2487 3157 2491
rect 3151 2486 3157 2487
rect 3255 2491 3261 2492
rect 3255 2487 3256 2491
rect 3260 2490 3261 2491
rect 3290 2491 3296 2492
rect 3290 2490 3291 2491
rect 3260 2488 3291 2490
rect 3260 2487 3261 2488
rect 3255 2486 3261 2487
rect 3290 2487 3291 2488
rect 3295 2487 3296 2491
rect 3290 2486 3296 2487
rect 3351 2491 3357 2492
rect 3351 2487 3352 2491
rect 3356 2490 3357 2491
rect 3386 2491 3392 2492
rect 3386 2490 3387 2491
rect 3356 2488 3387 2490
rect 3356 2487 3357 2488
rect 3351 2486 3357 2487
rect 3386 2487 3387 2488
rect 3391 2487 3392 2491
rect 3386 2486 3392 2487
rect 3410 2491 3416 2492
rect 3410 2487 3411 2491
rect 3415 2490 3416 2491
rect 3455 2491 3461 2492
rect 3455 2490 3456 2491
rect 3415 2488 3456 2490
rect 3415 2487 3416 2488
rect 3410 2486 3416 2487
rect 3455 2487 3456 2488
rect 3460 2487 3461 2491
rect 3455 2486 3461 2487
rect 3535 2491 3541 2492
rect 3535 2487 3536 2491
rect 3540 2490 3541 2491
rect 3570 2491 3576 2492
rect 3570 2490 3571 2491
rect 3540 2488 3571 2490
rect 3540 2487 3541 2488
rect 3535 2486 3541 2487
rect 3570 2487 3571 2488
rect 3575 2487 3576 2491
rect 3570 2486 3576 2487
rect 2884 2480 3050 2482
rect 2884 2479 2885 2480
rect 2879 2478 2885 2479
rect 2426 2474 2432 2475
rect 2028 2468 2046 2470
rect 2050 2471 2056 2472
rect 2028 2467 2029 2468
rect 2023 2466 2029 2467
rect 2050 2467 2051 2471
rect 2055 2470 2056 2471
rect 2151 2471 2157 2472
rect 2151 2470 2152 2471
rect 2055 2468 2152 2470
rect 2055 2467 2056 2468
rect 2050 2466 2056 2467
rect 2151 2467 2152 2468
rect 2156 2467 2157 2471
rect 2151 2466 2157 2467
rect 2178 2471 2184 2472
rect 2178 2467 2179 2471
rect 2183 2470 2184 2471
rect 2287 2471 2293 2472
rect 2287 2470 2288 2471
rect 2183 2468 2288 2470
rect 2183 2467 2184 2468
rect 2178 2466 2184 2467
rect 2287 2467 2288 2468
rect 2292 2467 2293 2471
rect 2287 2466 2293 2467
rect 2314 2471 2320 2472
rect 2314 2467 2315 2471
rect 2319 2470 2320 2471
rect 2431 2471 2437 2472
rect 2431 2470 2432 2471
rect 2319 2468 2432 2470
rect 2319 2467 2320 2468
rect 2314 2466 2320 2467
rect 2431 2467 2432 2468
rect 2436 2467 2437 2471
rect 2431 2466 2437 2467
rect 2458 2471 2464 2472
rect 2458 2467 2459 2471
rect 2463 2470 2464 2471
rect 2575 2471 2581 2472
rect 2575 2470 2576 2471
rect 2463 2468 2576 2470
rect 2463 2467 2464 2468
rect 2458 2466 2464 2467
rect 2575 2467 2576 2468
rect 2580 2467 2581 2471
rect 2575 2466 2581 2467
rect 2727 2471 2733 2472
rect 2727 2467 2728 2471
rect 2732 2470 2733 2471
rect 2802 2471 2808 2472
rect 2802 2470 2803 2471
rect 2732 2468 2803 2470
rect 2732 2467 2733 2468
rect 2727 2466 2733 2467
rect 2802 2467 2803 2468
rect 2807 2467 2808 2471
rect 2802 2466 2808 2467
rect 2810 2471 2816 2472
rect 2810 2467 2811 2471
rect 2815 2470 2816 2471
rect 2887 2471 2893 2472
rect 2887 2470 2888 2471
rect 2815 2468 2888 2470
rect 2815 2467 2816 2468
rect 2810 2466 2816 2467
rect 2887 2467 2888 2468
rect 2892 2467 2893 2471
rect 2887 2466 2893 2467
rect 3047 2471 3053 2472
rect 3047 2467 3048 2471
rect 3052 2470 3053 2471
rect 3074 2471 3080 2472
rect 3074 2470 3075 2471
rect 3052 2468 3075 2470
rect 3052 2467 3053 2468
rect 3047 2466 3053 2467
rect 3074 2467 3075 2468
rect 3079 2467 3080 2471
rect 3074 2466 3080 2467
rect 3127 2471 3133 2472
rect 3127 2467 3128 2471
rect 3132 2470 3133 2471
rect 3215 2471 3221 2472
rect 3215 2470 3216 2471
rect 3132 2468 3216 2470
rect 3132 2467 3133 2468
rect 3127 2466 3133 2467
rect 3215 2467 3216 2468
rect 3220 2467 3221 2471
rect 3215 2466 3221 2467
rect 3383 2471 3389 2472
rect 3383 2467 3384 2471
rect 3388 2470 3389 2471
rect 3418 2471 3424 2472
rect 3418 2470 3419 2471
rect 3388 2468 3419 2470
rect 3388 2467 3389 2468
rect 3383 2466 3389 2467
rect 3418 2467 3419 2468
rect 3423 2467 3424 2471
rect 3418 2466 3424 2467
rect 3535 2471 3541 2472
rect 3535 2467 3536 2471
rect 3540 2470 3541 2471
rect 3562 2471 3568 2472
rect 3562 2470 3563 2471
rect 3540 2468 3563 2470
rect 3540 2467 3541 2468
rect 3535 2466 3541 2467
rect 3562 2467 3563 2468
rect 3567 2467 3568 2471
rect 3562 2466 3568 2467
rect 214 2463 220 2464
rect 214 2462 215 2463
rect 197 2460 215 2462
rect 214 2459 215 2460
rect 219 2459 220 2463
rect 214 2458 220 2459
rect 274 2463 280 2464
rect 274 2459 275 2463
rect 279 2459 280 2463
rect 274 2458 280 2459
rect 354 2463 360 2464
rect 354 2459 355 2463
rect 359 2459 360 2463
rect 354 2458 360 2459
rect 442 2463 448 2464
rect 442 2459 443 2463
rect 447 2459 448 2463
rect 442 2458 448 2459
rect 562 2463 568 2464
rect 562 2459 563 2463
rect 567 2459 568 2463
rect 562 2458 568 2459
rect 698 2463 704 2464
rect 698 2459 699 2463
rect 703 2459 704 2463
rect 698 2458 704 2459
rect 834 2463 840 2464
rect 834 2459 835 2463
rect 839 2459 840 2463
rect 834 2458 840 2459
rect 934 2463 940 2464
rect 934 2459 935 2463
rect 939 2459 940 2463
rect 1142 2463 1148 2464
rect 1142 2462 1143 2463
rect 1117 2460 1143 2462
rect 934 2458 940 2459
rect 1142 2459 1143 2460
rect 1147 2459 1148 2463
rect 1142 2458 1148 2459
rect 1242 2463 1248 2464
rect 1242 2459 1243 2463
rect 1247 2459 1248 2463
rect 1422 2463 1428 2464
rect 1422 2462 1423 2463
rect 1365 2460 1423 2462
rect 1242 2458 1248 2459
rect 1422 2459 1423 2460
rect 1427 2459 1428 2463
rect 1422 2458 1428 2459
rect 1482 2463 1488 2464
rect 1482 2459 1483 2463
rect 1487 2459 1488 2463
rect 1482 2458 1488 2459
rect 1602 2463 1608 2464
rect 1602 2459 1603 2463
rect 1607 2459 1608 2463
rect 1602 2458 1608 2459
rect 1702 2463 1708 2464
rect 1702 2459 1703 2463
rect 1707 2459 1708 2463
rect 1702 2458 1708 2459
rect 1998 2462 2004 2463
rect 1998 2458 1999 2462
rect 2003 2458 2004 2462
rect 1998 2457 2004 2458
rect 2126 2462 2132 2463
rect 2126 2458 2127 2462
rect 2131 2458 2132 2462
rect 2126 2457 2132 2458
rect 2262 2462 2268 2463
rect 2262 2458 2263 2462
rect 2267 2458 2268 2462
rect 2262 2457 2268 2458
rect 2406 2462 2412 2463
rect 2406 2458 2407 2462
rect 2411 2458 2412 2462
rect 2406 2457 2412 2458
rect 2550 2462 2556 2463
rect 2550 2458 2551 2462
rect 2555 2458 2556 2462
rect 2550 2457 2556 2458
rect 2702 2462 2708 2463
rect 2702 2458 2703 2462
rect 2707 2458 2708 2462
rect 2702 2457 2708 2458
rect 2862 2462 2868 2463
rect 2862 2458 2863 2462
rect 2867 2458 2868 2462
rect 2862 2457 2868 2458
rect 3022 2462 3028 2463
rect 3022 2458 3023 2462
rect 3027 2458 3028 2462
rect 3022 2457 3028 2458
rect 3190 2462 3196 2463
rect 3190 2458 3191 2462
rect 3195 2458 3196 2462
rect 3190 2457 3196 2458
rect 3358 2462 3364 2463
rect 3358 2458 3359 2462
rect 3363 2458 3364 2462
rect 3358 2457 3364 2458
rect 3510 2462 3516 2463
rect 3510 2458 3511 2462
rect 3515 2458 3516 2462
rect 3510 2457 3516 2458
rect 110 2455 116 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 1830 2455 1836 2456
rect 110 2450 116 2451
rect 134 2452 140 2453
rect 134 2448 135 2452
rect 139 2448 140 2452
rect 134 2447 140 2448
rect 214 2452 220 2453
rect 214 2448 215 2452
rect 219 2448 220 2452
rect 214 2447 220 2448
rect 294 2452 300 2453
rect 294 2448 295 2452
rect 299 2448 300 2452
rect 294 2447 300 2448
rect 382 2452 388 2453
rect 382 2448 383 2452
rect 387 2448 388 2452
rect 382 2447 388 2448
rect 502 2452 508 2453
rect 502 2448 503 2452
rect 507 2448 508 2452
rect 502 2447 508 2448
rect 638 2452 644 2453
rect 638 2448 639 2452
rect 643 2448 644 2452
rect 638 2447 644 2448
rect 774 2452 780 2453
rect 774 2448 775 2452
rect 779 2448 780 2452
rect 774 2447 780 2448
rect 918 2452 924 2453
rect 918 2448 919 2452
rect 923 2448 924 2452
rect 918 2447 924 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1302 2452 1308 2453
rect 1302 2448 1303 2452
rect 1307 2448 1308 2452
rect 1302 2447 1308 2448
rect 1422 2452 1428 2453
rect 1422 2448 1423 2452
rect 1427 2448 1428 2452
rect 1422 2447 1428 2448
rect 1542 2452 1548 2453
rect 1542 2448 1543 2452
rect 1547 2448 1548 2452
rect 1542 2447 1548 2448
rect 1662 2452 1668 2453
rect 1662 2448 1663 2452
rect 1667 2448 1668 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1830 2450 1836 2451
rect 1662 2447 1668 2448
rect 1870 2444 1876 2445
rect 1870 2440 1871 2444
rect 1875 2440 1876 2444
rect 1870 2439 1876 2440
rect 3590 2444 3596 2445
rect 3590 2440 3591 2444
rect 3595 2440 3596 2444
rect 3590 2439 3596 2440
rect 2050 2435 2056 2436
rect 2050 2431 2051 2435
rect 2055 2431 2056 2435
rect 2050 2430 2056 2431
rect 2178 2435 2184 2436
rect 2178 2431 2179 2435
rect 2183 2431 2184 2435
rect 2178 2430 2184 2431
rect 2314 2435 2320 2436
rect 2314 2431 2315 2435
rect 2319 2431 2320 2435
rect 2314 2430 2320 2431
rect 2458 2435 2464 2436
rect 2458 2431 2459 2435
rect 2463 2431 2464 2435
rect 2810 2435 2816 2436
rect 2810 2434 2811 2435
rect 2757 2432 2811 2434
rect 2458 2430 2464 2431
rect 2810 2431 2811 2432
rect 2815 2431 2816 2435
rect 2810 2430 2816 2431
rect 2914 2435 2920 2436
rect 2914 2431 2915 2435
rect 2919 2431 2920 2435
rect 3127 2435 3133 2436
rect 3127 2434 3128 2435
rect 3077 2432 3128 2434
rect 2914 2430 2920 2431
rect 3127 2431 3128 2432
rect 3132 2431 3133 2435
rect 3127 2430 3133 2431
rect 3198 2435 3204 2436
rect 3198 2431 3199 2435
rect 3203 2431 3204 2435
rect 3198 2430 3204 2431
rect 3410 2435 3416 2436
rect 3410 2431 3411 2435
rect 3415 2431 3416 2435
rect 3410 2430 3416 2431
rect 3534 2435 3540 2436
rect 3534 2431 3535 2435
rect 3539 2431 3540 2435
rect 3534 2430 3540 2431
rect 1870 2427 1876 2428
rect 1870 2423 1871 2427
rect 1875 2423 1876 2427
rect 3590 2427 3596 2428
rect 1870 2422 1876 2423
rect 1990 2424 1996 2425
rect 1990 2420 1991 2424
rect 1995 2420 1996 2424
rect 1990 2419 1996 2420
rect 2118 2424 2124 2425
rect 2118 2420 2119 2424
rect 2123 2420 2124 2424
rect 2118 2419 2124 2420
rect 2254 2424 2260 2425
rect 2254 2420 2255 2424
rect 2259 2420 2260 2424
rect 2254 2419 2260 2420
rect 2398 2424 2404 2425
rect 2398 2420 2399 2424
rect 2403 2420 2404 2424
rect 2398 2419 2404 2420
rect 2542 2424 2548 2425
rect 2542 2420 2543 2424
rect 2547 2420 2548 2424
rect 2542 2419 2548 2420
rect 2694 2424 2700 2425
rect 2694 2420 2695 2424
rect 2699 2420 2700 2424
rect 2694 2419 2700 2420
rect 2854 2424 2860 2425
rect 2854 2420 2855 2424
rect 2859 2420 2860 2424
rect 2854 2419 2860 2420
rect 3014 2424 3020 2425
rect 3014 2420 3015 2424
rect 3019 2420 3020 2424
rect 3014 2419 3020 2420
rect 3182 2424 3188 2425
rect 3182 2420 3183 2424
rect 3187 2420 3188 2424
rect 3182 2419 3188 2420
rect 3350 2424 3356 2425
rect 3350 2420 3351 2424
rect 3355 2420 3356 2424
rect 3350 2419 3356 2420
rect 3502 2424 3508 2425
rect 3502 2420 3503 2424
rect 3507 2420 3508 2424
rect 3590 2423 3591 2427
rect 3595 2423 3596 2427
rect 3590 2422 3596 2423
rect 3502 2419 3508 2420
rect 2478 2407 2484 2408
rect 2478 2403 2479 2407
rect 2483 2406 2484 2407
rect 2559 2407 2565 2408
rect 2559 2406 2560 2407
rect 2483 2404 2560 2406
rect 2483 2403 2484 2404
rect 2478 2402 2484 2403
rect 2559 2403 2560 2404
rect 2564 2403 2565 2407
rect 2559 2402 2565 2403
rect 1062 2396 1068 2397
rect 110 2393 116 2394
rect 110 2389 111 2393
rect 115 2389 116 2393
rect 1062 2392 1063 2396
rect 1067 2392 1068 2396
rect 1062 2391 1068 2392
rect 1142 2396 1148 2397
rect 1142 2392 1143 2396
rect 1147 2392 1148 2396
rect 1142 2391 1148 2392
rect 1222 2396 1228 2397
rect 1222 2392 1223 2396
rect 1227 2392 1228 2396
rect 1222 2391 1228 2392
rect 1302 2396 1308 2397
rect 1302 2392 1303 2396
rect 1307 2392 1308 2396
rect 1302 2391 1308 2392
rect 1382 2396 1388 2397
rect 1382 2392 1383 2396
rect 1387 2392 1388 2396
rect 1382 2391 1388 2392
rect 1462 2396 1468 2397
rect 1462 2392 1463 2396
rect 1467 2392 1468 2396
rect 1462 2391 1468 2392
rect 1830 2393 1836 2394
rect 110 2388 116 2389
rect 1830 2389 1831 2393
rect 1835 2389 1836 2393
rect 1830 2388 1836 2389
rect 1134 2387 1140 2388
rect 1134 2386 1135 2387
rect 1125 2384 1135 2386
rect 1134 2383 1135 2384
rect 1139 2383 1140 2387
rect 1210 2387 1216 2388
rect 1210 2386 1211 2387
rect 1205 2384 1211 2386
rect 1134 2382 1140 2383
rect 1210 2383 1211 2384
rect 1215 2383 1216 2387
rect 1290 2387 1296 2388
rect 1290 2386 1291 2387
rect 1285 2384 1291 2386
rect 1210 2382 1216 2383
rect 1290 2383 1291 2384
rect 1295 2383 1296 2387
rect 1370 2387 1376 2388
rect 1370 2386 1371 2387
rect 1365 2384 1371 2386
rect 1290 2382 1296 2383
rect 1370 2383 1371 2384
rect 1375 2383 1376 2387
rect 1450 2387 1456 2388
rect 1450 2386 1451 2387
rect 1445 2384 1451 2386
rect 1370 2382 1376 2383
rect 1450 2383 1451 2384
rect 1455 2383 1456 2387
rect 1450 2382 1456 2383
rect 1470 2383 1476 2384
rect 1470 2379 1471 2383
rect 1475 2382 1476 2383
rect 1480 2382 1482 2385
rect 1475 2380 1482 2382
rect 1475 2379 1476 2380
rect 1470 2378 1476 2379
rect 110 2376 116 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 1830 2376 1836 2377
rect 1830 2372 1831 2376
rect 1835 2372 1836 2376
rect 2142 2376 2148 2377
rect 1830 2371 1836 2372
rect 1870 2373 1876 2374
rect 1870 2369 1871 2373
rect 1875 2369 1876 2373
rect 2142 2372 2143 2376
rect 2147 2372 2148 2376
rect 2142 2371 2148 2372
rect 2238 2376 2244 2377
rect 2238 2372 2239 2376
rect 2243 2372 2244 2376
rect 2238 2371 2244 2372
rect 2342 2376 2348 2377
rect 2342 2372 2343 2376
rect 2347 2372 2348 2376
rect 2342 2371 2348 2372
rect 2454 2376 2460 2377
rect 2454 2372 2455 2376
rect 2459 2372 2460 2376
rect 2454 2371 2460 2372
rect 2574 2376 2580 2377
rect 2574 2372 2575 2376
rect 2579 2372 2580 2376
rect 2574 2371 2580 2372
rect 2702 2376 2708 2377
rect 2702 2372 2703 2376
rect 2707 2372 2708 2376
rect 2702 2371 2708 2372
rect 2846 2376 2852 2377
rect 2846 2372 2847 2376
rect 2851 2372 2852 2376
rect 2846 2371 2852 2372
rect 3006 2376 3012 2377
rect 3006 2372 3007 2376
rect 3011 2372 3012 2376
rect 3006 2371 3012 2372
rect 3174 2376 3180 2377
rect 3174 2372 3175 2376
rect 3179 2372 3180 2376
rect 3174 2371 3180 2372
rect 3350 2376 3356 2377
rect 3350 2372 3351 2376
rect 3355 2372 3356 2376
rect 3350 2371 3356 2372
rect 3502 2376 3508 2377
rect 3502 2372 3503 2376
rect 3507 2372 3508 2376
rect 3502 2371 3508 2372
rect 3590 2373 3596 2374
rect 1870 2368 1876 2369
rect 3590 2369 3591 2373
rect 3595 2369 3596 2373
rect 3590 2368 3596 2369
rect 2214 2367 2220 2368
rect 2214 2366 2215 2367
rect 2205 2364 2215 2366
rect 2214 2363 2215 2364
rect 2219 2363 2220 2367
rect 2311 2367 2317 2368
rect 2311 2366 2312 2367
rect 2301 2364 2312 2366
rect 2214 2362 2220 2363
rect 2311 2363 2312 2364
rect 2316 2363 2317 2367
rect 2423 2367 2429 2368
rect 2423 2366 2424 2367
rect 2405 2364 2424 2366
rect 2311 2362 2317 2363
rect 2423 2363 2424 2364
rect 2428 2363 2429 2367
rect 2538 2367 2544 2368
rect 2538 2366 2539 2367
rect 2517 2364 2539 2366
rect 2423 2362 2429 2363
rect 2538 2363 2539 2364
rect 2543 2363 2544 2367
rect 2770 2367 2776 2368
rect 2538 2362 2544 2363
rect 2306 2359 2312 2360
rect 1070 2358 1076 2359
rect 1070 2354 1071 2358
rect 1075 2354 1076 2358
rect 1070 2353 1076 2354
rect 1150 2358 1156 2359
rect 1150 2354 1151 2358
rect 1155 2354 1156 2358
rect 1150 2353 1156 2354
rect 1230 2358 1236 2359
rect 1230 2354 1231 2358
rect 1235 2354 1236 2358
rect 1230 2353 1236 2354
rect 1310 2358 1316 2359
rect 1310 2354 1311 2358
rect 1315 2354 1316 2358
rect 1310 2353 1316 2354
rect 1390 2358 1396 2359
rect 1390 2354 1391 2358
rect 1395 2354 1396 2358
rect 1390 2353 1396 2354
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1870 2356 1876 2357
rect 1870 2352 1871 2356
rect 1875 2352 1876 2356
rect 2306 2355 2307 2359
rect 2311 2358 2312 2359
rect 2592 2358 2594 2365
rect 2311 2356 2594 2358
rect 2764 2358 2766 2365
rect 2770 2363 2771 2367
rect 2775 2366 2776 2367
rect 3114 2367 3120 2368
rect 3114 2366 3115 2367
rect 2775 2364 2865 2366
rect 3069 2364 3115 2366
rect 2775 2363 2776 2364
rect 2770 2362 2776 2363
rect 3114 2363 3115 2364
rect 3119 2363 3120 2367
rect 3114 2362 3120 2363
rect 3122 2367 3128 2368
rect 3122 2363 3123 2367
rect 3127 2366 3128 2367
rect 3418 2367 3424 2368
rect 3418 2366 3419 2367
rect 3127 2364 3193 2366
rect 3413 2364 3419 2366
rect 3127 2363 3128 2364
rect 3122 2362 3128 2363
rect 3418 2363 3419 2364
rect 3423 2363 3424 2367
rect 3570 2367 3576 2368
rect 3570 2366 3571 2367
rect 3565 2364 3571 2366
rect 3418 2362 3424 2363
rect 3570 2363 3571 2364
rect 3575 2363 3576 2367
rect 3570 2362 3576 2363
rect 2775 2359 2781 2360
rect 2775 2358 2776 2359
rect 2764 2356 2776 2358
rect 2311 2355 2312 2356
rect 2306 2354 2312 2355
rect 2775 2355 2776 2356
rect 2780 2355 2781 2359
rect 2775 2354 2781 2355
rect 3590 2356 3596 2357
rect 1870 2351 1876 2352
rect 3590 2352 3591 2356
rect 3595 2352 3596 2356
rect 3590 2351 3596 2352
rect 1095 2347 1101 2348
rect 1095 2343 1096 2347
rect 1100 2346 1101 2347
rect 1134 2347 1140 2348
rect 1100 2344 1130 2346
rect 1100 2343 1101 2344
rect 1095 2342 1101 2343
rect 1128 2338 1130 2344
rect 1134 2343 1135 2347
rect 1139 2346 1140 2347
rect 1175 2347 1181 2348
rect 1175 2346 1176 2347
rect 1139 2344 1176 2346
rect 1139 2343 1140 2344
rect 1134 2342 1140 2343
rect 1175 2343 1176 2344
rect 1180 2343 1181 2347
rect 1175 2342 1181 2343
rect 1210 2347 1216 2348
rect 1210 2343 1211 2347
rect 1215 2346 1216 2347
rect 1255 2347 1261 2348
rect 1255 2346 1256 2347
rect 1215 2344 1256 2346
rect 1215 2343 1216 2344
rect 1210 2342 1216 2343
rect 1255 2343 1256 2344
rect 1260 2343 1261 2347
rect 1255 2342 1261 2343
rect 1290 2347 1296 2348
rect 1290 2343 1291 2347
rect 1295 2346 1296 2347
rect 1335 2347 1341 2348
rect 1335 2346 1336 2347
rect 1295 2344 1336 2346
rect 1295 2343 1296 2344
rect 1290 2342 1296 2343
rect 1335 2343 1336 2344
rect 1340 2343 1341 2347
rect 1335 2342 1341 2343
rect 1370 2347 1376 2348
rect 1370 2343 1371 2347
rect 1375 2346 1376 2347
rect 1415 2347 1421 2348
rect 1415 2346 1416 2347
rect 1375 2344 1416 2346
rect 1375 2343 1376 2344
rect 1370 2342 1376 2343
rect 1415 2343 1416 2344
rect 1420 2343 1421 2347
rect 1415 2342 1421 2343
rect 1450 2347 1456 2348
rect 1450 2343 1451 2347
rect 1455 2346 1456 2347
rect 1495 2347 1501 2348
rect 1495 2346 1496 2347
rect 1455 2344 1496 2346
rect 1455 2343 1456 2344
rect 1450 2342 1456 2343
rect 1495 2343 1496 2344
rect 1500 2343 1501 2347
rect 1495 2342 1501 2343
rect 1326 2339 1332 2340
rect 1326 2338 1327 2339
rect 1128 2336 1327 2338
rect 926 2335 932 2336
rect 926 2334 927 2335
rect 856 2332 927 2334
rect 383 2327 389 2328
rect 383 2323 384 2327
rect 388 2326 389 2327
rect 446 2327 452 2328
rect 446 2326 447 2327
rect 388 2324 447 2326
rect 388 2323 389 2324
rect 383 2322 389 2323
rect 446 2323 447 2324
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 463 2327 469 2328
rect 463 2323 464 2327
rect 468 2326 469 2327
rect 526 2327 532 2328
rect 526 2326 527 2327
rect 468 2324 527 2326
rect 468 2323 469 2324
rect 463 2322 469 2323
rect 526 2323 527 2324
rect 531 2323 532 2327
rect 526 2322 532 2323
rect 543 2327 549 2328
rect 543 2323 544 2327
rect 548 2326 549 2327
rect 606 2327 612 2328
rect 606 2326 607 2327
rect 548 2324 607 2326
rect 548 2323 549 2324
rect 543 2322 549 2323
rect 606 2323 607 2324
rect 611 2323 612 2327
rect 606 2322 612 2323
rect 623 2327 629 2328
rect 623 2323 624 2327
rect 628 2326 629 2327
rect 686 2327 692 2328
rect 686 2326 687 2327
rect 628 2324 687 2326
rect 628 2323 629 2324
rect 623 2322 629 2323
rect 686 2323 687 2324
rect 691 2323 692 2327
rect 686 2322 692 2323
rect 703 2327 709 2328
rect 703 2323 704 2327
rect 708 2326 709 2327
rect 766 2327 772 2328
rect 766 2326 767 2327
rect 708 2324 767 2326
rect 708 2323 709 2324
rect 703 2322 709 2323
rect 766 2323 767 2324
rect 771 2323 772 2327
rect 766 2322 772 2323
rect 783 2327 789 2328
rect 783 2323 784 2327
rect 788 2326 789 2327
rect 856 2326 858 2332
rect 926 2331 927 2332
rect 931 2331 932 2335
rect 1326 2335 1327 2336
rect 1331 2335 1332 2339
rect 1326 2334 1332 2335
rect 2150 2338 2156 2339
rect 2150 2334 2151 2338
rect 2155 2334 2156 2338
rect 2150 2333 2156 2334
rect 2246 2338 2252 2339
rect 2246 2334 2247 2338
rect 2251 2334 2252 2338
rect 2246 2333 2252 2334
rect 2350 2338 2356 2339
rect 2350 2334 2351 2338
rect 2355 2334 2356 2338
rect 2350 2333 2356 2334
rect 2462 2338 2468 2339
rect 2462 2334 2463 2338
rect 2467 2334 2468 2338
rect 2462 2333 2468 2334
rect 2582 2338 2588 2339
rect 2582 2334 2583 2338
rect 2587 2334 2588 2338
rect 2582 2333 2588 2334
rect 2710 2338 2716 2339
rect 2710 2334 2711 2338
rect 2715 2334 2716 2338
rect 2710 2333 2716 2334
rect 2854 2338 2860 2339
rect 2854 2334 2855 2338
rect 2859 2334 2860 2338
rect 2854 2333 2860 2334
rect 3014 2338 3020 2339
rect 3014 2334 3015 2338
rect 3019 2334 3020 2338
rect 3014 2333 3020 2334
rect 3182 2338 3188 2339
rect 3182 2334 3183 2338
rect 3187 2334 3188 2338
rect 3182 2333 3188 2334
rect 3358 2338 3364 2339
rect 3358 2334 3359 2338
rect 3363 2334 3364 2338
rect 3358 2333 3364 2334
rect 3510 2338 3516 2339
rect 3510 2334 3511 2338
rect 3515 2334 3516 2338
rect 3510 2333 3516 2334
rect 926 2330 932 2331
rect 788 2324 858 2326
rect 862 2327 869 2328
rect 788 2323 789 2324
rect 783 2322 789 2323
rect 862 2323 863 2327
rect 868 2323 869 2327
rect 862 2322 869 2323
rect 890 2327 896 2328
rect 890 2323 891 2327
rect 895 2326 896 2327
rect 943 2327 949 2328
rect 943 2326 944 2327
rect 895 2324 944 2326
rect 895 2323 896 2324
rect 890 2322 896 2323
rect 943 2323 944 2324
rect 948 2323 949 2327
rect 943 2322 949 2323
rect 1023 2327 1029 2328
rect 1023 2323 1024 2327
rect 1028 2326 1029 2327
rect 1042 2327 1048 2328
rect 1042 2326 1043 2327
rect 1028 2324 1043 2326
rect 1028 2323 1029 2324
rect 1023 2322 1029 2323
rect 1042 2323 1043 2324
rect 1047 2323 1048 2327
rect 1042 2322 1048 2323
rect 1050 2327 1056 2328
rect 1050 2323 1051 2327
rect 1055 2326 1056 2327
rect 1103 2327 1109 2328
rect 1103 2326 1104 2327
rect 1055 2324 1104 2326
rect 1055 2323 1056 2324
rect 1050 2322 1056 2323
rect 1103 2323 1104 2324
rect 1108 2323 1109 2327
rect 1103 2322 1109 2323
rect 1130 2327 1136 2328
rect 1130 2323 1131 2327
rect 1135 2326 1136 2327
rect 1183 2327 1189 2328
rect 1183 2326 1184 2327
rect 1135 2324 1184 2326
rect 1135 2323 1136 2324
rect 1130 2322 1136 2323
rect 1183 2323 1184 2324
rect 1188 2323 1189 2327
rect 1183 2322 1189 2323
rect 1210 2327 1216 2328
rect 1210 2323 1211 2327
rect 1215 2326 1216 2327
rect 1263 2327 1269 2328
rect 1263 2326 1264 2327
rect 1215 2324 1264 2326
rect 1215 2323 1216 2324
rect 1210 2322 1216 2323
rect 1263 2323 1264 2324
rect 1268 2323 1269 2327
rect 1263 2322 1269 2323
rect 1290 2327 1296 2328
rect 1290 2323 1291 2327
rect 1295 2326 1296 2327
rect 1343 2327 1349 2328
rect 1343 2326 1344 2327
rect 1295 2324 1344 2326
rect 1295 2323 1296 2324
rect 1290 2322 1296 2323
rect 1343 2323 1344 2324
rect 1348 2323 1349 2327
rect 1343 2322 1349 2323
rect 2175 2327 2184 2328
rect 2175 2323 2176 2327
rect 2183 2323 2184 2327
rect 2175 2322 2184 2323
rect 2214 2327 2220 2328
rect 2214 2323 2215 2327
rect 2219 2326 2220 2327
rect 2271 2327 2277 2328
rect 2271 2326 2272 2327
rect 2219 2324 2272 2326
rect 2219 2323 2220 2324
rect 2214 2322 2220 2323
rect 2271 2323 2272 2324
rect 2276 2323 2277 2327
rect 2271 2322 2277 2323
rect 2311 2327 2317 2328
rect 2311 2323 2312 2327
rect 2316 2326 2317 2327
rect 2375 2327 2381 2328
rect 2375 2326 2376 2327
rect 2316 2324 2376 2326
rect 2316 2323 2317 2324
rect 2311 2322 2317 2323
rect 2375 2323 2376 2324
rect 2380 2323 2381 2327
rect 2375 2322 2381 2323
rect 2423 2327 2429 2328
rect 2423 2323 2424 2327
rect 2428 2326 2429 2327
rect 2487 2327 2493 2328
rect 2487 2326 2488 2327
rect 2428 2324 2488 2326
rect 2428 2323 2429 2324
rect 2423 2322 2429 2323
rect 2487 2323 2488 2324
rect 2492 2323 2493 2327
rect 2487 2322 2493 2323
rect 2538 2327 2544 2328
rect 2538 2323 2539 2327
rect 2543 2326 2544 2327
rect 2607 2327 2613 2328
rect 2607 2326 2608 2327
rect 2543 2324 2608 2326
rect 2543 2323 2544 2324
rect 2538 2322 2544 2323
rect 2607 2323 2608 2324
rect 2612 2323 2613 2327
rect 2607 2322 2613 2323
rect 2735 2327 2741 2328
rect 2735 2323 2736 2327
rect 2740 2326 2741 2327
rect 2770 2327 2776 2328
rect 2770 2326 2771 2327
rect 2740 2324 2771 2326
rect 2740 2323 2741 2324
rect 2735 2322 2741 2323
rect 2770 2323 2771 2324
rect 2775 2323 2776 2327
rect 2770 2322 2776 2323
rect 2879 2327 2888 2328
rect 2879 2323 2880 2327
rect 2887 2323 2888 2327
rect 2879 2322 2888 2323
rect 2914 2327 2920 2328
rect 2914 2323 2915 2327
rect 2919 2326 2920 2327
rect 3039 2327 3045 2328
rect 3039 2326 3040 2327
rect 2919 2324 3040 2326
rect 2919 2323 2920 2324
rect 2914 2322 2920 2323
rect 3039 2323 3040 2324
rect 3044 2323 3045 2327
rect 3039 2322 3045 2323
rect 3114 2327 3120 2328
rect 3114 2323 3115 2327
rect 3119 2326 3120 2327
rect 3207 2327 3213 2328
rect 3207 2326 3208 2327
rect 3119 2324 3208 2326
rect 3119 2323 3120 2324
rect 3114 2322 3120 2323
rect 3207 2323 3208 2324
rect 3212 2323 3213 2327
rect 3207 2322 3213 2323
rect 3383 2327 3389 2328
rect 3383 2323 3384 2327
rect 3388 2326 3389 2327
rect 3418 2327 3424 2328
rect 3418 2326 3419 2327
rect 3388 2324 3419 2326
rect 3388 2323 3389 2324
rect 3383 2322 3389 2323
rect 3418 2323 3419 2324
rect 3423 2323 3424 2327
rect 3418 2322 3424 2323
rect 3534 2327 3541 2328
rect 3534 2323 3535 2327
rect 3540 2323 3541 2327
rect 3534 2322 3541 2323
rect 2942 2319 2948 2320
rect 358 2318 364 2319
rect 358 2314 359 2318
rect 363 2314 364 2318
rect 358 2313 364 2314
rect 438 2318 444 2319
rect 438 2314 439 2318
rect 443 2314 444 2318
rect 438 2313 444 2314
rect 518 2318 524 2319
rect 518 2314 519 2318
rect 523 2314 524 2318
rect 518 2313 524 2314
rect 598 2318 604 2319
rect 598 2314 599 2318
rect 603 2314 604 2318
rect 598 2313 604 2314
rect 678 2318 684 2319
rect 678 2314 679 2318
rect 683 2314 684 2318
rect 678 2313 684 2314
rect 758 2318 764 2319
rect 758 2314 759 2318
rect 763 2314 764 2318
rect 758 2313 764 2314
rect 838 2318 844 2319
rect 838 2314 839 2318
rect 843 2314 844 2318
rect 838 2313 844 2314
rect 918 2318 924 2319
rect 918 2314 919 2318
rect 923 2314 924 2318
rect 918 2313 924 2314
rect 998 2318 1004 2319
rect 998 2314 999 2318
rect 1003 2314 1004 2318
rect 998 2313 1004 2314
rect 1078 2318 1084 2319
rect 1078 2314 1079 2318
rect 1083 2314 1084 2318
rect 1078 2313 1084 2314
rect 1158 2318 1164 2319
rect 1158 2314 1159 2318
rect 1163 2314 1164 2318
rect 1158 2313 1164 2314
rect 1238 2318 1244 2319
rect 1238 2314 1239 2318
rect 1243 2314 1244 2318
rect 1238 2313 1244 2314
rect 1318 2318 1324 2319
rect 2942 2318 2943 2319
rect 1318 2314 1319 2318
rect 1323 2314 1324 2318
rect 1318 2313 1324 2314
rect 2768 2316 2943 2318
rect 2303 2311 2312 2312
rect 2303 2307 2304 2311
rect 2311 2307 2312 2311
rect 2303 2306 2312 2307
rect 2330 2311 2336 2312
rect 2330 2307 2331 2311
rect 2335 2310 2336 2311
rect 2383 2311 2389 2312
rect 2383 2310 2384 2311
rect 2335 2308 2384 2310
rect 2335 2307 2336 2308
rect 2330 2306 2336 2307
rect 2383 2307 2384 2308
rect 2388 2307 2389 2311
rect 2383 2306 2389 2307
rect 2410 2311 2416 2312
rect 2410 2307 2411 2311
rect 2415 2310 2416 2311
rect 2463 2311 2469 2312
rect 2463 2310 2464 2311
rect 2415 2308 2464 2310
rect 2415 2307 2416 2308
rect 2410 2306 2416 2307
rect 2463 2307 2464 2308
rect 2468 2307 2469 2311
rect 2463 2306 2469 2307
rect 2490 2311 2496 2312
rect 2490 2307 2491 2311
rect 2495 2310 2496 2311
rect 2543 2311 2549 2312
rect 2543 2310 2544 2311
rect 2495 2308 2544 2310
rect 2495 2307 2496 2308
rect 2490 2306 2496 2307
rect 2543 2307 2544 2308
rect 2548 2307 2549 2311
rect 2543 2306 2549 2307
rect 2623 2311 2629 2312
rect 2623 2307 2624 2311
rect 2628 2310 2629 2311
rect 2686 2311 2692 2312
rect 2686 2310 2687 2311
rect 2628 2308 2687 2310
rect 2628 2307 2629 2308
rect 2623 2306 2629 2307
rect 2686 2307 2687 2308
rect 2691 2307 2692 2311
rect 2686 2306 2692 2307
rect 2703 2311 2709 2312
rect 2703 2307 2704 2311
rect 2708 2310 2709 2311
rect 2768 2310 2770 2316
rect 2942 2315 2943 2316
rect 2947 2315 2948 2319
rect 2942 2314 2948 2315
rect 2708 2308 2770 2310
rect 2775 2311 2781 2312
rect 2708 2307 2709 2308
rect 2703 2306 2709 2307
rect 2775 2307 2776 2311
rect 2780 2310 2781 2311
rect 2783 2311 2789 2312
rect 2783 2310 2784 2311
rect 2780 2308 2784 2310
rect 2780 2307 2781 2308
rect 2775 2306 2781 2307
rect 2783 2307 2784 2308
rect 2788 2307 2789 2311
rect 2783 2306 2789 2307
rect 2810 2311 2816 2312
rect 2810 2307 2811 2311
rect 2815 2310 2816 2311
rect 2871 2311 2877 2312
rect 2871 2310 2872 2311
rect 2815 2308 2872 2310
rect 2815 2307 2816 2308
rect 2810 2306 2816 2307
rect 2871 2307 2872 2308
rect 2876 2307 2877 2311
rect 2871 2306 2877 2307
rect 2898 2311 2904 2312
rect 2898 2307 2899 2311
rect 2903 2310 2904 2311
rect 2959 2311 2965 2312
rect 2959 2310 2960 2311
rect 2903 2308 2960 2310
rect 2903 2307 2904 2308
rect 2898 2306 2904 2307
rect 2959 2307 2960 2308
rect 2964 2307 2965 2311
rect 2959 2306 2965 2307
rect 2278 2302 2284 2303
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 110 2295 116 2296
rect 1830 2300 1836 2301
rect 1830 2296 1831 2300
rect 1835 2296 1836 2300
rect 2278 2298 2279 2302
rect 2283 2298 2284 2302
rect 2278 2297 2284 2298
rect 2358 2302 2364 2303
rect 2358 2298 2359 2302
rect 2363 2298 2364 2302
rect 2358 2297 2364 2298
rect 2438 2302 2444 2303
rect 2438 2298 2439 2302
rect 2443 2298 2444 2302
rect 2438 2297 2444 2298
rect 2518 2302 2524 2303
rect 2518 2298 2519 2302
rect 2523 2298 2524 2302
rect 2518 2297 2524 2298
rect 2598 2302 2604 2303
rect 2598 2298 2599 2302
rect 2603 2298 2604 2302
rect 2598 2297 2604 2298
rect 2678 2302 2684 2303
rect 2678 2298 2679 2302
rect 2683 2298 2684 2302
rect 2678 2297 2684 2298
rect 2758 2302 2764 2303
rect 2758 2298 2759 2302
rect 2763 2298 2764 2302
rect 2758 2297 2764 2298
rect 2846 2302 2852 2303
rect 2846 2298 2847 2302
rect 2851 2298 2852 2302
rect 2846 2297 2852 2298
rect 2934 2302 2940 2303
rect 2934 2298 2935 2302
rect 2939 2298 2940 2302
rect 2934 2297 2940 2298
rect 1830 2295 1836 2296
rect 406 2291 412 2292
rect 406 2287 407 2291
rect 411 2287 412 2291
rect 406 2286 412 2287
rect 446 2291 452 2292
rect 446 2287 447 2291
rect 451 2287 452 2291
rect 446 2286 452 2287
rect 526 2291 532 2292
rect 526 2287 527 2291
rect 531 2287 532 2291
rect 526 2286 532 2287
rect 606 2291 612 2292
rect 606 2287 607 2291
rect 611 2287 612 2291
rect 606 2286 612 2287
rect 686 2291 692 2292
rect 686 2287 687 2291
rect 691 2287 692 2291
rect 686 2286 692 2287
rect 766 2291 772 2292
rect 766 2287 767 2291
rect 771 2287 772 2291
rect 766 2286 772 2287
rect 890 2291 896 2292
rect 890 2287 891 2291
rect 895 2287 896 2291
rect 890 2286 896 2287
rect 926 2291 932 2292
rect 926 2287 927 2291
rect 931 2287 932 2291
rect 926 2286 932 2287
rect 1050 2291 1056 2292
rect 1050 2287 1051 2291
rect 1055 2287 1056 2291
rect 1050 2286 1056 2287
rect 1130 2291 1136 2292
rect 1130 2287 1131 2291
rect 1135 2287 1136 2291
rect 1130 2286 1136 2287
rect 1210 2291 1216 2292
rect 1210 2287 1211 2291
rect 1215 2287 1216 2291
rect 1210 2286 1216 2287
rect 1290 2291 1296 2292
rect 1290 2287 1291 2291
rect 1295 2287 1296 2291
rect 1290 2286 1296 2287
rect 1326 2291 1332 2292
rect 1326 2287 1327 2291
rect 1331 2287 1332 2291
rect 1326 2286 1332 2287
rect 1870 2284 1876 2285
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 1830 2283 1836 2284
rect 110 2278 116 2279
rect 350 2280 356 2281
rect 350 2276 351 2280
rect 355 2276 356 2280
rect 350 2275 356 2276
rect 430 2280 436 2281
rect 430 2276 431 2280
rect 435 2276 436 2280
rect 430 2275 436 2276
rect 510 2280 516 2281
rect 510 2276 511 2280
rect 515 2276 516 2280
rect 510 2275 516 2276
rect 590 2280 596 2281
rect 590 2276 591 2280
rect 595 2276 596 2280
rect 590 2275 596 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 750 2280 756 2281
rect 750 2276 751 2280
rect 755 2276 756 2280
rect 750 2275 756 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 1070 2280 1076 2281
rect 1070 2276 1071 2280
rect 1075 2276 1076 2280
rect 1070 2275 1076 2276
rect 1150 2280 1156 2281
rect 1150 2276 1151 2280
rect 1155 2276 1156 2280
rect 1150 2275 1156 2276
rect 1230 2280 1236 2281
rect 1230 2276 1231 2280
rect 1235 2276 1236 2280
rect 1230 2275 1236 2276
rect 1310 2280 1316 2281
rect 1310 2276 1311 2280
rect 1315 2276 1316 2280
rect 1830 2279 1831 2283
rect 1835 2279 1836 2283
rect 1870 2280 1871 2284
rect 1875 2280 1876 2284
rect 1870 2279 1876 2280
rect 3590 2284 3596 2285
rect 3590 2280 3591 2284
rect 3595 2280 3596 2284
rect 3590 2279 3596 2280
rect 1830 2278 1836 2279
rect 1310 2275 1316 2276
rect 2330 2275 2336 2276
rect 2330 2271 2331 2275
rect 2335 2271 2336 2275
rect 2330 2270 2336 2271
rect 2410 2275 2416 2276
rect 2410 2271 2411 2275
rect 2415 2271 2416 2275
rect 2410 2270 2416 2271
rect 2490 2275 2496 2276
rect 2490 2271 2491 2275
rect 2495 2271 2496 2275
rect 2490 2270 2496 2271
rect 2630 2275 2636 2276
rect 2630 2271 2631 2275
rect 2635 2271 2636 2275
rect 2630 2270 2636 2271
rect 2686 2275 2692 2276
rect 2686 2271 2687 2275
rect 2691 2271 2692 2275
rect 2686 2270 2692 2271
rect 2810 2275 2816 2276
rect 2810 2271 2811 2275
rect 2815 2271 2816 2275
rect 2810 2270 2816 2271
rect 2898 2275 2904 2276
rect 2898 2271 2899 2275
rect 2903 2271 2904 2275
rect 2898 2270 2904 2271
rect 2942 2275 2948 2276
rect 2942 2271 2943 2275
rect 2947 2271 2948 2275
rect 2942 2270 2948 2271
rect 1870 2267 1876 2268
rect 1870 2263 1871 2267
rect 1875 2263 1876 2267
rect 3590 2267 3596 2268
rect 1870 2262 1876 2263
rect 2270 2264 2276 2265
rect 2270 2260 2271 2264
rect 2275 2260 2276 2264
rect 1042 2259 1048 2260
rect 1042 2255 1043 2259
rect 1047 2258 1048 2259
rect 1242 2259 1248 2260
rect 2270 2259 2276 2260
rect 2350 2264 2356 2265
rect 2350 2260 2351 2264
rect 2355 2260 2356 2264
rect 2350 2259 2356 2260
rect 2430 2264 2436 2265
rect 2430 2260 2431 2264
rect 2435 2260 2436 2264
rect 2430 2259 2436 2260
rect 2510 2264 2516 2265
rect 2510 2260 2511 2264
rect 2515 2260 2516 2264
rect 2510 2259 2516 2260
rect 2590 2264 2596 2265
rect 2590 2260 2591 2264
rect 2595 2260 2596 2264
rect 2590 2259 2596 2260
rect 2670 2264 2676 2265
rect 2670 2260 2671 2264
rect 2675 2260 2676 2264
rect 2670 2259 2676 2260
rect 2750 2264 2756 2265
rect 2750 2260 2751 2264
rect 2755 2260 2756 2264
rect 2750 2259 2756 2260
rect 2838 2264 2844 2265
rect 2838 2260 2839 2264
rect 2843 2260 2844 2264
rect 2838 2259 2844 2260
rect 2926 2264 2932 2265
rect 2926 2260 2927 2264
rect 2931 2260 2932 2264
rect 3590 2263 3591 2267
rect 3595 2263 3596 2267
rect 3590 2262 3596 2263
rect 2926 2259 2932 2260
rect 1242 2258 1243 2259
rect 1047 2256 1243 2258
rect 1047 2255 1048 2256
rect 1042 2254 1048 2255
rect 1242 2255 1243 2256
rect 1247 2255 1248 2259
rect 1242 2254 1248 2255
rect 2358 2247 2364 2248
rect 2358 2243 2359 2247
rect 2363 2246 2364 2247
rect 2527 2247 2533 2248
rect 2527 2246 2528 2247
rect 2363 2244 2528 2246
rect 2363 2243 2364 2244
rect 2358 2242 2364 2243
rect 2527 2243 2528 2244
rect 2532 2243 2533 2247
rect 2527 2242 2533 2243
rect 374 2236 380 2237
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 374 2232 375 2236
rect 379 2232 380 2236
rect 374 2231 380 2232
rect 454 2236 460 2237
rect 454 2232 455 2236
rect 459 2232 460 2236
rect 454 2231 460 2232
rect 534 2236 540 2237
rect 534 2232 535 2236
rect 539 2232 540 2236
rect 534 2231 540 2232
rect 614 2236 620 2237
rect 614 2232 615 2236
rect 619 2232 620 2236
rect 614 2231 620 2232
rect 694 2236 700 2237
rect 694 2232 695 2236
rect 699 2232 700 2236
rect 694 2231 700 2232
rect 774 2236 780 2237
rect 774 2232 775 2236
rect 779 2232 780 2236
rect 774 2231 780 2232
rect 854 2236 860 2237
rect 854 2232 855 2236
rect 859 2232 860 2236
rect 854 2231 860 2232
rect 934 2236 940 2237
rect 934 2232 935 2236
rect 939 2232 940 2236
rect 934 2231 940 2232
rect 1014 2236 1020 2237
rect 1014 2232 1015 2236
rect 1019 2232 1020 2236
rect 1014 2231 1020 2232
rect 1094 2236 1100 2237
rect 1094 2232 1095 2236
rect 1099 2232 1100 2236
rect 1094 2231 1100 2232
rect 1174 2236 1180 2237
rect 1174 2232 1175 2236
rect 1179 2232 1180 2236
rect 1174 2231 1180 2232
rect 1254 2236 1260 2237
rect 1254 2232 1255 2236
rect 1259 2232 1260 2236
rect 1254 2231 1260 2232
rect 1830 2233 1836 2234
rect 110 2228 116 2229
rect 1830 2229 1831 2233
rect 1835 2229 1836 2233
rect 1830 2228 1836 2229
rect 442 2227 448 2228
rect 442 2226 443 2227
rect 437 2224 443 2226
rect 442 2223 443 2224
rect 447 2223 448 2227
rect 526 2227 532 2228
rect 442 2222 448 2223
rect 516 2220 518 2225
rect 526 2223 527 2227
rect 531 2226 532 2227
rect 682 2227 688 2228
rect 682 2226 683 2227
rect 531 2224 553 2226
rect 677 2224 683 2226
rect 531 2223 532 2224
rect 526 2222 532 2223
rect 682 2223 683 2224
rect 687 2223 688 2227
rect 762 2227 768 2228
rect 762 2226 763 2227
rect 757 2224 763 2226
rect 682 2222 688 2223
rect 762 2223 763 2224
rect 767 2223 768 2227
rect 922 2227 928 2228
rect 922 2226 923 2227
rect 762 2222 768 2223
rect 836 2222 838 2225
rect 917 2224 923 2226
rect 862 2223 868 2224
rect 862 2222 863 2223
rect 836 2220 863 2222
rect 514 2219 520 2220
rect 110 2216 116 2217
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 514 2215 515 2219
rect 519 2215 520 2219
rect 862 2219 863 2220
rect 867 2219 868 2223
rect 922 2223 923 2224
rect 927 2223 928 2227
rect 1002 2227 1008 2228
rect 1002 2226 1003 2227
rect 997 2224 1003 2226
rect 922 2222 928 2223
rect 1002 2223 1003 2224
rect 1007 2223 1008 2227
rect 1082 2227 1088 2228
rect 1082 2226 1083 2227
rect 1077 2224 1083 2226
rect 1002 2222 1008 2223
rect 1082 2223 1083 2224
rect 1087 2223 1088 2227
rect 1167 2227 1173 2228
rect 1167 2226 1168 2227
rect 1157 2224 1168 2226
rect 1082 2222 1088 2223
rect 1167 2223 1168 2224
rect 1172 2223 1173 2227
rect 1242 2227 1248 2228
rect 1167 2222 1173 2223
rect 1236 2220 1238 2225
rect 1242 2223 1243 2227
rect 1247 2226 1248 2227
rect 1247 2224 1273 2226
rect 1247 2223 1248 2224
rect 1242 2222 1248 2223
rect 2310 2220 2316 2221
rect 862 2218 868 2219
rect 1234 2219 1240 2220
rect 514 2214 520 2215
rect 1234 2215 1235 2219
rect 1239 2215 1240 2219
rect 1870 2217 1876 2218
rect 1234 2214 1240 2215
rect 1830 2216 1836 2217
rect 110 2211 116 2212
rect 1830 2212 1831 2216
rect 1835 2212 1836 2216
rect 1870 2213 1871 2217
rect 1875 2213 1876 2217
rect 2310 2216 2311 2220
rect 2315 2216 2316 2220
rect 2310 2215 2316 2216
rect 2398 2220 2404 2221
rect 2398 2216 2399 2220
rect 2403 2216 2404 2220
rect 2398 2215 2404 2216
rect 2494 2220 2500 2221
rect 2494 2216 2495 2220
rect 2499 2216 2500 2220
rect 2494 2215 2500 2216
rect 2598 2220 2604 2221
rect 2598 2216 2599 2220
rect 2603 2216 2604 2220
rect 2598 2215 2604 2216
rect 2718 2220 2724 2221
rect 2718 2216 2719 2220
rect 2723 2216 2724 2220
rect 2718 2215 2724 2216
rect 2854 2220 2860 2221
rect 2854 2216 2855 2220
rect 2859 2216 2860 2220
rect 2854 2215 2860 2216
rect 3006 2220 3012 2221
rect 3006 2216 3007 2220
rect 3011 2216 3012 2220
rect 3006 2215 3012 2216
rect 3174 2220 3180 2221
rect 3174 2216 3175 2220
rect 3179 2216 3180 2220
rect 3174 2215 3180 2216
rect 3350 2220 3356 2221
rect 3350 2216 3351 2220
rect 3355 2216 3356 2220
rect 3350 2215 3356 2216
rect 3502 2220 3508 2221
rect 3502 2216 3503 2220
rect 3507 2216 3508 2220
rect 3502 2215 3508 2216
rect 3590 2217 3596 2218
rect 1870 2212 1876 2213
rect 3590 2213 3591 2217
rect 3595 2213 3596 2217
rect 3590 2212 3596 2213
rect 1830 2211 1836 2212
rect 2378 2211 2384 2212
rect 2378 2210 2379 2211
rect 2373 2208 2379 2210
rect 2378 2207 2379 2208
rect 2383 2207 2384 2211
rect 2470 2211 2476 2212
rect 2470 2210 2471 2211
rect 2461 2208 2471 2210
rect 2378 2206 2384 2207
rect 2470 2207 2471 2208
rect 2475 2207 2476 2211
rect 2562 2211 2568 2212
rect 2562 2210 2563 2211
rect 2557 2208 2563 2210
rect 2470 2206 2476 2207
rect 2562 2207 2563 2208
rect 2567 2207 2568 2211
rect 2678 2211 2684 2212
rect 2678 2210 2679 2211
rect 2661 2208 2679 2210
rect 2562 2206 2568 2207
rect 2678 2207 2679 2208
rect 2683 2207 2684 2211
rect 2786 2211 2792 2212
rect 2786 2210 2787 2211
rect 2781 2208 2787 2210
rect 2678 2206 2684 2207
rect 2786 2207 2787 2208
rect 2791 2207 2792 2211
rect 2927 2211 2933 2212
rect 2927 2210 2928 2211
rect 2917 2208 2928 2210
rect 2786 2206 2792 2207
rect 2927 2207 2928 2208
rect 2932 2207 2933 2211
rect 3074 2211 3080 2212
rect 3074 2210 3075 2211
rect 3069 2208 3075 2210
rect 2927 2206 2933 2207
rect 3074 2207 3075 2208
rect 3079 2207 3080 2211
rect 3074 2206 3080 2207
rect 3082 2211 3088 2212
rect 3082 2207 3083 2211
rect 3087 2210 3088 2211
rect 3418 2211 3424 2212
rect 3418 2210 3419 2211
rect 3087 2208 3193 2210
rect 3413 2208 3419 2210
rect 3087 2207 3088 2208
rect 3082 2206 3088 2207
rect 3418 2207 3419 2208
rect 3423 2207 3424 2211
rect 3418 2206 3424 2207
rect 3564 2204 3566 2209
rect 3562 2203 3568 2204
rect 1870 2200 1876 2201
rect 382 2198 388 2199
rect 382 2194 383 2198
rect 387 2194 388 2198
rect 382 2193 388 2194
rect 462 2198 468 2199
rect 462 2194 463 2198
rect 467 2194 468 2198
rect 462 2193 468 2194
rect 542 2198 548 2199
rect 542 2194 543 2198
rect 547 2194 548 2198
rect 542 2193 548 2194
rect 622 2198 628 2199
rect 622 2194 623 2198
rect 627 2194 628 2198
rect 622 2193 628 2194
rect 702 2198 708 2199
rect 702 2194 703 2198
rect 707 2194 708 2198
rect 702 2193 708 2194
rect 782 2198 788 2199
rect 782 2194 783 2198
rect 787 2194 788 2198
rect 782 2193 788 2194
rect 862 2198 868 2199
rect 862 2194 863 2198
rect 867 2194 868 2198
rect 862 2193 868 2194
rect 942 2198 948 2199
rect 942 2194 943 2198
rect 947 2194 948 2198
rect 942 2193 948 2194
rect 1022 2198 1028 2199
rect 1022 2194 1023 2198
rect 1027 2194 1028 2198
rect 1022 2193 1028 2194
rect 1102 2198 1108 2199
rect 1102 2194 1103 2198
rect 1107 2194 1108 2198
rect 1102 2193 1108 2194
rect 1182 2198 1188 2199
rect 1182 2194 1183 2198
rect 1187 2194 1188 2198
rect 1182 2193 1188 2194
rect 1262 2198 1268 2199
rect 1262 2194 1263 2198
rect 1267 2194 1268 2198
rect 1870 2196 1871 2200
rect 1875 2196 1876 2200
rect 3562 2199 3563 2203
rect 3567 2199 3568 2203
rect 3562 2198 3568 2199
rect 3590 2200 3596 2201
rect 1870 2195 1876 2196
rect 3590 2196 3591 2200
rect 3595 2196 3596 2200
rect 3590 2195 3596 2196
rect 1262 2193 1268 2194
rect 406 2187 413 2188
rect 406 2183 407 2187
rect 412 2183 413 2187
rect 406 2182 413 2183
rect 442 2187 448 2188
rect 442 2183 443 2187
rect 447 2186 448 2187
rect 487 2187 493 2188
rect 487 2186 488 2187
rect 447 2184 488 2186
rect 447 2183 448 2184
rect 442 2182 448 2183
rect 487 2183 488 2184
rect 492 2183 493 2187
rect 487 2182 493 2183
rect 514 2187 520 2188
rect 514 2183 515 2187
rect 519 2186 520 2187
rect 567 2187 573 2188
rect 567 2186 568 2187
rect 519 2184 568 2186
rect 519 2183 520 2184
rect 514 2182 520 2183
rect 567 2183 568 2184
rect 572 2183 573 2187
rect 567 2182 573 2183
rect 647 2187 653 2188
rect 647 2183 648 2187
rect 652 2186 653 2187
rect 682 2187 688 2188
rect 652 2184 678 2186
rect 652 2183 653 2184
rect 647 2182 653 2183
rect 676 2178 678 2184
rect 682 2183 683 2187
rect 687 2186 688 2187
rect 727 2187 733 2188
rect 727 2186 728 2187
rect 687 2184 728 2186
rect 687 2183 688 2184
rect 682 2182 688 2183
rect 727 2183 728 2184
rect 732 2183 733 2187
rect 727 2182 733 2183
rect 762 2187 768 2188
rect 762 2183 763 2187
rect 767 2186 768 2187
rect 807 2187 813 2188
rect 807 2186 808 2187
rect 767 2184 808 2186
rect 767 2183 768 2184
rect 762 2182 768 2183
rect 807 2183 808 2184
rect 812 2183 813 2187
rect 807 2182 813 2183
rect 886 2187 893 2188
rect 886 2183 887 2187
rect 892 2183 893 2187
rect 886 2182 893 2183
rect 922 2187 928 2188
rect 922 2183 923 2187
rect 927 2186 928 2187
rect 967 2187 973 2188
rect 967 2186 968 2187
rect 927 2184 968 2186
rect 927 2183 928 2184
rect 922 2182 928 2183
rect 967 2183 968 2184
rect 972 2183 973 2187
rect 967 2182 973 2183
rect 1002 2187 1008 2188
rect 1002 2183 1003 2187
rect 1007 2186 1008 2187
rect 1047 2187 1053 2188
rect 1047 2186 1048 2187
rect 1007 2184 1048 2186
rect 1007 2183 1008 2184
rect 1002 2182 1008 2183
rect 1047 2183 1048 2184
rect 1052 2183 1053 2187
rect 1047 2182 1053 2183
rect 1082 2187 1088 2188
rect 1082 2183 1083 2187
rect 1087 2186 1088 2187
rect 1127 2187 1133 2188
rect 1127 2186 1128 2187
rect 1087 2184 1128 2186
rect 1087 2183 1088 2184
rect 1082 2182 1088 2183
rect 1127 2183 1128 2184
rect 1132 2183 1133 2187
rect 1127 2182 1133 2183
rect 1167 2187 1173 2188
rect 1167 2183 1168 2187
rect 1172 2186 1173 2187
rect 1207 2187 1213 2188
rect 1207 2186 1208 2187
rect 1172 2184 1208 2186
rect 1172 2183 1173 2184
rect 1167 2182 1173 2183
rect 1207 2183 1208 2184
rect 1212 2183 1213 2187
rect 1207 2182 1213 2183
rect 1234 2187 1240 2188
rect 1234 2183 1235 2187
rect 1239 2186 1240 2187
rect 1287 2187 1293 2188
rect 1287 2186 1288 2187
rect 1239 2184 1288 2186
rect 1239 2183 1240 2184
rect 1234 2182 1240 2183
rect 1287 2183 1288 2184
rect 1292 2183 1293 2187
rect 1287 2182 1293 2183
rect 2318 2182 2324 2183
rect 746 2179 752 2180
rect 746 2178 747 2179
rect 676 2176 747 2178
rect 746 2175 747 2176
rect 751 2175 752 2179
rect 2318 2178 2319 2182
rect 2323 2178 2324 2182
rect 2318 2177 2324 2178
rect 2406 2182 2412 2183
rect 2406 2178 2407 2182
rect 2411 2178 2412 2182
rect 2406 2177 2412 2178
rect 2502 2182 2508 2183
rect 2502 2178 2503 2182
rect 2507 2178 2508 2182
rect 2502 2177 2508 2178
rect 2606 2182 2612 2183
rect 2606 2178 2607 2182
rect 2611 2178 2612 2182
rect 2606 2177 2612 2178
rect 2726 2182 2732 2183
rect 2726 2178 2727 2182
rect 2731 2178 2732 2182
rect 2726 2177 2732 2178
rect 2862 2182 2868 2183
rect 2862 2178 2863 2182
rect 2867 2178 2868 2182
rect 2862 2177 2868 2178
rect 3014 2182 3020 2183
rect 3014 2178 3015 2182
rect 3019 2178 3020 2182
rect 3014 2177 3020 2178
rect 3182 2182 3188 2183
rect 3182 2178 3183 2182
rect 3187 2178 3188 2182
rect 3182 2177 3188 2178
rect 3358 2182 3364 2183
rect 3358 2178 3359 2182
rect 3363 2178 3364 2182
rect 3358 2177 3364 2178
rect 3510 2182 3516 2183
rect 3510 2178 3511 2182
rect 3515 2178 3516 2182
rect 3510 2177 3516 2178
rect 746 2174 752 2175
rect 2343 2171 2349 2172
rect 2343 2167 2344 2171
rect 2348 2170 2349 2171
rect 2358 2171 2364 2172
rect 2358 2170 2359 2171
rect 2348 2168 2359 2170
rect 2348 2167 2349 2168
rect 2343 2166 2349 2167
rect 2358 2167 2359 2168
rect 2363 2167 2364 2171
rect 2358 2166 2364 2167
rect 2378 2171 2384 2172
rect 2378 2167 2379 2171
rect 2383 2170 2384 2171
rect 2431 2171 2437 2172
rect 2431 2170 2432 2171
rect 2383 2168 2432 2170
rect 2383 2167 2384 2168
rect 2378 2166 2384 2167
rect 2431 2167 2432 2168
rect 2436 2167 2437 2171
rect 2431 2166 2437 2167
rect 2470 2171 2476 2172
rect 2470 2167 2471 2171
rect 2475 2170 2476 2171
rect 2527 2171 2533 2172
rect 2527 2170 2528 2171
rect 2475 2168 2528 2170
rect 2475 2167 2476 2168
rect 2470 2166 2476 2167
rect 2527 2167 2528 2168
rect 2532 2167 2533 2171
rect 2527 2166 2533 2167
rect 2630 2171 2637 2172
rect 2630 2167 2631 2171
rect 2636 2167 2637 2171
rect 2630 2166 2637 2167
rect 2678 2171 2684 2172
rect 2678 2167 2679 2171
rect 2683 2170 2684 2171
rect 2751 2171 2757 2172
rect 2751 2170 2752 2171
rect 2683 2168 2752 2170
rect 2683 2167 2684 2168
rect 2678 2166 2684 2167
rect 2751 2167 2752 2168
rect 2756 2167 2757 2171
rect 2751 2166 2757 2167
rect 2786 2171 2792 2172
rect 2786 2167 2787 2171
rect 2791 2170 2792 2171
rect 2887 2171 2893 2172
rect 2887 2170 2888 2171
rect 2791 2168 2888 2170
rect 2791 2167 2792 2168
rect 2786 2166 2792 2167
rect 2887 2167 2888 2168
rect 2892 2167 2893 2171
rect 2887 2166 2893 2167
rect 2927 2171 2933 2172
rect 2927 2167 2928 2171
rect 2932 2170 2933 2171
rect 3039 2171 3045 2172
rect 3039 2170 3040 2171
rect 2932 2168 3040 2170
rect 2932 2167 2933 2168
rect 2927 2166 2933 2167
rect 3039 2167 3040 2168
rect 3044 2167 3045 2171
rect 3039 2166 3045 2167
rect 3074 2171 3080 2172
rect 3074 2167 3075 2171
rect 3079 2170 3080 2171
rect 3207 2171 3213 2172
rect 3207 2170 3208 2171
rect 3079 2168 3208 2170
rect 3079 2167 3080 2168
rect 3074 2166 3080 2167
rect 3207 2167 3208 2168
rect 3212 2167 3213 2171
rect 3207 2166 3213 2167
rect 3383 2171 3392 2172
rect 3383 2167 3384 2171
rect 3391 2167 3392 2171
rect 3383 2166 3392 2167
rect 3535 2171 3541 2172
rect 3535 2167 3536 2171
rect 3540 2170 3541 2171
rect 3570 2171 3576 2172
rect 3570 2170 3571 2171
rect 3540 2168 3571 2170
rect 3540 2167 3541 2168
rect 3535 2166 3541 2167
rect 3570 2167 3571 2168
rect 3575 2167 3576 2171
rect 3570 2166 3576 2167
rect 335 2163 341 2164
rect 335 2159 336 2163
rect 340 2162 341 2163
rect 414 2163 420 2164
rect 414 2162 415 2163
rect 340 2160 415 2162
rect 340 2159 341 2160
rect 335 2158 341 2159
rect 414 2159 415 2160
rect 419 2159 420 2163
rect 414 2158 420 2159
rect 431 2163 437 2164
rect 431 2159 432 2163
rect 436 2162 437 2163
rect 510 2163 516 2164
rect 510 2162 511 2163
rect 436 2160 511 2162
rect 436 2159 437 2160
rect 431 2158 437 2159
rect 510 2159 511 2160
rect 515 2159 516 2163
rect 510 2158 516 2159
rect 526 2163 533 2164
rect 526 2159 527 2163
rect 532 2159 533 2163
rect 526 2158 533 2159
rect 623 2163 629 2164
rect 623 2159 624 2163
rect 628 2162 629 2163
rect 634 2163 640 2164
rect 634 2162 635 2163
rect 628 2160 635 2162
rect 628 2159 629 2160
rect 623 2158 629 2159
rect 634 2159 635 2160
rect 639 2159 640 2163
rect 634 2158 640 2159
rect 650 2163 656 2164
rect 650 2159 651 2163
rect 655 2162 656 2163
rect 711 2163 717 2164
rect 711 2162 712 2163
rect 655 2160 712 2162
rect 655 2159 656 2160
rect 650 2158 656 2159
rect 711 2159 712 2160
rect 716 2159 717 2163
rect 711 2158 717 2159
rect 738 2163 744 2164
rect 738 2159 739 2163
rect 743 2162 744 2163
rect 799 2163 805 2164
rect 799 2162 800 2163
rect 743 2160 800 2162
rect 743 2159 744 2160
rect 738 2158 744 2159
rect 799 2159 800 2160
rect 804 2159 805 2163
rect 799 2158 805 2159
rect 887 2163 893 2164
rect 887 2159 888 2163
rect 892 2162 893 2163
rect 958 2163 964 2164
rect 958 2162 959 2163
rect 892 2160 959 2162
rect 892 2159 893 2160
rect 887 2158 893 2159
rect 958 2159 959 2160
rect 963 2159 964 2163
rect 958 2158 964 2159
rect 975 2163 981 2164
rect 975 2159 976 2163
rect 980 2162 981 2163
rect 1046 2163 1052 2164
rect 1046 2162 1047 2163
rect 980 2160 1047 2162
rect 980 2159 981 2160
rect 975 2158 981 2159
rect 1046 2159 1047 2160
rect 1051 2159 1052 2163
rect 1046 2158 1052 2159
rect 1063 2163 1069 2164
rect 1063 2159 1064 2163
rect 1068 2162 1069 2163
rect 1134 2163 1140 2164
rect 1134 2162 1135 2163
rect 1068 2160 1135 2162
rect 1068 2159 1069 2160
rect 1063 2158 1069 2159
rect 1134 2159 1135 2160
rect 1139 2159 1140 2163
rect 1134 2158 1140 2159
rect 1151 2163 1157 2164
rect 1151 2159 1152 2163
rect 1156 2162 1157 2163
rect 1230 2163 1236 2164
rect 1230 2162 1231 2163
rect 1156 2160 1231 2162
rect 1156 2159 1157 2160
rect 1151 2158 1157 2159
rect 1230 2159 1231 2160
rect 1235 2159 1236 2163
rect 1230 2158 1236 2159
rect 1242 2163 1253 2164
rect 1242 2159 1243 2163
rect 1247 2159 1248 2163
rect 1252 2159 1253 2163
rect 2398 2163 2404 2164
rect 2398 2162 2399 2163
rect 1242 2158 1253 2159
rect 2044 2160 2399 2162
rect 1927 2155 1933 2156
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 406 2154 412 2155
rect 406 2150 407 2154
rect 411 2150 412 2154
rect 406 2149 412 2150
rect 502 2154 508 2155
rect 502 2150 503 2154
rect 507 2150 508 2154
rect 502 2149 508 2150
rect 598 2154 604 2155
rect 598 2150 599 2154
rect 603 2150 604 2154
rect 598 2149 604 2150
rect 686 2154 692 2155
rect 686 2150 687 2154
rect 691 2150 692 2154
rect 686 2149 692 2150
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 862 2154 868 2155
rect 862 2150 863 2154
rect 867 2150 868 2154
rect 862 2149 868 2150
rect 950 2154 956 2155
rect 950 2150 951 2154
rect 955 2150 956 2154
rect 950 2149 956 2150
rect 1038 2154 1044 2155
rect 1038 2150 1039 2154
rect 1043 2150 1044 2154
rect 1038 2149 1044 2150
rect 1126 2154 1132 2155
rect 1126 2150 1127 2154
rect 1131 2150 1132 2154
rect 1126 2149 1132 2150
rect 1222 2154 1228 2155
rect 1222 2150 1223 2154
rect 1227 2150 1228 2154
rect 1927 2151 1928 2155
rect 1932 2154 1933 2155
rect 1990 2155 1996 2156
rect 1990 2154 1991 2155
rect 1932 2152 1991 2154
rect 1932 2151 1933 2152
rect 1927 2150 1933 2151
rect 1990 2151 1991 2152
rect 1995 2151 1996 2155
rect 1990 2150 1996 2151
rect 2007 2155 2013 2156
rect 2007 2151 2008 2155
rect 2012 2154 2013 2155
rect 2044 2154 2046 2160
rect 2398 2159 2399 2160
rect 2403 2159 2404 2163
rect 2398 2158 2404 2159
rect 2012 2152 2046 2154
rect 2050 2155 2056 2156
rect 2012 2151 2013 2152
rect 2007 2150 2013 2151
rect 2050 2151 2051 2155
rect 2055 2154 2056 2155
rect 2135 2155 2141 2156
rect 2135 2154 2136 2155
rect 2055 2152 2136 2154
rect 2055 2151 2056 2152
rect 2050 2150 2056 2151
rect 2135 2151 2136 2152
rect 2140 2151 2141 2155
rect 2135 2150 2141 2151
rect 2162 2155 2168 2156
rect 2162 2151 2163 2155
rect 2167 2154 2168 2155
rect 2271 2155 2277 2156
rect 2271 2154 2272 2155
rect 2167 2152 2272 2154
rect 2167 2151 2168 2152
rect 2162 2150 2168 2151
rect 2271 2151 2272 2152
rect 2276 2151 2277 2155
rect 2271 2150 2277 2151
rect 2298 2155 2304 2156
rect 2298 2151 2299 2155
rect 2303 2154 2304 2155
rect 2415 2155 2421 2156
rect 2415 2154 2416 2155
rect 2303 2152 2416 2154
rect 2303 2151 2304 2152
rect 2298 2150 2304 2151
rect 2415 2151 2416 2152
rect 2420 2151 2421 2155
rect 2415 2150 2421 2151
rect 2562 2155 2573 2156
rect 2562 2151 2563 2155
rect 2567 2151 2568 2155
rect 2572 2151 2573 2155
rect 2562 2150 2573 2151
rect 2719 2155 2725 2156
rect 2719 2151 2720 2155
rect 2724 2154 2725 2155
rect 2734 2155 2740 2156
rect 2734 2154 2735 2155
rect 2724 2152 2735 2154
rect 2724 2151 2725 2152
rect 2719 2150 2725 2151
rect 2734 2151 2735 2152
rect 2739 2151 2740 2155
rect 2734 2150 2740 2151
rect 2746 2155 2752 2156
rect 2746 2151 2747 2155
rect 2751 2154 2752 2155
rect 2871 2155 2877 2156
rect 2871 2154 2872 2155
rect 2751 2152 2872 2154
rect 2751 2151 2752 2152
rect 2746 2150 2752 2151
rect 2871 2151 2872 2152
rect 2876 2151 2877 2155
rect 2871 2150 2877 2151
rect 2898 2155 2904 2156
rect 2898 2151 2899 2155
rect 2903 2154 2904 2155
rect 3031 2155 3037 2156
rect 3031 2154 3032 2155
rect 2903 2152 3032 2154
rect 2903 2151 2904 2152
rect 2898 2150 2904 2151
rect 3031 2151 3032 2152
rect 3036 2151 3037 2155
rect 3031 2150 3037 2151
rect 3058 2155 3064 2156
rect 3058 2151 3059 2155
rect 3063 2154 3064 2155
rect 3199 2155 3205 2156
rect 3199 2154 3200 2155
rect 3063 2152 3200 2154
rect 3063 2151 3064 2152
rect 3058 2150 3064 2151
rect 3199 2151 3200 2152
rect 3204 2151 3205 2155
rect 3199 2150 3205 2151
rect 3226 2155 3232 2156
rect 3226 2151 3227 2155
rect 3231 2154 3232 2155
rect 3375 2155 3381 2156
rect 3375 2154 3376 2155
rect 3231 2152 3376 2154
rect 3231 2151 3232 2152
rect 3226 2150 3232 2151
rect 3375 2151 3376 2152
rect 3380 2151 3381 2155
rect 3375 2150 3381 2151
rect 3535 2155 3541 2156
rect 3535 2151 3536 2155
rect 3540 2154 3541 2155
rect 3562 2155 3568 2156
rect 3562 2154 3563 2155
rect 3540 2152 3563 2154
rect 3540 2151 3541 2152
rect 3535 2150 3541 2151
rect 3562 2151 3563 2152
rect 3567 2151 3568 2155
rect 3562 2150 3568 2151
rect 1222 2149 1228 2150
rect 1902 2146 1908 2147
rect 1902 2142 1903 2146
rect 1907 2142 1908 2146
rect 1902 2141 1908 2142
rect 1982 2146 1988 2147
rect 1982 2142 1983 2146
rect 1987 2142 1988 2146
rect 1982 2141 1988 2142
rect 2110 2146 2116 2147
rect 2110 2142 2111 2146
rect 2115 2142 2116 2146
rect 2110 2141 2116 2142
rect 2246 2146 2252 2147
rect 2246 2142 2247 2146
rect 2251 2142 2252 2146
rect 2246 2141 2252 2142
rect 2390 2146 2396 2147
rect 2390 2142 2391 2146
rect 2395 2142 2396 2146
rect 2390 2141 2396 2142
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2694 2146 2700 2147
rect 2694 2142 2695 2146
rect 2699 2142 2700 2146
rect 2694 2141 2700 2142
rect 2846 2146 2852 2147
rect 2846 2142 2847 2146
rect 2851 2142 2852 2146
rect 2846 2141 2852 2142
rect 3006 2146 3012 2147
rect 3006 2142 3007 2146
rect 3011 2142 3012 2146
rect 3006 2141 3012 2142
rect 3174 2146 3180 2147
rect 3174 2142 3175 2146
rect 3179 2142 3180 2146
rect 3174 2141 3180 2142
rect 3350 2146 3356 2147
rect 3350 2142 3351 2146
rect 3355 2142 3356 2146
rect 3350 2141 3356 2142
rect 3510 2146 3516 2147
rect 3510 2142 3511 2146
rect 3515 2142 3516 2146
rect 3510 2141 3516 2142
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 1830 2136 1836 2137
rect 1830 2132 1831 2136
rect 1835 2132 1836 2136
rect 1830 2131 1836 2132
rect 1870 2128 1876 2129
rect 414 2127 420 2128
rect 414 2123 415 2127
rect 419 2123 420 2127
rect 414 2122 420 2123
rect 510 2127 516 2128
rect 510 2123 511 2127
rect 515 2123 516 2127
rect 510 2122 516 2123
rect 650 2127 656 2128
rect 650 2123 651 2127
rect 655 2123 656 2127
rect 650 2122 656 2123
rect 738 2127 744 2128
rect 738 2123 739 2127
rect 743 2123 744 2127
rect 738 2122 744 2123
rect 746 2127 752 2128
rect 746 2123 747 2127
rect 751 2126 752 2127
rect 886 2127 892 2128
rect 751 2124 785 2126
rect 751 2123 752 2124
rect 746 2122 752 2123
rect 886 2123 887 2127
rect 891 2123 892 2127
rect 886 2122 892 2123
rect 958 2127 964 2128
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 958 2122 964 2123
rect 1046 2127 1052 2128
rect 1046 2123 1047 2127
rect 1051 2123 1052 2127
rect 1046 2122 1052 2123
rect 1134 2127 1140 2128
rect 1134 2123 1135 2127
rect 1139 2123 1140 2127
rect 1134 2122 1140 2123
rect 1230 2127 1236 2128
rect 1230 2123 1231 2127
rect 1235 2123 1236 2127
rect 1870 2124 1871 2128
rect 1875 2124 1876 2128
rect 1870 2123 1876 2124
rect 3590 2128 3596 2129
rect 3590 2124 3591 2128
rect 3595 2124 3596 2128
rect 3590 2123 3596 2124
rect 1230 2122 1236 2123
rect 110 2119 116 2120
rect 110 2115 111 2119
rect 115 2115 116 2119
rect 1830 2119 1836 2120
rect 110 2114 116 2115
rect 302 2116 308 2117
rect 302 2112 303 2116
rect 307 2112 308 2116
rect 302 2111 308 2112
rect 398 2116 404 2117
rect 398 2112 399 2116
rect 403 2112 404 2116
rect 398 2111 404 2112
rect 494 2116 500 2117
rect 494 2112 495 2116
rect 499 2112 500 2116
rect 494 2111 500 2112
rect 590 2116 596 2117
rect 590 2112 591 2116
rect 595 2112 596 2116
rect 590 2111 596 2112
rect 678 2116 684 2117
rect 678 2112 679 2116
rect 683 2112 684 2116
rect 678 2111 684 2112
rect 766 2116 772 2117
rect 766 2112 767 2116
rect 771 2112 772 2116
rect 766 2111 772 2112
rect 854 2116 860 2117
rect 854 2112 855 2116
rect 859 2112 860 2116
rect 854 2111 860 2112
rect 942 2116 948 2117
rect 942 2112 943 2116
rect 947 2112 948 2116
rect 942 2111 948 2112
rect 1030 2116 1036 2117
rect 1030 2112 1031 2116
rect 1035 2112 1036 2116
rect 1030 2111 1036 2112
rect 1118 2116 1124 2117
rect 1118 2112 1119 2116
rect 1123 2112 1124 2116
rect 1118 2111 1124 2112
rect 1214 2116 1220 2117
rect 1214 2112 1215 2116
rect 1219 2112 1220 2116
rect 1830 2115 1831 2119
rect 1835 2115 1836 2119
rect 1830 2114 1836 2115
rect 1990 2119 1996 2120
rect 1990 2115 1991 2119
rect 1995 2115 1996 2119
rect 1990 2114 1996 2115
rect 2162 2119 2168 2120
rect 2162 2115 2163 2119
rect 2167 2115 2168 2119
rect 2162 2114 2168 2115
rect 2298 2119 2304 2120
rect 2298 2115 2299 2119
rect 2303 2115 2304 2119
rect 2298 2114 2304 2115
rect 2398 2119 2404 2120
rect 2398 2115 2399 2119
rect 2403 2115 2404 2119
rect 2398 2114 2404 2115
rect 2746 2119 2752 2120
rect 2746 2115 2747 2119
rect 2751 2115 2752 2119
rect 2746 2114 2752 2115
rect 2898 2119 2904 2120
rect 2898 2115 2899 2119
rect 2903 2115 2904 2119
rect 2898 2114 2904 2115
rect 3058 2119 3064 2120
rect 3058 2115 3059 2119
rect 3063 2115 3064 2119
rect 3058 2114 3064 2115
rect 3226 2119 3232 2120
rect 3226 2115 3227 2119
rect 3231 2115 3232 2119
rect 3226 2114 3232 2115
rect 3534 2119 3540 2120
rect 3534 2115 3535 2119
rect 3539 2115 3540 2119
rect 3534 2114 3540 2115
rect 1214 2111 1220 2112
rect 1870 2111 1876 2112
rect 1870 2107 1871 2111
rect 1875 2107 1876 2111
rect 3590 2111 3596 2112
rect 1870 2106 1876 2107
rect 1894 2108 1900 2109
rect 1894 2104 1895 2108
rect 1899 2104 1900 2108
rect 1894 2103 1900 2104
rect 1974 2108 1980 2109
rect 1974 2104 1975 2108
rect 1979 2104 1980 2108
rect 1974 2103 1980 2104
rect 2102 2108 2108 2109
rect 2102 2104 2103 2108
rect 2107 2104 2108 2108
rect 2102 2103 2108 2104
rect 2238 2108 2244 2109
rect 2238 2104 2239 2108
rect 2243 2104 2244 2108
rect 2238 2103 2244 2104
rect 2382 2108 2388 2109
rect 2382 2104 2383 2108
rect 2387 2104 2388 2108
rect 2382 2103 2388 2104
rect 2534 2108 2540 2109
rect 2534 2104 2535 2108
rect 2539 2104 2540 2108
rect 2534 2103 2540 2104
rect 2686 2108 2692 2109
rect 2686 2104 2687 2108
rect 2691 2104 2692 2108
rect 2686 2103 2692 2104
rect 2838 2108 2844 2109
rect 2838 2104 2839 2108
rect 2843 2104 2844 2108
rect 2838 2103 2844 2104
rect 2998 2108 3004 2109
rect 2998 2104 2999 2108
rect 3003 2104 3004 2108
rect 2998 2103 3004 2104
rect 3166 2108 3172 2109
rect 3166 2104 3167 2108
rect 3171 2104 3172 2108
rect 3166 2103 3172 2104
rect 3342 2108 3348 2109
rect 3342 2104 3343 2108
rect 3347 2104 3348 2108
rect 3342 2103 3348 2104
rect 3502 2108 3508 2109
rect 3502 2104 3503 2108
rect 3507 2104 3508 2108
rect 3590 2107 3591 2111
rect 3595 2107 3596 2111
rect 3590 2106 3596 2107
rect 3502 2103 3508 2104
rect 242 2099 248 2100
rect 242 2095 243 2099
rect 247 2098 248 2099
rect 319 2099 325 2100
rect 319 2098 320 2099
rect 247 2096 320 2098
rect 247 2095 248 2096
rect 242 2094 248 2095
rect 319 2095 320 2096
rect 324 2095 325 2099
rect 319 2094 325 2095
rect 1778 2091 1784 2092
rect 1778 2087 1779 2091
rect 1783 2090 1784 2091
rect 1911 2091 1917 2092
rect 1911 2090 1912 2091
rect 1783 2088 1912 2090
rect 1783 2087 1784 2088
rect 1778 2086 1784 2087
rect 1911 2087 1912 2088
rect 1916 2087 1917 2091
rect 1911 2086 1917 2087
rect 2482 2091 2488 2092
rect 2482 2087 2483 2091
rect 2487 2090 2488 2091
rect 2551 2091 2557 2092
rect 2551 2090 2552 2091
rect 2487 2088 2552 2090
rect 2487 2087 2488 2088
rect 2482 2086 2488 2087
rect 2551 2087 2552 2088
rect 2556 2087 2557 2091
rect 2551 2086 2557 2087
rect 3306 2091 3312 2092
rect 3306 2087 3307 2091
rect 3311 2090 3312 2091
rect 3359 2091 3365 2092
rect 3359 2090 3360 2091
rect 3311 2088 3360 2090
rect 3311 2087 3312 2088
rect 3306 2086 3312 2087
rect 3359 2087 3360 2088
rect 3364 2087 3365 2091
rect 3359 2086 3365 2087
rect 206 2060 212 2061
rect 110 2057 116 2058
rect 110 2053 111 2057
rect 115 2053 116 2057
rect 206 2056 207 2060
rect 211 2056 212 2060
rect 206 2055 212 2056
rect 326 2060 332 2061
rect 326 2056 327 2060
rect 331 2056 332 2060
rect 326 2055 332 2056
rect 446 2060 452 2061
rect 446 2056 447 2060
rect 451 2056 452 2060
rect 446 2055 452 2056
rect 574 2060 580 2061
rect 574 2056 575 2060
rect 579 2056 580 2060
rect 574 2055 580 2056
rect 702 2060 708 2061
rect 702 2056 703 2060
rect 707 2056 708 2060
rect 702 2055 708 2056
rect 822 2060 828 2061
rect 822 2056 823 2060
rect 827 2056 828 2060
rect 822 2055 828 2056
rect 942 2060 948 2061
rect 942 2056 943 2060
rect 947 2056 948 2060
rect 942 2055 948 2056
rect 1062 2060 1068 2061
rect 1062 2056 1063 2060
rect 1067 2056 1068 2060
rect 1062 2055 1068 2056
rect 1174 2060 1180 2061
rect 1174 2056 1175 2060
rect 1179 2056 1180 2060
rect 1174 2055 1180 2056
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1374 2060 1380 2061
rect 1374 2056 1375 2060
rect 1379 2056 1380 2060
rect 1374 2055 1380 2056
rect 1470 2060 1476 2061
rect 1470 2056 1471 2060
rect 1475 2056 1476 2060
rect 1470 2055 1476 2056
rect 1566 2060 1572 2061
rect 1566 2056 1567 2060
rect 1571 2056 1572 2060
rect 1566 2055 1572 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 1830 2057 1836 2058
rect 110 2052 116 2053
rect 1830 2053 1831 2057
rect 1835 2053 1836 2057
rect 1966 2056 1972 2057
rect 1830 2052 1836 2053
rect 1870 2053 1876 2054
rect 274 2051 280 2052
rect 274 2050 275 2051
rect 269 2048 275 2050
rect 274 2047 275 2048
rect 279 2047 280 2051
rect 394 2051 400 2052
rect 274 2046 280 2047
rect 388 2044 390 2049
rect 394 2047 395 2051
rect 399 2050 400 2051
rect 642 2051 648 2052
rect 399 2048 465 2050
rect 399 2047 400 2048
rect 394 2046 400 2047
rect 636 2044 638 2049
rect 642 2047 643 2051
rect 647 2050 648 2051
rect 770 2051 776 2052
rect 647 2048 721 2050
rect 647 2047 648 2048
rect 642 2046 648 2047
rect 770 2047 771 2051
rect 775 2050 776 2051
rect 1030 2051 1036 2052
rect 1030 2050 1031 2051
rect 775 2048 841 2050
rect 1005 2048 1031 2050
rect 775 2047 776 2048
rect 770 2046 776 2047
rect 1030 2047 1031 2048
rect 1035 2047 1036 2051
rect 1130 2051 1136 2052
rect 1130 2050 1131 2051
rect 1125 2048 1131 2050
rect 1030 2046 1036 2047
rect 1130 2047 1131 2048
rect 1135 2047 1136 2051
rect 1242 2051 1248 2052
rect 1242 2050 1243 2051
rect 1237 2048 1243 2050
rect 1130 2046 1136 2047
rect 1242 2047 1243 2048
rect 1247 2047 1248 2051
rect 1346 2051 1352 2052
rect 1242 2046 1248 2047
rect 1340 2044 1342 2049
rect 1346 2047 1347 2051
rect 1351 2050 1352 2051
rect 1442 2051 1448 2052
rect 1351 2048 1393 2050
rect 1351 2047 1352 2048
rect 1346 2046 1352 2047
rect 1442 2047 1443 2051
rect 1447 2050 1448 2051
rect 1538 2051 1544 2052
rect 1447 2048 1489 2050
rect 1447 2047 1448 2048
rect 1442 2046 1448 2047
rect 1538 2047 1539 2051
rect 1543 2050 1544 2051
rect 1634 2051 1640 2052
rect 1543 2048 1585 2050
rect 1543 2047 1544 2048
rect 1538 2046 1544 2047
rect 1634 2047 1635 2051
rect 1639 2050 1640 2051
rect 1730 2051 1736 2052
rect 1639 2048 1681 2050
rect 1639 2047 1640 2048
rect 1634 2046 1640 2047
rect 1730 2047 1731 2051
rect 1735 2050 1736 2051
rect 1735 2048 1761 2050
rect 1870 2049 1871 2053
rect 1875 2049 1876 2053
rect 1966 2052 1967 2056
rect 1971 2052 1972 2056
rect 1966 2051 1972 2052
rect 2214 2056 2220 2057
rect 2214 2052 2215 2056
rect 2219 2052 2220 2056
rect 2214 2051 2220 2052
rect 2446 2056 2452 2057
rect 2446 2052 2447 2056
rect 2451 2052 2452 2056
rect 2446 2051 2452 2052
rect 2654 2056 2660 2057
rect 2654 2052 2655 2056
rect 2659 2052 2660 2056
rect 2654 2051 2660 2052
rect 2838 2056 2844 2057
rect 2838 2052 2839 2056
rect 2843 2052 2844 2056
rect 2838 2051 2844 2052
rect 2998 2056 3004 2057
rect 2998 2052 2999 2056
rect 3003 2052 3004 2056
rect 2998 2051 3004 2052
rect 3142 2056 3148 2057
rect 3142 2052 3143 2056
rect 3147 2052 3148 2056
rect 3142 2051 3148 2052
rect 3270 2056 3276 2057
rect 3270 2052 3271 2056
rect 3275 2052 3276 2056
rect 3270 2051 3276 2052
rect 3398 2056 3404 2057
rect 3398 2052 3399 2056
rect 3403 2052 3404 2056
rect 3398 2051 3404 2052
rect 3502 2056 3508 2057
rect 3502 2052 3503 2056
rect 3507 2052 3508 2056
rect 3502 2051 3508 2052
rect 3590 2053 3596 2054
rect 1870 2048 1876 2049
rect 3590 2049 3591 2053
rect 3595 2049 3596 2053
rect 3590 2048 3596 2049
rect 1735 2047 1736 2048
rect 1730 2046 1736 2047
rect 2050 2047 2056 2048
rect 2050 2046 2051 2047
rect 2029 2044 2051 2046
rect 386 2043 392 2044
rect 110 2040 116 2041
rect 110 2036 111 2040
rect 115 2036 116 2040
rect 386 2039 387 2043
rect 391 2039 392 2043
rect 386 2038 392 2039
rect 634 2043 640 2044
rect 634 2039 635 2043
rect 639 2039 640 2043
rect 634 2038 640 2039
rect 1338 2043 1344 2044
rect 1338 2039 1339 2043
rect 1343 2039 1344 2043
rect 2050 2043 2051 2044
rect 2055 2043 2056 2047
rect 2282 2047 2288 2048
rect 2050 2042 2056 2043
rect 1338 2038 1344 2039
rect 1830 2040 1836 2041
rect 2276 2040 2278 2045
rect 2282 2043 2283 2047
rect 2287 2046 2288 2047
rect 2754 2047 2760 2048
rect 2754 2046 2755 2047
rect 2287 2044 2465 2046
rect 2717 2044 2755 2046
rect 2287 2043 2288 2044
rect 2282 2042 2288 2043
rect 2754 2043 2755 2044
rect 2759 2043 2760 2047
rect 2942 2047 2948 2048
rect 2942 2046 2943 2047
rect 2901 2044 2943 2046
rect 2754 2042 2760 2043
rect 2942 2043 2943 2044
rect 2947 2043 2948 2047
rect 3078 2047 3084 2048
rect 3078 2046 3079 2047
rect 3061 2044 3079 2046
rect 2942 2042 2948 2043
rect 3078 2043 3079 2044
rect 3083 2043 3084 2047
rect 3078 2042 3084 2043
rect 3086 2047 3092 2048
rect 3086 2043 3087 2047
rect 3091 2046 3092 2047
rect 3210 2047 3216 2048
rect 3091 2044 3161 2046
rect 3091 2043 3092 2044
rect 3086 2042 3092 2043
rect 3210 2043 3211 2047
rect 3215 2046 3216 2047
rect 3386 2047 3392 2048
rect 3215 2044 3289 2046
rect 3215 2043 3216 2044
rect 3210 2042 3216 2043
rect 3386 2043 3387 2047
rect 3391 2046 3392 2047
rect 3391 2044 3417 2046
rect 3391 2043 3392 2044
rect 3386 2042 3392 2043
rect 3564 2040 3566 2045
rect 110 2035 116 2036
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 2274 2039 2280 2040
rect 1830 2035 1836 2036
rect 1870 2036 1876 2037
rect 1870 2032 1871 2036
rect 1875 2032 1876 2036
rect 2274 2035 2275 2039
rect 2279 2035 2280 2039
rect 2274 2034 2280 2035
rect 3562 2039 3568 2040
rect 3562 2035 3563 2039
rect 3567 2035 3568 2039
rect 3562 2034 3568 2035
rect 3590 2036 3596 2037
rect 1870 2031 1876 2032
rect 3590 2032 3591 2036
rect 3595 2032 3596 2036
rect 3590 2031 3596 2032
rect 214 2022 220 2023
rect 214 2018 215 2022
rect 219 2018 220 2022
rect 214 2017 220 2018
rect 334 2022 340 2023
rect 334 2018 335 2022
rect 339 2018 340 2022
rect 334 2017 340 2018
rect 454 2022 460 2023
rect 454 2018 455 2022
rect 459 2018 460 2022
rect 454 2017 460 2018
rect 582 2022 588 2023
rect 582 2018 583 2022
rect 587 2018 588 2022
rect 582 2017 588 2018
rect 710 2022 716 2023
rect 710 2018 711 2022
rect 715 2018 716 2022
rect 710 2017 716 2018
rect 830 2022 836 2023
rect 830 2018 831 2022
rect 835 2018 836 2022
rect 830 2017 836 2018
rect 950 2022 956 2023
rect 950 2018 951 2022
rect 955 2018 956 2022
rect 950 2017 956 2018
rect 1070 2022 1076 2023
rect 1070 2018 1071 2022
rect 1075 2018 1076 2022
rect 1070 2017 1076 2018
rect 1182 2022 1188 2023
rect 1182 2018 1183 2022
rect 1187 2018 1188 2022
rect 1182 2017 1188 2018
rect 1286 2022 1292 2023
rect 1286 2018 1287 2022
rect 1291 2018 1292 2022
rect 1286 2017 1292 2018
rect 1382 2022 1388 2023
rect 1382 2018 1383 2022
rect 1387 2018 1388 2022
rect 1382 2017 1388 2018
rect 1478 2022 1484 2023
rect 1478 2018 1479 2022
rect 1483 2018 1484 2022
rect 1478 2017 1484 2018
rect 1574 2022 1580 2023
rect 1574 2018 1575 2022
rect 1579 2018 1580 2022
rect 1574 2017 1580 2018
rect 1670 2022 1676 2023
rect 1670 2018 1671 2022
rect 1675 2018 1676 2022
rect 1670 2017 1676 2018
rect 1750 2022 1756 2023
rect 1750 2018 1751 2022
rect 1755 2018 1756 2022
rect 1750 2017 1756 2018
rect 1974 2018 1980 2019
rect 1974 2014 1975 2018
rect 1979 2014 1980 2018
rect 1974 2013 1980 2014
rect 2222 2018 2228 2019
rect 2222 2014 2223 2018
rect 2227 2014 2228 2018
rect 2222 2013 2228 2014
rect 2454 2018 2460 2019
rect 2454 2014 2455 2018
rect 2459 2014 2460 2018
rect 2454 2013 2460 2014
rect 2662 2018 2668 2019
rect 2662 2014 2663 2018
rect 2667 2014 2668 2018
rect 2662 2013 2668 2014
rect 2846 2018 2852 2019
rect 2846 2014 2847 2018
rect 2851 2014 2852 2018
rect 2846 2013 2852 2014
rect 3006 2018 3012 2019
rect 3006 2014 3007 2018
rect 3011 2014 3012 2018
rect 3006 2013 3012 2014
rect 3150 2018 3156 2019
rect 3150 2014 3151 2018
rect 3155 2014 3156 2018
rect 3150 2013 3156 2014
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3406 2018 3412 2019
rect 3406 2014 3407 2018
rect 3411 2014 3412 2018
rect 3406 2013 3412 2014
rect 3510 2018 3516 2019
rect 3510 2014 3511 2018
rect 3515 2014 3516 2018
rect 3510 2013 3516 2014
rect 239 2011 248 2012
rect 239 2007 240 2011
rect 247 2007 248 2011
rect 239 2006 248 2007
rect 274 2011 280 2012
rect 274 2007 275 2011
rect 279 2010 280 2011
rect 359 2011 365 2012
rect 359 2010 360 2011
rect 279 2008 360 2010
rect 279 2007 280 2008
rect 274 2006 280 2007
rect 359 2007 360 2008
rect 364 2007 365 2011
rect 359 2006 365 2007
rect 386 2011 392 2012
rect 386 2007 387 2011
rect 391 2010 392 2011
rect 479 2011 485 2012
rect 479 2010 480 2011
rect 391 2008 480 2010
rect 391 2007 392 2008
rect 386 2006 392 2007
rect 479 2007 480 2008
rect 484 2007 485 2011
rect 479 2006 485 2007
rect 607 2011 613 2012
rect 607 2007 608 2011
rect 612 2010 613 2011
rect 642 2011 648 2012
rect 642 2010 643 2011
rect 612 2008 643 2010
rect 612 2007 613 2008
rect 607 2006 613 2007
rect 642 2007 643 2008
rect 647 2007 648 2011
rect 642 2006 648 2007
rect 735 2011 741 2012
rect 735 2007 736 2011
rect 740 2010 741 2011
rect 770 2011 776 2012
rect 770 2010 771 2011
rect 740 2008 771 2010
rect 740 2007 741 2008
rect 735 2006 741 2007
rect 770 2007 771 2008
rect 775 2007 776 2011
rect 770 2006 776 2007
rect 854 2011 861 2012
rect 854 2007 855 2011
rect 860 2007 861 2011
rect 854 2006 861 2007
rect 975 2011 981 2012
rect 975 2007 976 2011
rect 980 2010 981 2011
rect 1022 2011 1028 2012
rect 1022 2010 1023 2011
rect 980 2008 1023 2010
rect 980 2007 981 2008
rect 975 2006 981 2007
rect 1022 2007 1023 2008
rect 1027 2007 1028 2011
rect 1022 2006 1028 2007
rect 1030 2011 1036 2012
rect 1030 2007 1031 2011
rect 1035 2010 1036 2011
rect 1095 2011 1101 2012
rect 1095 2010 1096 2011
rect 1035 2008 1096 2010
rect 1035 2007 1036 2008
rect 1030 2006 1036 2007
rect 1095 2007 1096 2008
rect 1100 2007 1101 2011
rect 1095 2006 1101 2007
rect 1130 2011 1136 2012
rect 1130 2007 1131 2011
rect 1135 2010 1136 2011
rect 1207 2011 1213 2012
rect 1207 2010 1208 2011
rect 1135 2008 1208 2010
rect 1135 2007 1136 2008
rect 1130 2006 1136 2007
rect 1207 2007 1208 2008
rect 1212 2007 1213 2011
rect 1207 2006 1213 2007
rect 1311 2011 1317 2012
rect 1311 2007 1312 2011
rect 1316 2010 1317 2011
rect 1346 2011 1352 2012
rect 1346 2010 1347 2011
rect 1316 2008 1347 2010
rect 1316 2007 1317 2008
rect 1311 2006 1317 2007
rect 1346 2007 1347 2008
rect 1351 2007 1352 2011
rect 1346 2006 1352 2007
rect 1407 2011 1413 2012
rect 1407 2007 1408 2011
rect 1412 2010 1413 2011
rect 1442 2011 1448 2012
rect 1442 2010 1443 2011
rect 1412 2008 1443 2010
rect 1412 2007 1413 2008
rect 1407 2006 1413 2007
rect 1442 2007 1443 2008
rect 1447 2007 1448 2011
rect 1442 2006 1448 2007
rect 1503 2011 1509 2012
rect 1503 2007 1504 2011
rect 1508 2010 1509 2011
rect 1538 2011 1544 2012
rect 1538 2010 1539 2011
rect 1508 2008 1539 2010
rect 1508 2007 1509 2008
rect 1503 2006 1509 2007
rect 1538 2007 1539 2008
rect 1543 2007 1544 2011
rect 1538 2006 1544 2007
rect 1599 2011 1605 2012
rect 1599 2007 1600 2011
rect 1604 2010 1605 2011
rect 1634 2011 1640 2012
rect 1634 2010 1635 2011
rect 1604 2008 1635 2010
rect 1604 2007 1605 2008
rect 1599 2006 1605 2007
rect 1634 2007 1635 2008
rect 1639 2007 1640 2011
rect 1634 2006 1640 2007
rect 1695 2011 1701 2012
rect 1695 2007 1696 2011
rect 1700 2010 1701 2011
rect 1730 2011 1736 2012
rect 1730 2010 1731 2011
rect 1700 2008 1731 2010
rect 1700 2007 1701 2008
rect 1695 2006 1701 2007
rect 1730 2007 1731 2008
rect 1735 2007 1736 2011
rect 1730 2006 1736 2007
rect 1775 2011 1784 2012
rect 1775 2007 1776 2011
rect 1783 2007 1784 2011
rect 1775 2006 1784 2007
rect 1998 2007 2005 2008
rect 1998 2003 1999 2007
rect 2004 2003 2005 2007
rect 1998 2002 2005 2003
rect 2247 2007 2253 2008
rect 2247 2003 2248 2007
rect 2252 2006 2253 2007
rect 2282 2007 2288 2008
rect 2282 2006 2283 2007
rect 2252 2004 2283 2006
rect 2252 2003 2253 2004
rect 2247 2002 2253 2003
rect 2282 2003 2283 2004
rect 2287 2003 2288 2007
rect 2282 2002 2288 2003
rect 2479 2007 2488 2008
rect 2479 2003 2480 2007
rect 2487 2003 2488 2007
rect 2479 2002 2488 2003
rect 2686 2007 2693 2008
rect 2686 2003 2687 2007
rect 2692 2003 2693 2007
rect 2686 2002 2693 2003
rect 2754 2007 2760 2008
rect 2754 2003 2755 2007
rect 2759 2006 2760 2007
rect 2871 2007 2877 2008
rect 2871 2006 2872 2007
rect 2759 2004 2872 2006
rect 2759 2003 2760 2004
rect 2754 2002 2760 2003
rect 2871 2003 2872 2004
rect 2876 2003 2877 2007
rect 2871 2002 2877 2003
rect 2942 2007 2948 2008
rect 2942 2003 2943 2007
rect 2947 2006 2948 2007
rect 3031 2007 3037 2008
rect 3031 2006 3032 2007
rect 2947 2004 3032 2006
rect 2947 2003 2948 2004
rect 2942 2002 2948 2003
rect 3031 2003 3032 2004
rect 3036 2003 3037 2007
rect 3175 2007 3181 2008
rect 3031 2002 3037 2003
rect 3166 2003 3172 2004
rect 3166 2002 3167 2003
rect 3072 2000 3167 2002
rect 215 1995 221 1996
rect 215 1991 216 1995
rect 220 1994 221 1995
rect 358 1995 364 1996
rect 358 1994 359 1995
rect 220 1992 359 1994
rect 220 1991 221 1992
rect 215 1990 221 1991
rect 358 1991 359 1992
rect 363 1991 364 1995
rect 358 1990 364 1991
rect 375 1995 381 1996
rect 375 1991 376 1995
rect 380 1994 381 1995
rect 394 1995 400 1996
rect 394 1994 395 1995
rect 380 1992 395 1994
rect 380 1991 381 1992
rect 375 1990 381 1991
rect 394 1991 395 1992
rect 399 1991 400 1995
rect 394 1990 400 1991
rect 534 1995 540 1996
rect 534 1991 535 1995
rect 539 1994 540 1995
rect 543 1995 549 1996
rect 543 1994 544 1995
rect 539 1992 544 1994
rect 539 1991 540 1992
rect 534 1990 540 1991
rect 543 1991 544 1992
rect 548 1991 549 1995
rect 543 1990 549 1991
rect 570 1995 576 1996
rect 570 1991 571 1995
rect 575 1994 576 1995
rect 711 1995 717 1996
rect 711 1994 712 1995
rect 575 1992 712 1994
rect 575 1991 576 1992
rect 570 1990 576 1991
rect 711 1991 712 1992
rect 716 1991 717 1995
rect 711 1990 717 1991
rect 738 1995 744 1996
rect 738 1991 739 1995
rect 743 1994 744 1995
rect 879 1995 885 1996
rect 879 1994 880 1995
rect 743 1992 880 1994
rect 743 1991 744 1992
rect 738 1990 744 1991
rect 879 1991 880 1992
rect 884 1991 885 1995
rect 879 1990 885 1991
rect 1039 1995 1045 1996
rect 1039 1991 1040 1995
rect 1044 1994 1045 1995
rect 1174 1995 1180 1996
rect 1174 1994 1175 1995
rect 1044 1992 1175 1994
rect 1044 1991 1045 1992
rect 1039 1990 1045 1991
rect 1174 1991 1175 1992
rect 1179 1991 1180 1995
rect 1174 1990 1180 1991
rect 1191 1995 1197 1996
rect 1191 1991 1192 1995
rect 1196 1994 1197 1995
rect 1218 1995 1224 1996
rect 1218 1994 1219 1995
rect 1196 1992 1219 1994
rect 1196 1991 1197 1992
rect 1191 1990 1197 1991
rect 1218 1991 1219 1992
rect 1223 1991 1224 1995
rect 1218 1990 1224 1991
rect 1335 1995 1344 1996
rect 1335 1991 1336 1995
rect 1343 1991 1344 1995
rect 1335 1990 1344 1991
rect 1362 1995 1368 1996
rect 1362 1991 1363 1995
rect 1367 1994 1368 1995
rect 1471 1995 1477 1996
rect 1471 1994 1472 1995
rect 1367 1992 1472 1994
rect 1367 1991 1368 1992
rect 1362 1990 1368 1991
rect 1471 1991 1472 1992
rect 1476 1991 1477 1995
rect 1471 1990 1477 1991
rect 1498 1995 1504 1996
rect 1498 1991 1499 1995
rect 1503 1994 1504 1995
rect 1607 1995 1613 1996
rect 1607 1994 1608 1995
rect 1503 1992 1608 1994
rect 1503 1991 1504 1992
rect 1498 1990 1504 1991
rect 1607 1991 1608 1992
rect 1612 1991 1613 1995
rect 1607 1990 1613 1991
rect 1634 1995 1640 1996
rect 1634 1991 1635 1995
rect 1639 1994 1640 1995
rect 1743 1995 1749 1996
rect 1743 1994 1744 1995
rect 1639 1992 1744 1994
rect 1639 1991 1640 1992
rect 1634 1990 1640 1991
rect 1743 1991 1744 1992
rect 1748 1991 1749 1995
rect 1743 1990 1749 1991
rect 1983 1995 1989 1996
rect 1983 1991 1984 1995
rect 1988 1994 1989 1995
rect 2086 1995 2092 1996
rect 2086 1994 2087 1995
rect 1988 1992 2087 1994
rect 1988 1991 1989 1992
rect 1983 1990 1989 1991
rect 2086 1991 2087 1992
rect 2091 1991 2092 1995
rect 2086 1990 2092 1991
rect 2103 1995 2109 1996
rect 2103 1991 2104 1995
rect 2108 1994 2109 1995
rect 2206 1995 2212 1996
rect 2206 1994 2207 1995
rect 2108 1992 2207 1994
rect 2108 1991 2109 1992
rect 2103 1990 2109 1991
rect 2206 1991 2207 1992
rect 2211 1991 2212 1995
rect 2223 1995 2229 1996
rect 2223 1992 2224 1995
rect 2206 1990 2212 1991
rect 2222 1991 2224 1992
rect 2228 1991 2229 1995
rect 2222 1987 2223 1991
rect 2227 1990 2229 1991
rect 2274 1995 2280 1996
rect 2274 1991 2275 1995
rect 2279 1994 2280 1995
rect 2343 1995 2349 1996
rect 2343 1994 2344 1995
rect 2279 1992 2344 1994
rect 2279 1991 2280 1992
rect 2274 1990 2280 1991
rect 2343 1991 2344 1992
rect 2348 1991 2349 1995
rect 2343 1990 2349 1991
rect 2471 1995 2477 1996
rect 2471 1991 2472 1995
rect 2476 1994 2477 1995
rect 2590 1995 2596 1996
rect 2590 1994 2591 1995
rect 2476 1992 2591 1994
rect 2476 1991 2477 1992
rect 2471 1990 2477 1991
rect 2590 1991 2591 1992
rect 2595 1991 2596 1995
rect 2590 1990 2596 1991
rect 2607 1995 2613 1996
rect 2607 1991 2608 1995
rect 2612 1994 2613 1995
rect 2750 1995 2756 1996
rect 2750 1994 2751 1995
rect 2612 1992 2751 1994
rect 2612 1991 2613 1992
rect 2607 1990 2613 1991
rect 2750 1991 2751 1992
rect 2755 1991 2756 1995
rect 2750 1990 2756 1991
rect 2767 1995 2773 1996
rect 2767 1991 2768 1995
rect 2772 1994 2773 1995
rect 2926 1995 2932 1996
rect 2926 1994 2927 1995
rect 2772 1992 2927 1994
rect 2772 1991 2773 1992
rect 2767 1990 2773 1991
rect 2926 1991 2927 1992
rect 2931 1991 2932 1995
rect 2926 1990 2932 1991
rect 2943 1995 2949 1996
rect 2943 1991 2944 1995
rect 2948 1994 2949 1995
rect 3072 1994 3074 2000
rect 3166 1999 3167 2000
rect 3171 1999 3172 2003
rect 3175 2003 3176 2007
rect 3180 2006 3181 2007
rect 3210 2007 3216 2008
rect 3210 2006 3211 2007
rect 3180 2004 3211 2006
rect 3180 2003 3181 2004
rect 3175 2002 3181 2003
rect 3210 2003 3211 2004
rect 3215 2003 3216 2007
rect 3210 2002 3216 2003
rect 3303 2007 3312 2008
rect 3303 2003 3304 2007
rect 3311 2003 3312 2007
rect 3303 2002 3312 2003
rect 3431 2007 3437 2008
rect 3431 2003 3432 2007
rect 3436 2006 3437 2007
rect 3450 2007 3456 2008
rect 3450 2006 3451 2007
rect 3436 2004 3451 2006
rect 3436 2003 3437 2004
rect 3431 2002 3437 2003
rect 3450 2003 3451 2004
rect 3455 2003 3456 2007
rect 3450 2002 3456 2003
rect 3534 2007 3541 2008
rect 3534 2003 3535 2007
rect 3540 2003 3541 2007
rect 3534 2002 3541 2003
rect 3166 1998 3172 1999
rect 2948 1992 3074 1994
rect 3078 1995 3084 1996
rect 2948 1991 2949 1992
rect 2943 1990 2949 1991
rect 3078 1991 3079 1995
rect 3083 1994 3084 1995
rect 3143 1995 3149 1996
rect 3143 1994 3144 1995
rect 3083 1992 3144 1994
rect 3083 1991 3084 1992
rect 3078 1990 3084 1991
rect 3143 1991 3144 1992
rect 3148 1991 3149 1995
rect 3143 1990 3149 1991
rect 3170 1995 3176 1996
rect 3170 1991 3171 1995
rect 3175 1994 3176 1995
rect 3351 1995 3357 1996
rect 3351 1994 3352 1995
rect 3175 1992 3352 1994
rect 3175 1991 3176 1992
rect 3170 1990 3176 1991
rect 3351 1991 3352 1992
rect 3356 1991 3357 1995
rect 3351 1990 3357 1991
rect 3535 1995 3541 1996
rect 3535 1991 3536 1995
rect 3540 1994 3541 1995
rect 3562 1995 3568 1996
rect 3562 1994 3563 1995
rect 3540 1992 3563 1994
rect 3540 1991 3541 1992
rect 3535 1990 3541 1991
rect 3562 1991 3563 1992
rect 3567 1991 3568 1995
rect 3562 1990 3568 1991
rect 2227 1987 2228 1990
rect 190 1986 196 1987
rect 190 1982 191 1986
rect 195 1982 196 1986
rect 190 1981 196 1982
rect 350 1986 356 1987
rect 350 1982 351 1986
rect 355 1982 356 1986
rect 350 1981 356 1982
rect 518 1986 524 1987
rect 518 1982 519 1986
rect 523 1982 524 1986
rect 518 1981 524 1982
rect 686 1986 692 1987
rect 686 1982 687 1986
rect 691 1982 692 1986
rect 686 1981 692 1982
rect 854 1986 860 1987
rect 854 1982 855 1986
rect 859 1982 860 1986
rect 854 1981 860 1982
rect 1014 1986 1020 1987
rect 1014 1982 1015 1986
rect 1019 1982 1020 1986
rect 1014 1981 1020 1982
rect 1166 1986 1172 1987
rect 1166 1982 1167 1986
rect 1171 1982 1172 1986
rect 1166 1981 1172 1982
rect 1310 1986 1316 1987
rect 1310 1982 1311 1986
rect 1315 1982 1316 1986
rect 1310 1981 1316 1982
rect 1446 1986 1452 1987
rect 1446 1982 1447 1986
rect 1451 1982 1452 1986
rect 1446 1981 1452 1982
rect 1582 1986 1588 1987
rect 1582 1982 1583 1986
rect 1587 1982 1588 1986
rect 1582 1981 1588 1982
rect 1718 1986 1724 1987
rect 1718 1982 1719 1986
rect 1723 1982 1724 1986
rect 1718 1981 1724 1982
rect 1958 1986 1964 1987
rect 1958 1982 1959 1986
rect 1963 1982 1964 1986
rect 1958 1981 1964 1982
rect 2078 1986 2084 1987
rect 2078 1982 2079 1986
rect 2083 1982 2084 1986
rect 2078 1981 2084 1982
rect 2198 1986 2204 1987
rect 2222 1986 2228 1987
rect 2318 1986 2324 1987
rect 2198 1982 2199 1986
rect 2203 1982 2204 1986
rect 2198 1981 2204 1982
rect 2318 1982 2319 1986
rect 2323 1982 2324 1986
rect 2318 1981 2324 1982
rect 2446 1986 2452 1987
rect 2446 1982 2447 1986
rect 2451 1982 2452 1986
rect 2446 1981 2452 1982
rect 2582 1986 2588 1987
rect 2582 1982 2583 1986
rect 2587 1982 2588 1986
rect 2582 1981 2588 1982
rect 2742 1986 2748 1987
rect 2742 1982 2743 1986
rect 2747 1982 2748 1986
rect 2742 1981 2748 1982
rect 2918 1986 2924 1987
rect 2918 1982 2919 1986
rect 2923 1982 2924 1986
rect 2918 1981 2924 1982
rect 3118 1986 3124 1987
rect 3118 1982 3119 1986
rect 3123 1982 3124 1986
rect 3118 1981 3124 1982
rect 3326 1986 3332 1987
rect 3326 1982 3327 1986
rect 3331 1982 3332 1986
rect 3326 1981 3332 1982
rect 3510 1986 3516 1987
rect 3510 1982 3511 1986
rect 3515 1982 3516 1986
rect 3510 1981 3516 1982
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 1830 1968 1836 1969
rect 1830 1964 1831 1968
rect 1835 1964 1836 1968
rect 1830 1963 1836 1964
rect 1870 1968 1876 1969
rect 1870 1964 1871 1968
rect 1875 1964 1876 1968
rect 1870 1963 1876 1964
rect 3590 1968 3596 1969
rect 3590 1964 3591 1968
rect 3595 1964 3596 1968
rect 3590 1963 3596 1964
rect 358 1959 364 1960
rect 358 1955 359 1959
rect 363 1955 364 1959
rect 358 1954 364 1955
rect 570 1959 576 1960
rect 570 1955 571 1959
rect 575 1955 576 1959
rect 570 1954 576 1955
rect 738 1959 744 1960
rect 738 1955 739 1959
rect 743 1955 744 1959
rect 738 1954 744 1955
rect 862 1959 868 1960
rect 862 1955 863 1959
rect 867 1955 868 1959
rect 862 1954 868 1955
rect 1022 1959 1028 1960
rect 1022 1955 1023 1959
rect 1027 1955 1028 1959
rect 1022 1954 1028 1955
rect 1174 1959 1180 1960
rect 1174 1955 1175 1959
rect 1179 1955 1180 1959
rect 1174 1954 1180 1955
rect 1362 1959 1368 1960
rect 1362 1955 1363 1959
rect 1367 1955 1368 1959
rect 1362 1954 1368 1955
rect 1498 1959 1504 1960
rect 1498 1955 1499 1959
rect 1503 1955 1504 1959
rect 1498 1954 1504 1955
rect 1634 1959 1640 1960
rect 1634 1955 1635 1959
rect 1639 1955 1640 1959
rect 1634 1954 1640 1955
rect 1998 1959 2004 1960
rect 1998 1955 1999 1959
rect 2003 1955 2004 1959
rect 1998 1954 2004 1955
rect 2086 1959 2092 1960
rect 2086 1955 2087 1959
rect 2091 1955 2092 1959
rect 2086 1954 2092 1955
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 2590 1959 2596 1960
rect 2590 1955 2591 1959
rect 2595 1955 2596 1959
rect 2590 1954 2596 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2926 1959 2932 1960
rect 2926 1955 2927 1959
rect 2931 1955 2932 1959
rect 2926 1954 2932 1955
rect 3170 1959 3176 1960
rect 3170 1955 3171 1959
rect 3175 1955 3176 1959
rect 3170 1954 3176 1955
rect 3178 1959 3184 1960
rect 3178 1955 3179 1959
rect 3183 1958 3184 1959
rect 3534 1959 3540 1960
rect 3183 1956 3337 1958
rect 3183 1955 3184 1956
rect 3178 1954 3184 1955
rect 3534 1955 3535 1959
rect 3539 1955 3540 1959
rect 3534 1954 3540 1955
rect 110 1951 116 1952
rect 110 1947 111 1951
rect 115 1947 116 1951
rect 1830 1951 1836 1952
rect 110 1946 116 1947
rect 182 1948 188 1949
rect 182 1944 183 1948
rect 187 1944 188 1948
rect 182 1943 188 1944
rect 342 1948 348 1949
rect 342 1944 343 1948
rect 347 1944 348 1948
rect 342 1943 348 1944
rect 510 1948 516 1949
rect 510 1944 511 1948
rect 515 1944 516 1948
rect 510 1943 516 1944
rect 678 1948 684 1949
rect 678 1944 679 1948
rect 683 1944 684 1948
rect 678 1943 684 1944
rect 846 1948 852 1949
rect 846 1944 847 1948
rect 851 1944 852 1948
rect 846 1943 852 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1158 1948 1164 1949
rect 1158 1944 1159 1948
rect 1163 1944 1164 1948
rect 1158 1943 1164 1944
rect 1302 1948 1308 1949
rect 1302 1944 1303 1948
rect 1307 1944 1308 1948
rect 1302 1943 1308 1944
rect 1438 1948 1444 1949
rect 1438 1944 1439 1948
rect 1443 1944 1444 1948
rect 1438 1943 1444 1944
rect 1574 1948 1580 1949
rect 1574 1944 1575 1948
rect 1579 1944 1580 1948
rect 1574 1943 1580 1944
rect 1710 1948 1716 1949
rect 1710 1944 1711 1948
rect 1715 1944 1716 1948
rect 1830 1947 1831 1951
rect 1835 1947 1836 1951
rect 1830 1946 1836 1947
rect 1870 1951 1876 1952
rect 1870 1947 1871 1951
rect 1875 1947 1876 1951
rect 3590 1951 3596 1952
rect 1870 1946 1876 1947
rect 1950 1948 1956 1949
rect 1710 1943 1716 1944
rect 1950 1944 1951 1948
rect 1955 1944 1956 1948
rect 1950 1943 1956 1944
rect 2070 1948 2076 1949
rect 2070 1944 2071 1948
rect 2075 1944 2076 1948
rect 2070 1943 2076 1944
rect 2190 1948 2196 1949
rect 2190 1944 2191 1948
rect 2195 1944 2196 1948
rect 2190 1943 2196 1944
rect 2310 1948 2316 1949
rect 2310 1944 2311 1948
rect 2315 1944 2316 1948
rect 2310 1943 2316 1944
rect 2438 1948 2444 1949
rect 2438 1944 2439 1948
rect 2443 1944 2444 1948
rect 2438 1943 2444 1944
rect 2574 1948 2580 1949
rect 2574 1944 2575 1948
rect 2579 1944 2580 1948
rect 2574 1943 2580 1944
rect 2734 1948 2740 1949
rect 2734 1944 2735 1948
rect 2739 1944 2740 1948
rect 2734 1943 2740 1944
rect 2910 1948 2916 1949
rect 2910 1944 2911 1948
rect 2915 1944 2916 1948
rect 2910 1943 2916 1944
rect 3110 1948 3116 1949
rect 3110 1944 3111 1948
rect 3115 1944 3116 1948
rect 3110 1943 3116 1944
rect 3318 1948 3324 1949
rect 3318 1944 3319 1948
rect 3323 1944 3324 1948
rect 3318 1943 3324 1944
rect 3502 1948 3508 1949
rect 3502 1944 3503 1948
rect 3507 1944 3508 1948
rect 3590 1947 3591 1951
rect 3595 1947 3596 1951
rect 3590 1946 3596 1947
rect 3502 1943 3508 1944
rect 198 1931 205 1932
rect 198 1927 199 1931
rect 204 1927 205 1931
rect 198 1926 205 1927
rect 1726 1931 1733 1932
rect 1726 1927 1727 1931
rect 1732 1927 1733 1931
rect 1726 1926 1733 1927
rect 2302 1931 2308 1932
rect 2302 1927 2303 1931
rect 2307 1930 2308 1931
rect 2327 1931 2333 1932
rect 2327 1930 2328 1931
rect 2307 1928 2328 1930
rect 2307 1927 2308 1928
rect 2302 1926 2308 1927
rect 2327 1927 2328 1928
rect 2332 1927 2333 1931
rect 2327 1926 2333 1927
rect 2378 1931 2384 1932
rect 2378 1927 2379 1931
rect 2383 1930 2384 1931
rect 2455 1931 2461 1932
rect 2455 1930 2456 1931
rect 2383 1928 2456 1930
rect 2383 1927 2384 1928
rect 2378 1926 2384 1927
rect 2455 1927 2456 1928
rect 2460 1927 2461 1931
rect 2455 1926 2461 1927
rect 134 1900 140 1901
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 134 1896 135 1900
rect 139 1896 140 1900
rect 134 1895 140 1896
rect 238 1900 244 1901
rect 238 1896 239 1900
rect 243 1896 244 1900
rect 238 1895 244 1896
rect 374 1900 380 1901
rect 374 1896 375 1900
rect 379 1896 380 1900
rect 374 1895 380 1896
rect 526 1900 532 1901
rect 526 1896 527 1900
rect 531 1896 532 1900
rect 526 1895 532 1896
rect 686 1900 692 1901
rect 686 1896 687 1900
rect 691 1896 692 1900
rect 686 1895 692 1896
rect 846 1900 852 1901
rect 846 1896 847 1900
rect 851 1896 852 1900
rect 846 1895 852 1896
rect 1006 1900 1012 1901
rect 1006 1896 1007 1900
rect 1011 1896 1012 1900
rect 1006 1895 1012 1896
rect 1158 1900 1164 1901
rect 1158 1896 1159 1900
rect 1163 1896 1164 1900
rect 1158 1895 1164 1896
rect 1302 1900 1308 1901
rect 1302 1896 1303 1900
rect 1307 1896 1308 1900
rect 1302 1895 1308 1896
rect 1454 1900 1460 1901
rect 1454 1896 1455 1900
rect 1459 1896 1460 1900
rect 1454 1895 1460 1896
rect 1606 1900 1612 1901
rect 1606 1896 1607 1900
rect 1611 1896 1612 1900
rect 1606 1895 1612 1896
rect 1830 1897 1836 1898
rect 110 1892 116 1893
rect 1830 1893 1831 1897
rect 1835 1893 1836 1897
rect 2062 1896 2068 1897
rect 1830 1892 1836 1893
rect 1870 1893 1876 1894
rect 210 1891 216 1892
rect 210 1890 211 1891
rect 197 1888 211 1890
rect 210 1887 211 1888
rect 215 1887 216 1891
rect 306 1891 312 1892
rect 306 1890 307 1891
rect 301 1888 307 1890
rect 210 1886 216 1887
rect 306 1887 307 1888
rect 311 1887 312 1891
rect 306 1886 312 1887
rect 354 1891 360 1892
rect 354 1887 355 1891
rect 359 1890 360 1891
rect 594 1891 600 1892
rect 359 1888 393 1890
rect 536 1888 545 1890
rect 359 1887 360 1888
rect 354 1886 360 1887
rect 534 1887 540 1888
rect 534 1883 535 1887
rect 539 1883 540 1887
rect 594 1887 595 1891
rect 599 1890 600 1891
rect 754 1891 760 1892
rect 599 1888 705 1890
rect 599 1887 600 1888
rect 594 1886 600 1887
rect 754 1887 755 1891
rect 759 1890 760 1891
rect 1078 1891 1084 1892
rect 1078 1890 1079 1891
rect 759 1888 865 1890
rect 1069 1888 1079 1890
rect 759 1887 760 1888
rect 754 1886 760 1887
rect 1078 1887 1079 1888
rect 1083 1887 1084 1891
rect 1226 1891 1232 1892
rect 1078 1886 1084 1887
rect 1220 1884 1222 1889
rect 1226 1887 1227 1891
rect 1231 1890 1232 1891
rect 1370 1891 1376 1892
rect 1231 1888 1321 1890
rect 1231 1887 1232 1888
rect 1226 1886 1232 1887
rect 1370 1887 1371 1891
rect 1375 1890 1376 1891
rect 1522 1891 1528 1892
rect 1375 1888 1473 1890
rect 1375 1887 1376 1888
rect 1370 1886 1376 1887
rect 1522 1887 1523 1891
rect 1527 1890 1528 1891
rect 1527 1888 1625 1890
rect 1870 1889 1871 1893
rect 1875 1889 1876 1893
rect 2062 1892 2063 1896
rect 2067 1892 2068 1896
rect 2062 1891 2068 1892
rect 2150 1896 2156 1897
rect 2150 1892 2151 1896
rect 2155 1892 2156 1896
rect 2150 1891 2156 1892
rect 2238 1896 2244 1897
rect 2238 1892 2239 1896
rect 2243 1892 2244 1896
rect 2238 1891 2244 1892
rect 2318 1896 2324 1897
rect 2318 1892 2319 1896
rect 2323 1892 2324 1896
rect 2318 1891 2324 1892
rect 2398 1896 2404 1897
rect 2398 1892 2399 1896
rect 2403 1892 2404 1896
rect 2398 1891 2404 1892
rect 2486 1896 2492 1897
rect 2486 1892 2487 1896
rect 2491 1892 2492 1896
rect 2486 1891 2492 1892
rect 2574 1896 2580 1897
rect 2574 1892 2575 1896
rect 2579 1892 2580 1896
rect 2574 1891 2580 1892
rect 2662 1896 2668 1897
rect 2662 1892 2663 1896
rect 2667 1892 2668 1896
rect 2662 1891 2668 1892
rect 2758 1896 2764 1897
rect 2758 1892 2759 1896
rect 2763 1892 2764 1896
rect 2758 1891 2764 1892
rect 2870 1896 2876 1897
rect 2870 1892 2871 1896
rect 2875 1892 2876 1896
rect 2870 1891 2876 1892
rect 2990 1896 2996 1897
rect 2990 1892 2991 1896
rect 2995 1892 2996 1896
rect 2990 1891 2996 1892
rect 3118 1896 3124 1897
rect 3118 1892 3119 1896
rect 3123 1892 3124 1896
rect 3118 1891 3124 1892
rect 3246 1896 3252 1897
rect 3246 1892 3247 1896
rect 3251 1892 3252 1896
rect 3246 1891 3252 1892
rect 3382 1896 3388 1897
rect 3382 1892 3383 1896
rect 3387 1892 3388 1896
rect 3382 1891 3388 1892
rect 3502 1896 3508 1897
rect 3502 1892 3503 1896
rect 3507 1892 3508 1896
rect 3502 1891 3508 1892
rect 3590 1893 3596 1894
rect 1870 1888 1876 1889
rect 3590 1889 3591 1893
rect 3595 1889 3596 1893
rect 3590 1888 3596 1889
rect 1527 1887 1528 1888
rect 1522 1886 1528 1887
rect 2130 1887 2136 1888
rect 2130 1886 2131 1887
rect 2125 1884 2131 1886
rect 534 1882 540 1883
rect 1218 1883 1224 1884
rect 110 1880 116 1881
rect 110 1876 111 1880
rect 115 1876 116 1880
rect 1218 1879 1219 1883
rect 1223 1879 1224 1883
rect 2130 1883 2131 1884
rect 2135 1883 2136 1887
rect 2222 1887 2228 1888
rect 2222 1886 2223 1887
rect 2213 1884 2223 1886
rect 2130 1882 2136 1883
rect 2222 1883 2223 1884
rect 2227 1883 2228 1887
rect 2386 1887 2392 1888
rect 2386 1886 2387 1887
rect 2222 1882 2228 1883
rect 1218 1878 1224 1879
rect 1830 1880 1836 1881
rect 110 1875 116 1876
rect 1830 1876 1831 1880
rect 1835 1876 1836 1880
rect 2300 1878 2302 1885
rect 2381 1884 2387 1886
rect 2386 1883 2387 1884
rect 2391 1883 2392 1887
rect 2466 1887 2472 1888
rect 2466 1886 2467 1887
rect 2461 1884 2467 1886
rect 2386 1882 2392 1883
rect 2466 1883 2467 1884
rect 2471 1883 2472 1887
rect 2554 1887 2560 1888
rect 2554 1886 2555 1887
rect 2549 1884 2555 1886
rect 2466 1882 2472 1883
rect 2554 1883 2555 1884
rect 2559 1883 2560 1887
rect 2642 1887 2648 1888
rect 2642 1886 2643 1887
rect 2637 1884 2643 1886
rect 2554 1882 2560 1883
rect 2642 1883 2643 1884
rect 2647 1883 2648 1887
rect 2734 1887 2740 1888
rect 2734 1886 2735 1887
rect 2725 1884 2735 1886
rect 2642 1882 2648 1883
rect 2734 1883 2735 1884
rect 2739 1883 2740 1887
rect 2863 1887 2869 1888
rect 2863 1886 2864 1887
rect 2821 1884 2864 1886
rect 2734 1882 2740 1883
rect 2863 1883 2864 1884
rect 2868 1883 2869 1887
rect 2954 1887 2960 1888
rect 2954 1886 2955 1887
rect 2933 1884 2955 1886
rect 2863 1882 2869 1883
rect 2954 1883 2955 1884
rect 2959 1883 2960 1887
rect 3078 1887 3084 1888
rect 3078 1886 3079 1887
rect 3053 1884 3079 1886
rect 2954 1882 2960 1883
rect 3078 1883 3079 1884
rect 3083 1883 3084 1887
rect 3194 1887 3200 1888
rect 3194 1886 3195 1887
rect 3181 1884 3195 1886
rect 3078 1882 3084 1883
rect 3194 1883 3195 1884
rect 3199 1883 3200 1887
rect 3194 1882 3200 1883
rect 3202 1887 3208 1888
rect 3202 1883 3203 1887
rect 3207 1886 3208 1887
rect 3450 1887 3456 1888
rect 3450 1886 3451 1887
rect 3207 1884 3265 1886
rect 3445 1884 3451 1886
rect 3207 1883 3208 1884
rect 3202 1882 3208 1883
rect 3450 1883 3451 1884
rect 3455 1883 3456 1887
rect 3450 1882 3456 1883
rect 3458 1887 3464 1888
rect 3458 1883 3459 1887
rect 3463 1886 3464 1887
rect 3463 1884 3521 1886
rect 3463 1883 3464 1884
rect 3458 1882 3464 1883
rect 2458 1879 2464 1880
rect 2458 1878 2459 1879
rect 1830 1875 1836 1876
rect 1870 1876 1876 1877
rect 2300 1876 2459 1878
rect 1870 1872 1871 1876
rect 1875 1872 1876 1876
rect 2458 1875 2459 1876
rect 2463 1875 2464 1879
rect 2458 1874 2464 1875
rect 3590 1876 3596 1877
rect 1870 1871 1876 1872
rect 3590 1872 3591 1876
rect 3595 1872 3596 1876
rect 3590 1871 3596 1872
rect 142 1862 148 1863
rect 142 1858 143 1862
rect 147 1858 148 1862
rect 142 1857 148 1858
rect 246 1862 252 1863
rect 246 1858 247 1862
rect 251 1858 252 1862
rect 246 1857 252 1858
rect 382 1862 388 1863
rect 382 1858 383 1862
rect 387 1858 388 1862
rect 382 1857 388 1858
rect 534 1862 540 1863
rect 534 1858 535 1862
rect 539 1858 540 1862
rect 534 1857 540 1858
rect 694 1862 700 1863
rect 694 1858 695 1862
rect 699 1858 700 1862
rect 694 1857 700 1858
rect 854 1862 860 1863
rect 854 1858 855 1862
rect 859 1858 860 1862
rect 854 1857 860 1858
rect 1014 1862 1020 1863
rect 1014 1858 1015 1862
rect 1019 1858 1020 1862
rect 1014 1857 1020 1858
rect 1166 1862 1172 1863
rect 1166 1858 1167 1862
rect 1171 1858 1172 1862
rect 1166 1857 1172 1858
rect 1310 1862 1316 1863
rect 1310 1858 1311 1862
rect 1315 1858 1316 1862
rect 1310 1857 1316 1858
rect 1462 1862 1468 1863
rect 1462 1858 1463 1862
rect 1467 1858 1468 1862
rect 1462 1857 1468 1858
rect 1614 1862 1620 1863
rect 1614 1858 1615 1862
rect 1619 1858 1620 1862
rect 1614 1857 1620 1858
rect 2070 1858 2076 1859
rect 2070 1854 2071 1858
rect 2075 1854 2076 1858
rect 2070 1853 2076 1854
rect 2158 1858 2164 1859
rect 2158 1854 2159 1858
rect 2163 1854 2164 1858
rect 2158 1853 2164 1854
rect 2246 1858 2252 1859
rect 2246 1854 2247 1858
rect 2251 1854 2252 1858
rect 2246 1853 2252 1854
rect 2326 1858 2332 1859
rect 2326 1854 2327 1858
rect 2331 1854 2332 1858
rect 2326 1853 2332 1854
rect 2406 1858 2412 1859
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2494 1858 2500 1859
rect 2494 1854 2495 1858
rect 2499 1854 2500 1858
rect 2494 1853 2500 1854
rect 2582 1858 2588 1859
rect 2582 1854 2583 1858
rect 2587 1854 2588 1858
rect 2582 1853 2588 1854
rect 2670 1858 2676 1859
rect 2670 1854 2671 1858
rect 2675 1854 2676 1858
rect 2670 1853 2676 1854
rect 2766 1858 2772 1859
rect 2766 1854 2767 1858
rect 2771 1854 2772 1858
rect 2766 1853 2772 1854
rect 2878 1858 2884 1859
rect 2878 1854 2879 1858
rect 2883 1854 2884 1858
rect 2878 1853 2884 1854
rect 2998 1858 3004 1859
rect 2998 1854 2999 1858
rect 3003 1854 3004 1858
rect 2998 1853 3004 1854
rect 3126 1858 3132 1859
rect 3126 1854 3127 1858
rect 3131 1854 3132 1858
rect 3126 1853 3132 1854
rect 3254 1858 3260 1859
rect 3254 1854 3255 1858
rect 3259 1854 3260 1858
rect 3254 1853 3260 1854
rect 3390 1858 3396 1859
rect 3390 1854 3391 1858
rect 3395 1854 3396 1858
rect 3390 1853 3396 1854
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 167 1851 173 1852
rect 167 1847 168 1851
rect 172 1850 173 1851
rect 198 1851 204 1852
rect 198 1850 199 1851
rect 172 1848 199 1850
rect 172 1847 173 1848
rect 167 1846 173 1847
rect 198 1847 199 1848
rect 203 1847 204 1851
rect 198 1846 204 1847
rect 210 1851 216 1852
rect 210 1847 211 1851
rect 215 1850 216 1851
rect 271 1851 277 1852
rect 271 1850 272 1851
rect 215 1848 272 1850
rect 215 1847 216 1848
rect 210 1846 216 1847
rect 271 1847 272 1848
rect 276 1847 277 1851
rect 271 1846 277 1847
rect 306 1851 312 1852
rect 306 1847 307 1851
rect 311 1850 312 1851
rect 407 1851 413 1852
rect 407 1850 408 1851
rect 311 1848 408 1850
rect 311 1847 312 1848
rect 306 1846 312 1847
rect 407 1847 408 1848
rect 412 1847 413 1851
rect 407 1846 413 1847
rect 559 1851 565 1852
rect 559 1847 560 1851
rect 564 1850 565 1851
rect 594 1851 600 1852
rect 594 1850 595 1851
rect 564 1848 595 1850
rect 564 1847 565 1848
rect 559 1846 565 1847
rect 594 1847 595 1848
rect 599 1847 600 1851
rect 594 1846 600 1847
rect 719 1851 725 1852
rect 719 1847 720 1851
rect 724 1850 725 1851
rect 754 1851 760 1852
rect 754 1850 755 1851
rect 724 1848 755 1850
rect 724 1847 725 1848
rect 719 1846 725 1847
rect 754 1847 755 1848
rect 759 1847 760 1851
rect 754 1846 760 1847
rect 878 1851 885 1852
rect 878 1847 879 1851
rect 884 1847 885 1851
rect 878 1846 885 1847
rect 1038 1851 1045 1852
rect 1038 1847 1039 1851
rect 1044 1847 1045 1851
rect 1038 1846 1045 1847
rect 1078 1851 1084 1852
rect 1078 1847 1079 1851
rect 1083 1850 1084 1851
rect 1191 1851 1197 1852
rect 1191 1850 1192 1851
rect 1083 1848 1192 1850
rect 1083 1847 1084 1848
rect 1078 1846 1084 1847
rect 1191 1847 1192 1848
rect 1196 1847 1197 1851
rect 1191 1846 1197 1847
rect 1335 1851 1341 1852
rect 1335 1847 1336 1851
rect 1340 1850 1341 1851
rect 1370 1851 1376 1852
rect 1370 1850 1371 1851
rect 1340 1848 1371 1850
rect 1340 1847 1341 1848
rect 1335 1846 1341 1847
rect 1370 1847 1371 1848
rect 1375 1847 1376 1851
rect 1370 1846 1376 1847
rect 1487 1851 1493 1852
rect 1487 1847 1488 1851
rect 1492 1850 1493 1851
rect 1522 1851 1528 1852
rect 1522 1850 1523 1851
rect 1492 1848 1523 1850
rect 1492 1847 1493 1848
rect 1487 1846 1493 1847
rect 1522 1847 1523 1848
rect 1527 1847 1528 1851
rect 1522 1846 1528 1847
rect 1639 1851 1645 1852
rect 1639 1847 1640 1851
rect 1644 1850 1645 1851
rect 1726 1851 1732 1852
rect 1726 1850 1727 1851
rect 1644 1848 1727 1850
rect 1644 1847 1645 1848
rect 1639 1846 1645 1847
rect 1726 1847 1727 1848
rect 1731 1847 1732 1851
rect 1726 1846 1732 1847
rect 2094 1847 2101 1848
rect 2094 1843 2095 1847
rect 2100 1843 2101 1847
rect 2094 1842 2101 1843
rect 2130 1847 2136 1848
rect 2130 1843 2131 1847
rect 2135 1846 2136 1847
rect 2183 1847 2189 1848
rect 2183 1846 2184 1847
rect 2135 1844 2184 1846
rect 2135 1843 2136 1844
rect 2130 1842 2136 1843
rect 2183 1843 2184 1844
rect 2188 1843 2189 1847
rect 2183 1842 2189 1843
rect 2271 1847 2277 1848
rect 2271 1843 2272 1847
rect 2276 1846 2277 1847
rect 2302 1847 2308 1848
rect 2302 1846 2303 1847
rect 2276 1844 2303 1846
rect 2276 1843 2277 1844
rect 2271 1842 2277 1843
rect 2302 1843 2303 1844
rect 2307 1843 2308 1847
rect 2302 1842 2308 1843
rect 2351 1847 2357 1848
rect 2351 1843 2352 1847
rect 2356 1846 2357 1847
rect 2378 1847 2384 1848
rect 2378 1846 2379 1847
rect 2356 1844 2379 1846
rect 2356 1843 2357 1844
rect 2351 1842 2357 1843
rect 2378 1843 2379 1844
rect 2383 1843 2384 1847
rect 2378 1842 2384 1843
rect 2386 1847 2392 1848
rect 2386 1843 2387 1847
rect 2391 1846 2392 1847
rect 2431 1847 2437 1848
rect 2431 1846 2432 1847
rect 2391 1844 2432 1846
rect 2391 1843 2392 1844
rect 2386 1842 2392 1843
rect 2431 1843 2432 1844
rect 2436 1843 2437 1847
rect 2431 1842 2437 1843
rect 2466 1847 2472 1848
rect 2466 1843 2467 1847
rect 2471 1846 2472 1847
rect 2519 1847 2525 1848
rect 2519 1846 2520 1847
rect 2471 1844 2520 1846
rect 2471 1843 2472 1844
rect 2466 1842 2472 1843
rect 2519 1843 2520 1844
rect 2524 1843 2525 1847
rect 2519 1842 2525 1843
rect 2554 1847 2560 1848
rect 2554 1843 2555 1847
rect 2559 1846 2560 1847
rect 2607 1847 2613 1848
rect 2607 1846 2608 1847
rect 2559 1844 2608 1846
rect 2559 1843 2560 1844
rect 2554 1842 2560 1843
rect 2607 1843 2608 1844
rect 2612 1843 2613 1847
rect 2607 1842 2613 1843
rect 2642 1847 2648 1848
rect 2642 1843 2643 1847
rect 2647 1846 2648 1847
rect 2695 1847 2701 1848
rect 2695 1846 2696 1847
rect 2647 1844 2696 1846
rect 2647 1843 2648 1844
rect 2642 1842 2648 1843
rect 2695 1843 2696 1844
rect 2700 1843 2701 1847
rect 2695 1842 2701 1843
rect 2734 1847 2740 1848
rect 2734 1843 2735 1847
rect 2739 1846 2740 1847
rect 2791 1847 2797 1848
rect 2791 1846 2792 1847
rect 2739 1844 2792 1846
rect 2739 1843 2740 1844
rect 2734 1842 2740 1843
rect 2791 1843 2792 1844
rect 2796 1843 2797 1847
rect 2791 1842 2797 1843
rect 2863 1847 2869 1848
rect 2863 1843 2864 1847
rect 2868 1846 2869 1847
rect 2903 1847 2909 1848
rect 2903 1846 2904 1847
rect 2868 1844 2904 1846
rect 2868 1843 2869 1844
rect 2863 1842 2869 1843
rect 2903 1843 2904 1844
rect 2908 1843 2909 1847
rect 2903 1842 2909 1843
rect 2954 1847 2960 1848
rect 2954 1843 2955 1847
rect 2959 1846 2960 1847
rect 3023 1847 3029 1848
rect 3023 1846 3024 1847
rect 2959 1844 3024 1846
rect 2959 1843 2960 1844
rect 2954 1842 2960 1843
rect 3023 1843 3024 1844
rect 3028 1843 3029 1847
rect 3023 1842 3029 1843
rect 3078 1847 3084 1848
rect 3078 1843 3079 1847
rect 3083 1846 3084 1847
rect 3151 1847 3157 1848
rect 3151 1846 3152 1847
rect 3083 1844 3152 1846
rect 3083 1843 3084 1844
rect 3078 1842 3084 1843
rect 3151 1843 3152 1844
rect 3156 1843 3157 1847
rect 3151 1842 3157 1843
rect 3194 1847 3200 1848
rect 3194 1843 3195 1847
rect 3199 1846 3200 1847
rect 3279 1847 3285 1848
rect 3279 1846 3280 1847
rect 3199 1844 3280 1846
rect 3199 1843 3200 1844
rect 3194 1842 3200 1843
rect 3279 1843 3280 1844
rect 3284 1843 3285 1847
rect 3279 1842 3285 1843
rect 3415 1847 3421 1848
rect 3415 1843 3416 1847
rect 3420 1846 3421 1847
rect 3458 1847 3464 1848
rect 3458 1846 3459 1847
rect 3420 1844 3459 1846
rect 3420 1843 3421 1844
rect 3415 1842 3421 1843
rect 3458 1843 3459 1844
rect 3463 1843 3464 1847
rect 3458 1842 3464 1843
rect 3534 1847 3541 1848
rect 3534 1843 3535 1847
rect 3540 1843 3541 1847
rect 3534 1842 3541 1843
rect 167 1835 173 1836
rect 167 1831 168 1835
rect 172 1834 173 1835
rect 294 1835 300 1836
rect 294 1834 295 1835
rect 172 1832 295 1834
rect 172 1831 173 1832
rect 167 1830 173 1831
rect 294 1831 295 1832
rect 299 1831 300 1835
rect 294 1830 300 1831
rect 311 1835 317 1836
rect 311 1831 312 1835
rect 316 1834 317 1835
rect 354 1835 360 1836
rect 354 1834 355 1835
rect 316 1832 355 1834
rect 316 1831 317 1832
rect 311 1830 317 1831
rect 354 1831 355 1832
rect 359 1831 360 1835
rect 354 1830 360 1831
rect 486 1835 492 1836
rect 486 1831 487 1835
rect 491 1834 492 1835
rect 495 1835 501 1836
rect 495 1834 496 1835
rect 491 1832 496 1834
rect 491 1831 492 1832
rect 486 1830 492 1831
rect 495 1831 496 1832
rect 500 1831 501 1835
rect 495 1830 501 1831
rect 522 1835 528 1836
rect 522 1831 523 1835
rect 527 1834 528 1835
rect 687 1835 693 1836
rect 687 1834 688 1835
rect 527 1832 688 1834
rect 527 1831 528 1832
rect 522 1830 528 1831
rect 687 1831 688 1832
rect 692 1831 693 1835
rect 687 1830 693 1831
rect 714 1835 720 1836
rect 714 1831 715 1835
rect 719 1834 720 1835
rect 871 1835 877 1836
rect 871 1834 872 1835
rect 719 1832 872 1834
rect 719 1831 720 1832
rect 714 1830 720 1831
rect 871 1831 872 1832
rect 876 1831 877 1835
rect 871 1830 877 1831
rect 1047 1835 1053 1836
rect 1047 1831 1048 1835
rect 1052 1834 1053 1835
rect 1102 1835 1108 1836
rect 1102 1834 1103 1835
rect 1052 1832 1103 1834
rect 1052 1831 1053 1832
rect 1047 1830 1053 1831
rect 1102 1831 1103 1832
rect 1107 1831 1108 1835
rect 1102 1830 1108 1831
rect 1215 1835 1221 1836
rect 1215 1831 1216 1835
rect 1220 1834 1221 1835
rect 1226 1835 1232 1836
rect 1226 1834 1227 1835
rect 1220 1832 1227 1834
rect 1220 1831 1221 1832
rect 1215 1830 1221 1831
rect 1226 1831 1227 1832
rect 1231 1831 1232 1835
rect 1226 1830 1232 1831
rect 1242 1835 1248 1836
rect 1242 1831 1243 1835
rect 1247 1834 1248 1835
rect 1375 1835 1381 1836
rect 1375 1834 1376 1835
rect 1247 1832 1376 1834
rect 1247 1831 1248 1832
rect 1242 1830 1248 1831
rect 1375 1831 1376 1832
rect 1380 1831 1381 1835
rect 1375 1830 1381 1831
rect 1402 1835 1408 1836
rect 1402 1831 1403 1835
rect 1407 1834 1408 1835
rect 1535 1835 1541 1836
rect 1535 1834 1536 1835
rect 1407 1832 1536 1834
rect 1407 1831 1408 1832
rect 1402 1830 1408 1831
rect 1535 1831 1536 1832
rect 1540 1831 1541 1835
rect 1535 1830 1541 1831
rect 1562 1835 1568 1836
rect 1562 1831 1563 1835
rect 1567 1834 1568 1835
rect 1703 1835 1709 1836
rect 1703 1834 1704 1835
rect 1567 1832 1704 1834
rect 1567 1831 1568 1832
rect 1562 1830 1568 1831
rect 1703 1831 1704 1832
rect 1708 1831 1709 1835
rect 1703 1830 1709 1831
rect 142 1826 148 1827
rect 142 1822 143 1826
rect 147 1822 148 1826
rect 142 1821 148 1822
rect 286 1826 292 1827
rect 286 1822 287 1826
rect 291 1822 292 1826
rect 286 1821 292 1822
rect 470 1826 476 1827
rect 470 1822 471 1826
rect 475 1822 476 1826
rect 470 1821 476 1822
rect 662 1826 668 1827
rect 662 1822 663 1826
rect 667 1822 668 1826
rect 662 1821 668 1822
rect 846 1826 852 1827
rect 846 1822 847 1826
rect 851 1822 852 1826
rect 846 1821 852 1822
rect 1022 1826 1028 1827
rect 1022 1822 1023 1826
rect 1027 1822 1028 1826
rect 1022 1821 1028 1822
rect 1190 1826 1196 1827
rect 1190 1822 1191 1826
rect 1195 1822 1196 1826
rect 1190 1821 1196 1822
rect 1350 1826 1356 1827
rect 1350 1822 1351 1826
rect 1355 1822 1356 1826
rect 1350 1821 1356 1822
rect 1510 1826 1516 1827
rect 1510 1822 1511 1826
rect 1515 1822 1516 1826
rect 1510 1821 1516 1822
rect 1678 1826 1684 1827
rect 1678 1822 1679 1826
rect 1683 1822 1684 1826
rect 1678 1821 1684 1822
rect 2119 1819 2125 1820
rect 2119 1815 2120 1819
rect 2124 1818 2125 1819
rect 2167 1819 2173 1820
rect 2167 1818 2168 1819
rect 2124 1816 2168 1818
rect 2124 1815 2125 1816
rect 2119 1814 2125 1815
rect 2167 1815 2168 1816
rect 2172 1815 2173 1819
rect 2167 1814 2173 1815
rect 2263 1819 2269 1820
rect 2263 1815 2264 1819
rect 2268 1818 2269 1819
rect 2334 1819 2340 1820
rect 2334 1818 2335 1819
rect 2268 1816 2335 1818
rect 2268 1815 2269 1816
rect 2263 1814 2269 1815
rect 2334 1815 2335 1816
rect 2339 1815 2340 1819
rect 2334 1814 2340 1815
rect 2423 1819 2429 1820
rect 2423 1815 2424 1819
rect 2428 1818 2429 1819
rect 2450 1819 2456 1820
rect 2450 1818 2451 1819
rect 2428 1816 2451 1818
rect 2428 1815 2429 1816
rect 2423 1814 2429 1815
rect 2450 1815 2451 1816
rect 2455 1815 2456 1819
rect 2450 1814 2456 1815
rect 2458 1819 2464 1820
rect 2458 1815 2459 1819
rect 2463 1818 2464 1819
rect 2583 1819 2589 1820
rect 2583 1818 2584 1819
rect 2463 1816 2584 1818
rect 2463 1815 2464 1816
rect 2458 1814 2464 1815
rect 2583 1815 2584 1816
rect 2588 1815 2589 1819
rect 2583 1814 2589 1815
rect 2610 1819 2616 1820
rect 2610 1815 2611 1819
rect 2615 1818 2616 1819
rect 2743 1819 2749 1820
rect 2743 1818 2744 1819
rect 2615 1816 2744 1818
rect 2615 1815 2616 1816
rect 2610 1814 2616 1815
rect 2743 1815 2744 1816
rect 2748 1815 2749 1819
rect 2743 1814 2749 1815
rect 2903 1819 2909 1820
rect 2903 1815 2904 1819
rect 2908 1818 2909 1819
rect 3038 1819 3044 1820
rect 3038 1818 3039 1819
rect 2908 1816 3039 1818
rect 2908 1815 2909 1816
rect 2903 1814 2909 1815
rect 3038 1815 3039 1816
rect 3043 1815 3044 1819
rect 3038 1814 3044 1815
rect 3055 1819 3061 1820
rect 3055 1815 3056 1819
rect 3060 1818 3061 1819
rect 3118 1819 3124 1820
rect 3118 1818 3119 1819
rect 3060 1816 3119 1818
rect 3060 1815 3061 1816
rect 3055 1814 3061 1815
rect 3118 1815 3119 1816
rect 3123 1815 3124 1819
rect 3118 1814 3124 1815
rect 3199 1819 3208 1820
rect 3199 1815 3200 1819
rect 3207 1815 3208 1819
rect 3199 1814 3208 1815
rect 3226 1819 3232 1820
rect 3226 1815 3227 1819
rect 3231 1818 3232 1819
rect 3343 1819 3349 1820
rect 3343 1818 3344 1819
rect 3231 1816 3344 1818
rect 3231 1815 3232 1816
rect 3226 1814 3232 1815
rect 3343 1815 3344 1816
rect 3348 1815 3349 1819
rect 3343 1814 3349 1815
rect 3370 1819 3376 1820
rect 3370 1815 3371 1819
rect 3375 1818 3376 1819
rect 3495 1819 3501 1820
rect 3495 1818 3496 1819
rect 3375 1816 3496 1818
rect 3375 1815 3376 1816
rect 3370 1814 3376 1815
rect 3495 1815 3496 1816
rect 3500 1815 3501 1819
rect 3495 1814 3501 1815
rect 2094 1810 2100 1811
rect 110 1808 116 1809
rect 110 1804 111 1808
rect 115 1804 116 1808
rect 110 1803 116 1804
rect 1830 1808 1836 1809
rect 1830 1804 1831 1808
rect 1835 1804 1836 1808
rect 2094 1806 2095 1810
rect 2099 1806 2100 1810
rect 2094 1805 2100 1806
rect 2238 1810 2244 1811
rect 2238 1806 2239 1810
rect 2243 1806 2244 1810
rect 2238 1805 2244 1806
rect 2398 1810 2404 1811
rect 2398 1806 2399 1810
rect 2403 1806 2404 1810
rect 2398 1805 2404 1806
rect 2558 1810 2564 1811
rect 2558 1806 2559 1810
rect 2563 1806 2564 1810
rect 2558 1805 2564 1806
rect 2718 1810 2724 1811
rect 2718 1806 2719 1810
rect 2723 1806 2724 1810
rect 2718 1805 2724 1806
rect 2878 1810 2884 1811
rect 2878 1806 2879 1810
rect 2883 1806 2884 1810
rect 2878 1805 2884 1806
rect 3030 1810 3036 1811
rect 3030 1806 3031 1810
rect 3035 1806 3036 1810
rect 3030 1805 3036 1806
rect 3174 1810 3180 1811
rect 3174 1806 3175 1810
rect 3179 1806 3180 1810
rect 3174 1805 3180 1806
rect 3318 1810 3324 1811
rect 3318 1806 3319 1810
rect 3323 1806 3324 1810
rect 3318 1805 3324 1806
rect 3470 1810 3476 1811
rect 3470 1806 3471 1810
rect 3475 1806 3476 1810
rect 3470 1805 3476 1806
rect 1830 1803 1836 1804
rect 166 1799 172 1800
rect 166 1795 167 1799
rect 171 1795 172 1799
rect 166 1794 172 1795
rect 294 1799 300 1800
rect 294 1795 295 1799
rect 299 1795 300 1799
rect 294 1794 300 1795
rect 522 1799 528 1800
rect 522 1795 523 1799
rect 527 1795 528 1799
rect 522 1794 528 1795
rect 714 1799 720 1800
rect 714 1795 715 1799
rect 719 1795 720 1799
rect 714 1794 720 1795
rect 878 1799 884 1800
rect 878 1795 879 1799
rect 883 1795 884 1799
rect 878 1794 884 1795
rect 1038 1799 1044 1800
rect 1038 1795 1039 1799
rect 1043 1795 1044 1799
rect 1038 1794 1044 1795
rect 1242 1799 1248 1800
rect 1242 1795 1243 1799
rect 1247 1795 1248 1799
rect 1242 1794 1248 1795
rect 1402 1799 1408 1800
rect 1402 1795 1403 1799
rect 1407 1795 1408 1799
rect 1402 1794 1408 1795
rect 1562 1799 1568 1800
rect 1562 1795 1563 1799
rect 1567 1795 1568 1799
rect 1562 1794 1568 1795
rect 1870 1792 1876 1793
rect 110 1791 116 1792
rect 110 1787 111 1791
rect 115 1787 116 1791
rect 1830 1791 1836 1792
rect 110 1786 116 1787
rect 134 1788 140 1789
rect 134 1784 135 1788
rect 139 1784 140 1788
rect 134 1783 140 1784
rect 278 1788 284 1789
rect 278 1784 279 1788
rect 283 1784 284 1788
rect 278 1783 284 1784
rect 462 1788 468 1789
rect 462 1784 463 1788
rect 467 1784 468 1788
rect 462 1783 468 1784
rect 654 1788 660 1789
rect 654 1784 655 1788
rect 659 1784 660 1788
rect 654 1783 660 1784
rect 838 1788 844 1789
rect 838 1784 839 1788
rect 843 1784 844 1788
rect 838 1783 844 1784
rect 1014 1788 1020 1789
rect 1014 1784 1015 1788
rect 1019 1784 1020 1788
rect 1014 1783 1020 1784
rect 1182 1788 1188 1789
rect 1182 1784 1183 1788
rect 1187 1784 1188 1788
rect 1182 1783 1188 1784
rect 1342 1788 1348 1789
rect 1342 1784 1343 1788
rect 1347 1784 1348 1788
rect 1342 1783 1348 1784
rect 1502 1788 1508 1789
rect 1502 1784 1503 1788
rect 1507 1784 1508 1788
rect 1502 1783 1508 1784
rect 1670 1788 1676 1789
rect 1670 1784 1671 1788
rect 1675 1784 1676 1788
rect 1830 1787 1831 1791
rect 1835 1787 1836 1791
rect 1870 1788 1871 1792
rect 1875 1788 1876 1792
rect 1870 1787 1876 1788
rect 3590 1792 3596 1793
rect 3590 1788 3591 1792
rect 3595 1788 3596 1792
rect 3590 1787 3596 1788
rect 1830 1786 1836 1787
rect 1670 1783 1676 1784
rect 2102 1783 2108 1784
rect 2102 1779 2103 1783
rect 2107 1779 2108 1783
rect 2102 1778 2108 1779
rect 2167 1783 2173 1784
rect 2167 1779 2168 1783
rect 2172 1782 2173 1783
rect 2334 1783 2340 1784
rect 2172 1780 2249 1782
rect 2172 1779 2173 1780
rect 2167 1778 2173 1779
rect 2334 1779 2335 1783
rect 2339 1782 2340 1783
rect 2610 1783 2616 1784
rect 2339 1780 2409 1782
rect 2339 1779 2340 1780
rect 2334 1778 2340 1779
rect 2610 1779 2611 1783
rect 2615 1779 2616 1783
rect 2610 1778 2616 1779
rect 3038 1783 3044 1784
rect 3038 1779 3039 1783
rect 3043 1779 3044 1783
rect 3038 1778 3044 1779
rect 3226 1783 3232 1784
rect 3226 1779 3227 1783
rect 3231 1779 3232 1783
rect 3226 1778 3232 1779
rect 3370 1783 3376 1784
rect 3370 1779 3371 1783
rect 3375 1779 3376 1783
rect 3370 1778 3376 1779
rect 1870 1775 1876 1776
rect 1354 1771 1360 1772
rect 1354 1767 1355 1771
rect 1359 1770 1360 1771
rect 1687 1771 1693 1772
rect 1687 1770 1688 1771
rect 1359 1768 1688 1770
rect 1359 1767 1360 1768
rect 1354 1766 1360 1767
rect 1687 1767 1688 1768
rect 1692 1767 1693 1771
rect 1870 1771 1871 1775
rect 1875 1771 1876 1775
rect 3590 1775 3596 1776
rect 1870 1770 1876 1771
rect 2086 1772 2092 1773
rect 2086 1768 2087 1772
rect 2091 1768 2092 1772
rect 2086 1767 2092 1768
rect 2230 1772 2236 1773
rect 2230 1768 2231 1772
rect 2235 1768 2236 1772
rect 2230 1767 2236 1768
rect 2390 1772 2396 1773
rect 2390 1768 2391 1772
rect 2395 1768 2396 1772
rect 2390 1767 2396 1768
rect 2550 1772 2556 1773
rect 2550 1768 2551 1772
rect 2555 1768 2556 1772
rect 2550 1767 2556 1768
rect 2710 1772 2716 1773
rect 2710 1768 2711 1772
rect 2715 1768 2716 1772
rect 2710 1767 2716 1768
rect 2870 1772 2876 1773
rect 2870 1768 2871 1772
rect 2875 1768 2876 1772
rect 2870 1767 2876 1768
rect 3022 1772 3028 1773
rect 3022 1768 3023 1772
rect 3027 1768 3028 1772
rect 3022 1767 3028 1768
rect 3166 1772 3172 1773
rect 3166 1768 3167 1772
rect 3171 1768 3172 1772
rect 3166 1767 3172 1768
rect 3310 1772 3316 1773
rect 3310 1768 3311 1772
rect 3315 1768 3316 1772
rect 3310 1767 3316 1768
rect 3462 1772 3468 1773
rect 3462 1768 3463 1772
rect 3467 1768 3468 1772
rect 3590 1771 3591 1775
rect 3595 1771 3596 1775
rect 3590 1770 3596 1771
rect 3462 1767 3468 1768
rect 1687 1766 1693 1767
rect 2698 1755 2704 1756
rect 2698 1751 2699 1755
rect 2703 1754 2704 1755
rect 2727 1755 2733 1756
rect 2727 1754 2728 1755
rect 2703 1752 2728 1754
rect 2703 1751 2704 1752
rect 2698 1750 2704 1751
rect 2727 1751 2728 1752
rect 2732 1751 2733 1755
rect 2727 1750 2733 1751
rect 2834 1755 2840 1756
rect 2834 1751 2835 1755
rect 2839 1754 2840 1755
rect 2887 1755 2893 1756
rect 2887 1754 2888 1755
rect 2839 1752 2888 1754
rect 2839 1751 2840 1752
rect 2834 1750 2840 1751
rect 2887 1751 2888 1752
rect 2892 1751 2893 1755
rect 2887 1750 2893 1751
rect 3426 1755 3432 1756
rect 3426 1751 3427 1755
rect 3431 1754 3432 1755
rect 3479 1755 3485 1756
rect 3479 1754 3480 1755
rect 3431 1752 3480 1754
rect 3431 1751 3432 1752
rect 3426 1750 3432 1751
rect 3479 1751 3480 1752
rect 3484 1751 3485 1755
rect 3479 1750 3485 1751
rect 134 1736 140 1737
rect 110 1733 116 1734
rect 110 1729 111 1733
rect 115 1729 116 1733
rect 134 1732 135 1736
rect 139 1732 140 1736
rect 134 1731 140 1732
rect 214 1736 220 1737
rect 214 1732 215 1736
rect 219 1732 220 1736
rect 214 1731 220 1732
rect 342 1736 348 1737
rect 342 1732 343 1736
rect 347 1732 348 1736
rect 342 1731 348 1732
rect 494 1736 500 1737
rect 494 1732 495 1736
rect 499 1732 500 1736
rect 494 1731 500 1732
rect 662 1736 668 1737
rect 662 1732 663 1736
rect 667 1732 668 1736
rect 662 1731 668 1732
rect 838 1736 844 1737
rect 838 1732 839 1736
rect 843 1732 844 1736
rect 838 1731 844 1732
rect 1006 1736 1012 1737
rect 1006 1732 1007 1736
rect 1011 1732 1012 1736
rect 1006 1731 1012 1732
rect 1166 1736 1172 1737
rect 1166 1732 1167 1736
rect 1171 1732 1172 1736
rect 1166 1731 1172 1732
rect 1318 1736 1324 1737
rect 1318 1732 1319 1736
rect 1323 1732 1324 1736
rect 1318 1731 1324 1732
rect 1462 1736 1468 1737
rect 1462 1732 1463 1736
rect 1467 1732 1468 1736
rect 1462 1731 1468 1732
rect 1606 1736 1612 1737
rect 1606 1732 1607 1736
rect 1611 1732 1612 1736
rect 1606 1731 1612 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 1742 1731 1748 1732
rect 1830 1733 1836 1734
rect 110 1728 116 1729
rect 1830 1729 1831 1733
rect 1835 1729 1836 1733
rect 1830 1728 1836 1729
rect 202 1727 208 1728
rect 202 1726 203 1727
rect 197 1724 203 1726
rect 202 1723 203 1724
rect 207 1723 208 1727
rect 282 1727 288 1728
rect 282 1726 283 1727
rect 277 1724 283 1726
rect 202 1722 208 1723
rect 282 1723 283 1724
rect 287 1723 288 1727
rect 282 1722 288 1723
rect 327 1727 333 1728
rect 327 1723 328 1727
rect 332 1726 333 1727
rect 486 1727 492 1728
rect 332 1724 361 1726
rect 332 1723 333 1724
rect 327 1722 333 1723
rect 486 1723 487 1727
rect 491 1726 492 1727
rect 562 1727 568 1728
rect 491 1724 513 1726
rect 491 1723 492 1724
rect 486 1722 492 1723
rect 562 1723 563 1727
rect 567 1726 568 1727
rect 730 1727 736 1728
rect 567 1724 681 1726
rect 567 1723 568 1724
rect 562 1722 568 1723
rect 730 1723 731 1727
rect 735 1726 736 1727
rect 1090 1727 1096 1728
rect 1090 1726 1091 1727
rect 735 1724 857 1726
rect 1069 1724 1091 1726
rect 735 1723 736 1724
rect 730 1722 736 1723
rect 1090 1723 1091 1724
rect 1095 1723 1096 1727
rect 1090 1722 1096 1723
rect 1102 1727 1108 1728
rect 1102 1723 1103 1727
rect 1107 1726 1108 1727
rect 1410 1727 1416 1728
rect 1410 1726 1411 1727
rect 1107 1724 1185 1726
rect 1381 1724 1411 1726
rect 1107 1723 1108 1724
rect 1102 1722 1108 1723
rect 1410 1723 1411 1724
rect 1415 1723 1416 1727
rect 1554 1727 1560 1728
rect 1554 1726 1555 1727
rect 1525 1724 1555 1726
rect 1410 1722 1416 1723
rect 1554 1723 1555 1724
rect 1559 1723 1560 1727
rect 1690 1727 1696 1728
rect 1690 1726 1691 1727
rect 1669 1724 1691 1726
rect 1554 1722 1560 1723
rect 1690 1723 1691 1724
rect 1695 1723 1696 1727
rect 1690 1722 1696 1723
rect 1706 1727 1712 1728
rect 1706 1723 1707 1727
rect 1711 1726 1712 1727
rect 1711 1724 1761 1726
rect 2102 1724 2108 1725
rect 1711 1723 1712 1724
rect 1706 1722 1712 1723
rect 1870 1721 1876 1722
rect 1870 1717 1871 1721
rect 1875 1717 1876 1721
rect 2102 1720 2103 1724
rect 2107 1720 2108 1724
rect 2102 1719 2108 1720
rect 2238 1724 2244 1725
rect 2238 1720 2239 1724
rect 2243 1720 2244 1724
rect 2238 1719 2244 1720
rect 2382 1724 2388 1725
rect 2382 1720 2383 1724
rect 2387 1720 2388 1724
rect 2382 1719 2388 1720
rect 2526 1724 2532 1725
rect 2526 1720 2527 1724
rect 2531 1720 2532 1724
rect 2526 1719 2532 1720
rect 2662 1724 2668 1725
rect 2662 1720 2663 1724
rect 2667 1720 2668 1724
rect 2662 1719 2668 1720
rect 2798 1724 2804 1725
rect 2798 1720 2799 1724
rect 2803 1720 2804 1724
rect 2798 1719 2804 1720
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3046 1724 3052 1725
rect 3046 1720 3047 1724
rect 3051 1720 3052 1724
rect 3046 1719 3052 1720
rect 3158 1724 3164 1725
rect 3158 1720 3159 1724
rect 3163 1720 3164 1724
rect 3158 1719 3164 1720
rect 3270 1724 3276 1725
rect 3270 1720 3271 1724
rect 3275 1720 3276 1724
rect 3270 1719 3276 1720
rect 3390 1724 3396 1725
rect 3390 1720 3391 1724
rect 3395 1720 3396 1724
rect 3390 1719 3396 1720
rect 3502 1724 3508 1725
rect 3502 1720 3503 1724
rect 3507 1720 3508 1724
rect 3502 1719 3508 1720
rect 3590 1721 3596 1722
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 110 1711 116 1712
rect 1830 1716 1836 1717
rect 1870 1716 1876 1717
rect 3590 1717 3591 1721
rect 3595 1717 3596 1721
rect 3590 1716 3596 1717
rect 1830 1712 1831 1716
rect 1835 1712 1836 1716
rect 2186 1715 2192 1716
rect 2186 1714 2187 1715
rect 2165 1712 2187 1714
rect 1830 1711 1836 1712
rect 2186 1711 2187 1712
rect 2191 1711 2192 1715
rect 2330 1715 2336 1716
rect 2330 1714 2331 1715
rect 2301 1712 2331 1714
rect 2186 1710 2192 1711
rect 2330 1711 2331 1712
rect 2335 1711 2336 1715
rect 2450 1715 2456 1716
rect 2450 1714 2451 1715
rect 2445 1712 2451 1714
rect 2330 1710 2336 1711
rect 2450 1711 2451 1712
rect 2455 1711 2456 1715
rect 2594 1715 2600 1716
rect 2450 1710 2456 1711
rect 2588 1706 2590 1713
rect 2594 1711 2595 1715
rect 2599 1714 2600 1715
rect 2898 1715 2904 1716
rect 2898 1714 2899 1715
rect 2599 1712 2681 1714
rect 2861 1712 2899 1714
rect 2599 1711 2600 1712
rect 2594 1710 2600 1711
rect 2898 1711 2899 1712
rect 2903 1711 2904 1715
rect 3002 1715 3008 1716
rect 3002 1714 3003 1715
rect 2989 1712 3003 1714
rect 2898 1710 2904 1711
rect 3002 1711 3003 1712
rect 3007 1711 3008 1715
rect 3118 1715 3124 1716
rect 3002 1710 3008 1711
rect 3108 1708 3110 1713
rect 3118 1711 3119 1715
rect 3123 1714 3124 1715
rect 3226 1715 3232 1716
rect 3123 1712 3177 1714
rect 3123 1711 3124 1712
rect 3118 1710 3124 1711
rect 3226 1711 3227 1715
rect 3231 1714 3232 1715
rect 3458 1715 3464 1716
rect 3458 1714 3459 1715
rect 3231 1712 3289 1714
rect 3453 1712 3459 1714
rect 3231 1711 3232 1712
rect 3226 1710 3232 1711
rect 3458 1711 3459 1712
rect 3463 1711 3464 1715
rect 3458 1710 3464 1711
rect 3564 1708 3566 1713
rect 2654 1707 2660 1708
rect 2654 1706 2655 1707
rect 1870 1704 1876 1705
rect 2588 1704 2655 1706
rect 1870 1700 1871 1704
rect 1875 1700 1876 1704
rect 2654 1703 2655 1704
rect 2659 1703 2660 1707
rect 2654 1702 2660 1703
rect 3106 1707 3112 1708
rect 3106 1703 3107 1707
rect 3111 1703 3112 1707
rect 3106 1702 3112 1703
rect 3562 1707 3568 1708
rect 3562 1703 3563 1707
rect 3567 1703 3568 1707
rect 3562 1702 3568 1703
rect 3590 1704 3596 1705
rect 1870 1699 1876 1700
rect 3590 1700 3591 1704
rect 3595 1700 3596 1704
rect 3590 1699 3596 1700
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 222 1698 228 1699
rect 222 1694 223 1698
rect 227 1694 228 1698
rect 222 1693 228 1694
rect 350 1698 356 1699
rect 350 1694 351 1698
rect 355 1694 356 1698
rect 350 1693 356 1694
rect 502 1698 508 1699
rect 502 1694 503 1698
rect 507 1694 508 1698
rect 502 1693 508 1694
rect 670 1698 676 1699
rect 670 1694 671 1698
rect 675 1694 676 1698
rect 670 1693 676 1694
rect 846 1698 852 1699
rect 846 1694 847 1698
rect 851 1694 852 1698
rect 846 1693 852 1694
rect 1014 1698 1020 1699
rect 1014 1694 1015 1698
rect 1019 1694 1020 1698
rect 1014 1693 1020 1694
rect 1174 1698 1180 1699
rect 1174 1694 1175 1698
rect 1179 1694 1180 1698
rect 1174 1693 1180 1694
rect 1326 1698 1332 1699
rect 1326 1694 1327 1698
rect 1331 1694 1332 1698
rect 1326 1693 1332 1694
rect 1470 1698 1476 1699
rect 1470 1694 1471 1698
rect 1475 1694 1476 1698
rect 1470 1693 1476 1694
rect 1614 1698 1620 1699
rect 1614 1694 1615 1698
rect 1619 1694 1620 1698
rect 1614 1693 1620 1694
rect 1750 1698 1756 1699
rect 1750 1694 1751 1698
rect 1755 1694 1756 1698
rect 1750 1693 1756 1694
rect 166 1687 173 1688
rect 166 1683 167 1687
rect 172 1683 173 1687
rect 166 1682 173 1683
rect 202 1687 208 1688
rect 202 1683 203 1687
rect 207 1686 208 1687
rect 247 1687 253 1688
rect 247 1686 248 1687
rect 207 1684 248 1686
rect 207 1683 208 1684
rect 202 1682 208 1683
rect 247 1683 248 1684
rect 252 1683 253 1687
rect 247 1682 253 1683
rect 282 1687 288 1688
rect 282 1683 283 1687
rect 287 1686 288 1687
rect 375 1687 381 1688
rect 375 1686 376 1687
rect 287 1684 376 1686
rect 287 1683 288 1684
rect 282 1682 288 1683
rect 375 1683 376 1684
rect 380 1683 381 1687
rect 375 1682 381 1683
rect 527 1687 533 1688
rect 527 1683 528 1687
rect 532 1686 533 1687
rect 562 1687 568 1688
rect 562 1686 563 1687
rect 532 1684 563 1686
rect 532 1683 533 1684
rect 527 1682 533 1683
rect 562 1683 563 1684
rect 567 1683 568 1687
rect 562 1682 568 1683
rect 695 1687 701 1688
rect 695 1683 696 1687
rect 700 1686 701 1687
rect 730 1687 736 1688
rect 730 1686 731 1687
rect 700 1684 731 1686
rect 700 1683 701 1684
rect 695 1682 701 1683
rect 730 1683 731 1684
rect 735 1683 736 1687
rect 730 1682 736 1683
rect 814 1687 820 1688
rect 814 1683 815 1687
rect 819 1686 820 1687
rect 871 1687 877 1688
rect 871 1686 872 1687
rect 819 1684 872 1686
rect 819 1683 820 1684
rect 814 1682 820 1683
rect 871 1683 872 1684
rect 876 1683 877 1687
rect 871 1682 877 1683
rect 1038 1687 1045 1688
rect 1038 1683 1039 1687
rect 1044 1683 1045 1687
rect 1038 1682 1045 1683
rect 1090 1687 1096 1688
rect 1090 1683 1091 1687
rect 1095 1686 1096 1687
rect 1199 1687 1205 1688
rect 1199 1686 1200 1687
rect 1095 1684 1200 1686
rect 1095 1683 1096 1684
rect 1090 1682 1096 1683
rect 1199 1683 1200 1684
rect 1204 1683 1205 1687
rect 1199 1682 1205 1683
rect 1351 1687 1360 1688
rect 1351 1683 1352 1687
rect 1359 1683 1360 1687
rect 1351 1682 1360 1683
rect 1410 1687 1416 1688
rect 1410 1683 1411 1687
rect 1415 1686 1416 1687
rect 1495 1687 1501 1688
rect 1495 1686 1496 1687
rect 1415 1684 1496 1686
rect 1415 1683 1416 1684
rect 1410 1682 1416 1683
rect 1495 1683 1496 1684
rect 1500 1683 1501 1687
rect 1495 1682 1501 1683
rect 1554 1687 1560 1688
rect 1554 1683 1555 1687
rect 1559 1686 1560 1687
rect 1639 1687 1645 1688
rect 1639 1686 1640 1687
rect 1559 1684 1640 1686
rect 1559 1683 1560 1684
rect 1554 1682 1560 1683
rect 1639 1683 1640 1684
rect 1644 1683 1645 1687
rect 1639 1682 1645 1683
rect 1690 1687 1696 1688
rect 1690 1683 1691 1687
rect 1695 1686 1696 1687
rect 1775 1687 1781 1688
rect 1775 1686 1776 1687
rect 1695 1684 1776 1686
rect 1695 1683 1696 1684
rect 1690 1682 1696 1683
rect 1775 1683 1776 1684
rect 1780 1683 1781 1687
rect 1775 1682 1781 1683
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2246 1686 2252 1687
rect 2246 1682 2247 1686
rect 2251 1682 2252 1686
rect 2246 1681 2252 1682
rect 2390 1686 2396 1687
rect 2390 1682 2391 1686
rect 2395 1682 2396 1686
rect 2390 1681 2396 1682
rect 2534 1686 2540 1687
rect 2534 1682 2535 1686
rect 2539 1682 2540 1686
rect 2534 1681 2540 1682
rect 2670 1686 2676 1687
rect 2670 1682 2671 1686
rect 2675 1682 2676 1686
rect 2670 1681 2676 1682
rect 2806 1686 2812 1687
rect 2806 1682 2807 1686
rect 2811 1682 2812 1686
rect 2806 1681 2812 1682
rect 2934 1686 2940 1687
rect 2934 1682 2935 1686
rect 2939 1682 2940 1686
rect 2934 1681 2940 1682
rect 3054 1686 3060 1687
rect 3054 1682 3055 1686
rect 3059 1682 3060 1686
rect 3054 1681 3060 1682
rect 3166 1686 3172 1687
rect 3166 1682 3167 1686
rect 3171 1682 3172 1686
rect 3166 1681 3172 1682
rect 3278 1686 3284 1687
rect 3278 1682 3279 1686
rect 3283 1682 3284 1686
rect 3278 1681 3284 1682
rect 3398 1686 3404 1687
rect 3398 1682 3399 1686
rect 3403 1682 3404 1686
rect 3398 1681 3404 1682
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 862 1679 868 1680
rect 862 1678 863 1679
rect 524 1676 863 1678
rect 167 1671 173 1672
rect 167 1667 168 1671
rect 172 1670 173 1671
rect 302 1671 308 1672
rect 302 1670 303 1671
rect 172 1668 303 1670
rect 172 1667 173 1668
rect 167 1666 173 1667
rect 302 1667 303 1668
rect 307 1667 308 1671
rect 302 1666 308 1667
rect 319 1671 325 1672
rect 319 1667 320 1671
rect 324 1670 325 1671
rect 327 1671 333 1672
rect 327 1670 328 1671
rect 324 1668 328 1670
rect 324 1667 325 1668
rect 319 1666 325 1667
rect 327 1667 328 1668
rect 332 1667 333 1671
rect 327 1666 333 1667
rect 503 1671 509 1672
rect 503 1667 504 1671
rect 508 1670 509 1671
rect 524 1670 526 1676
rect 862 1675 863 1676
rect 867 1675 868 1679
rect 862 1674 868 1675
rect 2135 1675 2141 1676
rect 508 1668 526 1670
rect 530 1671 536 1672
rect 508 1667 509 1668
rect 503 1666 509 1667
rect 530 1667 531 1671
rect 535 1670 536 1671
rect 695 1671 701 1672
rect 695 1670 696 1671
rect 535 1668 696 1670
rect 535 1667 536 1668
rect 530 1666 536 1667
rect 695 1667 696 1668
rect 700 1667 701 1671
rect 695 1666 701 1667
rect 879 1671 885 1672
rect 879 1667 880 1671
rect 884 1670 885 1671
rect 914 1671 920 1672
rect 914 1670 915 1671
rect 884 1668 915 1670
rect 884 1667 885 1668
rect 879 1666 885 1667
rect 914 1667 915 1668
rect 919 1667 920 1671
rect 914 1666 920 1667
rect 1055 1671 1064 1672
rect 1055 1667 1056 1671
rect 1063 1667 1064 1671
rect 1055 1666 1064 1667
rect 1223 1671 1229 1672
rect 1223 1667 1224 1671
rect 1228 1670 1229 1671
rect 1366 1671 1372 1672
rect 1366 1670 1367 1671
rect 1228 1668 1367 1670
rect 1228 1667 1229 1668
rect 1223 1666 1229 1667
rect 1366 1667 1367 1668
rect 1371 1667 1372 1671
rect 1366 1666 1372 1667
rect 1383 1671 1389 1672
rect 1383 1667 1384 1671
rect 1388 1670 1389 1671
rect 1526 1671 1532 1672
rect 1526 1670 1527 1671
rect 1388 1668 1527 1670
rect 1388 1667 1389 1668
rect 1383 1666 1389 1667
rect 1526 1667 1527 1668
rect 1531 1667 1532 1671
rect 1526 1666 1532 1667
rect 1543 1671 1549 1672
rect 1543 1667 1544 1671
rect 1548 1670 1549 1671
rect 1686 1671 1692 1672
rect 1686 1670 1687 1671
rect 1548 1668 1687 1670
rect 1548 1667 1549 1668
rect 1543 1666 1549 1667
rect 1686 1667 1687 1668
rect 1691 1667 1692 1671
rect 1686 1666 1692 1667
rect 1703 1671 1712 1672
rect 1703 1667 1704 1671
rect 1711 1667 1712 1671
rect 2135 1671 2136 1675
rect 2140 1674 2141 1675
rect 2186 1675 2192 1676
rect 2140 1672 2182 1674
rect 2140 1671 2141 1672
rect 2135 1670 2141 1671
rect 1703 1666 1712 1667
rect 2180 1666 2182 1672
rect 2186 1671 2187 1675
rect 2191 1674 2192 1675
rect 2271 1675 2277 1676
rect 2271 1674 2272 1675
rect 2191 1672 2272 1674
rect 2191 1671 2192 1672
rect 2186 1670 2192 1671
rect 2271 1671 2272 1672
rect 2276 1671 2277 1675
rect 2271 1670 2277 1671
rect 2330 1675 2336 1676
rect 2330 1671 2331 1675
rect 2335 1674 2336 1675
rect 2415 1675 2421 1676
rect 2415 1674 2416 1675
rect 2335 1672 2416 1674
rect 2335 1671 2336 1672
rect 2330 1670 2336 1671
rect 2415 1671 2416 1672
rect 2420 1671 2421 1675
rect 2415 1670 2421 1671
rect 2559 1675 2565 1676
rect 2559 1671 2560 1675
rect 2564 1674 2565 1675
rect 2594 1675 2600 1676
rect 2594 1674 2595 1675
rect 2564 1672 2595 1674
rect 2564 1671 2565 1672
rect 2559 1670 2565 1671
rect 2594 1671 2595 1672
rect 2599 1671 2600 1675
rect 2594 1670 2600 1671
rect 2695 1675 2704 1676
rect 2695 1671 2696 1675
rect 2703 1671 2704 1675
rect 2695 1670 2704 1671
rect 2831 1675 2840 1676
rect 2831 1671 2832 1675
rect 2839 1671 2840 1675
rect 2831 1670 2840 1671
rect 2898 1675 2904 1676
rect 2898 1671 2899 1675
rect 2903 1674 2904 1675
rect 2959 1675 2965 1676
rect 2959 1674 2960 1675
rect 2903 1672 2960 1674
rect 2903 1671 2904 1672
rect 2898 1670 2904 1671
rect 2959 1671 2960 1672
rect 2964 1671 2965 1675
rect 2959 1670 2965 1671
rect 3002 1675 3008 1676
rect 3002 1671 3003 1675
rect 3007 1674 3008 1675
rect 3079 1675 3085 1676
rect 3079 1674 3080 1675
rect 3007 1672 3080 1674
rect 3007 1671 3008 1672
rect 3002 1670 3008 1671
rect 3079 1671 3080 1672
rect 3084 1671 3085 1675
rect 3079 1670 3085 1671
rect 3191 1675 3197 1676
rect 3191 1671 3192 1675
rect 3196 1674 3197 1675
rect 3226 1675 3232 1676
rect 3226 1674 3227 1675
rect 3196 1672 3227 1674
rect 3196 1671 3197 1672
rect 3191 1670 3197 1671
rect 3226 1671 3227 1672
rect 3231 1671 3232 1675
rect 3226 1670 3232 1671
rect 3303 1675 3309 1676
rect 3303 1671 3304 1675
rect 3308 1674 3309 1675
rect 3382 1675 3388 1676
rect 3382 1674 3383 1675
rect 3308 1672 3383 1674
rect 3308 1671 3309 1672
rect 3303 1670 3309 1671
rect 3382 1671 3383 1672
rect 3387 1671 3388 1675
rect 3382 1670 3388 1671
rect 3423 1675 3432 1676
rect 3423 1671 3424 1675
rect 3431 1671 3432 1675
rect 3423 1670 3432 1671
rect 3458 1675 3464 1676
rect 3458 1671 3459 1675
rect 3463 1674 3464 1675
rect 3535 1675 3541 1676
rect 3535 1674 3536 1675
rect 3463 1672 3536 1674
rect 3463 1671 3464 1672
rect 3458 1670 3464 1671
rect 3535 1671 3536 1672
rect 3540 1671 3541 1675
rect 3535 1670 3541 1671
rect 2358 1667 2364 1668
rect 2358 1666 2359 1667
rect 2180 1664 2359 1666
rect 2358 1663 2359 1664
rect 2363 1663 2364 1667
rect 142 1662 148 1663
rect 142 1658 143 1662
rect 147 1658 148 1662
rect 142 1657 148 1658
rect 294 1662 300 1663
rect 294 1658 295 1662
rect 299 1658 300 1662
rect 294 1657 300 1658
rect 478 1662 484 1663
rect 478 1658 479 1662
rect 483 1658 484 1662
rect 478 1657 484 1658
rect 670 1662 676 1663
rect 670 1658 671 1662
rect 675 1658 676 1662
rect 670 1657 676 1658
rect 854 1662 860 1663
rect 854 1658 855 1662
rect 859 1658 860 1662
rect 854 1657 860 1658
rect 1030 1662 1036 1663
rect 1030 1658 1031 1662
rect 1035 1658 1036 1662
rect 1030 1657 1036 1658
rect 1198 1662 1204 1663
rect 1198 1658 1199 1662
rect 1203 1658 1204 1662
rect 1198 1657 1204 1658
rect 1358 1662 1364 1663
rect 1358 1658 1359 1662
rect 1363 1658 1364 1662
rect 1358 1657 1364 1658
rect 1518 1662 1524 1663
rect 1518 1658 1519 1662
rect 1523 1658 1524 1662
rect 1518 1657 1524 1658
rect 1678 1662 1684 1663
rect 2358 1662 2364 1663
rect 1678 1658 1679 1662
rect 1683 1658 1684 1662
rect 1678 1657 1684 1658
rect 1974 1659 1980 1660
rect 1974 1655 1975 1659
rect 1979 1658 1980 1659
rect 1991 1659 1997 1660
rect 1991 1658 1992 1659
rect 1979 1656 1992 1658
rect 1979 1655 1980 1656
rect 1974 1654 1980 1655
rect 1991 1655 1992 1656
rect 1996 1655 1997 1659
rect 1991 1654 1997 1655
rect 2018 1659 2024 1660
rect 2018 1655 2019 1659
rect 2023 1658 2024 1659
rect 2111 1659 2117 1660
rect 2111 1658 2112 1659
rect 2023 1656 2112 1658
rect 2023 1655 2024 1656
rect 2018 1654 2024 1655
rect 2111 1655 2112 1656
rect 2116 1655 2117 1659
rect 2111 1654 2117 1655
rect 2138 1659 2144 1660
rect 2138 1655 2139 1659
rect 2143 1658 2144 1659
rect 2239 1659 2245 1660
rect 2239 1658 2240 1659
rect 2143 1656 2240 1658
rect 2143 1655 2144 1656
rect 2138 1654 2144 1655
rect 2239 1655 2240 1656
rect 2244 1655 2245 1659
rect 2239 1654 2245 1655
rect 2266 1659 2272 1660
rect 2266 1655 2267 1659
rect 2271 1658 2272 1659
rect 2375 1659 2381 1660
rect 2375 1658 2376 1659
rect 2271 1656 2376 1658
rect 2271 1655 2272 1656
rect 2266 1654 2272 1655
rect 2375 1655 2376 1656
rect 2380 1655 2381 1659
rect 2375 1654 2381 1655
rect 2519 1659 2525 1660
rect 2519 1655 2520 1659
rect 2524 1658 2525 1659
rect 2646 1659 2652 1660
rect 2646 1658 2647 1659
rect 2524 1656 2647 1658
rect 2524 1655 2525 1656
rect 2519 1654 2525 1655
rect 2646 1655 2647 1656
rect 2651 1655 2652 1659
rect 2646 1654 2652 1655
rect 2654 1659 2660 1660
rect 2654 1655 2655 1659
rect 2659 1658 2660 1659
rect 2663 1659 2669 1660
rect 2663 1658 2664 1659
rect 2659 1656 2664 1658
rect 2659 1655 2660 1656
rect 2654 1654 2660 1655
rect 2663 1655 2664 1656
rect 2668 1655 2669 1659
rect 2663 1654 2669 1655
rect 2807 1659 2813 1660
rect 2807 1655 2808 1659
rect 2812 1658 2813 1659
rect 2887 1659 2893 1660
rect 2887 1658 2888 1659
rect 2812 1656 2888 1658
rect 2812 1655 2813 1656
rect 2807 1654 2813 1655
rect 2887 1655 2888 1656
rect 2892 1655 2893 1659
rect 2887 1654 2893 1655
rect 2951 1659 2957 1660
rect 2951 1655 2952 1659
rect 2956 1658 2957 1659
rect 3078 1659 3084 1660
rect 3078 1658 3079 1659
rect 2956 1656 3079 1658
rect 2956 1655 2957 1656
rect 2951 1654 2957 1655
rect 3078 1655 3079 1656
rect 3083 1655 3084 1659
rect 3078 1654 3084 1655
rect 3095 1659 3101 1660
rect 3095 1655 3096 1659
rect 3100 1658 3101 1659
rect 3106 1659 3112 1660
rect 3106 1658 3107 1659
rect 3100 1656 3107 1658
rect 3100 1655 3101 1656
rect 3095 1654 3101 1655
rect 3106 1655 3107 1656
rect 3111 1655 3112 1659
rect 3106 1654 3112 1655
rect 3178 1659 3184 1660
rect 3178 1655 3179 1659
rect 3183 1658 3184 1659
rect 3247 1659 3253 1660
rect 3247 1658 3248 1659
rect 3183 1656 3248 1658
rect 3183 1655 3184 1656
rect 3178 1654 3184 1655
rect 3247 1655 3248 1656
rect 3252 1655 3253 1659
rect 3247 1654 3253 1655
rect 3330 1659 3336 1660
rect 3330 1655 3331 1659
rect 3335 1658 3336 1659
rect 3399 1659 3405 1660
rect 3399 1658 3400 1659
rect 3335 1656 3400 1658
rect 3335 1655 3336 1656
rect 3330 1654 3336 1655
rect 3399 1655 3400 1656
rect 3404 1655 3405 1659
rect 3399 1654 3405 1655
rect 3535 1659 3541 1660
rect 3535 1655 3536 1659
rect 3540 1658 3541 1659
rect 3562 1659 3568 1660
rect 3562 1658 3563 1659
rect 3540 1656 3563 1658
rect 3540 1655 3541 1656
rect 3535 1654 3541 1655
rect 3562 1655 3563 1656
rect 3567 1655 3568 1659
rect 3562 1654 3568 1655
rect 1966 1650 1972 1651
rect 1966 1646 1967 1650
rect 1971 1646 1972 1650
rect 1966 1645 1972 1646
rect 2086 1650 2092 1651
rect 2086 1646 2087 1650
rect 2091 1646 2092 1650
rect 2086 1645 2092 1646
rect 2214 1650 2220 1651
rect 2214 1646 2215 1650
rect 2219 1646 2220 1650
rect 2214 1645 2220 1646
rect 2350 1650 2356 1651
rect 2350 1646 2351 1650
rect 2355 1646 2356 1650
rect 2350 1645 2356 1646
rect 2494 1650 2500 1651
rect 2494 1646 2495 1650
rect 2499 1646 2500 1650
rect 2494 1645 2500 1646
rect 2638 1650 2644 1651
rect 2638 1646 2639 1650
rect 2643 1646 2644 1650
rect 2638 1645 2644 1646
rect 2782 1650 2788 1651
rect 2782 1646 2783 1650
rect 2787 1646 2788 1650
rect 2782 1645 2788 1646
rect 2926 1650 2932 1651
rect 2926 1646 2927 1650
rect 2931 1646 2932 1650
rect 2926 1645 2932 1646
rect 3070 1650 3076 1651
rect 3070 1646 3071 1650
rect 3075 1646 3076 1650
rect 3070 1645 3076 1646
rect 3222 1650 3228 1651
rect 3222 1646 3223 1650
rect 3227 1646 3228 1650
rect 3222 1645 3228 1646
rect 3374 1650 3380 1651
rect 3374 1646 3375 1650
rect 3379 1646 3380 1650
rect 3374 1645 3380 1646
rect 3510 1650 3516 1651
rect 3510 1646 3511 1650
rect 3515 1646 3516 1650
rect 3510 1645 3516 1646
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 110 1639 116 1640
rect 1830 1644 1836 1645
rect 1830 1640 1831 1644
rect 1835 1640 1836 1644
rect 1830 1639 1836 1640
rect 190 1635 196 1636
rect 190 1631 191 1635
rect 195 1631 196 1635
rect 190 1630 196 1631
rect 302 1635 308 1636
rect 302 1631 303 1635
rect 307 1631 308 1635
rect 302 1630 308 1631
rect 530 1635 536 1636
rect 530 1631 531 1635
rect 535 1631 536 1635
rect 814 1635 820 1636
rect 814 1634 815 1635
rect 725 1632 815 1634
rect 530 1630 536 1631
rect 814 1631 815 1632
rect 819 1631 820 1635
rect 814 1630 820 1631
rect 862 1635 868 1636
rect 862 1631 863 1635
rect 867 1631 868 1635
rect 862 1630 868 1631
rect 1038 1635 1044 1636
rect 1038 1631 1039 1635
rect 1043 1631 1044 1635
rect 1262 1635 1268 1636
rect 1262 1634 1263 1635
rect 1253 1632 1263 1634
rect 1038 1630 1044 1631
rect 1262 1631 1263 1632
rect 1267 1631 1268 1635
rect 1262 1630 1268 1631
rect 1366 1635 1372 1636
rect 1366 1631 1367 1635
rect 1371 1631 1372 1635
rect 1366 1630 1372 1631
rect 1526 1635 1532 1636
rect 1526 1631 1527 1635
rect 1531 1631 1532 1635
rect 1526 1630 1532 1631
rect 1686 1635 1692 1636
rect 1686 1631 1687 1635
rect 1691 1631 1692 1635
rect 1686 1630 1692 1631
rect 1870 1632 1876 1633
rect 1870 1628 1871 1632
rect 1875 1628 1876 1632
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 1830 1627 1836 1628
rect 1870 1627 1876 1628
rect 3590 1632 3596 1633
rect 3590 1628 3591 1632
rect 3595 1628 3596 1632
rect 3590 1627 3596 1628
rect 110 1622 116 1623
rect 134 1624 140 1625
rect 134 1620 135 1624
rect 139 1620 140 1624
rect 134 1619 140 1620
rect 286 1624 292 1625
rect 286 1620 287 1624
rect 291 1620 292 1624
rect 286 1619 292 1620
rect 470 1624 476 1625
rect 470 1620 471 1624
rect 475 1620 476 1624
rect 470 1619 476 1620
rect 662 1624 668 1625
rect 662 1620 663 1624
rect 667 1620 668 1624
rect 662 1619 668 1620
rect 846 1624 852 1625
rect 846 1620 847 1624
rect 851 1620 852 1624
rect 846 1619 852 1620
rect 1022 1624 1028 1625
rect 1022 1620 1023 1624
rect 1027 1620 1028 1624
rect 1022 1619 1028 1620
rect 1190 1624 1196 1625
rect 1190 1620 1191 1624
rect 1195 1620 1196 1624
rect 1190 1619 1196 1620
rect 1350 1624 1356 1625
rect 1350 1620 1351 1624
rect 1355 1620 1356 1624
rect 1350 1619 1356 1620
rect 1510 1624 1516 1625
rect 1510 1620 1511 1624
rect 1515 1620 1516 1624
rect 1510 1619 1516 1620
rect 1670 1624 1676 1625
rect 1670 1620 1671 1624
rect 1675 1620 1676 1624
rect 1830 1623 1831 1627
rect 1835 1623 1836 1627
rect 1830 1622 1836 1623
rect 2018 1623 2024 1624
rect 1670 1619 1676 1620
rect 2018 1619 2019 1623
rect 2023 1619 2024 1623
rect 2018 1618 2024 1619
rect 2138 1623 2144 1624
rect 2138 1619 2139 1623
rect 2143 1619 2144 1623
rect 2138 1618 2144 1619
rect 2266 1623 2272 1624
rect 2266 1619 2267 1623
rect 2271 1619 2272 1623
rect 2266 1618 2272 1619
rect 2358 1623 2364 1624
rect 2358 1619 2359 1623
rect 2363 1619 2364 1623
rect 2358 1618 2364 1619
rect 2546 1623 2552 1624
rect 2546 1619 2547 1623
rect 2551 1619 2552 1623
rect 2546 1618 2552 1619
rect 2646 1623 2652 1624
rect 2646 1619 2647 1623
rect 2651 1619 2652 1623
rect 2646 1618 2652 1619
rect 2887 1623 2893 1624
rect 2887 1619 2888 1623
rect 2892 1622 2893 1623
rect 3078 1623 3084 1624
rect 2892 1620 2937 1622
rect 2892 1619 2893 1620
rect 2887 1618 2893 1619
rect 3078 1619 3079 1623
rect 3083 1619 3084 1623
rect 3330 1623 3336 1624
rect 3330 1622 3331 1623
rect 3277 1620 3331 1622
rect 3078 1618 3084 1619
rect 3330 1619 3331 1620
rect 3335 1619 3336 1623
rect 3330 1618 3336 1619
rect 3382 1623 3388 1624
rect 3382 1619 3383 1623
rect 3387 1619 3388 1623
rect 3382 1618 3388 1619
rect 3534 1623 3540 1624
rect 3534 1619 3535 1623
rect 3539 1619 3540 1623
rect 3534 1618 3540 1619
rect 1870 1615 1876 1616
rect 1870 1611 1871 1615
rect 1875 1611 1876 1615
rect 3590 1615 3596 1616
rect 1870 1610 1876 1611
rect 1958 1612 1964 1613
rect 1958 1608 1959 1612
rect 1963 1608 1964 1612
rect 1958 1607 1964 1608
rect 2078 1612 2084 1613
rect 2078 1608 2079 1612
rect 2083 1608 2084 1612
rect 2078 1607 2084 1608
rect 2206 1612 2212 1613
rect 2206 1608 2207 1612
rect 2211 1608 2212 1612
rect 2206 1607 2212 1608
rect 2342 1612 2348 1613
rect 2342 1608 2343 1612
rect 2347 1608 2348 1612
rect 2342 1607 2348 1608
rect 2486 1612 2492 1613
rect 2486 1608 2487 1612
rect 2491 1608 2492 1612
rect 2486 1607 2492 1608
rect 2630 1612 2636 1613
rect 2630 1608 2631 1612
rect 2635 1608 2636 1612
rect 2630 1607 2636 1608
rect 2774 1612 2780 1613
rect 2774 1608 2775 1612
rect 2779 1608 2780 1612
rect 2774 1607 2780 1608
rect 2918 1612 2924 1613
rect 2918 1608 2919 1612
rect 2923 1608 2924 1612
rect 2918 1607 2924 1608
rect 3062 1612 3068 1613
rect 3062 1608 3063 1612
rect 3067 1608 3068 1612
rect 3062 1607 3068 1608
rect 3214 1612 3220 1613
rect 3214 1608 3215 1612
rect 3219 1608 3220 1612
rect 3214 1607 3220 1608
rect 3366 1612 3372 1613
rect 3366 1608 3367 1612
rect 3371 1608 3372 1612
rect 3366 1607 3372 1608
rect 3502 1612 3508 1613
rect 3502 1608 3503 1612
rect 3507 1608 3508 1612
rect 3590 1611 3591 1615
rect 3595 1611 3596 1615
rect 3590 1610 3596 1611
rect 3502 1607 3508 1608
rect 2722 1595 2728 1596
rect 2722 1591 2723 1595
rect 2727 1594 2728 1595
rect 2791 1595 2797 1596
rect 2791 1594 2792 1595
rect 2727 1592 2792 1594
rect 2727 1591 2728 1592
rect 2722 1590 2728 1591
rect 2791 1591 2792 1592
rect 2796 1591 2797 1595
rect 2791 1590 2797 1591
rect 158 1580 164 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 158 1576 159 1580
rect 163 1576 164 1580
rect 158 1575 164 1576
rect 286 1580 292 1581
rect 286 1576 287 1580
rect 291 1576 292 1580
rect 286 1575 292 1576
rect 422 1580 428 1581
rect 422 1576 423 1580
rect 427 1576 428 1580
rect 422 1575 428 1576
rect 566 1580 572 1581
rect 566 1576 567 1580
rect 571 1576 572 1580
rect 566 1575 572 1576
rect 710 1580 716 1581
rect 710 1576 711 1580
rect 715 1576 716 1580
rect 710 1575 716 1576
rect 846 1580 852 1581
rect 846 1576 847 1580
rect 851 1576 852 1580
rect 846 1575 852 1576
rect 982 1580 988 1581
rect 982 1576 983 1580
rect 987 1576 988 1580
rect 982 1575 988 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1246 1580 1252 1581
rect 1246 1576 1247 1580
rect 1251 1576 1252 1580
rect 1246 1575 1252 1576
rect 1374 1580 1380 1581
rect 1374 1576 1375 1580
rect 1379 1576 1380 1580
rect 1374 1575 1380 1576
rect 1510 1580 1516 1581
rect 1510 1576 1511 1580
rect 1515 1576 1516 1580
rect 1510 1575 1516 1576
rect 1830 1577 1836 1578
rect 110 1572 116 1573
rect 1830 1573 1831 1577
rect 1835 1573 1836 1577
rect 1830 1572 1836 1573
rect 230 1571 236 1572
rect 230 1570 231 1571
rect 221 1568 231 1570
rect 230 1567 231 1568
rect 235 1567 236 1571
rect 230 1566 236 1567
rect 258 1571 264 1572
rect 258 1567 259 1571
rect 263 1570 264 1571
rect 534 1571 540 1572
rect 534 1570 535 1571
rect 263 1568 305 1570
rect 485 1568 535 1570
rect 263 1567 264 1568
rect 258 1566 264 1567
rect 534 1567 535 1568
rect 539 1567 540 1571
rect 658 1571 664 1572
rect 658 1570 659 1571
rect 629 1568 659 1570
rect 534 1566 540 1567
rect 658 1567 659 1568
rect 663 1567 664 1571
rect 802 1571 808 1572
rect 802 1570 803 1571
rect 773 1568 803 1570
rect 658 1566 664 1567
rect 802 1567 803 1568
rect 807 1567 808 1571
rect 914 1571 920 1572
rect 914 1570 915 1571
rect 909 1568 915 1570
rect 802 1566 808 1567
rect 914 1567 915 1568
rect 919 1567 920 1571
rect 1050 1571 1056 1572
rect 1050 1570 1051 1571
rect 1045 1568 1051 1570
rect 914 1566 920 1567
rect 1050 1567 1051 1568
rect 1055 1567 1056 1571
rect 1050 1566 1056 1567
rect 1058 1571 1064 1572
rect 1058 1567 1059 1571
rect 1063 1570 1064 1571
rect 1330 1571 1336 1572
rect 1330 1570 1331 1571
rect 1063 1568 1137 1570
rect 1309 1568 1331 1570
rect 1063 1567 1064 1568
rect 1058 1566 1064 1567
rect 1330 1567 1331 1568
rect 1335 1567 1336 1571
rect 1442 1571 1448 1572
rect 1442 1570 1443 1571
rect 1437 1568 1443 1570
rect 1330 1566 1336 1567
rect 1442 1567 1443 1568
rect 1447 1567 1448 1571
rect 1442 1566 1448 1567
rect 1450 1571 1456 1572
rect 1450 1567 1451 1571
rect 1455 1570 1456 1571
rect 1455 1568 1529 1570
rect 1455 1567 1456 1568
rect 1450 1566 1456 1567
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 110 1555 116 1556
rect 1830 1560 1836 1561
rect 1830 1556 1831 1560
rect 1835 1556 1836 1560
rect 1894 1560 1900 1561
rect 1830 1555 1836 1556
rect 1870 1557 1876 1558
rect 1870 1553 1871 1557
rect 1875 1553 1876 1557
rect 1894 1556 1895 1560
rect 1899 1556 1900 1560
rect 1894 1555 1900 1556
rect 2046 1560 2052 1561
rect 2046 1556 2047 1560
rect 2051 1556 2052 1560
rect 2046 1555 2052 1556
rect 2206 1560 2212 1561
rect 2206 1556 2207 1560
rect 2211 1556 2212 1560
rect 2206 1555 2212 1556
rect 2366 1560 2372 1561
rect 2366 1556 2367 1560
rect 2371 1556 2372 1560
rect 2366 1555 2372 1556
rect 2526 1560 2532 1561
rect 2526 1556 2527 1560
rect 2531 1556 2532 1560
rect 2526 1555 2532 1556
rect 2686 1560 2692 1561
rect 2686 1556 2687 1560
rect 2691 1556 2692 1560
rect 2686 1555 2692 1556
rect 2838 1560 2844 1561
rect 2838 1556 2839 1560
rect 2843 1556 2844 1560
rect 2838 1555 2844 1556
rect 2982 1560 2988 1561
rect 2982 1556 2983 1560
rect 2987 1556 2988 1560
rect 2982 1555 2988 1556
rect 3118 1560 3124 1561
rect 3118 1556 3119 1560
rect 3123 1556 3124 1560
rect 3118 1555 3124 1556
rect 3254 1560 3260 1561
rect 3254 1556 3255 1560
rect 3259 1556 3260 1560
rect 3254 1555 3260 1556
rect 3390 1560 3396 1561
rect 3390 1556 3391 1560
rect 3395 1556 3396 1560
rect 3390 1555 3396 1556
rect 3502 1560 3508 1561
rect 3502 1556 3503 1560
rect 3507 1556 3508 1560
rect 3502 1555 3508 1556
rect 3590 1557 3596 1558
rect 1870 1552 1876 1553
rect 3590 1553 3591 1557
rect 3595 1553 3596 1557
rect 3590 1552 3596 1553
rect 1962 1551 1968 1552
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 294 1542 300 1543
rect 294 1538 295 1542
rect 299 1538 300 1542
rect 294 1537 300 1538
rect 430 1542 436 1543
rect 430 1538 431 1542
rect 435 1538 436 1542
rect 430 1537 436 1538
rect 574 1542 580 1543
rect 574 1538 575 1542
rect 579 1538 580 1542
rect 574 1537 580 1538
rect 718 1542 724 1543
rect 718 1538 719 1542
rect 723 1538 724 1542
rect 718 1537 724 1538
rect 854 1542 860 1543
rect 854 1538 855 1542
rect 859 1538 860 1542
rect 854 1537 860 1538
rect 990 1542 996 1543
rect 990 1538 991 1542
rect 995 1538 996 1542
rect 990 1537 996 1538
rect 1126 1542 1132 1543
rect 1126 1538 1127 1542
rect 1131 1538 1132 1542
rect 1126 1537 1132 1538
rect 1254 1542 1260 1543
rect 1254 1538 1255 1542
rect 1259 1538 1260 1542
rect 1254 1537 1260 1538
rect 1382 1542 1388 1543
rect 1382 1538 1383 1542
rect 1387 1538 1388 1542
rect 1382 1537 1388 1538
rect 1518 1542 1524 1543
rect 1518 1538 1519 1542
rect 1523 1538 1524 1542
rect 1956 1542 1958 1549
rect 1962 1547 1963 1551
rect 1967 1550 1968 1551
rect 2114 1551 2120 1552
rect 1967 1548 2065 1550
rect 1967 1547 1968 1548
rect 1962 1546 1968 1547
rect 2114 1547 2115 1551
rect 2119 1550 2120 1551
rect 2434 1551 2440 1552
rect 2119 1548 2225 1550
rect 2119 1547 2120 1548
rect 2114 1546 2120 1547
rect 1974 1543 1980 1544
rect 1974 1542 1975 1543
rect 1518 1537 1524 1538
rect 1870 1540 1876 1541
rect 1956 1540 1975 1542
rect 1870 1536 1871 1540
rect 1875 1536 1876 1540
rect 1974 1539 1975 1540
rect 1979 1539 1980 1543
rect 2428 1542 2430 1549
rect 2434 1547 2435 1551
rect 2439 1550 2440 1551
rect 2754 1551 2760 1552
rect 2754 1550 2755 1551
rect 2439 1548 2545 1550
rect 2749 1548 2755 1550
rect 2439 1547 2440 1548
rect 2434 1546 2440 1547
rect 2754 1547 2755 1548
rect 2759 1547 2760 1551
rect 2930 1551 2936 1552
rect 2930 1550 2931 1551
rect 2901 1548 2931 1550
rect 2754 1546 2760 1547
rect 2930 1547 2931 1548
rect 2935 1547 2936 1551
rect 3054 1551 3060 1552
rect 3054 1550 3055 1551
rect 3045 1548 3055 1550
rect 2930 1546 2936 1547
rect 3054 1547 3055 1548
rect 3059 1547 3060 1551
rect 3186 1551 3192 1552
rect 3054 1546 3060 1547
rect 3180 1544 3182 1549
rect 3186 1547 3187 1551
rect 3191 1550 3192 1551
rect 3322 1551 3328 1552
rect 3191 1548 3273 1550
rect 3191 1547 3192 1548
rect 3186 1546 3192 1547
rect 3322 1547 3323 1551
rect 3327 1550 3328 1551
rect 3327 1548 3409 1550
rect 3327 1547 3328 1548
rect 3322 1546 3328 1547
rect 3564 1544 3566 1549
rect 2442 1543 2448 1544
rect 2442 1542 2443 1543
rect 2428 1540 2443 1542
rect 1974 1538 1980 1539
rect 2442 1539 2443 1540
rect 2447 1539 2448 1543
rect 2442 1538 2448 1539
rect 3178 1543 3184 1544
rect 3178 1539 3179 1543
rect 3183 1539 3184 1543
rect 3178 1538 3184 1539
rect 3562 1543 3568 1544
rect 3562 1539 3563 1543
rect 3567 1539 3568 1543
rect 3562 1538 3568 1539
rect 3590 1540 3596 1541
rect 1870 1535 1876 1536
rect 3590 1536 3591 1540
rect 3595 1536 3596 1540
rect 3590 1535 3596 1536
rect 190 1531 197 1532
rect 190 1527 191 1531
rect 196 1527 197 1531
rect 190 1526 197 1527
rect 230 1531 236 1532
rect 230 1527 231 1531
rect 235 1530 236 1531
rect 319 1531 325 1532
rect 319 1530 320 1531
rect 235 1528 320 1530
rect 235 1527 236 1528
rect 230 1526 236 1527
rect 319 1527 320 1528
rect 324 1527 325 1531
rect 319 1526 325 1527
rect 455 1531 461 1532
rect 455 1527 456 1531
rect 460 1530 461 1531
rect 526 1531 532 1532
rect 526 1530 527 1531
rect 460 1528 527 1530
rect 460 1527 461 1528
rect 455 1526 461 1527
rect 526 1527 527 1528
rect 531 1527 532 1531
rect 526 1526 532 1527
rect 534 1531 540 1532
rect 534 1527 535 1531
rect 539 1530 540 1531
rect 599 1531 605 1532
rect 599 1530 600 1531
rect 539 1528 600 1530
rect 539 1527 540 1528
rect 534 1526 540 1527
rect 599 1527 600 1528
rect 604 1527 605 1531
rect 599 1526 605 1527
rect 658 1531 664 1532
rect 658 1527 659 1531
rect 663 1530 664 1531
rect 743 1531 749 1532
rect 743 1530 744 1531
rect 663 1528 744 1530
rect 663 1527 664 1528
rect 658 1526 664 1527
rect 743 1527 744 1528
rect 748 1527 749 1531
rect 743 1526 749 1527
rect 802 1531 808 1532
rect 802 1527 803 1531
rect 807 1530 808 1531
rect 879 1531 885 1532
rect 879 1530 880 1531
rect 807 1528 880 1530
rect 807 1527 808 1528
rect 802 1526 808 1527
rect 879 1527 880 1528
rect 884 1527 885 1531
rect 879 1526 885 1527
rect 1014 1531 1021 1532
rect 1014 1527 1015 1531
rect 1020 1527 1021 1531
rect 1014 1526 1021 1527
rect 1050 1531 1056 1532
rect 1050 1527 1051 1531
rect 1055 1530 1056 1531
rect 1151 1531 1157 1532
rect 1151 1530 1152 1531
rect 1055 1528 1152 1530
rect 1055 1527 1056 1528
rect 1050 1526 1056 1527
rect 1151 1527 1152 1528
rect 1156 1527 1157 1531
rect 1151 1526 1157 1527
rect 1262 1531 1268 1532
rect 1262 1527 1263 1531
rect 1267 1530 1268 1531
rect 1279 1531 1285 1532
rect 1279 1530 1280 1531
rect 1267 1528 1280 1530
rect 1267 1527 1268 1528
rect 1262 1526 1268 1527
rect 1279 1527 1280 1528
rect 1284 1527 1285 1531
rect 1279 1526 1285 1527
rect 1330 1531 1336 1532
rect 1330 1527 1331 1531
rect 1335 1530 1336 1531
rect 1407 1531 1413 1532
rect 1407 1530 1408 1531
rect 1335 1528 1408 1530
rect 1335 1527 1336 1528
rect 1330 1526 1336 1527
rect 1407 1527 1408 1528
rect 1412 1527 1413 1531
rect 1407 1526 1413 1527
rect 1442 1531 1448 1532
rect 1442 1527 1443 1531
rect 1447 1530 1448 1531
rect 1543 1531 1549 1532
rect 1543 1530 1544 1531
rect 1447 1528 1544 1530
rect 1447 1527 1448 1528
rect 1442 1526 1448 1527
rect 1543 1527 1544 1528
rect 1548 1527 1549 1531
rect 1543 1526 1549 1527
rect 790 1523 796 1524
rect 790 1522 791 1523
rect 668 1520 791 1522
rect 255 1515 264 1516
rect 255 1511 256 1515
rect 263 1511 264 1515
rect 255 1510 264 1511
rect 282 1515 288 1516
rect 282 1511 283 1515
rect 287 1514 288 1515
rect 399 1515 405 1516
rect 399 1514 400 1515
rect 287 1512 400 1514
rect 287 1511 288 1512
rect 282 1510 288 1511
rect 399 1511 400 1512
rect 404 1511 405 1515
rect 399 1510 405 1511
rect 543 1515 549 1516
rect 543 1511 544 1515
rect 548 1514 549 1515
rect 668 1514 670 1520
rect 790 1519 791 1520
rect 795 1519 796 1523
rect 790 1518 796 1519
rect 1902 1522 1908 1523
rect 1902 1518 1903 1522
rect 1907 1518 1908 1522
rect 1902 1517 1908 1518
rect 2054 1522 2060 1523
rect 2054 1518 2055 1522
rect 2059 1518 2060 1522
rect 2054 1517 2060 1518
rect 2214 1522 2220 1523
rect 2214 1518 2215 1522
rect 2219 1518 2220 1522
rect 2214 1517 2220 1518
rect 2374 1522 2380 1523
rect 2374 1518 2375 1522
rect 2379 1518 2380 1522
rect 2374 1517 2380 1518
rect 2534 1522 2540 1523
rect 2534 1518 2535 1522
rect 2539 1518 2540 1522
rect 2534 1517 2540 1518
rect 2694 1522 2700 1523
rect 2694 1518 2695 1522
rect 2699 1518 2700 1522
rect 2694 1517 2700 1518
rect 2846 1522 2852 1523
rect 2846 1518 2847 1522
rect 2851 1518 2852 1522
rect 2846 1517 2852 1518
rect 2990 1522 2996 1523
rect 2990 1518 2991 1522
rect 2995 1518 2996 1522
rect 2990 1517 2996 1518
rect 3126 1522 3132 1523
rect 3126 1518 3127 1522
rect 3131 1518 3132 1522
rect 3126 1517 3132 1518
rect 3262 1522 3268 1523
rect 3262 1518 3263 1522
rect 3267 1518 3268 1522
rect 3262 1517 3268 1518
rect 3398 1522 3404 1523
rect 3398 1518 3399 1522
rect 3403 1518 3404 1522
rect 3398 1517 3404 1518
rect 3510 1522 3516 1523
rect 3510 1518 3511 1522
rect 3515 1518 3516 1522
rect 3510 1517 3516 1518
rect 548 1512 670 1514
rect 679 1515 685 1516
rect 548 1511 549 1512
rect 543 1510 549 1511
rect 679 1511 680 1515
rect 684 1514 685 1515
rect 698 1515 704 1516
rect 698 1514 699 1515
rect 684 1512 699 1514
rect 684 1511 685 1512
rect 679 1510 685 1511
rect 698 1511 699 1512
rect 703 1511 704 1515
rect 698 1510 704 1511
rect 706 1515 712 1516
rect 706 1511 707 1515
rect 711 1514 712 1515
rect 807 1515 813 1516
rect 807 1514 808 1515
rect 711 1512 808 1514
rect 711 1511 712 1512
rect 706 1510 712 1511
rect 807 1511 808 1512
rect 812 1511 813 1515
rect 807 1510 813 1511
rect 926 1515 933 1516
rect 926 1511 927 1515
rect 932 1511 933 1515
rect 926 1510 933 1511
rect 954 1515 960 1516
rect 954 1511 955 1515
rect 959 1514 960 1515
rect 1039 1515 1045 1516
rect 1039 1514 1040 1515
rect 959 1512 1040 1514
rect 959 1511 960 1512
rect 954 1510 960 1511
rect 1039 1511 1040 1512
rect 1044 1511 1045 1515
rect 1039 1510 1045 1511
rect 1143 1515 1149 1516
rect 1143 1511 1144 1515
rect 1148 1514 1149 1515
rect 1154 1515 1160 1516
rect 1154 1514 1155 1515
rect 1148 1512 1155 1514
rect 1148 1511 1149 1512
rect 1143 1510 1149 1511
rect 1154 1511 1155 1512
rect 1159 1511 1160 1515
rect 1154 1510 1160 1511
rect 1170 1515 1176 1516
rect 1170 1511 1171 1515
rect 1175 1514 1176 1515
rect 1239 1515 1245 1516
rect 1239 1514 1240 1515
rect 1175 1512 1240 1514
rect 1175 1511 1176 1512
rect 1170 1510 1176 1511
rect 1239 1511 1240 1512
rect 1244 1511 1245 1515
rect 1239 1510 1245 1511
rect 1266 1515 1272 1516
rect 1266 1511 1267 1515
rect 1271 1514 1272 1515
rect 1343 1515 1349 1516
rect 1343 1514 1344 1515
rect 1271 1512 1344 1514
rect 1271 1511 1272 1512
rect 1266 1510 1272 1511
rect 1343 1511 1344 1512
rect 1348 1511 1349 1515
rect 1343 1510 1349 1511
rect 1447 1515 1456 1516
rect 1447 1511 1448 1515
rect 1455 1511 1456 1515
rect 1447 1510 1456 1511
rect 1927 1511 1933 1512
rect 1927 1507 1928 1511
rect 1932 1510 1933 1511
rect 1962 1511 1968 1512
rect 1962 1510 1963 1511
rect 1932 1508 1963 1510
rect 1932 1507 1933 1508
rect 230 1506 236 1507
rect 230 1502 231 1506
rect 235 1502 236 1506
rect 230 1501 236 1502
rect 374 1506 380 1507
rect 374 1502 375 1506
rect 379 1502 380 1506
rect 374 1501 380 1502
rect 518 1506 524 1507
rect 518 1502 519 1506
rect 523 1502 524 1506
rect 518 1501 524 1502
rect 654 1506 660 1507
rect 654 1502 655 1506
rect 659 1502 660 1506
rect 654 1501 660 1502
rect 782 1506 788 1507
rect 782 1502 783 1506
rect 787 1502 788 1506
rect 782 1501 788 1502
rect 902 1506 908 1507
rect 902 1502 903 1506
rect 907 1502 908 1506
rect 902 1501 908 1502
rect 1014 1506 1020 1507
rect 1014 1502 1015 1506
rect 1019 1502 1020 1506
rect 1014 1501 1020 1502
rect 1118 1506 1124 1507
rect 1118 1502 1119 1506
rect 1123 1502 1124 1506
rect 1118 1501 1124 1502
rect 1214 1506 1220 1507
rect 1214 1502 1215 1506
rect 1219 1502 1220 1506
rect 1214 1501 1220 1502
rect 1318 1506 1324 1507
rect 1318 1502 1319 1506
rect 1323 1502 1324 1506
rect 1318 1501 1324 1502
rect 1422 1506 1428 1507
rect 1927 1506 1933 1507
rect 1962 1507 1963 1508
rect 1967 1507 1968 1511
rect 1962 1506 1968 1507
rect 2079 1511 2085 1512
rect 2079 1507 2080 1511
rect 2084 1510 2085 1511
rect 2114 1511 2120 1512
rect 2114 1510 2115 1511
rect 2084 1508 2115 1510
rect 2084 1507 2085 1508
rect 2079 1506 2085 1507
rect 2114 1507 2115 1508
rect 2119 1507 2120 1511
rect 2114 1506 2120 1507
rect 2186 1511 2192 1512
rect 2186 1507 2187 1511
rect 2191 1510 2192 1511
rect 2239 1511 2245 1512
rect 2239 1510 2240 1511
rect 2191 1508 2240 1510
rect 2191 1507 2192 1508
rect 2186 1506 2192 1507
rect 2239 1507 2240 1508
rect 2244 1507 2245 1511
rect 2239 1506 2245 1507
rect 2399 1511 2405 1512
rect 2399 1507 2400 1511
rect 2404 1510 2405 1511
rect 2434 1511 2440 1512
rect 2434 1510 2435 1511
rect 2404 1508 2435 1510
rect 2404 1507 2405 1508
rect 2399 1506 2405 1507
rect 2434 1507 2435 1508
rect 2439 1507 2440 1511
rect 2434 1506 2440 1507
rect 2546 1511 2552 1512
rect 2546 1507 2547 1511
rect 2551 1510 2552 1511
rect 2559 1511 2565 1512
rect 2559 1510 2560 1511
rect 2551 1508 2560 1510
rect 2551 1507 2552 1508
rect 2546 1506 2552 1507
rect 2559 1507 2560 1508
rect 2564 1507 2565 1511
rect 2559 1506 2565 1507
rect 2719 1511 2728 1512
rect 2719 1507 2720 1511
rect 2727 1507 2728 1511
rect 2719 1506 2728 1507
rect 2754 1511 2760 1512
rect 2754 1507 2755 1511
rect 2759 1510 2760 1511
rect 2871 1511 2877 1512
rect 2871 1510 2872 1511
rect 2759 1508 2872 1510
rect 2759 1507 2760 1508
rect 2754 1506 2760 1507
rect 2871 1507 2872 1508
rect 2876 1507 2877 1511
rect 2871 1506 2877 1507
rect 2930 1511 2936 1512
rect 2930 1507 2931 1511
rect 2935 1510 2936 1511
rect 3015 1511 3021 1512
rect 3015 1510 3016 1511
rect 2935 1508 3016 1510
rect 2935 1507 2936 1508
rect 2930 1506 2936 1507
rect 3015 1507 3016 1508
rect 3020 1507 3021 1511
rect 3015 1506 3021 1507
rect 3151 1511 3157 1512
rect 3151 1507 3152 1511
rect 3156 1510 3157 1511
rect 3186 1511 3192 1512
rect 3186 1510 3187 1511
rect 3156 1508 3187 1510
rect 3156 1507 3157 1508
rect 3151 1506 3157 1507
rect 3186 1507 3187 1508
rect 3191 1507 3192 1511
rect 3186 1506 3192 1507
rect 3287 1511 3293 1512
rect 3287 1507 3288 1511
rect 3292 1510 3293 1511
rect 3322 1511 3328 1512
rect 3322 1510 3323 1511
rect 3292 1508 3323 1510
rect 3292 1507 3293 1508
rect 3287 1506 3293 1507
rect 3322 1507 3323 1508
rect 3327 1507 3328 1511
rect 3322 1506 3328 1507
rect 3418 1511 3429 1512
rect 3418 1507 3419 1511
rect 3423 1507 3424 1511
rect 3428 1507 3429 1511
rect 3418 1506 3429 1507
rect 3534 1511 3541 1512
rect 3534 1507 3535 1511
rect 3540 1507 3541 1511
rect 3534 1506 3541 1507
rect 1422 1502 1423 1506
rect 1427 1502 1428 1506
rect 1422 1501 1428 1502
rect 3518 1499 3524 1500
rect 3518 1498 3519 1499
rect 3244 1496 3519 1498
rect 1927 1491 1933 1492
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 110 1483 116 1484
rect 1830 1488 1836 1489
rect 1830 1484 1831 1488
rect 1835 1484 1836 1488
rect 1927 1487 1928 1491
rect 1932 1490 1933 1491
rect 1962 1491 1968 1492
rect 1962 1490 1963 1491
rect 1932 1488 1963 1490
rect 1932 1487 1933 1488
rect 1927 1486 1933 1487
rect 1962 1487 1963 1488
rect 1967 1487 1968 1491
rect 1962 1486 1968 1487
rect 1970 1491 1976 1492
rect 1970 1487 1971 1491
rect 1975 1490 1976 1491
rect 2031 1491 2037 1492
rect 2031 1490 2032 1491
rect 1975 1488 2032 1490
rect 1975 1487 1976 1488
rect 1970 1486 1976 1487
rect 2031 1487 2032 1488
rect 2036 1487 2037 1491
rect 2031 1486 2037 1487
rect 2126 1491 2132 1492
rect 2126 1487 2127 1491
rect 2131 1490 2132 1491
rect 2159 1491 2165 1492
rect 2159 1490 2160 1491
rect 2131 1488 2160 1490
rect 2131 1487 2132 1488
rect 2126 1486 2132 1487
rect 2159 1487 2160 1488
rect 2164 1487 2165 1491
rect 2159 1486 2165 1487
rect 2295 1491 2301 1492
rect 2295 1487 2296 1491
rect 2300 1490 2301 1491
rect 2422 1491 2428 1492
rect 2422 1490 2423 1491
rect 2300 1488 2423 1490
rect 2300 1487 2301 1488
rect 2295 1486 2301 1487
rect 2422 1487 2423 1488
rect 2427 1487 2428 1491
rect 2422 1486 2428 1487
rect 2439 1491 2448 1492
rect 2439 1487 2440 1491
rect 2447 1487 2448 1491
rect 2439 1486 2448 1487
rect 2591 1491 2597 1492
rect 2591 1487 2592 1491
rect 2596 1490 2597 1491
rect 2726 1491 2732 1492
rect 2726 1490 2727 1491
rect 2596 1488 2727 1490
rect 2596 1487 2597 1488
rect 2591 1486 2597 1487
rect 2726 1487 2727 1488
rect 2731 1487 2732 1491
rect 2726 1486 2732 1487
rect 2743 1491 2749 1492
rect 2743 1487 2744 1491
rect 2748 1490 2749 1491
rect 2886 1491 2892 1492
rect 2886 1490 2887 1491
rect 2748 1488 2887 1490
rect 2748 1487 2749 1488
rect 2743 1486 2749 1487
rect 2886 1487 2887 1488
rect 2891 1487 2892 1491
rect 2886 1486 2892 1487
rect 2903 1491 2909 1492
rect 2903 1487 2904 1491
rect 2908 1490 2909 1491
rect 3046 1491 3052 1492
rect 3046 1490 3047 1491
rect 2908 1488 3047 1490
rect 2908 1487 2909 1488
rect 2903 1486 2909 1487
rect 3046 1487 3047 1488
rect 3051 1487 3052 1491
rect 3046 1486 3052 1487
rect 3054 1491 3060 1492
rect 3054 1487 3055 1491
rect 3059 1490 3060 1491
rect 3063 1491 3069 1492
rect 3063 1490 3064 1491
rect 3059 1488 3064 1490
rect 3059 1487 3060 1488
rect 3054 1486 3060 1487
rect 3063 1487 3064 1488
rect 3068 1487 3069 1491
rect 3063 1486 3069 1487
rect 3223 1491 3229 1492
rect 3223 1487 3224 1491
rect 3228 1490 3229 1491
rect 3244 1490 3246 1496
rect 3518 1495 3519 1496
rect 3523 1495 3524 1499
rect 3518 1494 3524 1495
rect 3228 1488 3246 1490
rect 3250 1491 3256 1492
rect 3228 1487 3229 1488
rect 3223 1486 3229 1487
rect 3250 1487 3251 1491
rect 3255 1490 3256 1491
rect 3391 1491 3397 1492
rect 3391 1490 3392 1491
rect 3255 1488 3392 1490
rect 3255 1487 3256 1488
rect 3250 1486 3256 1487
rect 3391 1487 3392 1488
rect 3396 1487 3397 1491
rect 3391 1486 3397 1487
rect 3535 1491 3541 1492
rect 3535 1487 3536 1491
rect 3540 1490 3541 1491
rect 3562 1491 3568 1492
rect 3562 1490 3563 1491
rect 3540 1488 3563 1490
rect 3540 1487 3541 1488
rect 3535 1486 3541 1487
rect 3562 1487 3563 1488
rect 3567 1487 3568 1491
rect 3562 1486 3568 1487
rect 1830 1483 1836 1484
rect 1902 1482 1908 1483
rect 282 1479 288 1480
rect 282 1475 283 1479
rect 287 1475 288 1479
rect 282 1474 288 1475
rect 426 1479 432 1480
rect 426 1475 427 1479
rect 431 1475 432 1479
rect 426 1474 432 1475
rect 526 1479 532 1480
rect 526 1475 527 1479
rect 531 1475 532 1479
rect 526 1474 532 1475
rect 706 1479 712 1480
rect 706 1475 707 1479
rect 711 1475 712 1479
rect 706 1474 712 1475
rect 790 1479 796 1480
rect 790 1475 791 1479
rect 795 1475 796 1479
rect 790 1474 796 1475
rect 954 1479 960 1480
rect 954 1475 955 1479
rect 959 1475 960 1479
rect 954 1474 960 1475
rect 1022 1479 1028 1480
rect 1022 1475 1023 1479
rect 1027 1475 1028 1479
rect 1022 1474 1028 1475
rect 1170 1479 1176 1480
rect 1170 1475 1171 1479
rect 1175 1475 1176 1479
rect 1170 1474 1176 1475
rect 1266 1479 1272 1480
rect 1266 1475 1267 1479
rect 1271 1475 1272 1479
rect 1266 1474 1272 1475
rect 1370 1479 1376 1480
rect 1370 1475 1371 1479
rect 1375 1475 1376 1479
rect 1370 1474 1376 1475
rect 1430 1479 1436 1480
rect 1430 1475 1431 1479
rect 1435 1475 1436 1479
rect 1902 1478 1903 1482
rect 1907 1478 1908 1482
rect 1902 1477 1908 1478
rect 2006 1482 2012 1483
rect 2006 1478 2007 1482
rect 2011 1478 2012 1482
rect 2006 1477 2012 1478
rect 2134 1482 2140 1483
rect 2134 1478 2135 1482
rect 2139 1478 2140 1482
rect 2134 1477 2140 1478
rect 2270 1482 2276 1483
rect 2270 1478 2271 1482
rect 2275 1478 2276 1482
rect 2270 1477 2276 1478
rect 2414 1482 2420 1483
rect 2414 1478 2415 1482
rect 2419 1478 2420 1482
rect 2414 1477 2420 1478
rect 2566 1482 2572 1483
rect 2566 1478 2567 1482
rect 2571 1478 2572 1482
rect 2566 1477 2572 1478
rect 2718 1482 2724 1483
rect 2718 1478 2719 1482
rect 2723 1478 2724 1482
rect 2718 1477 2724 1478
rect 2878 1482 2884 1483
rect 2878 1478 2879 1482
rect 2883 1478 2884 1482
rect 2878 1477 2884 1478
rect 3038 1482 3044 1483
rect 3038 1478 3039 1482
rect 3043 1478 3044 1482
rect 3038 1477 3044 1478
rect 3198 1482 3204 1483
rect 3198 1478 3199 1482
rect 3203 1478 3204 1482
rect 3198 1477 3204 1478
rect 3366 1482 3372 1483
rect 3366 1478 3367 1482
rect 3371 1478 3372 1482
rect 3366 1477 3372 1478
rect 3510 1482 3516 1483
rect 3510 1478 3511 1482
rect 3515 1478 3516 1482
rect 3510 1477 3516 1478
rect 1430 1474 1436 1475
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 1830 1471 1836 1472
rect 110 1466 116 1467
rect 222 1468 228 1469
rect 222 1464 223 1468
rect 227 1464 228 1468
rect 222 1463 228 1464
rect 366 1468 372 1469
rect 366 1464 367 1468
rect 371 1464 372 1468
rect 366 1463 372 1464
rect 510 1468 516 1469
rect 510 1464 511 1468
rect 515 1464 516 1468
rect 510 1463 516 1464
rect 646 1468 652 1469
rect 646 1464 647 1468
rect 651 1464 652 1468
rect 646 1463 652 1464
rect 774 1468 780 1469
rect 774 1464 775 1468
rect 779 1464 780 1468
rect 774 1463 780 1464
rect 894 1468 900 1469
rect 894 1464 895 1468
rect 899 1464 900 1468
rect 894 1463 900 1464
rect 1006 1468 1012 1469
rect 1006 1464 1007 1468
rect 1011 1464 1012 1468
rect 1006 1463 1012 1464
rect 1110 1468 1116 1469
rect 1110 1464 1111 1468
rect 1115 1464 1116 1468
rect 1110 1463 1116 1464
rect 1206 1468 1212 1469
rect 1206 1464 1207 1468
rect 1211 1464 1212 1468
rect 1206 1463 1212 1464
rect 1310 1468 1316 1469
rect 1310 1464 1311 1468
rect 1315 1464 1316 1468
rect 1310 1463 1316 1464
rect 1414 1468 1420 1469
rect 1414 1464 1415 1468
rect 1419 1464 1420 1468
rect 1830 1467 1831 1471
rect 1835 1467 1836 1471
rect 1830 1466 1836 1467
rect 1414 1463 1420 1464
rect 1870 1464 1876 1465
rect 1870 1460 1871 1464
rect 1875 1460 1876 1464
rect 1870 1459 1876 1460
rect 3590 1464 3596 1465
rect 3590 1460 3591 1464
rect 3595 1460 3596 1464
rect 3590 1459 3596 1460
rect 1970 1455 1976 1456
rect 1970 1454 1971 1455
rect 1957 1452 1971 1454
rect 1970 1451 1971 1452
rect 1975 1451 1976 1455
rect 2126 1455 2132 1456
rect 2126 1454 2127 1455
rect 2061 1452 2127 1454
rect 1970 1450 1976 1451
rect 2126 1451 2127 1452
rect 2131 1451 2132 1455
rect 2126 1450 2132 1451
rect 2186 1455 2192 1456
rect 2186 1451 2187 1455
rect 2191 1451 2192 1455
rect 2186 1450 2192 1451
rect 2422 1455 2428 1456
rect 2422 1451 2423 1455
rect 2427 1451 2428 1455
rect 2422 1450 2428 1451
rect 2726 1455 2732 1456
rect 2726 1451 2727 1455
rect 2731 1451 2732 1455
rect 2726 1450 2732 1451
rect 2886 1455 2892 1456
rect 2886 1451 2887 1455
rect 2891 1451 2892 1455
rect 2886 1450 2892 1451
rect 3046 1455 3052 1456
rect 3046 1451 3047 1455
rect 3051 1451 3052 1455
rect 3046 1450 3052 1451
rect 3250 1455 3256 1456
rect 3250 1451 3251 1455
rect 3255 1451 3256 1455
rect 3250 1450 3256 1451
rect 3418 1455 3424 1456
rect 3418 1451 3419 1455
rect 3423 1451 3424 1455
rect 3418 1450 3424 1451
rect 3518 1455 3524 1456
rect 3518 1451 3519 1455
rect 3523 1451 3524 1455
rect 3518 1450 3524 1451
rect 1870 1447 1876 1448
rect 1870 1443 1871 1447
rect 1875 1443 1876 1447
rect 3590 1447 3596 1448
rect 1870 1442 1876 1443
rect 1894 1444 1900 1445
rect 1894 1440 1895 1444
rect 1899 1440 1900 1444
rect 1894 1439 1900 1440
rect 1998 1444 2004 1445
rect 1998 1440 1999 1444
rect 2003 1440 2004 1444
rect 1998 1439 2004 1440
rect 2126 1444 2132 1445
rect 2126 1440 2127 1444
rect 2131 1440 2132 1444
rect 2126 1439 2132 1440
rect 2262 1444 2268 1445
rect 2262 1440 2263 1444
rect 2267 1440 2268 1444
rect 2262 1439 2268 1440
rect 2406 1444 2412 1445
rect 2406 1440 2407 1444
rect 2411 1440 2412 1444
rect 2406 1439 2412 1440
rect 2558 1444 2564 1445
rect 2558 1440 2559 1444
rect 2563 1440 2564 1444
rect 2558 1439 2564 1440
rect 2710 1444 2716 1445
rect 2710 1440 2711 1444
rect 2715 1440 2716 1444
rect 2710 1439 2716 1440
rect 2870 1444 2876 1445
rect 2870 1440 2871 1444
rect 2875 1440 2876 1444
rect 2870 1439 2876 1440
rect 3030 1444 3036 1445
rect 3030 1440 3031 1444
rect 3035 1440 3036 1444
rect 3030 1439 3036 1440
rect 3190 1444 3196 1445
rect 3190 1440 3191 1444
rect 3195 1440 3196 1444
rect 3190 1439 3196 1440
rect 3358 1444 3364 1445
rect 3358 1440 3359 1444
rect 3363 1440 3364 1444
rect 3358 1439 3364 1440
rect 3502 1444 3508 1445
rect 3502 1440 3503 1444
rect 3507 1440 3508 1444
rect 3590 1443 3591 1447
rect 3595 1443 3596 1447
rect 3590 1442 3596 1443
rect 3502 1439 3508 1440
rect 2058 1427 2064 1428
rect 2058 1423 2059 1427
rect 2063 1426 2064 1427
rect 2279 1427 2285 1428
rect 2279 1426 2280 1427
rect 2063 1424 2280 1426
rect 2063 1423 2064 1424
rect 2058 1422 2064 1423
rect 2279 1423 2280 1424
rect 2284 1423 2285 1427
rect 2279 1422 2285 1423
rect 2466 1427 2472 1428
rect 2466 1423 2467 1427
rect 2471 1426 2472 1427
rect 2575 1427 2581 1428
rect 2575 1426 2576 1427
rect 2471 1424 2576 1426
rect 2471 1423 2472 1424
rect 2466 1422 2472 1423
rect 2575 1423 2576 1424
rect 2580 1423 2581 1427
rect 2575 1422 2581 1423
rect 254 1416 260 1417
rect 110 1413 116 1414
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 254 1412 255 1416
rect 259 1412 260 1416
rect 254 1411 260 1412
rect 350 1416 356 1417
rect 350 1412 351 1416
rect 355 1412 356 1416
rect 350 1411 356 1412
rect 446 1416 452 1417
rect 446 1412 447 1416
rect 451 1412 452 1416
rect 446 1411 452 1412
rect 542 1416 548 1417
rect 542 1412 543 1416
rect 547 1412 548 1416
rect 542 1411 548 1412
rect 630 1416 636 1417
rect 630 1412 631 1416
rect 635 1412 636 1416
rect 630 1411 636 1412
rect 718 1416 724 1417
rect 718 1412 719 1416
rect 723 1412 724 1416
rect 718 1411 724 1412
rect 806 1416 812 1417
rect 806 1412 807 1416
rect 811 1412 812 1416
rect 806 1411 812 1412
rect 918 1416 924 1417
rect 918 1412 919 1416
rect 923 1412 924 1416
rect 918 1411 924 1412
rect 1046 1416 1052 1417
rect 1046 1412 1047 1416
rect 1051 1412 1052 1416
rect 1046 1411 1052 1412
rect 1206 1416 1212 1417
rect 1206 1412 1207 1416
rect 1211 1412 1212 1416
rect 1206 1411 1212 1412
rect 1382 1416 1388 1417
rect 1382 1412 1383 1416
rect 1387 1412 1388 1416
rect 1382 1411 1388 1412
rect 1574 1416 1580 1417
rect 1574 1412 1575 1416
rect 1579 1412 1580 1416
rect 1574 1411 1580 1412
rect 1742 1416 1748 1417
rect 1742 1412 1743 1416
rect 1747 1412 1748 1416
rect 1742 1411 1748 1412
rect 1830 1413 1836 1414
rect 110 1408 116 1409
rect 1830 1409 1831 1413
rect 1835 1409 1836 1413
rect 1830 1408 1836 1409
rect 342 1407 348 1408
rect 316 1400 318 1405
rect 342 1403 343 1407
rect 347 1406 348 1407
rect 418 1407 424 1408
rect 347 1404 369 1406
rect 347 1403 348 1404
rect 342 1402 348 1403
rect 418 1403 419 1407
rect 423 1406 424 1407
rect 610 1407 616 1408
rect 610 1406 611 1407
rect 423 1404 465 1406
rect 605 1404 611 1406
rect 423 1403 424 1404
rect 418 1402 424 1403
rect 610 1403 611 1404
rect 615 1403 616 1407
rect 698 1407 704 1408
rect 698 1406 699 1407
rect 693 1404 699 1406
rect 610 1402 616 1403
rect 698 1403 699 1404
rect 703 1403 704 1407
rect 786 1407 792 1408
rect 698 1402 704 1403
rect 314 1399 320 1400
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 314 1395 315 1399
rect 319 1395 320 1399
rect 314 1394 320 1395
rect 602 1399 608 1400
rect 602 1395 603 1399
rect 607 1398 608 1399
rect 736 1398 738 1405
rect 786 1403 787 1407
rect 791 1406 792 1407
rect 986 1407 992 1408
rect 791 1404 825 1406
rect 791 1403 792 1404
rect 786 1402 792 1403
rect 926 1403 932 1404
rect 926 1399 927 1403
rect 931 1402 932 1403
rect 936 1402 938 1405
rect 986 1403 987 1407
rect 991 1406 992 1407
rect 1114 1407 1120 1408
rect 991 1404 1065 1406
rect 991 1403 992 1404
rect 986 1402 992 1403
rect 1114 1403 1115 1407
rect 1119 1406 1120 1407
rect 1502 1407 1508 1408
rect 1502 1406 1503 1407
rect 1119 1404 1225 1406
rect 1445 1404 1503 1406
rect 1119 1403 1120 1404
rect 1114 1402 1120 1403
rect 1502 1403 1503 1404
rect 1507 1403 1508 1407
rect 1502 1402 1508 1403
rect 1518 1407 1524 1408
rect 1518 1403 1519 1407
rect 1523 1406 1524 1407
rect 1810 1407 1816 1408
rect 1810 1406 1811 1407
rect 1523 1404 1593 1406
rect 1805 1404 1811 1406
rect 1523 1403 1524 1404
rect 1518 1402 1524 1403
rect 1810 1403 1811 1404
rect 1815 1403 1816 1407
rect 1810 1402 1816 1403
rect 931 1400 938 1402
rect 1894 1400 1900 1401
rect 931 1399 932 1400
rect 926 1398 932 1399
rect 607 1396 738 1398
rect 1870 1397 1876 1398
rect 1830 1396 1836 1397
rect 607 1395 608 1396
rect 602 1394 608 1395
rect 110 1391 116 1392
rect 1830 1392 1831 1396
rect 1835 1392 1836 1396
rect 1870 1393 1871 1397
rect 1875 1393 1876 1397
rect 1894 1396 1895 1400
rect 1899 1396 1900 1400
rect 1894 1395 1900 1396
rect 2022 1400 2028 1401
rect 2022 1396 2023 1400
rect 2027 1396 2028 1400
rect 2022 1395 2028 1396
rect 2166 1400 2172 1401
rect 2166 1396 2167 1400
rect 2171 1396 2172 1400
rect 2166 1395 2172 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2430 1400 2436 1401
rect 2430 1396 2431 1400
rect 2435 1396 2436 1400
rect 2430 1395 2436 1396
rect 2550 1400 2556 1401
rect 2550 1396 2551 1400
rect 2555 1396 2556 1400
rect 2550 1395 2556 1396
rect 2670 1400 2676 1401
rect 2670 1396 2671 1400
rect 2675 1396 2676 1400
rect 2670 1395 2676 1396
rect 2790 1400 2796 1401
rect 2790 1396 2791 1400
rect 2795 1396 2796 1400
rect 2790 1395 2796 1396
rect 2910 1400 2916 1401
rect 2910 1396 2911 1400
rect 2915 1396 2916 1400
rect 2910 1395 2916 1396
rect 3590 1397 3596 1398
rect 1870 1392 1876 1393
rect 3590 1393 3591 1397
rect 3595 1393 3596 1397
rect 3590 1392 3596 1393
rect 1830 1391 1836 1392
rect 1962 1391 1968 1392
rect 1962 1390 1963 1391
rect 1957 1388 1963 1390
rect 870 1387 876 1388
rect 870 1383 871 1387
rect 875 1386 876 1387
rect 986 1387 992 1388
rect 986 1386 987 1387
rect 875 1384 987 1386
rect 875 1383 876 1384
rect 870 1382 876 1383
rect 986 1383 987 1384
rect 991 1383 992 1387
rect 1962 1387 1963 1388
rect 1967 1387 1968 1391
rect 2114 1391 2120 1392
rect 2114 1390 2115 1391
rect 2085 1388 2115 1390
rect 1962 1386 1968 1387
rect 2114 1387 2115 1388
rect 2119 1387 2120 1391
rect 2258 1391 2264 1392
rect 2258 1390 2259 1391
rect 2229 1388 2259 1390
rect 2114 1386 2120 1387
rect 2258 1387 2259 1388
rect 2263 1387 2264 1391
rect 2378 1391 2384 1392
rect 2378 1390 2379 1391
rect 2365 1388 2379 1390
rect 2258 1386 2264 1387
rect 2378 1387 2379 1388
rect 2383 1387 2384 1391
rect 2514 1391 2520 1392
rect 2514 1390 2515 1391
rect 2493 1388 2515 1390
rect 2378 1386 2384 1387
rect 2514 1387 2515 1388
rect 2519 1387 2520 1391
rect 2634 1391 2640 1392
rect 2634 1390 2635 1391
rect 2613 1388 2635 1390
rect 2514 1386 2520 1387
rect 2634 1387 2635 1388
rect 2639 1387 2640 1391
rect 2754 1391 2760 1392
rect 2754 1390 2755 1391
rect 2733 1388 2755 1390
rect 2634 1386 2640 1387
rect 2754 1387 2755 1388
rect 2759 1387 2760 1391
rect 2866 1391 2872 1392
rect 2866 1390 2867 1391
rect 2853 1388 2867 1390
rect 2754 1386 2760 1387
rect 2866 1387 2867 1388
rect 2871 1387 2872 1391
rect 2866 1386 2872 1387
rect 2874 1391 2880 1392
rect 2874 1387 2875 1391
rect 2879 1390 2880 1391
rect 2879 1388 2929 1390
rect 2879 1387 2880 1388
rect 2874 1386 2880 1387
rect 986 1382 992 1383
rect 1870 1380 1876 1381
rect 262 1378 268 1379
rect 262 1374 263 1378
rect 267 1374 268 1378
rect 262 1373 268 1374
rect 358 1378 364 1379
rect 358 1374 359 1378
rect 363 1374 364 1378
rect 358 1373 364 1374
rect 454 1378 460 1379
rect 454 1374 455 1378
rect 459 1374 460 1378
rect 454 1373 460 1374
rect 550 1378 556 1379
rect 550 1374 551 1378
rect 555 1374 556 1378
rect 550 1373 556 1374
rect 638 1378 644 1379
rect 638 1374 639 1378
rect 643 1374 644 1378
rect 638 1373 644 1374
rect 726 1378 732 1379
rect 726 1374 727 1378
rect 731 1374 732 1378
rect 726 1373 732 1374
rect 814 1378 820 1379
rect 814 1374 815 1378
rect 819 1374 820 1378
rect 814 1373 820 1374
rect 926 1378 932 1379
rect 926 1374 927 1378
rect 931 1374 932 1378
rect 926 1373 932 1374
rect 1054 1378 1060 1379
rect 1054 1374 1055 1378
rect 1059 1374 1060 1378
rect 1054 1373 1060 1374
rect 1214 1378 1220 1379
rect 1214 1374 1215 1378
rect 1219 1374 1220 1378
rect 1214 1373 1220 1374
rect 1390 1378 1396 1379
rect 1390 1374 1391 1378
rect 1395 1374 1396 1378
rect 1390 1373 1396 1374
rect 1582 1378 1588 1379
rect 1582 1374 1583 1378
rect 1587 1374 1588 1378
rect 1582 1373 1588 1374
rect 1750 1378 1756 1379
rect 1750 1374 1751 1378
rect 1755 1374 1756 1378
rect 1870 1376 1871 1380
rect 1875 1376 1876 1380
rect 1870 1375 1876 1376
rect 3590 1380 3596 1381
rect 3590 1376 3591 1380
rect 3595 1376 3596 1380
rect 3590 1375 3596 1376
rect 1750 1373 1756 1374
rect 287 1367 293 1368
rect 287 1363 288 1367
rect 292 1366 293 1367
rect 342 1367 348 1368
rect 342 1366 343 1367
rect 292 1364 343 1366
rect 292 1363 293 1364
rect 287 1362 293 1363
rect 342 1363 343 1364
rect 347 1363 348 1367
rect 342 1362 348 1363
rect 383 1367 389 1368
rect 383 1363 384 1367
rect 388 1366 389 1367
rect 418 1367 424 1368
rect 418 1366 419 1367
rect 388 1364 419 1366
rect 388 1363 389 1364
rect 383 1362 389 1363
rect 418 1363 419 1364
rect 423 1363 424 1367
rect 418 1362 424 1363
rect 426 1367 432 1368
rect 426 1363 427 1367
rect 431 1366 432 1367
rect 479 1367 485 1368
rect 479 1366 480 1367
rect 431 1364 480 1366
rect 431 1363 432 1364
rect 426 1362 432 1363
rect 479 1363 480 1364
rect 484 1363 485 1367
rect 479 1362 485 1363
rect 575 1367 581 1368
rect 575 1363 576 1367
rect 580 1366 581 1367
rect 602 1367 608 1368
rect 602 1366 603 1367
rect 580 1364 603 1366
rect 580 1363 581 1364
rect 575 1362 581 1363
rect 602 1363 603 1364
rect 607 1363 608 1367
rect 602 1362 608 1363
rect 610 1367 616 1368
rect 610 1363 611 1367
rect 615 1366 616 1367
rect 663 1367 669 1368
rect 663 1366 664 1367
rect 615 1364 664 1366
rect 615 1363 616 1364
rect 610 1362 616 1363
rect 663 1363 664 1364
rect 668 1363 669 1367
rect 663 1362 669 1363
rect 751 1367 757 1368
rect 751 1363 752 1367
rect 756 1366 757 1367
rect 786 1367 792 1368
rect 786 1366 787 1367
rect 756 1364 787 1366
rect 756 1363 757 1364
rect 751 1362 757 1363
rect 786 1363 787 1364
rect 791 1363 792 1367
rect 786 1362 792 1363
rect 839 1367 845 1368
rect 839 1363 840 1367
rect 844 1366 845 1367
rect 870 1367 876 1368
rect 870 1366 871 1367
rect 844 1364 871 1366
rect 844 1363 845 1364
rect 839 1362 845 1363
rect 870 1363 871 1364
rect 875 1363 876 1367
rect 870 1362 876 1363
rect 914 1367 920 1368
rect 914 1363 915 1367
rect 919 1366 920 1367
rect 951 1367 957 1368
rect 951 1366 952 1367
rect 919 1364 952 1366
rect 919 1363 920 1364
rect 914 1362 920 1363
rect 951 1363 952 1364
rect 956 1363 957 1367
rect 951 1362 957 1363
rect 1079 1367 1085 1368
rect 1079 1363 1080 1367
rect 1084 1366 1085 1367
rect 1114 1367 1120 1368
rect 1114 1366 1115 1367
rect 1084 1364 1115 1366
rect 1084 1363 1085 1364
rect 1079 1362 1085 1363
rect 1114 1363 1115 1364
rect 1119 1363 1120 1367
rect 1114 1362 1120 1363
rect 1239 1367 1248 1368
rect 1239 1363 1240 1367
rect 1247 1363 1248 1367
rect 1239 1362 1248 1363
rect 1370 1367 1376 1368
rect 1370 1363 1371 1367
rect 1375 1366 1376 1367
rect 1415 1367 1421 1368
rect 1415 1366 1416 1367
rect 1375 1364 1416 1366
rect 1375 1363 1376 1364
rect 1370 1362 1376 1363
rect 1415 1363 1416 1364
rect 1420 1363 1421 1367
rect 1415 1362 1421 1363
rect 1502 1367 1508 1368
rect 1502 1363 1503 1367
rect 1507 1366 1508 1367
rect 1607 1367 1613 1368
rect 1607 1366 1608 1367
rect 1507 1364 1608 1366
rect 1507 1363 1508 1364
rect 1502 1362 1508 1363
rect 1607 1363 1608 1364
rect 1612 1363 1613 1367
rect 1607 1362 1613 1363
rect 1774 1367 1781 1368
rect 1774 1363 1775 1367
rect 1780 1363 1781 1367
rect 1774 1362 1781 1363
rect 1902 1362 1908 1363
rect 1902 1358 1903 1362
rect 1907 1358 1908 1362
rect 1902 1357 1908 1358
rect 2030 1362 2036 1363
rect 2030 1358 2031 1362
rect 2035 1358 2036 1362
rect 2030 1357 2036 1358
rect 2174 1362 2180 1363
rect 2174 1358 2175 1362
rect 2179 1358 2180 1362
rect 2174 1357 2180 1358
rect 2310 1362 2316 1363
rect 2310 1358 2311 1362
rect 2315 1358 2316 1362
rect 2310 1357 2316 1358
rect 2438 1362 2444 1363
rect 2438 1358 2439 1362
rect 2443 1358 2444 1362
rect 2438 1357 2444 1358
rect 2558 1362 2564 1363
rect 2558 1358 2559 1362
rect 2563 1358 2564 1362
rect 2558 1357 2564 1358
rect 2678 1362 2684 1363
rect 2678 1358 2679 1362
rect 2683 1358 2684 1362
rect 2678 1357 2684 1358
rect 2798 1362 2804 1363
rect 2798 1358 2799 1362
rect 2803 1358 2804 1362
rect 2798 1357 2804 1358
rect 2918 1362 2924 1363
rect 2918 1358 2919 1362
rect 2923 1358 2924 1362
rect 2918 1357 2924 1358
rect 314 1355 320 1356
rect 314 1351 315 1355
rect 319 1354 320 1355
rect 383 1355 389 1356
rect 383 1354 384 1355
rect 319 1352 384 1354
rect 319 1351 320 1352
rect 314 1350 320 1351
rect 383 1351 384 1352
rect 388 1351 389 1355
rect 383 1350 389 1351
rect 410 1355 416 1356
rect 410 1351 411 1355
rect 415 1354 416 1355
rect 495 1355 501 1356
rect 495 1354 496 1355
rect 415 1352 496 1354
rect 415 1351 416 1352
rect 410 1350 416 1351
rect 495 1351 496 1352
rect 500 1351 501 1355
rect 495 1350 501 1351
rect 522 1355 528 1356
rect 522 1351 523 1355
rect 527 1354 528 1355
rect 615 1355 621 1356
rect 615 1354 616 1355
rect 527 1352 616 1354
rect 527 1351 528 1352
rect 522 1350 528 1351
rect 615 1351 616 1352
rect 620 1351 621 1355
rect 615 1350 621 1351
rect 718 1355 724 1356
rect 718 1351 719 1355
rect 723 1354 724 1355
rect 751 1355 757 1356
rect 751 1354 752 1355
rect 723 1352 752 1354
rect 723 1351 724 1352
rect 718 1350 724 1351
rect 751 1351 752 1352
rect 756 1351 757 1355
rect 751 1350 757 1351
rect 887 1355 893 1356
rect 887 1351 888 1355
rect 892 1354 893 1355
rect 1014 1355 1020 1356
rect 1014 1354 1015 1355
rect 892 1352 1015 1354
rect 892 1351 893 1352
rect 887 1350 893 1351
rect 1014 1351 1015 1352
rect 1019 1351 1020 1355
rect 1014 1350 1020 1351
rect 1031 1355 1037 1356
rect 1031 1351 1032 1355
rect 1036 1354 1037 1355
rect 1150 1355 1156 1356
rect 1150 1354 1151 1355
rect 1036 1352 1151 1354
rect 1036 1351 1037 1352
rect 1031 1350 1037 1351
rect 1150 1351 1151 1352
rect 1155 1351 1156 1355
rect 1150 1350 1156 1351
rect 1167 1355 1176 1356
rect 1167 1351 1168 1355
rect 1175 1351 1176 1355
rect 1167 1350 1176 1351
rect 1303 1355 1312 1356
rect 1303 1351 1304 1355
rect 1311 1351 1312 1355
rect 1303 1350 1312 1351
rect 1330 1355 1336 1356
rect 1330 1351 1331 1355
rect 1335 1354 1336 1355
rect 1431 1355 1437 1356
rect 1431 1354 1432 1355
rect 1335 1352 1432 1354
rect 1335 1351 1336 1352
rect 1330 1350 1336 1351
rect 1431 1351 1432 1352
rect 1436 1351 1437 1355
rect 1431 1350 1437 1351
rect 1458 1355 1464 1356
rect 1458 1351 1459 1355
rect 1463 1354 1464 1355
rect 1551 1355 1557 1356
rect 1551 1354 1552 1355
rect 1463 1352 1552 1354
rect 1463 1351 1464 1352
rect 1458 1350 1464 1351
rect 1551 1351 1552 1352
rect 1556 1351 1557 1355
rect 1551 1350 1557 1351
rect 1615 1355 1621 1356
rect 1615 1351 1616 1355
rect 1620 1354 1621 1355
rect 1671 1355 1677 1356
rect 1671 1354 1672 1355
rect 1620 1352 1672 1354
rect 1620 1351 1621 1352
rect 1615 1350 1621 1351
rect 1671 1351 1672 1352
rect 1676 1351 1677 1355
rect 1671 1350 1677 1351
rect 1698 1355 1704 1356
rect 1698 1351 1699 1355
rect 1703 1354 1704 1355
rect 1775 1355 1781 1356
rect 1775 1354 1776 1355
rect 1703 1352 1776 1354
rect 1703 1351 1704 1352
rect 1698 1350 1704 1351
rect 1775 1351 1776 1352
rect 1780 1351 1781 1355
rect 1775 1350 1781 1351
rect 1810 1351 1816 1352
rect 1810 1347 1811 1351
rect 1815 1350 1816 1351
rect 1927 1351 1933 1352
rect 1927 1350 1928 1351
rect 1815 1348 1928 1350
rect 1815 1347 1816 1348
rect 358 1346 364 1347
rect 358 1342 359 1346
rect 363 1342 364 1346
rect 358 1341 364 1342
rect 470 1346 476 1347
rect 470 1342 471 1346
rect 475 1342 476 1346
rect 470 1341 476 1342
rect 590 1346 596 1347
rect 590 1342 591 1346
rect 595 1342 596 1346
rect 590 1341 596 1342
rect 726 1346 732 1347
rect 726 1342 727 1346
rect 731 1342 732 1346
rect 726 1341 732 1342
rect 862 1346 868 1347
rect 862 1342 863 1346
rect 867 1342 868 1346
rect 862 1341 868 1342
rect 1006 1346 1012 1347
rect 1006 1342 1007 1346
rect 1011 1342 1012 1346
rect 1006 1341 1012 1342
rect 1142 1346 1148 1347
rect 1142 1342 1143 1346
rect 1147 1342 1148 1346
rect 1142 1341 1148 1342
rect 1278 1346 1284 1347
rect 1278 1342 1279 1346
rect 1283 1342 1284 1346
rect 1278 1341 1284 1342
rect 1406 1346 1412 1347
rect 1406 1342 1407 1346
rect 1411 1342 1412 1346
rect 1406 1341 1412 1342
rect 1526 1346 1532 1347
rect 1526 1342 1527 1346
rect 1531 1342 1532 1346
rect 1526 1341 1532 1342
rect 1646 1346 1652 1347
rect 1646 1342 1647 1346
rect 1651 1342 1652 1346
rect 1646 1341 1652 1342
rect 1750 1346 1756 1347
rect 1810 1346 1816 1347
rect 1927 1347 1928 1348
rect 1932 1347 1933 1351
rect 1927 1346 1933 1347
rect 2055 1351 2064 1352
rect 2055 1347 2056 1351
rect 2063 1347 2064 1351
rect 2055 1346 2064 1347
rect 2114 1351 2120 1352
rect 2114 1347 2115 1351
rect 2119 1350 2120 1351
rect 2199 1351 2205 1352
rect 2199 1350 2200 1351
rect 2119 1348 2200 1350
rect 2119 1347 2120 1348
rect 2114 1346 2120 1347
rect 2199 1347 2200 1348
rect 2204 1347 2205 1351
rect 2199 1346 2205 1347
rect 2258 1351 2264 1352
rect 2258 1347 2259 1351
rect 2263 1350 2264 1351
rect 2335 1351 2341 1352
rect 2335 1350 2336 1351
rect 2263 1348 2336 1350
rect 2263 1347 2264 1348
rect 2258 1346 2264 1347
rect 2335 1347 2336 1348
rect 2340 1347 2341 1351
rect 2335 1346 2341 1347
rect 2463 1351 2472 1352
rect 2463 1347 2464 1351
rect 2471 1347 2472 1351
rect 2463 1346 2472 1347
rect 2514 1351 2520 1352
rect 2514 1347 2515 1351
rect 2519 1350 2520 1351
rect 2583 1351 2589 1352
rect 2583 1350 2584 1351
rect 2519 1348 2584 1350
rect 2519 1347 2520 1348
rect 2514 1346 2520 1347
rect 2583 1347 2584 1348
rect 2588 1347 2589 1351
rect 2583 1346 2589 1347
rect 2634 1351 2640 1352
rect 2634 1347 2635 1351
rect 2639 1350 2640 1351
rect 2703 1351 2709 1352
rect 2703 1350 2704 1351
rect 2639 1348 2704 1350
rect 2639 1347 2640 1348
rect 2634 1346 2640 1347
rect 2703 1347 2704 1348
rect 2708 1347 2709 1351
rect 2703 1346 2709 1347
rect 2754 1351 2760 1352
rect 2754 1347 2755 1351
rect 2759 1350 2760 1351
rect 2823 1351 2829 1352
rect 2823 1350 2824 1351
rect 2759 1348 2824 1350
rect 2759 1347 2760 1348
rect 2754 1346 2760 1347
rect 2823 1347 2824 1348
rect 2828 1347 2829 1351
rect 2823 1346 2829 1347
rect 2866 1351 2872 1352
rect 2866 1347 2867 1351
rect 2871 1350 2872 1351
rect 2943 1351 2949 1352
rect 2943 1350 2944 1351
rect 2871 1348 2944 1350
rect 2871 1347 2872 1348
rect 2866 1346 2872 1347
rect 2943 1347 2944 1348
rect 2948 1347 2949 1351
rect 2943 1346 2949 1347
rect 1750 1342 1751 1346
rect 1755 1342 1756 1346
rect 1750 1341 1756 1342
rect 2378 1339 2384 1340
rect 2378 1335 2379 1339
rect 2383 1338 2384 1339
rect 2383 1336 2474 1338
rect 2383 1335 2384 1336
rect 2378 1334 2384 1335
rect 1951 1331 1957 1332
rect 110 1328 116 1329
rect 110 1324 111 1328
rect 115 1324 116 1328
rect 110 1323 116 1324
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1951 1327 1952 1331
rect 1956 1330 1957 1331
rect 1978 1331 1984 1332
rect 1956 1328 1974 1330
rect 1956 1327 1957 1328
rect 1951 1326 1957 1327
rect 1830 1323 1836 1324
rect 1926 1322 1932 1323
rect 410 1319 416 1320
rect 410 1315 411 1319
rect 415 1315 416 1319
rect 410 1314 416 1315
rect 522 1319 528 1320
rect 522 1315 523 1319
rect 527 1315 528 1319
rect 718 1319 724 1320
rect 718 1318 719 1319
rect 645 1316 719 1318
rect 522 1314 528 1315
rect 718 1315 719 1316
rect 723 1315 724 1319
rect 718 1314 724 1315
rect 914 1319 920 1320
rect 914 1315 915 1319
rect 919 1315 920 1319
rect 914 1314 920 1315
rect 1014 1319 1020 1320
rect 1014 1315 1015 1319
rect 1019 1315 1020 1319
rect 1014 1314 1020 1315
rect 1150 1319 1156 1320
rect 1150 1315 1151 1319
rect 1155 1315 1156 1319
rect 1150 1314 1156 1315
rect 1330 1319 1336 1320
rect 1330 1315 1331 1319
rect 1335 1315 1336 1319
rect 1330 1314 1336 1315
rect 1458 1319 1464 1320
rect 1458 1315 1459 1319
rect 1463 1315 1464 1319
rect 1615 1319 1621 1320
rect 1615 1318 1616 1319
rect 1581 1316 1616 1318
rect 1458 1314 1464 1315
rect 1615 1315 1616 1316
rect 1620 1315 1621 1319
rect 1615 1314 1621 1315
rect 1698 1319 1704 1320
rect 1698 1315 1699 1319
rect 1703 1315 1704 1319
rect 1698 1314 1704 1315
rect 1774 1319 1780 1320
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1926 1318 1927 1322
rect 1931 1318 1932 1322
rect 1972 1322 1974 1328
rect 1978 1327 1979 1331
rect 1983 1330 1984 1331
rect 2071 1331 2077 1332
rect 2071 1330 2072 1331
rect 1983 1328 2072 1330
rect 1983 1327 1984 1328
rect 1978 1326 1984 1327
rect 2071 1327 2072 1328
rect 2076 1327 2077 1331
rect 2071 1326 2077 1327
rect 2098 1331 2104 1332
rect 2098 1327 2099 1331
rect 2103 1330 2104 1331
rect 2207 1331 2213 1332
rect 2207 1330 2208 1331
rect 2103 1328 2208 1330
rect 2103 1327 2104 1328
rect 2098 1326 2104 1327
rect 2207 1327 2208 1328
rect 2212 1327 2213 1331
rect 2207 1326 2213 1327
rect 2343 1331 2349 1332
rect 2343 1327 2344 1331
rect 2348 1330 2349 1331
rect 2462 1331 2468 1332
rect 2462 1330 2463 1331
rect 2348 1328 2463 1330
rect 2348 1327 2349 1328
rect 2343 1326 2349 1327
rect 2462 1327 2463 1328
rect 2467 1327 2468 1331
rect 2472 1330 2474 1336
rect 2479 1331 2485 1332
rect 2479 1330 2480 1331
rect 2472 1328 2480 1330
rect 2462 1326 2468 1327
rect 2479 1327 2480 1328
rect 2484 1327 2485 1331
rect 2479 1326 2485 1327
rect 2615 1331 2624 1332
rect 2615 1327 2616 1331
rect 2623 1327 2624 1331
rect 2615 1326 2624 1327
rect 2642 1331 2648 1332
rect 2642 1327 2643 1331
rect 2647 1330 2648 1331
rect 2743 1331 2749 1332
rect 2743 1330 2744 1331
rect 2647 1328 2744 1330
rect 2647 1327 2648 1328
rect 2642 1326 2648 1327
rect 2743 1327 2744 1328
rect 2748 1327 2749 1331
rect 2743 1326 2749 1327
rect 2770 1331 2776 1332
rect 2770 1327 2771 1331
rect 2775 1330 2776 1331
rect 2863 1331 2869 1332
rect 2863 1330 2864 1331
rect 2775 1328 2864 1330
rect 2775 1327 2776 1328
rect 2770 1326 2776 1327
rect 2863 1327 2864 1328
rect 2868 1327 2869 1331
rect 2863 1326 2869 1327
rect 2890 1331 2896 1332
rect 2890 1327 2891 1331
rect 2895 1330 2896 1331
rect 2975 1331 2981 1332
rect 2975 1330 2976 1331
rect 2895 1328 2976 1330
rect 2895 1327 2896 1328
rect 2890 1326 2896 1327
rect 2975 1327 2976 1328
rect 2980 1327 2981 1331
rect 2975 1326 2981 1327
rect 3002 1331 3008 1332
rect 3002 1327 3003 1331
rect 3007 1330 3008 1331
rect 3087 1331 3093 1332
rect 3087 1330 3088 1331
rect 3007 1328 3088 1330
rect 3007 1327 3008 1328
rect 3002 1326 3008 1327
rect 3087 1327 3088 1328
rect 3092 1327 3093 1331
rect 3087 1326 3093 1327
rect 3114 1331 3120 1332
rect 3114 1327 3115 1331
rect 3119 1330 3120 1331
rect 3207 1331 3213 1332
rect 3207 1330 3208 1331
rect 3119 1328 3208 1330
rect 3119 1327 3120 1328
rect 3114 1326 3120 1327
rect 3207 1327 3208 1328
rect 3212 1327 3213 1331
rect 3207 1326 3213 1327
rect 1986 1323 1992 1324
rect 1986 1322 1987 1323
rect 1972 1320 1987 1322
rect 1986 1319 1987 1320
rect 1991 1319 1992 1323
rect 1986 1318 1992 1319
rect 2046 1322 2052 1323
rect 2046 1318 2047 1322
rect 2051 1318 2052 1322
rect 1926 1317 1932 1318
rect 2046 1317 2052 1318
rect 2182 1322 2188 1323
rect 2182 1318 2183 1322
rect 2187 1318 2188 1322
rect 2182 1317 2188 1318
rect 2318 1322 2324 1323
rect 2318 1318 2319 1322
rect 2323 1318 2324 1322
rect 2318 1317 2324 1318
rect 2454 1322 2460 1323
rect 2454 1318 2455 1322
rect 2459 1318 2460 1322
rect 2454 1317 2460 1318
rect 2590 1322 2596 1323
rect 2590 1318 2591 1322
rect 2595 1318 2596 1322
rect 2590 1317 2596 1318
rect 2718 1322 2724 1323
rect 2718 1318 2719 1322
rect 2723 1318 2724 1322
rect 2718 1317 2724 1318
rect 2838 1322 2844 1323
rect 2838 1318 2839 1322
rect 2843 1318 2844 1322
rect 2838 1317 2844 1318
rect 2950 1322 2956 1323
rect 2950 1318 2951 1322
rect 2955 1318 2956 1322
rect 2950 1317 2956 1318
rect 3062 1322 3068 1323
rect 3062 1318 3063 1322
rect 3067 1318 3068 1322
rect 3062 1317 3068 1318
rect 3182 1322 3188 1323
rect 3182 1318 3183 1322
rect 3187 1318 3188 1322
rect 3182 1317 3188 1318
rect 1774 1314 1780 1315
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 1830 1311 1836 1312
rect 110 1306 116 1307
rect 350 1308 356 1309
rect 350 1304 351 1308
rect 355 1304 356 1308
rect 350 1303 356 1304
rect 462 1308 468 1309
rect 462 1304 463 1308
rect 467 1304 468 1308
rect 462 1303 468 1304
rect 582 1308 588 1309
rect 582 1304 583 1308
rect 587 1304 588 1308
rect 582 1303 588 1304
rect 718 1308 724 1309
rect 718 1304 719 1308
rect 723 1304 724 1308
rect 718 1303 724 1304
rect 854 1308 860 1309
rect 854 1304 855 1308
rect 859 1304 860 1308
rect 854 1303 860 1304
rect 998 1308 1004 1309
rect 998 1304 999 1308
rect 1003 1304 1004 1308
rect 998 1303 1004 1304
rect 1134 1308 1140 1309
rect 1134 1304 1135 1308
rect 1139 1304 1140 1308
rect 1134 1303 1140 1304
rect 1270 1308 1276 1309
rect 1270 1304 1271 1308
rect 1275 1304 1276 1308
rect 1270 1303 1276 1304
rect 1398 1308 1404 1309
rect 1398 1304 1399 1308
rect 1403 1304 1404 1308
rect 1398 1303 1404 1304
rect 1518 1308 1524 1309
rect 1518 1304 1519 1308
rect 1523 1304 1524 1308
rect 1518 1303 1524 1304
rect 1638 1308 1644 1309
rect 1638 1304 1639 1308
rect 1643 1304 1644 1308
rect 1638 1303 1644 1304
rect 1742 1308 1748 1309
rect 1742 1304 1743 1308
rect 1747 1304 1748 1308
rect 1830 1307 1831 1311
rect 1835 1307 1836 1311
rect 1830 1306 1836 1307
rect 1742 1303 1748 1304
rect 1870 1304 1876 1305
rect 1870 1300 1871 1304
rect 1875 1300 1876 1304
rect 1870 1299 1876 1300
rect 3590 1304 3596 1305
rect 3590 1300 3591 1304
rect 3595 1300 3596 1304
rect 3590 1299 3596 1300
rect 1978 1295 1984 1296
rect 706 1291 712 1292
rect 706 1287 707 1291
rect 711 1290 712 1291
rect 735 1291 741 1292
rect 735 1290 736 1291
rect 711 1288 736 1290
rect 711 1287 712 1288
rect 706 1286 712 1287
rect 735 1287 736 1288
rect 740 1287 741 1291
rect 1978 1291 1979 1295
rect 1983 1291 1984 1295
rect 1978 1290 1984 1291
rect 2098 1295 2104 1296
rect 2098 1291 2099 1295
rect 2103 1291 2104 1295
rect 2098 1290 2104 1291
rect 2234 1295 2240 1296
rect 2234 1291 2235 1295
rect 2239 1291 2240 1295
rect 2234 1290 2240 1291
rect 2326 1295 2332 1296
rect 2326 1291 2327 1295
rect 2331 1291 2332 1295
rect 2326 1290 2332 1291
rect 2462 1295 2468 1296
rect 2462 1291 2463 1295
rect 2467 1291 2468 1295
rect 2462 1290 2468 1291
rect 2642 1295 2648 1296
rect 2642 1291 2643 1295
rect 2647 1291 2648 1295
rect 2642 1290 2648 1291
rect 2770 1295 2776 1296
rect 2770 1291 2771 1295
rect 2775 1291 2776 1295
rect 2770 1290 2776 1291
rect 2890 1295 2896 1296
rect 2890 1291 2891 1295
rect 2895 1291 2896 1295
rect 2890 1290 2896 1291
rect 3002 1295 3008 1296
rect 3002 1291 3003 1295
rect 3007 1291 3008 1295
rect 3002 1290 3008 1291
rect 3114 1295 3120 1296
rect 3114 1291 3115 1295
rect 3119 1291 3120 1295
rect 3114 1290 3120 1291
rect 735 1286 741 1287
rect 1870 1287 1876 1288
rect 1870 1283 1871 1287
rect 1875 1283 1876 1287
rect 3590 1287 3596 1288
rect 1870 1282 1876 1283
rect 1918 1284 1924 1285
rect 1918 1280 1919 1284
rect 1923 1280 1924 1284
rect 1918 1279 1924 1280
rect 2038 1284 2044 1285
rect 2038 1280 2039 1284
rect 2043 1280 2044 1284
rect 2038 1279 2044 1280
rect 2174 1284 2180 1285
rect 2174 1280 2175 1284
rect 2179 1280 2180 1284
rect 2174 1279 2180 1280
rect 2310 1284 2316 1285
rect 2310 1280 2311 1284
rect 2315 1280 2316 1284
rect 2310 1279 2316 1280
rect 2446 1284 2452 1285
rect 2446 1280 2447 1284
rect 2451 1280 2452 1284
rect 2446 1279 2452 1280
rect 2582 1284 2588 1285
rect 2582 1280 2583 1284
rect 2587 1280 2588 1284
rect 2582 1279 2588 1280
rect 2710 1284 2716 1285
rect 2710 1280 2711 1284
rect 2715 1280 2716 1284
rect 2710 1279 2716 1280
rect 2830 1284 2836 1285
rect 2830 1280 2831 1284
rect 2835 1280 2836 1284
rect 2830 1279 2836 1280
rect 2942 1284 2948 1285
rect 2942 1280 2943 1284
rect 2947 1280 2948 1284
rect 2942 1279 2948 1280
rect 3054 1284 3060 1285
rect 3054 1280 3055 1284
rect 3059 1280 3060 1284
rect 3054 1279 3060 1280
rect 3174 1284 3180 1285
rect 3174 1280 3175 1284
rect 3179 1280 3180 1284
rect 3590 1283 3591 1287
rect 3595 1283 3596 1287
rect 3590 1282 3596 1283
rect 3174 1279 3180 1280
rect 3062 1267 3068 1268
rect 3062 1263 3063 1267
rect 3067 1266 3068 1267
rect 3191 1267 3197 1268
rect 3191 1266 3192 1267
rect 3067 1264 3192 1266
rect 3067 1263 3068 1264
rect 3062 1262 3068 1263
rect 3191 1263 3192 1264
rect 3196 1263 3197 1267
rect 3191 1262 3197 1263
rect 310 1260 316 1261
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 310 1256 311 1260
rect 315 1256 316 1260
rect 310 1255 316 1256
rect 414 1260 420 1261
rect 414 1256 415 1260
rect 419 1256 420 1260
rect 414 1255 420 1256
rect 534 1260 540 1261
rect 534 1256 535 1260
rect 539 1256 540 1260
rect 534 1255 540 1256
rect 670 1260 676 1261
rect 670 1256 671 1260
rect 675 1256 676 1260
rect 670 1255 676 1256
rect 814 1260 820 1261
rect 814 1256 815 1260
rect 819 1256 820 1260
rect 814 1255 820 1256
rect 958 1260 964 1261
rect 958 1256 959 1260
rect 963 1256 964 1260
rect 958 1255 964 1256
rect 1102 1260 1108 1261
rect 1102 1256 1103 1260
rect 1107 1256 1108 1260
rect 1102 1255 1108 1256
rect 1238 1260 1244 1261
rect 1238 1256 1239 1260
rect 1243 1256 1244 1260
rect 1238 1255 1244 1256
rect 1374 1260 1380 1261
rect 1374 1256 1375 1260
rect 1379 1256 1380 1260
rect 1374 1255 1380 1256
rect 1502 1260 1508 1261
rect 1502 1256 1503 1260
rect 1507 1256 1508 1260
rect 1502 1255 1508 1256
rect 1630 1260 1636 1261
rect 1630 1256 1631 1260
rect 1635 1256 1636 1260
rect 1630 1255 1636 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1742 1255 1748 1256
rect 1830 1257 1836 1258
rect 110 1252 116 1253
rect 1830 1253 1831 1257
rect 1835 1253 1836 1257
rect 1830 1252 1836 1253
rect 266 1251 272 1252
rect 266 1247 267 1251
rect 271 1250 272 1251
rect 378 1251 384 1252
rect 271 1248 329 1250
rect 271 1247 272 1248
rect 266 1246 272 1247
rect 378 1247 379 1251
rect 383 1250 384 1251
rect 482 1251 488 1252
rect 383 1248 433 1250
rect 383 1247 384 1248
rect 378 1246 384 1247
rect 482 1247 483 1251
rect 487 1250 488 1251
rect 602 1251 608 1252
rect 487 1248 553 1250
rect 487 1247 488 1248
rect 482 1246 488 1247
rect 602 1247 603 1251
rect 607 1250 608 1251
rect 906 1251 912 1252
rect 906 1250 907 1251
rect 607 1248 689 1250
rect 877 1248 907 1250
rect 607 1247 608 1248
rect 602 1246 608 1247
rect 906 1247 907 1248
rect 911 1247 912 1251
rect 1050 1251 1056 1252
rect 1050 1250 1051 1251
rect 1021 1248 1051 1250
rect 906 1246 912 1247
rect 1050 1247 1051 1248
rect 1055 1247 1056 1251
rect 1170 1251 1176 1252
rect 1170 1250 1171 1251
rect 1165 1248 1171 1250
rect 1050 1246 1056 1247
rect 1170 1247 1171 1248
rect 1175 1247 1176 1251
rect 1330 1251 1336 1252
rect 1330 1250 1331 1251
rect 1301 1248 1331 1250
rect 1170 1246 1176 1247
rect 1330 1247 1331 1248
rect 1335 1247 1336 1251
rect 1462 1251 1468 1252
rect 1462 1250 1463 1251
rect 1437 1248 1463 1250
rect 1330 1246 1336 1247
rect 1462 1247 1463 1248
rect 1467 1247 1468 1251
rect 1590 1251 1596 1252
rect 1590 1250 1591 1251
rect 1565 1248 1591 1250
rect 1462 1246 1468 1247
rect 1590 1247 1591 1248
rect 1595 1247 1596 1251
rect 1590 1246 1596 1247
rect 1598 1251 1604 1252
rect 1598 1247 1599 1251
rect 1603 1250 1604 1251
rect 1603 1248 1649 1250
rect 1603 1247 1604 1248
rect 1598 1246 1604 1247
rect 1804 1244 1806 1249
rect 1802 1243 1808 1244
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 1802 1239 1803 1243
rect 1807 1239 1808 1243
rect 1802 1238 1808 1239
rect 1830 1240 1836 1241
rect 110 1235 116 1236
rect 1830 1236 1831 1240
rect 1835 1236 1836 1240
rect 1830 1235 1836 1236
rect 1894 1232 1900 1233
rect 1870 1229 1876 1230
rect 1870 1225 1871 1229
rect 1875 1225 1876 1229
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 1894 1227 1900 1228
rect 2070 1232 2076 1233
rect 2070 1228 2071 1232
rect 2075 1228 2076 1232
rect 2070 1227 2076 1228
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2470 1232 2476 1233
rect 2470 1228 2471 1232
rect 2475 1228 2476 1232
rect 2470 1227 2476 1228
rect 2662 1232 2668 1233
rect 2662 1228 2663 1232
rect 2667 1228 2668 1232
rect 2662 1227 2668 1228
rect 2846 1232 2852 1233
rect 2846 1228 2847 1232
rect 2851 1228 2852 1232
rect 2846 1227 2852 1228
rect 3022 1232 3028 1233
rect 3022 1228 3023 1232
rect 3027 1228 3028 1232
rect 3022 1227 3028 1228
rect 3190 1232 3196 1233
rect 3190 1228 3191 1232
rect 3195 1228 3196 1232
rect 3190 1227 3196 1228
rect 3358 1232 3364 1233
rect 3358 1228 3359 1232
rect 3363 1228 3364 1232
rect 3358 1227 3364 1228
rect 3502 1232 3508 1233
rect 3502 1228 3503 1232
rect 3507 1228 3508 1232
rect 3502 1227 3508 1228
rect 3590 1229 3596 1230
rect 1870 1224 1876 1225
rect 3590 1225 3591 1229
rect 3595 1225 3596 1229
rect 3590 1224 3596 1225
rect 2138 1223 2144 1224
rect 318 1222 324 1223
rect 318 1218 319 1222
rect 323 1218 324 1222
rect 318 1217 324 1218
rect 422 1222 428 1223
rect 422 1218 423 1222
rect 427 1218 428 1222
rect 422 1217 428 1218
rect 542 1222 548 1223
rect 542 1218 543 1222
rect 547 1218 548 1222
rect 542 1217 548 1218
rect 678 1222 684 1223
rect 678 1218 679 1222
rect 683 1218 684 1222
rect 678 1217 684 1218
rect 822 1222 828 1223
rect 822 1218 823 1222
rect 827 1218 828 1222
rect 822 1217 828 1218
rect 966 1222 972 1223
rect 966 1218 967 1222
rect 971 1218 972 1222
rect 966 1217 972 1218
rect 1110 1222 1116 1223
rect 1110 1218 1111 1222
rect 1115 1218 1116 1222
rect 1110 1217 1116 1218
rect 1246 1222 1252 1223
rect 1246 1218 1247 1222
rect 1251 1218 1252 1222
rect 1246 1217 1252 1218
rect 1382 1222 1388 1223
rect 1382 1218 1383 1222
rect 1387 1218 1388 1222
rect 1382 1217 1388 1218
rect 1510 1222 1516 1223
rect 1510 1218 1511 1222
rect 1515 1218 1516 1222
rect 1510 1217 1516 1218
rect 1638 1222 1644 1223
rect 1638 1218 1639 1222
rect 1643 1218 1644 1222
rect 1638 1217 1644 1218
rect 1750 1222 1756 1223
rect 1750 1218 1751 1222
rect 1755 1218 1756 1222
rect 1750 1217 1756 1218
rect 1956 1216 1958 1221
rect 1964 1220 2089 1222
rect 1954 1215 1960 1216
rect 1870 1212 1876 1213
rect 343 1211 349 1212
rect 343 1207 344 1211
rect 348 1210 349 1211
rect 378 1211 384 1212
rect 378 1210 379 1211
rect 348 1208 379 1210
rect 348 1207 349 1208
rect 343 1206 349 1207
rect 378 1207 379 1208
rect 383 1207 384 1211
rect 378 1206 384 1207
rect 447 1211 453 1212
rect 447 1207 448 1211
rect 452 1210 453 1211
rect 482 1211 488 1212
rect 482 1210 483 1211
rect 452 1208 483 1210
rect 452 1207 453 1208
rect 447 1206 453 1207
rect 482 1207 483 1208
rect 487 1207 488 1211
rect 482 1206 488 1207
rect 567 1211 573 1212
rect 567 1207 568 1211
rect 572 1210 573 1211
rect 602 1211 608 1212
rect 602 1210 603 1211
rect 572 1208 603 1210
rect 572 1207 573 1208
rect 567 1206 573 1207
rect 602 1207 603 1208
rect 607 1207 608 1211
rect 602 1206 608 1207
rect 703 1211 712 1212
rect 703 1207 704 1211
rect 711 1207 712 1211
rect 703 1206 712 1207
rect 810 1211 816 1212
rect 810 1207 811 1211
rect 815 1210 816 1211
rect 847 1211 853 1212
rect 847 1210 848 1211
rect 815 1208 848 1210
rect 815 1207 816 1208
rect 810 1206 816 1207
rect 847 1207 848 1208
rect 852 1207 853 1211
rect 847 1206 853 1207
rect 906 1211 912 1212
rect 906 1207 907 1211
rect 911 1210 912 1211
rect 991 1211 997 1212
rect 991 1210 992 1211
rect 911 1208 992 1210
rect 911 1207 912 1208
rect 906 1206 912 1207
rect 991 1207 992 1208
rect 996 1207 997 1211
rect 991 1206 997 1207
rect 1050 1211 1056 1212
rect 1050 1207 1051 1211
rect 1055 1210 1056 1211
rect 1135 1211 1141 1212
rect 1135 1210 1136 1211
rect 1055 1208 1136 1210
rect 1055 1207 1056 1208
rect 1050 1206 1056 1207
rect 1135 1207 1136 1208
rect 1140 1207 1141 1211
rect 1135 1206 1141 1207
rect 1271 1211 1277 1212
rect 1271 1207 1272 1211
rect 1276 1210 1277 1211
rect 1287 1211 1293 1212
rect 1287 1210 1288 1211
rect 1276 1208 1288 1210
rect 1276 1207 1277 1208
rect 1271 1206 1277 1207
rect 1287 1207 1288 1208
rect 1292 1207 1293 1211
rect 1287 1206 1293 1207
rect 1330 1211 1336 1212
rect 1330 1207 1331 1211
rect 1335 1210 1336 1211
rect 1407 1211 1413 1212
rect 1407 1210 1408 1211
rect 1335 1208 1408 1210
rect 1335 1207 1336 1208
rect 1330 1206 1336 1207
rect 1407 1207 1408 1208
rect 1412 1207 1413 1211
rect 1407 1206 1413 1207
rect 1462 1211 1468 1212
rect 1462 1207 1463 1211
rect 1467 1210 1468 1211
rect 1535 1211 1541 1212
rect 1535 1210 1536 1211
rect 1467 1208 1536 1210
rect 1467 1207 1468 1208
rect 1462 1206 1468 1207
rect 1535 1207 1536 1208
rect 1540 1207 1541 1211
rect 1535 1206 1541 1207
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1210 1596 1211
rect 1663 1211 1669 1212
rect 1663 1210 1664 1211
rect 1595 1208 1664 1210
rect 1595 1207 1596 1208
rect 1590 1206 1596 1207
rect 1663 1207 1664 1208
rect 1668 1207 1669 1211
rect 1663 1206 1669 1207
rect 1775 1211 1781 1212
rect 1775 1207 1776 1211
rect 1780 1210 1781 1211
rect 1780 1208 1866 1210
rect 1780 1207 1781 1208
rect 1775 1206 1781 1207
rect 1864 1202 1866 1208
rect 1870 1208 1871 1212
rect 1875 1208 1876 1212
rect 1954 1211 1955 1215
rect 1959 1211 1960 1215
rect 1954 1210 1960 1211
rect 1870 1207 1876 1208
rect 1964 1202 1966 1220
rect 2138 1219 2139 1223
rect 2143 1222 2144 1223
rect 2590 1223 2596 1224
rect 2590 1222 2591 1223
rect 2143 1220 2289 1222
rect 2533 1220 2591 1222
rect 2143 1219 2144 1220
rect 2138 1218 2144 1219
rect 2590 1219 2591 1220
rect 2595 1219 2596 1223
rect 2778 1223 2784 1224
rect 2590 1218 2596 1219
rect 2724 1216 2726 1221
rect 2778 1219 2779 1223
rect 2783 1222 2784 1223
rect 2914 1223 2920 1224
rect 2783 1220 2865 1222
rect 2783 1219 2784 1220
rect 2778 1218 2784 1219
rect 2914 1219 2915 1223
rect 2919 1222 2920 1223
rect 3262 1223 3268 1224
rect 3262 1222 3263 1223
rect 2919 1220 3041 1222
rect 3253 1220 3263 1222
rect 2919 1219 2920 1220
rect 2914 1218 2920 1219
rect 3262 1219 3263 1220
rect 3267 1219 3268 1223
rect 3450 1223 3456 1224
rect 3450 1222 3451 1223
rect 3421 1220 3451 1222
rect 3262 1218 3268 1219
rect 3450 1219 3451 1220
rect 3455 1219 3456 1223
rect 3450 1218 3456 1219
rect 3564 1216 3566 1221
rect 2722 1215 2728 1216
rect 2722 1211 2723 1215
rect 2727 1211 2728 1215
rect 2722 1210 2728 1211
rect 3562 1215 3568 1216
rect 3562 1211 3563 1215
rect 3567 1211 3568 1215
rect 3562 1210 3568 1211
rect 3590 1212 3596 1213
rect 3590 1208 3591 1212
rect 3595 1208 3596 1212
rect 3590 1207 3596 1208
rect 1864 1200 1966 1202
rect 263 1199 272 1200
rect 263 1195 264 1199
rect 271 1195 272 1199
rect 263 1194 272 1195
rect 290 1199 296 1200
rect 290 1195 291 1199
rect 295 1198 296 1199
rect 439 1199 445 1200
rect 439 1198 440 1199
rect 295 1196 440 1198
rect 295 1195 296 1196
rect 290 1194 296 1195
rect 439 1195 440 1196
rect 444 1195 445 1199
rect 439 1194 445 1195
rect 466 1199 472 1200
rect 466 1195 467 1199
rect 471 1198 472 1199
rect 615 1199 621 1200
rect 615 1198 616 1199
rect 471 1196 616 1198
rect 471 1195 472 1196
rect 466 1194 472 1195
rect 615 1195 616 1196
rect 620 1195 621 1199
rect 615 1194 621 1195
rect 783 1199 789 1200
rect 783 1195 784 1199
rect 788 1198 789 1199
rect 934 1199 940 1200
rect 934 1198 935 1199
rect 788 1196 935 1198
rect 788 1195 789 1196
rect 783 1194 789 1195
rect 934 1195 935 1196
rect 939 1195 940 1199
rect 934 1194 940 1195
rect 942 1199 948 1200
rect 942 1195 943 1199
rect 947 1198 948 1199
rect 951 1199 957 1200
rect 951 1198 952 1199
rect 947 1196 952 1198
rect 947 1195 948 1196
rect 942 1194 948 1195
rect 951 1195 952 1196
rect 956 1195 957 1199
rect 951 1194 957 1195
rect 1103 1199 1109 1200
rect 1103 1195 1104 1199
rect 1108 1198 1109 1199
rect 1122 1199 1128 1200
rect 1122 1198 1123 1199
rect 1108 1196 1123 1198
rect 1108 1195 1109 1196
rect 1103 1194 1109 1195
rect 1122 1195 1123 1196
rect 1127 1195 1128 1199
rect 1122 1194 1128 1195
rect 1130 1199 1136 1200
rect 1130 1195 1131 1199
rect 1135 1198 1136 1199
rect 1247 1199 1253 1200
rect 1247 1198 1248 1199
rect 1135 1196 1248 1198
rect 1135 1195 1136 1196
rect 1130 1194 1136 1195
rect 1247 1195 1248 1196
rect 1252 1195 1253 1199
rect 1247 1194 1253 1195
rect 1274 1199 1280 1200
rect 1274 1195 1275 1199
rect 1279 1198 1280 1199
rect 1391 1199 1397 1200
rect 1391 1198 1392 1199
rect 1279 1196 1392 1198
rect 1279 1195 1280 1196
rect 1274 1194 1280 1195
rect 1391 1195 1392 1196
rect 1396 1195 1397 1199
rect 1391 1194 1397 1195
rect 1418 1199 1424 1200
rect 1418 1195 1419 1199
rect 1423 1198 1424 1199
rect 1527 1199 1533 1200
rect 1527 1198 1528 1199
rect 1423 1196 1528 1198
rect 1423 1195 1424 1196
rect 1418 1194 1424 1195
rect 1527 1195 1528 1196
rect 1532 1195 1533 1199
rect 1527 1194 1533 1195
rect 1554 1199 1560 1200
rect 1554 1195 1555 1199
rect 1559 1198 1560 1199
rect 1663 1199 1669 1200
rect 1663 1198 1664 1199
rect 1559 1196 1664 1198
rect 1559 1195 1560 1196
rect 1554 1194 1560 1195
rect 1663 1195 1664 1196
rect 1668 1195 1669 1199
rect 1663 1194 1669 1195
rect 1775 1199 1781 1200
rect 1775 1195 1776 1199
rect 1780 1198 1781 1199
rect 1802 1199 1808 1200
rect 1802 1198 1803 1199
rect 1780 1196 1803 1198
rect 1780 1195 1781 1196
rect 1775 1194 1781 1195
rect 1802 1195 1803 1196
rect 1807 1195 1808 1199
rect 1802 1194 1808 1195
rect 1902 1194 1908 1195
rect 238 1190 244 1191
rect 238 1186 239 1190
rect 243 1186 244 1190
rect 238 1185 244 1186
rect 414 1190 420 1191
rect 414 1186 415 1190
rect 419 1186 420 1190
rect 414 1185 420 1186
rect 590 1190 596 1191
rect 590 1186 591 1190
rect 595 1186 596 1190
rect 590 1185 596 1186
rect 758 1190 764 1191
rect 758 1186 759 1190
rect 763 1186 764 1190
rect 758 1185 764 1186
rect 926 1190 932 1191
rect 926 1186 927 1190
rect 931 1186 932 1190
rect 926 1185 932 1186
rect 1078 1190 1084 1191
rect 1078 1186 1079 1190
rect 1083 1186 1084 1190
rect 1078 1185 1084 1186
rect 1222 1190 1228 1191
rect 1222 1186 1223 1190
rect 1227 1186 1228 1190
rect 1222 1185 1228 1186
rect 1366 1190 1372 1191
rect 1366 1186 1367 1190
rect 1371 1186 1372 1190
rect 1366 1185 1372 1186
rect 1502 1190 1508 1191
rect 1502 1186 1503 1190
rect 1507 1186 1508 1190
rect 1502 1185 1508 1186
rect 1638 1190 1644 1191
rect 1638 1186 1639 1190
rect 1643 1186 1644 1190
rect 1638 1185 1644 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1902 1190 1903 1194
rect 1907 1190 1908 1194
rect 1902 1189 1908 1190
rect 2078 1194 2084 1195
rect 2078 1190 2079 1194
rect 2083 1190 2084 1194
rect 2078 1189 2084 1190
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2478 1194 2484 1195
rect 2478 1190 2479 1194
rect 2483 1190 2484 1194
rect 2478 1189 2484 1190
rect 2670 1194 2676 1195
rect 2670 1190 2671 1194
rect 2675 1190 2676 1194
rect 2670 1189 2676 1190
rect 2854 1194 2860 1195
rect 2854 1190 2855 1194
rect 2859 1190 2860 1194
rect 2854 1189 2860 1190
rect 3030 1194 3036 1195
rect 3030 1190 3031 1194
rect 3035 1190 3036 1194
rect 3030 1189 3036 1190
rect 3198 1194 3204 1195
rect 3198 1190 3199 1194
rect 3203 1190 3204 1194
rect 3198 1189 3204 1190
rect 3366 1194 3372 1195
rect 3366 1190 3367 1194
rect 3371 1190 3372 1194
rect 3366 1189 3372 1190
rect 3510 1194 3516 1195
rect 3510 1190 3511 1194
rect 3515 1190 3516 1194
rect 3510 1189 3516 1190
rect 1750 1185 1756 1186
rect 1802 1183 1808 1184
rect 1802 1179 1803 1183
rect 1807 1182 1808 1183
rect 1927 1183 1933 1184
rect 1927 1182 1928 1183
rect 1807 1180 1928 1182
rect 1807 1179 1808 1180
rect 1802 1178 1808 1179
rect 1927 1179 1928 1180
rect 1932 1179 1933 1183
rect 1927 1178 1933 1179
rect 2103 1183 2109 1184
rect 2103 1179 2104 1183
rect 2108 1182 2109 1183
rect 2138 1183 2144 1184
rect 2138 1182 2139 1183
rect 2108 1180 2139 1182
rect 2108 1179 2109 1180
rect 2103 1178 2109 1179
rect 2138 1179 2139 1180
rect 2143 1179 2144 1183
rect 2138 1178 2144 1179
rect 2234 1183 2240 1184
rect 2234 1179 2235 1183
rect 2239 1182 2240 1183
rect 2303 1183 2309 1184
rect 2303 1182 2304 1183
rect 2239 1180 2304 1182
rect 2239 1179 2240 1180
rect 2234 1178 2240 1179
rect 2303 1179 2304 1180
rect 2308 1179 2309 1183
rect 2303 1178 2309 1179
rect 2503 1183 2512 1184
rect 2503 1179 2504 1183
rect 2511 1179 2512 1183
rect 2503 1178 2512 1179
rect 2590 1183 2596 1184
rect 2590 1179 2591 1183
rect 2595 1182 2596 1183
rect 2695 1183 2701 1184
rect 2695 1182 2696 1183
rect 2595 1180 2696 1182
rect 2595 1179 2596 1180
rect 2590 1178 2596 1179
rect 2695 1179 2696 1180
rect 2700 1179 2701 1183
rect 2695 1178 2701 1179
rect 2879 1183 2885 1184
rect 2879 1179 2880 1183
rect 2884 1182 2885 1183
rect 2914 1183 2920 1184
rect 2914 1182 2915 1183
rect 2884 1180 2915 1182
rect 2884 1179 2885 1180
rect 2879 1178 2885 1179
rect 2914 1179 2915 1180
rect 2919 1179 2920 1183
rect 2914 1178 2920 1179
rect 3055 1183 3061 1184
rect 3055 1179 3056 1183
rect 3060 1179 3061 1183
rect 3055 1178 3061 1179
rect 3223 1183 3229 1184
rect 3223 1179 3224 1183
rect 3228 1182 3229 1183
rect 3262 1183 3268 1184
rect 3228 1180 3258 1182
rect 3228 1179 3229 1180
rect 3223 1178 3229 1179
rect 3256 1174 3258 1180
rect 3262 1179 3263 1183
rect 3267 1182 3268 1183
rect 3391 1183 3397 1184
rect 3391 1182 3392 1183
rect 3267 1180 3392 1182
rect 3267 1179 3268 1180
rect 3262 1178 3268 1179
rect 3391 1179 3392 1180
rect 3396 1179 3397 1183
rect 3391 1178 3397 1179
rect 3450 1183 3456 1184
rect 3450 1179 3451 1183
rect 3455 1182 3456 1183
rect 3535 1183 3541 1184
rect 3535 1182 3536 1183
rect 3455 1180 3536 1182
rect 3455 1179 3456 1180
rect 3450 1178 3456 1179
rect 3535 1179 3536 1180
rect 3540 1179 3541 1183
rect 3535 1178 3541 1179
rect 3406 1175 3412 1176
rect 3406 1174 3407 1175
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 1830 1172 1836 1173
rect 3256 1172 3407 1174
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 3406 1171 3407 1172
rect 3411 1171 3412 1175
rect 3406 1170 3412 1171
rect 1830 1167 1836 1168
rect 1927 1167 1933 1168
rect 290 1163 296 1164
rect 290 1159 291 1163
rect 295 1159 296 1163
rect 290 1158 296 1159
rect 466 1163 472 1164
rect 466 1159 467 1163
rect 471 1159 472 1163
rect 466 1158 472 1159
rect 810 1163 816 1164
rect 810 1159 811 1163
rect 815 1159 816 1163
rect 810 1158 816 1159
rect 934 1163 940 1164
rect 934 1159 935 1163
rect 939 1159 940 1163
rect 934 1158 940 1159
rect 1130 1163 1136 1164
rect 1130 1159 1131 1163
rect 1135 1159 1136 1163
rect 1130 1158 1136 1159
rect 1274 1163 1280 1164
rect 1274 1159 1275 1163
rect 1279 1159 1280 1163
rect 1274 1158 1280 1159
rect 1418 1163 1424 1164
rect 1418 1159 1419 1163
rect 1423 1159 1424 1163
rect 1418 1158 1424 1159
rect 1554 1163 1560 1164
rect 1554 1159 1555 1163
rect 1559 1159 1560 1163
rect 1554 1158 1560 1159
rect 1802 1163 1808 1164
rect 1802 1159 1803 1163
rect 1807 1159 1808 1163
rect 1927 1163 1928 1167
rect 1932 1166 1933 1167
rect 1954 1167 1960 1168
rect 1954 1166 1955 1167
rect 1932 1164 1955 1166
rect 1932 1163 1933 1164
rect 1927 1162 1933 1163
rect 1954 1163 1955 1164
rect 1959 1163 1960 1167
rect 1954 1162 1960 1163
rect 1962 1167 1968 1168
rect 1962 1163 1963 1167
rect 1967 1166 1968 1167
rect 2007 1167 2013 1168
rect 2007 1166 2008 1167
rect 1967 1164 2008 1166
rect 1967 1163 1968 1164
rect 1962 1162 1968 1163
rect 2007 1163 2008 1164
rect 2012 1163 2013 1167
rect 2007 1162 2013 1163
rect 2034 1167 2040 1168
rect 2034 1163 2035 1167
rect 2039 1166 2040 1167
rect 2111 1167 2117 1168
rect 2111 1166 2112 1167
rect 2039 1164 2112 1166
rect 2039 1163 2040 1164
rect 2034 1162 2040 1163
rect 2111 1163 2112 1164
rect 2116 1163 2117 1167
rect 2111 1162 2117 1163
rect 2138 1167 2144 1168
rect 2138 1163 2139 1167
rect 2143 1166 2144 1167
rect 2239 1167 2245 1168
rect 2239 1166 2240 1167
rect 2143 1164 2240 1166
rect 2143 1163 2144 1164
rect 2138 1162 2144 1163
rect 2239 1163 2240 1164
rect 2244 1163 2245 1167
rect 2239 1162 2245 1163
rect 2266 1167 2272 1168
rect 2266 1163 2267 1167
rect 2271 1166 2272 1167
rect 2391 1167 2397 1168
rect 2391 1166 2392 1167
rect 2271 1164 2392 1166
rect 2271 1163 2272 1164
rect 2266 1162 2272 1163
rect 2391 1163 2392 1164
rect 2396 1163 2397 1167
rect 2391 1162 2397 1163
rect 2418 1167 2424 1168
rect 2418 1163 2419 1167
rect 2423 1166 2424 1167
rect 2551 1167 2557 1168
rect 2551 1166 2552 1167
rect 2423 1164 2552 1166
rect 2423 1163 2424 1164
rect 2418 1162 2424 1163
rect 2551 1163 2552 1164
rect 2556 1163 2557 1167
rect 2551 1162 2557 1163
rect 2711 1167 2717 1168
rect 2711 1163 2712 1167
rect 2716 1166 2717 1167
rect 2722 1167 2728 1168
rect 2722 1166 2723 1167
rect 2716 1164 2723 1166
rect 2716 1163 2717 1164
rect 2711 1162 2717 1163
rect 2722 1163 2723 1164
rect 2727 1163 2728 1167
rect 2722 1162 2728 1163
rect 2738 1167 2744 1168
rect 2738 1163 2739 1167
rect 2743 1166 2744 1167
rect 2863 1167 2869 1168
rect 2863 1166 2864 1167
rect 2743 1164 2864 1166
rect 2743 1163 2744 1164
rect 2738 1162 2744 1163
rect 2863 1163 2864 1164
rect 2868 1163 2869 1167
rect 2863 1162 2869 1163
rect 3007 1167 3016 1168
rect 3007 1163 3008 1167
rect 3015 1163 3016 1167
rect 3007 1162 3016 1163
rect 3087 1167 3093 1168
rect 3087 1163 3088 1167
rect 3092 1166 3093 1167
rect 3151 1167 3157 1168
rect 3151 1166 3152 1167
rect 3092 1164 3152 1166
rect 3092 1163 3093 1164
rect 3087 1162 3093 1163
rect 3151 1163 3152 1164
rect 3156 1163 3157 1167
rect 3151 1162 3157 1163
rect 3178 1167 3184 1168
rect 3178 1163 3179 1167
rect 3183 1166 3184 1167
rect 3287 1167 3293 1168
rect 3287 1166 3288 1167
rect 3183 1164 3288 1166
rect 3183 1163 3184 1164
rect 3178 1162 3184 1163
rect 3287 1163 3288 1164
rect 3292 1163 3293 1167
rect 3287 1162 3293 1163
rect 3314 1167 3320 1168
rect 3314 1163 3315 1167
rect 3319 1166 3320 1167
rect 3423 1167 3429 1168
rect 3423 1166 3424 1167
rect 3319 1164 3424 1166
rect 3319 1163 3320 1164
rect 3314 1162 3320 1163
rect 3423 1163 3424 1164
rect 3428 1163 3429 1167
rect 3423 1162 3429 1163
rect 3535 1167 3541 1168
rect 3535 1163 3536 1167
rect 3540 1166 3541 1167
rect 3562 1167 3568 1168
rect 3562 1166 3563 1167
rect 3540 1164 3563 1166
rect 3540 1163 3541 1164
rect 3535 1162 3541 1163
rect 3562 1163 3563 1164
rect 3567 1163 3568 1167
rect 3562 1162 3568 1163
rect 1802 1158 1808 1159
rect 1902 1158 1908 1159
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 1830 1155 1836 1156
rect 110 1150 116 1151
rect 230 1152 236 1153
rect 230 1148 231 1152
rect 235 1148 236 1152
rect 230 1147 236 1148
rect 406 1152 412 1153
rect 406 1148 407 1152
rect 411 1148 412 1152
rect 406 1147 412 1148
rect 582 1152 588 1153
rect 582 1148 583 1152
rect 587 1148 588 1152
rect 582 1147 588 1148
rect 750 1152 756 1153
rect 750 1148 751 1152
rect 755 1148 756 1152
rect 750 1147 756 1148
rect 918 1152 924 1153
rect 918 1148 919 1152
rect 923 1148 924 1152
rect 918 1147 924 1148
rect 1070 1152 1076 1153
rect 1070 1148 1071 1152
rect 1075 1148 1076 1152
rect 1070 1147 1076 1148
rect 1214 1152 1220 1153
rect 1214 1148 1215 1152
rect 1219 1148 1220 1152
rect 1214 1147 1220 1148
rect 1358 1152 1364 1153
rect 1358 1148 1359 1152
rect 1363 1148 1364 1152
rect 1358 1147 1364 1148
rect 1494 1152 1500 1153
rect 1494 1148 1495 1152
rect 1499 1148 1500 1152
rect 1494 1147 1500 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1902 1154 1903 1158
rect 1907 1154 1908 1158
rect 1902 1153 1908 1154
rect 1982 1158 1988 1159
rect 1982 1154 1983 1158
rect 1987 1154 1988 1158
rect 1982 1153 1988 1154
rect 2086 1158 2092 1159
rect 2086 1154 2087 1158
rect 2091 1154 2092 1158
rect 2086 1153 2092 1154
rect 2214 1158 2220 1159
rect 2214 1154 2215 1158
rect 2219 1154 2220 1158
rect 2214 1153 2220 1154
rect 2366 1158 2372 1159
rect 2366 1154 2367 1158
rect 2371 1154 2372 1158
rect 2366 1153 2372 1154
rect 2526 1158 2532 1159
rect 2526 1154 2527 1158
rect 2531 1154 2532 1158
rect 2526 1153 2532 1154
rect 2686 1158 2692 1159
rect 2686 1154 2687 1158
rect 2691 1154 2692 1158
rect 2686 1153 2692 1154
rect 2838 1158 2844 1159
rect 2838 1154 2839 1158
rect 2843 1154 2844 1158
rect 2838 1153 2844 1154
rect 2982 1158 2988 1159
rect 2982 1154 2983 1158
rect 2987 1154 2988 1158
rect 2982 1153 2988 1154
rect 3126 1158 3132 1159
rect 3126 1154 3127 1158
rect 3131 1154 3132 1158
rect 3126 1153 3132 1154
rect 3262 1158 3268 1159
rect 3262 1154 3263 1158
rect 3267 1154 3268 1158
rect 3262 1153 3268 1154
rect 3398 1158 3404 1159
rect 3398 1154 3399 1158
rect 3403 1154 3404 1158
rect 3398 1153 3404 1154
rect 3510 1158 3516 1159
rect 3510 1154 3511 1158
rect 3515 1154 3516 1158
rect 3510 1153 3516 1154
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 1870 1140 1876 1141
rect 1870 1136 1871 1140
rect 1875 1136 1876 1140
rect 458 1135 464 1136
rect 458 1131 459 1135
rect 463 1134 464 1135
rect 599 1135 605 1136
rect 599 1134 600 1135
rect 463 1132 600 1134
rect 463 1131 464 1132
rect 458 1130 464 1131
rect 599 1131 600 1132
rect 604 1131 605 1135
rect 599 1130 605 1131
rect 1287 1135 1293 1136
rect 1287 1131 1288 1135
rect 1292 1134 1293 1135
rect 1647 1135 1653 1136
rect 1870 1135 1876 1136
rect 3590 1140 3596 1141
rect 3590 1136 3591 1140
rect 3595 1136 3596 1140
rect 3590 1135 3596 1136
rect 1647 1134 1648 1135
rect 1292 1132 1648 1134
rect 1292 1131 1293 1132
rect 1287 1130 1293 1131
rect 1647 1131 1648 1132
rect 1652 1131 1653 1135
rect 1647 1130 1653 1131
rect 1962 1131 1968 1132
rect 1962 1130 1963 1131
rect 1957 1128 1963 1130
rect 1122 1127 1128 1128
rect 1122 1123 1123 1127
rect 1127 1126 1128 1127
rect 1438 1127 1444 1128
rect 1438 1126 1439 1127
rect 1127 1124 1439 1126
rect 1127 1123 1128 1124
rect 1122 1122 1128 1123
rect 1438 1123 1439 1124
rect 1443 1123 1444 1127
rect 1962 1127 1963 1128
rect 1967 1127 1968 1131
rect 1962 1126 1968 1127
rect 2034 1131 2040 1132
rect 2034 1127 2035 1131
rect 2039 1127 2040 1131
rect 2034 1126 2040 1127
rect 2138 1131 2144 1132
rect 2138 1127 2139 1131
rect 2143 1127 2144 1131
rect 2138 1126 2144 1127
rect 2266 1131 2272 1132
rect 2266 1127 2267 1131
rect 2271 1127 2272 1131
rect 2266 1126 2272 1127
rect 2418 1131 2424 1132
rect 2418 1127 2419 1131
rect 2423 1127 2424 1131
rect 2418 1126 2424 1127
rect 2738 1131 2744 1132
rect 2738 1127 2739 1131
rect 2743 1127 2744 1131
rect 2918 1131 2924 1132
rect 2918 1130 2919 1131
rect 2893 1128 2919 1130
rect 2738 1126 2744 1127
rect 2918 1127 2919 1128
rect 2923 1127 2924 1131
rect 3087 1131 3093 1132
rect 3087 1130 3088 1131
rect 3037 1128 3088 1130
rect 2918 1126 2924 1127
rect 3087 1127 3088 1128
rect 3092 1127 3093 1131
rect 3087 1126 3093 1127
rect 3178 1131 3184 1132
rect 3178 1127 3179 1131
rect 3183 1127 3184 1131
rect 3178 1126 3184 1127
rect 3314 1131 3320 1132
rect 3314 1127 3315 1131
rect 3319 1127 3320 1131
rect 3314 1126 3320 1127
rect 3406 1131 3412 1132
rect 3406 1127 3407 1131
rect 3411 1127 3412 1131
rect 3406 1126 3412 1127
rect 3534 1131 3540 1132
rect 3534 1127 3535 1131
rect 3539 1127 3540 1131
rect 3534 1126 3540 1127
rect 1438 1122 1444 1123
rect 1870 1123 1876 1124
rect 1870 1119 1871 1123
rect 1875 1119 1876 1123
rect 3590 1123 3596 1124
rect 1870 1118 1876 1119
rect 1894 1120 1900 1121
rect 1894 1116 1895 1120
rect 1899 1116 1900 1120
rect 1894 1115 1900 1116
rect 1974 1120 1980 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 2078 1120 2084 1121
rect 2078 1116 2079 1120
rect 2083 1116 2084 1120
rect 2078 1115 2084 1116
rect 2206 1120 2212 1121
rect 2206 1116 2207 1120
rect 2211 1116 2212 1120
rect 2206 1115 2212 1116
rect 2358 1120 2364 1121
rect 2358 1116 2359 1120
rect 2363 1116 2364 1120
rect 2358 1115 2364 1116
rect 2518 1120 2524 1121
rect 2518 1116 2519 1120
rect 2523 1116 2524 1120
rect 2518 1115 2524 1116
rect 2678 1120 2684 1121
rect 2678 1116 2679 1120
rect 2683 1116 2684 1120
rect 2678 1115 2684 1116
rect 2830 1120 2836 1121
rect 2830 1116 2831 1120
rect 2835 1116 2836 1120
rect 2830 1115 2836 1116
rect 2974 1120 2980 1121
rect 2974 1116 2975 1120
rect 2979 1116 2980 1120
rect 2974 1115 2980 1116
rect 3118 1120 3124 1121
rect 3118 1116 3119 1120
rect 3123 1116 3124 1120
rect 3118 1115 3124 1116
rect 3254 1120 3260 1121
rect 3254 1116 3255 1120
rect 3259 1116 3260 1120
rect 3254 1115 3260 1116
rect 3390 1120 3396 1121
rect 3390 1116 3391 1120
rect 3395 1116 3396 1120
rect 3390 1115 3396 1116
rect 3502 1120 3508 1121
rect 3502 1116 3503 1120
rect 3507 1116 3508 1120
rect 3590 1119 3591 1123
rect 3595 1119 3596 1123
rect 3590 1118 3596 1119
rect 3502 1115 3508 1116
rect 142 1104 148 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 142 1100 143 1104
rect 147 1100 148 1104
rect 142 1099 148 1100
rect 278 1104 284 1105
rect 278 1100 279 1104
rect 283 1100 284 1104
rect 278 1099 284 1100
rect 422 1104 428 1105
rect 422 1100 423 1104
rect 427 1100 428 1104
rect 422 1099 428 1100
rect 566 1104 572 1105
rect 566 1100 567 1104
rect 571 1100 572 1104
rect 566 1099 572 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 846 1104 852 1105
rect 846 1100 847 1104
rect 851 1100 852 1104
rect 846 1099 852 1100
rect 974 1104 980 1105
rect 974 1100 975 1104
rect 979 1100 980 1104
rect 974 1099 980 1100
rect 1102 1104 1108 1105
rect 1102 1100 1103 1104
rect 1107 1100 1108 1104
rect 1102 1099 1108 1100
rect 1222 1104 1228 1105
rect 1222 1100 1223 1104
rect 1227 1100 1228 1104
rect 1222 1099 1228 1100
rect 1342 1104 1348 1105
rect 1342 1100 1343 1104
rect 1347 1100 1348 1104
rect 1342 1099 1348 1100
rect 1470 1104 1476 1105
rect 1470 1100 1471 1104
rect 1475 1100 1476 1104
rect 2214 1103 2220 1104
rect 1470 1099 1476 1100
rect 1830 1101 1836 1102
rect 110 1096 116 1097
rect 1830 1097 1831 1101
rect 1835 1097 1836 1101
rect 2214 1099 2215 1103
rect 2219 1102 2220 1103
rect 2535 1103 2541 1104
rect 2535 1102 2536 1103
rect 2219 1100 2536 1102
rect 2219 1099 2220 1100
rect 2214 1098 2220 1099
rect 2535 1099 2536 1100
rect 2540 1099 2541 1103
rect 2535 1098 2541 1099
rect 1830 1096 1836 1097
rect 210 1095 216 1096
rect 204 1088 206 1093
rect 210 1091 211 1095
rect 215 1094 216 1095
rect 346 1095 352 1096
rect 215 1092 297 1094
rect 215 1091 216 1092
rect 210 1090 216 1091
rect 346 1091 347 1095
rect 351 1094 352 1095
rect 634 1095 640 1096
rect 634 1094 635 1095
rect 351 1092 441 1094
rect 629 1092 635 1094
rect 351 1091 352 1092
rect 346 1090 352 1091
rect 634 1091 635 1092
rect 639 1091 640 1095
rect 802 1095 808 1096
rect 802 1094 803 1095
rect 773 1092 803 1094
rect 634 1090 640 1091
rect 802 1091 803 1092
rect 807 1091 808 1095
rect 942 1095 948 1096
rect 942 1094 943 1095
rect 909 1092 943 1094
rect 802 1090 808 1091
rect 942 1091 943 1092
rect 947 1091 948 1095
rect 1062 1095 1068 1096
rect 1062 1094 1063 1095
rect 1037 1092 1063 1094
rect 942 1090 948 1091
rect 1062 1091 1063 1092
rect 1067 1091 1068 1095
rect 1186 1095 1192 1096
rect 1186 1094 1187 1095
rect 1165 1092 1187 1094
rect 1062 1090 1068 1091
rect 1186 1091 1187 1092
rect 1191 1091 1192 1095
rect 1306 1095 1312 1096
rect 1306 1094 1307 1095
rect 1285 1092 1307 1094
rect 1186 1090 1192 1091
rect 1306 1091 1307 1092
rect 1311 1091 1312 1095
rect 1430 1095 1436 1096
rect 1430 1094 1431 1095
rect 1405 1092 1431 1094
rect 1306 1090 1312 1091
rect 1430 1091 1431 1092
rect 1435 1091 1436 1095
rect 1430 1090 1436 1091
rect 1438 1095 1444 1096
rect 1438 1091 1439 1095
rect 1443 1094 1444 1095
rect 1443 1092 1489 1094
rect 1443 1091 1444 1092
rect 1438 1090 1444 1091
rect 202 1087 208 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 202 1083 203 1087
rect 207 1083 208 1087
rect 202 1082 208 1083
rect 1830 1084 1836 1085
rect 110 1079 116 1080
rect 1830 1080 1831 1084
rect 1835 1080 1836 1084
rect 1830 1079 1836 1080
rect 2166 1068 2172 1069
rect 150 1066 156 1067
rect 150 1062 151 1066
rect 155 1062 156 1066
rect 150 1061 156 1062
rect 286 1066 292 1067
rect 286 1062 287 1066
rect 291 1062 292 1066
rect 286 1061 292 1062
rect 430 1066 436 1067
rect 430 1062 431 1066
rect 435 1062 436 1066
rect 430 1061 436 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 718 1066 724 1067
rect 718 1062 719 1066
rect 723 1062 724 1066
rect 718 1061 724 1062
rect 854 1066 860 1067
rect 854 1062 855 1066
rect 859 1062 860 1066
rect 854 1061 860 1062
rect 982 1066 988 1067
rect 982 1062 983 1066
rect 987 1062 988 1066
rect 982 1061 988 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1230 1066 1236 1067
rect 1230 1062 1231 1066
rect 1235 1062 1236 1066
rect 1230 1061 1236 1062
rect 1350 1066 1356 1067
rect 1350 1062 1351 1066
rect 1355 1062 1356 1066
rect 1350 1061 1356 1062
rect 1478 1066 1484 1067
rect 1478 1062 1479 1066
rect 1483 1062 1484 1066
rect 1478 1061 1484 1062
rect 1870 1065 1876 1066
rect 1870 1061 1871 1065
rect 1875 1061 1876 1065
rect 2166 1064 2167 1068
rect 2171 1064 2172 1068
rect 2166 1063 2172 1064
rect 2254 1068 2260 1069
rect 2254 1064 2255 1068
rect 2259 1064 2260 1068
rect 2254 1063 2260 1064
rect 2358 1068 2364 1069
rect 2358 1064 2359 1068
rect 2363 1064 2364 1068
rect 2358 1063 2364 1064
rect 2478 1068 2484 1069
rect 2478 1064 2479 1068
rect 2483 1064 2484 1068
rect 2478 1063 2484 1064
rect 2606 1068 2612 1069
rect 2606 1064 2607 1068
rect 2611 1064 2612 1068
rect 2606 1063 2612 1064
rect 2750 1068 2756 1069
rect 2750 1064 2751 1068
rect 2755 1064 2756 1068
rect 2750 1063 2756 1064
rect 2894 1068 2900 1069
rect 2894 1064 2895 1068
rect 2899 1064 2900 1068
rect 2894 1063 2900 1064
rect 3046 1068 3052 1069
rect 3046 1064 3047 1068
rect 3051 1064 3052 1068
rect 3046 1063 3052 1064
rect 3206 1068 3212 1069
rect 3206 1064 3207 1068
rect 3211 1064 3212 1068
rect 3206 1063 3212 1064
rect 3366 1068 3372 1069
rect 3366 1064 3367 1068
rect 3371 1064 3372 1068
rect 3366 1063 3372 1064
rect 3502 1068 3508 1069
rect 3502 1064 3503 1068
rect 3507 1064 3508 1068
rect 3502 1063 3508 1064
rect 3590 1065 3596 1066
rect 1870 1060 1876 1061
rect 3590 1061 3591 1065
rect 3595 1061 3596 1065
rect 3590 1060 3596 1061
rect 2234 1059 2240 1060
rect 2234 1058 2235 1059
rect 2229 1056 2235 1058
rect 175 1055 181 1056
rect 175 1051 176 1055
rect 180 1054 181 1055
rect 210 1055 216 1056
rect 210 1054 211 1055
rect 180 1052 211 1054
rect 180 1051 181 1052
rect 175 1050 181 1051
rect 210 1051 211 1052
rect 215 1051 216 1055
rect 210 1050 216 1051
rect 311 1055 317 1056
rect 311 1051 312 1055
rect 316 1054 317 1055
rect 346 1055 352 1056
rect 346 1054 347 1055
rect 316 1052 347 1054
rect 316 1051 317 1052
rect 311 1050 317 1051
rect 346 1051 347 1052
rect 351 1051 352 1055
rect 346 1050 352 1051
rect 455 1055 464 1056
rect 455 1051 456 1055
rect 463 1051 464 1055
rect 455 1050 464 1051
rect 598 1055 605 1056
rect 598 1051 599 1055
rect 604 1051 605 1055
rect 598 1050 605 1051
rect 634 1055 640 1056
rect 634 1051 635 1055
rect 639 1054 640 1055
rect 743 1055 749 1056
rect 743 1054 744 1055
rect 639 1052 744 1054
rect 639 1051 640 1052
rect 634 1050 640 1051
rect 743 1051 744 1052
rect 748 1051 749 1055
rect 743 1050 749 1051
rect 802 1055 808 1056
rect 802 1051 803 1055
rect 807 1054 808 1055
rect 879 1055 885 1056
rect 879 1054 880 1055
rect 807 1052 880 1054
rect 807 1051 808 1052
rect 802 1050 808 1051
rect 879 1051 880 1052
rect 884 1051 885 1055
rect 879 1050 885 1051
rect 1007 1055 1013 1056
rect 1007 1051 1008 1055
rect 1012 1054 1013 1055
rect 1054 1055 1060 1056
rect 1054 1054 1055 1055
rect 1012 1052 1055 1054
rect 1012 1051 1013 1052
rect 1007 1050 1013 1051
rect 1054 1051 1055 1052
rect 1059 1051 1060 1055
rect 1054 1050 1060 1051
rect 1062 1055 1068 1056
rect 1062 1051 1063 1055
rect 1067 1054 1068 1055
rect 1135 1055 1141 1056
rect 1135 1054 1136 1055
rect 1067 1052 1136 1054
rect 1067 1051 1068 1052
rect 1062 1050 1068 1051
rect 1135 1051 1136 1052
rect 1140 1051 1141 1055
rect 1135 1050 1141 1051
rect 1186 1055 1192 1056
rect 1186 1051 1187 1055
rect 1191 1054 1192 1055
rect 1255 1055 1261 1056
rect 1255 1054 1256 1055
rect 1191 1052 1256 1054
rect 1191 1051 1192 1052
rect 1186 1050 1192 1051
rect 1255 1051 1256 1052
rect 1260 1051 1261 1055
rect 1255 1050 1261 1051
rect 1306 1055 1312 1056
rect 1306 1051 1307 1055
rect 1311 1054 1312 1055
rect 1375 1055 1381 1056
rect 1375 1054 1376 1055
rect 1311 1052 1376 1054
rect 1311 1051 1312 1052
rect 1306 1050 1312 1051
rect 1375 1051 1376 1052
rect 1380 1051 1381 1055
rect 1375 1050 1381 1051
rect 1430 1055 1436 1056
rect 1430 1051 1431 1055
rect 1435 1054 1436 1055
rect 1503 1055 1509 1056
rect 1503 1054 1504 1055
rect 1435 1052 1504 1054
rect 1435 1051 1436 1052
rect 1430 1050 1436 1051
rect 1503 1051 1504 1052
rect 1508 1051 1509 1055
rect 2234 1055 2235 1056
rect 2239 1055 2240 1059
rect 2330 1059 2336 1060
rect 2330 1058 2331 1059
rect 2317 1056 2331 1058
rect 2234 1054 2240 1055
rect 2330 1055 2331 1056
rect 2335 1055 2336 1059
rect 2434 1059 2440 1060
rect 2434 1058 2435 1059
rect 2421 1056 2435 1058
rect 2330 1054 2336 1055
rect 2434 1055 2435 1056
rect 2439 1055 2440 1059
rect 2554 1059 2560 1060
rect 2554 1058 2555 1059
rect 2541 1056 2555 1058
rect 2434 1054 2440 1055
rect 2554 1055 2555 1056
rect 2559 1055 2560 1059
rect 2554 1054 2560 1055
rect 2562 1059 2568 1060
rect 2562 1055 2563 1059
rect 2567 1058 2568 1059
rect 2818 1059 2824 1060
rect 2567 1056 2625 1058
rect 2567 1055 2568 1056
rect 2562 1054 2568 1055
rect 2812 1052 2814 1057
rect 2818 1055 2819 1059
rect 2823 1058 2824 1059
rect 3010 1059 3016 1060
rect 2823 1056 2913 1058
rect 2823 1055 2824 1056
rect 2818 1054 2824 1055
rect 3010 1055 3011 1059
rect 3015 1058 3016 1059
rect 3114 1059 3120 1060
rect 3015 1056 3065 1058
rect 3015 1055 3016 1056
rect 3010 1054 3016 1055
rect 3114 1055 3115 1059
rect 3119 1058 3120 1059
rect 3274 1059 3280 1060
rect 3119 1056 3225 1058
rect 3119 1055 3120 1056
rect 3114 1054 3120 1055
rect 3274 1055 3275 1059
rect 3279 1058 3280 1059
rect 3279 1056 3385 1058
rect 3279 1055 3280 1056
rect 3274 1054 3280 1055
rect 3564 1052 3566 1057
rect 1503 1050 1509 1051
rect 2810 1051 2816 1052
rect 1870 1048 1876 1049
rect 1870 1044 1871 1048
rect 1875 1044 1876 1048
rect 2810 1047 2811 1051
rect 2815 1047 2816 1051
rect 2810 1046 2816 1047
rect 3562 1051 3568 1052
rect 3562 1047 3563 1051
rect 3567 1047 3568 1051
rect 3562 1046 3568 1047
rect 3590 1048 3596 1049
rect 414 1043 420 1044
rect 1870 1043 1876 1044
rect 3590 1044 3591 1048
rect 3595 1044 3596 1048
rect 3590 1043 3596 1044
rect 414 1042 415 1043
rect 196 1040 415 1042
rect 167 1035 173 1036
rect 167 1031 168 1035
rect 172 1034 173 1035
rect 196 1034 198 1040
rect 414 1039 415 1040
rect 419 1039 420 1043
rect 414 1038 420 1039
rect 172 1032 198 1034
rect 202 1035 208 1036
rect 172 1031 173 1032
rect 167 1030 173 1031
rect 202 1031 203 1035
rect 207 1034 208 1035
rect 287 1035 293 1036
rect 287 1034 288 1035
rect 207 1032 288 1034
rect 207 1031 208 1032
rect 202 1030 208 1031
rect 287 1031 288 1032
rect 292 1031 293 1035
rect 287 1030 293 1031
rect 314 1035 320 1036
rect 314 1031 315 1035
rect 319 1034 320 1035
rect 431 1035 437 1036
rect 431 1034 432 1035
rect 319 1032 432 1034
rect 319 1031 320 1032
rect 314 1030 320 1031
rect 431 1031 432 1032
rect 436 1031 437 1035
rect 431 1030 437 1031
rect 575 1035 581 1036
rect 575 1031 576 1035
rect 580 1034 581 1035
rect 694 1035 700 1036
rect 694 1034 695 1035
rect 580 1032 695 1034
rect 580 1031 581 1032
rect 575 1030 581 1031
rect 694 1031 695 1032
rect 699 1031 700 1035
rect 694 1030 700 1031
rect 711 1035 717 1036
rect 711 1031 712 1035
rect 716 1034 717 1035
rect 754 1035 760 1036
rect 754 1034 755 1035
rect 716 1032 755 1034
rect 716 1031 717 1032
rect 711 1030 717 1031
rect 754 1031 755 1032
rect 759 1031 760 1035
rect 754 1030 760 1031
rect 791 1035 797 1036
rect 791 1031 792 1035
rect 796 1034 797 1035
rect 831 1035 837 1036
rect 831 1034 832 1035
rect 796 1032 832 1034
rect 796 1031 797 1032
rect 791 1030 797 1031
rect 831 1031 832 1032
rect 836 1031 837 1035
rect 831 1030 837 1031
rect 918 1035 924 1036
rect 918 1031 919 1035
rect 923 1034 924 1035
rect 951 1035 957 1036
rect 951 1034 952 1035
rect 923 1032 952 1034
rect 923 1031 924 1032
rect 918 1030 924 1031
rect 951 1031 952 1032
rect 956 1031 957 1035
rect 951 1030 957 1031
rect 1030 1035 1036 1036
rect 1030 1031 1031 1035
rect 1035 1034 1036 1035
rect 1063 1035 1069 1036
rect 1063 1034 1064 1035
rect 1035 1032 1064 1034
rect 1035 1031 1036 1032
rect 1030 1030 1036 1031
rect 1063 1031 1064 1032
rect 1068 1031 1069 1035
rect 1063 1030 1069 1031
rect 1090 1035 1096 1036
rect 1090 1031 1091 1035
rect 1095 1034 1096 1035
rect 1167 1035 1173 1036
rect 1167 1034 1168 1035
rect 1095 1032 1168 1034
rect 1095 1031 1096 1032
rect 1090 1030 1096 1031
rect 1167 1031 1168 1032
rect 1172 1031 1173 1035
rect 1167 1030 1173 1031
rect 1194 1035 1200 1036
rect 1194 1031 1195 1035
rect 1199 1034 1200 1035
rect 1271 1035 1277 1036
rect 1271 1034 1272 1035
rect 1199 1032 1272 1034
rect 1199 1031 1200 1032
rect 1194 1030 1200 1031
rect 1271 1031 1272 1032
rect 1276 1031 1277 1035
rect 1271 1030 1277 1031
rect 1298 1035 1304 1036
rect 1298 1031 1299 1035
rect 1303 1034 1304 1035
rect 1383 1035 1389 1036
rect 1383 1034 1384 1035
rect 1303 1032 1384 1034
rect 1303 1031 1304 1032
rect 1298 1030 1304 1031
rect 1383 1031 1384 1032
rect 1388 1031 1389 1035
rect 1383 1030 1389 1031
rect 2174 1030 2180 1031
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 262 1026 268 1027
rect 262 1022 263 1026
rect 267 1022 268 1026
rect 262 1021 268 1022
rect 406 1026 412 1027
rect 406 1022 407 1026
rect 411 1022 412 1026
rect 406 1021 412 1022
rect 550 1026 556 1027
rect 550 1022 551 1026
rect 555 1022 556 1026
rect 550 1021 556 1022
rect 686 1026 692 1027
rect 686 1022 687 1026
rect 691 1022 692 1026
rect 686 1021 692 1022
rect 806 1026 812 1027
rect 806 1022 807 1026
rect 811 1022 812 1026
rect 806 1021 812 1022
rect 926 1026 932 1027
rect 926 1022 927 1026
rect 931 1022 932 1026
rect 926 1021 932 1022
rect 1038 1026 1044 1027
rect 1038 1022 1039 1026
rect 1043 1022 1044 1026
rect 1038 1021 1044 1022
rect 1142 1026 1148 1027
rect 1142 1022 1143 1026
rect 1147 1022 1148 1026
rect 1142 1021 1148 1022
rect 1246 1026 1252 1027
rect 1246 1022 1247 1026
rect 1251 1022 1252 1026
rect 1246 1021 1252 1022
rect 1358 1026 1364 1027
rect 1358 1022 1359 1026
rect 1363 1022 1364 1026
rect 2174 1026 2175 1030
rect 2179 1026 2180 1030
rect 2174 1025 2180 1026
rect 2262 1030 2268 1031
rect 2262 1026 2263 1030
rect 2267 1026 2268 1030
rect 2262 1025 2268 1026
rect 2366 1030 2372 1031
rect 2366 1026 2367 1030
rect 2371 1026 2372 1030
rect 2366 1025 2372 1026
rect 2486 1030 2492 1031
rect 2486 1026 2487 1030
rect 2491 1026 2492 1030
rect 2486 1025 2492 1026
rect 2614 1030 2620 1031
rect 2614 1026 2615 1030
rect 2619 1026 2620 1030
rect 2614 1025 2620 1026
rect 2758 1030 2764 1031
rect 2758 1026 2759 1030
rect 2763 1026 2764 1030
rect 2758 1025 2764 1026
rect 2902 1030 2908 1031
rect 2902 1026 2903 1030
rect 2907 1026 2908 1030
rect 2902 1025 2908 1026
rect 3054 1030 3060 1031
rect 3054 1026 3055 1030
rect 3059 1026 3060 1030
rect 3054 1025 3060 1026
rect 3214 1030 3220 1031
rect 3214 1026 3215 1030
rect 3219 1026 3220 1030
rect 3214 1025 3220 1026
rect 3374 1030 3380 1031
rect 3374 1026 3375 1030
rect 3379 1026 3380 1030
rect 3374 1025 3380 1026
rect 3510 1030 3516 1031
rect 3510 1026 3511 1030
rect 3515 1026 3516 1030
rect 3510 1025 3516 1026
rect 1358 1021 1364 1022
rect 2199 1019 2205 1020
rect 2199 1015 2200 1019
rect 2204 1018 2205 1019
rect 2214 1019 2220 1020
rect 2214 1018 2215 1019
rect 2204 1016 2215 1018
rect 2204 1015 2205 1016
rect 2199 1014 2205 1015
rect 2214 1015 2215 1016
rect 2219 1015 2220 1019
rect 2214 1014 2220 1015
rect 2234 1019 2240 1020
rect 2234 1015 2235 1019
rect 2239 1018 2240 1019
rect 2287 1019 2293 1020
rect 2287 1018 2288 1019
rect 2239 1016 2288 1018
rect 2239 1015 2240 1016
rect 2234 1014 2240 1015
rect 2287 1015 2288 1016
rect 2292 1015 2293 1019
rect 2287 1014 2293 1015
rect 2330 1019 2336 1020
rect 2330 1015 2331 1019
rect 2335 1018 2336 1019
rect 2391 1019 2397 1020
rect 2391 1018 2392 1019
rect 2335 1016 2392 1018
rect 2335 1015 2336 1016
rect 2330 1014 2336 1015
rect 2391 1015 2392 1016
rect 2396 1015 2397 1019
rect 2391 1014 2397 1015
rect 2434 1019 2440 1020
rect 2434 1015 2435 1019
rect 2439 1018 2440 1019
rect 2511 1019 2517 1020
rect 2511 1018 2512 1019
rect 2439 1016 2512 1018
rect 2439 1015 2440 1016
rect 2434 1014 2440 1015
rect 2511 1015 2512 1016
rect 2516 1015 2517 1019
rect 2511 1014 2517 1015
rect 2554 1019 2560 1020
rect 2554 1015 2555 1019
rect 2559 1018 2560 1019
rect 2639 1019 2645 1020
rect 2639 1018 2640 1019
rect 2559 1016 2640 1018
rect 2559 1015 2560 1016
rect 2554 1014 2560 1015
rect 2639 1015 2640 1016
rect 2644 1015 2645 1019
rect 2639 1014 2645 1015
rect 2783 1019 2789 1020
rect 2783 1015 2784 1019
rect 2788 1018 2789 1019
rect 2818 1019 2824 1020
rect 2818 1018 2819 1019
rect 2788 1016 2819 1018
rect 2788 1015 2789 1016
rect 2783 1014 2789 1015
rect 2818 1015 2819 1016
rect 2823 1015 2824 1019
rect 2818 1014 2824 1015
rect 2918 1019 2924 1020
rect 2918 1015 2919 1019
rect 2923 1018 2924 1019
rect 2927 1019 2933 1020
rect 2927 1018 2928 1019
rect 2923 1016 2928 1018
rect 2923 1015 2924 1016
rect 2918 1014 2924 1015
rect 2927 1015 2928 1016
rect 2932 1015 2933 1019
rect 2927 1014 2933 1015
rect 3079 1019 3085 1020
rect 3079 1015 3080 1019
rect 3084 1018 3085 1019
rect 3114 1019 3120 1020
rect 3114 1018 3115 1019
rect 3084 1016 3115 1018
rect 3084 1015 3085 1016
rect 3079 1014 3085 1015
rect 3114 1015 3115 1016
rect 3119 1015 3120 1019
rect 3114 1014 3120 1015
rect 3239 1019 3245 1020
rect 3239 1015 3240 1019
rect 3244 1018 3245 1019
rect 3274 1019 3280 1020
rect 3274 1018 3275 1019
rect 3244 1016 3275 1018
rect 3244 1015 3245 1016
rect 3239 1014 3245 1015
rect 3274 1015 3275 1016
rect 3279 1015 3280 1019
rect 3274 1014 3280 1015
rect 3398 1019 3405 1020
rect 3398 1015 3399 1019
rect 3404 1015 3405 1019
rect 3398 1014 3405 1015
rect 3534 1019 3541 1020
rect 3534 1015 3535 1019
rect 3540 1015 3541 1019
rect 3534 1014 3541 1015
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 2327 1007 2333 1008
rect 2327 1003 2328 1007
rect 2332 1006 2333 1007
rect 2346 1007 2352 1008
rect 2346 1006 2347 1007
rect 2332 1004 2347 1006
rect 2332 1003 2333 1004
rect 2327 1002 2333 1003
rect 2346 1003 2347 1004
rect 2351 1003 2352 1007
rect 2346 1002 2352 1003
rect 2354 1007 2360 1008
rect 2354 1003 2355 1007
rect 2359 1006 2360 1007
rect 2407 1007 2413 1008
rect 2407 1006 2408 1007
rect 2359 1004 2408 1006
rect 2359 1003 2360 1004
rect 2354 1002 2360 1003
rect 2407 1003 2408 1004
rect 2412 1003 2413 1007
rect 2407 1002 2413 1003
rect 2434 1007 2440 1008
rect 2434 1003 2435 1007
rect 2439 1006 2440 1007
rect 2495 1007 2501 1008
rect 2495 1006 2496 1007
rect 2439 1004 2496 1006
rect 2439 1003 2440 1004
rect 2434 1002 2440 1003
rect 2495 1003 2496 1004
rect 2500 1003 2501 1007
rect 2495 1002 2501 1003
rect 2522 1007 2528 1008
rect 2522 1003 2523 1007
rect 2527 1006 2528 1007
rect 2591 1007 2597 1008
rect 2591 1006 2592 1007
rect 2527 1004 2592 1006
rect 2527 1003 2528 1004
rect 2522 1002 2528 1003
rect 2591 1003 2592 1004
rect 2596 1003 2597 1007
rect 2591 1002 2597 1003
rect 2631 1007 2637 1008
rect 2631 1003 2632 1007
rect 2636 1006 2637 1007
rect 2695 1007 2701 1008
rect 2695 1006 2696 1007
rect 2636 1004 2696 1006
rect 2636 1003 2637 1004
rect 2631 1002 2637 1003
rect 2695 1003 2696 1004
rect 2700 1003 2701 1007
rect 2695 1002 2701 1003
rect 2807 1007 2816 1008
rect 2807 1003 2808 1007
rect 2815 1003 2816 1007
rect 2807 1002 2816 1003
rect 2834 1007 2840 1008
rect 2834 1003 2835 1007
rect 2839 1006 2840 1007
rect 2935 1007 2941 1008
rect 2935 1006 2936 1007
rect 2839 1004 2936 1006
rect 2839 1003 2840 1004
rect 2834 1002 2840 1003
rect 2935 1003 2936 1004
rect 2940 1003 2941 1007
rect 2935 1002 2941 1003
rect 3074 1007 3085 1008
rect 3074 1003 3075 1007
rect 3079 1003 3080 1007
rect 3084 1003 3085 1007
rect 3074 1002 3085 1003
rect 3106 1007 3112 1008
rect 3106 1003 3107 1007
rect 3111 1006 3112 1007
rect 3231 1007 3237 1008
rect 3231 1006 3232 1007
rect 3111 1004 3232 1006
rect 3111 1003 3112 1004
rect 3106 1002 3112 1003
rect 3231 1003 3232 1004
rect 3236 1003 3237 1007
rect 3231 1002 3237 1003
rect 3258 1007 3264 1008
rect 3258 1003 3259 1007
rect 3263 1006 3264 1007
rect 3391 1007 3397 1008
rect 3391 1006 3392 1007
rect 3263 1004 3392 1006
rect 3263 1003 3264 1004
rect 3258 1002 3264 1003
rect 3391 1003 3392 1004
rect 3396 1003 3397 1007
rect 3391 1002 3397 1003
rect 3535 1007 3541 1008
rect 3535 1003 3536 1007
rect 3540 1006 3541 1007
rect 3562 1007 3568 1008
rect 3562 1006 3563 1007
rect 3540 1004 3563 1006
rect 3540 1003 3541 1004
rect 3535 1002 3541 1003
rect 3562 1003 3563 1004
rect 3567 1003 3568 1007
rect 3562 1002 3568 1003
rect 166 999 172 1000
rect 166 995 167 999
rect 171 995 172 999
rect 166 994 172 995
rect 314 999 320 1000
rect 314 995 315 999
rect 319 995 320 999
rect 314 994 320 995
rect 414 999 420 1000
rect 414 995 415 999
rect 419 995 420 999
rect 414 994 420 995
rect 598 999 604 1000
rect 598 995 599 999
rect 603 995 604 999
rect 598 994 604 995
rect 694 999 700 1000
rect 694 995 695 999
rect 699 995 700 999
rect 918 999 924 1000
rect 918 998 919 999
rect 861 996 919 998
rect 694 994 700 995
rect 918 995 919 996
rect 923 995 924 999
rect 1030 999 1036 1000
rect 1030 998 1031 999
rect 981 996 1031 998
rect 918 994 924 995
rect 1030 995 1031 996
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1090 999 1096 1000
rect 1090 995 1091 999
rect 1095 995 1096 999
rect 1090 994 1096 995
rect 1194 999 1200 1000
rect 1194 995 1195 999
rect 1199 995 1200 999
rect 1194 994 1200 995
rect 1298 999 1304 1000
rect 1298 995 1299 999
rect 1303 995 1304 999
rect 1298 994 1304 995
rect 1366 999 1372 1000
rect 1366 995 1367 999
rect 1371 995 1372 999
rect 1366 994 1372 995
rect 2302 998 2308 999
rect 2302 994 2303 998
rect 2307 994 2308 998
rect 2302 993 2308 994
rect 2382 998 2388 999
rect 2382 994 2383 998
rect 2387 994 2388 998
rect 2382 993 2388 994
rect 2470 998 2476 999
rect 2470 994 2471 998
rect 2475 994 2476 998
rect 2470 993 2476 994
rect 2566 998 2572 999
rect 2566 994 2567 998
rect 2571 994 2572 998
rect 2566 993 2572 994
rect 2670 998 2676 999
rect 2670 994 2671 998
rect 2675 994 2676 998
rect 2670 993 2676 994
rect 2782 998 2788 999
rect 2782 994 2783 998
rect 2787 994 2788 998
rect 2782 993 2788 994
rect 2910 998 2916 999
rect 2910 994 2911 998
rect 2915 994 2916 998
rect 2910 993 2916 994
rect 3054 998 3060 999
rect 3054 994 3055 998
rect 3059 994 3060 998
rect 3054 993 3060 994
rect 3206 998 3212 999
rect 3206 994 3207 998
rect 3211 994 3212 998
rect 3206 993 3212 994
rect 3366 998 3372 999
rect 3366 994 3367 998
rect 3371 994 3372 998
rect 3366 993 3372 994
rect 3510 998 3516 999
rect 3510 994 3511 998
rect 3515 994 3516 998
rect 3510 993 3516 994
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1830 991 1836 992
rect 110 986 116 987
rect 134 988 140 989
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 254 988 260 989
rect 254 984 255 988
rect 259 984 260 988
rect 254 983 260 984
rect 398 988 404 989
rect 398 984 399 988
rect 403 984 404 988
rect 398 983 404 984
rect 542 988 548 989
rect 542 984 543 988
rect 547 984 548 988
rect 542 983 548 984
rect 678 988 684 989
rect 678 984 679 988
rect 683 984 684 988
rect 678 983 684 984
rect 798 988 804 989
rect 798 984 799 988
rect 803 984 804 988
rect 798 983 804 984
rect 918 988 924 989
rect 918 984 919 988
rect 923 984 924 988
rect 918 983 924 984
rect 1030 988 1036 989
rect 1030 984 1031 988
rect 1035 984 1036 988
rect 1030 983 1036 984
rect 1134 988 1140 989
rect 1134 984 1135 988
rect 1139 984 1140 988
rect 1134 983 1140 984
rect 1238 988 1244 989
rect 1238 984 1239 988
rect 1243 984 1244 988
rect 1238 983 1244 984
rect 1350 988 1356 989
rect 1350 984 1351 988
rect 1355 984 1356 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1350 983 1356 984
rect 1870 980 1876 981
rect 1870 976 1871 980
rect 1875 976 1876 980
rect 1870 975 1876 976
rect 3590 980 3596 981
rect 3590 976 3591 980
rect 3595 976 3596 980
rect 3590 975 3596 976
rect 2354 971 2360 972
rect 2354 967 2355 971
rect 2359 967 2360 971
rect 2354 966 2360 967
rect 2434 971 2440 972
rect 2434 967 2435 971
rect 2439 967 2440 971
rect 2434 966 2440 967
rect 2522 971 2528 972
rect 2522 967 2523 971
rect 2527 967 2528 971
rect 2631 971 2637 972
rect 2631 970 2632 971
rect 2621 968 2632 970
rect 2522 966 2528 967
rect 2631 967 2632 968
rect 2636 967 2637 971
rect 2631 966 2637 967
rect 2722 971 2728 972
rect 2722 967 2723 971
rect 2727 967 2728 971
rect 2722 966 2728 967
rect 2834 971 2840 972
rect 2834 967 2835 971
rect 2839 967 2840 971
rect 2834 966 2840 967
rect 3106 971 3112 972
rect 3106 967 3107 971
rect 3111 967 3112 971
rect 3106 966 3112 967
rect 3258 971 3264 972
rect 3258 967 3259 971
rect 3263 967 3264 971
rect 3258 966 3264 967
rect 3398 971 3404 972
rect 3398 967 3399 971
rect 3403 967 3404 971
rect 3398 966 3404 967
rect 3534 971 3540 972
rect 3534 967 3535 971
rect 3539 967 3540 971
rect 3534 966 3540 967
rect 1870 963 1876 964
rect 1870 959 1871 963
rect 1875 959 1876 963
rect 3590 963 3596 964
rect 1870 958 1876 959
rect 2294 960 2300 961
rect 2294 956 2295 960
rect 2299 956 2300 960
rect 2294 955 2300 956
rect 2374 960 2380 961
rect 2374 956 2375 960
rect 2379 956 2380 960
rect 2374 955 2380 956
rect 2462 960 2468 961
rect 2462 956 2463 960
rect 2467 956 2468 960
rect 2462 955 2468 956
rect 2558 960 2564 961
rect 2558 956 2559 960
rect 2563 956 2564 960
rect 2558 955 2564 956
rect 2662 960 2668 961
rect 2662 956 2663 960
rect 2667 956 2668 960
rect 2662 955 2668 956
rect 2774 960 2780 961
rect 2774 956 2775 960
rect 2779 956 2780 960
rect 2774 955 2780 956
rect 2902 960 2908 961
rect 2902 956 2903 960
rect 2907 956 2908 960
rect 2902 955 2908 956
rect 3046 960 3052 961
rect 3046 956 3047 960
rect 3051 956 3052 960
rect 3046 955 3052 956
rect 3198 960 3204 961
rect 3198 956 3199 960
rect 3203 956 3204 960
rect 3198 955 3204 956
rect 3358 960 3364 961
rect 3358 956 3359 960
rect 3363 956 3364 960
rect 3358 955 3364 956
rect 3502 960 3508 961
rect 3502 956 3503 960
rect 3507 956 3508 960
rect 3590 959 3591 963
rect 3595 959 3596 963
rect 3590 958 3596 959
rect 3502 955 3508 956
rect 2842 943 2848 944
rect 2842 939 2843 943
rect 2847 942 2848 943
rect 2919 943 2925 944
rect 2919 942 2920 943
rect 2847 940 2920 942
rect 2847 939 2848 940
rect 2842 938 2848 939
rect 2919 939 2920 940
rect 2924 939 2925 943
rect 2919 938 2925 939
rect 134 936 140 937
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 214 936 220 937
rect 214 932 215 936
rect 219 932 220 936
rect 214 931 220 932
rect 326 936 332 937
rect 326 932 327 936
rect 331 932 332 936
rect 326 931 332 932
rect 446 936 452 937
rect 446 932 447 936
rect 451 932 452 936
rect 446 931 452 932
rect 566 936 572 937
rect 566 932 567 936
rect 571 932 572 936
rect 566 931 572 932
rect 686 936 692 937
rect 686 932 687 936
rect 691 932 692 936
rect 686 931 692 932
rect 798 936 804 937
rect 798 932 799 936
rect 803 932 804 936
rect 798 931 804 932
rect 910 936 916 937
rect 910 932 911 936
rect 915 932 916 936
rect 910 931 916 932
rect 1014 936 1020 937
rect 1014 932 1015 936
rect 1019 932 1020 936
rect 1014 931 1020 932
rect 1118 936 1124 937
rect 1118 932 1119 936
rect 1123 932 1124 936
rect 1118 931 1124 932
rect 1222 936 1228 937
rect 1222 932 1223 936
rect 1227 932 1228 936
rect 1222 931 1228 932
rect 1326 936 1332 937
rect 1326 932 1327 936
rect 1331 932 1332 936
rect 1326 931 1332 932
rect 1830 933 1836 934
rect 110 928 116 929
rect 1830 929 1831 933
rect 1835 929 1836 933
rect 1830 928 1836 929
rect 202 927 208 928
rect 202 926 203 927
rect 197 924 203 926
rect 202 923 203 924
rect 207 923 208 927
rect 282 927 288 928
rect 282 926 283 927
rect 277 924 283 926
rect 202 922 208 923
rect 282 923 283 924
rect 287 923 288 927
rect 398 927 404 928
rect 398 926 399 927
rect 389 924 399 926
rect 282 922 288 923
rect 398 923 399 924
rect 403 923 404 927
rect 398 922 404 923
rect 426 927 432 928
rect 426 923 427 927
rect 431 926 432 927
rect 650 927 656 928
rect 650 926 651 927
rect 431 924 465 926
rect 629 924 651 926
rect 431 923 432 924
rect 426 922 432 923
rect 650 923 651 924
rect 655 923 656 927
rect 754 927 760 928
rect 754 926 755 927
rect 749 924 755 926
rect 650 922 656 923
rect 754 923 755 924
rect 759 923 760 927
rect 754 922 760 923
rect 791 927 797 928
rect 791 923 792 927
rect 796 926 797 927
rect 866 927 872 928
rect 796 924 817 926
rect 796 923 797 924
rect 791 922 797 923
rect 866 923 867 927
rect 871 926 872 927
rect 978 927 984 928
rect 871 924 929 926
rect 871 923 872 924
rect 866 922 872 923
rect 978 923 979 927
rect 983 926 984 927
rect 1082 927 1088 928
rect 983 924 1033 926
rect 983 923 984 924
rect 978 922 984 923
rect 1082 923 1083 927
rect 1087 926 1088 927
rect 1298 927 1304 928
rect 1298 926 1299 927
rect 1087 924 1137 926
rect 1285 924 1299 926
rect 1087 923 1088 924
rect 1082 922 1088 923
rect 1298 923 1299 924
rect 1303 923 1304 927
rect 1298 922 1304 923
rect 1194 919 1200 920
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 1194 915 1195 919
rect 1199 918 1200 919
rect 1344 918 1346 925
rect 1199 916 1346 918
rect 1830 916 1836 917
rect 1199 915 1200 916
rect 1194 914 1200 915
rect 110 911 116 912
rect 1830 912 1831 916
rect 1835 912 1836 916
rect 1830 911 1836 912
rect 2278 908 2284 909
rect 1870 905 1876 906
rect 1870 901 1871 905
rect 1875 901 1876 905
rect 2278 904 2279 908
rect 2283 904 2284 908
rect 2278 903 2284 904
rect 2358 908 2364 909
rect 2358 904 2359 908
rect 2363 904 2364 908
rect 2358 903 2364 904
rect 2438 908 2444 909
rect 2438 904 2439 908
rect 2443 904 2444 908
rect 2438 903 2444 904
rect 2518 908 2524 909
rect 2518 904 2519 908
rect 2523 904 2524 908
rect 2518 903 2524 904
rect 2606 908 2612 909
rect 2606 904 2607 908
rect 2611 904 2612 908
rect 2606 903 2612 904
rect 2702 908 2708 909
rect 2702 904 2703 908
rect 2707 904 2708 908
rect 2702 903 2708 904
rect 2806 908 2812 909
rect 2806 904 2807 908
rect 2811 904 2812 908
rect 2806 903 2812 904
rect 2910 908 2916 909
rect 2910 904 2911 908
rect 2915 904 2916 908
rect 2910 903 2916 904
rect 3014 908 3020 909
rect 3014 904 3015 908
rect 3019 904 3020 908
rect 3014 903 3020 904
rect 3110 908 3116 909
rect 3110 904 3111 908
rect 3115 904 3116 908
rect 3110 903 3116 904
rect 3214 908 3220 909
rect 3214 904 3215 908
rect 3219 904 3220 908
rect 3214 903 3220 904
rect 3318 908 3324 909
rect 3318 904 3319 908
rect 3323 904 3324 908
rect 3318 903 3324 904
rect 3422 908 3428 909
rect 3422 904 3423 908
rect 3427 904 3428 908
rect 3422 903 3428 904
rect 3502 908 3508 909
rect 3502 904 3503 908
rect 3507 904 3508 908
rect 3502 903 3508 904
rect 3590 905 3596 906
rect 1870 900 1876 901
rect 3590 901 3591 905
rect 3595 901 3596 905
rect 3590 900 3596 901
rect 2346 899 2352 900
rect 142 898 148 899
rect 142 894 143 898
rect 147 894 148 898
rect 142 893 148 894
rect 222 898 228 899
rect 222 894 223 898
rect 227 894 228 898
rect 222 893 228 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 454 898 460 899
rect 454 894 455 898
rect 459 894 460 898
rect 454 893 460 894
rect 574 898 580 899
rect 574 894 575 898
rect 579 894 580 898
rect 574 893 580 894
rect 694 898 700 899
rect 694 894 695 898
rect 699 894 700 898
rect 694 893 700 894
rect 806 898 812 899
rect 806 894 807 898
rect 811 894 812 898
rect 806 893 812 894
rect 918 898 924 899
rect 918 894 919 898
rect 923 894 924 898
rect 918 893 924 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1126 898 1132 899
rect 1126 894 1127 898
rect 1131 894 1132 898
rect 1126 893 1132 894
rect 1230 898 1236 899
rect 1230 894 1231 898
rect 1235 894 1236 898
rect 1230 893 1236 894
rect 1334 898 1340 899
rect 2346 898 2347 899
rect 1334 894 1335 898
rect 1339 894 1340 898
rect 2341 896 2347 898
rect 2346 895 2347 896
rect 2351 895 2352 899
rect 2430 899 2436 900
rect 2430 898 2431 899
rect 2421 896 2431 898
rect 2346 894 2352 895
rect 2430 895 2431 896
rect 2435 895 2436 899
rect 2506 899 2512 900
rect 2430 894 2436 895
rect 1334 893 1340 894
rect 2338 891 2344 892
rect 1870 888 1876 889
rect 166 887 173 888
rect 166 883 167 887
rect 172 883 173 887
rect 166 882 173 883
rect 202 887 208 888
rect 202 883 203 887
rect 207 886 208 887
rect 247 887 253 888
rect 247 886 248 887
rect 207 884 248 886
rect 207 883 208 884
rect 202 882 208 883
rect 247 883 248 884
rect 252 883 253 887
rect 247 882 253 883
rect 282 887 288 888
rect 282 883 283 887
rect 287 886 288 887
rect 359 887 365 888
rect 359 886 360 887
rect 287 884 360 886
rect 287 883 288 884
rect 282 882 288 883
rect 359 883 360 884
rect 364 883 365 887
rect 359 882 365 883
rect 398 887 404 888
rect 398 883 399 887
rect 403 886 404 887
rect 479 887 485 888
rect 479 886 480 887
rect 403 884 480 886
rect 403 883 404 884
rect 398 882 404 883
rect 479 883 480 884
rect 484 883 485 887
rect 479 882 485 883
rect 598 887 605 888
rect 598 883 599 887
rect 604 883 605 887
rect 598 882 605 883
rect 650 887 656 888
rect 650 883 651 887
rect 655 886 656 887
rect 719 887 725 888
rect 719 886 720 887
rect 655 884 720 886
rect 655 883 656 884
rect 650 882 656 883
rect 719 883 720 884
rect 724 883 725 887
rect 719 882 725 883
rect 831 887 837 888
rect 831 883 832 887
rect 836 886 837 887
rect 866 887 872 888
rect 866 886 867 887
rect 836 884 867 886
rect 836 883 837 884
rect 831 882 837 883
rect 866 883 867 884
rect 871 883 872 887
rect 866 882 872 883
rect 943 887 949 888
rect 943 883 944 887
rect 948 886 949 887
rect 978 887 984 888
rect 978 886 979 887
rect 948 884 979 886
rect 948 883 949 884
rect 943 882 949 883
rect 978 883 979 884
rect 983 883 984 887
rect 978 882 984 883
rect 1047 887 1053 888
rect 1047 883 1048 887
rect 1052 886 1053 887
rect 1082 887 1088 888
rect 1082 886 1083 887
rect 1052 884 1083 886
rect 1052 883 1053 884
rect 1047 882 1053 883
rect 1082 883 1083 884
rect 1087 883 1088 887
rect 1082 882 1088 883
rect 1151 887 1157 888
rect 1151 883 1152 887
rect 1156 886 1157 887
rect 1194 887 1200 888
rect 1194 886 1195 887
rect 1156 884 1195 886
rect 1156 883 1157 884
rect 1151 882 1157 883
rect 1194 883 1195 884
rect 1199 883 1200 887
rect 1194 882 1200 883
rect 1202 887 1208 888
rect 1202 883 1203 887
rect 1207 886 1208 887
rect 1255 887 1261 888
rect 1255 886 1256 887
rect 1207 884 1256 886
rect 1207 883 1208 884
rect 1202 882 1208 883
rect 1255 883 1256 884
rect 1260 883 1261 887
rect 1255 882 1261 883
rect 1298 887 1304 888
rect 1298 883 1299 887
rect 1303 886 1304 887
rect 1359 887 1365 888
rect 1359 886 1360 887
rect 1303 884 1360 886
rect 1303 883 1304 884
rect 1298 882 1304 883
rect 1359 883 1360 884
rect 1364 883 1365 887
rect 1870 884 1871 888
rect 1875 884 1876 888
rect 2338 887 2339 891
rect 2343 890 2344 891
rect 2456 890 2458 897
rect 2506 895 2507 899
rect 2511 898 2512 899
rect 2586 899 2592 900
rect 2511 896 2537 898
rect 2511 895 2512 896
rect 2506 894 2512 895
rect 2586 895 2587 899
rect 2591 898 2592 899
rect 2674 899 2680 900
rect 2591 896 2625 898
rect 2591 895 2592 896
rect 2586 894 2592 895
rect 2674 895 2675 899
rect 2679 898 2680 899
rect 2890 899 2896 900
rect 2890 898 2891 899
rect 2679 896 2721 898
rect 2869 896 2891 898
rect 2679 895 2680 896
rect 2674 894 2680 895
rect 2890 895 2891 896
rect 2895 895 2896 899
rect 3082 899 3088 900
rect 2920 896 2929 898
rect 2890 894 2896 895
rect 2918 895 2924 896
rect 2918 891 2919 895
rect 2923 891 2924 895
rect 3076 892 3078 897
rect 3082 895 3083 899
rect 3087 898 3088 899
rect 3178 899 3184 900
rect 3087 896 3129 898
rect 3087 895 3088 896
rect 3082 894 3088 895
rect 3178 895 3179 899
rect 3183 898 3184 899
rect 3282 899 3288 900
rect 3183 896 3233 898
rect 3183 895 3184 896
rect 3178 894 3184 895
rect 3282 895 3283 899
rect 3287 898 3288 899
rect 3490 899 3496 900
rect 3287 896 3337 898
rect 3287 895 3288 896
rect 3282 894 3288 895
rect 3484 892 3486 897
rect 3490 895 3491 899
rect 3495 898 3496 899
rect 3495 896 3521 898
rect 3495 895 3496 896
rect 3490 894 3496 895
rect 2918 890 2924 891
rect 3074 891 3080 892
rect 2343 888 2458 890
rect 2343 887 2344 888
rect 2338 886 2344 887
rect 3074 887 3075 891
rect 3079 887 3080 891
rect 3074 886 3080 887
rect 3482 891 3488 892
rect 3482 887 3483 891
rect 3487 887 3488 891
rect 3482 886 3488 887
rect 3590 888 3596 889
rect 1870 883 1876 884
rect 3590 884 3591 888
rect 3595 884 3596 888
rect 3590 883 3596 884
rect 1359 882 1365 883
rect 1286 875 1292 876
rect 1286 874 1287 875
rect 1159 872 1287 874
rect 1159 870 1161 872
rect 1286 871 1287 872
rect 1291 871 1292 875
rect 1286 870 1292 871
rect 2286 870 2292 871
rect 1100 868 1161 870
rect 167 867 173 868
rect 167 863 168 867
rect 172 866 173 867
rect 262 867 268 868
rect 262 866 263 867
rect 172 864 263 866
rect 172 863 173 864
rect 167 862 173 863
rect 262 863 263 864
rect 267 863 268 867
rect 262 862 268 863
rect 279 867 285 868
rect 279 863 280 867
rect 284 866 285 867
rect 406 867 412 868
rect 406 866 407 867
rect 284 864 407 866
rect 284 863 285 864
rect 279 862 285 863
rect 406 863 407 864
rect 411 863 412 867
rect 406 862 412 863
rect 423 867 432 868
rect 423 863 424 867
rect 431 863 432 867
rect 423 862 432 863
rect 583 867 589 868
rect 583 863 584 867
rect 588 866 589 867
rect 726 867 732 868
rect 726 866 727 867
rect 588 864 727 866
rect 588 863 589 864
rect 583 862 589 863
rect 726 863 727 864
rect 731 863 732 867
rect 726 862 732 863
rect 743 867 749 868
rect 743 863 744 867
rect 748 866 749 867
rect 878 867 884 868
rect 878 866 879 867
rect 748 864 879 866
rect 748 863 749 864
rect 743 862 749 863
rect 878 863 879 864
rect 883 863 884 867
rect 878 862 884 863
rect 886 867 892 868
rect 886 863 887 867
rect 891 866 892 867
rect 895 867 901 868
rect 895 866 896 867
rect 891 864 896 866
rect 891 863 892 864
rect 886 862 892 863
rect 895 863 896 864
rect 900 863 901 867
rect 895 862 901 863
rect 1039 867 1045 868
rect 1039 863 1040 867
rect 1044 866 1045 867
rect 1100 866 1102 868
rect 1175 867 1181 868
rect 1175 866 1176 867
rect 1044 864 1102 866
rect 1108 864 1176 866
rect 1044 863 1045 864
rect 1039 862 1045 863
rect 1106 863 1112 864
rect 1106 859 1107 863
rect 1111 859 1112 863
rect 1175 863 1176 864
rect 1180 863 1181 867
rect 1175 862 1181 863
rect 1303 867 1309 868
rect 1303 863 1304 867
rect 1308 866 1309 867
rect 1406 867 1412 868
rect 1406 866 1407 867
rect 1308 864 1407 866
rect 1308 863 1309 864
rect 1303 862 1309 863
rect 1406 863 1407 864
rect 1411 863 1412 867
rect 1406 862 1412 863
rect 1423 867 1429 868
rect 1423 863 1424 867
rect 1428 866 1429 867
rect 1526 867 1532 868
rect 1526 866 1527 867
rect 1428 864 1527 866
rect 1428 863 1429 864
rect 1423 862 1429 863
rect 1526 863 1527 864
rect 1531 863 1532 867
rect 1526 862 1532 863
rect 1543 867 1549 868
rect 1543 863 1544 867
rect 1548 866 1549 867
rect 1654 867 1660 868
rect 1654 866 1655 867
rect 1548 864 1655 866
rect 1548 863 1549 864
rect 1543 862 1549 863
rect 1654 863 1655 864
rect 1659 863 1660 867
rect 1654 862 1660 863
rect 1671 867 1677 868
rect 1671 863 1672 867
rect 1676 866 1677 867
rect 1710 867 1716 868
rect 1710 866 1711 867
rect 1676 864 1711 866
rect 1676 863 1677 864
rect 1671 862 1677 863
rect 1710 863 1711 864
rect 1715 863 1716 867
rect 2286 866 2287 870
rect 2291 866 2292 870
rect 2286 865 2292 866
rect 2366 870 2372 871
rect 2366 866 2367 870
rect 2371 866 2372 870
rect 2366 865 2372 866
rect 2446 870 2452 871
rect 2446 866 2447 870
rect 2451 866 2452 870
rect 2446 865 2452 866
rect 2526 870 2532 871
rect 2526 866 2527 870
rect 2531 866 2532 870
rect 2526 865 2532 866
rect 2614 870 2620 871
rect 2614 866 2615 870
rect 2619 866 2620 870
rect 2614 865 2620 866
rect 2710 870 2716 871
rect 2710 866 2711 870
rect 2715 866 2716 870
rect 2710 865 2716 866
rect 2814 870 2820 871
rect 2814 866 2815 870
rect 2819 866 2820 870
rect 2814 865 2820 866
rect 2918 870 2924 871
rect 2918 866 2919 870
rect 2923 866 2924 870
rect 2918 865 2924 866
rect 3022 870 3028 871
rect 3022 866 3023 870
rect 3027 866 3028 870
rect 3022 865 3028 866
rect 3118 870 3124 871
rect 3118 866 3119 870
rect 3123 866 3124 870
rect 3118 865 3124 866
rect 3222 870 3228 871
rect 3222 866 3223 870
rect 3227 866 3228 870
rect 3222 865 3228 866
rect 3326 870 3332 871
rect 3326 866 3327 870
rect 3331 866 3332 870
rect 3326 865 3332 866
rect 3430 870 3436 871
rect 3430 866 3431 870
rect 3435 866 3436 870
rect 3430 865 3436 866
rect 3510 870 3516 871
rect 3510 866 3511 870
rect 3515 866 3516 870
rect 3510 865 3516 866
rect 1710 862 1716 863
rect 2311 859 2317 860
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 254 858 260 859
rect 254 854 255 858
rect 259 854 260 858
rect 254 853 260 854
rect 398 858 404 859
rect 398 854 399 858
rect 403 854 404 858
rect 398 853 404 854
rect 558 858 564 859
rect 558 854 559 858
rect 563 854 564 858
rect 558 853 564 854
rect 718 858 724 859
rect 718 854 719 858
rect 723 854 724 858
rect 718 853 724 854
rect 870 858 876 859
rect 870 854 871 858
rect 875 854 876 858
rect 870 853 876 854
rect 1014 858 1020 859
rect 1106 858 1112 859
rect 1150 858 1156 859
rect 1014 854 1015 858
rect 1019 854 1020 858
rect 1014 853 1020 854
rect 1150 854 1151 858
rect 1155 854 1156 858
rect 1150 853 1156 854
rect 1278 858 1284 859
rect 1278 854 1279 858
rect 1283 854 1284 858
rect 1278 853 1284 854
rect 1398 858 1404 859
rect 1398 854 1399 858
rect 1403 854 1404 858
rect 1398 853 1404 854
rect 1518 858 1524 859
rect 1518 854 1519 858
rect 1523 854 1524 858
rect 1518 853 1524 854
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 2311 855 2312 859
rect 2316 858 2317 859
rect 2338 859 2344 860
rect 2338 858 2339 859
rect 2316 856 2339 858
rect 2316 855 2317 856
rect 2311 854 2317 855
rect 2338 855 2339 856
rect 2343 855 2344 859
rect 2338 854 2344 855
rect 2346 859 2352 860
rect 2346 855 2347 859
rect 2351 858 2352 859
rect 2391 859 2397 860
rect 2391 858 2392 859
rect 2351 856 2392 858
rect 2351 855 2352 856
rect 2346 854 2352 855
rect 2391 855 2392 856
rect 2396 855 2397 859
rect 2391 854 2397 855
rect 2471 859 2477 860
rect 2471 855 2472 859
rect 2476 858 2477 859
rect 2506 859 2512 860
rect 2506 858 2507 859
rect 2476 856 2507 858
rect 2476 855 2477 856
rect 2471 854 2477 855
rect 2506 855 2507 856
rect 2511 855 2512 859
rect 2506 854 2512 855
rect 2551 859 2557 860
rect 2551 855 2552 859
rect 2556 858 2557 859
rect 2586 859 2592 860
rect 2586 858 2587 859
rect 2556 856 2587 858
rect 2556 855 2557 856
rect 2551 854 2557 855
rect 2586 855 2587 856
rect 2591 855 2592 859
rect 2586 854 2592 855
rect 2639 859 2645 860
rect 2639 855 2640 859
rect 2644 858 2645 859
rect 2674 859 2680 860
rect 2674 858 2675 859
rect 2644 856 2675 858
rect 2644 855 2645 856
rect 2639 854 2645 855
rect 2674 855 2675 856
rect 2679 855 2680 859
rect 2674 854 2680 855
rect 2722 859 2728 860
rect 2722 855 2723 859
rect 2727 858 2728 859
rect 2735 859 2741 860
rect 2735 858 2736 859
rect 2727 856 2736 858
rect 2727 855 2728 856
rect 2722 854 2728 855
rect 2735 855 2736 856
rect 2740 855 2741 859
rect 2735 854 2741 855
rect 2839 859 2848 860
rect 2839 855 2840 859
rect 2847 855 2848 859
rect 2839 854 2848 855
rect 2890 859 2896 860
rect 2890 855 2891 859
rect 2895 858 2896 859
rect 2943 859 2949 860
rect 2943 858 2944 859
rect 2895 856 2944 858
rect 2895 855 2896 856
rect 2890 854 2896 855
rect 2943 855 2944 856
rect 2948 855 2949 859
rect 2943 854 2949 855
rect 3047 859 3053 860
rect 3047 855 3048 859
rect 3052 858 3053 859
rect 3082 859 3088 860
rect 3082 858 3083 859
rect 3052 856 3083 858
rect 3052 855 3053 856
rect 3047 854 3053 855
rect 3082 855 3083 856
rect 3087 855 3088 859
rect 3082 854 3088 855
rect 3143 859 3149 860
rect 3143 855 3144 859
rect 3148 858 3149 859
rect 3178 859 3184 860
rect 3178 858 3179 859
rect 3148 856 3179 858
rect 3148 855 3149 856
rect 3143 854 3149 855
rect 3178 855 3179 856
rect 3183 855 3184 859
rect 3178 854 3184 855
rect 3247 859 3253 860
rect 3247 855 3248 859
rect 3252 858 3253 859
rect 3282 859 3288 860
rect 3282 858 3283 859
rect 3252 856 3283 858
rect 3252 855 3253 856
rect 3247 854 3253 855
rect 3282 855 3283 856
rect 3287 855 3288 859
rect 3282 854 3288 855
rect 3351 859 3357 860
rect 3351 855 3352 859
rect 3356 858 3357 859
rect 3414 859 3420 860
rect 3414 858 3415 859
rect 3356 856 3415 858
rect 3356 855 3357 856
rect 3351 854 3357 855
rect 3414 855 3415 856
rect 3419 855 3420 859
rect 3414 854 3420 855
rect 3455 859 3461 860
rect 3455 855 3456 859
rect 3460 858 3461 859
rect 3490 859 3496 860
rect 3490 858 3491 859
rect 3460 856 3491 858
rect 3460 855 3461 856
rect 3455 854 3461 855
rect 3490 855 3491 856
rect 3495 855 3496 859
rect 3490 854 3496 855
rect 3534 859 3541 860
rect 3534 855 3535 859
rect 3540 855 3541 859
rect 3534 854 3541 855
rect 1646 853 1652 854
rect 2334 843 2340 844
rect 2334 842 2335 843
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 2212 840 2335 842
rect 1830 835 1836 836
rect 2191 835 2197 836
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 262 831 268 832
rect 262 827 263 831
rect 267 827 268 831
rect 262 826 268 827
rect 406 831 412 832
rect 406 827 407 831
rect 411 827 412 831
rect 406 826 412 827
rect 598 831 604 832
rect 598 827 599 831
rect 603 827 604 831
rect 598 826 604 827
rect 726 831 732 832
rect 726 827 727 831
rect 731 827 732 831
rect 726 826 732 827
rect 878 831 884 832
rect 878 827 879 831
rect 883 827 884 831
rect 1106 831 1112 832
rect 1106 830 1107 831
rect 1069 828 1107 830
rect 878 826 884 827
rect 1106 827 1107 828
rect 1111 827 1112 831
rect 1106 826 1112 827
rect 1202 831 1208 832
rect 1202 827 1203 831
rect 1207 827 1208 831
rect 1202 826 1208 827
rect 1286 831 1292 832
rect 1286 827 1287 831
rect 1291 827 1292 831
rect 1286 826 1292 827
rect 1406 831 1412 832
rect 1406 827 1407 831
rect 1411 827 1412 831
rect 1406 826 1412 827
rect 1526 831 1532 832
rect 1526 827 1527 831
rect 1531 827 1532 831
rect 1526 826 1532 827
rect 1654 831 1660 832
rect 1654 827 1655 831
rect 1659 827 1660 831
rect 2191 831 2192 835
rect 2196 834 2197 835
rect 2212 834 2214 840
rect 2334 839 2335 840
rect 2339 839 2340 843
rect 2662 843 2668 844
rect 2662 842 2663 843
rect 2334 838 2340 839
rect 2424 840 2663 842
rect 2196 832 2214 834
rect 2218 835 2224 836
rect 2196 831 2197 832
rect 2191 830 2197 831
rect 2218 831 2219 835
rect 2223 834 2224 835
rect 2271 835 2277 836
rect 2271 834 2272 835
rect 2223 832 2272 834
rect 2223 831 2224 832
rect 2218 830 2224 831
rect 2271 831 2272 832
rect 2276 831 2277 835
rect 2271 830 2277 831
rect 2351 835 2357 836
rect 2351 831 2352 835
rect 2356 834 2357 835
rect 2424 834 2426 840
rect 2662 839 2663 840
rect 2667 839 2668 843
rect 2662 838 2668 839
rect 2356 832 2426 834
rect 2430 835 2436 836
rect 2356 831 2357 832
rect 2351 830 2357 831
rect 2430 831 2431 835
rect 2435 834 2436 835
rect 2447 835 2453 836
rect 2447 834 2448 835
rect 2435 832 2448 834
rect 2435 831 2436 832
rect 2430 830 2436 831
rect 2447 831 2448 832
rect 2452 831 2453 835
rect 2447 830 2453 831
rect 2474 835 2480 836
rect 2474 831 2475 835
rect 2479 834 2480 835
rect 2559 835 2565 836
rect 2559 834 2560 835
rect 2479 832 2560 834
rect 2479 831 2480 832
rect 2474 830 2480 831
rect 2559 831 2560 832
rect 2564 831 2565 835
rect 2559 830 2565 831
rect 2586 835 2592 836
rect 2586 831 2587 835
rect 2591 834 2592 835
rect 2679 835 2685 836
rect 2679 834 2680 835
rect 2591 832 2680 834
rect 2591 831 2592 832
rect 2586 830 2592 831
rect 2679 831 2680 832
rect 2684 831 2685 835
rect 2679 830 2685 831
rect 2807 835 2813 836
rect 2807 831 2808 835
rect 2812 834 2813 835
rect 2858 835 2864 836
rect 2858 834 2859 835
rect 2812 832 2859 834
rect 2812 831 2813 832
rect 2807 830 2813 831
rect 2858 831 2859 832
rect 2863 831 2864 835
rect 2858 830 2864 831
rect 2926 835 2932 836
rect 2926 831 2927 835
rect 2931 834 2932 835
rect 2935 835 2941 836
rect 2935 834 2936 835
rect 2931 832 2936 834
rect 2931 831 2932 832
rect 2926 830 2932 831
rect 2935 831 2936 832
rect 2940 831 2941 835
rect 2935 830 2941 831
rect 3054 835 3060 836
rect 3054 831 3055 835
rect 3059 834 3060 835
rect 3063 835 3069 836
rect 3063 834 3064 835
rect 3059 832 3064 834
rect 3059 831 3060 832
rect 3054 830 3060 831
rect 3063 831 3064 832
rect 3068 831 3069 835
rect 3063 830 3069 831
rect 3090 835 3096 836
rect 3090 831 3091 835
rect 3095 834 3096 835
rect 3183 835 3189 836
rect 3183 834 3184 835
rect 3095 832 3184 834
rect 3095 831 3096 832
rect 3090 830 3096 831
rect 3183 831 3184 832
rect 3188 831 3189 835
rect 3183 830 3189 831
rect 3210 835 3216 836
rect 3210 831 3211 835
rect 3215 834 3216 835
rect 3303 835 3309 836
rect 3303 834 3304 835
rect 3215 832 3304 834
rect 3215 831 3216 832
rect 3210 830 3216 831
rect 3303 831 3304 832
rect 3308 831 3309 835
rect 3303 830 3309 831
rect 3394 835 3400 836
rect 3394 831 3395 835
rect 3399 834 3400 835
rect 3431 835 3437 836
rect 3431 834 3432 835
rect 3399 832 3432 834
rect 3399 831 3400 832
rect 3394 830 3400 831
rect 3431 831 3432 832
rect 3436 831 3437 835
rect 3431 830 3437 831
rect 3482 835 3488 836
rect 3482 831 3483 835
rect 3487 834 3488 835
rect 3535 835 3541 836
rect 3535 834 3536 835
rect 3487 832 3536 834
rect 3487 831 3488 832
rect 3482 830 3488 831
rect 3535 831 3536 832
rect 3540 831 3541 835
rect 3535 830 3541 831
rect 1654 826 1660 827
rect 2166 826 2172 827
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 1830 823 1836 824
rect 110 818 116 819
rect 134 820 140 821
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 246 820 252 821
rect 246 816 247 820
rect 251 816 252 820
rect 246 815 252 816
rect 390 820 396 821
rect 390 816 391 820
rect 395 816 396 820
rect 390 815 396 816
rect 550 820 556 821
rect 550 816 551 820
rect 555 816 556 820
rect 550 815 556 816
rect 710 820 716 821
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 1006 820 1012 821
rect 1006 816 1007 820
rect 1011 816 1012 820
rect 1006 815 1012 816
rect 1142 820 1148 821
rect 1142 816 1143 820
rect 1147 816 1148 820
rect 1142 815 1148 816
rect 1270 820 1276 821
rect 1270 816 1271 820
rect 1275 816 1276 820
rect 1270 815 1276 816
rect 1390 820 1396 821
rect 1390 816 1391 820
rect 1395 816 1396 820
rect 1390 815 1396 816
rect 1510 820 1516 821
rect 1510 816 1511 820
rect 1515 816 1516 820
rect 1510 815 1516 816
rect 1638 820 1644 821
rect 1638 816 1639 820
rect 1643 816 1644 820
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 2166 822 2167 826
rect 2171 822 2172 826
rect 2166 821 2172 822
rect 2246 826 2252 827
rect 2246 822 2247 826
rect 2251 822 2252 826
rect 2246 821 2252 822
rect 2326 826 2332 827
rect 2326 822 2327 826
rect 2331 822 2332 826
rect 2326 821 2332 822
rect 2422 826 2428 827
rect 2422 822 2423 826
rect 2427 822 2428 826
rect 2422 821 2428 822
rect 2534 826 2540 827
rect 2534 822 2535 826
rect 2539 822 2540 826
rect 2534 821 2540 822
rect 2654 826 2660 827
rect 2654 822 2655 826
rect 2659 822 2660 826
rect 2654 821 2660 822
rect 2782 826 2788 827
rect 2782 822 2783 826
rect 2787 822 2788 826
rect 2782 821 2788 822
rect 2910 826 2916 827
rect 2910 822 2911 826
rect 2915 822 2916 826
rect 2910 821 2916 822
rect 3038 826 3044 827
rect 3038 822 3039 826
rect 3043 822 3044 826
rect 3038 821 3044 822
rect 3158 826 3164 827
rect 3158 822 3159 826
rect 3163 822 3164 826
rect 3158 821 3164 822
rect 3278 826 3284 827
rect 3278 822 3279 826
rect 3283 822 3284 826
rect 3278 821 3284 822
rect 3406 826 3412 827
rect 3406 822 3407 826
rect 3411 822 3412 826
rect 3406 821 3412 822
rect 3510 826 3516 827
rect 3510 822 3511 826
rect 3515 822 3516 826
rect 3510 821 3516 822
rect 1830 818 1836 819
rect 1638 815 1644 816
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 3590 808 3596 809
rect 3590 804 3591 808
rect 3595 804 3596 808
rect 3590 803 3596 804
rect 2218 799 2224 800
rect 2218 795 2219 799
rect 2223 795 2224 799
rect 2218 794 2224 795
rect 2298 799 2304 800
rect 2298 795 2299 799
rect 2303 795 2304 799
rect 2298 794 2304 795
rect 2334 799 2340 800
rect 2334 795 2335 799
rect 2339 795 2340 799
rect 2334 794 2340 795
rect 2474 799 2480 800
rect 2474 795 2475 799
rect 2479 795 2480 799
rect 2474 794 2480 795
rect 2586 799 2592 800
rect 2586 795 2587 799
rect 2591 795 2592 799
rect 2586 794 2592 795
rect 2662 799 2668 800
rect 2662 795 2663 799
rect 2667 795 2668 799
rect 2662 794 2668 795
rect 2834 799 2840 800
rect 2834 795 2835 799
rect 2839 795 2840 799
rect 2834 794 2840 795
rect 2858 799 2864 800
rect 2858 795 2859 799
rect 2863 798 2864 799
rect 3090 799 3096 800
rect 2863 796 2921 798
rect 2863 795 2864 796
rect 2858 794 2864 795
rect 3090 795 3091 799
rect 3095 795 3096 799
rect 3090 794 3096 795
rect 3210 799 3216 800
rect 3210 795 3211 799
rect 3215 795 3216 799
rect 3394 799 3400 800
rect 3394 798 3395 799
rect 3333 796 3395 798
rect 3210 794 3216 795
rect 3394 795 3395 796
rect 3399 795 3400 799
rect 3394 794 3400 795
rect 3414 799 3420 800
rect 3414 795 3415 799
rect 3419 795 3420 799
rect 3414 794 3420 795
rect 3534 799 3540 800
rect 3534 795 3535 799
rect 3539 795 3540 799
rect 3534 794 3540 795
rect 1870 791 1876 792
rect 1870 787 1871 791
rect 1875 787 1876 791
rect 3590 791 3596 792
rect 1870 786 1876 787
rect 2158 788 2164 789
rect 2158 784 2159 788
rect 2163 784 2164 788
rect 2158 783 2164 784
rect 2238 788 2244 789
rect 2238 784 2239 788
rect 2243 784 2244 788
rect 2238 783 2244 784
rect 2318 788 2324 789
rect 2318 784 2319 788
rect 2323 784 2324 788
rect 2318 783 2324 784
rect 2414 788 2420 789
rect 2414 784 2415 788
rect 2419 784 2420 788
rect 2414 783 2420 784
rect 2526 788 2532 789
rect 2526 784 2527 788
rect 2531 784 2532 788
rect 2526 783 2532 784
rect 2646 788 2652 789
rect 2646 784 2647 788
rect 2651 784 2652 788
rect 2646 783 2652 784
rect 2774 788 2780 789
rect 2774 784 2775 788
rect 2779 784 2780 788
rect 2774 783 2780 784
rect 2902 788 2908 789
rect 2902 784 2903 788
rect 2907 784 2908 788
rect 2902 783 2908 784
rect 3030 788 3036 789
rect 3030 784 3031 788
rect 3035 784 3036 788
rect 3030 783 3036 784
rect 3150 788 3156 789
rect 3150 784 3151 788
rect 3155 784 3156 788
rect 3150 783 3156 784
rect 3270 788 3276 789
rect 3270 784 3271 788
rect 3275 784 3276 788
rect 3270 783 3276 784
rect 3398 788 3404 789
rect 3398 784 3399 788
rect 3403 784 3404 788
rect 3398 783 3404 784
rect 3502 788 3508 789
rect 3502 784 3503 788
rect 3507 784 3508 788
rect 3590 787 3591 791
rect 3595 787 3596 791
rect 3590 786 3596 787
rect 3502 783 3508 784
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 262 764 268 765
rect 262 760 263 764
rect 267 760 268 764
rect 262 759 268 760
rect 430 764 436 765
rect 430 760 431 764
rect 435 760 436 764
rect 430 759 436 760
rect 606 764 612 765
rect 606 760 607 764
rect 611 760 612 764
rect 606 759 612 760
rect 782 764 788 765
rect 782 760 783 764
rect 787 760 788 764
rect 782 759 788 760
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1102 764 1108 765
rect 1102 760 1103 764
rect 1107 760 1108 764
rect 1102 759 1108 760
rect 1246 764 1252 765
rect 1246 760 1247 764
rect 1251 760 1252 764
rect 1246 759 1252 760
rect 1382 764 1388 765
rect 1382 760 1383 764
rect 1387 760 1388 764
rect 1382 759 1388 760
rect 1510 764 1516 765
rect 1510 760 1511 764
rect 1515 760 1516 764
rect 1510 759 1516 760
rect 1638 764 1644 765
rect 1638 760 1639 764
rect 1643 760 1644 764
rect 1638 759 1644 760
rect 1742 764 1748 765
rect 1742 760 1743 764
rect 1747 760 1748 764
rect 1742 759 1748 760
rect 1830 761 1836 762
rect 110 756 116 757
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1830 756 1836 757
rect 218 755 224 756
rect 218 754 219 755
rect 197 752 219 754
rect 218 751 219 752
rect 223 751 224 755
rect 330 755 336 756
rect 330 754 331 755
rect 325 752 331 754
rect 218 750 224 751
rect 330 751 331 752
rect 335 751 336 755
rect 535 755 541 756
rect 535 754 536 755
rect 493 752 536 754
rect 330 750 336 751
rect 535 751 536 752
rect 540 751 541 755
rect 850 755 856 756
rect 535 750 541 751
rect 322 747 328 748
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 322 743 323 747
rect 327 746 328 747
rect 624 746 626 753
rect 327 744 626 746
rect 844 746 846 753
rect 850 751 851 755
rect 855 754 856 755
rect 1210 755 1216 756
rect 1210 754 1211 755
rect 855 752 969 754
rect 1165 752 1211 754
rect 855 751 856 752
rect 850 750 856 751
rect 1210 751 1211 752
rect 1215 751 1216 755
rect 1338 755 1344 756
rect 1338 754 1339 755
rect 1309 752 1339 754
rect 1210 750 1216 751
rect 1338 751 1339 752
rect 1343 751 1344 755
rect 1470 755 1476 756
rect 1470 754 1471 755
rect 1445 752 1471 754
rect 1338 750 1344 751
rect 1470 751 1471 752
rect 1475 751 1476 755
rect 1598 755 1604 756
rect 1598 754 1599 755
rect 1573 752 1599 754
rect 1470 750 1476 751
rect 1598 751 1599 752
rect 1603 751 1604 755
rect 1710 755 1716 756
rect 1598 750 1604 751
rect 1700 748 1702 753
rect 1710 751 1711 755
rect 1715 754 1716 755
rect 1715 752 1761 754
rect 1715 751 1716 752
rect 1710 750 1716 751
rect 886 747 892 748
rect 886 746 887 747
rect 844 744 887 746
rect 327 743 328 744
rect 322 742 328 743
rect 886 743 887 744
rect 891 743 892 747
rect 886 742 892 743
rect 1698 747 1704 748
rect 1698 743 1699 747
rect 1703 743 1704 747
rect 1698 742 1704 743
rect 1830 744 1836 745
rect 110 739 116 740
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1894 736 1900 737
rect 1870 733 1876 734
rect 1870 729 1871 733
rect 1875 729 1876 733
rect 1894 732 1895 736
rect 1899 732 1900 736
rect 1894 731 1900 732
rect 1974 736 1980 737
rect 1974 732 1975 736
rect 1979 732 1980 736
rect 1974 731 1980 732
rect 2070 736 2076 737
rect 2070 732 2071 736
rect 2075 732 2076 736
rect 2070 731 2076 732
rect 2182 736 2188 737
rect 2182 732 2183 736
rect 2187 732 2188 736
rect 2182 731 2188 732
rect 2310 736 2316 737
rect 2310 732 2311 736
rect 2315 732 2316 736
rect 2310 731 2316 732
rect 2446 736 2452 737
rect 2446 732 2447 736
rect 2451 732 2452 736
rect 2446 731 2452 732
rect 2590 736 2596 737
rect 2590 732 2591 736
rect 2595 732 2596 736
rect 2590 731 2596 732
rect 2742 736 2748 737
rect 2742 732 2743 736
rect 2747 732 2748 736
rect 2742 731 2748 732
rect 2894 736 2900 737
rect 2894 732 2895 736
rect 2899 732 2900 736
rect 2894 731 2900 732
rect 3046 736 3052 737
rect 3046 732 3047 736
rect 3051 732 3052 736
rect 3046 731 3052 732
rect 3198 736 3204 737
rect 3198 732 3199 736
rect 3203 732 3204 736
rect 3198 731 3204 732
rect 3358 736 3364 737
rect 3358 732 3359 736
rect 3363 732 3364 736
rect 3358 731 3364 732
rect 3502 736 3508 737
rect 3502 732 3503 736
rect 3507 732 3508 736
rect 3502 731 3508 732
rect 3590 733 3596 734
rect 1870 728 1876 729
rect 3590 729 3591 733
rect 3595 729 3596 733
rect 3590 728 3596 729
rect 2050 727 2056 728
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 270 726 276 727
rect 270 722 271 726
rect 275 722 276 726
rect 270 721 276 722
rect 438 726 444 727
rect 438 722 439 726
rect 443 722 444 726
rect 438 721 444 722
rect 614 726 620 727
rect 614 722 615 726
rect 619 722 620 726
rect 614 721 620 722
rect 790 726 796 727
rect 790 722 791 726
rect 795 722 796 726
rect 790 721 796 722
rect 958 726 964 727
rect 958 722 959 726
rect 963 722 964 726
rect 958 721 964 722
rect 1110 726 1116 727
rect 1110 722 1111 726
rect 1115 722 1116 726
rect 1110 721 1116 722
rect 1254 726 1260 727
rect 1254 722 1255 726
rect 1259 722 1260 726
rect 1254 721 1260 722
rect 1390 726 1396 727
rect 1390 722 1391 726
rect 1395 722 1396 726
rect 1390 721 1396 722
rect 1518 726 1524 727
rect 1518 722 1519 726
rect 1523 722 1524 726
rect 1518 721 1524 722
rect 1646 726 1652 727
rect 1646 722 1647 726
rect 1651 722 1652 726
rect 1646 721 1652 722
rect 1750 726 1756 727
rect 2050 726 2051 727
rect 1750 722 1751 726
rect 1755 722 1756 726
rect 1750 721 1756 722
rect 1956 722 1958 725
rect 2037 724 2051 726
rect 1970 723 1976 724
rect 1970 722 1971 723
rect 1956 720 1971 722
rect 1970 719 1971 720
rect 1975 719 1976 723
rect 2050 723 2051 724
rect 2055 723 2056 727
rect 2138 727 2144 728
rect 2050 722 2056 723
rect 2132 720 2134 725
rect 2138 723 2139 727
rect 2143 726 2144 727
rect 2402 727 2408 728
rect 2402 726 2403 727
rect 2143 724 2201 726
rect 2373 724 2403 726
rect 2143 723 2144 724
rect 2138 722 2144 723
rect 2402 723 2403 724
rect 2407 723 2408 727
rect 2514 727 2520 728
rect 2402 722 2408 723
rect 1970 718 1976 719
rect 2130 719 2136 720
rect 1870 716 1876 717
rect 166 715 173 716
rect 166 711 167 715
rect 172 711 173 715
rect 166 710 173 711
rect 218 715 224 716
rect 218 711 219 715
rect 223 714 224 715
rect 295 715 301 716
rect 295 714 296 715
rect 223 712 296 714
rect 223 711 224 712
rect 218 710 224 711
rect 295 711 296 712
rect 300 711 301 715
rect 295 710 301 711
rect 330 715 336 716
rect 330 711 331 715
rect 335 714 336 715
rect 463 715 469 716
rect 463 714 464 715
rect 335 712 464 714
rect 335 711 336 712
rect 330 710 336 711
rect 463 711 464 712
rect 468 711 469 715
rect 463 710 469 711
rect 535 715 541 716
rect 535 711 536 715
rect 540 714 541 715
rect 639 715 645 716
rect 639 714 640 715
rect 540 712 640 714
rect 540 711 541 712
rect 535 710 541 711
rect 639 711 640 712
rect 644 711 645 715
rect 639 710 645 711
rect 815 715 821 716
rect 815 711 816 715
rect 820 714 821 715
rect 850 715 856 716
rect 850 714 851 715
rect 820 712 851 714
rect 820 711 821 712
rect 815 710 821 711
rect 850 711 851 712
rect 855 711 856 715
rect 850 710 856 711
rect 966 715 972 716
rect 966 711 967 715
rect 971 714 972 715
rect 983 715 989 716
rect 983 714 984 715
rect 971 712 984 714
rect 971 711 972 712
rect 966 710 972 711
rect 983 711 984 712
rect 988 711 989 715
rect 983 710 989 711
rect 1135 715 1141 716
rect 1135 711 1136 715
rect 1140 714 1141 715
rect 1198 715 1204 716
rect 1198 714 1199 715
rect 1140 712 1199 714
rect 1140 711 1141 712
rect 1135 710 1141 711
rect 1198 711 1199 712
rect 1203 711 1204 715
rect 1198 710 1204 711
rect 1210 715 1216 716
rect 1210 711 1211 715
rect 1215 714 1216 715
rect 1279 715 1285 716
rect 1279 714 1280 715
rect 1215 712 1280 714
rect 1215 711 1216 712
rect 1210 710 1216 711
rect 1279 711 1280 712
rect 1284 711 1285 715
rect 1279 710 1285 711
rect 1338 715 1344 716
rect 1338 711 1339 715
rect 1343 714 1344 715
rect 1415 715 1421 716
rect 1415 714 1416 715
rect 1343 712 1416 714
rect 1343 711 1344 712
rect 1338 710 1344 711
rect 1415 711 1416 712
rect 1420 711 1421 715
rect 1415 710 1421 711
rect 1470 715 1476 716
rect 1470 711 1471 715
rect 1475 714 1476 715
rect 1543 715 1549 716
rect 1543 714 1544 715
rect 1475 712 1544 714
rect 1475 711 1476 712
rect 1470 710 1476 711
rect 1543 711 1544 712
rect 1548 711 1549 715
rect 1543 710 1549 711
rect 1598 715 1604 716
rect 1598 711 1599 715
rect 1603 714 1604 715
rect 1671 715 1677 716
rect 1671 714 1672 715
rect 1603 712 1672 714
rect 1603 711 1604 712
rect 1598 710 1604 711
rect 1671 711 1672 712
rect 1676 711 1677 715
rect 1671 710 1677 711
rect 1698 715 1704 716
rect 1698 711 1699 715
rect 1703 714 1704 715
rect 1775 715 1781 716
rect 1775 714 1776 715
rect 1703 712 1776 714
rect 1703 711 1704 712
rect 1698 710 1704 711
rect 1775 711 1776 712
rect 1780 711 1781 715
rect 1870 712 1871 716
rect 1875 712 1876 716
rect 2130 715 2131 719
rect 2135 715 2136 719
rect 2130 714 2136 715
rect 2262 719 2268 720
rect 2262 715 2263 719
rect 2267 718 2268 719
rect 2464 718 2466 725
rect 2514 723 2515 727
rect 2519 726 2520 727
rect 2658 727 2664 728
rect 2519 724 2609 726
rect 2519 723 2520 724
rect 2514 722 2520 723
rect 2658 723 2659 727
rect 2663 726 2664 727
rect 2810 727 2816 728
rect 2663 724 2761 726
rect 2663 723 2664 724
rect 2658 722 2664 723
rect 2810 723 2811 727
rect 2815 726 2816 727
rect 3114 727 3120 728
rect 2815 724 2913 726
rect 2815 723 2816 724
rect 2810 722 2816 723
rect 3054 723 3060 724
rect 3054 719 3055 723
rect 3059 722 3060 723
rect 3064 722 3066 725
rect 3114 723 3115 727
rect 3119 726 3120 727
rect 3266 727 3272 728
rect 3119 724 3217 726
rect 3119 723 3120 724
rect 3114 722 3120 723
rect 3266 723 3267 727
rect 3271 726 3272 727
rect 3271 724 3377 726
rect 3271 723 3272 724
rect 3266 722 3272 723
rect 3059 720 3066 722
rect 3564 720 3566 725
rect 3059 719 3060 720
rect 3054 718 3060 719
rect 3562 719 3568 720
rect 2267 716 2466 718
rect 2267 715 2268 716
rect 2262 714 2268 715
rect 3562 715 3563 719
rect 3567 715 3568 719
rect 3562 714 3568 715
rect 3590 716 3596 717
rect 1870 711 1876 712
rect 3590 712 3591 716
rect 3595 712 3596 716
rect 3590 711 3596 712
rect 1775 710 1781 711
rect 1902 698 1908 699
rect 1902 694 1903 698
rect 1907 694 1908 698
rect 1902 693 1908 694
rect 1982 698 1988 699
rect 1982 694 1983 698
rect 1987 694 1988 698
rect 1982 693 1988 694
rect 2078 698 2084 699
rect 2078 694 2079 698
rect 2083 694 2084 698
rect 2078 693 2084 694
rect 2190 698 2196 699
rect 2190 694 2191 698
rect 2195 694 2196 698
rect 2190 693 2196 694
rect 2318 698 2324 699
rect 2318 694 2319 698
rect 2323 694 2324 698
rect 2318 693 2324 694
rect 2454 698 2460 699
rect 2454 694 2455 698
rect 2459 694 2460 698
rect 2454 693 2460 694
rect 2598 698 2604 699
rect 2598 694 2599 698
rect 2603 694 2604 698
rect 2598 693 2604 694
rect 2750 698 2756 699
rect 2750 694 2751 698
rect 2755 694 2756 698
rect 2750 693 2756 694
rect 2902 698 2908 699
rect 2902 694 2903 698
rect 2907 694 2908 698
rect 2902 693 2908 694
rect 3054 698 3060 699
rect 3054 694 3055 698
rect 3059 694 3060 698
rect 3054 693 3060 694
rect 3206 698 3212 699
rect 3206 694 3207 698
rect 3211 694 3212 698
rect 3206 693 3212 694
rect 3366 698 3372 699
rect 3366 694 3367 698
rect 3371 694 3372 698
rect 3366 693 3372 694
rect 3510 698 3516 699
rect 3510 694 3511 698
rect 3515 694 3516 698
rect 3510 693 3516 694
rect 319 691 328 692
rect 319 687 320 691
rect 327 687 328 691
rect 319 686 328 687
rect 346 691 352 692
rect 346 687 347 691
rect 351 690 352 691
rect 431 691 437 692
rect 431 690 432 691
rect 351 688 432 690
rect 351 687 352 688
rect 346 686 352 687
rect 431 687 432 688
rect 436 687 437 691
rect 431 686 437 687
rect 458 691 464 692
rect 458 687 459 691
rect 463 690 464 691
rect 551 691 557 692
rect 551 690 552 691
rect 463 688 552 690
rect 463 687 464 688
rect 458 686 464 687
rect 551 687 552 688
rect 556 687 557 691
rect 551 686 557 687
rect 679 691 685 692
rect 679 687 680 691
rect 684 690 685 691
rect 714 691 720 692
rect 714 690 715 691
rect 684 688 715 690
rect 684 687 685 688
rect 679 686 685 687
rect 714 687 715 688
rect 719 687 720 691
rect 714 686 720 687
rect 774 691 780 692
rect 774 687 775 691
rect 779 690 780 691
rect 807 691 813 692
rect 807 690 808 691
rect 779 688 808 690
rect 779 687 780 688
rect 774 686 780 687
rect 807 687 808 688
rect 812 687 813 691
rect 807 686 813 687
rect 834 691 840 692
rect 834 687 835 691
rect 839 690 840 691
rect 927 691 933 692
rect 927 690 928 691
rect 839 688 928 690
rect 839 687 840 688
rect 834 686 840 687
rect 927 687 928 688
rect 932 687 933 691
rect 927 686 933 687
rect 1047 691 1053 692
rect 1047 687 1048 691
rect 1052 690 1053 691
rect 1058 691 1064 692
rect 1058 690 1059 691
rect 1052 688 1059 690
rect 1052 687 1053 688
rect 1047 686 1053 687
rect 1058 687 1059 688
rect 1063 687 1064 691
rect 1058 686 1064 687
rect 1074 691 1080 692
rect 1074 687 1075 691
rect 1079 690 1080 691
rect 1159 691 1165 692
rect 1159 690 1160 691
rect 1079 688 1160 690
rect 1079 687 1080 688
rect 1074 686 1080 687
rect 1159 687 1160 688
rect 1164 687 1165 691
rect 1159 686 1165 687
rect 1186 691 1192 692
rect 1186 687 1187 691
rect 1191 690 1192 691
rect 1271 691 1277 692
rect 1271 690 1272 691
rect 1191 688 1272 690
rect 1191 687 1192 688
rect 1186 686 1192 687
rect 1271 687 1272 688
rect 1276 687 1277 691
rect 1271 686 1277 687
rect 1298 691 1304 692
rect 1298 687 1299 691
rect 1303 690 1304 691
rect 1375 691 1381 692
rect 1375 690 1376 691
rect 1303 688 1376 690
rect 1303 687 1304 688
rect 1298 686 1304 687
rect 1375 687 1376 688
rect 1380 687 1381 691
rect 1375 686 1381 687
rect 1402 691 1408 692
rect 1402 687 1403 691
rect 1407 690 1408 691
rect 1479 691 1485 692
rect 1479 690 1480 691
rect 1407 688 1480 690
rect 1407 687 1408 688
rect 1402 686 1408 687
rect 1479 687 1480 688
rect 1484 687 1485 691
rect 1479 686 1485 687
rect 1506 691 1512 692
rect 1506 687 1507 691
rect 1511 690 1512 691
rect 1583 691 1589 692
rect 1583 690 1584 691
rect 1511 688 1584 690
rect 1511 687 1512 688
rect 1506 686 1512 687
rect 1583 687 1584 688
rect 1588 687 1589 691
rect 1583 686 1589 687
rect 1687 691 1693 692
rect 1687 687 1688 691
rect 1692 690 1693 691
rect 1706 691 1712 692
rect 1706 690 1707 691
rect 1692 688 1707 690
rect 1692 687 1693 688
rect 1687 686 1693 687
rect 1706 687 1707 688
rect 1711 687 1712 691
rect 1706 686 1712 687
rect 1714 691 1720 692
rect 1714 687 1715 691
rect 1719 690 1720 691
rect 1775 691 1781 692
rect 1775 690 1776 691
rect 1719 688 1776 690
rect 1719 687 1720 688
rect 1714 686 1720 687
rect 1775 687 1776 688
rect 1780 687 1781 691
rect 1775 686 1781 687
rect 1927 687 1933 688
rect 1927 683 1928 687
rect 1932 686 1933 687
rect 1970 687 1976 688
rect 1932 684 1966 686
rect 1932 683 1933 684
rect 294 682 300 683
rect 294 678 295 682
rect 299 678 300 682
rect 294 677 300 678
rect 406 682 412 683
rect 406 678 407 682
rect 411 678 412 682
rect 406 677 412 678
rect 526 682 532 683
rect 526 678 527 682
rect 531 678 532 682
rect 526 677 532 678
rect 654 682 660 683
rect 654 678 655 682
rect 659 678 660 682
rect 654 677 660 678
rect 782 682 788 683
rect 782 678 783 682
rect 787 678 788 682
rect 782 677 788 678
rect 902 682 908 683
rect 902 678 903 682
rect 907 678 908 682
rect 902 677 908 678
rect 1022 682 1028 683
rect 1022 678 1023 682
rect 1027 678 1028 682
rect 1022 677 1028 678
rect 1134 682 1140 683
rect 1134 678 1135 682
rect 1139 678 1140 682
rect 1134 677 1140 678
rect 1246 682 1252 683
rect 1246 678 1247 682
rect 1251 678 1252 682
rect 1246 677 1252 678
rect 1350 682 1356 683
rect 1350 678 1351 682
rect 1355 678 1356 682
rect 1350 677 1356 678
rect 1454 682 1460 683
rect 1454 678 1455 682
rect 1459 678 1460 682
rect 1454 677 1460 678
rect 1558 682 1564 683
rect 1558 678 1559 682
rect 1563 678 1564 682
rect 1558 677 1564 678
rect 1662 682 1668 683
rect 1662 678 1663 682
rect 1667 678 1668 682
rect 1662 677 1668 678
rect 1750 682 1756 683
rect 1927 682 1933 683
rect 1750 678 1751 682
rect 1755 678 1756 682
rect 1750 677 1756 678
rect 1964 678 1966 684
rect 1970 683 1971 687
rect 1975 686 1976 687
rect 2007 687 2013 688
rect 2007 686 2008 687
rect 1975 684 2008 686
rect 1975 683 1976 684
rect 1970 682 1976 683
rect 2007 683 2008 684
rect 2012 683 2013 687
rect 2007 682 2013 683
rect 2050 687 2056 688
rect 2050 683 2051 687
rect 2055 686 2056 687
rect 2103 687 2109 688
rect 2103 686 2104 687
rect 2055 684 2104 686
rect 2055 683 2056 684
rect 2050 682 2056 683
rect 2103 683 2104 684
rect 2108 683 2109 687
rect 2103 682 2109 683
rect 2215 687 2221 688
rect 2215 683 2216 687
rect 2220 686 2221 687
rect 2262 687 2268 688
rect 2262 686 2263 687
rect 2220 684 2263 686
rect 2220 683 2221 684
rect 2215 682 2221 683
rect 2262 683 2263 684
rect 2267 683 2268 687
rect 2262 682 2268 683
rect 2298 687 2304 688
rect 2298 683 2299 687
rect 2303 686 2304 687
rect 2343 687 2349 688
rect 2343 686 2344 687
rect 2303 684 2344 686
rect 2303 683 2304 684
rect 2298 682 2304 683
rect 2343 683 2344 684
rect 2348 683 2349 687
rect 2343 682 2349 683
rect 2402 687 2408 688
rect 2402 683 2403 687
rect 2407 686 2408 687
rect 2479 687 2485 688
rect 2479 686 2480 687
rect 2407 684 2480 686
rect 2407 683 2408 684
rect 2402 682 2408 683
rect 2479 683 2480 684
rect 2484 683 2485 687
rect 2479 682 2485 683
rect 2623 687 2629 688
rect 2623 683 2624 687
rect 2628 686 2629 687
rect 2658 687 2664 688
rect 2658 686 2659 687
rect 2628 684 2659 686
rect 2628 683 2629 684
rect 2623 682 2629 683
rect 2658 683 2659 684
rect 2663 683 2664 687
rect 2658 682 2664 683
rect 2775 687 2781 688
rect 2775 683 2776 687
rect 2780 686 2781 687
rect 2810 687 2816 688
rect 2810 686 2811 687
rect 2780 684 2811 686
rect 2780 683 2781 684
rect 2775 682 2781 683
rect 2810 683 2811 684
rect 2815 683 2816 687
rect 2810 682 2816 683
rect 2834 687 2840 688
rect 2834 683 2835 687
rect 2839 686 2840 687
rect 2927 687 2933 688
rect 2927 686 2928 687
rect 2839 684 2928 686
rect 2839 683 2840 684
rect 2834 682 2840 683
rect 2927 683 2928 684
rect 2932 683 2933 687
rect 2927 682 2933 683
rect 3079 687 3085 688
rect 3079 683 3080 687
rect 3084 686 3085 687
rect 3114 687 3120 688
rect 3114 686 3115 687
rect 3084 684 3115 686
rect 3084 683 3085 684
rect 3079 682 3085 683
rect 3114 683 3115 684
rect 3119 683 3120 687
rect 3114 682 3120 683
rect 3231 687 3237 688
rect 3231 683 3232 687
rect 3236 686 3237 687
rect 3266 687 3272 688
rect 3266 686 3267 687
rect 3236 684 3267 686
rect 3236 683 3237 684
rect 3231 682 3237 683
rect 3266 683 3267 684
rect 3271 683 3272 687
rect 3266 682 3272 683
rect 3390 687 3397 688
rect 3390 683 3391 687
rect 3396 683 3397 687
rect 3390 682 3397 683
rect 3534 687 3541 688
rect 3534 683 3535 687
rect 3540 683 3541 687
rect 3534 682 3541 683
rect 2138 679 2144 680
rect 2138 678 2139 679
rect 1964 676 2139 678
rect 2138 675 2139 676
rect 2143 675 2144 679
rect 2138 674 2144 675
rect 1927 671 1933 672
rect 1927 670 1928 671
rect 1804 668 1928 670
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 346 655 352 656
rect 346 651 347 655
rect 351 651 352 655
rect 346 650 352 651
rect 458 655 464 656
rect 458 651 459 655
rect 463 651 464 655
rect 458 650 464 651
rect 578 655 584 656
rect 578 651 579 655
rect 583 651 584 655
rect 774 655 780 656
rect 774 654 775 655
rect 709 652 775 654
rect 578 650 584 651
rect 774 651 775 652
rect 779 651 780 655
rect 774 650 780 651
rect 834 655 840 656
rect 834 651 835 655
rect 839 651 840 655
rect 966 655 972 656
rect 966 654 967 655
rect 957 652 967 654
rect 834 650 840 651
rect 966 651 967 652
rect 971 651 972 655
rect 966 650 972 651
rect 1074 655 1080 656
rect 1074 651 1075 655
rect 1079 651 1080 655
rect 1074 650 1080 651
rect 1186 655 1192 656
rect 1186 651 1187 655
rect 1191 651 1192 655
rect 1186 650 1192 651
rect 1298 655 1304 656
rect 1298 651 1299 655
rect 1303 651 1304 655
rect 1298 650 1304 651
rect 1402 655 1408 656
rect 1402 651 1403 655
rect 1407 651 1408 655
rect 1402 650 1408 651
rect 1506 655 1512 656
rect 1506 651 1507 655
rect 1511 651 1512 655
rect 1506 650 1512 651
rect 1566 655 1572 656
rect 1566 651 1567 655
rect 1571 651 1572 655
rect 1566 650 1572 651
rect 1714 655 1720 656
rect 1714 651 1715 655
rect 1719 651 1720 655
rect 1804 653 1806 668
rect 1927 667 1928 668
rect 1932 667 1933 671
rect 1927 666 1933 667
rect 2119 671 2125 672
rect 2119 667 2120 671
rect 2124 670 2125 671
rect 2130 671 2136 672
rect 2130 670 2131 671
rect 2124 668 2131 670
rect 2124 667 2125 668
rect 2119 666 2125 667
rect 2130 667 2131 668
rect 2135 667 2136 671
rect 2130 666 2136 667
rect 2146 671 2152 672
rect 2146 667 2147 671
rect 2151 670 2152 671
rect 2319 671 2325 672
rect 2319 670 2320 671
rect 2151 668 2320 670
rect 2151 667 2152 668
rect 2146 666 2152 667
rect 2319 667 2320 668
rect 2324 667 2325 671
rect 2319 666 2325 667
rect 2503 671 2509 672
rect 2503 667 2504 671
rect 2508 670 2509 671
rect 2514 671 2520 672
rect 2514 670 2515 671
rect 2508 668 2515 670
rect 2508 667 2509 668
rect 2503 666 2509 667
rect 2514 667 2515 668
rect 2519 667 2520 671
rect 2514 666 2520 667
rect 2530 671 2536 672
rect 2530 667 2531 671
rect 2535 670 2536 671
rect 2679 671 2685 672
rect 2679 670 2680 671
rect 2535 668 2680 670
rect 2535 667 2536 668
rect 2530 666 2536 667
rect 2679 667 2680 668
rect 2684 667 2685 671
rect 2679 666 2685 667
rect 2855 671 2861 672
rect 2855 667 2856 671
rect 2860 670 2861 671
rect 2874 671 2880 672
rect 2874 670 2875 671
rect 2860 668 2875 670
rect 2860 667 2861 668
rect 2855 666 2861 667
rect 2874 667 2875 668
rect 2879 667 2880 671
rect 2874 666 2880 667
rect 2882 671 2888 672
rect 2882 667 2883 671
rect 2887 670 2888 671
rect 3031 671 3037 672
rect 3031 670 3032 671
rect 2887 668 3032 670
rect 2887 667 2888 668
rect 2882 666 2888 667
rect 3031 667 3032 668
rect 3036 667 3037 671
rect 3031 666 3037 667
rect 3174 671 3180 672
rect 3174 667 3175 671
rect 3179 670 3180 671
rect 3207 671 3213 672
rect 3207 670 3208 671
rect 3179 668 3208 670
rect 3179 667 3180 668
rect 3174 666 3180 667
rect 3207 667 3208 668
rect 3212 667 3213 671
rect 3207 666 3213 667
rect 3234 671 3240 672
rect 3234 667 3235 671
rect 3239 670 3240 671
rect 3383 671 3389 672
rect 3383 670 3384 671
rect 3239 668 3384 670
rect 3239 667 3240 668
rect 3234 666 3240 667
rect 3383 667 3384 668
rect 3388 667 3389 671
rect 3383 666 3389 667
rect 3535 671 3541 672
rect 3535 667 3536 671
rect 3540 670 3541 671
rect 3562 671 3568 672
rect 3562 670 3563 671
rect 3540 668 3563 670
rect 3540 667 3541 668
rect 3535 666 3541 667
rect 3562 667 3563 668
rect 3567 667 3568 671
rect 3562 666 3568 667
rect 1830 664 1836 665
rect 1830 660 1831 664
rect 1835 660 1836 664
rect 1830 659 1836 660
rect 1902 662 1908 663
rect 1902 658 1903 662
rect 1907 658 1908 662
rect 1902 657 1908 658
rect 2094 662 2100 663
rect 2094 658 2095 662
rect 2099 658 2100 662
rect 2094 657 2100 658
rect 2294 662 2300 663
rect 2294 658 2295 662
rect 2299 658 2300 662
rect 2294 657 2300 658
rect 2478 662 2484 663
rect 2478 658 2479 662
rect 2483 658 2484 662
rect 2478 657 2484 658
rect 2654 662 2660 663
rect 2654 658 2655 662
rect 2659 658 2660 662
rect 2654 657 2660 658
rect 2830 662 2836 663
rect 2830 658 2831 662
rect 2835 658 2836 662
rect 2830 657 2836 658
rect 3006 662 3012 663
rect 3006 658 3007 662
rect 3011 658 3012 662
rect 3006 657 3012 658
rect 3182 662 3188 663
rect 3182 658 3183 662
rect 3187 658 3188 662
rect 3182 657 3188 658
rect 3358 662 3364 663
rect 3358 658 3359 662
rect 3363 658 3364 662
rect 3358 657 3364 658
rect 3510 662 3516 663
rect 3510 658 3511 662
rect 3515 658 3516 662
rect 3510 657 3516 658
rect 1714 650 1720 651
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 1830 647 1836 648
rect 110 642 116 643
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 518 644 524 645
rect 518 640 519 644
rect 523 640 524 644
rect 518 639 524 640
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 774 644 780 645
rect 774 640 775 644
rect 779 640 780 644
rect 774 639 780 640
rect 894 644 900 645
rect 894 640 895 644
rect 899 640 900 644
rect 894 639 900 640
rect 1014 644 1020 645
rect 1014 640 1015 644
rect 1019 640 1020 644
rect 1014 639 1020 640
rect 1126 644 1132 645
rect 1126 640 1127 644
rect 1131 640 1132 644
rect 1126 639 1132 640
rect 1238 644 1244 645
rect 1238 640 1239 644
rect 1243 640 1244 644
rect 1238 639 1244 640
rect 1342 644 1348 645
rect 1342 640 1343 644
rect 1347 640 1348 644
rect 1342 639 1348 640
rect 1446 644 1452 645
rect 1446 640 1447 644
rect 1451 640 1452 644
rect 1446 639 1452 640
rect 1550 644 1556 645
rect 1550 640 1551 644
rect 1555 640 1556 644
rect 1550 639 1556 640
rect 1654 644 1660 645
rect 1654 640 1655 644
rect 1659 640 1660 644
rect 1654 639 1660 640
rect 1742 644 1748 645
rect 1742 640 1743 644
rect 1747 640 1748 644
rect 1830 643 1831 647
rect 1835 643 1836 647
rect 1830 642 1836 643
rect 1870 644 1876 645
rect 1742 639 1748 640
rect 1870 640 1871 644
rect 1875 640 1876 644
rect 1870 639 1876 640
rect 3590 644 3596 645
rect 3590 640 3591 644
rect 3595 640 3596 644
rect 3590 639 3596 640
rect 1926 635 1932 636
rect 1926 631 1927 635
rect 1931 631 1932 635
rect 1926 630 1932 631
rect 2146 635 2152 636
rect 2146 631 2147 635
rect 2151 631 2152 635
rect 2146 630 2152 631
rect 2302 635 2308 636
rect 2302 631 2303 635
rect 2307 631 2308 635
rect 2302 630 2308 631
rect 2530 635 2536 636
rect 2530 631 2531 635
rect 2535 631 2536 635
rect 2530 630 2536 631
rect 2678 635 2684 636
rect 2678 631 2679 635
rect 2683 631 2684 635
rect 2678 630 2684 631
rect 2882 635 2888 636
rect 2882 631 2883 635
rect 2887 631 2888 635
rect 3174 635 3180 636
rect 3174 634 3175 635
rect 3061 632 3175 634
rect 2882 630 2888 631
rect 3174 631 3175 632
rect 3179 631 3180 635
rect 3174 630 3180 631
rect 3234 635 3240 636
rect 3234 631 3235 635
rect 3239 631 3240 635
rect 3234 630 3240 631
rect 3390 635 3396 636
rect 3390 631 3391 635
rect 3395 631 3396 635
rect 3390 630 3396 631
rect 3534 635 3540 636
rect 3534 631 3535 635
rect 3539 631 3540 635
rect 3534 630 3540 631
rect 1870 627 1876 628
rect 1870 623 1871 627
rect 1875 623 1876 627
rect 3590 627 3596 628
rect 1870 622 1876 623
rect 1894 624 1900 625
rect 1894 620 1895 624
rect 1899 620 1900 624
rect 1894 619 1900 620
rect 2086 624 2092 625
rect 2086 620 2087 624
rect 2091 620 2092 624
rect 2086 619 2092 620
rect 2286 624 2292 625
rect 2286 620 2287 624
rect 2291 620 2292 624
rect 2286 619 2292 620
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2646 624 2652 625
rect 2646 620 2647 624
rect 2651 620 2652 624
rect 2646 619 2652 620
rect 2822 624 2828 625
rect 2822 620 2823 624
rect 2827 620 2828 624
rect 2822 619 2828 620
rect 2998 624 3004 625
rect 2998 620 2999 624
rect 3003 620 3004 624
rect 2998 619 3004 620
rect 3174 624 3180 625
rect 3174 620 3175 624
rect 3179 620 3180 624
rect 3174 619 3180 620
rect 3350 624 3356 625
rect 3350 620 3351 624
rect 3355 620 3356 624
rect 3350 619 3356 620
rect 3502 624 3508 625
rect 3502 620 3503 624
rect 3507 620 3508 624
rect 3590 623 3591 627
rect 3595 623 3596 627
rect 3590 622 3596 623
rect 3502 619 3508 620
rect 310 596 316 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 310 592 311 596
rect 315 592 316 596
rect 310 591 316 592
rect 390 596 396 597
rect 390 592 391 596
rect 395 592 396 596
rect 390 591 396 592
rect 470 596 476 597
rect 470 592 471 596
rect 475 592 476 596
rect 470 591 476 592
rect 558 596 564 597
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 646 596 652 597
rect 646 592 647 596
rect 651 592 652 596
rect 646 591 652 592
rect 734 596 740 597
rect 734 592 735 596
rect 739 592 740 596
rect 734 591 740 592
rect 822 596 828 597
rect 822 592 823 596
rect 827 592 828 596
rect 822 591 828 592
rect 910 596 916 597
rect 910 592 911 596
rect 915 592 916 596
rect 910 591 916 592
rect 998 596 1004 597
rect 998 592 999 596
rect 1003 592 1004 596
rect 998 591 1004 592
rect 1086 596 1092 597
rect 1086 592 1087 596
rect 1091 592 1092 596
rect 1086 591 1092 592
rect 1174 596 1180 597
rect 1174 592 1175 596
rect 1179 592 1180 596
rect 1174 591 1180 592
rect 1262 596 1268 597
rect 1262 592 1263 596
rect 1267 592 1268 596
rect 1262 591 1268 592
rect 1830 593 1836 594
rect 110 588 116 589
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1830 588 1836 589
rect 266 587 272 588
rect 266 583 267 587
rect 271 586 272 587
rect 378 587 384 588
rect 271 584 329 586
rect 271 583 272 584
rect 266 582 272 583
rect 378 583 379 587
rect 383 586 384 587
rect 458 587 464 588
rect 383 584 409 586
rect 383 583 384 584
rect 378 582 384 583
rect 458 583 459 587
rect 463 586 464 587
rect 538 587 544 588
rect 463 584 489 586
rect 463 583 464 584
rect 458 582 464 583
rect 538 583 539 587
rect 543 586 544 587
rect 714 587 720 588
rect 543 584 577 586
rect 543 583 544 584
rect 538 582 544 583
rect 708 580 710 585
rect 714 583 715 587
rect 719 586 720 587
rect 890 587 896 588
rect 890 586 891 587
rect 719 584 753 586
rect 885 584 891 586
rect 719 583 720 584
rect 714 582 720 583
rect 890 583 891 584
rect 895 583 896 587
rect 978 587 984 588
rect 978 586 979 587
rect 973 584 979 586
rect 890 582 896 583
rect 978 583 979 584
rect 983 583 984 587
rect 1066 587 1072 588
rect 1066 586 1067 587
rect 1061 584 1067 586
rect 978 582 984 583
rect 1066 583 1067 584
rect 1071 583 1072 587
rect 1154 587 1160 588
rect 1154 586 1155 587
rect 1149 584 1155 586
rect 1066 582 1072 583
rect 1154 583 1155 584
rect 1159 583 1160 587
rect 1242 587 1248 588
rect 1242 586 1243 587
rect 1237 584 1243 586
rect 1154 582 1160 583
rect 1242 583 1243 584
rect 1247 583 1248 587
rect 1242 582 1248 583
rect 706 579 712 580
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 706 575 707 579
rect 711 575 712 579
rect 706 574 712 575
rect 1058 579 1064 580
rect 1058 575 1059 579
rect 1063 578 1064 579
rect 1280 578 1282 585
rect 1063 576 1282 578
rect 1830 576 1836 577
rect 1063 575 1064 576
rect 1058 574 1064 575
rect 110 571 116 572
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1894 576 1900 577
rect 1830 571 1836 572
rect 1870 573 1876 574
rect 1870 569 1871 573
rect 1875 569 1876 573
rect 1894 572 1895 576
rect 1899 572 1900 576
rect 1894 571 1900 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2086 576 2092 577
rect 2086 572 2087 576
rect 2091 572 2092 576
rect 2086 571 2092 572
rect 2214 576 2220 577
rect 2214 572 2215 576
rect 2219 572 2220 576
rect 2214 571 2220 572
rect 2350 576 2356 577
rect 2350 572 2351 576
rect 2355 572 2356 576
rect 2350 571 2356 572
rect 2494 576 2500 577
rect 2494 572 2495 576
rect 2499 572 2500 576
rect 2494 571 2500 572
rect 2646 576 2652 577
rect 2646 572 2647 576
rect 2651 572 2652 576
rect 2646 571 2652 572
rect 2806 576 2812 577
rect 2806 572 2807 576
rect 2811 572 2812 576
rect 2806 571 2812 572
rect 2974 576 2980 577
rect 2974 572 2975 576
rect 2979 572 2980 576
rect 2974 571 2980 572
rect 3150 576 3156 577
rect 3150 572 3151 576
rect 3155 572 3156 576
rect 3150 571 3156 572
rect 3334 576 3340 577
rect 3334 572 3335 576
rect 3339 572 3340 576
rect 3334 571 3340 572
rect 3502 576 3508 577
rect 3502 572 3503 576
rect 3507 572 3508 576
rect 3502 571 3508 572
rect 3590 573 3596 574
rect 1870 568 1876 569
rect 3590 569 3591 573
rect 3595 569 3596 573
rect 3590 568 3596 569
rect 1962 567 1968 568
rect 1962 566 1963 567
rect 1957 564 1963 566
rect 1962 563 1963 564
rect 1967 563 1968 567
rect 2058 567 2064 568
rect 2058 566 2059 567
rect 2037 564 2059 566
rect 1962 562 1968 563
rect 2058 563 2059 564
rect 2063 563 2064 567
rect 2162 567 2168 568
rect 2162 566 2163 567
rect 2149 564 2163 566
rect 2058 562 2064 563
rect 2162 563 2163 564
rect 2167 563 2168 567
rect 2298 567 2304 568
rect 2298 566 2299 567
rect 2277 564 2299 566
rect 2162 562 2168 563
rect 2298 563 2299 564
rect 2303 563 2304 567
rect 2442 567 2448 568
rect 2442 566 2443 567
rect 2413 564 2443 566
rect 2298 562 2304 563
rect 2442 563 2443 564
rect 2447 563 2448 567
rect 2442 562 2448 563
rect 2450 567 2456 568
rect 2450 563 2451 567
rect 2455 566 2456 567
rect 2746 567 2752 568
rect 2746 566 2747 567
rect 2455 564 2513 566
rect 2709 564 2747 566
rect 2455 563 2456 564
rect 2450 562 2456 563
rect 2746 563 2747 564
rect 2751 563 2752 567
rect 2874 567 2880 568
rect 2746 562 2752 563
rect 2868 560 2870 565
rect 2874 563 2875 567
rect 2879 566 2880 567
rect 3042 567 3048 568
rect 2879 564 2993 566
rect 2879 563 2880 564
rect 2874 562 2880 563
rect 3042 563 3043 567
rect 3047 566 3048 567
rect 3218 567 3224 568
rect 3047 564 3169 566
rect 3047 563 3048 564
rect 3042 562 3048 563
rect 3218 563 3219 567
rect 3223 566 3224 567
rect 3223 564 3353 566
rect 3223 563 3224 564
rect 3218 562 3224 563
rect 3564 560 3566 565
rect 2866 559 2872 560
rect 318 558 324 559
rect 318 554 319 558
rect 323 554 324 558
rect 318 553 324 554
rect 398 558 404 559
rect 398 554 399 558
rect 403 554 404 558
rect 398 553 404 554
rect 478 558 484 559
rect 478 554 479 558
rect 483 554 484 558
rect 478 553 484 554
rect 566 558 572 559
rect 566 554 567 558
rect 571 554 572 558
rect 566 553 572 554
rect 654 558 660 559
rect 654 554 655 558
rect 659 554 660 558
rect 654 553 660 554
rect 742 558 748 559
rect 742 554 743 558
rect 747 554 748 558
rect 742 553 748 554
rect 830 558 836 559
rect 830 554 831 558
rect 835 554 836 558
rect 830 553 836 554
rect 918 558 924 559
rect 918 554 919 558
rect 923 554 924 558
rect 918 553 924 554
rect 1006 558 1012 559
rect 1006 554 1007 558
rect 1011 554 1012 558
rect 1006 553 1012 554
rect 1094 558 1100 559
rect 1094 554 1095 558
rect 1099 554 1100 558
rect 1094 553 1100 554
rect 1182 558 1188 559
rect 1182 554 1183 558
rect 1187 554 1188 558
rect 1182 553 1188 554
rect 1270 558 1276 559
rect 1270 554 1271 558
rect 1275 554 1276 558
rect 1270 553 1276 554
rect 1870 556 1876 557
rect 1870 552 1871 556
rect 1875 552 1876 556
rect 2866 555 2867 559
rect 2871 555 2872 559
rect 2866 554 2872 555
rect 3562 559 3568 560
rect 3562 555 3563 559
rect 3567 555 3568 559
rect 3562 554 3568 555
rect 3590 556 3596 557
rect 1870 551 1876 552
rect 3590 552 3591 556
rect 3595 552 3596 556
rect 3590 551 3596 552
rect 343 547 349 548
rect 343 543 344 547
rect 348 546 349 547
rect 378 547 384 548
rect 378 546 379 547
rect 348 544 379 546
rect 348 543 349 544
rect 343 542 349 543
rect 378 543 379 544
rect 383 543 384 547
rect 378 542 384 543
rect 423 547 429 548
rect 423 543 424 547
rect 428 546 429 547
rect 458 547 464 548
rect 458 546 459 547
rect 428 544 459 546
rect 428 543 429 544
rect 423 542 429 543
rect 458 543 459 544
rect 463 543 464 547
rect 458 542 464 543
rect 503 547 509 548
rect 503 543 504 547
rect 508 546 509 547
rect 538 547 544 548
rect 538 546 539 547
rect 508 544 539 546
rect 508 543 509 544
rect 503 542 509 543
rect 538 543 539 544
rect 543 543 544 547
rect 538 542 544 543
rect 578 547 584 548
rect 578 543 579 547
rect 583 546 584 547
rect 591 547 597 548
rect 591 546 592 547
rect 583 544 592 546
rect 583 543 584 544
rect 578 542 584 543
rect 591 543 592 544
rect 596 543 597 547
rect 591 542 597 543
rect 622 547 628 548
rect 622 543 623 547
rect 627 546 628 547
rect 679 547 685 548
rect 679 546 680 547
rect 627 544 680 546
rect 627 543 628 544
rect 622 542 628 543
rect 679 543 680 544
rect 684 543 685 547
rect 679 542 685 543
rect 706 547 712 548
rect 706 543 707 547
rect 711 546 712 547
rect 767 547 773 548
rect 767 546 768 547
rect 711 544 768 546
rect 711 543 712 544
rect 706 542 712 543
rect 767 543 768 544
rect 772 543 773 547
rect 767 542 773 543
rect 855 547 861 548
rect 855 543 856 547
rect 860 546 861 547
rect 882 547 888 548
rect 882 546 883 547
rect 860 544 883 546
rect 860 543 861 544
rect 855 542 861 543
rect 882 543 883 544
rect 887 543 888 547
rect 882 542 888 543
rect 890 547 896 548
rect 890 543 891 547
rect 895 546 896 547
rect 943 547 949 548
rect 943 546 944 547
rect 895 544 944 546
rect 895 543 896 544
rect 890 542 896 543
rect 943 543 944 544
rect 948 543 949 547
rect 943 542 949 543
rect 978 547 984 548
rect 978 543 979 547
rect 983 546 984 547
rect 1031 547 1037 548
rect 1031 546 1032 547
rect 983 544 1032 546
rect 983 543 984 544
rect 978 542 984 543
rect 1031 543 1032 544
rect 1036 543 1037 547
rect 1031 542 1037 543
rect 1066 547 1072 548
rect 1066 543 1067 547
rect 1071 546 1072 547
rect 1119 547 1125 548
rect 1119 546 1120 547
rect 1071 544 1120 546
rect 1071 543 1072 544
rect 1066 542 1072 543
rect 1119 543 1120 544
rect 1124 543 1125 547
rect 1119 542 1125 543
rect 1154 547 1160 548
rect 1154 543 1155 547
rect 1159 546 1160 547
rect 1207 547 1213 548
rect 1207 546 1208 547
rect 1159 544 1208 546
rect 1159 543 1160 544
rect 1154 542 1160 543
rect 1207 543 1208 544
rect 1212 543 1213 547
rect 1207 542 1213 543
rect 1242 547 1248 548
rect 1242 543 1243 547
rect 1247 546 1248 547
rect 1295 547 1301 548
rect 1295 546 1296 547
rect 1247 544 1296 546
rect 1247 543 1248 544
rect 1242 542 1248 543
rect 1295 543 1296 544
rect 1300 543 1301 547
rect 1295 542 1301 543
rect 1902 538 1908 539
rect 1902 534 1903 538
rect 1907 534 1908 538
rect 1902 533 1908 534
rect 1982 538 1988 539
rect 1982 534 1983 538
rect 1987 534 1988 538
rect 1982 533 1988 534
rect 2094 538 2100 539
rect 2094 534 2095 538
rect 2099 534 2100 538
rect 2094 533 2100 534
rect 2222 538 2228 539
rect 2222 534 2223 538
rect 2227 534 2228 538
rect 2222 533 2228 534
rect 2358 538 2364 539
rect 2358 534 2359 538
rect 2363 534 2364 538
rect 2358 533 2364 534
rect 2502 538 2508 539
rect 2502 534 2503 538
rect 2507 534 2508 538
rect 2502 533 2508 534
rect 2654 538 2660 539
rect 2654 534 2655 538
rect 2659 534 2660 538
rect 2654 533 2660 534
rect 2814 538 2820 539
rect 2814 534 2815 538
rect 2819 534 2820 538
rect 2814 533 2820 534
rect 2982 538 2988 539
rect 2982 534 2983 538
rect 2987 534 2988 538
rect 2982 533 2988 534
rect 3158 538 3164 539
rect 3158 534 3159 538
rect 3163 534 3164 538
rect 3158 533 3164 534
rect 3342 538 3348 539
rect 3342 534 3343 538
rect 3347 534 3348 538
rect 3342 533 3348 534
rect 3510 538 3516 539
rect 3510 534 3511 538
rect 3515 534 3516 538
rect 3510 533 3516 534
rect 786 531 792 532
rect 786 530 787 531
rect 676 528 787 530
rect 263 523 272 524
rect 263 519 264 523
rect 271 519 272 523
rect 263 518 272 519
rect 290 523 296 524
rect 290 519 291 523
rect 295 522 296 523
rect 367 523 373 524
rect 367 522 368 523
rect 295 520 368 522
rect 295 519 296 520
rect 290 518 296 519
rect 367 519 368 520
rect 372 519 373 523
rect 367 518 373 519
rect 463 523 472 524
rect 463 519 464 523
rect 471 519 472 523
rect 463 518 472 519
rect 490 523 496 524
rect 490 519 491 523
rect 495 522 496 523
rect 559 523 565 524
rect 559 522 560 523
rect 495 520 560 522
rect 495 519 496 520
rect 490 518 496 519
rect 559 519 560 520
rect 564 519 565 523
rect 559 518 565 519
rect 655 523 661 524
rect 655 519 656 523
rect 660 522 661 523
rect 676 522 678 528
rect 786 527 787 528
rect 791 527 792 531
rect 786 526 792 527
rect 1926 527 1933 528
rect 660 520 678 522
rect 682 523 688 524
rect 660 519 661 520
rect 655 518 661 519
rect 682 519 683 523
rect 687 522 688 523
rect 743 523 749 524
rect 743 522 744 523
rect 687 520 744 522
rect 687 519 688 520
rect 682 518 688 519
rect 743 519 744 520
rect 748 519 749 523
rect 743 518 749 519
rect 770 523 776 524
rect 770 519 771 523
rect 775 522 776 523
rect 831 523 837 524
rect 831 522 832 523
rect 775 520 832 522
rect 775 519 776 520
rect 770 518 776 519
rect 831 519 832 520
rect 836 519 837 523
rect 831 518 837 519
rect 858 523 864 524
rect 858 519 859 523
rect 863 522 864 523
rect 919 523 925 524
rect 919 522 920 523
rect 863 520 920 522
rect 863 519 864 520
rect 858 518 864 519
rect 919 519 920 520
rect 924 519 925 523
rect 919 518 925 519
rect 946 523 952 524
rect 946 519 947 523
rect 951 522 952 523
rect 1007 523 1013 524
rect 1007 522 1008 523
rect 951 520 1008 522
rect 951 519 952 520
rect 946 518 952 519
rect 1007 519 1008 520
rect 1012 519 1013 523
rect 1007 518 1013 519
rect 1034 523 1040 524
rect 1034 519 1035 523
rect 1039 522 1040 523
rect 1095 523 1101 524
rect 1095 522 1096 523
rect 1039 520 1096 522
rect 1039 519 1040 520
rect 1034 518 1040 519
rect 1095 519 1096 520
rect 1100 519 1101 523
rect 1095 518 1101 519
rect 1122 523 1128 524
rect 1122 519 1123 523
rect 1127 522 1128 523
rect 1183 523 1189 524
rect 1183 522 1184 523
rect 1127 520 1184 522
rect 1127 519 1128 520
rect 1122 518 1128 519
rect 1183 519 1184 520
rect 1188 519 1189 523
rect 1183 518 1189 519
rect 1210 523 1216 524
rect 1210 519 1211 523
rect 1215 522 1216 523
rect 1271 523 1277 524
rect 1271 522 1272 523
rect 1215 520 1272 522
rect 1215 519 1216 520
rect 1210 518 1216 519
rect 1271 519 1272 520
rect 1276 519 1277 523
rect 1926 523 1927 527
rect 1932 523 1933 527
rect 1926 522 1933 523
rect 1962 527 1968 528
rect 1962 523 1963 527
rect 1967 526 1968 527
rect 2007 527 2013 528
rect 2007 526 2008 527
rect 1967 524 2008 526
rect 1967 523 1968 524
rect 1962 522 1968 523
rect 2007 523 2008 524
rect 2012 523 2013 527
rect 2007 522 2013 523
rect 2058 527 2064 528
rect 2058 523 2059 527
rect 2063 526 2064 527
rect 2119 527 2125 528
rect 2119 526 2120 527
rect 2063 524 2120 526
rect 2063 523 2064 524
rect 2058 522 2064 523
rect 2119 523 2120 524
rect 2124 523 2125 527
rect 2119 522 2125 523
rect 2162 527 2168 528
rect 2162 523 2163 527
rect 2167 526 2168 527
rect 2247 527 2253 528
rect 2247 526 2248 527
rect 2167 524 2248 526
rect 2167 523 2168 524
rect 2162 522 2168 523
rect 2247 523 2248 524
rect 2252 523 2253 527
rect 2247 522 2253 523
rect 2298 527 2304 528
rect 2298 523 2299 527
rect 2303 526 2304 527
rect 2383 527 2389 528
rect 2383 526 2384 527
rect 2303 524 2384 526
rect 2303 523 2304 524
rect 2298 522 2304 523
rect 2383 523 2384 524
rect 2388 523 2389 527
rect 2383 522 2389 523
rect 2442 527 2448 528
rect 2442 523 2443 527
rect 2447 526 2448 527
rect 2527 527 2533 528
rect 2527 526 2528 527
rect 2447 524 2528 526
rect 2447 523 2448 524
rect 2442 522 2448 523
rect 2527 523 2528 524
rect 2532 523 2533 527
rect 2527 522 2533 523
rect 2678 527 2685 528
rect 2678 523 2679 527
rect 2684 523 2685 527
rect 2678 522 2685 523
rect 2746 527 2752 528
rect 2746 523 2747 527
rect 2751 526 2752 527
rect 2839 527 2845 528
rect 2839 526 2840 527
rect 2751 524 2840 526
rect 2751 523 2752 524
rect 2746 522 2752 523
rect 2839 523 2840 524
rect 2844 523 2845 527
rect 2839 522 2845 523
rect 3007 527 3013 528
rect 3007 523 3008 527
rect 3012 526 3013 527
rect 3042 527 3048 528
rect 3042 526 3043 527
rect 3012 524 3043 526
rect 3012 523 3013 524
rect 3007 522 3013 523
rect 3042 523 3043 524
rect 3047 523 3048 527
rect 3042 522 3048 523
rect 3183 527 3189 528
rect 3183 523 3184 527
rect 3188 526 3189 527
rect 3218 527 3224 528
rect 3218 526 3219 527
rect 3188 524 3219 526
rect 3188 523 3189 524
rect 3183 522 3189 523
rect 3218 523 3219 524
rect 3223 523 3224 527
rect 3218 522 3224 523
rect 3366 527 3373 528
rect 3366 523 3367 527
rect 3372 523 3373 527
rect 3366 522 3373 523
rect 3534 527 3541 528
rect 3534 523 3535 527
rect 3540 523 3541 527
rect 3534 522 3541 523
rect 1271 518 1277 519
rect 2175 515 2184 516
rect 238 514 244 515
rect 238 510 239 514
rect 243 510 244 514
rect 238 509 244 510
rect 342 514 348 515
rect 342 510 343 514
rect 347 510 348 514
rect 342 509 348 510
rect 438 514 444 515
rect 438 510 439 514
rect 443 510 444 514
rect 438 509 444 510
rect 534 514 540 515
rect 534 510 535 514
rect 539 510 540 514
rect 534 509 540 510
rect 630 514 636 515
rect 630 510 631 514
rect 635 510 636 514
rect 630 509 636 510
rect 718 514 724 515
rect 718 510 719 514
rect 723 510 724 514
rect 718 509 724 510
rect 806 514 812 515
rect 806 510 807 514
rect 811 510 812 514
rect 806 509 812 510
rect 894 514 900 515
rect 894 510 895 514
rect 899 510 900 514
rect 894 509 900 510
rect 982 514 988 515
rect 982 510 983 514
rect 987 510 988 514
rect 982 509 988 510
rect 1070 514 1076 515
rect 1070 510 1071 514
rect 1075 510 1076 514
rect 1070 509 1076 510
rect 1158 514 1164 515
rect 1158 510 1159 514
rect 1163 510 1164 514
rect 1158 509 1164 510
rect 1246 514 1252 515
rect 1246 510 1247 514
rect 1251 510 1252 514
rect 2175 511 2176 515
rect 2183 511 2184 515
rect 2175 510 2184 511
rect 2202 515 2208 516
rect 2202 511 2203 515
rect 2207 514 2208 515
rect 2255 515 2261 516
rect 2255 514 2256 515
rect 2207 512 2256 514
rect 2207 511 2208 512
rect 2202 510 2208 511
rect 2255 511 2256 512
rect 2260 511 2261 515
rect 2255 510 2261 511
rect 2282 515 2288 516
rect 2282 511 2283 515
rect 2287 514 2288 515
rect 2351 515 2357 516
rect 2351 514 2352 515
rect 2287 512 2352 514
rect 2287 511 2288 512
rect 2282 510 2288 511
rect 2351 511 2352 512
rect 2356 511 2357 515
rect 2351 510 2357 511
rect 2378 515 2384 516
rect 2378 511 2379 515
rect 2383 514 2384 515
rect 2455 515 2461 516
rect 2455 514 2456 515
rect 2383 512 2456 514
rect 2383 511 2384 512
rect 2378 510 2384 511
rect 2455 511 2456 512
rect 2460 511 2461 515
rect 2455 510 2461 511
rect 2482 515 2488 516
rect 2482 511 2483 515
rect 2487 514 2488 515
rect 2575 515 2581 516
rect 2575 514 2576 515
rect 2487 512 2576 514
rect 2487 511 2488 512
rect 2482 510 2488 511
rect 2575 511 2576 512
rect 2580 511 2581 515
rect 2575 510 2581 511
rect 2602 515 2608 516
rect 2602 511 2603 515
rect 2607 514 2608 515
rect 2711 515 2717 516
rect 2711 514 2712 515
rect 2607 512 2712 514
rect 2607 511 2608 512
rect 2602 510 2608 511
rect 2711 511 2712 512
rect 2716 511 2717 515
rect 2711 510 2717 511
rect 2863 515 2872 516
rect 2863 511 2864 515
rect 2871 511 2872 515
rect 2863 510 2872 511
rect 2890 515 2896 516
rect 2890 511 2891 515
rect 2895 514 2896 515
rect 3023 515 3029 516
rect 3023 514 3024 515
rect 2895 512 3024 514
rect 2895 511 2896 512
rect 2890 510 2896 511
rect 3023 511 3024 512
rect 3028 511 3029 515
rect 3023 510 3029 511
rect 3199 515 3208 516
rect 3199 511 3200 515
rect 3207 511 3208 515
rect 3199 510 3208 511
rect 3226 515 3232 516
rect 3226 511 3227 515
rect 3231 514 3232 515
rect 3375 515 3381 516
rect 3375 514 3376 515
rect 3231 512 3376 514
rect 3231 511 3232 512
rect 3226 510 3232 511
rect 3375 511 3376 512
rect 3380 511 3381 515
rect 3375 510 3381 511
rect 3535 515 3541 516
rect 3535 511 3536 515
rect 3540 514 3541 515
rect 3562 515 3568 516
rect 3562 514 3563 515
rect 3540 512 3563 514
rect 3540 511 3541 512
rect 3535 510 3541 511
rect 3562 511 3563 512
rect 3567 511 3568 515
rect 3562 510 3568 511
rect 1246 509 1252 510
rect 2150 506 2156 507
rect 2150 502 2151 506
rect 2155 502 2156 506
rect 2150 501 2156 502
rect 2230 506 2236 507
rect 2230 502 2231 506
rect 2235 502 2236 506
rect 2230 501 2236 502
rect 2326 506 2332 507
rect 2326 502 2327 506
rect 2331 502 2332 506
rect 2326 501 2332 502
rect 2430 506 2436 507
rect 2430 502 2431 506
rect 2435 502 2436 506
rect 2430 501 2436 502
rect 2550 506 2556 507
rect 2550 502 2551 506
rect 2555 502 2556 506
rect 2550 501 2556 502
rect 2686 506 2692 507
rect 2686 502 2687 506
rect 2691 502 2692 506
rect 2686 501 2692 502
rect 2838 506 2844 507
rect 2838 502 2839 506
rect 2843 502 2844 506
rect 2838 501 2844 502
rect 2998 506 3004 507
rect 2998 502 2999 506
rect 3003 502 3004 506
rect 2998 501 3004 502
rect 3174 506 3180 507
rect 3174 502 3175 506
rect 3179 502 3180 506
rect 3174 501 3180 502
rect 3350 506 3356 507
rect 3350 502 3351 506
rect 3355 502 3356 506
rect 3350 501 3356 502
rect 3510 506 3516 507
rect 3510 502 3511 506
rect 3515 502 3516 506
rect 3510 501 3516 502
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 1870 488 1876 489
rect 290 487 296 488
rect 290 483 291 487
rect 295 483 296 487
rect 290 482 296 483
rect 394 487 400 488
rect 394 483 395 487
rect 399 483 400 487
rect 394 482 400 483
rect 490 487 496 488
rect 490 483 491 487
rect 495 483 496 487
rect 622 487 628 488
rect 622 486 623 487
rect 589 484 623 486
rect 490 482 496 483
rect 622 483 623 484
rect 627 483 628 487
rect 622 482 628 483
rect 682 487 688 488
rect 682 483 683 487
rect 687 483 688 487
rect 682 482 688 483
rect 770 487 776 488
rect 770 483 771 487
rect 775 483 776 487
rect 770 482 776 483
rect 858 487 864 488
rect 858 483 859 487
rect 863 483 864 487
rect 858 482 864 483
rect 946 487 952 488
rect 946 483 947 487
rect 951 483 952 487
rect 946 482 952 483
rect 1034 487 1040 488
rect 1034 483 1035 487
rect 1039 483 1040 487
rect 1034 482 1040 483
rect 1122 487 1128 488
rect 1122 483 1123 487
rect 1127 483 1128 487
rect 1122 482 1128 483
rect 1210 487 1216 488
rect 1210 483 1211 487
rect 1215 483 1216 487
rect 1210 482 1216 483
rect 1254 487 1260 488
rect 1254 483 1255 487
rect 1259 483 1260 487
rect 1870 484 1871 488
rect 1875 484 1876 488
rect 1870 483 1876 484
rect 3590 488 3596 489
rect 3590 484 3591 488
rect 3595 484 3596 488
rect 3590 483 3596 484
rect 1254 482 1260 483
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 1830 479 1836 480
rect 110 474 116 475
rect 230 476 236 477
rect 230 472 231 476
rect 235 472 236 476
rect 230 471 236 472
rect 334 476 340 477
rect 334 472 335 476
rect 339 472 340 476
rect 334 471 340 472
rect 430 476 436 477
rect 430 472 431 476
rect 435 472 436 476
rect 430 471 436 472
rect 526 476 532 477
rect 526 472 527 476
rect 531 472 532 476
rect 526 471 532 472
rect 622 476 628 477
rect 622 472 623 476
rect 627 472 628 476
rect 622 471 628 472
rect 710 476 716 477
rect 710 472 711 476
rect 715 472 716 476
rect 710 471 716 472
rect 798 476 804 477
rect 798 472 799 476
rect 803 472 804 476
rect 798 471 804 472
rect 886 476 892 477
rect 886 472 887 476
rect 891 472 892 476
rect 886 471 892 472
rect 974 476 980 477
rect 974 472 975 476
rect 979 472 980 476
rect 974 471 980 472
rect 1062 476 1068 477
rect 1062 472 1063 476
rect 1067 472 1068 476
rect 1062 471 1068 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1238 476 1244 477
rect 1238 472 1239 476
rect 1243 472 1244 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 2202 479 2208 480
rect 2202 475 2203 479
rect 2207 475 2208 479
rect 2202 474 2208 475
rect 2282 479 2288 480
rect 2282 475 2283 479
rect 2287 475 2288 479
rect 2282 474 2288 475
rect 2378 479 2384 480
rect 2378 475 2379 479
rect 2383 475 2384 479
rect 2378 474 2384 475
rect 2482 479 2488 480
rect 2482 475 2483 479
rect 2487 475 2488 479
rect 2482 474 2488 475
rect 2602 479 2608 480
rect 2602 475 2603 479
rect 2607 475 2608 479
rect 2602 474 2608 475
rect 2718 479 2724 480
rect 2718 475 2719 479
rect 2723 475 2724 479
rect 2718 474 2724 475
rect 2890 479 2896 480
rect 2890 475 2891 479
rect 2895 475 2896 479
rect 2890 474 2896 475
rect 3050 479 3056 480
rect 3050 475 3051 479
rect 3055 475 3056 479
rect 3050 474 3056 475
rect 3226 479 3232 480
rect 3226 475 3227 479
rect 3231 475 3232 479
rect 3226 474 3232 475
rect 3366 479 3372 480
rect 3366 475 3367 479
rect 3371 475 3372 479
rect 3366 474 3372 475
rect 3534 479 3540 480
rect 3534 475 3535 479
rect 3539 475 3540 479
rect 3534 474 3540 475
rect 1238 471 1244 472
rect 1870 471 1876 472
rect 1870 467 1871 471
rect 1875 467 1876 471
rect 3590 471 3596 472
rect 1870 466 1876 467
rect 2142 468 2148 469
rect 2142 464 2143 468
rect 2147 464 2148 468
rect 2142 463 2148 464
rect 2222 468 2228 469
rect 2222 464 2223 468
rect 2227 464 2228 468
rect 2222 463 2228 464
rect 2318 468 2324 469
rect 2318 464 2319 468
rect 2323 464 2324 468
rect 2318 463 2324 464
rect 2422 468 2428 469
rect 2422 464 2423 468
rect 2427 464 2428 468
rect 2422 463 2428 464
rect 2542 468 2548 469
rect 2542 464 2543 468
rect 2547 464 2548 468
rect 2542 463 2548 464
rect 2678 468 2684 469
rect 2678 464 2679 468
rect 2683 464 2684 468
rect 2678 463 2684 464
rect 2830 468 2836 469
rect 2830 464 2831 468
rect 2835 464 2836 468
rect 2830 463 2836 464
rect 2990 468 2996 469
rect 2990 464 2991 468
rect 2995 464 2996 468
rect 2990 463 2996 464
rect 3166 468 3172 469
rect 3166 464 3167 468
rect 3171 464 3172 468
rect 3166 463 3172 464
rect 3342 468 3348 469
rect 3342 464 3343 468
rect 3347 464 3348 468
rect 3342 463 3348 464
rect 3502 468 3508 469
rect 3502 464 3503 468
rect 3507 464 3508 468
rect 3590 467 3591 471
rect 3595 467 3596 471
rect 3590 466 3596 467
rect 3502 463 3508 464
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 246 424 252 425
rect 246 420 247 424
rect 251 420 252 424
rect 246 419 252 420
rect 374 424 380 425
rect 374 420 375 424
rect 379 420 380 424
rect 374 419 380 420
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 822 424 828 425
rect 822 420 823 424
rect 827 420 828 424
rect 822 419 828 420
rect 918 424 924 425
rect 918 420 919 424
rect 923 420 924 424
rect 918 419 924 420
rect 1006 424 1012 425
rect 1006 420 1007 424
rect 1011 420 1012 424
rect 1006 419 1012 420
rect 1102 424 1108 425
rect 1102 420 1103 424
rect 1107 420 1108 424
rect 1102 419 1108 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 110 416 116 417
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 2334 420 2340 421
rect 1830 416 1836 417
rect 1870 417 1876 418
rect 202 415 208 416
rect 196 408 198 413
rect 202 411 203 415
rect 207 414 208 415
rect 314 415 320 416
rect 207 412 265 414
rect 207 411 208 412
rect 202 410 208 411
rect 314 411 315 415
rect 319 414 320 415
rect 466 415 472 416
rect 319 412 393 414
rect 319 411 320 412
rect 314 410 320 411
rect 466 411 467 415
rect 471 414 472 415
rect 562 415 568 416
rect 471 412 513 414
rect 471 411 472 412
rect 466 410 472 411
rect 562 411 563 415
rect 567 414 568 415
rect 674 415 680 416
rect 567 412 625 414
rect 567 411 568 412
rect 562 410 568 411
rect 674 411 675 415
rect 679 414 680 415
rect 786 415 792 416
rect 679 412 737 414
rect 679 411 680 412
rect 674 410 680 411
rect 786 411 787 415
rect 791 414 792 415
rect 890 415 896 416
rect 791 412 841 414
rect 791 411 792 412
rect 786 410 792 411
rect 890 411 891 415
rect 895 414 896 415
rect 986 415 992 416
rect 895 412 937 414
rect 895 411 896 412
rect 890 410 896 411
rect 986 411 987 415
rect 991 414 992 415
rect 1074 415 1080 416
rect 991 412 1025 414
rect 991 411 992 412
rect 986 410 992 411
rect 1074 411 1075 415
rect 1079 414 1080 415
rect 1270 415 1276 416
rect 1270 414 1271 415
rect 1079 412 1121 414
rect 1261 412 1271 414
rect 1079 411 1080 412
rect 1074 410 1080 411
rect 1270 411 1271 412
rect 1275 411 1276 415
rect 1870 413 1871 417
rect 1875 413 1876 417
rect 2334 416 2335 420
rect 2339 416 2340 420
rect 2334 415 2340 416
rect 2414 420 2420 421
rect 2414 416 2415 420
rect 2419 416 2420 420
rect 2414 415 2420 416
rect 2494 420 2500 421
rect 2494 416 2495 420
rect 2499 416 2500 420
rect 2494 415 2500 416
rect 2582 420 2588 421
rect 2582 416 2583 420
rect 2587 416 2588 420
rect 2582 415 2588 416
rect 2686 420 2692 421
rect 2686 416 2687 420
rect 2691 416 2692 420
rect 2686 415 2692 416
rect 2798 420 2804 421
rect 2798 416 2799 420
rect 2803 416 2804 420
rect 2798 415 2804 416
rect 2926 420 2932 421
rect 2926 416 2927 420
rect 2931 416 2932 420
rect 2926 415 2932 416
rect 3070 420 3076 421
rect 3070 416 3071 420
rect 3075 416 3076 420
rect 3070 415 3076 416
rect 3214 420 3220 421
rect 3214 416 3215 420
rect 3219 416 3220 420
rect 3214 415 3220 416
rect 3366 420 3372 421
rect 3366 416 3367 420
rect 3371 416 3372 420
rect 3366 415 3372 416
rect 3502 420 3508 421
rect 3502 416 3503 420
rect 3507 416 3508 420
rect 3502 415 3508 416
rect 3590 417 3596 418
rect 1270 410 1276 411
rect 194 407 200 408
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 194 403 195 407
rect 199 403 200 407
rect 194 402 200 403
rect 1162 407 1168 408
rect 1162 403 1163 407
rect 1167 406 1168 407
rect 1312 406 1314 413
rect 1870 412 1876 413
rect 3590 413 3591 417
rect 3595 413 3596 417
rect 3590 412 3596 413
rect 2402 411 2408 412
rect 2402 410 2403 411
rect 2397 408 2403 410
rect 2402 407 2403 408
rect 2407 407 2408 411
rect 2482 411 2488 412
rect 2482 410 2483 411
rect 2477 408 2483 410
rect 2402 406 2408 407
rect 2482 407 2483 408
rect 2487 407 2488 411
rect 2562 411 2568 412
rect 2482 406 2488 407
rect 1167 404 1314 406
rect 1830 404 1836 405
rect 1167 403 1168 404
rect 1162 402 1168 403
rect 110 399 116 400
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 2394 403 2400 404
rect 1830 399 1836 400
rect 1870 400 1876 401
rect 1870 396 1871 400
rect 1875 396 1876 400
rect 2394 399 2395 403
rect 2399 402 2400 403
rect 2512 402 2514 409
rect 2562 407 2563 411
rect 2567 410 2568 411
rect 2650 411 2656 412
rect 2567 408 2601 410
rect 2567 407 2568 408
rect 2562 406 2568 407
rect 2650 407 2651 411
rect 2655 410 2656 411
rect 2866 411 2872 412
rect 2655 408 2705 410
rect 2800 408 2817 410
rect 2655 407 2656 408
rect 2650 406 2656 407
rect 2798 407 2804 408
rect 2798 403 2799 407
rect 2803 403 2804 407
rect 2866 407 2867 411
rect 2871 410 2872 411
rect 2994 411 3000 412
rect 2871 408 2945 410
rect 2871 407 2872 408
rect 2866 406 2872 407
rect 2994 407 2995 411
rect 2999 410 3000 411
rect 3202 411 3208 412
rect 2999 408 3089 410
rect 2999 407 3000 408
rect 2994 406 3000 407
rect 3202 407 3203 411
rect 3207 410 3208 411
rect 3282 411 3288 412
rect 3207 408 3233 410
rect 3207 407 3208 408
rect 3202 406 3208 407
rect 3282 407 3283 411
rect 3287 410 3288 411
rect 3434 411 3440 412
rect 3287 408 3385 410
rect 3287 407 3288 408
rect 3282 406 3288 407
rect 3434 407 3435 411
rect 3439 410 3440 411
rect 3439 408 3521 410
rect 3439 407 3440 408
rect 3434 406 3440 407
rect 2798 402 2804 403
rect 2399 400 2514 402
rect 3590 400 3596 401
rect 2399 399 2400 400
rect 2394 398 2400 399
rect 1870 395 1876 396
rect 3590 396 3591 400
rect 3595 396 3596 400
rect 3590 395 3596 396
rect 142 386 148 387
rect 142 382 143 386
rect 147 382 148 386
rect 142 381 148 382
rect 254 386 260 387
rect 254 382 255 386
rect 259 382 260 386
rect 254 381 260 382
rect 382 386 388 387
rect 382 382 383 386
rect 387 382 388 386
rect 382 381 388 382
rect 502 386 508 387
rect 502 382 503 386
rect 507 382 508 386
rect 502 381 508 382
rect 614 386 620 387
rect 614 382 615 386
rect 619 382 620 386
rect 614 381 620 382
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 926 386 932 387
rect 926 382 927 386
rect 931 382 932 386
rect 926 381 932 382
rect 1014 386 1020 387
rect 1014 382 1015 386
rect 1019 382 1020 386
rect 1014 381 1020 382
rect 1110 386 1116 387
rect 1110 382 1111 386
rect 1115 382 1116 386
rect 1110 381 1116 382
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 2342 382 2348 383
rect 2342 378 2343 382
rect 2347 378 2348 382
rect 2342 377 2348 378
rect 2422 382 2428 383
rect 2422 378 2423 382
rect 2427 378 2428 382
rect 2422 377 2428 378
rect 2502 382 2508 383
rect 2502 378 2503 382
rect 2507 378 2508 382
rect 2502 377 2508 378
rect 2590 382 2596 383
rect 2590 378 2591 382
rect 2595 378 2596 382
rect 2590 377 2596 378
rect 2694 382 2700 383
rect 2694 378 2695 382
rect 2699 378 2700 382
rect 2694 377 2700 378
rect 2806 382 2812 383
rect 2806 378 2807 382
rect 2811 378 2812 382
rect 2806 377 2812 378
rect 2934 382 2940 383
rect 2934 378 2935 382
rect 2939 378 2940 382
rect 2934 377 2940 378
rect 3078 382 3084 383
rect 3078 378 3079 382
rect 3083 378 3084 382
rect 3078 377 3084 378
rect 3222 382 3228 383
rect 3222 378 3223 382
rect 3227 378 3228 382
rect 3222 377 3228 378
rect 3374 382 3380 383
rect 3374 378 3375 382
rect 3379 378 3380 382
rect 3374 377 3380 378
rect 3510 382 3516 383
rect 3510 378 3511 382
rect 3515 378 3516 382
rect 3510 377 3516 378
rect 167 375 173 376
rect 167 371 168 375
rect 172 374 173 375
rect 202 375 208 376
rect 202 374 203 375
rect 172 372 203 374
rect 172 371 173 372
rect 167 370 173 371
rect 202 371 203 372
rect 207 371 208 375
rect 202 370 208 371
rect 279 375 285 376
rect 279 371 280 375
rect 284 374 285 375
rect 314 375 320 376
rect 314 374 315 375
rect 284 372 315 374
rect 284 371 285 372
rect 279 370 285 371
rect 314 371 315 372
rect 319 371 320 375
rect 314 370 320 371
rect 394 375 400 376
rect 394 371 395 375
rect 399 374 400 375
rect 407 375 413 376
rect 407 374 408 375
rect 399 372 408 374
rect 399 371 400 372
rect 394 370 400 371
rect 407 371 408 372
rect 412 371 413 375
rect 407 370 413 371
rect 527 375 533 376
rect 527 371 528 375
rect 532 374 533 375
rect 562 375 568 376
rect 562 374 563 375
rect 532 372 563 374
rect 532 371 533 372
rect 527 370 533 371
rect 562 371 563 372
rect 567 371 568 375
rect 562 370 568 371
rect 639 375 645 376
rect 639 371 640 375
rect 644 374 645 375
rect 674 375 680 376
rect 674 374 675 375
rect 644 372 675 374
rect 644 371 645 372
rect 639 370 645 371
rect 674 371 675 372
rect 679 371 680 375
rect 674 370 680 371
rect 751 375 757 376
rect 751 371 752 375
rect 756 374 757 375
rect 782 375 788 376
rect 782 374 783 375
rect 756 372 783 374
rect 756 371 757 372
rect 751 370 757 371
rect 782 371 783 372
rect 787 371 788 375
rect 782 370 788 371
rect 855 375 861 376
rect 855 371 856 375
rect 860 374 861 375
rect 890 375 896 376
rect 890 374 891 375
rect 860 372 891 374
rect 860 371 861 372
rect 855 370 861 371
rect 890 371 891 372
rect 895 371 896 375
rect 890 370 896 371
rect 951 375 957 376
rect 951 371 952 375
rect 956 374 957 375
rect 986 375 992 376
rect 986 374 987 375
rect 956 372 987 374
rect 956 371 957 372
rect 951 370 957 371
rect 986 371 987 372
rect 991 371 992 375
rect 986 370 992 371
rect 1039 375 1045 376
rect 1039 371 1040 375
rect 1044 374 1045 375
rect 1074 375 1080 376
rect 1074 374 1075 375
rect 1044 372 1075 374
rect 1044 371 1045 372
rect 1039 370 1045 371
rect 1074 371 1075 372
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1135 375 1141 376
rect 1135 371 1136 375
rect 1140 374 1141 375
rect 1162 375 1168 376
rect 1162 374 1163 375
rect 1140 372 1163 374
rect 1140 371 1141 372
rect 1135 370 1141 371
rect 1162 371 1163 372
rect 1167 371 1168 375
rect 1162 370 1168 371
rect 1170 375 1176 376
rect 1170 371 1171 375
rect 1175 374 1176 375
rect 1231 375 1237 376
rect 1231 374 1232 375
rect 1175 372 1232 374
rect 1175 371 1176 372
rect 1170 370 1176 371
rect 1231 371 1232 372
rect 1236 371 1237 375
rect 1231 370 1237 371
rect 1270 375 1276 376
rect 1270 371 1271 375
rect 1275 374 1276 375
rect 1327 375 1333 376
rect 1327 374 1328 375
rect 1275 372 1328 374
rect 1275 371 1276 372
rect 1270 370 1276 371
rect 1327 371 1328 372
rect 1332 371 1333 375
rect 2482 375 2488 376
rect 1327 370 1333 371
rect 2367 371 2373 372
rect 2367 367 2368 371
rect 2372 370 2373 371
rect 2394 371 2400 372
rect 2394 370 2395 371
rect 2372 368 2395 370
rect 2372 367 2373 368
rect 2367 366 2373 367
rect 2394 367 2395 368
rect 2399 367 2400 371
rect 2394 366 2400 367
rect 2402 371 2408 372
rect 2402 367 2403 371
rect 2407 370 2408 371
rect 2447 371 2453 372
rect 2447 370 2448 371
rect 2407 368 2448 370
rect 2407 367 2408 368
rect 2402 366 2408 367
rect 2447 367 2448 368
rect 2452 367 2453 371
rect 2482 371 2483 375
rect 2487 374 2488 375
rect 2518 375 2524 376
rect 2518 374 2519 375
rect 2487 372 2519 374
rect 2487 371 2488 372
rect 2482 370 2488 371
rect 2518 371 2519 372
rect 2523 371 2524 375
rect 2518 370 2524 371
rect 2527 371 2533 372
rect 2447 366 2453 367
rect 2527 367 2528 371
rect 2532 370 2533 371
rect 2562 371 2568 372
rect 2562 370 2563 371
rect 2532 368 2563 370
rect 2532 367 2533 368
rect 2527 366 2533 367
rect 2562 367 2563 368
rect 2567 367 2568 371
rect 2562 366 2568 367
rect 2615 371 2621 372
rect 2615 367 2616 371
rect 2620 370 2621 371
rect 2650 371 2656 372
rect 2650 370 2651 371
rect 2620 368 2651 370
rect 2620 367 2621 368
rect 2615 366 2621 367
rect 2650 367 2651 368
rect 2655 367 2656 371
rect 2650 366 2656 367
rect 2718 371 2725 372
rect 2718 367 2719 371
rect 2724 367 2725 371
rect 2718 366 2725 367
rect 2831 371 2837 372
rect 2831 367 2832 371
rect 2836 370 2837 371
rect 2866 371 2872 372
rect 2866 370 2867 371
rect 2836 368 2867 370
rect 2836 367 2837 368
rect 2831 366 2837 367
rect 2866 367 2867 368
rect 2871 367 2872 371
rect 2866 366 2872 367
rect 2959 371 2965 372
rect 2959 367 2960 371
rect 2964 370 2965 371
rect 2994 371 3000 372
rect 2994 370 2995 371
rect 2964 368 2995 370
rect 2964 367 2965 368
rect 2959 366 2965 367
rect 2994 367 2995 368
rect 2999 367 3000 371
rect 2994 366 3000 367
rect 3050 371 3056 372
rect 3050 367 3051 371
rect 3055 370 3056 371
rect 3103 371 3109 372
rect 3103 370 3104 371
rect 3055 368 3104 370
rect 3055 367 3056 368
rect 3050 366 3056 367
rect 3103 367 3104 368
rect 3108 367 3109 371
rect 3103 366 3109 367
rect 3247 371 3253 372
rect 3247 367 3248 371
rect 3252 370 3253 371
rect 3282 371 3288 372
rect 3282 370 3283 371
rect 3252 368 3283 370
rect 3252 367 3253 368
rect 3247 366 3253 367
rect 3282 367 3283 368
rect 3287 367 3288 371
rect 3282 366 3288 367
rect 3338 371 3344 372
rect 3338 367 3339 371
rect 3343 370 3344 371
rect 3399 371 3405 372
rect 3399 370 3400 371
rect 3343 368 3400 370
rect 3343 367 3344 368
rect 3338 366 3344 367
rect 3399 367 3400 368
rect 3404 367 3405 371
rect 3399 366 3405 367
rect 3534 371 3541 372
rect 3534 367 3535 371
rect 3540 367 3541 371
rect 3534 366 3541 367
rect 1230 359 1236 360
rect 1230 358 1231 359
rect 1024 356 1231 358
rect 167 351 173 352
rect 167 347 168 351
rect 172 350 173 351
rect 194 351 200 352
rect 194 350 195 351
rect 172 348 195 350
rect 172 347 173 348
rect 167 346 173 347
rect 194 347 195 348
rect 199 347 200 351
rect 194 346 200 347
rect 207 351 213 352
rect 207 347 208 351
rect 212 350 213 351
rect 271 351 277 352
rect 271 350 272 351
rect 212 348 272 350
rect 212 347 213 348
rect 207 346 213 347
rect 271 347 272 348
rect 276 347 277 351
rect 271 346 277 347
rect 298 351 304 352
rect 298 347 299 351
rect 303 350 304 351
rect 399 351 405 352
rect 399 350 400 351
rect 303 348 400 350
rect 303 347 304 348
rect 298 346 304 347
rect 399 347 400 348
rect 404 347 405 351
rect 399 346 405 347
rect 426 351 432 352
rect 426 347 427 351
rect 431 350 432 351
rect 535 351 541 352
rect 535 350 536 351
rect 431 348 536 350
rect 431 347 432 348
rect 426 346 432 347
rect 535 347 536 348
rect 540 347 541 351
rect 535 346 541 347
rect 662 351 668 352
rect 662 347 663 351
rect 667 350 668 351
rect 671 351 677 352
rect 671 350 672 351
rect 667 348 672 350
rect 667 347 668 348
rect 662 346 668 347
rect 671 347 672 348
rect 676 347 677 351
rect 671 346 677 347
rect 698 351 704 352
rect 698 347 699 351
rect 703 350 704 351
rect 799 351 805 352
rect 799 350 800 351
rect 703 348 800 350
rect 703 347 704 348
rect 698 346 704 347
rect 799 347 800 348
rect 804 347 805 351
rect 799 346 805 347
rect 919 351 925 352
rect 919 347 920 351
rect 924 350 925 351
rect 1024 350 1026 356
rect 1230 355 1231 356
rect 1235 355 1236 359
rect 1446 359 1452 360
rect 1446 358 1447 359
rect 1230 354 1236 355
rect 1336 356 1447 358
rect 924 348 1026 350
rect 1030 351 1037 352
rect 924 347 925 348
rect 919 346 925 347
rect 1030 347 1031 351
rect 1036 347 1037 351
rect 1030 346 1037 347
rect 1058 351 1064 352
rect 1058 347 1059 351
rect 1063 350 1064 351
rect 1143 351 1149 352
rect 1143 350 1144 351
rect 1063 348 1144 350
rect 1063 347 1064 348
rect 1058 346 1064 347
rect 1143 347 1144 348
rect 1148 347 1149 351
rect 1143 346 1149 347
rect 1247 351 1253 352
rect 1247 347 1248 351
rect 1252 350 1253 351
rect 1336 350 1338 356
rect 1446 355 1447 356
rect 1451 355 1452 359
rect 2270 359 2276 360
rect 2270 358 2271 359
rect 1446 354 1452 355
rect 2124 356 2271 358
rect 1252 348 1338 350
rect 1342 351 1348 352
rect 1252 347 1253 348
rect 1247 346 1253 347
rect 1342 347 1343 351
rect 1347 350 1348 351
rect 1351 351 1357 352
rect 1351 350 1352 351
rect 1347 348 1352 350
rect 1347 347 1348 348
rect 1342 346 1348 347
rect 1351 347 1352 348
rect 1356 347 1357 351
rect 1351 346 1357 347
rect 1378 351 1384 352
rect 1378 347 1379 351
rect 1383 350 1384 351
rect 1463 351 1469 352
rect 1463 350 1464 351
rect 1383 348 1464 350
rect 1383 347 1384 348
rect 1378 346 1384 347
rect 1463 347 1464 348
rect 1468 347 1469 351
rect 1463 346 1469 347
rect 2103 351 2109 352
rect 2103 347 2104 351
rect 2108 350 2109 351
rect 2124 350 2126 356
rect 2270 355 2271 356
rect 2275 355 2276 359
rect 2646 359 2652 360
rect 2646 358 2647 359
rect 2270 354 2276 355
rect 2520 356 2647 358
rect 2108 348 2126 350
rect 2130 351 2136 352
rect 2108 347 2109 348
rect 2103 346 2109 347
rect 2130 347 2131 351
rect 2135 350 2136 351
rect 2191 351 2197 352
rect 2191 350 2192 351
rect 2135 348 2192 350
rect 2135 347 2136 348
rect 2130 346 2136 347
rect 2191 347 2192 348
rect 2196 347 2197 351
rect 2191 346 2197 347
rect 2287 351 2293 352
rect 2287 347 2288 351
rect 2292 350 2293 351
rect 2382 351 2388 352
rect 2382 350 2383 351
rect 2292 348 2383 350
rect 2292 347 2293 348
rect 2287 346 2293 347
rect 2382 347 2383 348
rect 2387 347 2388 351
rect 2382 346 2388 347
rect 2399 351 2405 352
rect 2399 347 2400 351
rect 2404 350 2405 351
rect 2520 350 2522 356
rect 2646 355 2647 356
rect 2651 355 2652 359
rect 2646 354 2652 355
rect 2404 348 2522 350
rect 2526 351 2533 352
rect 2404 347 2405 348
rect 2399 346 2405 347
rect 2526 347 2527 351
rect 2532 347 2533 351
rect 2526 346 2533 347
rect 2554 351 2560 352
rect 2554 347 2555 351
rect 2559 350 2560 351
rect 2663 351 2669 352
rect 2663 350 2664 351
rect 2559 348 2664 350
rect 2559 347 2560 348
rect 2554 346 2560 347
rect 2663 347 2664 348
rect 2668 347 2669 351
rect 2663 346 2669 347
rect 2798 351 2805 352
rect 2798 347 2799 351
rect 2804 347 2805 351
rect 2798 346 2805 347
rect 2826 351 2832 352
rect 2826 347 2827 351
rect 2831 350 2832 351
rect 2935 351 2941 352
rect 2935 350 2936 351
rect 2831 348 2936 350
rect 2831 347 2832 348
rect 2826 346 2832 347
rect 2935 347 2936 348
rect 2940 347 2941 351
rect 2935 346 2941 347
rect 3063 351 3072 352
rect 3063 347 3064 351
rect 3071 347 3072 351
rect 3063 346 3072 347
rect 3090 351 3096 352
rect 3090 347 3091 351
rect 3095 350 3096 351
rect 3191 351 3197 352
rect 3191 350 3192 351
rect 3095 348 3192 350
rect 3095 347 3096 348
rect 3090 346 3096 347
rect 3191 347 3192 348
rect 3196 347 3197 351
rect 3191 346 3197 347
rect 3278 351 3284 352
rect 3278 347 3279 351
rect 3283 350 3284 351
rect 3311 351 3317 352
rect 3311 350 3312 351
rect 3283 348 3312 350
rect 3283 347 3284 348
rect 3278 346 3284 347
rect 3311 347 3312 348
rect 3316 347 3317 351
rect 3311 346 3317 347
rect 3431 351 3440 352
rect 3431 347 3432 351
rect 3439 347 3440 351
rect 3431 346 3440 347
rect 3458 351 3464 352
rect 3458 347 3459 351
rect 3463 350 3464 351
rect 3535 351 3541 352
rect 3535 350 3536 351
rect 3463 348 3536 350
rect 3463 347 3464 348
rect 3458 346 3464 347
rect 3535 347 3536 348
rect 3540 347 3541 351
rect 3535 346 3541 347
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 246 342 252 343
rect 246 338 247 342
rect 251 338 252 342
rect 246 337 252 338
rect 374 342 380 343
rect 374 338 375 342
rect 379 338 380 342
rect 374 337 380 338
rect 510 342 516 343
rect 510 338 511 342
rect 515 338 516 342
rect 510 337 516 338
rect 646 342 652 343
rect 646 338 647 342
rect 651 338 652 342
rect 646 337 652 338
rect 774 342 780 343
rect 774 338 775 342
rect 779 338 780 342
rect 774 337 780 338
rect 894 342 900 343
rect 894 338 895 342
rect 899 338 900 342
rect 894 337 900 338
rect 1006 342 1012 343
rect 1006 338 1007 342
rect 1011 338 1012 342
rect 1006 337 1012 338
rect 1118 342 1124 343
rect 1118 338 1119 342
rect 1123 338 1124 342
rect 1118 337 1124 338
rect 1222 342 1228 343
rect 1222 338 1223 342
rect 1227 338 1228 342
rect 1222 337 1228 338
rect 1326 342 1332 343
rect 1326 338 1327 342
rect 1331 338 1332 342
rect 1326 337 1332 338
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 2078 342 2084 343
rect 2078 338 2079 342
rect 2083 338 2084 342
rect 2078 337 2084 338
rect 2166 342 2172 343
rect 2166 338 2167 342
rect 2171 338 2172 342
rect 2166 337 2172 338
rect 2262 342 2268 343
rect 2262 338 2263 342
rect 2267 338 2268 342
rect 2262 337 2268 338
rect 2374 342 2380 343
rect 2374 338 2375 342
rect 2379 338 2380 342
rect 2374 337 2380 338
rect 2502 342 2508 343
rect 2502 338 2503 342
rect 2507 338 2508 342
rect 2502 337 2508 338
rect 2638 342 2644 343
rect 2638 338 2639 342
rect 2643 338 2644 342
rect 2638 337 2644 338
rect 2774 342 2780 343
rect 2774 338 2775 342
rect 2779 338 2780 342
rect 2774 337 2780 338
rect 2910 342 2916 343
rect 2910 338 2911 342
rect 2915 338 2916 342
rect 2910 337 2916 338
rect 3038 342 3044 343
rect 3038 338 3039 342
rect 3043 338 3044 342
rect 3038 337 3044 338
rect 3166 342 3172 343
rect 3166 338 3167 342
rect 3171 338 3172 342
rect 3166 337 3172 338
rect 3286 342 3292 343
rect 3286 338 3287 342
rect 3291 338 3292 342
rect 3286 337 3292 338
rect 3406 342 3412 343
rect 3406 338 3407 342
rect 3411 338 3412 342
rect 3406 337 3412 338
rect 3510 342 3516 343
rect 3510 338 3511 342
rect 3515 338 3516 342
rect 3510 337 3516 338
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1870 324 1876 325
rect 1870 320 1871 324
rect 1875 320 1876 324
rect 1870 319 1876 320
rect 3590 324 3596 325
rect 3590 320 3591 324
rect 3595 320 3596 324
rect 3590 319 3596 320
rect 207 315 213 316
rect 207 314 208 315
rect 197 312 208 314
rect 207 311 208 312
rect 212 311 213 315
rect 207 310 213 311
rect 298 315 304 316
rect 298 311 299 315
rect 303 311 304 315
rect 298 310 304 311
rect 426 315 432 316
rect 426 311 427 315
rect 431 311 432 315
rect 426 310 432 311
rect 698 315 704 316
rect 698 311 699 315
rect 703 311 704 315
rect 698 310 704 311
rect 782 315 788 316
rect 782 311 783 315
rect 787 311 788 315
rect 1006 315 1012 316
rect 1006 314 1007 315
rect 949 312 1007 314
rect 782 310 788 311
rect 1006 311 1007 312
rect 1011 311 1012 315
rect 1006 310 1012 311
rect 1058 315 1064 316
rect 1058 311 1059 315
rect 1063 311 1064 315
rect 1058 310 1064 311
rect 1170 315 1176 316
rect 1170 311 1171 315
rect 1175 311 1176 315
rect 1170 310 1176 311
rect 1230 315 1236 316
rect 1230 311 1231 315
rect 1235 311 1236 315
rect 1230 310 1236 311
rect 1378 315 1384 316
rect 1378 311 1379 315
rect 1383 311 1384 315
rect 1378 310 1384 311
rect 1446 315 1452 316
rect 1446 311 1447 315
rect 1451 311 1452 315
rect 1446 310 1452 311
rect 2130 315 2136 316
rect 2130 311 2131 315
rect 2135 311 2136 315
rect 2238 315 2244 316
rect 2238 314 2239 315
rect 2221 312 2239 314
rect 2130 310 2136 311
rect 2238 311 2239 312
rect 2243 311 2244 315
rect 2238 310 2244 311
rect 2270 315 2276 316
rect 2270 311 2271 315
rect 2275 311 2276 315
rect 2270 310 2276 311
rect 2382 315 2388 316
rect 2382 311 2383 315
rect 2387 311 2388 315
rect 2382 310 2388 311
rect 2554 315 2560 316
rect 2554 311 2555 315
rect 2559 311 2560 315
rect 2554 310 2560 311
rect 2646 315 2652 316
rect 2646 311 2647 315
rect 2651 311 2652 315
rect 2646 310 2652 311
rect 2826 315 2832 316
rect 2826 311 2827 315
rect 2831 311 2832 315
rect 2826 310 2832 311
rect 2962 315 2968 316
rect 2962 311 2963 315
rect 2967 311 2968 315
rect 2962 310 2968 311
rect 3090 315 3096 316
rect 3090 311 3091 315
rect 3095 311 3096 315
rect 3278 315 3284 316
rect 3278 314 3279 315
rect 3221 312 3279 314
rect 3090 310 3096 311
rect 3278 311 3279 312
rect 3283 311 3284 315
rect 3278 310 3284 311
rect 3338 315 3344 316
rect 3338 311 3339 315
rect 3343 311 3344 315
rect 3338 310 3344 311
rect 3458 315 3464 316
rect 3458 311 3459 315
rect 3463 311 3464 315
rect 3458 310 3464 311
rect 3534 315 3540 316
rect 3534 311 3535 315
rect 3539 311 3540 315
rect 3534 310 3540 311
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 1830 307 1836 308
rect 110 302 116 303
rect 134 304 140 305
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 238 304 244 305
rect 238 300 239 304
rect 243 300 244 304
rect 238 299 244 300
rect 366 304 372 305
rect 366 300 367 304
rect 371 300 372 304
rect 366 299 372 300
rect 502 304 508 305
rect 502 300 503 304
rect 507 300 508 304
rect 502 299 508 300
rect 638 304 644 305
rect 638 300 639 304
rect 643 300 644 304
rect 638 299 644 300
rect 766 304 772 305
rect 766 300 767 304
rect 771 300 772 304
rect 766 299 772 300
rect 886 304 892 305
rect 886 300 887 304
rect 891 300 892 304
rect 886 299 892 300
rect 998 304 1004 305
rect 998 300 999 304
rect 1003 300 1004 304
rect 998 299 1004 300
rect 1110 304 1116 305
rect 1110 300 1111 304
rect 1115 300 1116 304
rect 1110 299 1116 300
rect 1214 304 1220 305
rect 1214 300 1215 304
rect 1219 300 1220 304
rect 1214 299 1220 300
rect 1318 304 1324 305
rect 1318 300 1319 304
rect 1323 300 1324 304
rect 1318 299 1324 300
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1870 307 1876 308
rect 1870 303 1871 307
rect 1875 303 1876 307
rect 3590 307 3596 308
rect 1870 302 1876 303
rect 2070 304 2076 305
rect 1430 299 1436 300
rect 2070 300 2071 304
rect 2075 300 2076 304
rect 2070 299 2076 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2254 304 2260 305
rect 2254 300 2255 304
rect 2259 300 2260 304
rect 2254 299 2260 300
rect 2366 304 2372 305
rect 2366 300 2367 304
rect 2371 300 2372 304
rect 2366 299 2372 300
rect 2494 304 2500 305
rect 2494 300 2495 304
rect 2499 300 2500 304
rect 2494 299 2500 300
rect 2630 304 2636 305
rect 2630 300 2631 304
rect 2635 300 2636 304
rect 2630 299 2636 300
rect 2766 304 2772 305
rect 2766 300 2767 304
rect 2771 300 2772 304
rect 2766 299 2772 300
rect 2902 304 2908 305
rect 2902 300 2903 304
rect 2907 300 2908 304
rect 2902 299 2908 300
rect 3030 304 3036 305
rect 3030 300 3031 304
rect 3035 300 3036 304
rect 3030 299 3036 300
rect 3158 304 3164 305
rect 3158 300 3159 304
rect 3163 300 3164 304
rect 3158 299 3164 300
rect 3278 304 3284 305
rect 3278 300 3279 304
rect 3283 300 3284 304
rect 3278 299 3284 300
rect 3398 304 3404 305
rect 3398 300 3399 304
rect 3403 300 3404 304
rect 3398 299 3404 300
rect 3502 304 3508 305
rect 3502 300 3503 304
rect 3507 300 3508 304
rect 3590 303 3591 307
rect 3595 303 3596 307
rect 3590 302 3596 303
rect 3502 299 3508 300
rect 510 287 516 288
rect 510 283 511 287
rect 515 286 516 287
rect 519 287 525 288
rect 519 286 520 287
rect 515 284 520 286
rect 515 283 516 284
rect 510 282 516 283
rect 519 283 520 284
rect 524 283 525 287
rect 519 282 525 283
rect 222 252 228 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 222 248 223 252
rect 227 248 228 252
rect 222 247 228 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 598 252 604 253
rect 598 248 599 252
rect 603 248 604 252
rect 598 247 604 248
rect 734 252 740 253
rect 734 248 735 252
rect 739 248 740 252
rect 734 247 740 248
rect 870 252 876 253
rect 870 248 871 252
rect 875 248 876 252
rect 870 247 876 248
rect 1006 252 1012 253
rect 1006 248 1007 252
rect 1011 248 1012 252
rect 1006 247 1012 248
rect 1134 252 1140 253
rect 1134 248 1135 252
rect 1139 248 1140 252
rect 1134 247 1140 248
rect 1254 252 1260 253
rect 1254 248 1255 252
rect 1259 248 1260 252
rect 1254 247 1260 248
rect 1366 252 1372 253
rect 1366 248 1367 252
rect 1371 248 1372 252
rect 1366 247 1372 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1894 252 1900 253
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 110 244 116 245
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1870 249 1876 250
rect 1870 245 1871 249
rect 1875 245 1876 249
rect 1894 248 1895 252
rect 1899 248 1900 252
rect 1894 247 1900 248
rect 1982 252 1988 253
rect 1982 248 1983 252
rect 1987 248 1988 252
rect 1982 247 1988 248
rect 2094 252 2100 253
rect 2094 248 2095 252
rect 2099 248 2100 252
rect 2094 247 2100 248
rect 2222 252 2228 253
rect 2222 248 2223 252
rect 2227 248 2228 252
rect 2222 247 2228 248
rect 2358 252 2364 253
rect 2358 248 2359 252
rect 2363 248 2364 252
rect 2358 247 2364 248
rect 2502 252 2508 253
rect 2502 248 2503 252
rect 2507 248 2508 252
rect 2502 247 2508 248
rect 2646 252 2652 253
rect 2646 248 2647 252
rect 2651 248 2652 252
rect 2646 247 2652 248
rect 2790 252 2796 253
rect 2790 248 2791 252
rect 2795 248 2796 252
rect 2790 247 2796 248
rect 2934 252 2940 253
rect 2934 248 2935 252
rect 2939 248 2940 252
rect 2934 247 2940 248
rect 3078 252 3084 253
rect 3078 248 3079 252
rect 3083 248 3084 252
rect 3078 247 3084 248
rect 3222 252 3228 253
rect 3222 248 3223 252
rect 3227 248 3228 252
rect 3222 247 3228 248
rect 3374 252 3380 253
rect 3374 248 3375 252
rect 3379 248 3380 252
rect 3374 247 3380 248
rect 3502 252 3508 253
rect 3502 248 3503 252
rect 3507 248 3508 252
rect 3502 247 3508 248
rect 3590 249 3596 250
rect 1870 244 1876 245
rect 3590 245 3591 249
rect 3595 245 3596 249
rect 3590 244 3596 245
rect 186 243 192 244
rect 186 239 187 243
rect 191 242 192 243
rect 290 243 296 244
rect 191 240 241 242
rect 191 239 192 240
rect 186 238 192 239
rect 290 239 291 243
rect 295 242 296 243
rect 402 243 408 244
rect 295 240 353 242
rect 295 239 296 240
rect 290 238 296 239
rect 402 239 403 243
rect 407 242 408 243
rect 666 243 672 244
rect 407 240 481 242
rect 407 239 408 240
rect 402 238 408 239
rect 660 236 662 241
rect 666 239 667 243
rect 671 242 672 243
rect 802 243 808 244
rect 671 240 753 242
rect 671 239 672 240
rect 666 238 672 239
rect 802 239 803 243
rect 807 242 808 243
rect 1078 243 1084 244
rect 1078 242 1079 243
rect 807 240 889 242
rect 1069 240 1079 242
rect 807 239 808 240
rect 802 238 808 239
rect 1078 239 1079 240
rect 1083 239 1084 243
rect 1210 243 1216 244
rect 1210 242 1211 243
rect 1197 240 1211 242
rect 1078 238 1084 239
rect 1210 239 1211 240
rect 1215 239 1216 243
rect 1342 243 1348 244
rect 1342 242 1343 243
rect 1317 240 1343 242
rect 1210 238 1216 239
rect 1342 239 1343 240
rect 1347 239 1348 243
rect 1446 243 1452 244
rect 1446 242 1447 243
rect 1429 240 1447 242
rect 1342 238 1348 239
rect 1446 239 1447 240
rect 1451 239 1452 243
rect 1562 243 1568 244
rect 1562 242 1563 243
rect 1541 240 1563 242
rect 1446 238 1452 239
rect 1562 239 1563 240
rect 1567 239 1568 243
rect 1562 238 1568 239
rect 1570 243 1576 244
rect 1570 239 1571 243
rect 1575 242 1576 243
rect 1962 243 1968 244
rect 1962 242 1963 243
rect 1575 240 1617 242
rect 1957 240 1963 242
rect 1575 239 1576 240
rect 1570 238 1576 239
rect 1962 239 1963 240
rect 1967 239 1968 243
rect 2062 243 2068 244
rect 2062 242 2063 243
rect 2045 240 2063 242
rect 1962 238 1968 239
rect 2062 239 2063 240
rect 2067 239 2068 243
rect 2162 243 2168 244
rect 2162 242 2163 243
rect 2157 240 2163 242
rect 2062 238 2068 239
rect 2162 239 2163 240
rect 2167 239 2168 243
rect 2314 243 2320 244
rect 2314 242 2315 243
rect 2285 240 2315 242
rect 2162 238 2168 239
rect 2314 239 2315 240
rect 2319 239 2320 243
rect 2450 243 2456 244
rect 2450 242 2451 243
rect 2421 240 2451 242
rect 2314 238 2320 239
rect 2450 239 2451 240
rect 2455 239 2456 243
rect 2450 238 2456 239
rect 2458 243 2464 244
rect 2458 239 2459 243
rect 2463 242 2464 243
rect 2610 243 2616 244
rect 2463 240 2521 242
rect 2463 239 2464 240
rect 2458 238 2464 239
rect 2610 239 2611 243
rect 2615 242 2616 243
rect 2714 243 2720 244
rect 2615 240 2665 242
rect 2615 239 2616 240
rect 2610 238 2616 239
rect 2714 239 2715 243
rect 2719 242 2720 243
rect 2878 243 2884 244
rect 2719 240 2809 242
rect 2719 239 2720 240
rect 2714 238 2720 239
rect 2878 239 2879 243
rect 2883 242 2884 243
rect 3066 243 3072 244
rect 2883 240 2953 242
rect 2883 239 2884 240
rect 2878 238 2884 239
rect 3066 239 3067 243
rect 3071 242 3072 243
rect 3146 243 3152 244
rect 3071 240 3097 242
rect 3071 239 3072 240
rect 3066 238 3072 239
rect 3146 239 3147 243
rect 3151 242 3152 243
rect 3290 243 3296 244
rect 3151 240 3241 242
rect 3151 239 3152 240
rect 3146 238 3152 239
rect 3290 239 3291 243
rect 3295 242 3296 243
rect 3295 240 3393 242
rect 3295 239 3296 240
rect 3290 238 3296 239
rect 658 235 664 236
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 658 231 659 235
rect 663 231 664 235
rect 658 230 664 231
rect 1830 232 1836 233
rect 110 227 116 228
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 1870 232 1876 233
rect 1870 228 1871 232
rect 1875 228 1876 232
rect 1870 227 1876 228
rect 3590 232 3596 233
rect 3590 228 3591 232
rect 3595 228 3596 232
rect 3590 227 3596 228
rect 230 214 236 215
rect 230 210 231 214
rect 235 210 236 214
rect 230 209 236 210
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 606 214 612 215
rect 606 210 607 214
rect 611 210 612 214
rect 606 209 612 210
rect 742 214 748 215
rect 742 210 743 214
rect 747 210 748 214
rect 742 209 748 210
rect 878 214 884 215
rect 878 210 879 214
rect 883 210 884 214
rect 878 209 884 210
rect 1014 214 1020 215
rect 1014 210 1015 214
rect 1019 210 1020 214
rect 1014 209 1020 210
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1606 214 1612 215
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1902 214 1908 215
rect 1902 210 1903 214
rect 1907 210 1908 214
rect 1902 209 1908 210
rect 1990 214 1996 215
rect 1990 210 1991 214
rect 1995 210 1996 214
rect 1990 209 1996 210
rect 2102 214 2108 215
rect 2102 210 2103 214
rect 2107 210 2108 214
rect 2102 209 2108 210
rect 2230 214 2236 215
rect 2230 210 2231 214
rect 2235 210 2236 214
rect 2230 209 2236 210
rect 2366 214 2372 215
rect 2366 210 2367 214
rect 2371 210 2372 214
rect 2366 209 2372 210
rect 2510 214 2516 215
rect 2510 210 2511 214
rect 2515 210 2516 214
rect 2510 209 2516 210
rect 2654 214 2660 215
rect 2654 210 2655 214
rect 2659 210 2660 214
rect 2654 209 2660 210
rect 2798 214 2804 215
rect 2798 210 2799 214
rect 2803 210 2804 214
rect 2798 209 2804 210
rect 2942 214 2948 215
rect 2942 210 2943 214
rect 2947 210 2948 214
rect 2942 209 2948 210
rect 3086 214 3092 215
rect 3086 210 3087 214
rect 3091 210 3092 214
rect 3086 209 3092 210
rect 3230 214 3236 215
rect 3230 210 3231 214
rect 3235 210 3236 214
rect 3230 209 3236 210
rect 3382 214 3388 215
rect 3382 210 3383 214
rect 3387 210 3388 214
rect 3382 209 3388 210
rect 3510 214 3516 215
rect 3510 210 3511 214
rect 3515 210 3516 214
rect 3510 209 3516 210
rect 255 203 261 204
rect 255 199 256 203
rect 260 202 261 203
rect 290 203 296 204
rect 290 202 291 203
rect 260 200 291 202
rect 260 199 261 200
rect 255 198 261 199
rect 290 199 291 200
rect 295 199 296 203
rect 290 198 296 199
rect 367 203 373 204
rect 367 199 368 203
rect 372 202 373 203
rect 402 203 408 204
rect 402 202 403 203
rect 372 200 403 202
rect 372 199 373 200
rect 367 198 373 199
rect 402 199 403 200
rect 407 199 408 203
rect 402 198 408 199
rect 495 203 501 204
rect 495 199 496 203
rect 500 202 501 203
rect 510 203 516 204
rect 510 202 511 203
rect 500 200 511 202
rect 500 199 501 200
rect 495 198 501 199
rect 510 199 511 200
rect 515 199 516 203
rect 510 198 516 199
rect 631 203 637 204
rect 631 199 632 203
rect 636 202 637 203
rect 666 203 672 204
rect 666 202 667 203
rect 636 200 667 202
rect 636 199 637 200
rect 631 198 637 199
rect 666 199 667 200
rect 671 199 672 203
rect 666 198 672 199
rect 767 203 773 204
rect 767 199 768 203
rect 772 202 773 203
rect 802 203 808 204
rect 802 202 803 203
rect 772 200 803 202
rect 772 199 773 200
rect 767 198 773 199
rect 802 199 803 200
rect 807 199 808 203
rect 802 198 808 199
rect 902 203 909 204
rect 902 199 903 203
rect 908 199 909 203
rect 902 198 909 199
rect 1039 203 1048 204
rect 1039 199 1040 203
rect 1047 199 1048 203
rect 1039 198 1048 199
rect 1078 203 1084 204
rect 1078 199 1079 203
rect 1083 202 1084 203
rect 1167 203 1173 204
rect 1167 202 1168 203
rect 1083 200 1168 202
rect 1083 199 1084 200
rect 1078 198 1084 199
rect 1167 199 1168 200
rect 1172 199 1173 203
rect 1167 198 1173 199
rect 1210 203 1216 204
rect 1210 199 1211 203
rect 1215 202 1216 203
rect 1287 203 1293 204
rect 1287 202 1288 203
rect 1215 200 1288 202
rect 1215 199 1216 200
rect 1210 198 1216 199
rect 1287 199 1288 200
rect 1292 199 1293 203
rect 1399 203 1405 204
rect 1399 202 1400 203
rect 1287 198 1293 199
rect 1296 200 1400 202
rect 1158 195 1164 196
rect 1158 191 1159 195
rect 1163 194 1164 195
rect 1296 194 1298 200
rect 1399 199 1400 200
rect 1404 199 1405 203
rect 1399 198 1405 199
rect 1446 203 1452 204
rect 1446 199 1447 203
rect 1451 202 1452 203
rect 1511 203 1517 204
rect 1511 202 1512 203
rect 1451 200 1512 202
rect 1451 199 1452 200
rect 1446 198 1452 199
rect 1511 199 1512 200
rect 1516 199 1517 203
rect 1511 198 1517 199
rect 1562 203 1568 204
rect 1562 199 1563 203
rect 1567 202 1568 203
rect 1631 203 1637 204
rect 1631 202 1632 203
rect 1567 200 1632 202
rect 1567 199 1568 200
rect 1562 198 1568 199
rect 1631 199 1632 200
rect 1636 199 1637 203
rect 1631 198 1637 199
rect 1927 203 1936 204
rect 1927 199 1928 203
rect 1935 199 1936 203
rect 1927 198 1936 199
rect 1962 203 1968 204
rect 1962 199 1963 203
rect 1967 202 1968 203
rect 2015 203 2021 204
rect 2015 202 2016 203
rect 1967 200 2016 202
rect 1967 199 1968 200
rect 1962 198 1968 199
rect 2015 199 2016 200
rect 2020 199 2021 203
rect 2015 198 2021 199
rect 2062 203 2068 204
rect 2062 199 2063 203
rect 2067 202 2068 203
rect 2127 203 2133 204
rect 2127 202 2128 203
rect 2067 200 2128 202
rect 2067 199 2068 200
rect 2062 198 2068 199
rect 2127 199 2128 200
rect 2132 199 2133 203
rect 2127 198 2133 199
rect 2238 203 2244 204
rect 2238 199 2239 203
rect 2243 202 2244 203
rect 2255 203 2261 204
rect 2255 202 2256 203
rect 2243 200 2256 202
rect 2243 199 2244 200
rect 2238 198 2244 199
rect 2255 199 2256 200
rect 2260 199 2261 203
rect 2255 198 2261 199
rect 2314 203 2320 204
rect 2314 199 2315 203
rect 2319 202 2320 203
rect 2391 203 2397 204
rect 2391 202 2392 203
rect 2319 200 2392 202
rect 2319 199 2320 200
rect 2314 198 2320 199
rect 2391 199 2392 200
rect 2396 199 2397 203
rect 2391 198 2397 199
rect 2450 203 2456 204
rect 2450 199 2451 203
rect 2455 202 2456 203
rect 2535 203 2541 204
rect 2535 202 2536 203
rect 2455 200 2536 202
rect 2455 199 2456 200
rect 2450 198 2456 199
rect 2535 199 2536 200
rect 2540 199 2541 203
rect 2535 198 2541 199
rect 2679 203 2685 204
rect 2679 199 2680 203
rect 2684 202 2685 203
rect 2714 203 2720 204
rect 2714 202 2715 203
rect 2684 200 2715 202
rect 2684 199 2685 200
rect 2679 198 2685 199
rect 2714 199 2715 200
rect 2719 199 2720 203
rect 2714 198 2720 199
rect 2823 203 2829 204
rect 2823 199 2824 203
rect 2828 202 2829 203
rect 2878 203 2884 204
rect 2878 202 2879 203
rect 2828 200 2879 202
rect 2828 199 2829 200
rect 2823 198 2829 199
rect 2878 199 2879 200
rect 2883 199 2884 203
rect 2878 198 2884 199
rect 2962 203 2973 204
rect 2962 199 2963 203
rect 2967 199 2968 203
rect 2972 199 2973 203
rect 2962 198 2973 199
rect 3111 203 3117 204
rect 3111 199 3112 203
rect 3116 202 3117 203
rect 3146 203 3152 204
rect 3146 202 3147 203
rect 3116 200 3147 202
rect 3116 199 3117 200
rect 3111 198 3117 199
rect 3146 199 3147 200
rect 3151 199 3152 203
rect 3146 198 3152 199
rect 3255 203 3261 204
rect 3255 199 3256 203
rect 3260 202 3261 203
rect 3290 203 3296 204
rect 3290 202 3291 203
rect 3260 200 3291 202
rect 3260 199 3261 200
rect 3255 198 3261 199
rect 3290 199 3291 200
rect 3295 199 3296 203
rect 3290 198 3296 199
rect 3406 203 3413 204
rect 3406 199 3407 203
rect 3412 199 3413 203
rect 3406 198 3413 199
rect 3534 203 3541 204
rect 3534 199 3535 203
rect 3540 199 3541 203
rect 3534 198 3541 199
rect 1163 192 1298 194
rect 1163 191 1164 192
rect 1158 190 1164 191
rect 1927 179 1933 180
rect 1927 175 1928 179
rect 1932 178 1933 179
rect 1962 179 1968 180
rect 1962 178 1963 179
rect 1932 176 1963 178
rect 1932 175 1933 176
rect 1927 174 1933 175
rect 1962 175 1963 176
rect 1967 175 1968 179
rect 1962 174 1968 175
rect 2007 179 2013 180
rect 2007 175 2008 179
rect 2012 178 2013 179
rect 2094 179 2100 180
rect 2094 178 2095 179
rect 2012 176 2095 178
rect 2012 175 2013 176
rect 2007 174 2013 175
rect 2094 175 2095 176
rect 2099 175 2100 179
rect 2094 174 2100 175
rect 2111 179 2117 180
rect 2111 175 2112 179
rect 2116 178 2117 179
rect 2162 179 2168 180
rect 2116 176 2158 178
rect 2116 175 2117 176
rect 2111 174 2117 175
rect 2154 175 2160 176
rect 2154 171 2155 175
rect 2159 171 2160 175
rect 2162 175 2163 179
rect 2167 178 2168 179
rect 2231 179 2237 180
rect 2231 178 2232 179
rect 2167 176 2232 178
rect 2167 175 2168 176
rect 2162 174 2168 175
rect 2231 175 2232 176
rect 2236 175 2237 179
rect 2231 174 2237 175
rect 2258 179 2264 180
rect 2258 175 2259 179
rect 2263 178 2264 179
rect 2359 179 2365 180
rect 2359 178 2360 179
rect 2263 176 2360 178
rect 2263 175 2264 176
rect 2258 174 2264 175
rect 2359 175 2360 176
rect 2364 175 2365 179
rect 2359 174 2365 175
rect 2386 179 2392 180
rect 2386 175 2387 179
rect 2391 178 2392 179
rect 2487 179 2493 180
rect 2487 178 2488 179
rect 2391 176 2488 178
rect 2391 175 2392 176
rect 2386 174 2392 175
rect 2487 175 2488 176
rect 2492 175 2493 179
rect 2487 174 2493 175
rect 2607 179 2616 180
rect 2607 175 2608 179
rect 2615 175 2616 179
rect 2607 174 2616 175
rect 2634 179 2640 180
rect 2634 175 2635 179
rect 2639 178 2640 179
rect 2727 179 2733 180
rect 2727 178 2728 179
rect 2639 176 2728 178
rect 2639 175 2640 176
rect 2634 174 2640 175
rect 2727 175 2728 176
rect 2732 175 2733 179
rect 2727 174 2733 175
rect 2754 179 2760 180
rect 2754 175 2755 179
rect 2759 178 2760 179
rect 2839 179 2845 180
rect 2839 178 2840 179
rect 2759 176 2840 178
rect 2759 175 2760 176
rect 2754 174 2760 175
rect 2839 175 2840 176
rect 2844 175 2845 179
rect 2839 174 2845 175
rect 2866 179 2872 180
rect 2866 175 2867 179
rect 2871 178 2872 179
rect 2943 179 2949 180
rect 2943 178 2944 179
rect 2871 176 2944 178
rect 2871 175 2872 176
rect 2866 174 2872 175
rect 2943 175 2944 176
rect 2948 175 2949 179
rect 2943 174 2949 175
rect 2970 179 2976 180
rect 2970 175 2971 179
rect 2975 178 2976 179
rect 3039 179 3045 180
rect 3039 178 3040 179
rect 2975 176 3040 178
rect 2975 175 2976 176
rect 2970 174 2976 175
rect 3039 175 3040 176
rect 3044 175 3045 179
rect 3039 174 3045 175
rect 3066 179 3072 180
rect 3066 175 3067 179
rect 3071 178 3072 179
rect 3135 179 3141 180
rect 3135 178 3136 179
rect 3071 176 3136 178
rect 3071 175 3072 176
rect 3066 174 3072 175
rect 3135 175 3136 176
rect 3140 175 3141 179
rect 3135 174 3141 175
rect 3162 179 3168 180
rect 3162 175 3163 179
rect 3167 178 3168 179
rect 3231 179 3237 180
rect 3231 178 3232 179
rect 3167 176 3232 178
rect 3167 175 3168 176
rect 3162 174 3168 175
rect 3231 175 3232 176
rect 3236 175 3237 179
rect 3231 174 3237 175
rect 3258 179 3264 180
rect 3258 175 3259 179
rect 3263 178 3264 179
rect 3327 179 3333 180
rect 3327 178 3328 179
rect 3263 176 3328 178
rect 3263 175 3264 176
rect 3258 174 3264 175
rect 3327 175 3328 176
rect 3332 175 3333 179
rect 3327 174 3333 175
rect 3354 179 3360 180
rect 3354 175 3355 179
rect 3359 178 3360 179
rect 3423 179 3429 180
rect 3423 178 3424 179
rect 3359 176 3424 178
rect 3359 175 3360 176
rect 3354 174 3360 175
rect 3423 175 3424 176
rect 3428 175 3429 179
rect 3423 174 3429 175
rect 1902 170 1908 171
rect 1174 167 1180 168
rect 1174 166 1175 167
rect 1016 164 1175 166
rect 183 159 192 160
rect 183 155 184 159
rect 191 155 192 159
rect 183 154 192 155
rect 210 159 216 160
rect 210 155 211 159
rect 215 158 216 159
rect 263 159 269 160
rect 263 158 264 159
rect 215 156 264 158
rect 215 155 216 156
rect 210 154 216 155
rect 263 155 264 156
rect 268 155 269 159
rect 263 154 269 155
rect 290 159 296 160
rect 290 155 291 159
rect 295 158 296 159
rect 343 159 349 160
rect 343 158 344 159
rect 295 156 344 158
rect 295 155 296 156
rect 290 154 296 155
rect 343 155 344 156
rect 348 155 349 159
rect 343 154 349 155
rect 370 159 376 160
rect 370 155 371 159
rect 375 158 376 159
rect 423 159 429 160
rect 423 158 424 159
rect 375 156 424 158
rect 375 155 376 156
rect 370 154 376 155
rect 423 155 424 156
rect 428 155 429 159
rect 423 154 429 155
rect 450 159 456 160
rect 450 155 451 159
rect 455 158 456 159
rect 503 159 509 160
rect 503 158 504 159
rect 455 156 504 158
rect 455 155 456 156
rect 450 154 456 155
rect 503 155 504 156
rect 508 155 509 159
rect 503 154 509 155
rect 530 159 536 160
rect 530 155 531 159
rect 535 158 536 159
rect 583 159 589 160
rect 583 158 584 159
rect 535 156 584 158
rect 535 155 536 156
rect 530 154 536 155
rect 583 155 584 156
rect 588 155 589 159
rect 583 154 589 155
rect 638 159 644 160
rect 638 155 639 159
rect 643 158 644 159
rect 671 159 677 160
rect 671 158 672 159
rect 643 156 672 158
rect 643 155 644 156
rect 638 154 644 155
rect 671 155 672 156
rect 676 155 677 159
rect 671 154 677 155
rect 698 159 704 160
rect 698 155 699 159
rect 703 158 704 159
rect 759 159 765 160
rect 759 158 760 159
rect 703 156 760 158
rect 703 155 704 156
rect 698 154 704 155
rect 759 155 760 156
rect 764 155 765 159
rect 759 154 765 155
rect 786 159 792 160
rect 786 155 787 159
rect 791 158 792 159
rect 847 159 853 160
rect 847 158 848 159
rect 791 156 848 158
rect 791 155 792 156
rect 786 154 792 155
rect 847 155 848 156
rect 852 155 853 159
rect 847 154 853 155
rect 935 159 941 160
rect 935 155 936 159
rect 940 158 941 159
rect 1016 158 1018 164
rect 1174 163 1175 164
rect 1179 163 1180 167
rect 1902 166 1903 170
rect 1907 166 1908 170
rect 1902 165 1908 166
rect 1982 170 1988 171
rect 1982 166 1983 170
rect 1987 166 1988 170
rect 1982 165 1988 166
rect 2086 170 2092 171
rect 2154 170 2160 171
rect 2206 170 2212 171
rect 2086 166 2087 170
rect 2091 166 2092 170
rect 2086 165 2092 166
rect 2206 166 2207 170
rect 2211 166 2212 170
rect 2206 165 2212 166
rect 2334 170 2340 171
rect 2334 166 2335 170
rect 2339 166 2340 170
rect 2334 165 2340 166
rect 2462 170 2468 171
rect 2462 166 2463 170
rect 2467 166 2468 170
rect 2462 165 2468 166
rect 2582 170 2588 171
rect 2582 166 2583 170
rect 2587 166 2588 170
rect 2582 165 2588 166
rect 2702 170 2708 171
rect 2702 166 2703 170
rect 2707 166 2708 170
rect 2702 165 2708 166
rect 2814 170 2820 171
rect 2814 166 2815 170
rect 2819 166 2820 170
rect 2814 165 2820 166
rect 2918 170 2924 171
rect 2918 166 2919 170
rect 2923 166 2924 170
rect 2918 165 2924 166
rect 3014 170 3020 171
rect 3014 166 3015 170
rect 3019 166 3020 170
rect 3014 165 3020 166
rect 3110 170 3116 171
rect 3110 166 3111 170
rect 3115 166 3116 170
rect 3110 165 3116 166
rect 3206 170 3212 171
rect 3206 166 3207 170
rect 3211 166 3212 170
rect 3206 165 3212 166
rect 3302 170 3308 171
rect 3302 166 3303 170
rect 3307 166 3308 170
rect 3302 165 3308 166
rect 3398 170 3404 171
rect 3398 166 3399 170
rect 3403 166 3404 170
rect 3398 165 3404 166
rect 1174 162 1180 163
rect 940 156 1018 158
rect 1022 159 1029 160
rect 940 155 941 156
rect 935 154 941 155
rect 1022 155 1023 159
rect 1028 155 1029 159
rect 1022 154 1029 155
rect 1050 159 1056 160
rect 1050 155 1051 159
rect 1055 158 1056 159
rect 1111 159 1117 160
rect 1111 158 1112 159
rect 1055 156 1112 158
rect 1055 155 1056 156
rect 1050 154 1056 155
rect 1111 155 1112 156
rect 1116 155 1117 159
rect 1111 154 1117 155
rect 1191 159 1197 160
rect 1191 155 1192 159
rect 1196 158 1197 159
rect 1254 159 1260 160
rect 1254 158 1255 159
rect 1196 156 1255 158
rect 1196 155 1197 156
rect 1191 154 1197 155
rect 1254 155 1255 156
rect 1259 155 1260 159
rect 1254 154 1260 155
rect 1271 159 1277 160
rect 1271 155 1272 159
rect 1276 158 1277 159
rect 1342 159 1348 160
rect 1342 158 1343 159
rect 1276 156 1343 158
rect 1276 155 1277 156
rect 1271 154 1277 155
rect 1342 155 1343 156
rect 1347 155 1348 159
rect 1342 154 1348 155
rect 1359 159 1365 160
rect 1359 155 1360 159
rect 1364 158 1365 159
rect 1430 159 1436 160
rect 1430 158 1431 159
rect 1364 156 1431 158
rect 1364 155 1365 156
rect 1359 154 1365 155
rect 1430 155 1431 156
rect 1435 155 1436 159
rect 1430 154 1436 155
rect 1447 159 1453 160
rect 1447 155 1448 159
rect 1452 158 1453 159
rect 1518 159 1524 160
rect 1518 158 1519 159
rect 1452 156 1519 158
rect 1452 155 1453 156
rect 1447 154 1453 155
rect 1518 155 1519 156
rect 1523 155 1524 159
rect 1518 154 1524 155
rect 1535 159 1541 160
rect 1535 155 1536 159
rect 1540 158 1541 159
rect 1598 159 1604 160
rect 1598 158 1599 159
rect 1540 156 1599 158
rect 1540 155 1541 156
rect 1535 154 1541 155
rect 1598 155 1599 156
rect 1603 155 1604 159
rect 1598 154 1604 155
rect 1615 159 1621 160
rect 1615 155 1616 159
rect 1620 158 1621 159
rect 1678 159 1684 160
rect 1678 158 1679 159
rect 1620 156 1679 158
rect 1620 155 1621 156
rect 1615 154 1621 155
rect 1678 155 1679 156
rect 1683 155 1684 159
rect 1678 154 1684 155
rect 1695 159 1701 160
rect 1695 155 1696 159
rect 1700 158 1701 159
rect 1758 159 1764 160
rect 1758 158 1759 159
rect 1700 156 1759 158
rect 1700 155 1701 156
rect 1695 154 1701 155
rect 1758 155 1759 156
rect 1763 155 1764 159
rect 1758 154 1764 155
rect 1775 159 1781 160
rect 1775 155 1776 159
rect 1780 158 1781 159
rect 1780 156 1850 158
rect 1780 155 1781 156
rect 1775 154 1781 155
rect 158 150 164 151
rect 158 146 159 150
rect 163 146 164 150
rect 158 145 164 146
rect 238 150 244 151
rect 238 146 239 150
rect 243 146 244 150
rect 238 145 244 146
rect 318 150 324 151
rect 318 146 319 150
rect 323 146 324 150
rect 318 145 324 146
rect 398 150 404 151
rect 398 146 399 150
rect 403 146 404 150
rect 398 145 404 146
rect 478 150 484 151
rect 478 146 479 150
rect 483 146 484 150
rect 478 145 484 146
rect 558 150 564 151
rect 558 146 559 150
rect 563 146 564 150
rect 558 145 564 146
rect 646 150 652 151
rect 646 146 647 150
rect 651 146 652 150
rect 646 145 652 146
rect 734 150 740 151
rect 734 146 735 150
rect 739 146 740 150
rect 734 145 740 146
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 910 150 916 151
rect 910 146 911 150
rect 915 146 916 150
rect 910 145 916 146
rect 998 150 1004 151
rect 998 146 999 150
rect 1003 146 1004 150
rect 998 145 1004 146
rect 1086 150 1092 151
rect 1086 146 1087 150
rect 1091 146 1092 150
rect 1086 145 1092 146
rect 1166 150 1172 151
rect 1166 146 1167 150
rect 1171 146 1172 150
rect 1166 145 1172 146
rect 1246 150 1252 151
rect 1246 146 1247 150
rect 1251 146 1252 150
rect 1246 145 1252 146
rect 1334 150 1340 151
rect 1334 146 1335 150
rect 1339 146 1340 150
rect 1334 145 1340 146
rect 1422 150 1428 151
rect 1422 146 1423 150
rect 1427 146 1428 150
rect 1422 145 1428 146
rect 1510 150 1516 151
rect 1510 146 1511 150
rect 1515 146 1516 150
rect 1510 145 1516 146
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1670 150 1676 151
rect 1670 146 1671 150
rect 1675 146 1676 150
rect 1670 145 1676 146
rect 1750 150 1756 151
rect 1750 146 1751 150
rect 1755 146 1756 150
rect 1750 145 1756 146
rect 1848 142 1850 156
rect 1870 152 1876 153
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 3590 152 3596 153
rect 3590 148 3591 152
rect 3595 148 3596 152
rect 3590 147 3596 148
rect 1962 143 1968 144
rect 1848 140 1913 142
rect 1962 139 1963 143
rect 1967 142 1968 143
rect 2094 143 2100 144
rect 1967 140 1993 142
rect 1967 139 1968 140
rect 1962 138 1968 139
rect 2094 139 2095 143
rect 2099 139 2100 143
rect 2094 138 2100 139
rect 2258 143 2264 144
rect 2258 139 2259 143
rect 2263 139 2264 143
rect 2258 138 2264 139
rect 2386 143 2392 144
rect 2386 139 2387 143
rect 2391 139 2392 143
rect 2386 138 2392 139
rect 2470 143 2476 144
rect 2470 139 2471 143
rect 2475 139 2476 143
rect 2470 138 2476 139
rect 2634 143 2640 144
rect 2634 139 2635 143
rect 2639 139 2640 143
rect 2634 138 2640 139
rect 2754 143 2760 144
rect 2754 139 2755 143
rect 2759 139 2760 143
rect 2754 138 2760 139
rect 2866 143 2872 144
rect 2866 139 2867 143
rect 2871 139 2872 143
rect 2866 138 2872 139
rect 2970 143 2976 144
rect 2970 139 2971 143
rect 2975 139 2976 143
rect 2970 138 2976 139
rect 3066 143 3072 144
rect 3066 139 3067 143
rect 3071 139 3072 143
rect 3066 138 3072 139
rect 3162 143 3168 144
rect 3162 139 3163 143
rect 3167 139 3168 143
rect 3162 138 3168 139
rect 3258 143 3264 144
rect 3258 139 3259 143
rect 3263 139 3264 143
rect 3258 138 3264 139
rect 3354 143 3360 144
rect 3354 139 3355 143
rect 3359 139 3360 143
rect 3354 138 3360 139
rect 3406 143 3412 144
rect 3406 139 3407 143
rect 3411 139 3412 143
rect 3406 138 3412 139
rect 1870 135 1876 136
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1870 131 1871 135
rect 1875 131 1876 135
rect 3590 135 3596 136
rect 1870 130 1876 131
rect 1894 132 1900 133
rect 1830 127 1836 128
rect 1894 128 1895 132
rect 1899 128 1900 132
rect 1894 127 1900 128
rect 1974 132 1980 133
rect 1974 128 1975 132
rect 1979 128 1980 132
rect 1974 127 1980 128
rect 2078 132 2084 133
rect 2078 128 2079 132
rect 2083 128 2084 132
rect 2078 127 2084 128
rect 2198 132 2204 133
rect 2198 128 2199 132
rect 2203 128 2204 132
rect 2198 127 2204 128
rect 2326 132 2332 133
rect 2326 128 2327 132
rect 2331 128 2332 132
rect 2326 127 2332 128
rect 2454 132 2460 133
rect 2454 128 2455 132
rect 2459 128 2460 132
rect 2454 127 2460 128
rect 2574 132 2580 133
rect 2574 128 2575 132
rect 2579 128 2580 132
rect 2574 127 2580 128
rect 2694 132 2700 133
rect 2694 128 2695 132
rect 2699 128 2700 132
rect 2694 127 2700 128
rect 2806 132 2812 133
rect 2806 128 2807 132
rect 2811 128 2812 132
rect 2806 127 2812 128
rect 2910 132 2916 133
rect 2910 128 2911 132
rect 2915 128 2916 132
rect 2910 127 2916 128
rect 3006 132 3012 133
rect 3006 128 3007 132
rect 3011 128 3012 132
rect 3006 127 3012 128
rect 3102 132 3108 133
rect 3102 128 3103 132
rect 3107 128 3108 132
rect 3102 127 3108 128
rect 3198 132 3204 133
rect 3198 128 3199 132
rect 3203 128 3204 132
rect 3198 127 3204 128
rect 3294 132 3300 133
rect 3294 128 3295 132
rect 3299 128 3300 132
rect 3294 127 3300 128
rect 3390 132 3396 133
rect 3390 128 3391 132
rect 3395 128 3396 132
rect 3590 131 3591 135
rect 3595 131 3596 135
rect 3590 130 3596 131
rect 3390 127 3396 128
rect 210 123 216 124
rect 210 119 211 123
rect 215 119 216 123
rect 210 118 216 119
rect 290 123 296 124
rect 290 119 291 123
rect 295 119 296 123
rect 290 118 296 119
rect 370 123 376 124
rect 370 119 371 123
rect 375 119 376 123
rect 370 118 376 119
rect 450 123 456 124
rect 450 119 451 123
rect 455 119 456 123
rect 450 118 456 119
rect 530 123 536 124
rect 530 119 531 123
rect 535 119 536 123
rect 638 123 644 124
rect 638 122 639 123
rect 613 120 639 122
rect 530 118 536 119
rect 638 119 639 120
rect 643 119 644 123
rect 638 118 644 119
rect 698 123 704 124
rect 698 119 699 123
rect 703 119 704 123
rect 698 118 704 119
rect 786 123 792 124
rect 786 119 787 123
rect 791 119 792 123
rect 902 123 908 124
rect 902 122 903 123
rect 877 120 903 122
rect 786 118 792 119
rect 902 119 903 120
rect 907 119 908 123
rect 998 123 1004 124
rect 998 122 999 123
rect 965 120 999 122
rect 902 118 908 119
rect 998 119 999 120
rect 1003 119 1004 123
rect 998 118 1004 119
rect 1050 123 1056 124
rect 1050 119 1051 123
rect 1055 119 1056 123
rect 1158 123 1164 124
rect 1158 122 1159 123
rect 1141 120 1159 122
rect 1050 118 1056 119
rect 1158 119 1159 120
rect 1163 119 1164 123
rect 1158 118 1164 119
rect 1174 123 1180 124
rect 1174 119 1175 123
rect 1179 119 1180 123
rect 1174 118 1180 119
rect 1254 123 1260 124
rect 1254 119 1255 123
rect 1259 119 1260 123
rect 1254 118 1260 119
rect 1342 123 1348 124
rect 1342 119 1343 123
rect 1347 119 1348 123
rect 1342 118 1348 119
rect 1430 123 1436 124
rect 1430 119 1431 123
rect 1435 119 1436 123
rect 1430 118 1436 119
rect 1518 123 1524 124
rect 1518 119 1519 123
rect 1523 119 1524 123
rect 1518 118 1524 119
rect 1598 123 1604 124
rect 1598 119 1599 123
rect 1603 119 1604 123
rect 1598 118 1604 119
rect 1678 123 1684 124
rect 1678 119 1679 123
rect 1683 119 1684 123
rect 1678 118 1684 119
rect 1758 123 1764 124
rect 1758 119 1759 123
rect 1763 119 1764 123
rect 1758 118 1764 119
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 150 112 156 113
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 230 112 236 113
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 390 112 396 113
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 470 112 476 113
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 550 112 556 113
rect 550 108 551 112
rect 555 108 556 112
rect 550 107 556 108
rect 638 112 644 113
rect 638 108 639 112
rect 643 108 644 112
rect 638 107 644 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 902 112 908 113
rect 902 108 903 112
rect 907 108 908 112
rect 902 107 908 108
rect 990 112 996 113
rect 990 108 991 112
rect 995 108 996 112
rect 990 107 996 108
rect 1078 112 1084 113
rect 1078 108 1079 112
rect 1083 108 1084 112
rect 1078 107 1084 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1326 107 1332 108
rect 1414 112 1420 113
rect 1414 108 1415 112
rect 1419 108 1420 112
rect 1414 107 1420 108
rect 1502 112 1508 113
rect 1502 108 1503 112
rect 1507 108 1508 112
rect 1502 107 1508 108
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1662 112 1668 113
rect 1662 108 1663 112
rect 1667 108 1668 112
rect 1662 107 1668 108
rect 1742 112 1748 113
rect 1742 108 1743 112
rect 1747 108 1748 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1830 110 1836 111
rect 1742 107 1748 108
<< m3c >>
rect 1871 3641 1875 3645
rect 2151 3644 2155 3648
rect 2439 3644 2443 3648
rect 2727 3644 2731 3648
rect 3015 3644 3019 3648
rect 3591 3641 3595 3645
rect 195 3631 199 3635
rect 291 3631 295 3635
rect 419 3631 423 3635
rect 555 3631 559 3635
rect 803 3631 804 3635
rect 804 3631 807 3635
rect 827 3631 831 3635
rect 963 3631 967 3635
rect 1107 3631 1111 3635
rect 2243 3635 2247 3639
rect 2511 3635 2515 3639
rect 3087 3635 3091 3639
rect 143 3622 147 3626
rect 239 3622 243 3626
rect 367 3622 371 3626
rect 503 3622 507 3626
rect 639 3622 643 3626
rect 775 3622 779 3626
rect 911 3622 915 3626
rect 1055 3622 1059 3626
rect 1199 3622 1203 3626
rect 1871 3624 1875 3628
rect 3591 3624 3595 3628
rect 111 3604 115 3608
rect 1831 3604 1835 3608
rect 2159 3606 2163 3610
rect 2447 3606 2451 3610
rect 2735 3606 2739 3610
rect 3023 3606 3027 3610
rect 195 3595 199 3599
rect 291 3595 295 3599
rect 419 3595 423 3599
rect 555 3595 559 3599
rect 827 3595 831 3599
rect 963 3595 967 3599
rect 1107 3595 1111 3599
rect 2183 3595 2184 3599
rect 2184 3595 2187 3599
rect 2503 3595 2507 3599
rect 2511 3595 2515 3599
rect 111 3587 115 3591
rect 135 3584 139 3588
rect 231 3584 235 3588
rect 359 3584 363 3588
rect 495 3584 499 3588
rect 631 3584 635 3588
rect 767 3584 771 3588
rect 903 3584 907 3588
rect 1047 3584 1051 3588
rect 1191 3584 1195 3588
rect 1831 3587 1835 3591
rect 1931 3583 1932 3587
rect 1932 3583 1935 3587
rect 1955 3583 1959 3587
rect 2035 3583 2039 3587
rect 2123 3583 2127 3587
rect 2243 3583 2247 3587
rect 2347 3583 2351 3587
rect 2475 3583 2479 3587
rect 2731 3579 2735 3583
rect 2747 3583 2751 3587
rect 3271 3591 3275 3595
rect 3087 3583 3091 3587
rect 3171 3583 3175 3587
rect 1903 3574 1907 3578
rect 1983 3574 1987 3578
rect 2071 3574 2075 3578
rect 2175 3574 2179 3578
rect 2295 3574 2299 3578
rect 2423 3574 2427 3578
rect 2559 3574 2563 3578
rect 2695 3574 2699 3578
rect 2831 3574 2835 3578
rect 2975 3574 2979 3578
rect 3119 3574 3123 3578
rect 3263 3574 3267 3578
rect 451 3567 455 3571
rect 803 3567 807 3571
rect 911 3567 915 3571
rect 1055 3567 1059 3571
rect 1871 3556 1875 3560
rect 3591 3556 3595 3560
rect 1955 3547 1959 3551
rect 2035 3547 2039 3551
rect 2123 3547 2127 3551
rect 2183 3547 2187 3551
rect 2347 3547 2351 3551
rect 2475 3547 2479 3551
rect 2747 3547 2751 3551
rect 2839 3547 2843 3551
rect 3171 3547 3175 3551
rect 3271 3547 3275 3551
rect 111 3537 115 3541
rect 183 3540 187 3544
rect 303 3540 307 3544
rect 415 3540 419 3544
rect 527 3540 531 3544
rect 631 3540 635 3544
rect 735 3540 739 3544
rect 831 3540 835 3544
rect 919 3540 923 3544
rect 1007 3540 1011 3544
rect 1095 3540 1099 3544
rect 1183 3540 1187 3544
rect 1271 3540 1275 3544
rect 1359 3540 1363 3544
rect 1447 3540 1451 3544
rect 1831 3537 1835 3541
rect 1871 3539 1875 3543
rect 1895 3536 1899 3540
rect 259 3531 263 3535
rect 383 3531 387 3535
rect 111 3520 115 3524
rect 243 3523 247 3527
rect 603 3531 607 3535
rect 707 3531 711 3535
rect 807 3531 811 3535
rect 899 3531 903 3535
rect 911 3531 915 3535
rect 1075 3531 1079 3535
rect 1251 3531 1255 3535
rect 1339 3531 1343 3535
rect 1427 3531 1431 3535
rect 1975 3536 1979 3540
rect 2063 3536 2067 3540
rect 2167 3536 2171 3540
rect 2287 3536 2291 3540
rect 2415 3536 2419 3540
rect 2551 3536 2555 3540
rect 2687 3536 2691 3540
rect 2823 3536 2827 3540
rect 2967 3536 2971 3540
rect 3111 3536 3115 3540
rect 3255 3536 3259 3540
rect 3591 3539 3595 3543
rect 1435 3531 1439 3535
rect 1831 3520 1835 3524
rect 2559 3519 2563 3523
rect 2987 3519 2988 3523
rect 2988 3519 2991 3523
rect 191 3502 195 3506
rect 311 3502 315 3506
rect 423 3502 427 3506
rect 535 3502 539 3506
rect 639 3502 643 3506
rect 743 3502 747 3506
rect 839 3502 843 3506
rect 927 3502 931 3506
rect 1015 3502 1019 3506
rect 1103 3502 1107 3506
rect 1191 3502 1195 3506
rect 1279 3502 1283 3506
rect 1367 3502 1371 3506
rect 1455 3502 1459 3506
rect 243 3491 247 3495
rect 259 3491 263 3495
rect 451 3491 452 3495
rect 452 3491 455 3495
rect 603 3491 607 3495
rect 707 3491 711 3495
rect 807 3491 811 3495
rect 899 3491 903 3495
rect 1055 3491 1059 3495
rect 1075 3491 1079 3495
rect 1251 3491 1255 3495
rect 1339 3491 1343 3495
rect 1427 3491 1431 3495
rect 1871 3489 1875 3493
rect 1967 3492 1971 3496
rect 2151 3492 2155 3496
rect 2335 3492 2339 3496
rect 2511 3492 2515 3496
rect 2671 3492 2675 3496
rect 2823 3492 2827 3496
rect 2959 3492 2963 3496
rect 3079 3492 3083 3496
rect 3191 3492 3195 3496
rect 3303 3492 3307 3496
rect 3415 3492 3419 3496
rect 3503 3492 3507 3496
rect 3591 3489 3595 3493
rect 847 3483 851 3487
rect 1931 3483 1935 3487
rect 2035 3483 2039 3487
rect 2403 3483 2407 3487
rect 2739 3483 2743 3487
rect 3043 3483 3047 3487
rect 3159 3483 3163 3487
rect 3271 3483 3275 3487
rect 3383 3483 3387 3487
rect 3483 3483 3487 3487
rect 375 3471 379 3475
rect 383 3471 387 3475
rect 519 3471 523 3475
rect 555 3471 559 3475
rect 675 3471 679 3475
rect 787 3471 791 3475
rect 987 3471 991 3475
rect 995 3471 999 3475
rect 1091 3471 1095 3475
rect 1207 3471 1211 3475
rect 1871 3472 1875 3476
rect 2731 3475 2735 3479
rect 3563 3475 3567 3479
rect 3591 3472 3595 3476
rect 231 3462 235 3466
rect 367 3462 371 3466
rect 503 3462 507 3466
rect 623 3462 627 3466
rect 735 3462 739 3466
rect 839 3462 843 3466
rect 943 3462 947 3466
rect 1039 3462 1043 3466
rect 1135 3462 1139 3466
rect 1231 3462 1235 3466
rect 1327 3462 1331 3466
rect 1975 3454 1979 3458
rect 2159 3454 2163 3458
rect 2343 3454 2347 3458
rect 2519 3454 2523 3458
rect 2679 3454 2683 3458
rect 2831 3454 2835 3458
rect 2967 3454 2971 3458
rect 3087 3454 3091 3458
rect 3199 3454 3203 3458
rect 3311 3454 3315 3458
rect 3423 3454 3427 3458
rect 3511 3454 3515 3458
rect 111 3444 115 3448
rect 1831 3444 1835 3448
rect 2035 3443 2039 3447
rect 2179 3443 2183 3447
rect 2403 3443 2407 3447
rect 2559 3443 2563 3447
rect 2739 3443 2743 3447
rect 2855 3443 2856 3447
rect 2856 3443 2859 3447
rect 2987 3443 2991 3447
rect 3043 3443 3047 3447
rect 3159 3443 3163 3447
rect 3271 3443 3275 3447
rect 3383 3443 3387 3447
rect 3483 3443 3487 3447
rect 375 3435 379 3439
rect 555 3435 559 3439
rect 675 3435 679 3439
rect 787 3435 791 3439
rect 847 3435 851 3439
rect 995 3435 999 3439
rect 1091 3435 1095 3439
rect 1207 3435 1211 3439
rect 111 3427 115 3431
rect 223 3424 227 3428
rect 359 3424 363 3428
rect 495 3424 499 3428
rect 615 3424 619 3428
rect 727 3424 731 3428
rect 831 3424 835 3428
rect 935 3424 939 3428
rect 1031 3424 1035 3428
rect 1127 3424 1131 3428
rect 1223 3424 1227 3428
rect 1319 3424 1323 3428
rect 1831 3427 1835 3431
rect 2059 3431 2063 3435
rect 2263 3435 2267 3439
rect 2283 3431 2284 3435
rect 2284 3431 2287 3435
rect 2443 3431 2447 3435
rect 2587 3431 2591 3435
rect 3007 3431 3011 3435
rect 3175 3431 3179 3435
rect 3351 3431 3355 3435
rect 3359 3431 3363 3435
rect 3563 3431 3567 3435
rect 2007 3422 2011 3426
rect 2127 3422 2131 3426
rect 2255 3422 2259 3426
rect 2391 3422 2395 3426
rect 2535 3422 2539 3426
rect 2679 3422 2683 3426
rect 2831 3422 2835 3426
rect 2999 3422 3003 3426
rect 3167 3422 3171 3426
rect 3343 3422 3347 3426
rect 3511 3422 3515 3426
rect 243 3407 244 3411
rect 244 3407 247 3411
rect 1247 3407 1251 3411
rect 1871 3404 1875 3408
rect 3591 3404 3595 3408
rect 2059 3395 2063 3399
rect 2179 3395 2183 3399
rect 2263 3395 2267 3399
rect 2443 3395 2447 3399
rect 2587 3395 2591 3399
rect 2855 3395 2859 3399
rect 3007 3395 3011 3399
rect 3175 3395 3179 3399
rect 3351 3395 3355 3399
rect 3535 3395 3539 3399
rect 1871 3387 1875 3391
rect 1999 3384 2003 3388
rect 2119 3384 2123 3388
rect 2247 3384 2251 3388
rect 2383 3384 2387 3388
rect 2527 3384 2531 3388
rect 2671 3384 2675 3388
rect 2823 3384 2827 3388
rect 2991 3384 2995 3388
rect 3159 3384 3163 3388
rect 3335 3384 3339 3388
rect 3503 3384 3507 3388
rect 3591 3387 3595 3391
rect 111 3373 115 3377
rect 215 3376 219 3380
rect 367 3376 371 3380
rect 511 3376 515 3380
rect 647 3376 651 3380
rect 775 3376 779 3380
rect 895 3376 899 3380
rect 1015 3376 1019 3380
rect 1127 3376 1131 3380
rect 1239 3376 1243 3380
rect 1351 3376 1355 3380
rect 1831 3373 1835 3377
rect 283 3367 287 3371
rect 375 3363 379 3367
rect 519 3363 523 3367
rect 579 3367 583 3371
rect 715 3367 719 3371
rect 1095 3367 1099 3371
rect 1207 3367 1211 3371
rect 1319 3367 1323 3371
rect 1327 3367 1331 3371
rect 2619 3367 2623 3371
rect 111 3356 115 3360
rect 1831 3356 1835 3360
rect 223 3338 227 3342
rect 375 3338 379 3342
rect 519 3338 523 3342
rect 655 3338 659 3342
rect 783 3338 787 3342
rect 903 3338 907 3342
rect 1023 3338 1027 3342
rect 1135 3338 1139 3342
rect 1247 3338 1251 3342
rect 1359 3338 1363 3342
rect 1871 3337 1875 3341
rect 2015 3340 2019 3344
rect 2151 3340 2155 3344
rect 2295 3340 2299 3344
rect 2439 3340 2443 3344
rect 2583 3340 2587 3344
rect 2727 3340 2731 3344
rect 2871 3340 2875 3344
rect 3023 3340 3027 3344
rect 3183 3340 3187 3344
rect 3351 3340 3355 3344
rect 3503 3340 3507 3344
rect 3591 3337 3595 3341
rect 243 3327 247 3331
rect 283 3327 287 3331
rect 579 3327 583 3331
rect 715 3327 719 3331
rect 823 3327 827 3331
rect 927 3327 928 3331
rect 928 3327 931 3331
rect 1095 3327 1099 3331
rect 1207 3327 1211 3331
rect 1319 3327 1323 3331
rect 2107 3331 2111 3335
rect 2247 3331 2251 3335
rect 2283 3331 2287 3335
rect 2507 3331 2511 3335
rect 2795 3331 2799 3335
rect 2971 3331 2975 3335
rect 3127 3331 3131 3335
rect 3291 3331 3295 3335
rect 1871 3320 1875 3324
rect 2499 3323 2503 3327
rect 3359 3327 3363 3331
rect 3563 3323 3567 3327
rect 3591 3320 3595 3324
rect 299 3311 303 3315
rect 383 3311 387 3315
rect 547 3311 548 3315
rect 548 3311 551 3315
rect 571 3311 575 3315
rect 723 3311 727 3315
rect 979 3311 980 3315
rect 980 3311 983 3315
rect 1003 3311 1007 3315
rect 1167 3311 1171 3315
rect 1267 3311 1271 3315
rect 1395 3311 1399 3315
rect 207 3302 211 3306
rect 367 3302 371 3306
rect 519 3302 523 3306
rect 671 3302 675 3306
rect 815 3302 819 3306
rect 951 3302 955 3306
rect 1087 3302 1091 3306
rect 1215 3302 1219 3306
rect 1343 3302 1347 3306
rect 1471 3302 1475 3306
rect 2023 3302 2027 3306
rect 2159 3302 2163 3306
rect 2303 3302 2307 3306
rect 2447 3302 2451 3306
rect 2591 3302 2595 3306
rect 2735 3302 2739 3306
rect 2879 3302 2883 3306
rect 3031 3302 3035 3306
rect 3191 3302 3195 3306
rect 3359 3302 3363 3306
rect 3511 3302 3515 3306
rect 1979 3291 1983 3295
rect 2107 3291 2111 3295
rect 2247 3291 2251 3295
rect 2507 3291 2511 3295
rect 2619 3291 2620 3295
rect 2620 3291 2623 3295
rect 2787 3291 2791 3295
rect 2795 3291 2799 3295
rect 2971 3291 2975 3295
rect 3127 3291 3131 3295
rect 3291 3291 3295 3295
rect 3535 3291 3536 3295
rect 3536 3291 3539 3295
rect 111 3284 115 3288
rect 1831 3284 1835 3288
rect 259 3275 263 3279
rect 299 3275 303 3279
rect 571 3275 575 3279
rect 723 3275 727 3279
rect 823 3275 827 3279
rect 1003 3275 1007 3279
rect 1167 3275 1171 3279
rect 1267 3275 1271 3279
rect 1395 3275 1399 3279
rect 2071 3279 2075 3283
rect 2199 3279 2203 3283
rect 2211 3279 2215 3283
rect 2455 3279 2459 3283
rect 2499 3279 2503 3283
rect 2615 3279 2616 3283
rect 2616 3279 2619 3283
rect 2643 3279 2647 3283
rect 2795 3279 2799 3283
rect 2971 3279 2975 3283
rect 3163 3279 3167 3283
rect 3563 3279 3567 3283
rect 111 3267 115 3271
rect 199 3264 203 3268
rect 359 3264 363 3268
rect 511 3264 515 3268
rect 663 3264 667 3268
rect 807 3264 811 3268
rect 943 3264 947 3268
rect 1079 3264 1083 3268
rect 1207 3264 1211 3268
rect 1335 3264 1339 3268
rect 1463 3264 1467 3268
rect 1831 3267 1835 3271
rect 1927 3270 1931 3274
rect 2063 3270 2067 3274
rect 2191 3270 2195 3274
rect 2319 3270 2323 3274
rect 2447 3270 2451 3274
rect 2591 3270 2595 3274
rect 2743 3270 2747 3274
rect 2919 3270 2923 3274
rect 3111 3270 3115 3274
rect 3311 3270 3315 3274
rect 3511 3270 3515 3274
rect 1871 3252 1875 3256
rect 1399 3247 1403 3251
rect 3591 3252 3595 3256
rect 1979 3243 1983 3247
rect 2071 3243 2075 3247
rect 2199 3243 2203 3247
rect 2455 3243 2459 3247
rect 2643 3243 2647 3247
rect 2795 3243 2799 3247
rect 2971 3243 2975 3247
rect 3163 3243 3167 3247
rect 3319 3243 3323 3247
rect 3535 3243 3539 3247
rect 1871 3235 1875 3239
rect 1919 3232 1923 3236
rect 2055 3232 2059 3236
rect 2183 3232 2187 3236
rect 2311 3232 2315 3236
rect 2439 3232 2443 3236
rect 2583 3232 2587 3236
rect 2735 3232 2739 3236
rect 2911 3232 2915 3236
rect 3103 3232 3107 3236
rect 3303 3232 3307 3236
rect 3503 3232 3507 3236
rect 3591 3235 3595 3239
rect 111 3217 115 3221
rect 135 3220 139 3224
rect 271 3220 275 3224
rect 415 3220 419 3224
rect 575 3220 579 3224
rect 735 3220 739 3224
rect 895 3220 899 3224
rect 1047 3220 1051 3224
rect 1191 3220 1195 3224
rect 1327 3220 1331 3224
rect 1463 3220 1467 3224
rect 1607 3220 1611 3224
rect 1831 3217 1835 3221
rect 203 3211 207 3215
rect 111 3200 115 3204
rect 195 3203 199 3207
rect 547 3211 551 3215
rect 643 3211 647 3215
rect 803 3211 807 3215
rect 1115 3211 1119 3215
rect 1283 3211 1287 3215
rect 1419 3211 1423 3215
rect 1559 3211 1563 3215
rect 1587 3211 1591 3215
rect 2327 3215 2328 3219
rect 2328 3215 2331 3219
rect 1831 3200 1835 3204
rect 143 3182 147 3186
rect 279 3182 283 3186
rect 423 3182 427 3186
rect 583 3182 587 3186
rect 743 3182 747 3186
rect 903 3182 907 3186
rect 1055 3182 1059 3186
rect 1199 3182 1203 3186
rect 1335 3182 1339 3186
rect 1471 3182 1475 3186
rect 1615 3182 1619 3186
rect 1871 3185 1875 3189
rect 1895 3188 1899 3192
rect 2007 3188 2011 3192
rect 2143 3188 2147 3192
rect 2295 3188 2299 3192
rect 2455 3188 2459 3192
rect 2623 3188 2627 3192
rect 2799 3188 2803 3192
rect 2975 3188 2979 3192
rect 3151 3188 3155 3192
rect 3327 3188 3331 3192
rect 3503 3188 3507 3192
rect 3591 3185 3595 3189
rect 1963 3179 1967 3183
rect 2091 3179 2095 3183
rect 2211 3179 2215 3183
rect 2371 3179 2375 3183
rect 195 3171 199 3175
rect 259 3171 263 3175
rect 643 3171 647 3175
rect 803 3171 807 3175
rect 1079 3171 1080 3175
rect 1080 3171 1083 3175
rect 1115 3171 1119 3175
rect 1283 3171 1287 3175
rect 1419 3171 1423 3175
rect 1559 3171 1563 3175
rect 2463 3175 2467 3179
rect 2615 3179 2619 3183
rect 2691 3179 2695 3183
rect 2915 3179 2919 3183
rect 3263 3179 3267 3183
rect 3399 3179 3403 3183
rect 1871 3168 1875 3172
rect 3211 3171 3215 3175
rect 3591 3168 3595 3172
rect 203 3151 204 3155
rect 204 3151 207 3155
rect 227 3151 231 3155
rect 499 3151 503 3155
rect 515 3151 519 3155
rect 659 3151 663 3155
rect 911 3151 915 3155
rect 923 3151 927 3155
rect 1043 3151 1047 3155
rect 1155 3151 1159 3155
rect 1259 3151 1263 3155
rect 1363 3151 1367 3155
rect 1459 3151 1463 3155
rect 1547 3151 1551 3155
rect 1635 3151 1639 3155
rect 1723 3151 1727 3155
rect 1903 3150 1907 3154
rect 2015 3150 2019 3154
rect 2151 3150 2155 3154
rect 2303 3150 2307 3154
rect 2463 3150 2467 3154
rect 2631 3150 2635 3154
rect 2807 3150 2811 3154
rect 2983 3150 2987 3154
rect 3159 3150 3163 3154
rect 3335 3150 3339 3154
rect 3511 3150 3515 3154
rect 175 3142 179 3146
rect 319 3142 323 3146
rect 463 3142 467 3146
rect 607 3142 611 3146
rect 743 3142 747 3146
rect 871 3142 875 3146
rect 991 3142 995 3146
rect 1103 3142 1107 3146
rect 1207 3142 1211 3146
rect 1311 3142 1315 3146
rect 1407 3142 1411 3146
rect 1495 3142 1499 3146
rect 1583 3142 1587 3146
rect 1671 3142 1675 3146
rect 1751 3142 1755 3146
rect 1927 3139 1928 3143
rect 1928 3139 1931 3143
rect 1963 3139 1967 3143
rect 2091 3139 2095 3143
rect 2327 3139 2328 3143
rect 2328 3139 2331 3143
rect 2371 3139 2375 3143
rect 2691 3139 2695 3143
rect 2915 3139 2919 3143
rect 3007 3139 3008 3143
rect 3008 3139 3011 3143
rect 3211 3139 3215 3143
rect 3263 3139 3267 3143
rect 3535 3139 3536 3143
rect 3536 3139 3539 3143
rect 111 3124 115 3128
rect 1831 3124 1835 3128
rect 227 3115 231 3119
rect 359 3115 363 3119
rect 515 3115 519 3119
rect 659 3115 663 3119
rect 923 3115 927 3119
rect 1043 3115 1047 3119
rect 1155 3115 1159 3119
rect 1259 3115 1263 3119
rect 1363 3115 1367 3119
rect 1459 3115 1463 3119
rect 1547 3115 1551 3119
rect 1635 3115 1639 3119
rect 1723 3115 1727 3119
rect 2115 3127 2119 3131
rect 2123 3127 2127 3131
rect 2471 3127 2475 3131
rect 2683 3127 2687 3131
rect 2699 3127 2703 3131
rect 3043 3127 3044 3131
rect 3044 3127 3047 3131
rect 3067 3127 3071 3131
rect 3399 3127 3403 3131
rect 1903 3118 1907 3122
rect 2071 3118 2075 3122
rect 2263 3118 2267 3122
rect 2455 3118 2459 3122
rect 2647 3118 2651 3122
rect 2831 3118 2835 3122
rect 3015 3118 3019 3122
rect 3199 3118 3203 3122
rect 3391 3118 3395 3122
rect 111 3107 115 3111
rect 167 3104 171 3108
rect 311 3104 315 3108
rect 455 3104 459 3108
rect 599 3104 603 3108
rect 735 3104 739 3108
rect 863 3104 867 3108
rect 983 3104 987 3108
rect 1095 3104 1099 3108
rect 1199 3104 1203 3108
rect 1303 3104 1307 3108
rect 1399 3104 1403 3108
rect 1487 3104 1491 3108
rect 1575 3104 1579 3108
rect 1663 3104 1667 3108
rect 1743 3104 1747 3108
rect 1831 3107 1835 3111
rect 1871 3100 1875 3104
rect 3591 3100 3595 3104
rect 1927 3091 1931 3095
rect 2123 3091 2127 3095
rect 2315 3091 2319 3095
rect 2699 3091 2703 3095
rect 3007 3091 3011 3095
rect 3067 3091 3071 3095
rect 3283 3091 3287 3095
rect 1871 3083 1875 3087
rect 1895 3080 1899 3084
rect 2063 3080 2067 3084
rect 2255 3080 2259 3084
rect 2447 3080 2451 3084
rect 2639 3080 2643 3084
rect 2823 3080 2827 3084
rect 3007 3080 3011 3084
rect 3191 3080 3195 3084
rect 3383 3080 3387 3084
rect 3591 3083 3595 3087
rect 2115 3063 2119 3067
rect 3043 3063 3047 3067
rect 111 3045 115 3049
rect 135 3048 139 3052
rect 223 3048 227 3052
rect 327 3048 331 3052
rect 439 3048 443 3052
rect 551 3048 555 3052
rect 663 3048 667 3052
rect 1831 3045 1835 3049
rect 203 3039 207 3043
rect 291 3039 295 3043
rect 507 3039 511 3043
rect 619 3039 623 3043
rect 111 3028 115 3032
rect 195 3031 199 3035
rect 499 3031 503 3035
rect 1831 3028 1835 3032
rect 1871 3021 1875 3025
rect 2199 3024 2203 3028
rect 2335 3024 2339 3028
rect 2479 3024 2483 3028
rect 2623 3024 2627 3028
rect 2767 3024 2771 3028
rect 2903 3024 2907 3028
rect 3039 3024 3043 3028
rect 3183 3024 3187 3028
rect 3327 3024 3331 3028
rect 3591 3021 3595 3025
rect 143 3010 147 3014
rect 231 3010 235 3014
rect 335 3010 339 3014
rect 447 3010 451 3014
rect 559 3010 563 3014
rect 671 3010 675 3014
rect 2427 3015 2431 3019
rect 1871 3004 1875 3008
rect 2259 3007 2263 3011
rect 2267 3007 2271 3011
rect 2691 3015 2695 3019
rect 2835 3015 2839 3019
rect 3107 3015 3111 3019
rect 3251 3015 3255 3019
rect 2683 3007 2687 3011
rect 3099 3007 3103 3011
rect 203 2999 207 3003
rect 291 2999 295 3003
rect 359 2999 360 3003
rect 360 2999 363 3003
rect 507 2999 511 3003
rect 619 2999 623 3003
rect 3591 3004 3595 3008
rect 807 2999 811 3003
rect 195 2975 199 2979
rect 211 2975 215 2979
rect 531 2975 535 2979
rect 539 2975 543 2979
rect 699 2975 703 2979
rect 1263 2983 1267 2987
rect 2207 2986 2211 2990
rect 2343 2986 2347 2990
rect 2487 2986 2491 2990
rect 2631 2986 2635 2990
rect 2775 2986 2779 2990
rect 2911 2986 2915 2990
rect 3047 2986 3051 2990
rect 3191 2986 3195 2990
rect 3335 2986 3339 2990
rect 1071 2975 1075 2979
rect 1131 2975 1135 2979
rect 1251 2975 1255 2979
rect 1363 2975 1367 2979
rect 1475 2975 1479 2979
rect 1587 2975 1591 2979
rect 2267 2975 2271 2979
rect 2315 2975 2319 2979
rect 2427 2975 2431 2979
rect 2691 2975 2695 2979
rect 2835 2975 2839 2979
rect 3107 2975 3111 2979
rect 3251 2975 3255 2979
rect 3283 2975 3287 2979
rect 159 2966 163 2970
rect 319 2966 323 2970
rect 487 2966 491 2970
rect 647 2966 651 2970
rect 799 2966 803 2970
rect 943 2966 947 2970
rect 1079 2966 1083 2970
rect 1199 2966 1203 2970
rect 1311 2966 1315 2970
rect 1423 2966 1427 2970
rect 1535 2966 1539 2970
rect 1647 2966 1651 2970
rect 111 2948 115 2952
rect 1831 2948 1835 2952
rect 2215 2951 2219 2955
rect 2259 2951 2263 2955
rect 2315 2951 2316 2955
rect 2316 2951 2319 2955
rect 2351 2951 2355 2955
rect 2419 2951 2423 2955
rect 2499 2951 2503 2955
rect 2579 2951 2583 2955
rect 2659 2951 2663 2955
rect 2747 2951 2751 2955
rect 2947 2951 2951 2955
rect 2963 2951 2967 2955
rect 3099 2951 3103 2955
rect 3235 2951 3239 2955
rect 3439 2951 3443 2955
rect 211 2939 215 2943
rect 343 2939 347 2943
rect 539 2939 543 2943
rect 699 2939 703 2943
rect 807 2939 811 2943
rect 1071 2939 1075 2943
rect 1131 2939 1135 2943
rect 1251 2939 1255 2943
rect 1363 2939 1367 2943
rect 1475 2939 1479 2943
rect 1587 2939 1591 2943
rect 2127 2942 2131 2946
rect 2207 2942 2211 2946
rect 2287 2942 2291 2946
rect 2367 2942 2371 2946
rect 2447 2942 2451 2946
rect 2527 2942 2531 2946
rect 2607 2942 2611 2946
rect 2695 2942 2699 2946
rect 2791 2942 2795 2946
rect 2911 2942 2915 2946
rect 3039 2942 3043 2946
rect 3183 2942 3187 2946
rect 3335 2942 3339 2946
rect 3495 2942 3499 2946
rect 111 2931 115 2935
rect 151 2928 155 2932
rect 311 2928 315 2932
rect 479 2928 483 2932
rect 639 2928 643 2932
rect 791 2928 795 2932
rect 935 2928 939 2932
rect 1071 2928 1075 2932
rect 1191 2928 1195 2932
rect 1303 2928 1307 2932
rect 1415 2928 1419 2932
rect 1527 2928 1531 2932
rect 1639 2928 1643 2932
rect 1831 2931 1835 2935
rect 1871 2924 1875 2928
rect 3591 2924 3595 2928
rect 1427 2911 1431 2915
rect 2215 2915 2219 2919
rect 2351 2915 2355 2919
rect 2419 2915 2423 2919
rect 2499 2915 2503 2919
rect 2579 2915 2583 2919
rect 2659 2915 2663 2919
rect 2747 2915 2751 2919
rect 2963 2915 2967 2919
rect 3235 2915 3239 2919
rect 3535 2915 3539 2919
rect 1871 2907 1875 2911
rect 2119 2904 2123 2908
rect 2199 2904 2203 2908
rect 2279 2904 2283 2908
rect 2359 2904 2363 2908
rect 2439 2904 2443 2908
rect 2519 2904 2523 2908
rect 2599 2904 2603 2908
rect 2687 2904 2691 2908
rect 2783 2904 2787 2908
rect 2903 2904 2907 2908
rect 3031 2904 3035 2908
rect 3175 2904 3179 2908
rect 3327 2904 3331 2908
rect 3487 2904 3491 2908
rect 3591 2907 3595 2911
rect 111 2881 115 2885
rect 151 2884 155 2888
rect 311 2884 315 2888
rect 471 2884 475 2888
rect 631 2884 635 2888
rect 783 2884 787 2888
rect 927 2884 931 2888
rect 1055 2884 1059 2888
rect 1175 2884 1179 2888
rect 1287 2884 1291 2888
rect 1391 2884 1395 2888
rect 1487 2884 1491 2888
rect 1591 2884 1595 2888
rect 1695 2884 1699 2888
rect 2083 2887 2087 2891
rect 2627 2887 2631 2891
rect 3227 2887 3231 2891
rect 1831 2881 1835 2885
rect 151 2871 155 2875
rect 219 2875 223 2879
rect 539 2875 543 2879
rect 699 2875 703 2879
rect 1015 2875 1019 2879
rect 1123 2875 1127 2879
rect 1255 2875 1259 2879
rect 1263 2875 1267 2879
rect 1463 2875 1467 2879
rect 1563 2875 1567 2879
rect 1667 2875 1671 2879
rect 1675 2875 1679 2879
rect 111 2864 115 2868
rect 531 2867 535 2871
rect 1831 2864 1835 2868
rect 1871 2857 1875 2861
rect 2047 2860 2051 2864
rect 2135 2860 2139 2864
rect 2239 2860 2243 2864
rect 2343 2860 2347 2864
rect 2463 2860 2467 2864
rect 2591 2860 2595 2864
rect 2727 2860 2731 2864
rect 2879 2860 2883 2864
rect 3031 2860 3035 2864
rect 3191 2860 3195 2864
rect 3359 2860 3363 2864
rect 3503 2860 3507 2864
rect 3591 2857 3595 2861
rect 2115 2851 2119 2855
rect 159 2846 163 2850
rect 319 2846 323 2850
rect 479 2846 483 2850
rect 639 2846 643 2850
rect 791 2846 795 2850
rect 935 2846 939 2850
rect 1063 2846 1067 2850
rect 1183 2846 1187 2850
rect 1295 2846 1299 2850
rect 1399 2846 1403 2850
rect 1495 2846 1499 2850
rect 1599 2846 1603 2850
rect 1703 2846 1707 2850
rect 1871 2840 1875 2844
rect 2195 2843 2199 2847
rect 2307 2851 2311 2855
rect 2411 2851 2415 2855
rect 2683 2851 2687 2855
rect 2795 2851 2799 2855
rect 2947 2851 2951 2855
rect 2959 2851 2963 2855
rect 3099 2851 3103 2855
rect 3439 2851 3443 2855
rect 2315 2843 2319 2847
rect 3563 2843 3567 2847
rect 219 2835 223 2839
rect 343 2835 344 2839
rect 344 2835 347 2839
rect 539 2835 543 2839
rect 699 2835 703 2839
rect 855 2835 859 2839
rect 1007 2835 1011 2839
rect 1015 2835 1019 2839
rect 1123 2835 1127 2839
rect 1255 2835 1259 2839
rect 1427 2835 1428 2839
rect 1428 2835 1431 2839
rect 1463 2835 1467 2839
rect 1563 2835 1567 2839
rect 1667 2835 1671 2839
rect 3591 2840 3595 2844
rect 151 2819 155 2823
rect 195 2819 199 2823
rect 299 2819 303 2823
rect 571 2819 575 2823
rect 587 2819 591 2823
rect 739 2819 743 2823
rect 1287 2827 1291 2831
rect 1203 2819 1207 2823
rect 1231 2819 1235 2823
rect 1435 2819 1436 2823
rect 1436 2819 1439 2823
rect 1459 2819 1463 2823
rect 1579 2819 1583 2823
rect 1715 2819 1719 2823
rect 2055 2822 2059 2826
rect 2143 2822 2147 2826
rect 2247 2822 2251 2826
rect 2351 2822 2355 2826
rect 2471 2822 2475 2826
rect 2599 2822 2603 2826
rect 2735 2822 2739 2826
rect 2887 2822 2891 2826
rect 3039 2822 3043 2826
rect 3199 2822 3203 2826
rect 3367 2822 3371 2826
rect 3511 2822 3515 2826
rect 143 2810 147 2814
rect 247 2810 251 2814
rect 383 2810 387 2814
rect 535 2810 539 2814
rect 687 2810 691 2814
rect 847 2810 851 2814
rect 999 2810 1003 2814
rect 1143 2810 1147 2814
rect 1279 2810 1283 2814
rect 1407 2810 1411 2814
rect 1527 2810 1531 2814
rect 1647 2810 1651 2814
rect 1751 2810 1755 2814
rect 2083 2811 2084 2815
rect 2084 2811 2087 2815
rect 2115 2811 2119 2815
rect 2307 2811 2311 2815
rect 2411 2811 2415 2815
rect 2495 2811 2496 2815
rect 2496 2811 2499 2815
rect 2627 2811 2628 2815
rect 2628 2811 2631 2815
rect 2683 2811 2687 2815
rect 2795 2811 2799 2815
rect 3099 2811 3103 2815
rect 3227 2811 3228 2815
rect 3228 2811 3231 2815
rect 3391 2811 3392 2815
rect 3392 2811 3395 2815
rect 3535 2811 3536 2815
rect 3536 2811 3539 2815
rect 111 2792 115 2796
rect 1831 2792 1835 2796
rect 195 2783 199 2787
rect 299 2783 303 2787
rect 587 2783 591 2787
rect 739 2783 743 2787
rect 855 2783 859 2787
rect 1007 2783 1011 2787
rect 1231 2783 1235 2787
rect 1287 2783 1291 2787
rect 1459 2783 1463 2787
rect 1579 2783 1583 2787
rect 1715 2783 1719 2787
rect 2023 2795 2027 2799
rect 1955 2787 1959 2791
rect 2195 2787 2196 2791
rect 2196 2787 2199 2791
rect 2219 2787 2223 2791
rect 2419 2787 2423 2791
rect 2667 2787 2668 2791
rect 2668 2787 2671 2791
rect 2691 2787 2695 2791
rect 2843 2787 2847 2791
rect 2995 2787 2999 2791
rect 3139 2787 3143 2791
rect 3443 2787 3447 2791
rect 3563 2787 3567 2791
rect 111 2775 115 2779
rect 135 2772 139 2776
rect 239 2772 243 2776
rect 375 2772 379 2776
rect 527 2772 531 2776
rect 679 2772 683 2776
rect 839 2772 843 2776
rect 991 2772 995 2776
rect 1135 2772 1139 2776
rect 1271 2772 1275 2776
rect 1399 2772 1403 2776
rect 1519 2772 1523 2776
rect 1639 2772 1643 2776
rect 1743 2772 1747 2776
rect 1831 2775 1835 2779
rect 1903 2778 1907 2782
rect 2015 2778 2019 2782
rect 2167 2778 2171 2782
rect 2327 2778 2331 2782
rect 2487 2778 2491 2782
rect 2639 2778 2643 2782
rect 2791 2778 2795 2782
rect 2943 2778 2947 2782
rect 3087 2778 3091 2782
rect 3231 2778 3235 2782
rect 3383 2778 3387 2782
rect 3511 2778 3515 2782
rect 1871 2760 1875 2764
rect 395 2755 396 2759
rect 396 2755 399 2759
rect 1731 2755 1735 2759
rect 3591 2760 3595 2764
rect 1955 2751 1959 2755
rect 2067 2751 2071 2755
rect 2219 2751 2223 2755
rect 2359 2751 2363 2755
rect 2495 2751 2499 2755
rect 2691 2751 2695 2755
rect 2843 2751 2847 2755
rect 2995 2751 2999 2755
rect 3139 2751 3143 2755
rect 3391 2751 3395 2755
rect 3535 2751 3539 2755
rect 1871 2743 1875 2747
rect 1895 2740 1899 2744
rect 2007 2740 2011 2744
rect 2159 2740 2163 2744
rect 2319 2740 2323 2744
rect 2479 2740 2483 2744
rect 2631 2740 2635 2744
rect 2783 2740 2787 2744
rect 2935 2740 2939 2744
rect 3079 2740 3083 2744
rect 3223 2740 3227 2744
rect 3375 2740 3379 2744
rect 3503 2740 3507 2744
rect 3591 2743 3595 2747
rect 111 2721 115 2725
rect 135 2724 139 2728
rect 231 2724 235 2728
rect 367 2724 371 2728
rect 511 2724 515 2728
rect 663 2724 667 2728
rect 815 2724 819 2728
rect 975 2724 979 2728
rect 1135 2724 1139 2728
rect 1287 2724 1291 2728
rect 1447 2724 1451 2728
rect 1607 2724 1611 2728
rect 1743 2724 1747 2728
rect 1831 2721 1835 2725
rect 3139 2723 3143 2727
rect 203 2715 207 2719
rect 299 2715 303 2719
rect 579 2715 583 2719
rect 731 2715 735 2719
rect 1071 2715 1075 2719
rect 1203 2715 1207 2719
rect 1223 2715 1227 2719
rect 1355 2715 1359 2719
rect 111 2704 115 2708
rect 195 2707 199 2711
rect 571 2707 575 2711
rect 1739 2711 1743 2715
rect 1843 2715 1847 2719
rect 1831 2704 1835 2708
rect 1871 2693 1875 2697
rect 1895 2696 1899 2700
rect 2103 2696 2107 2700
rect 2327 2696 2331 2700
rect 2535 2696 2539 2700
rect 2735 2696 2739 2700
rect 2911 2696 2915 2700
rect 3071 2696 3075 2700
rect 3223 2696 3227 2700
rect 3375 2696 3379 2700
rect 3503 2696 3507 2700
rect 3591 2693 3595 2697
rect 143 2686 147 2690
rect 239 2686 243 2690
rect 375 2686 379 2690
rect 519 2686 523 2690
rect 671 2686 675 2690
rect 823 2686 827 2690
rect 983 2686 987 2690
rect 1143 2686 1147 2690
rect 1295 2686 1299 2690
rect 1455 2686 1459 2690
rect 1615 2686 1619 2690
rect 1751 2686 1755 2690
rect 203 2675 207 2679
rect 299 2675 303 2679
rect 395 2675 399 2679
rect 579 2675 583 2679
rect 731 2675 735 2679
rect 843 2675 847 2679
rect 1007 2675 1008 2679
rect 1008 2675 1011 2679
rect 1071 2675 1075 2679
rect 1355 2675 1359 2679
rect 1559 2675 1563 2679
rect 1731 2675 1735 2679
rect 1739 2675 1743 2679
rect 1871 2676 1875 2680
rect 2023 2679 2027 2683
rect 2455 2687 2459 2691
rect 2479 2687 2483 2691
rect 3015 2687 3019 2691
rect 3171 2687 3175 2691
rect 3323 2687 3327 2691
rect 3443 2687 3447 2691
rect 3571 2687 3575 2691
rect 3591 2676 3595 2680
rect 195 2655 199 2659
rect 331 2655 335 2659
rect 587 2655 591 2659
rect 991 2655 995 2659
rect 1003 2655 1007 2659
rect 1155 2655 1159 2659
rect 1391 2655 1395 2659
rect 1543 2655 1547 2659
rect 1903 2658 1907 2662
rect 2111 2658 2115 2662
rect 2335 2658 2339 2662
rect 2543 2658 2547 2662
rect 2743 2658 2747 2662
rect 2919 2658 2923 2662
rect 3079 2658 3083 2662
rect 3231 2658 3235 2662
rect 3383 2658 3387 2662
rect 3511 2658 3515 2662
rect 143 2646 147 2650
rect 279 2646 283 2650
rect 447 2646 451 2650
rect 623 2646 627 2650
rect 791 2646 795 2650
rect 951 2646 955 2650
rect 1103 2646 1107 2650
rect 1247 2646 1251 2650
rect 1399 2646 1403 2650
rect 1551 2646 1555 2650
rect 1843 2647 1847 2651
rect 2359 2647 2360 2651
rect 2360 2647 2363 2651
rect 2455 2647 2459 2651
rect 2771 2647 2772 2651
rect 2772 2647 2775 2651
rect 3015 2647 3019 2651
rect 3171 2647 3175 2651
rect 3323 2647 3327 2651
rect 3535 2647 3536 2651
rect 3536 2647 3539 2651
rect 111 2628 115 2632
rect 1831 2628 1835 2632
rect 1931 2627 1932 2631
rect 1932 2627 1935 2631
rect 1955 2627 1959 2631
rect 2255 2627 2259 2631
rect 2315 2627 2319 2631
rect 3295 2627 3299 2631
rect 3303 2627 3307 2631
rect 331 2619 335 2623
rect 843 2619 847 2623
rect 1003 2619 1007 2623
rect 1155 2619 1159 2623
rect 1391 2619 1395 2623
rect 1543 2619 1547 2623
rect 1559 2619 1563 2623
rect 1903 2618 1907 2622
rect 2055 2618 2059 2622
rect 2263 2618 2267 2622
rect 2495 2618 2499 2622
rect 2751 2618 2755 2622
rect 3015 2618 3019 2622
rect 3287 2618 3291 2622
rect 111 2611 115 2615
rect 135 2608 139 2612
rect 271 2608 275 2612
rect 439 2608 443 2612
rect 615 2608 619 2612
rect 783 2608 787 2612
rect 943 2608 947 2612
rect 1095 2608 1099 2612
rect 1239 2608 1243 2612
rect 1391 2608 1395 2612
rect 1543 2608 1547 2612
rect 1831 2611 1835 2615
rect 1871 2600 1875 2604
rect 3591 2600 3595 2604
rect 403 2591 407 2595
rect 1955 2591 1959 2595
rect 2255 2591 2259 2595
rect 2315 2591 2319 2595
rect 3039 2591 3043 2595
rect 3295 2591 3299 2595
rect 1871 2583 1875 2587
rect 1895 2580 1899 2584
rect 2047 2580 2051 2584
rect 2255 2580 2259 2584
rect 2487 2580 2491 2584
rect 2743 2580 2747 2584
rect 3007 2580 3011 2584
rect 3279 2580 3283 2584
rect 3591 2583 3595 2587
rect 111 2557 115 2561
rect 135 2560 139 2564
rect 223 2560 227 2564
rect 367 2560 371 2564
rect 527 2560 531 2564
rect 703 2560 707 2564
rect 879 2560 883 2564
rect 1047 2560 1051 2564
rect 1207 2560 1211 2564
rect 1359 2560 1363 2564
rect 1511 2560 1515 2564
rect 1671 2560 1675 2564
rect 2659 2563 2663 2567
rect 1831 2557 1835 2561
rect 203 2551 207 2555
rect 291 2551 295 2555
rect 595 2551 599 2555
rect 771 2551 775 2555
rect 991 2551 995 2555
rect 1115 2551 1119 2555
rect 1275 2551 1279 2555
rect 1427 2551 1431 2555
rect 1579 2551 1583 2555
rect 111 2540 115 2544
rect 195 2543 199 2547
rect 587 2543 591 2547
rect 1831 2540 1835 2544
rect 1871 2533 1875 2537
rect 1895 2536 1899 2540
rect 2007 2536 2011 2540
rect 2159 2536 2163 2540
rect 2319 2536 2323 2540
rect 2471 2536 2475 2540
rect 2623 2536 2627 2540
rect 2759 2536 2763 2540
rect 2887 2536 2891 2540
rect 3007 2536 3011 2540
rect 3119 2536 3123 2540
rect 3223 2536 3227 2540
rect 3319 2536 3323 2540
rect 3423 2536 3427 2540
rect 3503 2536 3507 2540
rect 3591 2533 3595 2537
rect 1963 2527 1967 2531
rect 143 2522 147 2526
rect 231 2522 235 2526
rect 375 2522 379 2526
rect 535 2522 539 2526
rect 711 2522 715 2526
rect 887 2522 891 2526
rect 1055 2522 1059 2526
rect 1215 2522 1219 2526
rect 1367 2522 1371 2526
rect 1519 2522 1523 2526
rect 2107 2527 2111 2531
rect 2263 2527 2267 2531
rect 2419 2527 2423 2531
rect 2427 2527 2431 2531
rect 2715 2527 2719 2531
rect 1679 2522 1683 2526
rect 1871 2516 1875 2520
rect 2683 2519 2687 2523
rect 2955 2527 2959 2531
rect 3075 2527 3079 2531
rect 3291 2527 3295 2531
rect 3387 2527 3391 2531
rect 3303 2519 3307 2523
rect 3563 2519 3567 2523
rect 203 2511 207 2515
rect 291 2511 295 2515
rect 403 2511 404 2515
rect 404 2511 407 2515
rect 595 2511 599 2515
rect 771 2511 775 2515
rect 935 2511 939 2515
rect 1115 2511 1119 2515
rect 1275 2511 1279 2515
rect 1427 2511 1431 2515
rect 1579 2511 1583 2515
rect 3591 2516 3595 2520
rect 1703 2511 1704 2515
rect 1704 2511 1707 2515
rect 195 2495 199 2499
rect 215 2495 219 2499
rect 275 2495 279 2499
rect 355 2495 359 2499
rect 443 2495 447 2499
rect 563 2495 567 2499
rect 699 2495 703 2499
rect 835 2495 839 2499
rect 1135 2495 1139 2499
rect 1143 2495 1147 2499
rect 1243 2495 1247 2499
rect 1423 2495 1427 2499
rect 1483 2495 1487 2499
rect 1603 2495 1607 2499
rect 1903 2498 1907 2502
rect 2015 2498 2019 2502
rect 2167 2498 2171 2502
rect 2327 2498 2331 2502
rect 2479 2498 2483 2502
rect 2631 2498 2635 2502
rect 2767 2498 2771 2502
rect 2895 2498 2899 2502
rect 3015 2498 3019 2502
rect 3127 2498 3131 2502
rect 3231 2498 3235 2502
rect 3327 2498 3331 2502
rect 3431 2498 3435 2502
rect 3511 2498 3515 2502
rect 143 2486 147 2490
rect 223 2486 227 2490
rect 303 2486 307 2490
rect 391 2486 395 2490
rect 511 2486 515 2490
rect 647 2486 651 2490
rect 783 2486 787 2490
rect 927 2486 931 2490
rect 1063 2486 1067 2490
rect 1191 2486 1195 2490
rect 1311 2486 1315 2490
rect 1431 2486 1435 2490
rect 1551 2486 1555 2490
rect 1671 2486 1675 2490
rect 1931 2487 1932 2491
rect 1932 2487 1935 2491
rect 1963 2487 1967 2491
rect 2107 2487 2111 2491
rect 2263 2487 2267 2491
rect 2419 2487 2423 2491
rect 2683 2487 2687 2491
rect 2715 2487 2719 2491
rect 2955 2487 2959 2491
rect 3039 2487 3040 2491
rect 3040 2487 3043 2491
rect 111 2468 115 2472
rect 1831 2468 1835 2472
rect 2427 2475 2431 2479
rect 3291 2487 3295 2491
rect 3387 2487 3391 2491
rect 3411 2487 3415 2491
rect 3571 2487 3575 2491
rect 2051 2467 2055 2471
rect 2179 2467 2183 2471
rect 2315 2467 2319 2471
rect 2459 2467 2463 2471
rect 2803 2467 2807 2471
rect 2811 2467 2815 2471
rect 3075 2467 3079 2471
rect 3419 2467 3423 2471
rect 3563 2467 3567 2471
rect 215 2459 219 2463
rect 275 2459 279 2463
rect 355 2459 359 2463
rect 443 2459 447 2463
rect 563 2459 567 2463
rect 699 2459 703 2463
rect 835 2459 839 2463
rect 935 2459 939 2463
rect 1143 2459 1147 2463
rect 1243 2459 1247 2463
rect 1423 2459 1427 2463
rect 1483 2459 1487 2463
rect 1603 2459 1607 2463
rect 1703 2459 1707 2463
rect 1999 2458 2003 2462
rect 2127 2458 2131 2462
rect 2263 2458 2267 2462
rect 2407 2458 2411 2462
rect 2551 2458 2555 2462
rect 2703 2458 2707 2462
rect 2863 2458 2867 2462
rect 3023 2458 3027 2462
rect 3191 2458 3195 2462
rect 3359 2458 3363 2462
rect 3511 2458 3515 2462
rect 111 2451 115 2455
rect 135 2448 139 2452
rect 215 2448 219 2452
rect 295 2448 299 2452
rect 383 2448 387 2452
rect 503 2448 507 2452
rect 639 2448 643 2452
rect 775 2448 779 2452
rect 919 2448 923 2452
rect 1055 2448 1059 2452
rect 1183 2448 1187 2452
rect 1303 2448 1307 2452
rect 1423 2448 1427 2452
rect 1543 2448 1547 2452
rect 1663 2448 1667 2452
rect 1831 2451 1835 2455
rect 1871 2440 1875 2444
rect 3591 2440 3595 2444
rect 2051 2431 2055 2435
rect 2179 2431 2183 2435
rect 2315 2431 2319 2435
rect 2459 2431 2463 2435
rect 2811 2431 2815 2435
rect 2915 2431 2919 2435
rect 3199 2431 3203 2435
rect 3411 2431 3415 2435
rect 3535 2431 3539 2435
rect 1871 2423 1875 2427
rect 1991 2420 1995 2424
rect 2119 2420 2123 2424
rect 2255 2420 2259 2424
rect 2399 2420 2403 2424
rect 2543 2420 2547 2424
rect 2695 2420 2699 2424
rect 2855 2420 2859 2424
rect 3015 2420 3019 2424
rect 3183 2420 3187 2424
rect 3351 2420 3355 2424
rect 3503 2420 3507 2424
rect 3591 2423 3595 2427
rect 2479 2403 2483 2407
rect 111 2389 115 2393
rect 1063 2392 1067 2396
rect 1143 2392 1147 2396
rect 1223 2392 1227 2396
rect 1303 2392 1307 2396
rect 1383 2392 1387 2396
rect 1463 2392 1467 2396
rect 1831 2389 1835 2393
rect 1135 2383 1139 2387
rect 1211 2383 1215 2387
rect 1291 2383 1295 2387
rect 1371 2383 1375 2387
rect 1451 2383 1455 2387
rect 1471 2379 1475 2383
rect 111 2372 115 2376
rect 1831 2372 1835 2376
rect 1871 2369 1875 2373
rect 2143 2372 2147 2376
rect 2239 2372 2243 2376
rect 2343 2372 2347 2376
rect 2455 2372 2459 2376
rect 2575 2372 2579 2376
rect 2703 2372 2707 2376
rect 2847 2372 2851 2376
rect 3007 2372 3011 2376
rect 3175 2372 3179 2376
rect 3351 2372 3355 2376
rect 3503 2372 3507 2376
rect 3591 2369 3595 2373
rect 2215 2363 2219 2367
rect 2539 2363 2543 2367
rect 1071 2354 1075 2358
rect 1151 2354 1155 2358
rect 1231 2354 1235 2358
rect 1311 2354 1315 2358
rect 1391 2354 1395 2358
rect 1471 2354 1475 2358
rect 1871 2352 1875 2356
rect 2307 2355 2311 2359
rect 2771 2363 2775 2367
rect 3115 2363 3119 2367
rect 3123 2363 3127 2367
rect 3419 2363 3423 2367
rect 3571 2363 3575 2367
rect 3591 2352 3595 2356
rect 1135 2343 1139 2347
rect 1211 2343 1215 2347
rect 1291 2343 1295 2347
rect 1371 2343 1375 2347
rect 1451 2343 1455 2347
rect 447 2323 451 2327
rect 527 2323 531 2327
rect 607 2323 611 2327
rect 687 2323 691 2327
rect 767 2323 771 2327
rect 927 2331 931 2335
rect 1327 2335 1331 2339
rect 2151 2334 2155 2338
rect 2247 2334 2251 2338
rect 2351 2334 2355 2338
rect 2463 2334 2467 2338
rect 2583 2334 2587 2338
rect 2711 2334 2715 2338
rect 2855 2334 2859 2338
rect 3015 2334 3019 2338
rect 3183 2334 3187 2338
rect 3359 2334 3363 2338
rect 3511 2334 3515 2338
rect 863 2323 864 2327
rect 864 2323 867 2327
rect 891 2323 895 2327
rect 1043 2323 1047 2327
rect 1051 2323 1055 2327
rect 1131 2323 1135 2327
rect 1211 2323 1215 2327
rect 1291 2323 1295 2327
rect 2179 2323 2180 2327
rect 2180 2323 2183 2327
rect 2215 2323 2219 2327
rect 2539 2323 2543 2327
rect 2771 2323 2775 2327
rect 2883 2323 2884 2327
rect 2884 2323 2887 2327
rect 2915 2323 2919 2327
rect 3115 2323 3119 2327
rect 3419 2323 3423 2327
rect 3535 2323 3536 2327
rect 3536 2323 3539 2327
rect 359 2314 363 2318
rect 439 2314 443 2318
rect 519 2314 523 2318
rect 599 2314 603 2318
rect 679 2314 683 2318
rect 759 2314 763 2318
rect 839 2314 843 2318
rect 919 2314 923 2318
rect 999 2314 1003 2318
rect 1079 2314 1083 2318
rect 1159 2314 1163 2318
rect 1239 2314 1243 2318
rect 1319 2314 1323 2318
rect 2307 2307 2308 2311
rect 2308 2307 2311 2311
rect 2331 2307 2335 2311
rect 2411 2307 2415 2311
rect 2491 2307 2495 2311
rect 2687 2307 2691 2311
rect 2943 2315 2947 2319
rect 2811 2307 2815 2311
rect 2899 2307 2903 2311
rect 111 2296 115 2300
rect 1831 2296 1835 2300
rect 2279 2298 2283 2302
rect 2359 2298 2363 2302
rect 2439 2298 2443 2302
rect 2519 2298 2523 2302
rect 2599 2298 2603 2302
rect 2679 2298 2683 2302
rect 2759 2298 2763 2302
rect 2847 2298 2851 2302
rect 2935 2298 2939 2302
rect 407 2287 411 2291
rect 447 2287 451 2291
rect 527 2287 531 2291
rect 607 2287 611 2291
rect 687 2287 691 2291
rect 767 2287 771 2291
rect 891 2287 895 2291
rect 927 2287 931 2291
rect 1051 2287 1055 2291
rect 1131 2287 1135 2291
rect 1211 2287 1215 2291
rect 1291 2287 1295 2291
rect 1327 2287 1331 2291
rect 111 2279 115 2283
rect 351 2276 355 2280
rect 431 2276 435 2280
rect 511 2276 515 2280
rect 591 2276 595 2280
rect 671 2276 675 2280
rect 751 2276 755 2280
rect 831 2276 835 2280
rect 911 2276 915 2280
rect 991 2276 995 2280
rect 1071 2276 1075 2280
rect 1151 2276 1155 2280
rect 1231 2276 1235 2280
rect 1311 2276 1315 2280
rect 1831 2279 1835 2283
rect 1871 2280 1875 2284
rect 3591 2280 3595 2284
rect 2331 2271 2335 2275
rect 2411 2271 2415 2275
rect 2491 2271 2495 2275
rect 2631 2271 2635 2275
rect 2687 2271 2691 2275
rect 2811 2271 2815 2275
rect 2899 2271 2903 2275
rect 2943 2271 2947 2275
rect 1871 2263 1875 2267
rect 2271 2260 2275 2264
rect 1043 2255 1047 2259
rect 2351 2260 2355 2264
rect 2431 2260 2435 2264
rect 2511 2260 2515 2264
rect 2591 2260 2595 2264
rect 2671 2260 2675 2264
rect 2751 2260 2755 2264
rect 2839 2260 2843 2264
rect 2927 2260 2931 2264
rect 3591 2263 3595 2267
rect 1243 2255 1247 2259
rect 2359 2243 2363 2247
rect 111 2229 115 2233
rect 375 2232 379 2236
rect 455 2232 459 2236
rect 535 2232 539 2236
rect 615 2232 619 2236
rect 695 2232 699 2236
rect 775 2232 779 2236
rect 855 2232 859 2236
rect 935 2232 939 2236
rect 1015 2232 1019 2236
rect 1095 2232 1099 2236
rect 1175 2232 1179 2236
rect 1255 2232 1259 2236
rect 1831 2229 1835 2233
rect 443 2223 447 2227
rect 527 2223 531 2227
rect 683 2223 687 2227
rect 763 2223 767 2227
rect 111 2212 115 2216
rect 515 2215 519 2219
rect 863 2219 867 2223
rect 923 2223 927 2227
rect 1003 2223 1007 2227
rect 1083 2223 1087 2227
rect 1243 2223 1247 2227
rect 1235 2215 1239 2219
rect 1831 2212 1835 2216
rect 1871 2213 1875 2217
rect 2311 2216 2315 2220
rect 2399 2216 2403 2220
rect 2495 2216 2499 2220
rect 2599 2216 2603 2220
rect 2719 2216 2723 2220
rect 2855 2216 2859 2220
rect 3007 2216 3011 2220
rect 3175 2216 3179 2220
rect 3351 2216 3355 2220
rect 3503 2216 3507 2220
rect 3591 2213 3595 2217
rect 2379 2207 2383 2211
rect 2471 2207 2475 2211
rect 2563 2207 2567 2211
rect 2679 2207 2683 2211
rect 2787 2207 2791 2211
rect 3075 2207 3079 2211
rect 3083 2207 3087 2211
rect 3419 2207 3423 2211
rect 383 2194 387 2198
rect 463 2194 467 2198
rect 543 2194 547 2198
rect 623 2194 627 2198
rect 703 2194 707 2198
rect 783 2194 787 2198
rect 863 2194 867 2198
rect 943 2194 947 2198
rect 1023 2194 1027 2198
rect 1103 2194 1107 2198
rect 1183 2194 1187 2198
rect 1263 2194 1267 2198
rect 1871 2196 1875 2200
rect 3563 2199 3567 2203
rect 3591 2196 3595 2200
rect 407 2183 408 2187
rect 408 2183 411 2187
rect 443 2183 447 2187
rect 515 2183 519 2187
rect 683 2183 687 2187
rect 763 2183 767 2187
rect 887 2183 888 2187
rect 888 2183 891 2187
rect 923 2183 927 2187
rect 1003 2183 1007 2187
rect 1083 2183 1087 2187
rect 1235 2183 1239 2187
rect 747 2175 751 2179
rect 2319 2178 2323 2182
rect 2407 2178 2411 2182
rect 2503 2178 2507 2182
rect 2607 2178 2611 2182
rect 2727 2178 2731 2182
rect 2863 2178 2867 2182
rect 3015 2178 3019 2182
rect 3183 2178 3187 2182
rect 3359 2178 3363 2182
rect 3511 2178 3515 2182
rect 2359 2167 2363 2171
rect 2379 2167 2383 2171
rect 2471 2167 2475 2171
rect 2631 2167 2632 2171
rect 2632 2167 2635 2171
rect 2679 2167 2683 2171
rect 2787 2167 2791 2171
rect 3075 2167 3079 2171
rect 3387 2167 3388 2171
rect 3388 2167 3391 2171
rect 3571 2167 3575 2171
rect 415 2159 419 2163
rect 511 2159 515 2163
rect 527 2159 528 2163
rect 528 2159 531 2163
rect 635 2159 639 2163
rect 651 2159 655 2163
rect 739 2159 743 2163
rect 959 2159 963 2163
rect 1047 2159 1051 2163
rect 1135 2159 1139 2163
rect 1231 2159 1235 2163
rect 1243 2159 1247 2163
rect 311 2150 315 2154
rect 407 2150 411 2154
rect 503 2150 507 2154
rect 599 2150 603 2154
rect 687 2150 691 2154
rect 775 2150 779 2154
rect 863 2150 867 2154
rect 951 2150 955 2154
rect 1039 2150 1043 2154
rect 1127 2150 1131 2154
rect 1223 2150 1227 2154
rect 1991 2151 1995 2155
rect 2399 2159 2403 2163
rect 2051 2151 2055 2155
rect 2163 2151 2167 2155
rect 2299 2151 2303 2155
rect 2563 2151 2567 2155
rect 2735 2151 2739 2155
rect 2747 2151 2751 2155
rect 2899 2151 2903 2155
rect 3059 2151 3063 2155
rect 3227 2151 3231 2155
rect 3563 2151 3567 2155
rect 1903 2142 1907 2146
rect 1983 2142 1987 2146
rect 2111 2142 2115 2146
rect 2247 2142 2251 2146
rect 2391 2142 2395 2146
rect 2543 2142 2547 2146
rect 2695 2142 2699 2146
rect 2847 2142 2851 2146
rect 3007 2142 3011 2146
rect 3175 2142 3179 2146
rect 3351 2142 3355 2146
rect 3511 2142 3515 2146
rect 111 2132 115 2136
rect 1831 2132 1835 2136
rect 415 2123 419 2127
rect 511 2123 515 2127
rect 651 2123 655 2127
rect 739 2123 743 2127
rect 747 2123 751 2127
rect 887 2123 891 2127
rect 959 2123 963 2127
rect 1047 2123 1051 2127
rect 1135 2123 1139 2127
rect 1231 2123 1235 2127
rect 1871 2124 1875 2128
rect 3591 2124 3595 2128
rect 111 2115 115 2119
rect 303 2112 307 2116
rect 399 2112 403 2116
rect 495 2112 499 2116
rect 591 2112 595 2116
rect 679 2112 683 2116
rect 767 2112 771 2116
rect 855 2112 859 2116
rect 943 2112 947 2116
rect 1031 2112 1035 2116
rect 1119 2112 1123 2116
rect 1215 2112 1219 2116
rect 1831 2115 1835 2119
rect 1991 2115 1995 2119
rect 2163 2115 2167 2119
rect 2299 2115 2303 2119
rect 2399 2115 2403 2119
rect 2747 2115 2751 2119
rect 2899 2115 2903 2119
rect 3059 2115 3063 2119
rect 3227 2115 3231 2119
rect 3535 2115 3539 2119
rect 1871 2107 1875 2111
rect 1895 2104 1899 2108
rect 1975 2104 1979 2108
rect 2103 2104 2107 2108
rect 2239 2104 2243 2108
rect 2383 2104 2387 2108
rect 2535 2104 2539 2108
rect 2687 2104 2691 2108
rect 2839 2104 2843 2108
rect 2999 2104 3003 2108
rect 3167 2104 3171 2108
rect 3343 2104 3347 2108
rect 3503 2104 3507 2108
rect 3591 2107 3595 2111
rect 243 2095 247 2099
rect 1779 2087 1783 2091
rect 2483 2087 2487 2091
rect 3307 2087 3311 2091
rect 111 2053 115 2057
rect 207 2056 211 2060
rect 327 2056 331 2060
rect 447 2056 451 2060
rect 575 2056 579 2060
rect 703 2056 707 2060
rect 823 2056 827 2060
rect 943 2056 947 2060
rect 1063 2056 1067 2060
rect 1175 2056 1179 2060
rect 1279 2056 1283 2060
rect 1375 2056 1379 2060
rect 1471 2056 1475 2060
rect 1567 2056 1571 2060
rect 1663 2056 1667 2060
rect 1743 2056 1747 2060
rect 1831 2053 1835 2057
rect 275 2047 279 2051
rect 395 2047 399 2051
rect 643 2047 647 2051
rect 771 2047 775 2051
rect 1031 2047 1035 2051
rect 1131 2047 1135 2051
rect 1243 2047 1247 2051
rect 1347 2047 1351 2051
rect 1443 2047 1447 2051
rect 1539 2047 1543 2051
rect 1635 2047 1639 2051
rect 1731 2047 1735 2051
rect 1871 2049 1875 2053
rect 1967 2052 1971 2056
rect 2215 2052 2219 2056
rect 2447 2052 2451 2056
rect 2655 2052 2659 2056
rect 2839 2052 2843 2056
rect 2999 2052 3003 2056
rect 3143 2052 3147 2056
rect 3271 2052 3275 2056
rect 3399 2052 3403 2056
rect 3503 2052 3507 2056
rect 3591 2049 3595 2053
rect 111 2036 115 2040
rect 387 2039 391 2043
rect 635 2039 639 2043
rect 1339 2039 1343 2043
rect 2051 2043 2055 2047
rect 2283 2043 2287 2047
rect 2755 2043 2759 2047
rect 2943 2043 2947 2047
rect 3079 2043 3083 2047
rect 3087 2043 3091 2047
rect 3211 2043 3215 2047
rect 3387 2043 3391 2047
rect 1831 2036 1835 2040
rect 1871 2032 1875 2036
rect 2275 2035 2279 2039
rect 3563 2035 3567 2039
rect 3591 2032 3595 2036
rect 215 2018 219 2022
rect 335 2018 339 2022
rect 455 2018 459 2022
rect 583 2018 587 2022
rect 711 2018 715 2022
rect 831 2018 835 2022
rect 951 2018 955 2022
rect 1071 2018 1075 2022
rect 1183 2018 1187 2022
rect 1287 2018 1291 2022
rect 1383 2018 1387 2022
rect 1479 2018 1483 2022
rect 1575 2018 1579 2022
rect 1671 2018 1675 2022
rect 1751 2018 1755 2022
rect 1975 2014 1979 2018
rect 2223 2014 2227 2018
rect 2455 2014 2459 2018
rect 2663 2014 2667 2018
rect 2847 2014 2851 2018
rect 3007 2014 3011 2018
rect 3151 2014 3155 2018
rect 3279 2014 3283 2018
rect 3407 2014 3411 2018
rect 3511 2014 3515 2018
rect 243 2007 244 2011
rect 244 2007 247 2011
rect 275 2007 279 2011
rect 387 2007 391 2011
rect 643 2007 647 2011
rect 771 2007 775 2011
rect 855 2007 856 2011
rect 856 2007 859 2011
rect 1023 2007 1027 2011
rect 1031 2007 1035 2011
rect 1131 2007 1135 2011
rect 1347 2007 1351 2011
rect 1443 2007 1447 2011
rect 1539 2007 1543 2011
rect 1635 2007 1639 2011
rect 1731 2007 1735 2011
rect 1779 2007 1780 2011
rect 1780 2007 1783 2011
rect 1999 2003 2000 2007
rect 2000 2003 2003 2007
rect 2283 2003 2287 2007
rect 2483 2003 2484 2007
rect 2484 2003 2487 2007
rect 2687 2003 2688 2007
rect 2688 2003 2691 2007
rect 2755 2003 2759 2007
rect 2943 2003 2947 2007
rect 359 1991 363 1995
rect 395 1991 399 1995
rect 535 1991 539 1995
rect 571 1991 575 1995
rect 739 1991 743 1995
rect 1175 1991 1179 1995
rect 1219 1991 1223 1995
rect 1339 1991 1340 1995
rect 1340 1991 1343 1995
rect 1363 1991 1367 1995
rect 1499 1991 1503 1995
rect 1635 1991 1639 1995
rect 2087 1991 2091 1995
rect 2207 1991 2211 1995
rect 2223 1987 2227 1991
rect 2275 1991 2279 1995
rect 2591 1991 2595 1995
rect 2751 1991 2755 1995
rect 2927 1991 2931 1995
rect 3167 1999 3171 2003
rect 3211 2003 3215 2007
rect 3307 2003 3308 2007
rect 3308 2003 3311 2007
rect 3451 2003 3455 2007
rect 3535 2003 3536 2007
rect 3536 2003 3539 2007
rect 3079 1991 3083 1995
rect 3171 1991 3175 1995
rect 3563 1991 3567 1995
rect 191 1982 195 1986
rect 351 1982 355 1986
rect 519 1982 523 1986
rect 687 1982 691 1986
rect 855 1982 859 1986
rect 1015 1982 1019 1986
rect 1167 1982 1171 1986
rect 1311 1982 1315 1986
rect 1447 1982 1451 1986
rect 1583 1982 1587 1986
rect 1719 1982 1723 1986
rect 1959 1982 1963 1986
rect 2079 1982 2083 1986
rect 2199 1982 2203 1986
rect 2319 1982 2323 1986
rect 2447 1982 2451 1986
rect 2583 1982 2587 1986
rect 2743 1982 2747 1986
rect 2919 1982 2923 1986
rect 3119 1982 3123 1986
rect 3327 1982 3331 1986
rect 3511 1982 3515 1986
rect 111 1964 115 1968
rect 1831 1964 1835 1968
rect 1871 1964 1875 1968
rect 3591 1964 3595 1968
rect 359 1955 363 1959
rect 571 1955 575 1959
rect 739 1955 743 1959
rect 863 1955 867 1959
rect 1023 1955 1027 1959
rect 1175 1955 1179 1959
rect 1363 1955 1367 1959
rect 1499 1955 1503 1959
rect 1635 1955 1639 1959
rect 1999 1955 2003 1959
rect 2087 1955 2091 1959
rect 2207 1955 2211 1959
rect 2591 1955 2595 1959
rect 2751 1955 2755 1959
rect 2927 1955 2931 1959
rect 3171 1955 3175 1959
rect 3179 1955 3183 1959
rect 3535 1955 3539 1959
rect 111 1947 115 1951
rect 183 1944 187 1948
rect 343 1944 347 1948
rect 511 1944 515 1948
rect 679 1944 683 1948
rect 847 1944 851 1948
rect 1007 1944 1011 1948
rect 1159 1944 1163 1948
rect 1303 1944 1307 1948
rect 1439 1944 1443 1948
rect 1575 1944 1579 1948
rect 1711 1944 1715 1948
rect 1831 1947 1835 1951
rect 1871 1947 1875 1951
rect 1951 1944 1955 1948
rect 2071 1944 2075 1948
rect 2191 1944 2195 1948
rect 2311 1944 2315 1948
rect 2439 1944 2443 1948
rect 2575 1944 2579 1948
rect 2735 1944 2739 1948
rect 2911 1944 2915 1948
rect 3111 1944 3115 1948
rect 3319 1944 3323 1948
rect 3503 1944 3507 1948
rect 3591 1947 3595 1951
rect 199 1927 200 1931
rect 200 1927 203 1931
rect 1727 1927 1728 1931
rect 1728 1927 1731 1931
rect 2303 1927 2307 1931
rect 2379 1927 2383 1931
rect 111 1893 115 1897
rect 135 1896 139 1900
rect 239 1896 243 1900
rect 375 1896 379 1900
rect 527 1896 531 1900
rect 687 1896 691 1900
rect 847 1896 851 1900
rect 1007 1896 1011 1900
rect 1159 1896 1163 1900
rect 1303 1896 1307 1900
rect 1455 1896 1459 1900
rect 1607 1896 1611 1900
rect 1831 1893 1835 1897
rect 211 1887 215 1891
rect 307 1887 311 1891
rect 355 1887 359 1891
rect 535 1883 539 1887
rect 595 1887 599 1891
rect 755 1887 759 1891
rect 1079 1887 1083 1891
rect 1227 1887 1231 1891
rect 1371 1887 1375 1891
rect 1523 1887 1527 1891
rect 1871 1889 1875 1893
rect 2063 1892 2067 1896
rect 2151 1892 2155 1896
rect 2239 1892 2243 1896
rect 2319 1892 2323 1896
rect 2399 1892 2403 1896
rect 2487 1892 2491 1896
rect 2575 1892 2579 1896
rect 2663 1892 2667 1896
rect 2759 1892 2763 1896
rect 2871 1892 2875 1896
rect 2991 1892 2995 1896
rect 3119 1892 3123 1896
rect 3247 1892 3251 1896
rect 3383 1892 3387 1896
rect 3503 1892 3507 1896
rect 3591 1889 3595 1893
rect 111 1876 115 1880
rect 1219 1879 1223 1883
rect 2131 1883 2135 1887
rect 2223 1883 2227 1887
rect 1831 1876 1835 1880
rect 2387 1883 2391 1887
rect 2467 1883 2471 1887
rect 2555 1883 2559 1887
rect 2643 1883 2647 1887
rect 2735 1883 2739 1887
rect 2955 1883 2959 1887
rect 3079 1883 3083 1887
rect 3195 1883 3199 1887
rect 3203 1883 3207 1887
rect 3451 1883 3455 1887
rect 3459 1883 3463 1887
rect 1871 1872 1875 1876
rect 2459 1875 2463 1879
rect 3591 1872 3595 1876
rect 143 1858 147 1862
rect 247 1858 251 1862
rect 383 1858 387 1862
rect 535 1858 539 1862
rect 695 1858 699 1862
rect 855 1858 859 1862
rect 1015 1858 1019 1862
rect 1167 1858 1171 1862
rect 1311 1858 1315 1862
rect 1463 1858 1467 1862
rect 1615 1858 1619 1862
rect 2071 1854 2075 1858
rect 2159 1854 2163 1858
rect 2247 1854 2251 1858
rect 2327 1854 2331 1858
rect 2407 1854 2411 1858
rect 2495 1854 2499 1858
rect 2583 1854 2587 1858
rect 2671 1854 2675 1858
rect 2767 1854 2771 1858
rect 2879 1854 2883 1858
rect 2999 1854 3003 1858
rect 3127 1854 3131 1858
rect 3255 1854 3259 1858
rect 3391 1854 3395 1858
rect 3511 1854 3515 1858
rect 199 1847 203 1851
rect 211 1847 215 1851
rect 307 1847 311 1851
rect 595 1847 599 1851
rect 755 1847 759 1851
rect 879 1847 880 1851
rect 880 1847 883 1851
rect 1039 1847 1040 1851
rect 1040 1847 1043 1851
rect 1079 1847 1083 1851
rect 1371 1847 1375 1851
rect 1523 1847 1527 1851
rect 1727 1847 1731 1851
rect 2095 1843 2096 1847
rect 2096 1843 2099 1847
rect 2131 1843 2135 1847
rect 2303 1843 2307 1847
rect 2379 1843 2383 1847
rect 2387 1843 2391 1847
rect 2467 1843 2471 1847
rect 2555 1843 2559 1847
rect 2643 1843 2647 1847
rect 2735 1843 2739 1847
rect 2955 1843 2959 1847
rect 3079 1843 3083 1847
rect 3195 1843 3199 1847
rect 3459 1843 3463 1847
rect 3535 1843 3536 1847
rect 3536 1843 3539 1847
rect 295 1831 299 1835
rect 355 1831 359 1835
rect 487 1831 491 1835
rect 523 1831 527 1835
rect 715 1831 719 1835
rect 1103 1831 1107 1835
rect 1227 1831 1231 1835
rect 1243 1831 1247 1835
rect 1403 1831 1407 1835
rect 1563 1831 1567 1835
rect 143 1822 147 1826
rect 287 1822 291 1826
rect 471 1822 475 1826
rect 663 1822 667 1826
rect 847 1822 851 1826
rect 1023 1822 1027 1826
rect 1191 1822 1195 1826
rect 1351 1822 1355 1826
rect 1511 1822 1515 1826
rect 1679 1822 1683 1826
rect 2335 1815 2339 1819
rect 2451 1815 2455 1819
rect 2459 1815 2463 1819
rect 2611 1815 2615 1819
rect 3039 1815 3043 1819
rect 3119 1815 3123 1819
rect 3203 1815 3204 1819
rect 3204 1815 3207 1819
rect 3227 1815 3231 1819
rect 3371 1815 3375 1819
rect 111 1804 115 1808
rect 1831 1804 1835 1808
rect 2095 1806 2099 1810
rect 2239 1806 2243 1810
rect 2399 1806 2403 1810
rect 2559 1806 2563 1810
rect 2719 1806 2723 1810
rect 2879 1806 2883 1810
rect 3031 1806 3035 1810
rect 3175 1806 3179 1810
rect 3319 1806 3323 1810
rect 3471 1806 3475 1810
rect 167 1795 171 1799
rect 295 1795 299 1799
rect 523 1795 527 1799
rect 715 1795 719 1799
rect 879 1795 883 1799
rect 1039 1795 1043 1799
rect 1243 1795 1247 1799
rect 1403 1795 1407 1799
rect 1563 1795 1567 1799
rect 111 1787 115 1791
rect 135 1784 139 1788
rect 279 1784 283 1788
rect 463 1784 467 1788
rect 655 1784 659 1788
rect 839 1784 843 1788
rect 1015 1784 1019 1788
rect 1183 1784 1187 1788
rect 1343 1784 1347 1788
rect 1503 1784 1507 1788
rect 1671 1784 1675 1788
rect 1831 1787 1835 1791
rect 1871 1788 1875 1792
rect 3591 1788 3595 1792
rect 2103 1779 2107 1783
rect 2335 1779 2339 1783
rect 2611 1779 2615 1783
rect 3039 1779 3043 1783
rect 3227 1779 3231 1783
rect 3371 1779 3375 1783
rect 1355 1767 1359 1771
rect 1871 1771 1875 1775
rect 2087 1768 2091 1772
rect 2231 1768 2235 1772
rect 2391 1768 2395 1772
rect 2551 1768 2555 1772
rect 2711 1768 2715 1772
rect 2871 1768 2875 1772
rect 3023 1768 3027 1772
rect 3167 1768 3171 1772
rect 3311 1768 3315 1772
rect 3463 1768 3467 1772
rect 3591 1771 3595 1775
rect 2699 1751 2703 1755
rect 2835 1751 2839 1755
rect 3427 1751 3431 1755
rect 111 1729 115 1733
rect 135 1732 139 1736
rect 215 1732 219 1736
rect 343 1732 347 1736
rect 495 1732 499 1736
rect 663 1732 667 1736
rect 839 1732 843 1736
rect 1007 1732 1011 1736
rect 1167 1732 1171 1736
rect 1319 1732 1323 1736
rect 1463 1732 1467 1736
rect 1607 1732 1611 1736
rect 1743 1732 1747 1736
rect 1831 1729 1835 1733
rect 203 1723 207 1727
rect 283 1723 287 1727
rect 487 1723 491 1727
rect 563 1723 567 1727
rect 731 1723 735 1727
rect 1091 1723 1095 1727
rect 1103 1723 1107 1727
rect 1411 1723 1415 1727
rect 1555 1723 1559 1727
rect 1691 1723 1695 1727
rect 1707 1723 1711 1727
rect 1871 1717 1875 1721
rect 2103 1720 2107 1724
rect 2239 1720 2243 1724
rect 2383 1720 2387 1724
rect 2527 1720 2531 1724
rect 2663 1720 2667 1724
rect 2799 1720 2803 1724
rect 2927 1720 2931 1724
rect 3047 1720 3051 1724
rect 3159 1720 3163 1724
rect 3271 1720 3275 1724
rect 3391 1720 3395 1724
rect 3503 1720 3507 1724
rect 111 1712 115 1716
rect 3591 1717 3595 1721
rect 1831 1712 1835 1716
rect 2187 1711 2191 1715
rect 2331 1711 2335 1715
rect 2451 1711 2455 1715
rect 2595 1711 2599 1715
rect 2899 1711 2903 1715
rect 3003 1711 3007 1715
rect 3119 1711 3123 1715
rect 3227 1711 3231 1715
rect 3459 1711 3463 1715
rect 1871 1700 1875 1704
rect 2655 1703 2659 1707
rect 3107 1703 3111 1707
rect 3563 1703 3567 1707
rect 3591 1700 3595 1704
rect 143 1694 147 1698
rect 223 1694 227 1698
rect 351 1694 355 1698
rect 503 1694 507 1698
rect 671 1694 675 1698
rect 847 1694 851 1698
rect 1015 1694 1019 1698
rect 1175 1694 1179 1698
rect 1327 1694 1331 1698
rect 1471 1694 1475 1698
rect 1615 1694 1619 1698
rect 1751 1694 1755 1698
rect 167 1683 168 1687
rect 168 1683 171 1687
rect 203 1683 207 1687
rect 283 1683 287 1687
rect 563 1683 567 1687
rect 731 1683 735 1687
rect 815 1683 819 1687
rect 1039 1683 1040 1687
rect 1040 1683 1043 1687
rect 1091 1683 1095 1687
rect 1355 1683 1356 1687
rect 1356 1683 1359 1687
rect 1411 1683 1415 1687
rect 1555 1683 1559 1687
rect 1691 1683 1695 1687
rect 2111 1682 2115 1686
rect 2247 1682 2251 1686
rect 2391 1682 2395 1686
rect 2535 1682 2539 1686
rect 2671 1682 2675 1686
rect 2807 1682 2811 1686
rect 2935 1682 2939 1686
rect 3055 1682 3059 1686
rect 3167 1682 3171 1686
rect 3279 1682 3283 1686
rect 3399 1682 3403 1686
rect 3511 1682 3515 1686
rect 303 1667 307 1671
rect 863 1675 867 1679
rect 531 1667 535 1671
rect 915 1667 919 1671
rect 1059 1667 1060 1671
rect 1060 1667 1063 1671
rect 1367 1667 1371 1671
rect 1527 1667 1531 1671
rect 1687 1667 1691 1671
rect 1707 1667 1708 1671
rect 1708 1667 1711 1671
rect 2187 1671 2191 1675
rect 2331 1671 2335 1675
rect 2595 1671 2599 1675
rect 2699 1671 2700 1675
rect 2700 1671 2703 1675
rect 2835 1671 2836 1675
rect 2836 1671 2839 1675
rect 2899 1671 2903 1675
rect 3003 1671 3007 1675
rect 3227 1671 3231 1675
rect 3383 1671 3387 1675
rect 3427 1671 3428 1675
rect 3428 1671 3431 1675
rect 3459 1671 3463 1675
rect 2359 1663 2363 1667
rect 143 1658 147 1662
rect 295 1658 299 1662
rect 479 1658 483 1662
rect 671 1658 675 1662
rect 855 1658 859 1662
rect 1031 1658 1035 1662
rect 1199 1658 1203 1662
rect 1359 1658 1363 1662
rect 1519 1658 1523 1662
rect 1679 1658 1683 1662
rect 1975 1655 1979 1659
rect 2019 1655 2023 1659
rect 2139 1655 2143 1659
rect 2267 1655 2271 1659
rect 2647 1655 2651 1659
rect 2655 1655 2659 1659
rect 3079 1655 3083 1659
rect 3107 1655 3111 1659
rect 3179 1655 3183 1659
rect 3331 1655 3335 1659
rect 3563 1655 3567 1659
rect 1967 1646 1971 1650
rect 2087 1646 2091 1650
rect 2215 1646 2219 1650
rect 2351 1646 2355 1650
rect 2495 1646 2499 1650
rect 2639 1646 2643 1650
rect 2783 1646 2787 1650
rect 2927 1646 2931 1650
rect 3071 1646 3075 1650
rect 3223 1646 3227 1650
rect 3375 1646 3379 1650
rect 3511 1646 3515 1650
rect 111 1640 115 1644
rect 1831 1640 1835 1644
rect 191 1631 195 1635
rect 303 1631 307 1635
rect 531 1631 535 1635
rect 815 1631 819 1635
rect 863 1631 867 1635
rect 1039 1631 1043 1635
rect 1263 1631 1267 1635
rect 1367 1631 1371 1635
rect 1527 1631 1531 1635
rect 1687 1631 1691 1635
rect 1871 1628 1875 1632
rect 111 1623 115 1627
rect 3591 1628 3595 1632
rect 135 1620 139 1624
rect 287 1620 291 1624
rect 471 1620 475 1624
rect 663 1620 667 1624
rect 847 1620 851 1624
rect 1023 1620 1027 1624
rect 1191 1620 1195 1624
rect 1351 1620 1355 1624
rect 1511 1620 1515 1624
rect 1671 1620 1675 1624
rect 1831 1623 1835 1627
rect 2019 1619 2023 1623
rect 2139 1619 2143 1623
rect 2267 1619 2271 1623
rect 2359 1619 2363 1623
rect 2547 1619 2551 1623
rect 2647 1619 2651 1623
rect 3079 1619 3083 1623
rect 3331 1619 3335 1623
rect 3383 1619 3387 1623
rect 3535 1619 3539 1623
rect 1871 1611 1875 1615
rect 1959 1608 1963 1612
rect 2079 1608 2083 1612
rect 2207 1608 2211 1612
rect 2343 1608 2347 1612
rect 2487 1608 2491 1612
rect 2631 1608 2635 1612
rect 2775 1608 2779 1612
rect 2919 1608 2923 1612
rect 3063 1608 3067 1612
rect 3215 1608 3219 1612
rect 3367 1608 3371 1612
rect 3503 1608 3507 1612
rect 3591 1611 3595 1615
rect 2723 1591 2727 1595
rect 111 1573 115 1577
rect 159 1576 163 1580
rect 287 1576 291 1580
rect 423 1576 427 1580
rect 567 1576 571 1580
rect 711 1576 715 1580
rect 847 1576 851 1580
rect 983 1576 987 1580
rect 1119 1576 1123 1580
rect 1247 1576 1251 1580
rect 1375 1576 1379 1580
rect 1511 1576 1515 1580
rect 1831 1573 1835 1577
rect 231 1567 235 1571
rect 259 1567 263 1571
rect 535 1567 539 1571
rect 659 1567 663 1571
rect 803 1567 807 1571
rect 915 1567 919 1571
rect 1051 1567 1055 1571
rect 1059 1567 1063 1571
rect 1331 1567 1335 1571
rect 1443 1567 1447 1571
rect 1451 1567 1455 1571
rect 111 1556 115 1560
rect 1831 1556 1835 1560
rect 1871 1553 1875 1557
rect 1895 1556 1899 1560
rect 2047 1556 2051 1560
rect 2207 1556 2211 1560
rect 2367 1556 2371 1560
rect 2527 1556 2531 1560
rect 2687 1556 2691 1560
rect 2839 1556 2843 1560
rect 2983 1556 2987 1560
rect 3119 1556 3123 1560
rect 3255 1556 3259 1560
rect 3391 1556 3395 1560
rect 3503 1556 3507 1560
rect 3591 1553 3595 1557
rect 167 1538 171 1542
rect 295 1538 299 1542
rect 431 1538 435 1542
rect 575 1538 579 1542
rect 719 1538 723 1542
rect 855 1538 859 1542
rect 991 1538 995 1542
rect 1127 1538 1131 1542
rect 1255 1538 1259 1542
rect 1383 1538 1387 1542
rect 1519 1538 1523 1542
rect 1963 1547 1967 1551
rect 2115 1547 2119 1551
rect 1871 1536 1875 1540
rect 1975 1539 1979 1543
rect 2435 1547 2439 1551
rect 2755 1547 2759 1551
rect 2931 1547 2935 1551
rect 3055 1547 3059 1551
rect 3187 1547 3191 1551
rect 3323 1547 3327 1551
rect 2443 1539 2447 1543
rect 3179 1539 3183 1543
rect 3563 1539 3567 1543
rect 3591 1536 3595 1540
rect 191 1527 192 1531
rect 192 1527 195 1531
rect 231 1527 235 1531
rect 527 1527 531 1531
rect 535 1527 539 1531
rect 659 1527 663 1531
rect 803 1527 807 1531
rect 1015 1527 1016 1531
rect 1016 1527 1019 1531
rect 1051 1527 1055 1531
rect 1263 1527 1267 1531
rect 1331 1527 1335 1531
rect 1443 1527 1447 1531
rect 259 1511 260 1515
rect 260 1511 263 1515
rect 283 1511 287 1515
rect 791 1519 795 1523
rect 1903 1518 1907 1522
rect 2055 1518 2059 1522
rect 2215 1518 2219 1522
rect 2375 1518 2379 1522
rect 2535 1518 2539 1522
rect 2695 1518 2699 1522
rect 2847 1518 2851 1522
rect 2991 1518 2995 1522
rect 3127 1518 3131 1522
rect 3263 1518 3267 1522
rect 3399 1518 3403 1522
rect 3511 1518 3515 1522
rect 699 1511 703 1515
rect 707 1511 711 1515
rect 927 1511 928 1515
rect 928 1511 931 1515
rect 955 1511 959 1515
rect 1155 1511 1159 1515
rect 1171 1511 1175 1515
rect 1267 1511 1271 1515
rect 1451 1511 1452 1515
rect 1452 1511 1455 1515
rect 231 1502 235 1506
rect 375 1502 379 1506
rect 519 1502 523 1506
rect 655 1502 659 1506
rect 783 1502 787 1506
rect 903 1502 907 1506
rect 1015 1502 1019 1506
rect 1119 1502 1123 1506
rect 1215 1502 1219 1506
rect 1319 1502 1323 1506
rect 1963 1507 1967 1511
rect 2115 1507 2119 1511
rect 2187 1507 2191 1511
rect 2435 1507 2439 1511
rect 2547 1507 2551 1511
rect 2723 1507 2724 1511
rect 2724 1507 2727 1511
rect 2755 1507 2759 1511
rect 2931 1507 2935 1511
rect 3187 1507 3191 1511
rect 3323 1507 3327 1511
rect 3419 1507 3423 1511
rect 3535 1507 3536 1511
rect 3536 1507 3539 1511
rect 1423 1502 1427 1506
rect 111 1484 115 1488
rect 1831 1484 1835 1488
rect 1963 1487 1967 1491
rect 1971 1487 1975 1491
rect 2127 1487 2131 1491
rect 2423 1487 2427 1491
rect 2443 1487 2444 1491
rect 2444 1487 2447 1491
rect 2727 1487 2731 1491
rect 2887 1487 2891 1491
rect 3047 1487 3051 1491
rect 3055 1487 3059 1491
rect 3519 1495 3523 1499
rect 3251 1487 3255 1491
rect 3563 1487 3567 1491
rect 283 1475 287 1479
rect 427 1475 431 1479
rect 527 1475 531 1479
rect 707 1475 711 1479
rect 791 1475 795 1479
rect 955 1475 959 1479
rect 1023 1475 1027 1479
rect 1171 1475 1175 1479
rect 1267 1475 1271 1479
rect 1371 1475 1375 1479
rect 1431 1475 1435 1479
rect 1903 1478 1907 1482
rect 2007 1478 2011 1482
rect 2135 1478 2139 1482
rect 2271 1478 2275 1482
rect 2415 1478 2419 1482
rect 2567 1478 2571 1482
rect 2719 1478 2723 1482
rect 2879 1478 2883 1482
rect 3039 1478 3043 1482
rect 3199 1478 3203 1482
rect 3367 1478 3371 1482
rect 3511 1478 3515 1482
rect 111 1467 115 1471
rect 223 1464 227 1468
rect 367 1464 371 1468
rect 511 1464 515 1468
rect 647 1464 651 1468
rect 775 1464 779 1468
rect 895 1464 899 1468
rect 1007 1464 1011 1468
rect 1111 1464 1115 1468
rect 1207 1464 1211 1468
rect 1311 1464 1315 1468
rect 1415 1464 1419 1468
rect 1831 1467 1835 1471
rect 1871 1460 1875 1464
rect 3591 1460 3595 1464
rect 1971 1451 1975 1455
rect 2127 1451 2131 1455
rect 2187 1451 2191 1455
rect 2423 1451 2427 1455
rect 2727 1451 2731 1455
rect 2887 1451 2891 1455
rect 3047 1451 3051 1455
rect 3251 1451 3255 1455
rect 3419 1451 3423 1455
rect 3519 1451 3523 1455
rect 1871 1443 1875 1447
rect 1895 1440 1899 1444
rect 1999 1440 2003 1444
rect 2127 1440 2131 1444
rect 2263 1440 2267 1444
rect 2407 1440 2411 1444
rect 2559 1440 2563 1444
rect 2711 1440 2715 1444
rect 2871 1440 2875 1444
rect 3031 1440 3035 1444
rect 3191 1440 3195 1444
rect 3359 1440 3363 1444
rect 3503 1440 3507 1444
rect 3591 1443 3595 1447
rect 2059 1423 2063 1427
rect 2467 1423 2471 1427
rect 111 1409 115 1413
rect 255 1412 259 1416
rect 351 1412 355 1416
rect 447 1412 451 1416
rect 543 1412 547 1416
rect 631 1412 635 1416
rect 719 1412 723 1416
rect 807 1412 811 1416
rect 919 1412 923 1416
rect 1047 1412 1051 1416
rect 1207 1412 1211 1416
rect 1383 1412 1387 1416
rect 1575 1412 1579 1416
rect 1743 1412 1747 1416
rect 1831 1409 1835 1413
rect 343 1403 347 1407
rect 419 1403 423 1407
rect 611 1403 615 1407
rect 699 1403 703 1407
rect 111 1392 115 1396
rect 315 1395 319 1399
rect 603 1395 607 1399
rect 787 1403 791 1407
rect 927 1399 931 1403
rect 987 1403 991 1407
rect 1115 1403 1119 1407
rect 1503 1403 1507 1407
rect 1519 1403 1523 1407
rect 1811 1403 1815 1407
rect 1831 1392 1835 1396
rect 1871 1393 1875 1397
rect 1895 1396 1899 1400
rect 2023 1396 2027 1400
rect 2167 1396 2171 1400
rect 2303 1396 2307 1400
rect 2431 1396 2435 1400
rect 2551 1396 2555 1400
rect 2671 1396 2675 1400
rect 2791 1396 2795 1400
rect 2911 1396 2915 1400
rect 3591 1393 3595 1397
rect 871 1383 875 1387
rect 987 1383 991 1387
rect 1963 1387 1967 1391
rect 2115 1387 2119 1391
rect 2259 1387 2263 1391
rect 2379 1387 2383 1391
rect 2515 1387 2519 1391
rect 2635 1387 2639 1391
rect 2755 1387 2759 1391
rect 2867 1387 2871 1391
rect 2875 1387 2879 1391
rect 263 1374 267 1378
rect 359 1374 363 1378
rect 455 1374 459 1378
rect 551 1374 555 1378
rect 639 1374 643 1378
rect 727 1374 731 1378
rect 815 1374 819 1378
rect 927 1374 931 1378
rect 1055 1374 1059 1378
rect 1215 1374 1219 1378
rect 1391 1374 1395 1378
rect 1583 1374 1587 1378
rect 1751 1374 1755 1378
rect 1871 1376 1875 1380
rect 3591 1376 3595 1380
rect 343 1363 347 1367
rect 419 1363 423 1367
rect 427 1363 431 1367
rect 603 1363 607 1367
rect 611 1363 615 1367
rect 787 1363 791 1367
rect 871 1363 875 1367
rect 915 1363 919 1367
rect 1115 1363 1119 1367
rect 1243 1363 1244 1367
rect 1244 1363 1247 1367
rect 1371 1363 1375 1367
rect 1503 1363 1507 1367
rect 1775 1363 1776 1367
rect 1776 1363 1779 1367
rect 1903 1358 1907 1362
rect 2031 1358 2035 1362
rect 2175 1358 2179 1362
rect 2311 1358 2315 1362
rect 2439 1358 2443 1362
rect 2559 1358 2563 1362
rect 2679 1358 2683 1362
rect 2799 1358 2803 1362
rect 2919 1358 2923 1362
rect 315 1351 319 1355
rect 411 1351 415 1355
rect 523 1351 527 1355
rect 719 1351 723 1355
rect 1015 1351 1019 1355
rect 1151 1351 1155 1355
rect 1171 1351 1172 1355
rect 1172 1351 1175 1355
rect 1307 1351 1308 1355
rect 1308 1351 1311 1355
rect 1331 1351 1335 1355
rect 1459 1351 1463 1355
rect 1699 1351 1703 1355
rect 1811 1347 1815 1351
rect 359 1342 363 1346
rect 471 1342 475 1346
rect 591 1342 595 1346
rect 727 1342 731 1346
rect 863 1342 867 1346
rect 1007 1342 1011 1346
rect 1143 1342 1147 1346
rect 1279 1342 1283 1346
rect 1407 1342 1411 1346
rect 1527 1342 1531 1346
rect 1647 1342 1651 1346
rect 2059 1347 2060 1351
rect 2060 1347 2063 1351
rect 2115 1347 2119 1351
rect 2259 1347 2263 1351
rect 2467 1347 2468 1351
rect 2468 1347 2471 1351
rect 2515 1347 2519 1351
rect 2635 1347 2639 1351
rect 2755 1347 2759 1351
rect 2867 1347 2871 1351
rect 1751 1342 1755 1346
rect 2379 1335 2383 1339
rect 111 1324 115 1328
rect 1831 1324 1835 1328
rect 411 1315 415 1319
rect 523 1315 527 1319
rect 719 1315 723 1319
rect 915 1315 919 1319
rect 1015 1315 1019 1319
rect 1151 1315 1155 1319
rect 1331 1315 1335 1319
rect 1459 1315 1463 1319
rect 1699 1315 1703 1319
rect 1775 1315 1779 1319
rect 1927 1318 1931 1322
rect 1979 1327 1983 1331
rect 2099 1327 2103 1331
rect 2463 1327 2467 1331
rect 2619 1327 2620 1331
rect 2620 1327 2623 1331
rect 2643 1327 2647 1331
rect 2771 1327 2775 1331
rect 2891 1327 2895 1331
rect 3003 1327 3007 1331
rect 3115 1327 3119 1331
rect 1987 1319 1991 1323
rect 2047 1318 2051 1322
rect 2183 1318 2187 1322
rect 2319 1318 2323 1322
rect 2455 1318 2459 1322
rect 2591 1318 2595 1322
rect 2719 1318 2723 1322
rect 2839 1318 2843 1322
rect 2951 1318 2955 1322
rect 3063 1318 3067 1322
rect 3183 1318 3187 1322
rect 111 1307 115 1311
rect 351 1304 355 1308
rect 463 1304 467 1308
rect 583 1304 587 1308
rect 719 1304 723 1308
rect 855 1304 859 1308
rect 999 1304 1003 1308
rect 1135 1304 1139 1308
rect 1271 1304 1275 1308
rect 1399 1304 1403 1308
rect 1519 1304 1523 1308
rect 1639 1304 1643 1308
rect 1743 1304 1747 1308
rect 1831 1307 1835 1311
rect 1871 1300 1875 1304
rect 3591 1300 3595 1304
rect 707 1287 711 1291
rect 1979 1291 1983 1295
rect 2099 1291 2103 1295
rect 2235 1291 2239 1295
rect 2327 1291 2331 1295
rect 2463 1291 2467 1295
rect 2643 1291 2647 1295
rect 2771 1291 2775 1295
rect 2891 1291 2895 1295
rect 3003 1291 3007 1295
rect 3115 1291 3119 1295
rect 1871 1283 1875 1287
rect 1919 1280 1923 1284
rect 2039 1280 2043 1284
rect 2175 1280 2179 1284
rect 2311 1280 2315 1284
rect 2447 1280 2451 1284
rect 2583 1280 2587 1284
rect 2711 1280 2715 1284
rect 2831 1280 2835 1284
rect 2943 1280 2947 1284
rect 3055 1280 3059 1284
rect 3175 1280 3179 1284
rect 3591 1283 3595 1287
rect 3063 1263 3067 1267
rect 111 1253 115 1257
rect 311 1256 315 1260
rect 415 1256 419 1260
rect 535 1256 539 1260
rect 671 1256 675 1260
rect 815 1256 819 1260
rect 959 1256 963 1260
rect 1103 1256 1107 1260
rect 1239 1256 1243 1260
rect 1375 1256 1379 1260
rect 1503 1256 1507 1260
rect 1631 1256 1635 1260
rect 1743 1256 1747 1260
rect 1831 1253 1835 1257
rect 267 1247 271 1251
rect 379 1247 383 1251
rect 483 1247 487 1251
rect 603 1247 607 1251
rect 907 1247 911 1251
rect 1051 1247 1055 1251
rect 1171 1247 1175 1251
rect 1331 1247 1335 1251
rect 1463 1247 1467 1251
rect 1591 1247 1595 1251
rect 1599 1247 1603 1251
rect 111 1236 115 1240
rect 1803 1239 1807 1243
rect 1831 1236 1835 1240
rect 1871 1225 1875 1229
rect 1895 1228 1899 1232
rect 2071 1228 2075 1232
rect 2271 1228 2275 1232
rect 2471 1228 2475 1232
rect 2663 1228 2667 1232
rect 2847 1228 2851 1232
rect 3023 1228 3027 1232
rect 3191 1228 3195 1232
rect 3359 1228 3363 1232
rect 3503 1228 3507 1232
rect 3591 1225 3595 1229
rect 319 1218 323 1222
rect 423 1218 427 1222
rect 543 1218 547 1222
rect 679 1218 683 1222
rect 823 1218 827 1222
rect 967 1218 971 1222
rect 1111 1218 1115 1222
rect 1247 1218 1251 1222
rect 1383 1218 1387 1222
rect 1511 1218 1515 1222
rect 1639 1218 1643 1222
rect 1751 1218 1755 1222
rect 379 1207 383 1211
rect 483 1207 487 1211
rect 603 1207 607 1211
rect 707 1207 708 1211
rect 708 1207 711 1211
rect 811 1207 815 1211
rect 907 1207 911 1211
rect 1051 1207 1055 1211
rect 1331 1207 1335 1211
rect 1463 1207 1467 1211
rect 1591 1207 1595 1211
rect 1871 1208 1875 1212
rect 1955 1211 1959 1215
rect 2139 1219 2143 1223
rect 2591 1219 2595 1223
rect 2779 1219 2783 1223
rect 2915 1219 2919 1223
rect 3263 1219 3267 1223
rect 3451 1219 3455 1223
rect 2723 1211 2727 1215
rect 3563 1211 3567 1215
rect 3591 1208 3595 1212
rect 267 1195 268 1199
rect 268 1195 271 1199
rect 291 1195 295 1199
rect 467 1195 471 1199
rect 935 1195 939 1199
rect 943 1195 947 1199
rect 1123 1195 1127 1199
rect 1131 1195 1135 1199
rect 1275 1195 1279 1199
rect 1419 1195 1423 1199
rect 1555 1195 1559 1199
rect 1803 1195 1807 1199
rect 239 1186 243 1190
rect 415 1186 419 1190
rect 591 1186 595 1190
rect 759 1186 763 1190
rect 927 1186 931 1190
rect 1079 1186 1083 1190
rect 1223 1186 1227 1190
rect 1367 1186 1371 1190
rect 1503 1186 1507 1190
rect 1639 1186 1643 1190
rect 1751 1186 1755 1190
rect 1903 1190 1907 1194
rect 2079 1190 2083 1194
rect 2279 1190 2283 1194
rect 2479 1190 2483 1194
rect 2671 1190 2675 1194
rect 2855 1190 2859 1194
rect 3031 1190 3035 1194
rect 3199 1190 3203 1194
rect 3367 1190 3371 1194
rect 3511 1190 3515 1194
rect 1803 1179 1807 1183
rect 2139 1179 2143 1183
rect 2235 1179 2239 1183
rect 2507 1179 2508 1183
rect 2508 1179 2511 1183
rect 2591 1179 2595 1183
rect 2915 1179 2919 1183
rect 3056 1179 3060 1183
rect 3263 1179 3267 1183
rect 3451 1179 3455 1183
rect 111 1168 115 1172
rect 1831 1168 1835 1172
rect 3407 1171 3411 1175
rect 291 1159 295 1163
rect 467 1159 471 1163
rect 811 1159 815 1163
rect 935 1159 939 1163
rect 1131 1159 1135 1163
rect 1275 1159 1279 1163
rect 1419 1159 1423 1163
rect 1555 1159 1559 1163
rect 1803 1159 1807 1163
rect 1955 1163 1959 1167
rect 1963 1163 1967 1167
rect 2035 1163 2039 1167
rect 2139 1163 2143 1167
rect 2267 1163 2271 1167
rect 2419 1163 2423 1167
rect 2723 1163 2727 1167
rect 2739 1163 2743 1167
rect 3011 1163 3012 1167
rect 3012 1163 3015 1167
rect 3179 1163 3183 1167
rect 3315 1163 3319 1167
rect 3563 1163 3567 1167
rect 111 1151 115 1155
rect 231 1148 235 1152
rect 407 1148 411 1152
rect 583 1148 587 1152
rect 751 1148 755 1152
rect 919 1148 923 1152
rect 1071 1148 1075 1152
rect 1215 1148 1219 1152
rect 1359 1148 1363 1152
rect 1495 1148 1499 1152
rect 1631 1148 1635 1152
rect 1743 1148 1747 1152
rect 1831 1151 1835 1155
rect 1903 1154 1907 1158
rect 1983 1154 1987 1158
rect 2087 1154 2091 1158
rect 2215 1154 2219 1158
rect 2367 1154 2371 1158
rect 2527 1154 2531 1158
rect 2687 1154 2691 1158
rect 2839 1154 2843 1158
rect 2983 1154 2987 1158
rect 3127 1154 3131 1158
rect 3263 1154 3267 1158
rect 3399 1154 3403 1158
rect 3511 1154 3515 1158
rect 1871 1136 1875 1140
rect 459 1131 463 1135
rect 3591 1136 3595 1140
rect 1123 1123 1127 1127
rect 1439 1123 1443 1127
rect 1963 1127 1967 1131
rect 2035 1127 2039 1131
rect 2139 1127 2143 1131
rect 2267 1127 2271 1131
rect 2419 1127 2423 1131
rect 2739 1127 2743 1131
rect 2919 1127 2923 1131
rect 3179 1127 3183 1131
rect 3315 1127 3319 1131
rect 3407 1127 3411 1131
rect 3535 1127 3539 1131
rect 1871 1119 1875 1123
rect 1895 1116 1899 1120
rect 1975 1116 1979 1120
rect 2079 1116 2083 1120
rect 2207 1116 2211 1120
rect 2359 1116 2363 1120
rect 2519 1116 2523 1120
rect 2679 1116 2683 1120
rect 2831 1116 2835 1120
rect 2975 1116 2979 1120
rect 3119 1116 3123 1120
rect 3255 1116 3259 1120
rect 3391 1116 3395 1120
rect 3503 1116 3507 1120
rect 3591 1119 3595 1123
rect 111 1097 115 1101
rect 143 1100 147 1104
rect 279 1100 283 1104
rect 423 1100 427 1104
rect 567 1100 571 1104
rect 711 1100 715 1104
rect 847 1100 851 1104
rect 975 1100 979 1104
rect 1103 1100 1107 1104
rect 1223 1100 1227 1104
rect 1343 1100 1347 1104
rect 1471 1100 1475 1104
rect 1831 1097 1835 1101
rect 2215 1099 2219 1103
rect 211 1091 215 1095
rect 347 1091 351 1095
rect 635 1091 639 1095
rect 803 1091 807 1095
rect 943 1091 947 1095
rect 1063 1091 1067 1095
rect 1187 1091 1191 1095
rect 1307 1091 1311 1095
rect 1431 1091 1435 1095
rect 1439 1091 1443 1095
rect 111 1080 115 1084
rect 203 1083 207 1087
rect 1831 1080 1835 1084
rect 151 1062 155 1066
rect 287 1062 291 1066
rect 431 1062 435 1066
rect 575 1062 579 1066
rect 719 1062 723 1066
rect 855 1062 859 1066
rect 983 1062 987 1066
rect 1111 1062 1115 1066
rect 1231 1062 1235 1066
rect 1351 1062 1355 1066
rect 1479 1062 1483 1066
rect 1871 1061 1875 1065
rect 2167 1064 2171 1068
rect 2255 1064 2259 1068
rect 2359 1064 2363 1068
rect 2479 1064 2483 1068
rect 2607 1064 2611 1068
rect 2751 1064 2755 1068
rect 2895 1064 2899 1068
rect 3047 1064 3051 1068
rect 3207 1064 3211 1068
rect 3367 1064 3371 1068
rect 3503 1064 3507 1068
rect 3591 1061 3595 1065
rect 211 1051 215 1055
rect 347 1051 351 1055
rect 459 1051 460 1055
rect 460 1051 463 1055
rect 599 1051 600 1055
rect 600 1051 603 1055
rect 635 1051 639 1055
rect 803 1051 807 1055
rect 1055 1051 1059 1055
rect 1063 1051 1067 1055
rect 1187 1051 1191 1055
rect 1307 1051 1311 1055
rect 1431 1051 1435 1055
rect 2235 1055 2239 1059
rect 2331 1055 2335 1059
rect 2435 1055 2439 1059
rect 2555 1055 2559 1059
rect 2563 1055 2567 1059
rect 2819 1055 2823 1059
rect 3011 1055 3015 1059
rect 3115 1055 3119 1059
rect 3275 1055 3279 1059
rect 1871 1044 1875 1048
rect 2811 1047 2815 1051
rect 3563 1047 3567 1051
rect 3591 1044 3595 1048
rect 415 1039 419 1043
rect 203 1031 207 1035
rect 315 1031 319 1035
rect 695 1031 699 1035
rect 755 1031 759 1035
rect 919 1031 923 1035
rect 1031 1031 1035 1035
rect 1091 1031 1095 1035
rect 1195 1031 1199 1035
rect 1299 1031 1303 1035
rect 143 1022 147 1026
rect 263 1022 267 1026
rect 407 1022 411 1026
rect 551 1022 555 1026
rect 687 1022 691 1026
rect 807 1022 811 1026
rect 927 1022 931 1026
rect 1039 1022 1043 1026
rect 1143 1022 1147 1026
rect 1247 1022 1251 1026
rect 1359 1022 1363 1026
rect 2175 1026 2179 1030
rect 2263 1026 2267 1030
rect 2367 1026 2371 1030
rect 2487 1026 2491 1030
rect 2615 1026 2619 1030
rect 2759 1026 2763 1030
rect 2903 1026 2907 1030
rect 3055 1026 3059 1030
rect 3215 1026 3219 1030
rect 3375 1026 3379 1030
rect 3511 1026 3515 1030
rect 2215 1015 2219 1019
rect 2235 1015 2239 1019
rect 2331 1015 2335 1019
rect 2435 1015 2439 1019
rect 2555 1015 2559 1019
rect 2819 1015 2823 1019
rect 2919 1015 2923 1019
rect 3115 1015 3119 1019
rect 3275 1015 3279 1019
rect 3399 1015 3400 1019
rect 3400 1015 3403 1019
rect 3535 1015 3536 1019
rect 3536 1015 3539 1019
rect 111 1004 115 1008
rect 1831 1004 1835 1008
rect 2347 1003 2351 1007
rect 2355 1003 2359 1007
rect 2435 1003 2439 1007
rect 2523 1003 2527 1007
rect 2811 1003 2812 1007
rect 2812 1003 2815 1007
rect 2835 1003 2839 1007
rect 3075 1003 3079 1007
rect 3107 1003 3111 1007
rect 3259 1003 3263 1007
rect 3563 1003 3567 1007
rect 167 995 171 999
rect 315 995 319 999
rect 415 995 419 999
rect 599 995 603 999
rect 695 995 699 999
rect 919 995 923 999
rect 1031 995 1035 999
rect 1091 995 1095 999
rect 1195 995 1199 999
rect 1299 995 1303 999
rect 1367 995 1371 999
rect 2303 994 2307 998
rect 2383 994 2387 998
rect 2471 994 2475 998
rect 2567 994 2571 998
rect 2671 994 2675 998
rect 2783 994 2787 998
rect 2911 994 2915 998
rect 3055 994 3059 998
rect 3207 994 3211 998
rect 3367 994 3371 998
rect 3511 994 3515 998
rect 111 987 115 991
rect 135 984 139 988
rect 255 984 259 988
rect 399 984 403 988
rect 543 984 547 988
rect 679 984 683 988
rect 799 984 803 988
rect 919 984 923 988
rect 1031 984 1035 988
rect 1135 984 1139 988
rect 1239 984 1243 988
rect 1351 984 1355 988
rect 1831 987 1835 991
rect 1871 976 1875 980
rect 3591 976 3595 980
rect 2355 967 2359 971
rect 2435 967 2439 971
rect 2523 967 2527 971
rect 2723 967 2727 971
rect 2835 967 2839 971
rect 3107 967 3111 971
rect 3259 967 3263 971
rect 3399 967 3403 971
rect 3535 967 3539 971
rect 1871 959 1875 963
rect 2295 956 2299 960
rect 2375 956 2379 960
rect 2463 956 2467 960
rect 2559 956 2563 960
rect 2663 956 2667 960
rect 2775 956 2779 960
rect 2903 956 2907 960
rect 3047 956 3051 960
rect 3199 956 3203 960
rect 3359 956 3363 960
rect 3503 956 3507 960
rect 3591 959 3595 963
rect 2843 939 2847 943
rect 111 929 115 933
rect 135 932 139 936
rect 215 932 219 936
rect 327 932 331 936
rect 447 932 451 936
rect 567 932 571 936
rect 687 932 691 936
rect 799 932 803 936
rect 911 932 915 936
rect 1015 932 1019 936
rect 1119 932 1123 936
rect 1223 932 1227 936
rect 1327 932 1331 936
rect 1831 929 1835 933
rect 203 923 207 927
rect 283 923 287 927
rect 399 923 403 927
rect 427 923 431 927
rect 651 923 655 927
rect 755 923 759 927
rect 867 923 871 927
rect 979 923 983 927
rect 1083 923 1087 927
rect 1299 923 1303 927
rect 111 912 115 916
rect 1195 915 1199 919
rect 1831 912 1835 916
rect 1871 901 1875 905
rect 2279 904 2283 908
rect 2359 904 2363 908
rect 2439 904 2443 908
rect 2519 904 2523 908
rect 2607 904 2611 908
rect 2703 904 2707 908
rect 2807 904 2811 908
rect 2911 904 2915 908
rect 3015 904 3019 908
rect 3111 904 3115 908
rect 3215 904 3219 908
rect 3319 904 3323 908
rect 3423 904 3427 908
rect 3503 904 3507 908
rect 3591 901 3595 905
rect 143 894 147 898
rect 223 894 227 898
rect 335 894 339 898
rect 455 894 459 898
rect 575 894 579 898
rect 695 894 699 898
rect 807 894 811 898
rect 919 894 923 898
rect 1023 894 1027 898
rect 1127 894 1131 898
rect 1231 894 1235 898
rect 1335 894 1339 898
rect 2347 895 2351 899
rect 2431 895 2435 899
rect 167 883 168 887
rect 168 883 171 887
rect 203 883 207 887
rect 283 883 287 887
rect 399 883 403 887
rect 599 883 600 887
rect 600 883 603 887
rect 651 883 655 887
rect 867 883 871 887
rect 979 883 983 887
rect 1083 883 1087 887
rect 1195 883 1199 887
rect 1203 883 1207 887
rect 1299 883 1303 887
rect 1871 884 1875 888
rect 2339 887 2343 891
rect 2507 895 2511 899
rect 2587 895 2591 899
rect 2675 895 2679 899
rect 2891 895 2895 899
rect 2919 891 2923 895
rect 3083 895 3087 899
rect 3179 895 3183 899
rect 3283 895 3287 899
rect 3491 895 3495 899
rect 3075 887 3079 891
rect 3483 887 3487 891
rect 3591 884 3595 888
rect 1287 871 1291 875
rect 263 863 267 867
rect 407 863 411 867
rect 427 863 428 867
rect 428 863 431 867
rect 727 863 731 867
rect 879 863 883 867
rect 887 863 891 867
rect 1107 859 1111 863
rect 1407 863 1411 867
rect 1527 863 1531 867
rect 1655 863 1659 867
rect 1711 863 1715 867
rect 2287 866 2291 870
rect 2367 866 2371 870
rect 2447 866 2451 870
rect 2527 866 2531 870
rect 2615 866 2619 870
rect 2711 866 2715 870
rect 2815 866 2819 870
rect 2919 866 2923 870
rect 3023 866 3027 870
rect 3119 866 3123 870
rect 3223 866 3227 870
rect 3327 866 3331 870
rect 3431 866 3435 870
rect 3511 866 3515 870
rect 143 854 147 858
rect 255 854 259 858
rect 399 854 403 858
rect 559 854 563 858
rect 719 854 723 858
rect 871 854 875 858
rect 1015 854 1019 858
rect 1151 854 1155 858
rect 1279 854 1283 858
rect 1399 854 1403 858
rect 1519 854 1523 858
rect 1647 854 1651 858
rect 2339 855 2343 859
rect 2347 855 2351 859
rect 2507 855 2511 859
rect 2587 855 2591 859
rect 2675 855 2679 859
rect 2723 855 2727 859
rect 2843 855 2844 859
rect 2844 855 2847 859
rect 2891 855 2895 859
rect 3083 855 3087 859
rect 3179 855 3183 859
rect 3283 855 3287 859
rect 3415 855 3419 859
rect 3491 855 3495 859
rect 3535 855 3536 859
rect 3536 855 3539 859
rect 111 836 115 840
rect 1831 836 1835 840
rect 167 827 171 831
rect 263 827 267 831
rect 407 827 411 831
rect 599 827 603 831
rect 727 827 731 831
rect 879 827 883 831
rect 1107 827 1111 831
rect 1203 827 1207 831
rect 1287 827 1291 831
rect 1407 827 1411 831
rect 1527 827 1531 831
rect 1655 827 1659 831
rect 2335 839 2339 843
rect 2219 831 2223 835
rect 2663 839 2667 843
rect 2431 831 2435 835
rect 2475 831 2479 835
rect 2587 831 2591 835
rect 2859 831 2863 835
rect 2927 831 2931 835
rect 3055 831 3059 835
rect 3091 831 3095 835
rect 3211 831 3215 835
rect 3395 831 3399 835
rect 3483 831 3487 835
rect 111 819 115 823
rect 135 816 139 820
rect 247 816 251 820
rect 391 816 395 820
rect 551 816 555 820
rect 711 816 715 820
rect 863 816 867 820
rect 1007 816 1011 820
rect 1143 816 1147 820
rect 1271 816 1275 820
rect 1391 816 1395 820
rect 1511 816 1515 820
rect 1639 816 1643 820
rect 1831 819 1835 823
rect 2167 822 2171 826
rect 2247 822 2251 826
rect 2327 822 2331 826
rect 2423 822 2427 826
rect 2535 822 2539 826
rect 2655 822 2659 826
rect 2783 822 2787 826
rect 2911 822 2915 826
rect 3039 822 3043 826
rect 3159 822 3163 826
rect 3279 822 3283 826
rect 3407 822 3411 826
rect 3511 822 3515 826
rect 1871 804 1875 808
rect 3591 804 3595 808
rect 2219 795 2223 799
rect 2299 795 2303 799
rect 2335 795 2339 799
rect 2475 795 2479 799
rect 2587 795 2591 799
rect 2663 795 2667 799
rect 2835 795 2839 799
rect 2859 795 2863 799
rect 3091 795 3095 799
rect 3211 795 3215 799
rect 3395 795 3399 799
rect 3415 795 3419 799
rect 3535 795 3539 799
rect 1871 787 1875 791
rect 2159 784 2163 788
rect 2239 784 2243 788
rect 2319 784 2323 788
rect 2415 784 2419 788
rect 2527 784 2531 788
rect 2647 784 2651 788
rect 2775 784 2779 788
rect 2903 784 2907 788
rect 3031 784 3035 788
rect 3151 784 3155 788
rect 3271 784 3275 788
rect 3399 784 3403 788
rect 3503 784 3507 788
rect 3591 787 3595 791
rect 111 757 115 761
rect 135 760 139 764
rect 263 760 267 764
rect 431 760 435 764
rect 607 760 611 764
rect 783 760 787 764
rect 951 760 955 764
rect 1103 760 1107 764
rect 1247 760 1251 764
rect 1383 760 1387 764
rect 1511 760 1515 764
rect 1639 760 1643 764
rect 1743 760 1747 764
rect 1831 757 1835 761
rect 219 751 223 755
rect 331 751 335 755
rect 111 740 115 744
rect 323 743 327 747
rect 851 751 855 755
rect 1211 751 1215 755
rect 1339 751 1343 755
rect 1471 751 1475 755
rect 1599 751 1603 755
rect 1711 751 1715 755
rect 887 743 891 747
rect 1699 743 1703 747
rect 1831 740 1835 744
rect 1871 729 1875 733
rect 1895 732 1899 736
rect 1975 732 1979 736
rect 2071 732 2075 736
rect 2183 732 2187 736
rect 2311 732 2315 736
rect 2447 732 2451 736
rect 2591 732 2595 736
rect 2743 732 2747 736
rect 2895 732 2899 736
rect 3047 732 3051 736
rect 3199 732 3203 736
rect 3359 732 3363 736
rect 3503 732 3507 736
rect 3591 729 3595 733
rect 143 722 147 726
rect 271 722 275 726
rect 439 722 443 726
rect 615 722 619 726
rect 791 722 795 726
rect 959 722 963 726
rect 1111 722 1115 726
rect 1255 722 1259 726
rect 1391 722 1395 726
rect 1519 722 1523 726
rect 1647 722 1651 726
rect 1751 722 1755 726
rect 1971 719 1975 723
rect 2051 723 2055 727
rect 2139 723 2143 727
rect 2403 723 2407 727
rect 167 711 168 715
rect 168 711 171 715
rect 219 711 223 715
rect 331 711 335 715
rect 851 711 855 715
rect 967 711 971 715
rect 1199 711 1203 715
rect 1211 711 1215 715
rect 1339 711 1343 715
rect 1471 711 1475 715
rect 1599 711 1603 715
rect 1699 711 1703 715
rect 1871 712 1875 716
rect 2131 715 2135 719
rect 2263 715 2267 719
rect 2515 723 2519 727
rect 2659 723 2663 727
rect 2811 723 2815 727
rect 3055 719 3059 723
rect 3115 723 3119 727
rect 3267 723 3271 727
rect 3563 715 3567 719
rect 3591 712 3595 716
rect 1903 694 1907 698
rect 1983 694 1987 698
rect 2079 694 2083 698
rect 2191 694 2195 698
rect 2319 694 2323 698
rect 2455 694 2459 698
rect 2599 694 2603 698
rect 2751 694 2755 698
rect 2903 694 2907 698
rect 3055 694 3059 698
rect 3207 694 3211 698
rect 3367 694 3371 698
rect 3511 694 3515 698
rect 323 687 324 691
rect 324 687 327 691
rect 347 687 351 691
rect 459 687 463 691
rect 715 687 719 691
rect 775 687 779 691
rect 835 687 839 691
rect 1059 687 1063 691
rect 1075 687 1079 691
rect 1187 687 1191 691
rect 1299 687 1303 691
rect 1403 687 1407 691
rect 1507 687 1511 691
rect 1707 687 1711 691
rect 1715 687 1719 691
rect 295 678 299 682
rect 407 678 411 682
rect 527 678 531 682
rect 655 678 659 682
rect 783 678 787 682
rect 903 678 907 682
rect 1023 678 1027 682
rect 1135 678 1139 682
rect 1247 678 1251 682
rect 1351 678 1355 682
rect 1455 678 1459 682
rect 1559 678 1563 682
rect 1663 678 1667 682
rect 1751 678 1755 682
rect 1971 683 1975 687
rect 2051 683 2055 687
rect 2263 683 2267 687
rect 2299 683 2303 687
rect 2403 683 2407 687
rect 2659 683 2663 687
rect 2811 683 2815 687
rect 2835 683 2839 687
rect 3115 683 3119 687
rect 3267 683 3271 687
rect 3391 683 3392 687
rect 3392 683 3395 687
rect 3535 683 3536 687
rect 3536 683 3539 687
rect 2139 675 2143 679
rect 111 660 115 664
rect 347 651 351 655
rect 459 651 463 655
rect 579 651 583 655
rect 775 651 779 655
rect 835 651 839 655
rect 967 651 971 655
rect 1075 651 1079 655
rect 1187 651 1191 655
rect 1299 651 1303 655
rect 1403 651 1407 655
rect 1507 651 1511 655
rect 1567 651 1571 655
rect 1715 651 1719 655
rect 2131 667 2135 671
rect 2147 667 2151 671
rect 2515 667 2519 671
rect 2531 667 2535 671
rect 2875 667 2879 671
rect 2883 667 2887 671
rect 3175 667 3179 671
rect 3235 667 3239 671
rect 3563 667 3567 671
rect 1831 660 1835 664
rect 1903 658 1907 662
rect 2095 658 2099 662
rect 2295 658 2299 662
rect 2479 658 2483 662
rect 2655 658 2659 662
rect 2831 658 2835 662
rect 3007 658 3011 662
rect 3183 658 3187 662
rect 3359 658 3363 662
rect 3511 658 3515 662
rect 111 643 115 647
rect 287 640 291 644
rect 399 640 403 644
rect 519 640 523 644
rect 647 640 651 644
rect 775 640 779 644
rect 895 640 899 644
rect 1015 640 1019 644
rect 1127 640 1131 644
rect 1239 640 1243 644
rect 1343 640 1347 644
rect 1447 640 1451 644
rect 1551 640 1555 644
rect 1655 640 1659 644
rect 1743 640 1747 644
rect 1831 643 1835 647
rect 1871 640 1875 644
rect 3591 640 3595 644
rect 1927 631 1931 635
rect 2147 631 2151 635
rect 2303 631 2307 635
rect 2531 631 2535 635
rect 2679 631 2683 635
rect 2883 631 2887 635
rect 3175 631 3179 635
rect 3235 631 3239 635
rect 3391 631 3395 635
rect 3535 631 3539 635
rect 1871 623 1875 627
rect 1895 620 1899 624
rect 2087 620 2091 624
rect 2287 620 2291 624
rect 2471 620 2475 624
rect 2647 620 2651 624
rect 2823 620 2827 624
rect 2999 620 3003 624
rect 3175 620 3179 624
rect 3351 620 3355 624
rect 3503 620 3507 624
rect 3591 623 3595 627
rect 111 589 115 593
rect 311 592 315 596
rect 391 592 395 596
rect 471 592 475 596
rect 559 592 563 596
rect 647 592 651 596
rect 735 592 739 596
rect 823 592 827 596
rect 911 592 915 596
rect 999 592 1003 596
rect 1087 592 1091 596
rect 1175 592 1179 596
rect 1263 592 1267 596
rect 1831 589 1835 593
rect 267 583 271 587
rect 379 583 383 587
rect 459 583 463 587
rect 539 583 543 587
rect 715 583 719 587
rect 891 583 895 587
rect 979 583 983 587
rect 1067 583 1071 587
rect 1155 583 1159 587
rect 1243 583 1247 587
rect 111 572 115 576
rect 707 575 711 579
rect 1059 575 1063 579
rect 1831 572 1835 576
rect 1871 569 1875 573
rect 1895 572 1899 576
rect 1975 572 1979 576
rect 2087 572 2091 576
rect 2215 572 2219 576
rect 2351 572 2355 576
rect 2495 572 2499 576
rect 2647 572 2651 576
rect 2807 572 2811 576
rect 2975 572 2979 576
rect 3151 572 3155 576
rect 3335 572 3339 576
rect 3503 572 3507 576
rect 3591 569 3595 573
rect 1963 563 1967 567
rect 2059 563 2063 567
rect 2163 563 2167 567
rect 2299 563 2303 567
rect 2443 563 2447 567
rect 2451 563 2455 567
rect 2747 563 2751 567
rect 2875 563 2879 567
rect 3043 563 3047 567
rect 3219 563 3223 567
rect 319 554 323 558
rect 399 554 403 558
rect 479 554 483 558
rect 567 554 571 558
rect 655 554 659 558
rect 743 554 747 558
rect 831 554 835 558
rect 919 554 923 558
rect 1007 554 1011 558
rect 1095 554 1099 558
rect 1183 554 1187 558
rect 1271 554 1275 558
rect 1871 552 1875 556
rect 2867 555 2871 559
rect 3563 555 3567 559
rect 3591 552 3595 556
rect 379 543 383 547
rect 459 543 463 547
rect 539 543 543 547
rect 579 543 583 547
rect 623 543 627 547
rect 707 543 711 547
rect 883 543 887 547
rect 891 543 895 547
rect 979 543 983 547
rect 1067 543 1071 547
rect 1155 543 1159 547
rect 1243 543 1247 547
rect 1903 534 1907 538
rect 1983 534 1987 538
rect 2095 534 2099 538
rect 2223 534 2227 538
rect 2359 534 2363 538
rect 2503 534 2507 538
rect 2655 534 2659 538
rect 2815 534 2819 538
rect 2983 534 2987 538
rect 3159 534 3163 538
rect 3343 534 3347 538
rect 3511 534 3515 538
rect 267 519 268 523
rect 268 519 271 523
rect 291 519 295 523
rect 467 519 468 523
rect 468 519 471 523
rect 491 519 495 523
rect 787 527 791 531
rect 683 519 687 523
rect 771 519 775 523
rect 859 519 863 523
rect 947 519 951 523
rect 1035 519 1039 523
rect 1123 519 1127 523
rect 1211 519 1215 523
rect 1927 523 1928 527
rect 1928 523 1931 527
rect 1963 523 1967 527
rect 2059 523 2063 527
rect 2163 523 2167 527
rect 2299 523 2303 527
rect 2443 523 2447 527
rect 2679 523 2680 527
rect 2680 523 2683 527
rect 2747 523 2751 527
rect 3043 523 3047 527
rect 3219 523 3223 527
rect 3367 523 3368 527
rect 3368 523 3371 527
rect 3535 523 3536 527
rect 3536 523 3539 527
rect 239 510 243 514
rect 343 510 347 514
rect 439 510 443 514
rect 535 510 539 514
rect 631 510 635 514
rect 719 510 723 514
rect 807 510 811 514
rect 895 510 899 514
rect 983 510 987 514
rect 1071 510 1075 514
rect 1159 510 1163 514
rect 1247 510 1251 514
rect 2179 511 2180 515
rect 2180 511 2183 515
rect 2203 511 2207 515
rect 2283 511 2287 515
rect 2379 511 2383 515
rect 2483 511 2487 515
rect 2603 511 2607 515
rect 2867 511 2868 515
rect 2868 511 2871 515
rect 2891 511 2895 515
rect 3203 511 3204 515
rect 3204 511 3207 515
rect 3227 511 3231 515
rect 3563 511 3567 515
rect 2151 502 2155 506
rect 2231 502 2235 506
rect 2327 502 2331 506
rect 2431 502 2435 506
rect 2551 502 2555 506
rect 2687 502 2691 506
rect 2839 502 2843 506
rect 2999 502 3003 506
rect 3175 502 3179 506
rect 3351 502 3355 506
rect 3511 502 3515 506
rect 111 492 115 496
rect 1831 492 1835 496
rect 291 483 295 487
rect 395 483 399 487
rect 491 483 495 487
rect 623 483 627 487
rect 683 483 687 487
rect 771 483 775 487
rect 859 483 863 487
rect 947 483 951 487
rect 1035 483 1039 487
rect 1123 483 1127 487
rect 1211 483 1215 487
rect 1255 483 1259 487
rect 1871 484 1875 488
rect 3591 484 3595 488
rect 111 475 115 479
rect 231 472 235 476
rect 335 472 339 476
rect 431 472 435 476
rect 527 472 531 476
rect 623 472 627 476
rect 711 472 715 476
rect 799 472 803 476
rect 887 472 891 476
rect 975 472 979 476
rect 1063 472 1067 476
rect 1151 472 1155 476
rect 1239 472 1243 476
rect 1831 475 1835 479
rect 2203 475 2207 479
rect 2283 475 2287 479
rect 2379 475 2383 479
rect 2483 475 2487 479
rect 2603 475 2607 479
rect 2719 475 2723 479
rect 2891 475 2895 479
rect 3051 475 3055 479
rect 3227 475 3231 479
rect 3367 475 3371 479
rect 3535 475 3539 479
rect 1871 467 1875 471
rect 2143 464 2147 468
rect 2223 464 2227 468
rect 2319 464 2323 468
rect 2423 464 2427 468
rect 2543 464 2547 468
rect 2679 464 2683 468
rect 2831 464 2835 468
rect 2991 464 2995 468
rect 3167 464 3171 468
rect 3343 464 3347 468
rect 3503 464 3507 468
rect 3591 467 3595 471
rect 111 417 115 421
rect 135 420 139 424
rect 247 420 251 424
rect 375 420 379 424
rect 495 420 499 424
rect 607 420 611 424
rect 719 420 723 424
rect 823 420 827 424
rect 919 420 923 424
rect 1007 420 1011 424
rect 1103 420 1107 424
rect 1199 420 1203 424
rect 1295 420 1299 424
rect 1831 417 1835 421
rect 203 411 207 415
rect 315 411 319 415
rect 467 411 471 415
rect 563 411 567 415
rect 675 411 679 415
rect 787 411 791 415
rect 891 411 895 415
rect 987 411 991 415
rect 1075 411 1079 415
rect 1271 411 1275 415
rect 1871 413 1875 417
rect 2335 416 2339 420
rect 2415 416 2419 420
rect 2495 416 2499 420
rect 2583 416 2587 420
rect 2687 416 2691 420
rect 2799 416 2803 420
rect 2927 416 2931 420
rect 3071 416 3075 420
rect 3215 416 3219 420
rect 3367 416 3371 420
rect 3503 416 3507 420
rect 111 400 115 404
rect 195 403 199 407
rect 1163 403 1167 407
rect 3591 413 3595 417
rect 2403 407 2407 411
rect 2483 407 2487 411
rect 1831 400 1835 404
rect 1871 396 1875 400
rect 2395 399 2399 403
rect 2563 407 2567 411
rect 2651 407 2655 411
rect 2799 403 2803 407
rect 2867 407 2871 411
rect 2995 407 2999 411
rect 3203 407 3207 411
rect 3283 407 3287 411
rect 3435 407 3439 411
rect 3591 396 3595 400
rect 143 382 147 386
rect 255 382 259 386
rect 383 382 387 386
rect 503 382 507 386
rect 615 382 619 386
rect 727 382 731 386
rect 831 382 835 386
rect 927 382 931 386
rect 1015 382 1019 386
rect 1111 382 1115 386
rect 1207 382 1211 386
rect 1303 382 1307 386
rect 2343 378 2347 382
rect 2423 378 2427 382
rect 2503 378 2507 382
rect 2591 378 2595 382
rect 2695 378 2699 382
rect 2807 378 2811 382
rect 2935 378 2939 382
rect 3079 378 3083 382
rect 3223 378 3227 382
rect 3375 378 3379 382
rect 3511 378 3515 382
rect 203 371 207 375
rect 315 371 319 375
rect 395 371 399 375
rect 563 371 567 375
rect 675 371 679 375
rect 783 371 787 375
rect 891 371 895 375
rect 987 371 991 375
rect 1075 371 1079 375
rect 1163 371 1167 375
rect 1171 371 1175 375
rect 1271 371 1275 375
rect 2395 367 2399 371
rect 2403 367 2407 371
rect 2483 371 2487 375
rect 2519 371 2523 375
rect 2563 367 2567 371
rect 2651 367 2655 371
rect 2719 367 2720 371
rect 2720 367 2723 371
rect 2867 367 2871 371
rect 2995 367 2999 371
rect 3051 367 3055 371
rect 3283 367 3287 371
rect 3339 367 3343 371
rect 3535 367 3536 371
rect 3536 367 3539 371
rect 195 347 199 351
rect 299 347 303 351
rect 427 347 431 351
rect 663 347 667 351
rect 699 347 703 351
rect 1231 355 1235 359
rect 1031 347 1032 351
rect 1032 347 1035 351
rect 1059 347 1063 351
rect 1447 355 1451 359
rect 1343 347 1347 351
rect 1379 347 1383 351
rect 2271 355 2275 359
rect 2131 347 2135 351
rect 2383 347 2387 351
rect 2647 355 2651 359
rect 2527 347 2528 351
rect 2528 347 2531 351
rect 2555 347 2559 351
rect 2799 347 2800 351
rect 2800 347 2803 351
rect 2827 347 2831 351
rect 3067 347 3068 351
rect 3068 347 3071 351
rect 3091 347 3095 351
rect 3279 347 3283 351
rect 3435 347 3436 351
rect 3436 347 3439 351
rect 3459 347 3463 351
rect 143 338 147 342
rect 247 338 251 342
rect 375 338 379 342
rect 511 338 515 342
rect 647 338 651 342
rect 775 338 779 342
rect 895 338 899 342
rect 1007 338 1011 342
rect 1119 338 1123 342
rect 1223 338 1227 342
rect 1327 338 1331 342
rect 1439 338 1443 342
rect 2079 338 2083 342
rect 2167 338 2171 342
rect 2263 338 2267 342
rect 2375 338 2379 342
rect 2503 338 2507 342
rect 2639 338 2643 342
rect 2775 338 2779 342
rect 2911 338 2915 342
rect 3039 338 3043 342
rect 3167 338 3171 342
rect 3287 338 3291 342
rect 3407 338 3411 342
rect 3511 338 3515 342
rect 111 320 115 324
rect 1831 320 1835 324
rect 1871 320 1875 324
rect 3591 320 3595 324
rect 299 311 303 315
rect 427 311 431 315
rect 699 311 703 315
rect 783 311 787 315
rect 1007 311 1011 315
rect 1059 311 1063 315
rect 1171 311 1175 315
rect 1231 311 1235 315
rect 1379 311 1383 315
rect 1447 311 1451 315
rect 2131 311 2135 315
rect 2239 311 2243 315
rect 2271 311 2275 315
rect 2383 311 2387 315
rect 2555 311 2559 315
rect 2647 311 2651 315
rect 2827 311 2831 315
rect 2963 311 2967 315
rect 3091 311 3095 315
rect 3279 311 3283 315
rect 3339 311 3343 315
rect 3459 311 3463 315
rect 3535 311 3539 315
rect 111 303 115 307
rect 135 300 139 304
rect 239 300 243 304
rect 367 300 371 304
rect 503 300 507 304
rect 639 300 643 304
rect 767 300 771 304
rect 887 300 891 304
rect 999 300 1003 304
rect 1111 300 1115 304
rect 1215 300 1219 304
rect 1319 300 1323 304
rect 1431 300 1435 304
rect 1831 303 1835 307
rect 1871 303 1875 307
rect 2071 300 2075 304
rect 2159 300 2163 304
rect 2255 300 2259 304
rect 2367 300 2371 304
rect 2495 300 2499 304
rect 2631 300 2635 304
rect 2767 300 2771 304
rect 2903 300 2907 304
rect 3031 300 3035 304
rect 3159 300 3163 304
rect 3279 300 3283 304
rect 3399 300 3403 304
rect 3503 300 3507 304
rect 3591 303 3595 307
rect 511 283 515 287
rect 111 245 115 249
rect 223 248 227 252
rect 335 248 339 252
rect 463 248 467 252
rect 599 248 603 252
rect 735 248 739 252
rect 871 248 875 252
rect 1007 248 1011 252
rect 1135 248 1139 252
rect 1255 248 1259 252
rect 1367 248 1371 252
rect 1479 248 1483 252
rect 1599 248 1603 252
rect 1831 245 1835 249
rect 1871 245 1875 249
rect 1895 248 1899 252
rect 1983 248 1987 252
rect 2095 248 2099 252
rect 2223 248 2227 252
rect 2359 248 2363 252
rect 2503 248 2507 252
rect 2647 248 2651 252
rect 2791 248 2795 252
rect 2935 248 2939 252
rect 3079 248 3083 252
rect 3223 248 3227 252
rect 3375 248 3379 252
rect 3503 248 3507 252
rect 3591 245 3595 249
rect 187 239 191 243
rect 291 239 295 243
rect 403 239 407 243
rect 667 239 671 243
rect 803 239 807 243
rect 1079 239 1083 243
rect 1211 239 1215 243
rect 1343 239 1347 243
rect 1447 239 1451 243
rect 1563 239 1567 243
rect 1571 239 1575 243
rect 1963 239 1967 243
rect 2063 239 2067 243
rect 2163 239 2167 243
rect 2315 239 2319 243
rect 2451 239 2455 243
rect 2459 239 2463 243
rect 2611 239 2615 243
rect 2715 239 2719 243
rect 2879 239 2883 243
rect 3067 239 3071 243
rect 3147 239 3151 243
rect 3291 239 3295 243
rect 111 228 115 232
rect 659 231 663 235
rect 1831 228 1835 232
rect 1871 228 1875 232
rect 3591 228 3595 232
rect 231 210 235 214
rect 343 210 347 214
rect 471 210 475 214
rect 607 210 611 214
rect 743 210 747 214
rect 879 210 883 214
rect 1015 210 1019 214
rect 1143 210 1147 214
rect 1263 210 1267 214
rect 1375 210 1379 214
rect 1487 210 1491 214
rect 1607 210 1611 214
rect 1903 210 1907 214
rect 1991 210 1995 214
rect 2103 210 2107 214
rect 2231 210 2235 214
rect 2367 210 2371 214
rect 2511 210 2515 214
rect 2655 210 2659 214
rect 2799 210 2803 214
rect 2943 210 2947 214
rect 3087 210 3091 214
rect 3231 210 3235 214
rect 3383 210 3387 214
rect 3511 210 3515 214
rect 291 199 295 203
rect 403 199 407 203
rect 511 199 515 203
rect 667 199 671 203
rect 803 199 807 203
rect 903 199 904 203
rect 904 199 907 203
rect 1043 199 1044 203
rect 1044 199 1047 203
rect 1079 199 1083 203
rect 1211 199 1215 203
rect 1159 191 1163 195
rect 1447 199 1451 203
rect 1563 199 1567 203
rect 1931 199 1932 203
rect 1932 199 1935 203
rect 1963 199 1967 203
rect 2063 199 2067 203
rect 2239 199 2243 203
rect 2315 199 2319 203
rect 2451 199 2455 203
rect 2715 199 2719 203
rect 2879 199 2883 203
rect 2963 199 2967 203
rect 3147 199 3151 203
rect 3291 199 3295 203
rect 3407 199 3408 203
rect 3408 199 3411 203
rect 3535 199 3536 203
rect 3536 199 3539 203
rect 1963 175 1967 179
rect 2095 175 2099 179
rect 2155 171 2159 175
rect 2163 175 2167 179
rect 2259 175 2263 179
rect 2387 175 2391 179
rect 2611 175 2612 179
rect 2612 175 2615 179
rect 2635 175 2639 179
rect 2755 175 2759 179
rect 2867 175 2871 179
rect 2971 175 2975 179
rect 3067 175 3071 179
rect 3163 175 3167 179
rect 3259 175 3263 179
rect 3355 175 3359 179
rect 187 155 188 159
rect 188 155 191 159
rect 211 155 215 159
rect 291 155 295 159
rect 371 155 375 159
rect 451 155 455 159
rect 531 155 535 159
rect 639 155 643 159
rect 699 155 703 159
rect 787 155 791 159
rect 1175 163 1179 167
rect 1903 166 1907 170
rect 1983 166 1987 170
rect 2087 166 2091 170
rect 2207 166 2211 170
rect 2335 166 2339 170
rect 2463 166 2467 170
rect 2583 166 2587 170
rect 2703 166 2707 170
rect 2815 166 2819 170
rect 2919 166 2923 170
rect 3015 166 3019 170
rect 3111 166 3115 170
rect 3207 166 3211 170
rect 3303 166 3307 170
rect 3399 166 3403 170
rect 1023 155 1024 159
rect 1024 155 1027 159
rect 1051 155 1055 159
rect 1255 155 1259 159
rect 1343 155 1347 159
rect 1431 155 1435 159
rect 1519 155 1523 159
rect 1599 155 1603 159
rect 1679 155 1683 159
rect 1759 155 1763 159
rect 159 146 163 150
rect 239 146 243 150
rect 319 146 323 150
rect 399 146 403 150
rect 479 146 483 150
rect 559 146 563 150
rect 647 146 651 150
rect 735 146 739 150
rect 823 146 827 150
rect 911 146 915 150
rect 999 146 1003 150
rect 1087 146 1091 150
rect 1167 146 1171 150
rect 1247 146 1251 150
rect 1335 146 1339 150
rect 1423 146 1427 150
rect 1511 146 1515 150
rect 1591 146 1595 150
rect 1671 146 1675 150
rect 1751 146 1755 150
rect 1871 148 1875 152
rect 3591 148 3595 152
rect 1963 139 1967 143
rect 2095 139 2099 143
rect 2259 139 2263 143
rect 2387 139 2391 143
rect 2471 139 2475 143
rect 2635 139 2639 143
rect 2755 139 2759 143
rect 2867 139 2871 143
rect 2971 139 2975 143
rect 3067 139 3071 143
rect 3163 139 3167 143
rect 3259 139 3263 143
rect 3355 139 3359 143
rect 3407 139 3411 143
rect 111 128 115 132
rect 1831 128 1835 132
rect 1871 131 1875 135
rect 1895 128 1899 132
rect 1975 128 1979 132
rect 2079 128 2083 132
rect 2199 128 2203 132
rect 2327 128 2331 132
rect 2455 128 2459 132
rect 2575 128 2579 132
rect 2695 128 2699 132
rect 2807 128 2811 132
rect 2911 128 2915 132
rect 3007 128 3011 132
rect 3103 128 3107 132
rect 3199 128 3203 132
rect 3295 128 3299 132
rect 3391 128 3395 132
rect 3591 131 3595 135
rect 211 119 215 123
rect 291 119 295 123
rect 371 119 375 123
rect 451 119 455 123
rect 531 119 535 123
rect 639 119 643 123
rect 699 119 703 123
rect 787 119 791 123
rect 903 119 907 123
rect 999 119 1003 123
rect 1051 119 1055 123
rect 1159 119 1163 123
rect 1175 119 1179 123
rect 1255 119 1259 123
rect 1343 119 1347 123
rect 1431 119 1435 123
rect 1519 119 1523 123
rect 1599 119 1603 123
rect 1679 119 1683 123
rect 1759 119 1763 123
rect 111 111 115 115
rect 151 108 155 112
rect 231 108 235 112
rect 311 108 315 112
rect 391 108 395 112
rect 471 108 475 112
rect 551 108 555 112
rect 639 108 643 112
rect 727 108 731 112
rect 815 108 819 112
rect 903 108 907 112
rect 991 108 995 112
rect 1079 108 1083 112
rect 1159 108 1163 112
rect 1239 108 1243 112
rect 1327 108 1331 112
rect 1415 108 1419 112
rect 1503 108 1507 112
rect 1583 108 1587 112
rect 1663 108 1667 112
rect 1743 108 1747 112
rect 1831 111 1835 115
<< m3 >>
rect 1871 3670 1875 3671
rect 1871 3665 1875 3666
rect 2151 3670 2155 3671
rect 2151 3665 2155 3666
rect 2439 3670 2443 3671
rect 2439 3665 2443 3666
rect 2727 3670 2731 3671
rect 2727 3665 2731 3666
rect 3015 3670 3019 3671
rect 3015 3665 3019 3666
rect 3591 3670 3595 3671
rect 3591 3665 3595 3666
rect 1872 3646 1874 3665
rect 2152 3649 2154 3665
rect 2440 3649 2442 3665
rect 2728 3649 2730 3665
rect 3016 3649 3018 3665
rect 2150 3648 2156 3649
rect 1870 3645 1876 3646
rect 111 3642 115 3643
rect 111 3637 115 3638
rect 143 3642 147 3643
rect 143 3637 147 3638
rect 239 3642 243 3643
rect 239 3637 243 3638
rect 367 3642 371 3643
rect 367 3637 371 3638
rect 503 3642 507 3643
rect 503 3637 507 3638
rect 639 3642 643 3643
rect 639 3637 643 3638
rect 775 3642 779 3643
rect 775 3637 779 3638
rect 911 3642 915 3643
rect 911 3637 915 3638
rect 1055 3642 1059 3643
rect 1055 3637 1059 3638
rect 1199 3642 1203 3643
rect 1199 3637 1203 3638
rect 1831 3642 1835 3643
rect 1870 3641 1871 3645
rect 1875 3641 1876 3645
rect 2150 3644 2151 3648
rect 2155 3644 2156 3648
rect 2150 3643 2156 3644
rect 2438 3648 2444 3649
rect 2438 3644 2439 3648
rect 2443 3644 2444 3648
rect 2438 3643 2444 3644
rect 2726 3648 2732 3649
rect 2726 3644 2727 3648
rect 2731 3644 2732 3648
rect 2726 3643 2732 3644
rect 3014 3648 3020 3649
rect 3014 3644 3015 3648
rect 3019 3644 3020 3648
rect 3592 3646 3594 3665
rect 3014 3643 3020 3644
rect 3590 3645 3596 3646
rect 1870 3640 1876 3641
rect 3590 3641 3591 3645
rect 3595 3641 3596 3645
rect 3590 3640 3596 3641
rect 1831 3637 1835 3638
rect 2242 3639 2248 3640
rect 112 3609 114 3637
rect 144 3627 146 3637
rect 194 3635 200 3636
rect 194 3631 195 3635
rect 199 3631 200 3635
rect 194 3630 200 3631
rect 142 3626 148 3627
rect 142 3622 143 3626
rect 147 3622 148 3626
rect 142 3621 148 3622
rect 110 3608 116 3609
rect 110 3604 111 3608
rect 115 3604 116 3608
rect 110 3603 116 3604
rect 196 3600 198 3630
rect 240 3627 242 3637
rect 290 3635 296 3636
rect 290 3631 291 3635
rect 295 3631 296 3635
rect 290 3630 296 3631
rect 238 3626 244 3627
rect 238 3622 239 3626
rect 243 3622 244 3626
rect 238 3621 244 3622
rect 292 3600 294 3630
rect 368 3627 370 3637
rect 418 3635 424 3636
rect 418 3631 419 3635
rect 423 3631 424 3635
rect 418 3630 424 3631
rect 366 3626 372 3627
rect 366 3622 367 3626
rect 371 3622 372 3626
rect 366 3621 372 3622
rect 420 3600 422 3630
rect 504 3627 506 3637
rect 554 3635 560 3636
rect 554 3631 555 3635
rect 559 3631 560 3635
rect 554 3630 560 3631
rect 502 3626 508 3627
rect 502 3622 503 3626
rect 507 3622 508 3626
rect 502 3621 508 3622
rect 556 3600 558 3630
rect 640 3627 642 3637
rect 776 3627 778 3637
rect 802 3635 808 3636
rect 802 3631 803 3635
rect 807 3631 808 3635
rect 802 3630 808 3631
rect 826 3635 832 3636
rect 826 3631 827 3635
rect 831 3631 832 3635
rect 826 3630 832 3631
rect 638 3626 644 3627
rect 638 3622 639 3626
rect 643 3622 644 3626
rect 638 3621 644 3622
rect 774 3626 780 3627
rect 774 3622 775 3626
rect 779 3622 780 3626
rect 774 3621 780 3622
rect 194 3599 200 3600
rect 194 3595 195 3599
rect 199 3595 200 3599
rect 194 3594 200 3595
rect 290 3599 296 3600
rect 290 3595 291 3599
rect 295 3595 296 3599
rect 290 3594 296 3595
rect 418 3599 424 3600
rect 418 3595 419 3599
rect 423 3595 424 3599
rect 418 3594 424 3595
rect 554 3599 560 3600
rect 554 3595 555 3599
rect 559 3595 560 3599
rect 554 3594 560 3595
rect 110 3591 116 3592
rect 110 3587 111 3591
rect 115 3587 116 3591
rect 110 3586 116 3587
rect 134 3588 140 3589
rect 112 3567 114 3586
rect 134 3584 135 3588
rect 139 3584 140 3588
rect 134 3583 140 3584
rect 230 3588 236 3589
rect 230 3584 231 3588
rect 235 3584 236 3588
rect 230 3583 236 3584
rect 358 3588 364 3589
rect 358 3584 359 3588
rect 363 3584 364 3588
rect 358 3583 364 3584
rect 494 3588 500 3589
rect 494 3584 495 3588
rect 499 3584 500 3588
rect 494 3583 500 3584
rect 630 3588 636 3589
rect 630 3584 631 3588
rect 635 3584 636 3588
rect 630 3583 636 3584
rect 766 3588 772 3589
rect 766 3584 767 3588
rect 771 3584 772 3588
rect 766 3583 772 3584
rect 136 3567 138 3583
rect 232 3567 234 3583
rect 360 3567 362 3583
rect 450 3571 456 3572
rect 450 3567 451 3571
rect 455 3567 456 3571
rect 496 3567 498 3583
rect 632 3567 634 3583
rect 768 3567 770 3583
rect 804 3572 806 3630
rect 828 3600 830 3630
rect 912 3627 914 3637
rect 962 3635 968 3636
rect 962 3631 963 3635
rect 967 3631 968 3635
rect 962 3630 968 3631
rect 910 3626 916 3627
rect 910 3622 911 3626
rect 915 3622 916 3626
rect 910 3621 916 3622
rect 964 3600 966 3630
rect 1056 3627 1058 3637
rect 1106 3635 1112 3636
rect 1106 3631 1107 3635
rect 1111 3631 1112 3635
rect 1106 3630 1112 3631
rect 1054 3626 1060 3627
rect 1054 3622 1055 3626
rect 1059 3622 1060 3626
rect 1054 3621 1060 3622
rect 1108 3600 1110 3630
rect 1200 3627 1202 3637
rect 1198 3626 1204 3627
rect 1198 3622 1199 3626
rect 1203 3622 1204 3626
rect 1198 3621 1204 3622
rect 1832 3609 1834 3637
rect 2242 3635 2243 3639
rect 2247 3635 2248 3639
rect 2242 3634 2248 3635
rect 2510 3639 2516 3640
rect 2510 3635 2511 3639
rect 2515 3635 2516 3639
rect 2510 3634 2516 3635
rect 3086 3639 3092 3640
rect 3086 3635 3087 3639
rect 3091 3635 3092 3639
rect 3086 3634 3092 3635
rect 1870 3628 1876 3629
rect 1870 3624 1871 3628
rect 1875 3624 1876 3628
rect 1870 3623 1876 3624
rect 1830 3608 1836 3609
rect 1830 3604 1831 3608
rect 1835 3604 1836 3608
rect 1830 3603 1836 3604
rect 826 3599 832 3600
rect 826 3595 827 3599
rect 831 3595 832 3599
rect 826 3594 832 3595
rect 962 3599 968 3600
rect 962 3595 963 3599
rect 967 3595 968 3599
rect 962 3594 968 3595
rect 1106 3599 1112 3600
rect 1106 3595 1107 3599
rect 1111 3595 1112 3599
rect 1872 3595 1874 3623
rect 2158 3610 2164 3611
rect 2158 3606 2159 3610
rect 2163 3606 2164 3610
rect 2158 3605 2164 3606
rect 2160 3595 2162 3605
rect 2182 3599 2188 3600
rect 2182 3595 2183 3599
rect 2187 3595 2188 3599
rect 1106 3594 1112 3595
rect 1871 3594 1875 3595
rect 1830 3591 1836 3592
rect 902 3588 908 3589
rect 902 3584 903 3588
rect 907 3584 908 3588
rect 902 3583 908 3584
rect 1046 3588 1052 3589
rect 1046 3584 1047 3588
rect 1051 3584 1052 3588
rect 1046 3583 1052 3584
rect 1190 3588 1196 3589
rect 1190 3584 1191 3588
rect 1195 3584 1196 3588
rect 1830 3587 1831 3591
rect 1835 3587 1836 3591
rect 1871 3589 1875 3590
rect 1903 3594 1907 3595
rect 1903 3589 1907 3590
rect 1983 3594 1987 3595
rect 1983 3589 1987 3590
rect 2071 3594 2075 3595
rect 2071 3589 2075 3590
rect 2159 3594 2163 3595
rect 2159 3589 2163 3590
rect 2175 3594 2179 3595
rect 2182 3594 2188 3595
rect 2175 3589 2179 3590
rect 1830 3586 1836 3587
rect 1190 3583 1196 3584
rect 802 3571 808 3572
rect 802 3567 803 3571
rect 807 3567 808 3571
rect 904 3567 906 3583
rect 910 3571 916 3572
rect 910 3567 911 3571
rect 915 3567 916 3571
rect 1048 3567 1050 3583
rect 1054 3571 1060 3572
rect 1054 3567 1055 3571
rect 1059 3567 1060 3571
rect 1192 3567 1194 3583
rect 1832 3567 1834 3586
rect 111 3566 115 3567
rect 111 3561 115 3562
rect 135 3566 139 3567
rect 135 3561 139 3562
rect 183 3566 187 3567
rect 183 3561 187 3562
rect 231 3566 235 3567
rect 231 3561 235 3562
rect 303 3566 307 3567
rect 303 3561 307 3562
rect 359 3566 363 3567
rect 359 3561 363 3562
rect 415 3566 419 3567
rect 450 3566 456 3567
rect 495 3566 499 3567
rect 415 3561 419 3562
rect 112 3542 114 3561
rect 184 3545 186 3561
rect 304 3545 306 3561
rect 416 3545 418 3561
rect 182 3544 188 3545
rect 110 3541 116 3542
rect 110 3537 111 3541
rect 115 3537 116 3541
rect 182 3540 183 3544
rect 187 3540 188 3544
rect 182 3539 188 3540
rect 302 3544 308 3545
rect 302 3540 303 3544
rect 307 3540 308 3544
rect 302 3539 308 3540
rect 414 3544 420 3545
rect 414 3540 415 3544
rect 419 3540 420 3544
rect 414 3539 420 3540
rect 110 3536 116 3537
rect 258 3535 264 3536
rect 258 3531 259 3535
rect 263 3531 264 3535
rect 258 3530 264 3531
rect 382 3535 388 3536
rect 382 3531 383 3535
rect 387 3531 388 3535
rect 382 3530 388 3531
rect 242 3527 248 3528
rect 110 3524 116 3525
rect 110 3520 111 3524
rect 115 3520 116 3524
rect 242 3523 243 3527
rect 247 3523 248 3527
rect 242 3522 248 3523
rect 110 3519 116 3520
rect 112 3483 114 3519
rect 190 3506 196 3507
rect 190 3502 191 3506
rect 195 3502 196 3506
rect 190 3501 196 3502
rect 192 3483 194 3501
rect 244 3496 246 3522
rect 260 3496 262 3530
rect 310 3506 316 3507
rect 310 3502 311 3506
rect 315 3502 316 3506
rect 310 3501 316 3502
rect 242 3495 248 3496
rect 242 3491 243 3495
rect 247 3491 248 3495
rect 242 3490 248 3491
rect 258 3495 264 3496
rect 258 3491 259 3495
rect 263 3491 264 3495
rect 258 3490 264 3491
rect 312 3483 314 3501
rect 111 3482 115 3483
rect 111 3477 115 3478
rect 191 3482 195 3483
rect 191 3477 195 3478
rect 231 3482 235 3483
rect 231 3477 235 3478
rect 311 3482 315 3483
rect 311 3477 315 3478
rect 367 3482 371 3483
rect 367 3477 371 3478
rect 112 3449 114 3477
rect 232 3467 234 3477
rect 368 3467 370 3477
rect 384 3476 386 3530
rect 422 3506 428 3507
rect 422 3502 423 3506
rect 427 3502 428 3506
rect 422 3501 428 3502
rect 424 3483 426 3501
rect 452 3496 454 3566
rect 495 3561 499 3562
rect 527 3566 531 3567
rect 527 3561 531 3562
rect 631 3566 635 3567
rect 631 3561 635 3562
rect 735 3566 739 3567
rect 735 3561 739 3562
rect 767 3566 771 3567
rect 802 3566 808 3567
rect 831 3566 835 3567
rect 767 3561 771 3562
rect 831 3561 835 3562
rect 903 3566 907 3567
rect 910 3566 916 3567
rect 919 3566 923 3567
rect 903 3561 907 3562
rect 528 3545 530 3561
rect 632 3545 634 3561
rect 736 3545 738 3561
rect 832 3545 834 3561
rect 526 3544 532 3545
rect 526 3540 527 3544
rect 531 3540 532 3544
rect 526 3539 532 3540
rect 630 3544 636 3545
rect 630 3540 631 3544
rect 635 3540 636 3544
rect 630 3539 636 3540
rect 734 3544 740 3545
rect 734 3540 735 3544
rect 739 3540 740 3544
rect 734 3539 740 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 912 3536 914 3566
rect 919 3561 923 3562
rect 1007 3566 1011 3567
rect 1007 3561 1011 3562
rect 1047 3566 1051 3567
rect 1054 3566 1060 3567
rect 1095 3566 1099 3567
rect 1047 3561 1051 3562
rect 920 3545 922 3561
rect 1008 3545 1010 3561
rect 918 3544 924 3545
rect 918 3540 919 3544
rect 923 3540 924 3544
rect 918 3539 924 3540
rect 1006 3544 1012 3545
rect 1006 3540 1007 3544
rect 1011 3540 1012 3544
rect 1006 3539 1012 3540
rect 602 3535 608 3536
rect 602 3531 603 3535
rect 607 3531 608 3535
rect 602 3530 608 3531
rect 706 3535 712 3536
rect 706 3531 707 3535
rect 711 3531 712 3535
rect 706 3530 712 3531
rect 806 3535 812 3536
rect 806 3531 807 3535
rect 811 3531 812 3535
rect 806 3530 812 3531
rect 898 3535 904 3536
rect 898 3531 899 3535
rect 903 3531 904 3535
rect 898 3530 904 3531
rect 910 3535 916 3536
rect 910 3531 911 3535
rect 915 3531 916 3535
rect 910 3530 916 3531
rect 534 3506 540 3507
rect 534 3502 535 3506
rect 539 3502 540 3506
rect 534 3501 540 3502
rect 450 3495 456 3496
rect 450 3491 451 3495
rect 455 3491 456 3495
rect 450 3490 456 3491
rect 536 3483 538 3501
rect 604 3496 606 3530
rect 638 3506 644 3507
rect 638 3502 639 3506
rect 643 3502 644 3506
rect 638 3501 644 3502
rect 602 3495 608 3496
rect 602 3491 603 3495
rect 607 3491 608 3495
rect 602 3490 608 3491
rect 640 3483 642 3501
rect 708 3496 710 3530
rect 742 3506 748 3507
rect 742 3502 743 3506
rect 747 3502 748 3506
rect 742 3501 748 3502
rect 706 3495 712 3496
rect 706 3491 707 3495
rect 711 3491 712 3495
rect 706 3490 712 3491
rect 744 3483 746 3501
rect 808 3496 810 3530
rect 838 3506 844 3507
rect 838 3502 839 3506
rect 843 3502 844 3506
rect 838 3501 844 3502
rect 806 3495 812 3496
rect 806 3491 807 3495
rect 811 3491 812 3495
rect 806 3490 812 3491
rect 840 3483 842 3501
rect 900 3496 902 3530
rect 987 3508 991 3509
rect 926 3506 932 3507
rect 926 3502 927 3506
rect 931 3502 932 3506
rect 987 3503 991 3504
rect 1014 3506 1020 3507
rect 926 3501 932 3502
rect 898 3495 904 3496
rect 898 3491 899 3495
rect 903 3491 904 3495
rect 898 3490 904 3491
rect 846 3487 852 3488
rect 846 3483 847 3487
rect 851 3483 852 3487
rect 928 3483 930 3501
rect 423 3482 427 3483
rect 423 3477 427 3478
rect 503 3482 507 3483
rect 503 3477 507 3478
rect 535 3482 539 3483
rect 535 3477 539 3478
rect 623 3482 627 3483
rect 623 3477 627 3478
rect 639 3482 643 3483
rect 639 3477 643 3478
rect 735 3482 739 3483
rect 735 3477 739 3478
rect 743 3482 747 3483
rect 743 3477 747 3478
rect 839 3482 843 3483
rect 846 3482 852 3483
rect 927 3482 931 3483
rect 839 3477 843 3478
rect 374 3475 380 3476
rect 374 3471 375 3475
rect 379 3471 380 3475
rect 374 3470 380 3471
rect 382 3475 388 3476
rect 382 3471 383 3475
rect 387 3471 388 3475
rect 382 3470 388 3471
rect 230 3466 236 3467
rect 230 3462 231 3466
rect 235 3462 236 3466
rect 230 3461 236 3462
rect 366 3466 372 3467
rect 366 3462 367 3466
rect 371 3462 372 3466
rect 366 3461 372 3462
rect 110 3448 116 3449
rect 110 3444 111 3448
rect 115 3444 116 3448
rect 110 3443 116 3444
rect 376 3440 378 3470
rect 504 3467 506 3477
rect 518 3475 524 3476
rect 518 3471 519 3475
rect 523 3471 524 3475
rect 518 3470 524 3471
rect 554 3475 560 3476
rect 554 3471 555 3475
rect 559 3471 560 3475
rect 554 3470 560 3471
rect 502 3466 508 3467
rect 502 3462 503 3466
rect 507 3462 508 3466
rect 502 3461 508 3462
rect 374 3439 380 3440
rect 374 3435 375 3439
rect 379 3435 380 3439
rect 374 3434 380 3435
rect 110 3431 116 3432
rect 110 3427 111 3431
rect 115 3427 116 3431
rect 110 3426 116 3427
rect 222 3428 228 3429
rect 112 3403 114 3426
rect 222 3424 223 3428
rect 227 3424 228 3428
rect 222 3423 228 3424
rect 358 3428 364 3429
rect 358 3424 359 3428
rect 363 3424 364 3428
rect 358 3423 364 3424
rect 494 3428 500 3429
rect 494 3424 495 3428
rect 499 3424 500 3428
rect 494 3423 500 3424
rect 224 3403 226 3423
rect 242 3411 248 3412
rect 242 3407 243 3411
rect 247 3407 248 3411
rect 242 3406 248 3407
rect 111 3402 115 3403
rect 111 3397 115 3398
rect 215 3402 219 3403
rect 215 3397 219 3398
rect 223 3402 227 3403
rect 223 3397 227 3398
rect 112 3378 114 3397
rect 216 3381 218 3397
rect 214 3380 220 3381
rect 110 3377 116 3378
rect 110 3373 111 3377
rect 115 3373 116 3377
rect 214 3376 215 3380
rect 219 3376 220 3380
rect 214 3375 220 3376
rect 110 3372 116 3373
rect 110 3360 116 3361
rect 110 3356 111 3360
rect 115 3356 116 3360
rect 110 3355 116 3356
rect 112 3323 114 3355
rect 222 3342 228 3343
rect 222 3338 223 3342
rect 227 3338 228 3342
rect 222 3337 228 3338
rect 224 3323 226 3337
rect 244 3332 246 3406
rect 360 3403 362 3423
rect 496 3403 498 3423
rect 359 3402 363 3403
rect 359 3397 363 3398
rect 367 3402 371 3403
rect 367 3397 371 3398
rect 495 3402 499 3403
rect 495 3397 499 3398
rect 511 3402 515 3403
rect 511 3397 515 3398
rect 368 3381 370 3397
rect 512 3381 514 3397
rect 366 3380 372 3381
rect 366 3376 367 3380
rect 371 3376 372 3380
rect 366 3375 372 3376
rect 510 3380 516 3381
rect 510 3376 511 3380
rect 515 3376 516 3380
rect 510 3375 516 3376
rect 282 3371 288 3372
rect 282 3367 283 3371
rect 287 3367 288 3371
rect 520 3368 522 3470
rect 556 3440 558 3470
rect 624 3467 626 3477
rect 674 3475 680 3476
rect 674 3471 675 3475
rect 679 3471 680 3475
rect 674 3470 680 3471
rect 622 3466 628 3467
rect 622 3462 623 3466
rect 627 3462 628 3466
rect 622 3461 628 3462
rect 676 3440 678 3470
rect 736 3467 738 3477
rect 786 3475 792 3476
rect 786 3471 787 3475
rect 791 3471 792 3475
rect 786 3470 792 3471
rect 734 3466 740 3467
rect 734 3462 735 3466
rect 739 3462 740 3466
rect 734 3461 740 3462
rect 788 3440 790 3470
rect 840 3467 842 3477
rect 838 3466 844 3467
rect 838 3462 839 3466
rect 843 3462 844 3466
rect 838 3461 844 3462
rect 848 3440 850 3482
rect 927 3477 931 3478
rect 943 3482 947 3483
rect 943 3477 947 3478
rect 944 3467 946 3477
rect 988 3476 990 3503
rect 1014 3502 1015 3506
rect 1019 3502 1020 3506
rect 1014 3501 1020 3502
rect 1016 3483 1018 3501
rect 1056 3496 1058 3566
rect 1095 3561 1099 3562
rect 1183 3566 1187 3567
rect 1183 3561 1187 3562
rect 1191 3566 1195 3567
rect 1191 3561 1195 3562
rect 1271 3566 1275 3567
rect 1271 3561 1275 3562
rect 1359 3566 1363 3567
rect 1359 3561 1363 3562
rect 1447 3566 1451 3567
rect 1447 3561 1451 3562
rect 1831 3566 1835 3567
rect 1831 3561 1835 3562
rect 1872 3561 1874 3589
rect 1904 3579 1906 3589
rect 1930 3587 1936 3588
rect 1930 3583 1931 3587
rect 1935 3583 1936 3587
rect 1930 3582 1936 3583
rect 1954 3587 1960 3588
rect 1954 3583 1955 3587
rect 1959 3583 1960 3587
rect 1954 3582 1960 3583
rect 1902 3578 1908 3579
rect 1902 3574 1903 3578
rect 1907 3574 1908 3578
rect 1902 3573 1908 3574
rect 1096 3545 1098 3561
rect 1184 3545 1186 3561
rect 1272 3545 1274 3561
rect 1360 3545 1362 3561
rect 1448 3545 1450 3561
rect 1094 3544 1100 3545
rect 1094 3540 1095 3544
rect 1099 3540 1100 3544
rect 1094 3539 1100 3540
rect 1182 3544 1188 3545
rect 1182 3540 1183 3544
rect 1187 3540 1188 3544
rect 1182 3539 1188 3540
rect 1270 3544 1276 3545
rect 1270 3540 1271 3544
rect 1275 3540 1276 3544
rect 1270 3539 1276 3540
rect 1358 3544 1364 3545
rect 1358 3540 1359 3544
rect 1363 3540 1364 3544
rect 1358 3539 1364 3540
rect 1446 3544 1452 3545
rect 1446 3540 1447 3544
rect 1451 3540 1452 3544
rect 1832 3542 1834 3561
rect 1870 3560 1876 3561
rect 1870 3556 1871 3560
rect 1875 3556 1876 3560
rect 1870 3555 1876 3556
rect 1870 3543 1876 3544
rect 1446 3539 1452 3540
rect 1830 3541 1836 3542
rect 1830 3537 1831 3541
rect 1835 3537 1836 3541
rect 1870 3539 1871 3543
rect 1875 3539 1876 3543
rect 1870 3538 1876 3539
rect 1894 3540 1900 3541
rect 1830 3536 1836 3537
rect 1074 3535 1080 3536
rect 1074 3531 1075 3535
rect 1079 3531 1080 3535
rect 1074 3530 1080 3531
rect 1250 3535 1256 3536
rect 1250 3531 1251 3535
rect 1255 3531 1256 3535
rect 1250 3530 1256 3531
rect 1338 3535 1344 3536
rect 1338 3531 1339 3535
rect 1343 3531 1344 3535
rect 1338 3530 1344 3531
rect 1426 3535 1432 3536
rect 1426 3531 1427 3535
rect 1431 3531 1432 3535
rect 1426 3530 1432 3531
rect 1434 3535 1440 3536
rect 1434 3531 1435 3535
rect 1439 3531 1440 3535
rect 1434 3530 1440 3531
rect 1076 3496 1078 3530
rect 1102 3506 1108 3507
rect 1102 3502 1103 3506
rect 1107 3502 1108 3506
rect 1102 3501 1108 3502
rect 1190 3506 1196 3507
rect 1190 3502 1191 3506
rect 1195 3502 1196 3506
rect 1190 3501 1196 3502
rect 1054 3495 1060 3496
rect 1054 3491 1055 3495
rect 1059 3491 1060 3495
rect 1054 3490 1060 3491
rect 1074 3495 1080 3496
rect 1074 3491 1075 3495
rect 1079 3491 1080 3495
rect 1074 3490 1080 3491
rect 1104 3483 1106 3501
rect 1192 3483 1194 3501
rect 1252 3496 1254 3530
rect 1278 3506 1284 3507
rect 1278 3502 1279 3506
rect 1283 3502 1284 3506
rect 1278 3501 1284 3502
rect 1250 3495 1256 3496
rect 1250 3491 1251 3495
rect 1255 3491 1256 3495
rect 1250 3490 1256 3491
rect 1280 3483 1282 3501
rect 1340 3496 1342 3530
rect 1366 3506 1372 3507
rect 1366 3502 1367 3506
rect 1371 3502 1372 3506
rect 1366 3501 1372 3502
rect 1338 3495 1344 3496
rect 1338 3491 1339 3495
rect 1343 3491 1344 3495
rect 1338 3490 1344 3491
rect 1368 3483 1370 3501
rect 1428 3496 1430 3530
rect 1436 3509 1438 3530
rect 1830 3524 1836 3525
rect 1830 3520 1831 3524
rect 1835 3520 1836 3524
rect 1830 3519 1836 3520
rect 1872 3519 1874 3538
rect 1894 3536 1895 3540
rect 1899 3536 1900 3540
rect 1894 3535 1900 3536
rect 1896 3519 1898 3535
rect 1435 3508 1439 3509
rect 1435 3503 1439 3504
rect 1454 3506 1460 3507
rect 1454 3502 1455 3506
rect 1459 3502 1460 3506
rect 1454 3501 1460 3502
rect 1426 3495 1432 3496
rect 1426 3491 1427 3495
rect 1431 3491 1432 3495
rect 1426 3490 1432 3491
rect 1456 3483 1458 3501
rect 1832 3483 1834 3519
rect 1871 3518 1875 3519
rect 1871 3513 1875 3514
rect 1895 3518 1899 3519
rect 1895 3513 1899 3514
rect 1872 3494 1874 3513
rect 1870 3493 1876 3494
rect 1870 3489 1871 3493
rect 1875 3489 1876 3493
rect 1870 3488 1876 3489
rect 1932 3488 1934 3582
rect 1956 3552 1958 3582
rect 1984 3579 1986 3589
rect 2034 3587 2040 3588
rect 2034 3583 2035 3587
rect 2039 3583 2040 3587
rect 2034 3582 2040 3583
rect 1982 3578 1988 3579
rect 1982 3574 1983 3578
rect 1987 3574 1988 3578
rect 1982 3573 1988 3574
rect 2036 3552 2038 3582
rect 2072 3579 2074 3589
rect 2122 3587 2128 3588
rect 2122 3583 2123 3587
rect 2127 3583 2128 3587
rect 2122 3582 2128 3583
rect 2070 3578 2076 3579
rect 2070 3574 2071 3578
rect 2075 3574 2076 3578
rect 2070 3573 2076 3574
rect 2124 3552 2126 3582
rect 2176 3579 2178 3589
rect 2174 3578 2180 3579
rect 2174 3574 2175 3578
rect 2179 3574 2180 3578
rect 2174 3573 2180 3574
rect 2184 3552 2186 3594
rect 2244 3588 2246 3634
rect 2446 3610 2452 3611
rect 2446 3606 2447 3610
rect 2451 3606 2452 3610
rect 2446 3605 2452 3606
rect 2448 3595 2450 3605
rect 2512 3600 2514 3634
rect 2734 3610 2740 3611
rect 2734 3606 2735 3610
rect 2739 3606 2740 3610
rect 2734 3605 2740 3606
rect 3022 3610 3028 3611
rect 3022 3606 3023 3610
rect 3027 3606 3028 3610
rect 3022 3605 3028 3606
rect 2502 3599 2508 3600
rect 2502 3595 2503 3599
rect 2507 3595 2508 3599
rect 2295 3594 2299 3595
rect 2295 3589 2299 3590
rect 2423 3594 2427 3595
rect 2423 3589 2427 3590
rect 2447 3594 2451 3595
rect 2502 3594 2508 3595
rect 2510 3599 2516 3600
rect 2510 3595 2511 3599
rect 2515 3595 2516 3599
rect 2736 3595 2738 3605
rect 3024 3595 3026 3605
rect 2510 3594 2516 3595
rect 2559 3594 2563 3595
rect 2447 3589 2451 3590
rect 2242 3587 2248 3588
rect 2242 3583 2243 3587
rect 2247 3583 2248 3587
rect 2242 3582 2248 3583
rect 2296 3579 2298 3589
rect 2346 3587 2352 3588
rect 2346 3583 2347 3587
rect 2351 3583 2352 3587
rect 2346 3582 2352 3583
rect 2294 3578 2300 3579
rect 2294 3574 2295 3578
rect 2299 3574 2300 3578
rect 2294 3573 2300 3574
rect 2348 3552 2350 3582
rect 2424 3579 2426 3589
rect 2474 3587 2480 3588
rect 2474 3583 2475 3587
rect 2479 3583 2480 3587
rect 2474 3582 2480 3583
rect 2422 3578 2428 3579
rect 2422 3574 2423 3578
rect 2427 3574 2428 3578
rect 2422 3573 2428 3574
rect 2476 3552 2478 3582
rect 2504 3573 2506 3594
rect 2559 3589 2563 3590
rect 2695 3594 2699 3595
rect 2695 3589 2699 3590
rect 2735 3594 2739 3595
rect 2735 3589 2739 3590
rect 2831 3594 2835 3595
rect 2831 3589 2835 3590
rect 2975 3594 2979 3595
rect 2975 3589 2979 3590
rect 3023 3594 3027 3595
rect 3023 3589 3027 3590
rect 2560 3579 2562 3589
rect 2696 3579 2698 3589
rect 2746 3587 2752 3588
rect 2730 3583 2736 3584
rect 2730 3579 2731 3583
rect 2735 3579 2736 3583
rect 2746 3583 2747 3587
rect 2751 3583 2752 3587
rect 2746 3582 2752 3583
rect 2558 3578 2564 3579
rect 2558 3574 2559 3578
rect 2563 3574 2564 3578
rect 2558 3573 2564 3574
rect 2694 3578 2700 3579
rect 2730 3578 2736 3579
rect 2694 3574 2695 3578
rect 2699 3574 2700 3578
rect 2694 3573 2700 3574
rect 2503 3572 2507 3573
rect 2503 3567 2507 3568
rect 1954 3551 1960 3552
rect 1954 3547 1955 3551
rect 1959 3547 1960 3551
rect 1954 3546 1960 3547
rect 2034 3551 2040 3552
rect 2034 3547 2035 3551
rect 2039 3547 2040 3551
rect 2034 3546 2040 3547
rect 2122 3551 2128 3552
rect 2122 3547 2123 3551
rect 2127 3547 2128 3551
rect 2122 3546 2128 3547
rect 2182 3551 2188 3552
rect 2182 3547 2183 3551
rect 2187 3547 2188 3551
rect 2182 3546 2188 3547
rect 2346 3551 2352 3552
rect 2346 3547 2347 3551
rect 2351 3547 2352 3551
rect 2346 3546 2352 3547
rect 2474 3551 2480 3552
rect 2474 3547 2475 3551
rect 2479 3547 2480 3551
rect 2474 3546 2480 3547
rect 1974 3540 1980 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 2062 3540 2068 3541
rect 2062 3536 2063 3540
rect 2067 3536 2068 3540
rect 2062 3535 2068 3536
rect 2166 3540 2172 3541
rect 2166 3536 2167 3540
rect 2171 3536 2172 3540
rect 2166 3535 2172 3536
rect 2286 3540 2292 3541
rect 2286 3536 2287 3540
rect 2291 3536 2292 3540
rect 2286 3535 2292 3536
rect 2414 3540 2420 3541
rect 2414 3536 2415 3540
rect 2419 3536 2420 3540
rect 2414 3535 2420 3536
rect 2550 3540 2556 3541
rect 2550 3536 2551 3540
rect 2555 3536 2556 3540
rect 2550 3535 2556 3536
rect 2686 3540 2692 3541
rect 2686 3536 2687 3540
rect 2691 3536 2692 3540
rect 2686 3535 2692 3536
rect 1976 3519 1978 3535
rect 2064 3519 2066 3535
rect 2168 3519 2170 3535
rect 2288 3519 2290 3535
rect 2416 3519 2418 3535
rect 2552 3519 2554 3535
rect 2558 3523 2564 3524
rect 2558 3519 2559 3523
rect 2563 3519 2564 3523
rect 2688 3519 2690 3535
rect 1967 3518 1971 3519
rect 1967 3513 1971 3514
rect 1975 3518 1979 3519
rect 1975 3513 1979 3514
rect 2063 3518 2067 3519
rect 2063 3513 2067 3514
rect 2151 3518 2155 3519
rect 2151 3513 2155 3514
rect 2167 3518 2171 3519
rect 2167 3513 2171 3514
rect 2287 3518 2291 3519
rect 2287 3513 2291 3514
rect 2335 3518 2339 3519
rect 2335 3513 2339 3514
rect 2415 3518 2419 3519
rect 2415 3513 2419 3514
rect 2511 3518 2515 3519
rect 2511 3513 2515 3514
rect 2551 3518 2555 3519
rect 2558 3518 2564 3519
rect 2671 3518 2675 3519
rect 2551 3513 2555 3514
rect 1968 3497 1970 3513
rect 2152 3497 2154 3513
rect 2336 3497 2338 3513
rect 2512 3497 2514 3513
rect 1966 3496 1972 3497
rect 1966 3492 1967 3496
rect 1971 3492 1972 3496
rect 1966 3491 1972 3492
rect 2150 3496 2156 3497
rect 2150 3492 2151 3496
rect 2155 3492 2156 3496
rect 2150 3491 2156 3492
rect 2334 3496 2340 3497
rect 2334 3492 2335 3496
rect 2339 3492 2340 3496
rect 2334 3491 2340 3492
rect 2510 3496 2516 3497
rect 2510 3492 2511 3496
rect 2515 3492 2516 3496
rect 2510 3491 2516 3492
rect 1930 3487 1936 3488
rect 1930 3483 1931 3487
rect 1935 3483 1936 3487
rect 1015 3482 1019 3483
rect 1015 3477 1019 3478
rect 1039 3482 1043 3483
rect 1039 3477 1043 3478
rect 1103 3482 1107 3483
rect 1103 3477 1107 3478
rect 1135 3482 1139 3483
rect 1135 3477 1139 3478
rect 1191 3482 1195 3483
rect 1191 3477 1195 3478
rect 1231 3482 1235 3483
rect 1231 3477 1235 3478
rect 1279 3482 1283 3483
rect 1279 3477 1283 3478
rect 1327 3482 1331 3483
rect 1327 3477 1331 3478
rect 1367 3482 1371 3483
rect 1367 3477 1371 3478
rect 1455 3482 1459 3483
rect 1455 3477 1459 3478
rect 1831 3482 1835 3483
rect 1930 3482 1936 3483
rect 2034 3487 2040 3488
rect 2034 3483 2035 3487
rect 2039 3483 2040 3487
rect 2034 3482 2040 3483
rect 2402 3487 2408 3488
rect 2402 3483 2403 3487
rect 2407 3483 2408 3487
rect 2402 3482 2408 3483
rect 1831 3477 1835 3478
rect 986 3475 992 3476
rect 986 3471 987 3475
rect 991 3471 992 3475
rect 986 3470 992 3471
rect 994 3475 1000 3476
rect 994 3471 995 3475
rect 999 3471 1000 3475
rect 994 3470 1000 3471
rect 942 3466 948 3467
rect 942 3462 943 3466
rect 947 3462 948 3466
rect 942 3461 948 3462
rect 996 3440 998 3470
rect 1040 3467 1042 3477
rect 1090 3475 1096 3476
rect 1090 3471 1091 3475
rect 1095 3471 1096 3475
rect 1090 3470 1096 3471
rect 1038 3466 1044 3467
rect 1038 3462 1039 3466
rect 1043 3462 1044 3466
rect 1038 3461 1044 3462
rect 1092 3440 1094 3470
rect 1136 3467 1138 3477
rect 1206 3475 1212 3476
rect 1206 3471 1207 3475
rect 1211 3471 1212 3475
rect 1206 3470 1212 3471
rect 1134 3466 1140 3467
rect 1134 3462 1135 3466
rect 1139 3462 1140 3466
rect 1134 3461 1140 3462
rect 1208 3440 1210 3470
rect 1232 3467 1234 3477
rect 1328 3467 1330 3477
rect 1230 3466 1236 3467
rect 1230 3462 1231 3466
rect 1235 3462 1236 3466
rect 1230 3461 1236 3462
rect 1326 3466 1332 3467
rect 1326 3462 1327 3466
rect 1331 3462 1332 3466
rect 1326 3461 1332 3462
rect 1832 3449 1834 3477
rect 1870 3476 1876 3477
rect 1870 3472 1871 3476
rect 1875 3472 1876 3476
rect 1870 3471 1876 3472
rect 1830 3448 1836 3449
rect 1830 3444 1831 3448
rect 1835 3444 1836 3448
rect 1830 3443 1836 3444
rect 1872 3443 1874 3471
rect 1974 3458 1980 3459
rect 1974 3454 1975 3458
rect 1979 3454 1980 3458
rect 1974 3453 1980 3454
rect 1976 3443 1978 3453
rect 2036 3448 2038 3482
rect 2158 3458 2164 3459
rect 2158 3454 2159 3458
rect 2163 3454 2164 3458
rect 2158 3453 2164 3454
rect 2342 3458 2348 3459
rect 2342 3454 2343 3458
rect 2347 3454 2348 3458
rect 2342 3453 2348 3454
rect 2034 3447 2040 3448
rect 2034 3443 2035 3447
rect 2039 3443 2040 3447
rect 2160 3443 2162 3453
rect 2178 3447 2184 3448
rect 2178 3443 2179 3447
rect 2183 3443 2184 3447
rect 2344 3443 2346 3453
rect 2404 3448 2406 3482
rect 2518 3458 2524 3459
rect 2518 3454 2519 3458
rect 2523 3454 2524 3458
rect 2518 3453 2524 3454
rect 2402 3447 2408 3448
rect 2402 3443 2403 3447
rect 2407 3443 2408 3447
rect 2520 3443 2522 3453
rect 2560 3448 2562 3518
rect 2671 3513 2675 3514
rect 2687 3518 2691 3519
rect 2687 3513 2691 3514
rect 2672 3497 2674 3513
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2732 3480 2734 3578
rect 2748 3552 2750 3582
rect 2832 3579 2834 3589
rect 2976 3579 2978 3589
rect 3088 3588 3090 3634
rect 3590 3628 3596 3629
rect 3590 3624 3591 3628
rect 3595 3624 3596 3628
rect 3590 3623 3596 3624
rect 3270 3595 3276 3596
rect 3592 3595 3594 3623
rect 3119 3594 3123 3595
rect 3119 3589 3123 3590
rect 3263 3594 3267 3595
rect 3270 3591 3271 3595
rect 3275 3591 3276 3595
rect 3270 3590 3276 3591
rect 3591 3594 3595 3595
rect 3263 3589 3267 3590
rect 3086 3587 3092 3588
rect 3086 3583 3087 3587
rect 3091 3583 3092 3587
rect 3086 3582 3092 3583
rect 3120 3579 3122 3589
rect 3170 3587 3176 3588
rect 3170 3583 3171 3587
rect 3175 3583 3176 3587
rect 3170 3582 3176 3583
rect 2830 3578 2836 3579
rect 2830 3574 2831 3578
rect 2835 3574 2836 3578
rect 2830 3573 2836 3574
rect 2974 3578 2980 3579
rect 2974 3574 2975 3578
rect 2979 3574 2980 3578
rect 2974 3573 2980 3574
rect 3118 3578 3124 3579
rect 3118 3574 3119 3578
rect 3123 3574 3124 3578
rect 3118 3573 3124 3574
rect 2839 3572 2843 3573
rect 2839 3567 2843 3568
rect 2840 3552 2842 3567
rect 3172 3552 3174 3582
rect 3264 3579 3266 3589
rect 3262 3578 3268 3579
rect 3262 3574 3263 3578
rect 3267 3574 3268 3578
rect 3262 3573 3268 3574
rect 3272 3552 3274 3590
rect 3591 3589 3595 3590
rect 3592 3561 3594 3589
rect 3590 3560 3596 3561
rect 3590 3556 3591 3560
rect 3595 3556 3596 3560
rect 3590 3555 3596 3556
rect 2746 3551 2752 3552
rect 2746 3547 2747 3551
rect 2751 3547 2752 3551
rect 2746 3546 2752 3547
rect 2838 3551 2844 3552
rect 2838 3547 2839 3551
rect 2843 3547 2844 3551
rect 2838 3546 2844 3547
rect 3170 3551 3176 3552
rect 3170 3547 3171 3551
rect 3175 3547 3176 3551
rect 3170 3546 3176 3547
rect 3270 3551 3276 3552
rect 3270 3547 3271 3551
rect 3275 3547 3276 3551
rect 3270 3546 3276 3547
rect 3590 3543 3596 3544
rect 2822 3540 2828 3541
rect 2822 3536 2823 3540
rect 2827 3536 2828 3540
rect 2822 3535 2828 3536
rect 2966 3540 2972 3541
rect 2966 3536 2967 3540
rect 2971 3536 2972 3540
rect 2966 3535 2972 3536
rect 3110 3540 3116 3541
rect 3110 3536 3111 3540
rect 3115 3536 3116 3540
rect 3110 3535 3116 3536
rect 3254 3540 3260 3541
rect 3254 3536 3255 3540
rect 3259 3536 3260 3540
rect 3590 3539 3591 3543
rect 3595 3539 3596 3543
rect 3590 3538 3596 3539
rect 3254 3535 3260 3536
rect 2824 3519 2826 3535
rect 2968 3519 2970 3535
rect 2986 3523 2992 3524
rect 2986 3519 2987 3523
rect 2991 3519 2992 3523
rect 3112 3519 3114 3535
rect 3256 3519 3258 3535
rect 3592 3519 3594 3538
rect 2823 3518 2827 3519
rect 2823 3513 2827 3514
rect 2959 3518 2963 3519
rect 2959 3513 2963 3514
rect 2967 3518 2971 3519
rect 2986 3518 2992 3519
rect 3079 3518 3083 3519
rect 2967 3513 2971 3514
rect 2824 3497 2826 3513
rect 2960 3497 2962 3513
rect 2822 3496 2828 3497
rect 2822 3492 2823 3496
rect 2827 3492 2828 3496
rect 2822 3491 2828 3492
rect 2958 3496 2964 3497
rect 2958 3492 2959 3496
rect 2963 3492 2964 3496
rect 2958 3491 2964 3492
rect 2738 3487 2744 3488
rect 2738 3483 2739 3487
rect 2743 3483 2744 3487
rect 2738 3482 2744 3483
rect 2730 3479 2736 3480
rect 2730 3475 2731 3479
rect 2735 3475 2736 3479
rect 2730 3474 2736 3475
rect 2678 3458 2684 3459
rect 2678 3454 2679 3458
rect 2683 3454 2684 3458
rect 2678 3453 2684 3454
rect 2558 3447 2564 3448
rect 2558 3443 2559 3447
rect 2563 3443 2564 3447
rect 2680 3443 2682 3453
rect 2740 3448 2742 3482
rect 2830 3458 2836 3459
rect 2830 3454 2831 3458
rect 2835 3454 2836 3458
rect 2830 3453 2836 3454
rect 2966 3458 2972 3459
rect 2966 3454 2967 3458
rect 2971 3454 2972 3458
rect 2966 3453 2972 3454
rect 2738 3447 2744 3448
rect 2738 3443 2739 3447
rect 2743 3443 2744 3447
rect 2832 3443 2834 3453
rect 2854 3447 2860 3448
rect 2854 3443 2855 3447
rect 2859 3443 2860 3447
rect 2968 3443 2970 3453
rect 2988 3448 2990 3518
rect 3079 3513 3083 3514
rect 3111 3518 3115 3519
rect 3111 3513 3115 3514
rect 3191 3518 3195 3519
rect 3191 3513 3195 3514
rect 3255 3518 3259 3519
rect 3255 3513 3259 3514
rect 3303 3518 3307 3519
rect 3303 3513 3307 3514
rect 3415 3518 3419 3519
rect 3415 3513 3419 3514
rect 3503 3518 3507 3519
rect 3503 3513 3507 3514
rect 3591 3518 3595 3519
rect 3591 3513 3595 3514
rect 3080 3497 3082 3513
rect 3192 3497 3194 3513
rect 3304 3497 3306 3513
rect 3416 3497 3418 3513
rect 3504 3497 3506 3513
rect 3078 3496 3084 3497
rect 3078 3492 3079 3496
rect 3083 3492 3084 3496
rect 3078 3491 3084 3492
rect 3190 3496 3196 3497
rect 3190 3492 3191 3496
rect 3195 3492 3196 3496
rect 3190 3491 3196 3492
rect 3302 3496 3308 3497
rect 3302 3492 3303 3496
rect 3307 3492 3308 3496
rect 3302 3491 3308 3492
rect 3414 3496 3420 3497
rect 3414 3492 3415 3496
rect 3419 3492 3420 3496
rect 3414 3491 3420 3492
rect 3502 3496 3508 3497
rect 3502 3492 3503 3496
rect 3507 3492 3508 3496
rect 3592 3494 3594 3513
rect 3502 3491 3508 3492
rect 3590 3493 3596 3494
rect 3590 3489 3591 3493
rect 3595 3489 3596 3493
rect 3590 3488 3596 3489
rect 3042 3487 3048 3488
rect 3042 3483 3043 3487
rect 3047 3483 3048 3487
rect 3042 3482 3048 3483
rect 3158 3487 3164 3488
rect 3158 3483 3159 3487
rect 3163 3483 3164 3487
rect 3158 3482 3164 3483
rect 3270 3487 3276 3488
rect 3270 3483 3271 3487
rect 3275 3483 3276 3487
rect 3270 3482 3276 3483
rect 3382 3487 3388 3488
rect 3382 3483 3383 3487
rect 3387 3483 3388 3487
rect 3382 3482 3388 3483
rect 3482 3487 3488 3488
rect 3482 3483 3483 3487
rect 3487 3483 3488 3487
rect 3482 3482 3488 3483
rect 3044 3448 3046 3482
rect 3086 3458 3092 3459
rect 3086 3454 3087 3458
rect 3091 3454 3092 3458
rect 3086 3453 3092 3454
rect 2986 3447 2992 3448
rect 2986 3443 2987 3447
rect 2991 3443 2992 3447
rect 3042 3447 3048 3448
rect 3042 3443 3043 3447
rect 3047 3443 3048 3447
rect 3088 3443 3090 3453
rect 3160 3448 3162 3482
rect 3198 3458 3204 3459
rect 3198 3454 3199 3458
rect 3203 3454 3204 3458
rect 3198 3453 3204 3454
rect 3158 3447 3164 3448
rect 3158 3443 3159 3447
rect 3163 3443 3164 3447
rect 3200 3443 3202 3453
rect 3272 3448 3274 3482
rect 3310 3458 3316 3459
rect 3310 3454 3311 3458
rect 3315 3454 3316 3458
rect 3310 3453 3316 3454
rect 3270 3447 3276 3448
rect 3270 3443 3271 3447
rect 3275 3443 3276 3447
rect 3312 3443 3314 3453
rect 3384 3448 3386 3482
rect 3422 3458 3428 3459
rect 3422 3454 3423 3458
rect 3427 3454 3428 3458
rect 3422 3453 3428 3454
rect 3382 3447 3388 3448
rect 3382 3443 3383 3447
rect 3387 3443 3388 3447
rect 3424 3443 3426 3453
rect 3484 3448 3486 3482
rect 3562 3479 3568 3480
rect 3562 3475 3563 3479
rect 3567 3475 3568 3479
rect 3562 3474 3568 3475
rect 3590 3476 3596 3477
rect 3510 3458 3516 3459
rect 3510 3454 3511 3458
rect 3515 3454 3516 3458
rect 3510 3453 3516 3454
rect 3482 3447 3488 3448
rect 3482 3443 3483 3447
rect 3487 3443 3488 3447
rect 3512 3443 3514 3453
rect 1871 3442 1875 3443
rect 554 3439 560 3440
rect 554 3435 555 3439
rect 559 3435 560 3439
rect 554 3434 560 3435
rect 674 3439 680 3440
rect 674 3435 675 3439
rect 679 3435 680 3439
rect 674 3434 680 3435
rect 786 3439 792 3440
rect 786 3435 787 3439
rect 791 3435 792 3439
rect 786 3434 792 3435
rect 846 3439 852 3440
rect 846 3435 847 3439
rect 851 3435 852 3439
rect 846 3434 852 3435
rect 994 3439 1000 3440
rect 994 3435 995 3439
rect 999 3435 1000 3439
rect 994 3434 1000 3435
rect 1090 3439 1096 3440
rect 1090 3435 1091 3439
rect 1095 3435 1096 3439
rect 1090 3434 1096 3435
rect 1206 3439 1212 3440
rect 1206 3435 1207 3439
rect 1211 3435 1212 3439
rect 1871 3437 1875 3438
rect 1975 3442 1979 3443
rect 1975 3437 1979 3438
rect 2007 3442 2011 3443
rect 2034 3442 2040 3443
rect 2127 3442 2131 3443
rect 2007 3437 2011 3438
rect 2127 3437 2131 3438
rect 2159 3442 2163 3443
rect 2178 3442 2184 3443
rect 2255 3442 2259 3443
rect 2159 3437 2163 3438
rect 1206 3434 1212 3435
rect 1830 3431 1836 3432
rect 614 3428 620 3429
rect 614 3424 615 3428
rect 619 3424 620 3428
rect 614 3423 620 3424
rect 726 3428 732 3429
rect 726 3424 727 3428
rect 731 3424 732 3428
rect 726 3423 732 3424
rect 830 3428 836 3429
rect 830 3424 831 3428
rect 835 3424 836 3428
rect 830 3423 836 3424
rect 934 3428 940 3429
rect 934 3424 935 3428
rect 939 3424 940 3428
rect 934 3423 940 3424
rect 1030 3428 1036 3429
rect 1030 3424 1031 3428
rect 1035 3424 1036 3428
rect 1030 3423 1036 3424
rect 1126 3428 1132 3429
rect 1126 3424 1127 3428
rect 1131 3424 1132 3428
rect 1126 3423 1132 3424
rect 1222 3428 1228 3429
rect 1222 3424 1223 3428
rect 1227 3424 1228 3428
rect 1222 3423 1228 3424
rect 1318 3428 1324 3429
rect 1318 3424 1319 3428
rect 1323 3424 1324 3428
rect 1830 3427 1831 3431
rect 1835 3427 1836 3431
rect 1830 3426 1836 3427
rect 1318 3423 1324 3424
rect 616 3403 618 3423
rect 728 3403 730 3423
rect 832 3403 834 3423
rect 936 3403 938 3423
rect 1032 3403 1034 3423
rect 1128 3403 1130 3423
rect 1224 3403 1226 3423
rect 1246 3411 1252 3412
rect 1246 3407 1247 3411
rect 1251 3407 1252 3411
rect 1246 3406 1252 3407
rect 615 3402 619 3403
rect 615 3397 619 3398
rect 647 3402 651 3403
rect 647 3397 651 3398
rect 727 3402 731 3403
rect 727 3397 731 3398
rect 775 3402 779 3403
rect 775 3397 779 3398
rect 831 3402 835 3403
rect 831 3397 835 3398
rect 895 3402 899 3403
rect 895 3397 899 3398
rect 935 3402 939 3403
rect 935 3397 939 3398
rect 1015 3402 1019 3403
rect 1015 3397 1019 3398
rect 1031 3402 1035 3403
rect 1031 3397 1035 3398
rect 1127 3402 1131 3403
rect 1127 3397 1131 3398
rect 1223 3402 1227 3403
rect 1223 3397 1227 3398
rect 1239 3402 1243 3403
rect 1239 3397 1243 3398
rect 648 3381 650 3397
rect 776 3381 778 3397
rect 896 3381 898 3397
rect 1016 3381 1018 3397
rect 1128 3381 1130 3397
rect 1240 3381 1242 3397
rect 646 3380 652 3381
rect 646 3376 647 3380
rect 651 3376 652 3380
rect 646 3375 652 3376
rect 774 3380 780 3381
rect 774 3376 775 3380
rect 779 3376 780 3380
rect 774 3375 780 3376
rect 894 3380 900 3381
rect 894 3376 895 3380
rect 899 3376 900 3380
rect 894 3375 900 3376
rect 1014 3380 1020 3381
rect 1014 3376 1015 3380
rect 1019 3376 1020 3380
rect 1014 3375 1020 3376
rect 1126 3380 1132 3381
rect 1126 3376 1127 3380
rect 1131 3376 1132 3380
rect 1126 3375 1132 3376
rect 1238 3380 1244 3381
rect 1238 3376 1239 3380
rect 1243 3376 1244 3380
rect 1238 3375 1244 3376
rect 578 3371 584 3372
rect 282 3366 288 3367
rect 374 3367 380 3368
rect 284 3332 286 3366
rect 374 3363 375 3367
rect 379 3363 380 3367
rect 374 3362 380 3363
rect 518 3367 524 3368
rect 518 3363 519 3367
rect 523 3363 524 3367
rect 578 3367 579 3371
rect 583 3367 584 3371
rect 578 3366 584 3367
rect 714 3371 720 3372
rect 714 3367 715 3371
rect 719 3367 720 3371
rect 714 3366 720 3367
rect 1094 3371 1100 3372
rect 1094 3367 1095 3371
rect 1099 3367 1100 3371
rect 1094 3366 1100 3367
rect 1206 3371 1212 3372
rect 1206 3367 1207 3371
rect 1211 3367 1212 3371
rect 1206 3366 1212 3367
rect 518 3362 524 3363
rect 376 3347 378 3362
rect 376 3345 386 3347
rect 374 3342 380 3343
rect 374 3338 375 3342
rect 379 3338 380 3342
rect 374 3337 380 3338
rect 242 3331 248 3332
rect 242 3327 243 3331
rect 247 3327 248 3331
rect 242 3326 248 3327
rect 282 3331 288 3332
rect 282 3327 283 3331
rect 287 3327 288 3331
rect 282 3326 288 3327
rect 376 3323 378 3337
rect 111 3322 115 3323
rect 111 3317 115 3318
rect 207 3322 211 3323
rect 207 3317 211 3318
rect 223 3322 227 3323
rect 223 3317 227 3318
rect 367 3322 371 3323
rect 367 3317 371 3318
rect 375 3322 379 3323
rect 375 3317 379 3318
rect 112 3289 114 3317
rect 208 3307 210 3317
rect 298 3315 304 3316
rect 298 3311 299 3315
rect 303 3311 304 3315
rect 298 3310 304 3311
rect 206 3306 212 3307
rect 206 3302 207 3306
rect 211 3302 212 3306
rect 206 3301 212 3302
rect 110 3288 116 3289
rect 110 3284 111 3288
rect 115 3284 116 3288
rect 110 3283 116 3284
rect 300 3280 302 3310
rect 368 3307 370 3317
rect 384 3316 386 3345
rect 518 3342 524 3343
rect 518 3338 519 3342
rect 523 3338 524 3342
rect 518 3337 524 3338
rect 520 3323 522 3337
rect 580 3332 582 3366
rect 654 3342 660 3343
rect 654 3338 655 3342
rect 659 3338 660 3342
rect 654 3337 660 3338
rect 578 3331 584 3332
rect 578 3327 579 3331
rect 583 3327 584 3331
rect 578 3326 584 3327
rect 656 3323 658 3337
rect 716 3332 718 3366
rect 927 3356 931 3357
rect 927 3351 931 3352
rect 782 3342 788 3343
rect 782 3338 783 3342
rect 787 3338 788 3342
rect 782 3337 788 3338
rect 902 3342 908 3343
rect 902 3338 903 3342
rect 907 3338 908 3342
rect 902 3337 908 3338
rect 714 3331 720 3332
rect 714 3327 715 3331
rect 719 3327 720 3331
rect 714 3326 720 3327
rect 784 3323 786 3337
rect 822 3331 828 3332
rect 822 3327 823 3331
rect 827 3327 828 3331
rect 822 3326 828 3327
rect 519 3322 523 3323
rect 519 3317 523 3318
rect 655 3322 659 3323
rect 655 3317 659 3318
rect 671 3322 675 3323
rect 671 3317 675 3318
rect 783 3322 787 3323
rect 783 3317 787 3318
rect 815 3322 819 3323
rect 815 3317 819 3318
rect 382 3315 388 3316
rect 382 3311 383 3315
rect 387 3311 388 3315
rect 382 3310 388 3311
rect 520 3307 522 3317
rect 546 3315 552 3316
rect 546 3311 547 3315
rect 551 3311 552 3315
rect 546 3310 552 3311
rect 570 3315 576 3316
rect 570 3311 571 3315
rect 575 3311 576 3315
rect 570 3310 576 3311
rect 366 3306 372 3307
rect 366 3302 367 3306
rect 371 3302 372 3306
rect 366 3301 372 3302
rect 518 3306 524 3307
rect 518 3302 519 3306
rect 523 3302 524 3306
rect 518 3301 524 3302
rect 258 3279 264 3280
rect 258 3275 259 3279
rect 263 3275 264 3279
rect 258 3274 264 3275
rect 298 3279 304 3280
rect 298 3275 299 3279
rect 303 3275 304 3279
rect 298 3274 304 3275
rect 110 3271 116 3272
rect 110 3267 111 3271
rect 115 3267 116 3271
rect 110 3266 116 3267
rect 198 3268 204 3269
rect 112 3247 114 3266
rect 198 3264 199 3268
rect 203 3264 204 3268
rect 198 3263 204 3264
rect 200 3247 202 3263
rect 111 3246 115 3247
rect 111 3241 115 3242
rect 135 3246 139 3247
rect 135 3241 139 3242
rect 199 3246 203 3247
rect 199 3241 203 3242
rect 112 3222 114 3241
rect 136 3225 138 3241
rect 134 3224 140 3225
rect 110 3221 116 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 134 3220 135 3224
rect 139 3220 140 3224
rect 134 3219 140 3220
rect 110 3216 116 3217
rect 202 3215 208 3216
rect 202 3211 203 3215
rect 207 3211 208 3215
rect 202 3210 208 3211
rect 194 3207 200 3208
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 194 3203 195 3207
rect 199 3203 200 3207
rect 194 3202 200 3203
rect 110 3199 116 3200
rect 112 3163 114 3199
rect 142 3186 148 3187
rect 142 3182 143 3186
rect 147 3182 148 3186
rect 142 3181 148 3182
rect 144 3163 146 3181
rect 196 3176 198 3202
rect 194 3175 200 3176
rect 194 3171 195 3175
rect 199 3171 200 3175
rect 194 3170 200 3171
rect 111 3162 115 3163
rect 111 3157 115 3158
rect 143 3162 147 3163
rect 143 3157 147 3158
rect 175 3162 179 3163
rect 175 3157 179 3158
rect 112 3129 114 3157
rect 176 3147 178 3157
rect 204 3156 206 3210
rect 260 3176 262 3274
rect 358 3268 364 3269
rect 358 3264 359 3268
rect 363 3264 364 3268
rect 358 3263 364 3264
rect 510 3268 516 3269
rect 510 3264 511 3268
rect 515 3264 516 3268
rect 510 3263 516 3264
rect 360 3247 362 3263
rect 512 3247 514 3263
rect 271 3246 275 3247
rect 271 3241 275 3242
rect 359 3246 363 3247
rect 359 3241 363 3242
rect 415 3246 419 3247
rect 415 3241 419 3242
rect 511 3246 515 3247
rect 511 3241 515 3242
rect 272 3225 274 3241
rect 416 3225 418 3241
rect 270 3224 276 3225
rect 270 3220 271 3224
rect 275 3220 276 3224
rect 270 3219 276 3220
rect 414 3224 420 3225
rect 414 3220 415 3224
rect 419 3220 420 3224
rect 414 3219 420 3220
rect 548 3216 550 3310
rect 572 3280 574 3310
rect 672 3307 674 3317
rect 722 3315 728 3316
rect 722 3311 723 3315
rect 727 3311 728 3315
rect 722 3310 728 3311
rect 670 3306 676 3307
rect 670 3302 671 3306
rect 675 3302 676 3306
rect 670 3301 676 3302
rect 724 3280 726 3310
rect 816 3307 818 3317
rect 814 3306 820 3307
rect 814 3302 815 3306
rect 819 3302 820 3306
rect 814 3301 820 3302
rect 824 3280 826 3326
rect 904 3323 906 3337
rect 928 3332 930 3351
rect 1022 3342 1028 3343
rect 979 3340 983 3341
rect 1022 3338 1023 3342
rect 1027 3338 1028 3342
rect 1022 3337 1028 3338
rect 979 3335 983 3336
rect 926 3331 932 3332
rect 926 3327 927 3331
rect 931 3327 932 3331
rect 926 3326 932 3327
rect 903 3322 907 3323
rect 903 3317 907 3318
rect 951 3322 955 3323
rect 951 3317 955 3318
rect 952 3307 954 3317
rect 980 3316 982 3335
rect 1024 3323 1026 3337
rect 1096 3332 1098 3366
rect 1134 3342 1140 3343
rect 1134 3338 1135 3342
rect 1139 3338 1140 3342
rect 1134 3337 1140 3338
rect 1094 3331 1100 3332
rect 1094 3327 1095 3331
rect 1099 3327 1100 3331
rect 1094 3326 1100 3327
rect 1136 3323 1138 3337
rect 1208 3332 1210 3366
rect 1248 3357 1250 3406
rect 1320 3403 1322 3423
rect 1832 3403 1834 3426
rect 1872 3409 1874 3437
rect 2008 3427 2010 3437
rect 2058 3435 2064 3436
rect 2058 3431 2059 3435
rect 2063 3431 2064 3435
rect 2058 3430 2064 3431
rect 2006 3426 2012 3427
rect 2006 3422 2007 3426
rect 2011 3422 2012 3426
rect 2006 3421 2012 3422
rect 1870 3408 1876 3409
rect 1870 3404 1871 3408
rect 1875 3404 1876 3408
rect 1870 3403 1876 3404
rect 1319 3402 1323 3403
rect 1319 3397 1323 3398
rect 1351 3402 1355 3403
rect 1351 3397 1355 3398
rect 1831 3402 1835 3403
rect 2060 3400 2062 3430
rect 2128 3427 2130 3437
rect 2126 3426 2132 3427
rect 2126 3422 2127 3426
rect 2131 3422 2132 3426
rect 2126 3421 2132 3422
rect 2180 3400 2182 3442
rect 2343 3442 2347 3443
rect 2255 3437 2259 3438
rect 2262 3439 2268 3440
rect 2256 3427 2258 3437
rect 2262 3435 2263 3439
rect 2267 3435 2268 3439
rect 2343 3437 2347 3438
rect 2391 3442 2395 3443
rect 2402 3442 2408 3443
rect 2519 3442 2523 3443
rect 2391 3437 2395 3438
rect 2519 3437 2523 3438
rect 2535 3442 2539 3443
rect 2558 3442 2564 3443
rect 2679 3442 2683 3443
rect 2738 3442 2744 3443
rect 2831 3442 2835 3443
rect 2854 3442 2860 3443
rect 2967 3442 2971 3443
rect 2986 3442 2992 3443
rect 2999 3442 3003 3443
rect 3042 3442 3048 3443
rect 3087 3442 3091 3443
rect 3158 3442 3164 3443
rect 3167 3442 3171 3443
rect 2535 3437 2539 3438
rect 2679 3437 2683 3438
rect 2831 3437 2835 3438
rect 2262 3434 2268 3435
rect 2282 3435 2288 3436
rect 2254 3426 2260 3427
rect 2254 3422 2255 3426
rect 2259 3422 2260 3426
rect 2254 3421 2260 3422
rect 2264 3400 2266 3434
rect 2282 3431 2283 3435
rect 2287 3431 2288 3435
rect 2282 3430 2288 3431
rect 1831 3397 1835 3398
rect 2058 3399 2064 3400
rect 1352 3381 1354 3397
rect 1350 3380 1356 3381
rect 1350 3376 1351 3380
rect 1355 3376 1356 3380
rect 1832 3378 1834 3397
rect 2058 3395 2059 3399
rect 2063 3395 2064 3399
rect 2058 3394 2064 3395
rect 2178 3399 2184 3400
rect 2178 3395 2179 3399
rect 2183 3395 2184 3399
rect 2178 3394 2184 3395
rect 2262 3399 2268 3400
rect 2262 3395 2263 3399
rect 2267 3395 2268 3399
rect 2262 3394 2268 3395
rect 1870 3391 1876 3392
rect 1870 3387 1871 3391
rect 1875 3387 1876 3391
rect 1870 3386 1876 3387
rect 1998 3388 2004 3389
rect 1350 3375 1356 3376
rect 1830 3377 1836 3378
rect 1830 3373 1831 3377
rect 1835 3373 1836 3377
rect 1830 3372 1836 3373
rect 1318 3371 1324 3372
rect 1318 3367 1319 3371
rect 1323 3367 1324 3371
rect 1318 3366 1324 3367
rect 1326 3371 1332 3372
rect 1326 3367 1327 3371
rect 1331 3367 1332 3371
rect 1872 3367 1874 3386
rect 1998 3384 1999 3388
rect 2003 3384 2004 3388
rect 1998 3383 2004 3384
rect 2118 3388 2124 3389
rect 2118 3384 2119 3388
rect 2123 3384 2124 3388
rect 2118 3383 2124 3384
rect 2246 3388 2252 3389
rect 2246 3384 2247 3388
rect 2251 3384 2252 3388
rect 2246 3383 2252 3384
rect 2000 3367 2002 3383
rect 2120 3367 2122 3383
rect 2248 3367 2250 3383
rect 1326 3366 1332 3367
rect 1871 3366 1875 3367
rect 1247 3356 1251 3357
rect 1247 3351 1251 3352
rect 1246 3342 1252 3343
rect 1246 3338 1247 3342
rect 1251 3338 1252 3342
rect 1246 3337 1252 3338
rect 1206 3331 1212 3332
rect 1206 3327 1207 3331
rect 1211 3327 1212 3331
rect 1206 3326 1212 3327
rect 1248 3323 1250 3337
rect 1320 3332 1322 3366
rect 1328 3341 1330 3366
rect 1871 3361 1875 3362
rect 1999 3366 2003 3367
rect 1999 3361 2003 3362
rect 2015 3366 2019 3367
rect 2015 3361 2019 3362
rect 2119 3366 2123 3367
rect 2119 3361 2123 3362
rect 2151 3366 2155 3367
rect 2151 3361 2155 3362
rect 2247 3366 2251 3367
rect 2247 3361 2251 3362
rect 1830 3360 1836 3361
rect 1830 3356 1831 3360
rect 1835 3356 1836 3360
rect 1830 3355 1836 3356
rect 1358 3342 1364 3343
rect 1327 3340 1331 3341
rect 1358 3338 1359 3342
rect 1363 3338 1364 3342
rect 1358 3337 1364 3338
rect 1327 3335 1331 3336
rect 1318 3331 1324 3332
rect 1318 3327 1319 3331
rect 1323 3327 1324 3331
rect 1318 3326 1324 3327
rect 1360 3323 1362 3337
rect 1832 3323 1834 3355
rect 1872 3342 1874 3361
rect 2016 3345 2018 3361
rect 2152 3345 2154 3361
rect 2014 3344 2020 3345
rect 1870 3341 1876 3342
rect 1870 3337 1871 3341
rect 1875 3337 1876 3341
rect 2014 3340 2015 3344
rect 2019 3340 2020 3344
rect 2014 3339 2020 3340
rect 2150 3344 2156 3345
rect 2150 3340 2151 3344
rect 2155 3340 2156 3344
rect 2150 3339 2156 3340
rect 1870 3336 1876 3337
rect 2284 3336 2286 3430
rect 2392 3427 2394 3437
rect 2442 3435 2448 3436
rect 2442 3431 2443 3435
rect 2447 3431 2448 3435
rect 2442 3430 2448 3431
rect 2390 3426 2396 3427
rect 2390 3422 2391 3426
rect 2395 3422 2396 3426
rect 2390 3421 2396 3422
rect 2444 3400 2446 3430
rect 2536 3427 2538 3437
rect 2586 3435 2592 3436
rect 2586 3431 2587 3435
rect 2591 3431 2592 3435
rect 2586 3430 2592 3431
rect 2534 3426 2540 3427
rect 2534 3422 2535 3426
rect 2539 3422 2540 3426
rect 2534 3421 2540 3422
rect 2588 3400 2590 3430
rect 2680 3427 2682 3437
rect 2832 3427 2834 3437
rect 2678 3426 2684 3427
rect 2678 3422 2679 3426
rect 2683 3422 2684 3426
rect 2678 3421 2684 3422
rect 2830 3426 2836 3427
rect 2830 3422 2831 3426
rect 2835 3422 2836 3426
rect 2830 3421 2836 3422
rect 2856 3400 2858 3442
rect 2967 3437 2971 3438
rect 2999 3437 3003 3438
rect 3087 3437 3091 3438
rect 3167 3437 3171 3438
rect 3199 3442 3203 3443
rect 3270 3442 3276 3443
rect 3311 3442 3315 3443
rect 3199 3437 3203 3438
rect 3311 3437 3315 3438
rect 3343 3442 3347 3443
rect 3382 3442 3388 3443
rect 3423 3442 3427 3443
rect 3482 3442 3488 3443
rect 3511 3442 3515 3443
rect 3343 3437 3347 3438
rect 3423 3437 3427 3438
rect 3511 3437 3515 3438
rect 3000 3427 3002 3437
rect 3006 3435 3012 3436
rect 3006 3431 3007 3435
rect 3011 3431 3012 3435
rect 3006 3430 3012 3431
rect 2998 3426 3004 3427
rect 2998 3422 2999 3426
rect 3003 3422 3004 3426
rect 2998 3421 3004 3422
rect 3008 3400 3010 3430
rect 3168 3427 3170 3437
rect 3174 3435 3180 3436
rect 3174 3431 3175 3435
rect 3179 3431 3180 3435
rect 3174 3430 3180 3431
rect 3166 3426 3172 3427
rect 3166 3422 3167 3426
rect 3171 3422 3172 3426
rect 3166 3421 3172 3422
rect 3176 3400 3178 3430
rect 3344 3427 3346 3437
rect 3350 3435 3356 3436
rect 3350 3431 3351 3435
rect 3355 3431 3356 3435
rect 3350 3430 3356 3431
rect 3358 3435 3364 3436
rect 3358 3431 3359 3435
rect 3363 3431 3364 3435
rect 3358 3430 3364 3431
rect 3342 3426 3348 3427
rect 3342 3422 3343 3426
rect 3347 3422 3348 3426
rect 3342 3421 3348 3422
rect 3352 3400 3354 3430
rect 2442 3399 2448 3400
rect 2442 3395 2443 3399
rect 2447 3395 2448 3399
rect 2442 3394 2448 3395
rect 2586 3399 2592 3400
rect 2586 3395 2587 3399
rect 2591 3395 2592 3399
rect 2586 3394 2592 3395
rect 2854 3399 2860 3400
rect 2854 3395 2855 3399
rect 2859 3395 2860 3399
rect 2854 3394 2860 3395
rect 3006 3399 3012 3400
rect 3006 3395 3007 3399
rect 3011 3395 3012 3399
rect 3006 3394 3012 3395
rect 3174 3399 3180 3400
rect 3174 3395 3175 3399
rect 3179 3395 3180 3399
rect 3174 3394 3180 3395
rect 3350 3399 3356 3400
rect 3350 3395 3351 3399
rect 3355 3395 3356 3399
rect 3350 3394 3356 3395
rect 2382 3388 2388 3389
rect 2382 3384 2383 3388
rect 2387 3384 2388 3388
rect 2382 3383 2388 3384
rect 2526 3388 2532 3389
rect 2526 3384 2527 3388
rect 2531 3384 2532 3388
rect 2526 3383 2532 3384
rect 2670 3388 2676 3389
rect 2670 3384 2671 3388
rect 2675 3384 2676 3388
rect 2670 3383 2676 3384
rect 2822 3388 2828 3389
rect 2822 3384 2823 3388
rect 2827 3384 2828 3388
rect 2822 3383 2828 3384
rect 2990 3388 2996 3389
rect 2990 3384 2991 3388
rect 2995 3384 2996 3388
rect 2990 3383 2996 3384
rect 3158 3388 3164 3389
rect 3158 3384 3159 3388
rect 3163 3384 3164 3388
rect 3158 3383 3164 3384
rect 3334 3388 3340 3389
rect 3334 3384 3335 3388
rect 3339 3384 3340 3388
rect 3334 3383 3340 3384
rect 2384 3367 2386 3383
rect 2528 3367 2530 3383
rect 2618 3371 2624 3372
rect 2618 3367 2619 3371
rect 2623 3367 2624 3371
rect 2672 3367 2674 3383
rect 2824 3367 2826 3383
rect 2992 3367 2994 3383
rect 3160 3367 3162 3383
rect 3336 3367 3338 3383
rect 2295 3366 2299 3367
rect 2295 3361 2299 3362
rect 2383 3366 2387 3367
rect 2383 3361 2387 3362
rect 2439 3366 2443 3367
rect 2439 3361 2443 3362
rect 2527 3366 2531 3367
rect 2527 3361 2531 3362
rect 2583 3366 2587 3367
rect 2618 3366 2624 3367
rect 2671 3366 2675 3367
rect 2583 3361 2587 3362
rect 2296 3345 2298 3361
rect 2440 3345 2442 3361
rect 2584 3345 2586 3361
rect 2294 3344 2300 3345
rect 2294 3340 2295 3344
rect 2299 3340 2300 3344
rect 2294 3339 2300 3340
rect 2438 3344 2444 3345
rect 2438 3340 2439 3344
rect 2443 3340 2444 3344
rect 2438 3339 2444 3340
rect 2582 3344 2588 3345
rect 2582 3340 2583 3344
rect 2587 3340 2588 3344
rect 2582 3339 2588 3340
rect 2106 3335 2112 3336
rect 2106 3331 2107 3335
rect 2111 3331 2112 3335
rect 2106 3330 2112 3331
rect 2246 3335 2252 3336
rect 2246 3331 2247 3335
rect 2251 3331 2252 3335
rect 2246 3330 2252 3331
rect 2282 3335 2288 3336
rect 2282 3331 2283 3335
rect 2287 3331 2288 3335
rect 2282 3330 2288 3331
rect 2506 3335 2512 3336
rect 2506 3331 2507 3335
rect 2511 3331 2512 3335
rect 2506 3330 2512 3331
rect 1870 3324 1876 3325
rect 1023 3322 1027 3323
rect 1023 3317 1027 3318
rect 1087 3322 1091 3323
rect 1087 3317 1091 3318
rect 1135 3322 1139 3323
rect 1135 3317 1139 3318
rect 1215 3322 1219 3323
rect 1215 3317 1219 3318
rect 1247 3322 1251 3323
rect 1247 3317 1251 3318
rect 1343 3322 1347 3323
rect 1343 3317 1347 3318
rect 1359 3322 1363 3323
rect 1359 3317 1363 3318
rect 1471 3322 1475 3323
rect 1471 3317 1475 3318
rect 1831 3322 1835 3323
rect 1870 3320 1871 3324
rect 1875 3320 1876 3324
rect 1870 3319 1876 3320
rect 1831 3317 1835 3318
rect 978 3315 984 3316
rect 978 3311 979 3315
rect 983 3311 984 3315
rect 978 3310 984 3311
rect 1002 3315 1008 3316
rect 1002 3311 1003 3315
rect 1007 3311 1008 3315
rect 1002 3310 1008 3311
rect 950 3306 956 3307
rect 950 3302 951 3306
rect 955 3302 956 3306
rect 950 3301 956 3302
rect 1004 3280 1006 3310
rect 1088 3307 1090 3317
rect 1166 3315 1172 3316
rect 1166 3311 1167 3315
rect 1171 3311 1172 3315
rect 1166 3310 1172 3311
rect 1086 3306 1092 3307
rect 1086 3302 1087 3306
rect 1091 3302 1092 3306
rect 1086 3301 1092 3302
rect 1168 3280 1170 3310
rect 1216 3307 1218 3317
rect 1266 3315 1272 3316
rect 1266 3311 1267 3315
rect 1271 3311 1272 3315
rect 1266 3310 1272 3311
rect 1214 3306 1220 3307
rect 1214 3302 1215 3306
rect 1219 3302 1220 3306
rect 1214 3301 1220 3302
rect 1268 3280 1270 3310
rect 1344 3307 1346 3317
rect 1394 3315 1400 3316
rect 1394 3311 1395 3315
rect 1399 3311 1400 3315
rect 1394 3310 1400 3311
rect 1342 3306 1348 3307
rect 1342 3302 1343 3306
rect 1347 3302 1348 3306
rect 1342 3301 1348 3302
rect 1396 3280 1398 3310
rect 1472 3307 1474 3317
rect 1470 3306 1476 3307
rect 1470 3302 1471 3306
rect 1475 3302 1476 3306
rect 1470 3301 1476 3302
rect 1832 3289 1834 3317
rect 1872 3291 1874 3319
rect 2022 3306 2028 3307
rect 2022 3302 2023 3306
rect 2027 3302 2028 3306
rect 2022 3301 2028 3302
rect 1978 3295 1984 3296
rect 1978 3291 1979 3295
rect 1983 3291 1984 3295
rect 2024 3291 2026 3301
rect 2108 3296 2110 3330
rect 2158 3306 2164 3307
rect 2158 3302 2159 3306
rect 2163 3302 2164 3306
rect 2158 3301 2164 3302
rect 2106 3295 2112 3296
rect 2106 3291 2107 3295
rect 2111 3291 2112 3295
rect 2160 3291 2162 3301
rect 2248 3296 2250 3330
rect 2498 3327 2504 3328
rect 2498 3323 2499 3327
rect 2503 3323 2504 3327
rect 2498 3322 2504 3323
rect 2302 3306 2308 3307
rect 2302 3302 2303 3306
rect 2307 3302 2308 3306
rect 2302 3301 2308 3302
rect 2446 3306 2452 3307
rect 2446 3302 2447 3306
rect 2451 3302 2452 3306
rect 2446 3301 2452 3302
rect 2246 3295 2252 3296
rect 2246 3291 2247 3295
rect 2251 3291 2252 3295
rect 2304 3291 2306 3301
rect 2448 3291 2450 3301
rect 1871 3290 1875 3291
rect 1830 3288 1836 3289
rect 1830 3284 1831 3288
rect 1835 3284 1836 3288
rect 1871 3285 1875 3286
rect 1927 3290 1931 3291
rect 1978 3290 1984 3291
rect 2023 3290 2027 3291
rect 1927 3285 1931 3286
rect 1830 3283 1836 3284
rect 570 3279 576 3280
rect 570 3275 571 3279
rect 575 3275 576 3279
rect 570 3274 576 3275
rect 722 3279 728 3280
rect 722 3275 723 3279
rect 727 3275 728 3279
rect 722 3274 728 3275
rect 822 3279 828 3280
rect 822 3275 823 3279
rect 827 3275 828 3279
rect 822 3274 828 3275
rect 1002 3279 1008 3280
rect 1002 3275 1003 3279
rect 1007 3275 1008 3279
rect 1002 3274 1008 3275
rect 1166 3279 1172 3280
rect 1166 3275 1167 3279
rect 1171 3275 1172 3279
rect 1166 3274 1172 3275
rect 1266 3279 1272 3280
rect 1266 3275 1267 3279
rect 1271 3275 1272 3279
rect 1266 3274 1272 3275
rect 1394 3279 1400 3280
rect 1394 3275 1395 3279
rect 1399 3275 1400 3279
rect 1394 3274 1400 3275
rect 1830 3271 1836 3272
rect 662 3268 668 3269
rect 662 3264 663 3268
rect 667 3264 668 3268
rect 662 3263 668 3264
rect 806 3268 812 3269
rect 806 3264 807 3268
rect 811 3264 812 3268
rect 806 3263 812 3264
rect 942 3268 948 3269
rect 942 3264 943 3268
rect 947 3264 948 3268
rect 942 3263 948 3264
rect 1078 3268 1084 3269
rect 1078 3264 1079 3268
rect 1083 3264 1084 3268
rect 1078 3263 1084 3264
rect 1206 3268 1212 3269
rect 1206 3264 1207 3268
rect 1211 3264 1212 3268
rect 1206 3263 1212 3264
rect 1334 3268 1340 3269
rect 1334 3264 1335 3268
rect 1339 3264 1340 3268
rect 1334 3263 1340 3264
rect 1462 3268 1468 3269
rect 1462 3264 1463 3268
rect 1467 3264 1468 3268
rect 1830 3267 1831 3271
rect 1835 3267 1836 3271
rect 1830 3266 1836 3267
rect 1462 3263 1468 3264
rect 664 3247 666 3263
rect 808 3247 810 3263
rect 944 3247 946 3263
rect 1080 3247 1082 3263
rect 1208 3247 1210 3263
rect 1336 3247 1338 3263
rect 1398 3251 1404 3252
rect 1398 3247 1399 3251
rect 1403 3247 1404 3251
rect 1464 3247 1466 3263
rect 1832 3247 1834 3266
rect 1872 3257 1874 3285
rect 1928 3275 1930 3285
rect 1926 3274 1932 3275
rect 1926 3270 1927 3274
rect 1931 3270 1932 3274
rect 1926 3269 1932 3270
rect 1870 3256 1876 3257
rect 1870 3252 1871 3256
rect 1875 3252 1876 3256
rect 1870 3251 1876 3252
rect 1980 3248 1982 3290
rect 2023 3285 2027 3286
rect 2063 3290 2067 3291
rect 2106 3290 2112 3291
rect 2159 3290 2163 3291
rect 2063 3285 2067 3286
rect 2159 3285 2163 3286
rect 2191 3290 2195 3291
rect 2246 3290 2252 3291
rect 2303 3290 2307 3291
rect 2191 3285 2195 3286
rect 2303 3285 2307 3286
rect 2319 3290 2323 3291
rect 2319 3285 2323 3286
rect 2447 3290 2451 3291
rect 2447 3285 2451 3286
rect 2064 3275 2066 3285
rect 2070 3283 2076 3284
rect 2070 3279 2071 3283
rect 2075 3279 2076 3283
rect 2070 3278 2076 3279
rect 2062 3274 2068 3275
rect 2062 3270 2063 3274
rect 2067 3270 2068 3274
rect 2062 3269 2068 3270
rect 2072 3248 2074 3278
rect 2192 3275 2194 3285
rect 2198 3283 2204 3284
rect 2198 3279 2199 3283
rect 2203 3279 2204 3283
rect 2198 3278 2204 3279
rect 2210 3283 2216 3284
rect 2210 3279 2211 3283
rect 2215 3279 2216 3283
rect 2210 3278 2216 3279
rect 2190 3274 2196 3275
rect 2190 3270 2191 3274
rect 2195 3270 2196 3274
rect 2190 3269 2196 3270
rect 2200 3248 2202 3278
rect 1978 3247 1984 3248
rect 575 3246 579 3247
rect 575 3241 579 3242
rect 663 3246 667 3247
rect 663 3241 667 3242
rect 735 3246 739 3247
rect 735 3241 739 3242
rect 807 3246 811 3247
rect 807 3241 811 3242
rect 895 3246 899 3247
rect 895 3241 899 3242
rect 943 3246 947 3247
rect 943 3241 947 3242
rect 1047 3246 1051 3247
rect 1047 3241 1051 3242
rect 1079 3246 1083 3247
rect 1079 3241 1083 3242
rect 1191 3246 1195 3247
rect 1191 3241 1195 3242
rect 1207 3246 1211 3247
rect 1207 3241 1211 3242
rect 1327 3246 1331 3247
rect 1327 3241 1331 3242
rect 1335 3246 1339 3247
rect 1398 3246 1404 3247
rect 1463 3246 1467 3247
rect 1335 3241 1339 3242
rect 576 3225 578 3241
rect 736 3225 738 3241
rect 896 3225 898 3241
rect 1048 3225 1050 3241
rect 1192 3225 1194 3241
rect 1328 3225 1330 3241
rect 574 3224 580 3225
rect 574 3220 575 3224
rect 579 3220 580 3224
rect 574 3219 580 3220
rect 734 3224 740 3225
rect 734 3220 735 3224
rect 739 3220 740 3224
rect 734 3219 740 3220
rect 894 3224 900 3225
rect 894 3220 895 3224
rect 899 3220 900 3224
rect 894 3219 900 3220
rect 1046 3224 1052 3225
rect 1046 3220 1047 3224
rect 1051 3220 1052 3224
rect 1046 3219 1052 3220
rect 1190 3224 1196 3225
rect 1190 3220 1191 3224
rect 1195 3220 1196 3224
rect 1190 3219 1196 3220
rect 1326 3224 1332 3225
rect 1326 3220 1327 3224
rect 1331 3220 1332 3224
rect 1326 3219 1332 3220
rect 546 3215 552 3216
rect 546 3211 547 3215
rect 551 3211 552 3215
rect 546 3210 552 3211
rect 642 3215 648 3216
rect 642 3211 643 3215
rect 647 3211 648 3215
rect 642 3210 648 3211
rect 802 3215 808 3216
rect 802 3211 803 3215
rect 807 3211 808 3215
rect 802 3210 808 3211
rect 1114 3215 1120 3216
rect 1114 3211 1115 3215
rect 1119 3211 1120 3215
rect 1114 3210 1120 3211
rect 1282 3215 1288 3216
rect 1282 3211 1283 3215
rect 1287 3211 1288 3215
rect 1282 3210 1288 3211
rect 278 3186 284 3187
rect 278 3182 279 3186
rect 283 3182 284 3186
rect 278 3181 284 3182
rect 422 3186 428 3187
rect 422 3182 423 3186
rect 427 3182 428 3186
rect 422 3181 428 3182
rect 582 3186 588 3187
rect 582 3182 583 3186
rect 587 3182 588 3186
rect 582 3181 588 3182
rect 258 3175 264 3176
rect 258 3171 259 3175
rect 263 3171 264 3175
rect 258 3170 264 3171
rect 280 3163 282 3181
rect 424 3163 426 3181
rect 584 3163 586 3181
rect 644 3176 646 3210
rect 742 3186 748 3187
rect 742 3182 743 3186
rect 747 3182 748 3186
rect 742 3181 748 3182
rect 642 3175 648 3176
rect 642 3171 643 3175
rect 647 3171 648 3175
rect 642 3170 648 3171
rect 744 3163 746 3181
rect 804 3176 806 3210
rect 902 3186 908 3187
rect 902 3182 903 3186
rect 907 3182 908 3186
rect 902 3181 908 3182
rect 1054 3186 1060 3187
rect 1054 3182 1055 3186
rect 1059 3182 1060 3186
rect 1054 3181 1060 3182
rect 802 3175 808 3176
rect 802 3171 803 3175
rect 807 3171 808 3175
rect 802 3170 808 3171
rect 904 3163 906 3181
rect 911 3172 915 3173
rect 911 3167 915 3168
rect 279 3162 283 3163
rect 279 3157 283 3158
rect 319 3162 323 3163
rect 319 3157 323 3158
rect 423 3162 427 3163
rect 423 3157 427 3158
rect 463 3162 467 3163
rect 463 3157 467 3158
rect 583 3162 587 3163
rect 583 3157 587 3158
rect 607 3162 611 3163
rect 607 3157 611 3158
rect 743 3162 747 3163
rect 743 3157 747 3158
rect 871 3162 875 3163
rect 871 3157 875 3158
rect 903 3162 907 3163
rect 903 3157 907 3158
rect 202 3155 208 3156
rect 202 3151 203 3155
rect 207 3151 208 3155
rect 202 3150 208 3151
rect 226 3155 232 3156
rect 226 3151 227 3155
rect 231 3151 232 3155
rect 226 3150 232 3151
rect 174 3146 180 3147
rect 174 3142 175 3146
rect 179 3142 180 3146
rect 174 3141 180 3142
rect 110 3128 116 3129
rect 110 3124 111 3128
rect 115 3124 116 3128
rect 110 3123 116 3124
rect 228 3120 230 3150
rect 320 3147 322 3157
rect 464 3147 466 3157
rect 498 3155 504 3156
rect 498 3151 499 3155
rect 503 3151 504 3155
rect 498 3150 504 3151
rect 514 3155 520 3156
rect 514 3151 515 3155
rect 519 3151 520 3155
rect 514 3150 520 3151
rect 318 3146 324 3147
rect 318 3142 319 3146
rect 323 3142 324 3146
rect 318 3141 324 3142
rect 462 3146 468 3147
rect 462 3142 463 3146
rect 467 3142 468 3146
rect 462 3141 468 3142
rect 226 3119 232 3120
rect 226 3115 227 3119
rect 231 3115 232 3119
rect 226 3114 232 3115
rect 358 3119 364 3120
rect 358 3115 359 3119
rect 363 3115 364 3119
rect 358 3114 364 3115
rect 110 3111 116 3112
rect 110 3107 111 3111
rect 115 3107 116 3111
rect 110 3106 116 3107
rect 166 3108 172 3109
rect 112 3075 114 3106
rect 166 3104 167 3108
rect 171 3104 172 3108
rect 166 3103 172 3104
rect 310 3108 316 3109
rect 310 3104 311 3108
rect 315 3104 316 3108
rect 310 3103 316 3104
rect 168 3075 170 3103
rect 312 3075 314 3103
rect 111 3074 115 3075
rect 111 3069 115 3070
rect 135 3074 139 3075
rect 135 3069 139 3070
rect 167 3074 171 3075
rect 167 3069 171 3070
rect 223 3074 227 3075
rect 223 3069 227 3070
rect 311 3074 315 3075
rect 311 3069 315 3070
rect 327 3074 331 3075
rect 327 3069 331 3070
rect 112 3050 114 3069
rect 136 3053 138 3069
rect 224 3053 226 3069
rect 328 3053 330 3069
rect 134 3052 140 3053
rect 110 3049 116 3050
rect 110 3045 111 3049
rect 115 3045 116 3049
rect 134 3048 135 3052
rect 139 3048 140 3052
rect 134 3047 140 3048
rect 222 3052 228 3053
rect 222 3048 223 3052
rect 227 3048 228 3052
rect 222 3047 228 3048
rect 326 3052 332 3053
rect 326 3048 327 3052
rect 331 3048 332 3052
rect 326 3047 332 3048
rect 110 3044 116 3045
rect 202 3043 208 3044
rect 202 3039 203 3043
rect 207 3039 208 3043
rect 202 3038 208 3039
rect 290 3043 296 3044
rect 290 3039 291 3043
rect 295 3039 296 3043
rect 290 3038 296 3039
rect 194 3035 200 3036
rect 110 3032 116 3033
rect 110 3028 111 3032
rect 115 3028 116 3032
rect 194 3031 195 3035
rect 199 3031 200 3035
rect 194 3030 200 3031
rect 110 3027 116 3028
rect 112 2987 114 3027
rect 142 3014 148 3015
rect 142 3010 143 3014
rect 147 3010 148 3014
rect 142 3009 148 3010
rect 144 2987 146 3009
rect 111 2986 115 2987
rect 111 2981 115 2982
rect 143 2986 147 2987
rect 143 2981 147 2982
rect 159 2986 163 2987
rect 159 2981 163 2982
rect 112 2953 114 2981
rect 160 2971 162 2981
rect 196 2980 198 3030
rect 204 3004 206 3038
rect 230 3014 236 3015
rect 230 3010 231 3014
rect 235 3010 236 3014
rect 230 3009 236 3010
rect 202 3003 208 3004
rect 202 2999 203 3003
rect 207 2999 208 3003
rect 202 2998 208 2999
rect 232 2987 234 3009
rect 292 3004 294 3038
rect 334 3014 340 3015
rect 334 3010 335 3014
rect 339 3010 340 3014
rect 334 3009 340 3010
rect 290 3003 296 3004
rect 290 2999 291 3003
rect 295 2999 296 3003
rect 290 2998 296 2999
rect 336 2987 338 3009
rect 360 3004 362 3114
rect 454 3108 460 3109
rect 454 3104 455 3108
rect 459 3104 460 3108
rect 454 3103 460 3104
rect 456 3075 458 3103
rect 439 3074 443 3075
rect 439 3069 443 3070
rect 455 3074 459 3075
rect 455 3069 459 3070
rect 440 3053 442 3069
rect 438 3052 444 3053
rect 438 3048 439 3052
rect 443 3048 444 3052
rect 438 3047 444 3048
rect 500 3036 502 3150
rect 516 3120 518 3150
rect 608 3147 610 3157
rect 658 3155 664 3156
rect 658 3151 659 3155
rect 663 3151 664 3155
rect 658 3150 664 3151
rect 606 3146 612 3147
rect 606 3142 607 3146
rect 611 3142 612 3146
rect 606 3141 612 3142
rect 660 3120 662 3150
rect 744 3147 746 3157
rect 872 3147 874 3157
rect 912 3156 914 3167
rect 1056 3163 1058 3181
rect 1079 3180 1083 3181
rect 1116 3176 1118 3210
rect 1198 3186 1204 3187
rect 1198 3182 1199 3186
rect 1203 3182 1204 3186
rect 1198 3181 1204 3182
rect 1078 3175 1084 3176
rect 1078 3171 1079 3175
rect 1083 3171 1084 3175
rect 1078 3170 1084 3171
rect 1114 3175 1120 3176
rect 1114 3171 1115 3175
rect 1119 3171 1120 3175
rect 1114 3170 1120 3171
rect 1200 3163 1202 3181
rect 1284 3176 1286 3210
rect 1334 3186 1340 3187
rect 1334 3182 1335 3186
rect 1339 3182 1340 3186
rect 1334 3181 1340 3182
rect 1400 3181 1402 3246
rect 1463 3241 1467 3242
rect 1607 3246 1611 3247
rect 1607 3241 1611 3242
rect 1831 3246 1835 3247
rect 1978 3243 1979 3247
rect 1983 3243 1984 3247
rect 1978 3242 1984 3243
rect 2070 3247 2076 3248
rect 2070 3243 2071 3247
rect 2075 3243 2076 3247
rect 2070 3242 2076 3243
rect 2198 3247 2204 3248
rect 2198 3243 2199 3247
rect 2203 3243 2204 3247
rect 2198 3242 2204 3243
rect 1831 3241 1835 3242
rect 1464 3225 1466 3241
rect 1608 3225 1610 3241
rect 1462 3224 1468 3225
rect 1462 3220 1463 3224
rect 1467 3220 1468 3224
rect 1462 3219 1468 3220
rect 1606 3224 1612 3225
rect 1606 3220 1607 3224
rect 1611 3220 1612 3224
rect 1832 3222 1834 3241
rect 1870 3239 1876 3240
rect 1870 3235 1871 3239
rect 1875 3235 1876 3239
rect 1870 3234 1876 3235
rect 1918 3236 1924 3237
rect 1606 3219 1612 3220
rect 1830 3221 1836 3222
rect 1830 3217 1831 3221
rect 1835 3217 1836 3221
rect 1830 3216 1836 3217
rect 1418 3215 1424 3216
rect 1418 3211 1419 3215
rect 1423 3211 1424 3215
rect 1418 3210 1424 3211
rect 1558 3215 1564 3216
rect 1558 3211 1559 3215
rect 1563 3211 1564 3215
rect 1558 3210 1564 3211
rect 1586 3215 1592 3216
rect 1872 3215 1874 3234
rect 1918 3232 1919 3236
rect 1923 3232 1924 3236
rect 1918 3231 1924 3232
rect 2054 3236 2060 3237
rect 2054 3232 2055 3236
rect 2059 3232 2060 3236
rect 2054 3231 2060 3232
rect 2182 3236 2188 3237
rect 2182 3232 2183 3236
rect 2187 3232 2188 3236
rect 2182 3231 2188 3232
rect 1920 3215 1922 3231
rect 2056 3215 2058 3231
rect 2184 3215 2186 3231
rect 1586 3211 1587 3215
rect 1591 3211 1592 3215
rect 1586 3210 1592 3211
rect 1871 3214 1875 3215
rect 1282 3175 1288 3176
rect 1282 3171 1283 3175
rect 1287 3171 1288 3175
rect 1282 3170 1288 3171
rect 1336 3163 1338 3181
rect 1399 3180 1403 3181
rect 1420 3176 1422 3210
rect 1470 3186 1476 3187
rect 1470 3182 1471 3186
rect 1475 3182 1476 3186
rect 1470 3181 1476 3182
rect 1399 3175 1403 3176
rect 1418 3175 1424 3176
rect 1418 3171 1419 3175
rect 1423 3171 1424 3175
rect 1418 3170 1424 3171
rect 1472 3163 1474 3181
rect 1560 3176 1562 3210
rect 1588 3197 1590 3210
rect 1871 3209 1875 3210
rect 1895 3214 1899 3215
rect 1895 3209 1899 3210
rect 1919 3214 1923 3215
rect 1919 3209 1923 3210
rect 2007 3214 2011 3215
rect 2007 3209 2011 3210
rect 2055 3214 2059 3215
rect 2055 3209 2059 3210
rect 2143 3214 2147 3215
rect 2143 3209 2147 3210
rect 2183 3214 2187 3215
rect 2183 3209 2187 3210
rect 1830 3204 1836 3205
rect 1830 3200 1831 3204
rect 1835 3200 1836 3204
rect 1830 3199 1836 3200
rect 1587 3196 1591 3197
rect 1587 3191 1591 3192
rect 1614 3186 1620 3187
rect 1614 3182 1615 3186
rect 1619 3182 1620 3186
rect 1614 3181 1620 3182
rect 1558 3175 1564 3176
rect 1558 3171 1559 3175
rect 1563 3171 1564 3175
rect 1558 3170 1564 3171
rect 1616 3163 1618 3181
rect 1832 3163 1834 3199
rect 1872 3190 1874 3209
rect 1896 3193 1898 3209
rect 2008 3193 2010 3209
rect 2144 3193 2146 3209
rect 1894 3192 1900 3193
rect 1870 3189 1876 3190
rect 1870 3185 1871 3189
rect 1875 3185 1876 3189
rect 1894 3188 1895 3192
rect 1899 3188 1900 3192
rect 1894 3187 1900 3188
rect 2006 3192 2012 3193
rect 2006 3188 2007 3192
rect 2011 3188 2012 3192
rect 2006 3187 2012 3188
rect 2142 3192 2148 3193
rect 2142 3188 2143 3192
rect 2147 3188 2148 3192
rect 2142 3187 2148 3188
rect 1870 3184 1876 3185
rect 2212 3184 2214 3278
rect 2320 3275 2322 3285
rect 2448 3275 2450 3285
rect 2500 3284 2502 3322
rect 2508 3296 2510 3330
rect 2590 3306 2596 3307
rect 2590 3302 2591 3306
rect 2595 3302 2596 3306
rect 2590 3301 2596 3302
rect 2506 3295 2512 3296
rect 2506 3291 2507 3295
rect 2511 3291 2512 3295
rect 2592 3291 2594 3301
rect 2620 3296 2622 3366
rect 2671 3361 2675 3362
rect 2727 3366 2731 3367
rect 2727 3361 2731 3362
rect 2823 3366 2827 3367
rect 2823 3361 2827 3362
rect 2871 3366 2875 3367
rect 2871 3361 2875 3362
rect 2991 3366 2995 3367
rect 2991 3361 2995 3362
rect 3023 3366 3027 3367
rect 3023 3361 3027 3362
rect 3159 3366 3163 3367
rect 3159 3361 3163 3362
rect 3183 3366 3187 3367
rect 3183 3361 3187 3362
rect 3335 3366 3339 3367
rect 3335 3361 3339 3362
rect 3351 3366 3355 3367
rect 3351 3361 3355 3362
rect 2728 3345 2730 3361
rect 2872 3345 2874 3361
rect 3024 3345 3026 3361
rect 3184 3345 3186 3361
rect 3352 3345 3354 3361
rect 2726 3344 2732 3345
rect 2726 3340 2727 3344
rect 2731 3340 2732 3344
rect 2726 3339 2732 3340
rect 2870 3344 2876 3345
rect 2870 3340 2871 3344
rect 2875 3340 2876 3344
rect 2870 3339 2876 3340
rect 3022 3344 3028 3345
rect 3022 3340 3023 3344
rect 3027 3340 3028 3344
rect 3022 3339 3028 3340
rect 3182 3344 3188 3345
rect 3182 3340 3183 3344
rect 3187 3340 3188 3344
rect 3182 3339 3188 3340
rect 3350 3344 3356 3345
rect 3350 3340 3351 3344
rect 3355 3340 3356 3344
rect 3350 3339 3356 3340
rect 2794 3335 2800 3336
rect 2794 3331 2795 3335
rect 2799 3331 2800 3335
rect 2794 3330 2800 3331
rect 2970 3335 2976 3336
rect 2970 3331 2971 3335
rect 2975 3331 2976 3335
rect 2970 3330 2976 3331
rect 3126 3335 3132 3336
rect 3126 3331 3127 3335
rect 3131 3331 3132 3335
rect 3126 3330 3132 3331
rect 3290 3335 3296 3336
rect 3290 3331 3291 3335
rect 3295 3331 3296 3335
rect 3360 3332 3362 3430
rect 3512 3427 3514 3437
rect 3564 3436 3566 3474
rect 3590 3472 3591 3476
rect 3595 3472 3596 3476
rect 3590 3471 3596 3472
rect 3592 3443 3594 3471
rect 3591 3442 3595 3443
rect 3591 3437 3595 3438
rect 3562 3435 3568 3436
rect 3562 3431 3563 3435
rect 3567 3431 3568 3435
rect 3562 3430 3568 3431
rect 3510 3426 3516 3427
rect 3510 3422 3511 3426
rect 3515 3422 3516 3426
rect 3510 3421 3516 3422
rect 3592 3409 3594 3437
rect 3590 3408 3596 3409
rect 3590 3404 3591 3408
rect 3595 3404 3596 3408
rect 3590 3403 3596 3404
rect 3534 3399 3540 3400
rect 3534 3395 3535 3399
rect 3539 3395 3540 3399
rect 3534 3394 3540 3395
rect 3502 3388 3508 3389
rect 3502 3384 3503 3388
rect 3507 3384 3508 3388
rect 3502 3383 3508 3384
rect 3504 3367 3506 3383
rect 3503 3366 3507 3367
rect 3503 3361 3507 3362
rect 3504 3345 3506 3361
rect 3502 3344 3508 3345
rect 3502 3340 3503 3344
rect 3507 3340 3508 3344
rect 3502 3339 3508 3340
rect 3290 3330 3296 3331
rect 3358 3331 3364 3332
rect 2734 3306 2740 3307
rect 2734 3302 2735 3306
rect 2739 3302 2740 3306
rect 2734 3301 2740 3302
rect 2618 3295 2624 3296
rect 2618 3291 2619 3295
rect 2623 3291 2624 3295
rect 2736 3291 2738 3301
rect 2796 3296 2798 3330
rect 2878 3306 2884 3307
rect 2878 3302 2879 3306
rect 2883 3302 2884 3306
rect 2878 3301 2884 3302
rect 2786 3295 2792 3296
rect 2786 3291 2787 3295
rect 2791 3291 2792 3295
rect 2506 3290 2512 3291
rect 2591 3290 2595 3291
rect 2618 3290 2624 3291
rect 2735 3290 2739 3291
rect 2591 3285 2595 3286
rect 2735 3285 2739 3286
rect 2743 3290 2747 3291
rect 2786 3290 2792 3291
rect 2794 3295 2800 3296
rect 2794 3291 2795 3295
rect 2799 3291 2800 3295
rect 2880 3291 2882 3301
rect 2972 3296 2974 3330
rect 3030 3306 3036 3307
rect 3030 3302 3031 3306
rect 3035 3302 3036 3306
rect 3030 3301 3036 3302
rect 2970 3295 2976 3296
rect 2970 3291 2971 3295
rect 2975 3291 2976 3295
rect 3032 3291 3034 3301
rect 3128 3296 3130 3330
rect 3190 3306 3196 3307
rect 3190 3302 3191 3306
rect 3195 3302 3196 3306
rect 3190 3301 3196 3302
rect 3126 3295 3132 3296
rect 3126 3291 3127 3295
rect 3131 3291 3132 3295
rect 3192 3291 3194 3301
rect 3292 3296 3294 3330
rect 3358 3327 3359 3331
rect 3363 3327 3364 3331
rect 3358 3326 3364 3327
rect 3358 3306 3364 3307
rect 3358 3302 3359 3306
rect 3363 3302 3364 3306
rect 3358 3301 3364 3302
rect 3510 3306 3516 3307
rect 3510 3302 3511 3306
rect 3515 3302 3516 3306
rect 3510 3301 3516 3302
rect 3290 3295 3296 3296
rect 3290 3291 3291 3295
rect 3295 3291 3296 3295
rect 3360 3291 3362 3301
rect 3512 3291 3514 3301
rect 3536 3296 3538 3394
rect 3590 3391 3596 3392
rect 3590 3387 3591 3391
rect 3595 3387 3596 3391
rect 3590 3386 3596 3387
rect 3592 3367 3594 3386
rect 3591 3366 3595 3367
rect 3591 3361 3595 3362
rect 3592 3342 3594 3361
rect 3590 3341 3596 3342
rect 3590 3337 3591 3341
rect 3595 3337 3596 3341
rect 3590 3336 3596 3337
rect 3562 3327 3568 3328
rect 3562 3323 3563 3327
rect 3567 3323 3568 3327
rect 3562 3322 3568 3323
rect 3590 3324 3596 3325
rect 3534 3295 3540 3296
rect 3534 3291 3535 3295
rect 3539 3291 3540 3295
rect 2794 3290 2800 3291
rect 2879 3290 2883 3291
rect 2743 3285 2747 3286
rect 2454 3283 2460 3284
rect 2454 3279 2455 3283
rect 2459 3279 2460 3283
rect 2454 3278 2460 3279
rect 2498 3283 2504 3284
rect 2498 3279 2499 3283
rect 2503 3279 2504 3283
rect 2498 3278 2504 3279
rect 2318 3274 2324 3275
rect 2318 3270 2319 3274
rect 2323 3270 2324 3274
rect 2318 3269 2324 3270
rect 2446 3274 2452 3275
rect 2446 3270 2447 3274
rect 2451 3270 2452 3274
rect 2446 3269 2452 3270
rect 2456 3248 2458 3278
rect 2592 3275 2594 3285
rect 2614 3283 2620 3284
rect 2614 3279 2615 3283
rect 2619 3279 2620 3283
rect 2614 3278 2620 3279
rect 2642 3283 2648 3284
rect 2642 3279 2643 3283
rect 2647 3279 2648 3283
rect 2642 3278 2648 3279
rect 2590 3274 2596 3275
rect 2590 3270 2591 3274
rect 2595 3270 2596 3274
rect 2590 3269 2596 3270
rect 2454 3247 2460 3248
rect 2454 3243 2455 3247
rect 2459 3243 2460 3247
rect 2454 3242 2460 3243
rect 2310 3236 2316 3237
rect 2310 3232 2311 3236
rect 2315 3232 2316 3236
rect 2310 3231 2316 3232
rect 2438 3236 2444 3237
rect 2438 3232 2439 3236
rect 2443 3232 2444 3236
rect 2438 3231 2444 3232
rect 2582 3236 2588 3237
rect 2582 3232 2583 3236
rect 2587 3232 2588 3236
rect 2582 3231 2588 3232
rect 2312 3215 2314 3231
rect 2326 3219 2332 3220
rect 2326 3215 2327 3219
rect 2331 3215 2332 3219
rect 2440 3215 2442 3231
rect 2584 3215 2586 3231
rect 2295 3214 2299 3215
rect 2295 3209 2299 3210
rect 2311 3214 2315 3215
rect 2326 3214 2332 3215
rect 2439 3214 2443 3215
rect 2311 3209 2315 3210
rect 2296 3193 2298 3209
rect 2294 3192 2300 3193
rect 2294 3188 2295 3192
rect 2299 3188 2300 3192
rect 2294 3187 2300 3188
rect 1962 3183 1968 3184
rect 1962 3179 1963 3183
rect 1967 3179 1968 3183
rect 1962 3178 1968 3179
rect 2090 3183 2096 3184
rect 2090 3179 2091 3183
rect 2095 3179 2096 3183
rect 2090 3178 2096 3179
rect 2210 3183 2216 3184
rect 2210 3179 2211 3183
rect 2215 3179 2216 3183
rect 2210 3178 2216 3179
rect 1870 3172 1876 3173
rect 1870 3168 1871 3172
rect 1875 3168 1876 3172
rect 1870 3167 1876 3168
rect 991 3162 995 3163
rect 991 3157 995 3158
rect 1055 3162 1059 3163
rect 1055 3157 1059 3158
rect 1103 3162 1107 3163
rect 1103 3157 1107 3158
rect 1199 3162 1203 3163
rect 1199 3157 1203 3158
rect 1207 3162 1211 3163
rect 1207 3157 1211 3158
rect 1311 3162 1315 3163
rect 1311 3157 1315 3158
rect 1335 3162 1339 3163
rect 1335 3157 1339 3158
rect 1407 3162 1411 3163
rect 1407 3157 1411 3158
rect 1471 3162 1475 3163
rect 1471 3157 1475 3158
rect 1495 3162 1499 3163
rect 1495 3157 1499 3158
rect 1583 3162 1587 3163
rect 1583 3157 1587 3158
rect 1615 3162 1619 3163
rect 1615 3157 1619 3158
rect 1671 3162 1675 3163
rect 1671 3157 1675 3158
rect 1751 3162 1755 3163
rect 1751 3157 1755 3158
rect 1831 3162 1835 3163
rect 1831 3157 1835 3158
rect 910 3155 916 3156
rect 910 3151 911 3155
rect 915 3151 916 3155
rect 910 3150 916 3151
rect 922 3155 928 3156
rect 922 3151 923 3155
rect 927 3151 928 3155
rect 922 3150 928 3151
rect 742 3146 748 3147
rect 742 3142 743 3146
rect 747 3142 748 3146
rect 742 3141 748 3142
rect 870 3146 876 3147
rect 870 3142 871 3146
rect 875 3142 876 3146
rect 870 3141 876 3142
rect 924 3120 926 3150
rect 992 3147 994 3157
rect 1042 3155 1048 3156
rect 1042 3151 1043 3155
rect 1047 3151 1048 3155
rect 1042 3150 1048 3151
rect 990 3146 996 3147
rect 990 3142 991 3146
rect 995 3142 996 3146
rect 990 3141 996 3142
rect 1044 3120 1046 3150
rect 1104 3147 1106 3157
rect 1154 3155 1160 3156
rect 1154 3151 1155 3155
rect 1159 3151 1160 3155
rect 1154 3150 1160 3151
rect 1102 3146 1108 3147
rect 1102 3142 1103 3146
rect 1107 3142 1108 3146
rect 1102 3141 1108 3142
rect 1156 3120 1158 3150
rect 1208 3147 1210 3157
rect 1258 3155 1264 3156
rect 1258 3151 1259 3155
rect 1263 3151 1264 3155
rect 1258 3150 1264 3151
rect 1206 3146 1212 3147
rect 1206 3142 1207 3146
rect 1211 3142 1212 3146
rect 1206 3141 1212 3142
rect 1260 3120 1262 3150
rect 1312 3147 1314 3157
rect 1362 3155 1368 3156
rect 1362 3151 1363 3155
rect 1367 3151 1368 3155
rect 1362 3150 1368 3151
rect 1310 3146 1316 3147
rect 1310 3142 1311 3146
rect 1315 3142 1316 3146
rect 1310 3141 1316 3142
rect 1364 3120 1366 3150
rect 1408 3147 1410 3157
rect 1458 3155 1464 3156
rect 1458 3151 1459 3155
rect 1463 3151 1464 3155
rect 1458 3150 1464 3151
rect 1406 3146 1412 3147
rect 1406 3142 1407 3146
rect 1411 3142 1412 3146
rect 1406 3141 1412 3142
rect 1460 3120 1462 3150
rect 1496 3147 1498 3157
rect 1546 3155 1552 3156
rect 1546 3151 1547 3155
rect 1551 3151 1552 3155
rect 1546 3150 1552 3151
rect 1494 3146 1500 3147
rect 1494 3142 1495 3146
rect 1499 3142 1500 3146
rect 1494 3141 1500 3142
rect 1548 3120 1550 3150
rect 1584 3147 1586 3157
rect 1634 3155 1640 3156
rect 1634 3151 1635 3155
rect 1639 3151 1640 3155
rect 1634 3150 1640 3151
rect 1582 3146 1588 3147
rect 1582 3142 1583 3146
rect 1587 3142 1588 3146
rect 1582 3141 1588 3142
rect 1636 3120 1638 3150
rect 1672 3147 1674 3157
rect 1722 3155 1728 3156
rect 1722 3151 1723 3155
rect 1727 3151 1728 3155
rect 1722 3150 1728 3151
rect 1670 3146 1676 3147
rect 1670 3142 1671 3146
rect 1675 3142 1676 3146
rect 1670 3141 1676 3142
rect 1724 3120 1726 3150
rect 1752 3147 1754 3157
rect 1750 3146 1756 3147
rect 1750 3142 1751 3146
rect 1755 3142 1756 3146
rect 1750 3141 1756 3142
rect 1832 3129 1834 3157
rect 1872 3139 1874 3167
rect 1902 3154 1908 3155
rect 1902 3150 1903 3154
rect 1907 3150 1908 3154
rect 1902 3149 1908 3150
rect 1904 3139 1906 3149
rect 1964 3144 1966 3178
rect 2014 3154 2020 3155
rect 2014 3150 2015 3154
rect 2019 3150 2020 3154
rect 2014 3149 2020 3150
rect 1926 3143 1932 3144
rect 1926 3139 1927 3143
rect 1931 3139 1932 3143
rect 1871 3138 1875 3139
rect 1871 3133 1875 3134
rect 1903 3138 1907 3139
rect 1926 3138 1932 3139
rect 1962 3143 1968 3144
rect 1962 3139 1963 3143
rect 1967 3139 1968 3143
rect 2016 3139 2018 3149
rect 2092 3144 2094 3178
rect 2150 3154 2156 3155
rect 2150 3150 2151 3154
rect 2155 3150 2156 3154
rect 2150 3149 2156 3150
rect 2302 3154 2308 3155
rect 2302 3150 2303 3154
rect 2307 3150 2308 3154
rect 2302 3149 2308 3150
rect 2090 3143 2096 3144
rect 2090 3139 2091 3143
rect 2095 3139 2096 3143
rect 2152 3139 2154 3149
rect 2304 3139 2306 3149
rect 2328 3144 2330 3214
rect 2439 3209 2443 3210
rect 2455 3214 2459 3215
rect 2455 3209 2459 3210
rect 2583 3214 2587 3215
rect 2583 3209 2587 3210
rect 2456 3193 2458 3209
rect 2454 3192 2460 3193
rect 2454 3188 2455 3192
rect 2459 3188 2460 3192
rect 2454 3187 2460 3188
rect 2616 3184 2618 3278
rect 2644 3248 2646 3278
rect 2744 3275 2746 3285
rect 2742 3274 2748 3275
rect 2742 3270 2743 3274
rect 2747 3270 2748 3274
rect 2742 3269 2748 3270
rect 2788 3269 2790 3290
rect 2879 3285 2883 3286
rect 2919 3290 2923 3291
rect 2970 3290 2976 3291
rect 3031 3290 3035 3291
rect 2919 3285 2923 3286
rect 3031 3285 3035 3286
rect 3111 3290 3115 3291
rect 3126 3290 3132 3291
rect 3191 3290 3195 3291
rect 3290 3290 3296 3291
rect 3311 3290 3315 3291
rect 3111 3285 3115 3286
rect 3191 3285 3195 3286
rect 3311 3285 3315 3286
rect 3359 3290 3363 3291
rect 3359 3285 3363 3286
rect 3511 3290 3515 3291
rect 3534 3290 3540 3291
rect 3511 3285 3515 3286
rect 2794 3283 2800 3284
rect 2794 3279 2795 3283
rect 2799 3279 2800 3283
rect 2794 3278 2800 3279
rect 2787 3268 2791 3269
rect 2787 3263 2791 3264
rect 2796 3248 2798 3278
rect 2920 3275 2922 3285
rect 2970 3283 2976 3284
rect 2970 3279 2971 3283
rect 2975 3279 2976 3283
rect 2970 3278 2976 3279
rect 2918 3274 2924 3275
rect 2918 3270 2919 3274
rect 2923 3270 2924 3274
rect 2918 3269 2924 3270
rect 2972 3248 2974 3278
rect 3112 3275 3114 3285
rect 3162 3283 3168 3284
rect 3162 3279 3163 3283
rect 3167 3279 3168 3283
rect 3162 3278 3168 3279
rect 3110 3274 3116 3275
rect 3110 3270 3111 3274
rect 3115 3270 3116 3274
rect 3110 3269 3116 3270
rect 3164 3248 3166 3278
rect 3312 3275 3314 3285
rect 3512 3275 3514 3285
rect 3564 3284 3566 3322
rect 3590 3320 3591 3324
rect 3595 3320 3596 3324
rect 3590 3319 3596 3320
rect 3592 3291 3594 3319
rect 3591 3290 3595 3291
rect 3591 3285 3595 3286
rect 3562 3283 3568 3284
rect 3562 3279 3563 3283
rect 3567 3279 3568 3283
rect 3562 3278 3568 3279
rect 3310 3274 3316 3275
rect 3310 3270 3311 3274
rect 3315 3270 3316 3274
rect 3310 3269 3316 3270
rect 3510 3274 3516 3275
rect 3510 3270 3511 3274
rect 3515 3270 3516 3274
rect 3510 3269 3516 3270
rect 3319 3268 3323 3269
rect 3319 3263 3323 3264
rect 3320 3248 3322 3263
rect 3592 3257 3594 3285
rect 3590 3256 3596 3257
rect 3590 3252 3591 3256
rect 3595 3252 3596 3256
rect 3590 3251 3596 3252
rect 2642 3247 2648 3248
rect 2642 3243 2643 3247
rect 2647 3243 2648 3247
rect 2642 3242 2648 3243
rect 2794 3247 2800 3248
rect 2794 3243 2795 3247
rect 2799 3243 2800 3247
rect 2794 3242 2800 3243
rect 2970 3247 2976 3248
rect 2970 3243 2971 3247
rect 2975 3243 2976 3247
rect 2970 3242 2976 3243
rect 3162 3247 3168 3248
rect 3162 3243 3163 3247
rect 3167 3243 3168 3247
rect 3162 3242 3168 3243
rect 3318 3247 3324 3248
rect 3318 3243 3319 3247
rect 3323 3243 3324 3247
rect 3318 3242 3324 3243
rect 3534 3247 3540 3248
rect 3534 3243 3535 3247
rect 3539 3243 3540 3247
rect 3534 3242 3540 3243
rect 2734 3236 2740 3237
rect 2734 3232 2735 3236
rect 2739 3232 2740 3236
rect 2734 3231 2740 3232
rect 2910 3236 2916 3237
rect 2910 3232 2911 3236
rect 2915 3232 2916 3236
rect 2910 3231 2916 3232
rect 3102 3236 3108 3237
rect 3102 3232 3103 3236
rect 3107 3232 3108 3236
rect 3102 3231 3108 3232
rect 3302 3236 3308 3237
rect 3302 3232 3303 3236
rect 3307 3232 3308 3236
rect 3302 3231 3308 3232
rect 3502 3236 3508 3237
rect 3502 3232 3503 3236
rect 3507 3232 3508 3236
rect 3502 3231 3508 3232
rect 2736 3215 2738 3231
rect 2912 3215 2914 3231
rect 3104 3215 3106 3231
rect 3304 3215 3306 3231
rect 3504 3215 3506 3231
rect 2623 3214 2627 3215
rect 2623 3209 2627 3210
rect 2735 3214 2739 3215
rect 2735 3209 2739 3210
rect 2799 3214 2803 3215
rect 2799 3209 2803 3210
rect 2911 3214 2915 3215
rect 2911 3209 2915 3210
rect 2975 3214 2979 3215
rect 2975 3209 2979 3210
rect 3103 3214 3107 3215
rect 3103 3209 3107 3210
rect 3151 3214 3155 3215
rect 3151 3209 3155 3210
rect 3303 3214 3307 3215
rect 3303 3209 3307 3210
rect 3327 3214 3331 3215
rect 3327 3209 3331 3210
rect 3503 3214 3507 3215
rect 3503 3209 3507 3210
rect 2624 3193 2626 3209
rect 2800 3193 2802 3209
rect 2976 3193 2978 3209
rect 3152 3193 3154 3209
rect 3328 3193 3330 3209
rect 3504 3193 3506 3209
rect 2622 3192 2628 3193
rect 2622 3188 2623 3192
rect 2627 3188 2628 3192
rect 2622 3187 2628 3188
rect 2798 3192 2804 3193
rect 2798 3188 2799 3192
rect 2803 3188 2804 3192
rect 2798 3187 2804 3188
rect 2974 3192 2980 3193
rect 2974 3188 2975 3192
rect 2979 3188 2980 3192
rect 2974 3187 2980 3188
rect 3150 3192 3156 3193
rect 3150 3188 3151 3192
rect 3155 3188 3156 3192
rect 3150 3187 3156 3188
rect 3326 3192 3332 3193
rect 3326 3188 3327 3192
rect 3331 3188 3332 3192
rect 3326 3187 3332 3188
rect 3502 3192 3508 3193
rect 3502 3188 3503 3192
rect 3507 3188 3508 3192
rect 3502 3187 3508 3188
rect 2370 3183 2376 3184
rect 2370 3179 2371 3183
rect 2375 3179 2376 3183
rect 2614 3183 2620 3184
rect 2370 3178 2376 3179
rect 2462 3179 2468 3180
rect 2372 3144 2374 3178
rect 2462 3175 2463 3179
rect 2467 3175 2468 3179
rect 2614 3179 2615 3183
rect 2619 3179 2620 3183
rect 2614 3178 2620 3179
rect 2690 3183 2696 3184
rect 2690 3179 2691 3183
rect 2695 3179 2696 3183
rect 2690 3178 2696 3179
rect 2914 3183 2920 3184
rect 2914 3179 2915 3183
rect 2919 3179 2920 3183
rect 2914 3178 2920 3179
rect 3262 3183 3268 3184
rect 3262 3179 3263 3183
rect 3267 3179 3268 3183
rect 3262 3178 3268 3179
rect 3398 3183 3404 3184
rect 3398 3179 3399 3183
rect 3403 3179 3404 3183
rect 3398 3178 3404 3179
rect 2462 3174 2468 3175
rect 2464 3163 2466 3174
rect 2464 3161 2474 3163
rect 2462 3154 2468 3155
rect 2462 3150 2463 3154
rect 2467 3150 2468 3154
rect 2462 3149 2468 3150
rect 2326 3143 2332 3144
rect 2326 3139 2327 3143
rect 2331 3139 2332 3143
rect 1962 3138 1968 3139
rect 2015 3138 2019 3139
rect 1903 3133 1907 3134
rect 1830 3128 1836 3129
rect 1830 3124 1831 3128
rect 1835 3124 1836 3128
rect 1830 3123 1836 3124
rect 514 3119 520 3120
rect 514 3115 515 3119
rect 519 3115 520 3119
rect 514 3114 520 3115
rect 658 3119 664 3120
rect 658 3115 659 3119
rect 663 3115 664 3119
rect 658 3114 664 3115
rect 922 3119 928 3120
rect 922 3115 923 3119
rect 927 3115 928 3119
rect 922 3114 928 3115
rect 1042 3119 1048 3120
rect 1042 3115 1043 3119
rect 1047 3115 1048 3119
rect 1042 3114 1048 3115
rect 1154 3119 1160 3120
rect 1154 3115 1155 3119
rect 1159 3115 1160 3119
rect 1154 3114 1160 3115
rect 1258 3119 1264 3120
rect 1258 3115 1259 3119
rect 1263 3115 1264 3119
rect 1258 3114 1264 3115
rect 1362 3119 1368 3120
rect 1362 3115 1363 3119
rect 1367 3115 1368 3119
rect 1362 3114 1368 3115
rect 1458 3119 1464 3120
rect 1458 3115 1459 3119
rect 1463 3115 1464 3119
rect 1458 3114 1464 3115
rect 1546 3119 1552 3120
rect 1546 3115 1547 3119
rect 1551 3115 1552 3119
rect 1546 3114 1552 3115
rect 1634 3119 1640 3120
rect 1634 3115 1635 3119
rect 1639 3115 1640 3119
rect 1634 3114 1640 3115
rect 1722 3119 1728 3120
rect 1722 3115 1723 3119
rect 1727 3115 1728 3119
rect 1722 3114 1728 3115
rect 1830 3111 1836 3112
rect 598 3108 604 3109
rect 598 3104 599 3108
rect 603 3104 604 3108
rect 598 3103 604 3104
rect 734 3108 740 3109
rect 734 3104 735 3108
rect 739 3104 740 3108
rect 734 3103 740 3104
rect 862 3108 868 3109
rect 862 3104 863 3108
rect 867 3104 868 3108
rect 862 3103 868 3104
rect 982 3108 988 3109
rect 982 3104 983 3108
rect 987 3104 988 3108
rect 982 3103 988 3104
rect 1094 3108 1100 3109
rect 1094 3104 1095 3108
rect 1099 3104 1100 3108
rect 1094 3103 1100 3104
rect 1198 3108 1204 3109
rect 1198 3104 1199 3108
rect 1203 3104 1204 3108
rect 1198 3103 1204 3104
rect 1302 3108 1308 3109
rect 1302 3104 1303 3108
rect 1307 3104 1308 3108
rect 1302 3103 1308 3104
rect 1398 3108 1404 3109
rect 1398 3104 1399 3108
rect 1403 3104 1404 3108
rect 1398 3103 1404 3104
rect 1486 3108 1492 3109
rect 1486 3104 1487 3108
rect 1491 3104 1492 3108
rect 1486 3103 1492 3104
rect 1574 3108 1580 3109
rect 1574 3104 1575 3108
rect 1579 3104 1580 3108
rect 1574 3103 1580 3104
rect 1662 3108 1668 3109
rect 1662 3104 1663 3108
rect 1667 3104 1668 3108
rect 1662 3103 1668 3104
rect 1742 3108 1748 3109
rect 1742 3104 1743 3108
rect 1747 3104 1748 3108
rect 1830 3107 1831 3111
rect 1835 3107 1836 3111
rect 1830 3106 1836 3107
rect 1742 3103 1748 3104
rect 600 3075 602 3103
rect 736 3075 738 3103
rect 864 3075 866 3103
rect 984 3075 986 3103
rect 1096 3075 1098 3103
rect 1200 3075 1202 3103
rect 1304 3075 1306 3103
rect 1400 3075 1402 3103
rect 1488 3075 1490 3103
rect 1576 3075 1578 3103
rect 1664 3075 1666 3103
rect 1744 3075 1746 3103
rect 1832 3075 1834 3106
rect 1872 3105 1874 3133
rect 1904 3123 1906 3133
rect 1902 3122 1908 3123
rect 1902 3118 1903 3122
rect 1907 3118 1908 3122
rect 1902 3117 1908 3118
rect 1870 3104 1876 3105
rect 1870 3100 1871 3104
rect 1875 3100 1876 3104
rect 1870 3099 1876 3100
rect 1928 3096 1930 3138
rect 2015 3133 2019 3134
rect 2071 3138 2075 3139
rect 2090 3138 2096 3139
rect 2151 3138 2155 3139
rect 2071 3133 2075 3134
rect 2151 3133 2155 3134
rect 2263 3138 2267 3139
rect 2263 3133 2267 3134
rect 2303 3138 2307 3139
rect 2326 3138 2332 3139
rect 2370 3143 2376 3144
rect 2370 3139 2371 3143
rect 2375 3139 2376 3143
rect 2464 3139 2466 3149
rect 2370 3138 2376 3139
rect 2455 3138 2459 3139
rect 2303 3133 2307 3134
rect 2455 3133 2459 3134
rect 2463 3138 2467 3139
rect 2463 3133 2467 3134
rect 2072 3123 2074 3133
rect 2114 3131 2120 3132
rect 2114 3127 2115 3131
rect 2119 3127 2120 3131
rect 2114 3126 2120 3127
rect 2122 3131 2128 3132
rect 2122 3127 2123 3131
rect 2127 3127 2128 3131
rect 2122 3126 2128 3127
rect 2070 3122 2076 3123
rect 2070 3118 2071 3122
rect 2075 3118 2076 3122
rect 2070 3117 2076 3118
rect 1926 3095 1932 3096
rect 1926 3091 1927 3095
rect 1931 3091 1932 3095
rect 1926 3090 1932 3091
rect 1870 3087 1876 3088
rect 1870 3083 1871 3087
rect 1875 3083 1876 3087
rect 1870 3082 1876 3083
rect 1894 3084 1900 3085
rect 551 3074 555 3075
rect 551 3069 555 3070
rect 599 3074 603 3075
rect 599 3069 603 3070
rect 663 3074 667 3075
rect 663 3069 667 3070
rect 735 3074 739 3075
rect 735 3069 739 3070
rect 863 3074 867 3075
rect 863 3069 867 3070
rect 983 3074 987 3075
rect 983 3069 987 3070
rect 1095 3074 1099 3075
rect 1095 3069 1099 3070
rect 1199 3074 1203 3075
rect 1199 3069 1203 3070
rect 1303 3074 1307 3075
rect 1303 3069 1307 3070
rect 1399 3074 1403 3075
rect 1399 3069 1403 3070
rect 1487 3074 1491 3075
rect 1487 3069 1491 3070
rect 1575 3074 1579 3075
rect 1575 3069 1579 3070
rect 1663 3074 1667 3075
rect 1663 3069 1667 3070
rect 1743 3074 1747 3075
rect 1743 3069 1747 3070
rect 1831 3074 1835 3075
rect 1831 3069 1835 3070
rect 552 3053 554 3069
rect 664 3053 666 3069
rect 550 3052 556 3053
rect 550 3048 551 3052
rect 555 3048 556 3052
rect 550 3047 556 3048
rect 662 3052 668 3053
rect 662 3048 663 3052
rect 667 3048 668 3052
rect 1832 3050 1834 3069
rect 1872 3051 1874 3082
rect 1894 3080 1895 3084
rect 1899 3080 1900 3084
rect 1894 3079 1900 3080
rect 2062 3084 2068 3085
rect 2062 3080 2063 3084
rect 2067 3080 2068 3084
rect 2062 3079 2068 3080
rect 1896 3051 1898 3079
rect 2064 3051 2066 3079
rect 2116 3068 2118 3126
rect 2124 3096 2126 3126
rect 2264 3123 2266 3133
rect 2456 3123 2458 3133
rect 2472 3132 2474 3161
rect 2630 3154 2636 3155
rect 2630 3150 2631 3154
rect 2635 3150 2636 3154
rect 2630 3149 2636 3150
rect 2632 3139 2634 3149
rect 2692 3144 2694 3178
rect 2806 3154 2812 3155
rect 2806 3150 2807 3154
rect 2811 3150 2812 3154
rect 2806 3149 2812 3150
rect 2690 3143 2696 3144
rect 2690 3139 2691 3143
rect 2695 3139 2696 3143
rect 2808 3139 2810 3149
rect 2916 3144 2918 3178
rect 3210 3175 3216 3176
rect 3210 3171 3211 3175
rect 3215 3171 3216 3175
rect 3210 3170 3216 3171
rect 2982 3154 2988 3155
rect 2982 3150 2983 3154
rect 2987 3150 2988 3154
rect 2982 3149 2988 3150
rect 3158 3154 3164 3155
rect 3158 3150 3159 3154
rect 3163 3150 3164 3154
rect 3158 3149 3164 3150
rect 2914 3143 2920 3144
rect 2914 3139 2915 3143
rect 2919 3139 2920 3143
rect 2984 3139 2986 3149
rect 3006 3143 3012 3144
rect 3006 3139 3007 3143
rect 3011 3139 3012 3143
rect 3160 3139 3162 3149
rect 3212 3144 3214 3170
rect 3264 3144 3266 3178
rect 3334 3154 3340 3155
rect 3334 3150 3335 3154
rect 3339 3150 3340 3154
rect 3334 3149 3340 3150
rect 3210 3143 3216 3144
rect 3210 3139 3211 3143
rect 3215 3139 3216 3143
rect 2631 3138 2635 3139
rect 2631 3133 2635 3134
rect 2647 3138 2651 3139
rect 2690 3138 2696 3139
rect 2807 3138 2811 3139
rect 2647 3133 2651 3134
rect 2807 3133 2811 3134
rect 2831 3138 2835 3139
rect 2914 3138 2920 3139
rect 2983 3138 2987 3139
rect 3006 3138 3012 3139
rect 3015 3138 3019 3139
rect 2831 3133 2835 3134
rect 2983 3133 2987 3134
rect 2470 3131 2476 3132
rect 2470 3127 2471 3131
rect 2475 3127 2476 3131
rect 2470 3126 2476 3127
rect 2648 3123 2650 3133
rect 2682 3131 2688 3132
rect 2682 3127 2683 3131
rect 2687 3127 2688 3131
rect 2682 3126 2688 3127
rect 2698 3131 2704 3132
rect 2698 3127 2699 3131
rect 2703 3127 2704 3131
rect 2698 3126 2704 3127
rect 2262 3122 2268 3123
rect 2262 3118 2263 3122
rect 2267 3118 2268 3122
rect 2262 3117 2268 3118
rect 2454 3122 2460 3123
rect 2454 3118 2455 3122
rect 2459 3118 2460 3122
rect 2454 3117 2460 3118
rect 2646 3122 2652 3123
rect 2646 3118 2647 3122
rect 2651 3118 2652 3122
rect 2646 3117 2652 3118
rect 2122 3095 2128 3096
rect 2122 3091 2123 3095
rect 2127 3091 2128 3095
rect 2122 3090 2128 3091
rect 2314 3095 2320 3096
rect 2314 3091 2315 3095
rect 2319 3091 2320 3095
rect 2314 3090 2320 3091
rect 2254 3084 2260 3085
rect 2254 3080 2255 3084
rect 2259 3080 2260 3084
rect 2254 3079 2260 3080
rect 2114 3067 2120 3068
rect 2114 3063 2115 3067
rect 2119 3063 2120 3067
rect 2114 3062 2120 3063
rect 2256 3051 2258 3079
rect 1871 3050 1875 3051
rect 662 3047 668 3048
rect 1830 3049 1836 3050
rect 1830 3045 1831 3049
rect 1835 3045 1836 3049
rect 1871 3045 1875 3046
rect 1895 3050 1899 3051
rect 1895 3045 1899 3046
rect 2063 3050 2067 3051
rect 2063 3045 2067 3046
rect 2199 3050 2203 3051
rect 2199 3045 2203 3046
rect 2255 3050 2259 3051
rect 2255 3045 2259 3046
rect 1830 3044 1836 3045
rect 506 3043 512 3044
rect 506 3039 507 3043
rect 511 3039 512 3043
rect 506 3038 512 3039
rect 618 3043 624 3044
rect 618 3039 619 3043
rect 623 3039 624 3043
rect 618 3038 624 3039
rect 498 3035 504 3036
rect 498 3031 499 3035
rect 503 3031 504 3035
rect 498 3030 504 3031
rect 446 3014 452 3015
rect 446 3010 447 3014
rect 451 3010 452 3014
rect 446 3009 452 3010
rect 358 3003 364 3004
rect 358 2999 359 3003
rect 363 2999 364 3003
rect 358 2998 364 2999
rect 448 2987 450 3009
rect 508 3004 510 3038
rect 558 3014 564 3015
rect 558 3010 559 3014
rect 563 3010 564 3014
rect 558 3009 564 3010
rect 506 3003 512 3004
rect 506 2999 507 3003
rect 511 2999 512 3003
rect 506 2998 512 2999
rect 560 2987 562 3009
rect 620 3004 622 3038
rect 1830 3032 1836 3033
rect 1830 3028 1831 3032
rect 1835 3028 1836 3032
rect 1830 3027 1836 3028
rect 670 3014 676 3015
rect 670 3010 671 3014
rect 675 3010 676 3014
rect 670 3009 676 3010
rect 618 3003 624 3004
rect 618 2999 619 3003
rect 623 2999 624 3003
rect 618 2998 624 2999
rect 672 2987 674 3009
rect 806 3003 812 3004
rect 806 2999 807 3003
rect 811 2999 812 3003
rect 806 2998 812 2999
rect 231 2986 235 2987
rect 231 2981 235 2982
rect 319 2986 323 2987
rect 319 2981 323 2982
rect 335 2986 339 2987
rect 335 2981 339 2982
rect 447 2986 451 2987
rect 447 2981 451 2982
rect 487 2986 491 2987
rect 487 2981 491 2982
rect 559 2986 563 2987
rect 559 2981 563 2982
rect 647 2986 651 2987
rect 647 2981 651 2982
rect 671 2986 675 2987
rect 671 2981 675 2982
rect 799 2986 803 2987
rect 799 2981 803 2982
rect 194 2979 200 2980
rect 194 2975 195 2979
rect 199 2975 200 2979
rect 194 2974 200 2975
rect 210 2979 216 2980
rect 210 2975 211 2979
rect 215 2975 216 2979
rect 210 2974 216 2975
rect 158 2970 164 2971
rect 158 2966 159 2970
rect 163 2966 164 2970
rect 158 2965 164 2966
rect 110 2952 116 2953
rect 110 2948 111 2952
rect 115 2948 116 2952
rect 110 2947 116 2948
rect 212 2944 214 2974
rect 320 2971 322 2981
rect 488 2971 490 2981
rect 530 2979 536 2980
rect 530 2975 531 2979
rect 535 2975 536 2979
rect 530 2974 536 2975
rect 538 2979 544 2980
rect 538 2975 539 2979
rect 543 2975 544 2979
rect 538 2974 544 2975
rect 318 2970 324 2971
rect 318 2966 319 2970
rect 323 2966 324 2970
rect 318 2965 324 2966
rect 486 2970 492 2971
rect 486 2966 487 2970
rect 491 2966 492 2970
rect 486 2965 492 2966
rect 210 2943 216 2944
rect 210 2939 211 2943
rect 215 2939 216 2943
rect 210 2938 216 2939
rect 342 2943 348 2944
rect 342 2939 343 2943
rect 347 2939 348 2943
rect 342 2938 348 2939
rect 110 2935 116 2936
rect 110 2931 111 2935
rect 115 2931 116 2935
rect 110 2930 116 2931
rect 150 2932 156 2933
rect 112 2911 114 2930
rect 150 2928 151 2932
rect 155 2928 156 2932
rect 150 2927 156 2928
rect 310 2932 316 2933
rect 310 2928 311 2932
rect 315 2928 316 2932
rect 310 2927 316 2928
rect 152 2911 154 2927
rect 312 2911 314 2927
rect 111 2910 115 2911
rect 111 2905 115 2906
rect 151 2910 155 2911
rect 151 2905 155 2906
rect 311 2910 315 2911
rect 311 2905 315 2906
rect 112 2886 114 2905
rect 152 2889 154 2905
rect 312 2889 314 2905
rect 150 2888 156 2889
rect 110 2885 116 2886
rect 110 2881 111 2885
rect 115 2881 116 2885
rect 150 2884 151 2888
rect 155 2884 156 2888
rect 150 2883 156 2884
rect 310 2888 316 2889
rect 310 2884 311 2888
rect 315 2884 316 2888
rect 310 2883 316 2884
rect 110 2880 116 2881
rect 218 2879 224 2880
rect 150 2875 156 2876
rect 150 2871 151 2875
rect 155 2871 156 2875
rect 218 2875 219 2879
rect 223 2875 224 2879
rect 218 2874 224 2875
rect 150 2870 156 2871
rect 110 2868 116 2869
rect 110 2864 111 2868
rect 115 2864 116 2868
rect 110 2863 116 2864
rect 112 2831 114 2863
rect 111 2830 115 2831
rect 111 2825 115 2826
rect 143 2830 147 2831
rect 143 2825 147 2826
rect 112 2797 114 2825
rect 144 2815 146 2825
rect 152 2824 154 2870
rect 158 2850 164 2851
rect 158 2846 159 2850
rect 163 2846 164 2850
rect 158 2845 164 2846
rect 160 2831 162 2845
rect 220 2840 222 2874
rect 318 2850 324 2851
rect 318 2846 319 2850
rect 323 2846 324 2850
rect 318 2845 324 2846
rect 218 2839 224 2840
rect 218 2835 219 2839
rect 223 2835 224 2839
rect 218 2834 224 2835
rect 320 2831 322 2845
rect 344 2840 346 2938
rect 478 2932 484 2933
rect 478 2928 479 2932
rect 483 2928 484 2932
rect 478 2927 484 2928
rect 480 2911 482 2927
rect 471 2910 475 2911
rect 471 2905 475 2906
rect 479 2910 483 2911
rect 479 2905 483 2906
rect 472 2889 474 2905
rect 470 2888 476 2889
rect 470 2884 471 2888
rect 475 2884 476 2888
rect 470 2883 476 2884
rect 532 2872 534 2974
rect 540 2944 542 2974
rect 648 2971 650 2981
rect 698 2979 704 2980
rect 698 2975 699 2979
rect 703 2975 704 2979
rect 698 2974 704 2975
rect 646 2970 652 2971
rect 646 2966 647 2970
rect 651 2966 652 2970
rect 646 2965 652 2966
rect 700 2944 702 2974
rect 800 2971 802 2981
rect 798 2970 804 2971
rect 798 2966 799 2970
rect 803 2966 804 2970
rect 798 2965 804 2966
rect 808 2944 810 2998
rect 1262 2987 1268 2988
rect 1832 2987 1834 3027
rect 1872 3026 1874 3045
rect 2200 3029 2202 3045
rect 2198 3028 2204 3029
rect 1870 3025 1876 3026
rect 1870 3021 1871 3025
rect 1875 3021 1876 3025
rect 2198 3024 2199 3028
rect 2203 3024 2204 3028
rect 2198 3023 2204 3024
rect 1870 3020 1876 3021
rect 2258 3011 2264 3012
rect 1870 3008 1876 3009
rect 1870 3004 1871 3008
rect 1875 3004 1876 3008
rect 2258 3007 2259 3011
rect 2263 3007 2264 3011
rect 2258 3006 2264 3007
rect 2266 3011 2272 3012
rect 2266 3007 2267 3011
rect 2271 3007 2272 3011
rect 2266 3006 2272 3007
rect 1870 3003 1876 3004
rect 943 2986 947 2987
rect 943 2981 947 2982
rect 1079 2986 1083 2987
rect 1079 2981 1083 2982
rect 1199 2986 1203 2987
rect 1262 2983 1263 2987
rect 1267 2983 1268 2987
rect 1262 2982 1268 2983
rect 1311 2986 1315 2987
rect 1199 2981 1203 2982
rect 944 2971 946 2981
rect 1070 2979 1076 2980
rect 1070 2975 1071 2979
rect 1075 2975 1076 2979
rect 1070 2974 1076 2975
rect 942 2970 948 2971
rect 942 2966 943 2970
rect 947 2966 948 2970
rect 942 2965 948 2966
rect 1072 2944 1074 2974
rect 1080 2971 1082 2981
rect 1130 2979 1136 2980
rect 1130 2975 1131 2979
rect 1135 2975 1136 2979
rect 1130 2974 1136 2975
rect 1078 2970 1084 2971
rect 1078 2966 1079 2970
rect 1083 2966 1084 2970
rect 1078 2965 1084 2966
rect 1132 2944 1134 2974
rect 1200 2971 1202 2981
rect 1250 2979 1256 2980
rect 1250 2975 1251 2979
rect 1255 2975 1256 2979
rect 1250 2974 1256 2975
rect 1198 2970 1204 2971
rect 1198 2966 1199 2970
rect 1203 2966 1204 2970
rect 1198 2965 1204 2966
rect 1252 2944 1254 2974
rect 538 2943 544 2944
rect 538 2939 539 2943
rect 543 2939 544 2943
rect 538 2938 544 2939
rect 698 2943 704 2944
rect 698 2939 699 2943
rect 703 2939 704 2943
rect 698 2938 704 2939
rect 806 2943 812 2944
rect 806 2939 807 2943
rect 811 2939 812 2943
rect 806 2938 812 2939
rect 1070 2943 1076 2944
rect 1070 2939 1071 2943
rect 1075 2939 1076 2943
rect 1070 2938 1076 2939
rect 1130 2943 1136 2944
rect 1130 2939 1131 2943
rect 1135 2939 1136 2943
rect 1130 2938 1136 2939
rect 1250 2943 1256 2944
rect 1250 2939 1251 2943
rect 1255 2939 1256 2943
rect 1250 2938 1256 2939
rect 638 2932 644 2933
rect 638 2928 639 2932
rect 643 2928 644 2932
rect 638 2927 644 2928
rect 790 2932 796 2933
rect 790 2928 791 2932
rect 795 2928 796 2932
rect 790 2927 796 2928
rect 934 2932 940 2933
rect 934 2928 935 2932
rect 939 2928 940 2932
rect 934 2927 940 2928
rect 1070 2932 1076 2933
rect 1070 2928 1071 2932
rect 1075 2928 1076 2932
rect 1070 2927 1076 2928
rect 1190 2932 1196 2933
rect 1190 2928 1191 2932
rect 1195 2928 1196 2932
rect 1190 2927 1196 2928
rect 640 2911 642 2927
rect 792 2911 794 2927
rect 936 2911 938 2927
rect 1072 2911 1074 2927
rect 1192 2911 1194 2927
rect 631 2910 635 2911
rect 631 2905 635 2906
rect 639 2910 643 2911
rect 639 2905 643 2906
rect 783 2910 787 2911
rect 783 2905 787 2906
rect 791 2910 795 2911
rect 791 2905 795 2906
rect 927 2910 931 2911
rect 927 2905 931 2906
rect 935 2910 939 2911
rect 935 2905 939 2906
rect 1055 2910 1059 2911
rect 1055 2905 1059 2906
rect 1071 2910 1075 2911
rect 1071 2905 1075 2906
rect 1175 2910 1179 2911
rect 1175 2905 1179 2906
rect 1191 2910 1195 2911
rect 1191 2905 1195 2906
rect 632 2889 634 2905
rect 784 2889 786 2905
rect 928 2889 930 2905
rect 1056 2889 1058 2905
rect 1176 2889 1178 2905
rect 630 2888 636 2889
rect 630 2884 631 2888
rect 635 2884 636 2888
rect 630 2883 636 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 926 2888 932 2889
rect 926 2884 927 2888
rect 931 2884 932 2888
rect 926 2883 932 2884
rect 1054 2888 1060 2889
rect 1054 2884 1055 2888
rect 1059 2884 1060 2888
rect 1054 2883 1060 2884
rect 1174 2888 1180 2889
rect 1174 2884 1175 2888
rect 1179 2884 1180 2888
rect 1174 2883 1180 2884
rect 1264 2880 1266 2982
rect 1311 2981 1315 2982
rect 1423 2986 1427 2987
rect 1423 2981 1427 2982
rect 1535 2986 1539 2987
rect 1535 2981 1539 2982
rect 1647 2986 1651 2987
rect 1647 2981 1651 2982
rect 1831 2986 1835 2987
rect 1831 2981 1835 2982
rect 1312 2971 1314 2981
rect 1362 2979 1368 2980
rect 1362 2975 1363 2979
rect 1367 2975 1368 2979
rect 1362 2974 1368 2975
rect 1310 2970 1316 2971
rect 1310 2966 1311 2970
rect 1315 2966 1316 2970
rect 1310 2965 1316 2966
rect 1364 2944 1366 2974
rect 1424 2971 1426 2981
rect 1474 2979 1480 2980
rect 1474 2975 1475 2979
rect 1479 2975 1480 2979
rect 1474 2974 1480 2975
rect 1422 2970 1428 2971
rect 1422 2966 1423 2970
rect 1427 2966 1428 2970
rect 1422 2965 1428 2966
rect 1476 2944 1478 2974
rect 1536 2971 1538 2981
rect 1586 2979 1592 2980
rect 1586 2975 1587 2979
rect 1591 2975 1592 2979
rect 1586 2974 1592 2975
rect 1534 2970 1540 2971
rect 1534 2966 1535 2970
rect 1539 2966 1540 2970
rect 1534 2965 1540 2966
rect 1588 2944 1590 2974
rect 1648 2971 1650 2981
rect 1646 2970 1652 2971
rect 1646 2966 1647 2970
rect 1651 2966 1652 2970
rect 1646 2965 1652 2966
rect 1832 2953 1834 2981
rect 1872 2963 1874 3003
rect 2206 2990 2212 2991
rect 2206 2986 2207 2990
rect 2211 2986 2212 2990
rect 2206 2985 2212 2986
rect 2208 2963 2210 2985
rect 1871 2962 1875 2963
rect 1871 2957 1875 2958
rect 2127 2962 2131 2963
rect 2127 2957 2131 2958
rect 2207 2962 2211 2963
rect 2207 2957 2211 2958
rect 1830 2952 1836 2953
rect 1830 2948 1831 2952
rect 1835 2948 1836 2952
rect 1830 2947 1836 2948
rect 1362 2943 1368 2944
rect 1362 2939 1363 2943
rect 1367 2939 1368 2943
rect 1362 2938 1368 2939
rect 1474 2943 1480 2944
rect 1474 2939 1475 2943
rect 1479 2939 1480 2943
rect 1474 2938 1480 2939
rect 1586 2943 1592 2944
rect 1586 2939 1587 2943
rect 1591 2939 1592 2943
rect 1586 2938 1592 2939
rect 1830 2935 1836 2936
rect 1302 2932 1308 2933
rect 1302 2928 1303 2932
rect 1307 2928 1308 2932
rect 1302 2927 1308 2928
rect 1414 2932 1420 2933
rect 1414 2928 1415 2932
rect 1419 2928 1420 2932
rect 1414 2927 1420 2928
rect 1526 2932 1532 2933
rect 1526 2928 1527 2932
rect 1531 2928 1532 2932
rect 1526 2927 1532 2928
rect 1638 2932 1644 2933
rect 1638 2928 1639 2932
rect 1643 2928 1644 2932
rect 1830 2931 1831 2935
rect 1835 2931 1836 2935
rect 1830 2930 1836 2931
rect 1638 2927 1644 2928
rect 1304 2911 1306 2927
rect 1416 2911 1418 2927
rect 1426 2915 1432 2916
rect 1426 2911 1427 2915
rect 1431 2911 1432 2915
rect 1528 2911 1530 2927
rect 1640 2911 1642 2927
rect 1832 2911 1834 2930
rect 1872 2929 1874 2957
rect 2128 2947 2130 2957
rect 2208 2947 2210 2957
rect 2260 2956 2262 3006
rect 2268 2980 2270 3006
rect 2316 2980 2318 3090
rect 2446 3084 2452 3085
rect 2446 3080 2447 3084
rect 2451 3080 2452 3084
rect 2446 3079 2452 3080
rect 2638 3084 2644 3085
rect 2638 3080 2639 3084
rect 2643 3080 2644 3084
rect 2638 3079 2644 3080
rect 2448 3051 2450 3079
rect 2640 3051 2642 3079
rect 2335 3050 2339 3051
rect 2335 3045 2339 3046
rect 2447 3050 2451 3051
rect 2447 3045 2451 3046
rect 2479 3050 2483 3051
rect 2479 3045 2483 3046
rect 2623 3050 2627 3051
rect 2623 3045 2627 3046
rect 2639 3050 2643 3051
rect 2639 3045 2643 3046
rect 2336 3029 2338 3045
rect 2480 3029 2482 3045
rect 2624 3029 2626 3045
rect 2334 3028 2340 3029
rect 2334 3024 2335 3028
rect 2339 3024 2340 3028
rect 2334 3023 2340 3024
rect 2478 3028 2484 3029
rect 2478 3024 2479 3028
rect 2483 3024 2484 3028
rect 2478 3023 2484 3024
rect 2622 3028 2628 3029
rect 2622 3024 2623 3028
rect 2627 3024 2628 3028
rect 2622 3023 2628 3024
rect 2426 3019 2432 3020
rect 2426 3015 2427 3019
rect 2431 3015 2432 3019
rect 2426 3014 2432 3015
rect 2342 2990 2348 2991
rect 2342 2986 2343 2990
rect 2347 2986 2348 2990
rect 2342 2985 2348 2986
rect 2266 2979 2272 2980
rect 2266 2975 2267 2979
rect 2271 2975 2272 2979
rect 2266 2974 2272 2975
rect 2314 2979 2320 2980
rect 2314 2975 2315 2979
rect 2319 2975 2320 2979
rect 2314 2974 2320 2975
rect 2344 2963 2346 2985
rect 2428 2980 2430 3014
rect 2684 3012 2686 3126
rect 2700 3096 2702 3126
rect 2832 3123 2834 3133
rect 2830 3122 2836 3123
rect 2830 3118 2831 3122
rect 2835 3118 2836 3122
rect 2830 3117 2836 3118
rect 3008 3096 3010 3138
rect 3015 3133 3019 3134
rect 3159 3138 3163 3139
rect 3159 3133 3163 3134
rect 3199 3138 3203 3139
rect 3210 3138 3216 3139
rect 3262 3143 3268 3144
rect 3262 3139 3263 3143
rect 3267 3139 3268 3143
rect 3336 3139 3338 3149
rect 3262 3138 3268 3139
rect 3335 3138 3339 3139
rect 3199 3133 3203 3134
rect 3335 3133 3339 3134
rect 3391 3138 3395 3139
rect 3391 3133 3395 3134
rect 3016 3123 3018 3133
rect 3042 3131 3048 3132
rect 3042 3127 3043 3131
rect 3047 3127 3048 3131
rect 3042 3126 3048 3127
rect 3066 3131 3072 3132
rect 3066 3127 3067 3131
rect 3071 3127 3072 3131
rect 3066 3126 3072 3127
rect 3014 3122 3020 3123
rect 3014 3118 3015 3122
rect 3019 3118 3020 3122
rect 3014 3117 3020 3118
rect 2698 3095 2704 3096
rect 2698 3091 2699 3095
rect 2703 3091 2704 3095
rect 2698 3090 2704 3091
rect 3006 3095 3012 3096
rect 3006 3091 3007 3095
rect 3011 3091 3012 3095
rect 3006 3090 3012 3091
rect 2822 3084 2828 3085
rect 2822 3080 2823 3084
rect 2827 3080 2828 3084
rect 2822 3079 2828 3080
rect 3006 3084 3012 3085
rect 3006 3080 3007 3084
rect 3011 3080 3012 3084
rect 3006 3079 3012 3080
rect 2824 3051 2826 3079
rect 3008 3051 3010 3079
rect 3044 3068 3046 3126
rect 3068 3096 3070 3126
rect 3200 3123 3202 3133
rect 3392 3123 3394 3133
rect 3400 3132 3402 3178
rect 3510 3154 3516 3155
rect 3510 3150 3511 3154
rect 3515 3150 3516 3154
rect 3510 3149 3516 3150
rect 3512 3139 3514 3149
rect 3536 3144 3538 3242
rect 3590 3239 3596 3240
rect 3590 3235 3591 3239
rect 3595 3235 3596 3239
rect 3590 3234 3596 3235
rect 3592 3215 3594 3234
rect 3591 3214 3595 3215
rect 3591 3209 3595 3210
rect 3592 3190 3594 3209
rect 3590 3189 3596 3190
rect 3590 3185 3591 3189
rect 3595 3185 3596 3189
rect 3590 3184 3596 3185
rect 3590 3172 3596 3173
rect 3590 3168 3591 3172
rect 3595 3168 3596 3172
rect 3590 3167 3596 3168
rect 3534 3143 3540 3144
rect 3534 3139 3535 3143
rect 3539 3139 3540 3143
rect 3592 3139 3594 3167
rect 3511 3138 3515 3139
rect 3534 3138 3540 3139
rect 3591 3138 3595 3139
rect 3511 3133 3515 3134
rect 3591 3133 3595 3134
rect 3398 3131 3404 3132
rect 3398 3127 3399 3131
rect 3403 3127 3404 3131
rect 3398 3126 3404 3127
rect 3198 3122 3204 3123
rect 3198 3118 3199 3122
rect 3203 3118 3204 3122
rect 3198 3117 3204 3118
rect 3390 3122 3396 3123
rect 3390 3118 3391 3122
rect 3395 3118 3396 3122
rect 3390 3117 3396 3118
rect 3592 3105 3594 3133
rect 3590 3104 3596 3105
rect 3590 3100 3591 3104
rect 3595 3100 3596 3104
rect 3590 3099 3596 3100
rect 3066 3095 3072 3096
rect 3066 3091 3067 3095
rect 3071 3091 3072 3095
rect 3066 3090 3072 3091
rect 3282 3095 3288 3096
rect 3282 3091 3283 3095
rect 3287 3091 3288 3095
rect 3282 3090 3288 3091
rect 3190 3084 3196 3085
rect 3190 3080 3191 3084
rect 3195 3080 3196 3084
rect 3190 3079 3196 3080
rect 3042 3067 3048 3068
rect 3042 3063 3043 3067
rect 3047 3063 3048 3067
rect 3042 3062 3048 3063
rect 3192 3051 3194 3079
rect 2767 3050 2771 3051
rect 2767 3045 2771 3046
rect 2823 3050 2827 3051
rect 2823 3045 2827 3046
rect 2903 3050 2907 3051
rect 2903 3045 2907 3046
rect 3007 3050 3011 3051
rect 3007 3045 3011 3046
rect 3039 3050 3043 3051
rect 3039 3045 3043 3046
rect 3183 3050 3187 3051
rect 3183 3045 3187 3046
rect 3191 3050 3195 3051
rect 3191 3045 3195 3046
rect 2768 3029 2770 3045
rect 2904 3029 2906 3045
rect 3040 3029 3042 3045
rect 3184 3029 3186 3045
rect 2766 3028 2772 3029
rect 2766 3024 2767 3028
rect 2771 3024 2772 3028
rect 2766 3023 2772 3024
rect 2902 3028 2908 3029
rect 2902 3024 2903 3028
rect 2907 3024 2908 3028
rect 2902 3023 2908 3024
rect 3038 3028 3044 3029
rect 3038 3024 3039 3028
rect 3043 3024 3044 3028
rect 3038 3023 3044 3024
rect 3182 3028 3188 3029
rect 3182 3024 3183 3028
rect 3187 3024 3188 3028
rect 3182 3023 3188 3024
rect 2690 3019 2696 3020
rect 2690 3015 2691 3019
rect 2695 3015 2696 3019
rect 2690 3014 2696 3015
rect 2834 3019 2840 3020
rect 2834 3015 2835 3019
rect 2839 3015 2840 3019
rect 2834 3014 2840 3015
rect 3106 3019 3112 3020
rect 3106 3015 3107 3019
rect 3111 3015 3112 3019
rect 3106 3014 3112 3015
rect 3250 3019 3256 3020
rect 3250 3015 3251 3019
rect 3255 3015 3256 3019
rect 3250 3014 3256 3015
rect 2682 3011 2688 3012
rect 2682 3007 2683 3011
rect 2687 3007 2688 3011
rect 2682 3006 2688 3007
rect 2486 2990 2492 2991
rect 2486 2986 2487 2990
rect 2491 2986 2492 2990
rect 2486 2985 2492 2986
rect 2630 2990 2636 2991
rect 2630 2986 2631 2990
rect 2635 2986 2636 2990
rect 2630 2985 2636 2986
rect 2426 2979 2432 2980
rect 2426 2975 2427 2979
rect 2431 2975 2432 2979
rect 2426 2974 2432 2975
rect 2488 2963 2490 2985
rect 2632 2963 2634 2985
rect 2692 2980 2694 3014
rect 2774 2990 2780 2991
rect 2774 2986 2775 2990
rect 2779 2986 2780 2990
rect 2774 2985 2780 2986
rect 2690 2979 2696 2980
rect 2690 2975 2691 2979
rect 2695 2975 2696 2979
rect 2690 2974 2696 2975
rect 2776 2963 2778 2985
rect 2836 2980 2838 3014
rect 3098 3011 3104 3012
rect 3098 3007 3099 3011
rect 3103 3007 3104 3011
rect 3098 3006 3104 3007
rect 2910 2990 2916 2991
rect 2910 2986 2911 2990
rect 2915 2986 2916 2990
rect 2910 2985 2916 2986
rect 3046 2990 3052 2991
rect 3046 2986 3047 2990
rect 3051 2986 3052 2990
rect 3046 2985 3052 2986
rect 2834 2979 2840 2980
rect 2834 2975 2835 2979
rect 2839 2975 2840 2979
rect 2834 2974 2840 2975
rect 2912 2963 2914 2985
rect 3048 2963 3050 2985
rect 2287 2962 2291 2963
rect 2287 2957 2291 2958
rect 2343 2962 2347 2963
rect 2343 2957 2347 2958
rect 2367 2962 2371 2963
rect 2367 2957 2371 2958
rect 2447 2962 2451 2963
rect 2447 2957 2451 2958
rect 2487 2962 2491 2963
rect 2487 2957 2491 2958
rect 2527 2962 2531 2963
rect 2527 2957 2531 2958
rect 2607 2962 2611 2963
rect 2607 2957 2611 2958
rect 2631 2962 2635 2963
rect 2631 2957 2635 2958
rect 2695 2962 2699 2963
rect 2695 2957 2699 2958
rect 2775 2962 2779 2963
rect 2775 2957 2779 2958
rect 2791 2962 2795 2963
rect 2791 2957 2795 2958
rect 2911 2962 2915 2963
rect 2911 2957 2915 2958
rect 3039 2962 3043 2963
rect 3039 2957 3043 2958
rect 3047 2962 3051 2963
rect 3047 2957 3051 2958
rect 2214 2955 2220 2956
rect 2214 2951 2215 2955
rect 2219 2951 2220 2955
rect 2214 2950 2220 2951
rect 2258 2955 2264 2956
rect 2258 2951 2259 2955
rect 2263 2951 2264 2955
rect 2258 2950 2264 2951
rect 2126 2946 2132 2947
rect 2126 2942 2127 2946
rect 2131 2942 2132 2946
rect 2126 2941 2132 2942
rect 2206 2946 2212 2947
rect 2206 2942 2207 2946
rect 2211 2942 2212 2946
rect 2206 2941 2212 2942
rect 1870 2928 1876 2929
rect 1870 2924 1871 2928
rect 1875 2924 1876 2928
rect 1870 2923 1876 2924
rect 2216 2920 2218 2950
rect 2288 2947 2290 2957
rect 2314 2955 2320 2956
rect 2314 2951 2315 2955
rect 2319 2951 2320 2955
rect 2314 2950 2320 2951
rect 2350 2955 2356 2956
rect 2350 2951 2351 2955
rect 2355 2951 2356 2955
rect 2350 2950 2356 2951
rect 2286 2946 2292 2947
rect 2286 2942 2287 2946
rect 2291 2942 2292 2946
rect 2286 2941 2292 2942
rect 2214 2919 2220 2920
rect 2214 2915 2215 2919
rect 2219 2915 2220 2919
rect 2214 2914 2220 2915
rect 1870 2911 1876 2912
rect 1287 2910 1291 2911
rect 1287 2905 1291 2906
rect 1303 2910 1307 2911
rect 1303 2905 1307 2906
rect 1391 2910 1395 2911
rect 1391 2905 1395 2906
rect 1415 2910 1419 2911
rect 1426 2910 1432 2911
rect 1487 2910 1491 2911
rect 1415 2905 1419 2906
rect 1288 2889 1290 2905
rect 1392 2889 1394 2905
rect 1286 2888 1292 2889
rect 1286 2884 1287 2888
rect 1291 2884 1292 2888
rect 1286 2883 1292 2884
rect 1390 2888 1396 2889
rect 1390 2884 1391 2888
rect 1395 2884 1396 2888
rect 1390 2883 1396 2884
rect 538 2879 544 2880
rect 538 2875 539 2879
rect 543 2875 544 2879
rect 538 2874 544 2875
rect 698 2879 704 2880
rect 698 2875 699 2879
rect 703 2875 704 2879
rect 698 2874 704 2875
rect 1014 2879 1020 2880
rect 1014 2875 1015 2879
rect 1019 2875 1020 2879
rect 1014 2874 1020 2875
rect 1122 2879 1128 2880
rect 1122 2875 1123 2879
rect 1127 2875 1128 2879
rect 1122 2874 1128 2875
rect 1254 2879 1260 2880
rect 1254 2875 1255 2879
rect 1259 2875 1260 2879
rect 1254 2874 1260 2875
rect 1262 2879 1268 2880
rect 1262 2875 1263 2879
rect 1267 2875 1268 2879
rect 1262 2874 1268 2875
rect 530 2871 536 2872
rect 530 2867 531 2871
rect 535 2867 536 2871
rect 530 2866 536 2867
rect 478 2850 484 2851
rect 478 2846 479 2850
rect 483 2846 484 2850
rect 478 2845 484 2846
rect 342 2839 348 2840
rect 342 2835 343 2839
rect 347 2835 348 2839
rect 342 2834 348 2835
rect 480 2831 482 2845
rect 540 2840 542 2874
rect 638 2850 644 2851
rect 638 2846 639 2850
rect 643 2846 644 2850
rect 638 2845 644 2846
rect 538 2839 544 2840
rect 538 2835 539 2839
rect 543 2835 544 2839
rect 538 2834 544 2835
rect 640 2831 642 2845
rect 700 2840 702 2874
rect 790 2850 796 2851
rect 790 2846 791 2850
rect 795 2846 796 2850
rect 790 2845 796 2846
rect 934 2850 940 2851
rect 934 2846 935 2850
rect 939 2846 940 2850
rect 934 2845 940 2846
rect 698 2839 704 2840
rect 698 2835 699 2839
rect 703 2835 704 2839
rect 698 2834 704 2835
rect 792 2831 794 2845
rect 854 2839 860 2840
rect 854 2835 855 2839
rect 859 2835 860 2839
rect 854 2834 860 2835
rect 159 2830 163 2831
rect 159 2825 163 2826
rect 247 2830 251 2831
rect 247 2825 251 2826
rect 319 2830 323 2831
rect 319 2825 323 2826
rect 383 2830 387 2831
rect 383 2825 387 2826
rect 479 2830 483 2831
rect 479 2825 483 2826
rect 535 2830 539 2831
rect 535 2825 539 2826
rect 639 2830 643 2831
rect 639 2825 643 2826
rect 687 2830 691 2831
rect 687 2825 691 2826
rect 791 2830 795 2831
rect 791 2825 795 2826
rect 847 2830 851 2831
rect 847 2825 851 2826
rect 150 2823 156 2824
rect 150 2819 151 2823
rect 155 2819 156 2823
rect 150 2818 156 2819
rect 194 2823 200 2824
rect 194 2819 195 2823
rect 199 2819 200 2823
rect 194 2818 200 2819
rect 142 2814 148 2815
rect 142 2810 143 2814
rect 147 2810 148 2814
rect 142 2809 148 2810
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 196 2788 198 2818
rect 248 2815 250 2825
rect 298 2823 304 2824
rect 298 2819 299 2823
rect 303 2819 304 2823
rect 298 2818 304 2819
rect 246 2814 252 2815
rect 246 2810 247 2814
rect 251 2810 252 2814
rect 246 2809 252 2810
rect 300 2788 302 2818
rect 384 2815 386 2825
rect 536 2815 538 2825
rect 570 2823 576 2824
rect 570 2819 571 2823
rect 575 2819 576 2823
rect 570 2818 576 2819
rect 586 2823 592 2824
rect 586 2819 587 2823
rect 591 2819 592 2823
rect 586 2818 592 2819
rect 382 2814 388 2815
rect 382 2810 383 2814
rect 387 2810 388 2814
rect 382 2809 388 2810
rect 534 2814 540 2815
rect 534 2810 535 2814
rect 539 2810 540 2814
rect 534 2809 540 2810
rect 194 2787 200 2788
rect 194 2783 195 2787
rect 199 2783 200 2787
rect 194 2782 200 2783
rect 298 2787 304 2788
rect 298 2783 299 2787
rect 303 2783 304 2787
rect 298 2782 304 2783
rect 110 2779 116 2780
rect 110 2775 111 2779
rect 115 2775 116 2779
rect 110 2774 116 2775
rect 134 2776 140 2777
rect 112 2751 114 2774
rect 134 2772 135 2776
rect 139 2772 140 2776
rect 134 2771 140 2772
rect 238 2776 244 2777
rect 238 2772 239 2776
rect 243 2772 244 2776
rect 238 2771 244 2772
rect 374 2776 380 2777
rect 374 2772 375 2776
rect 379 2772 380 2776
rect 374 2771 380 2772
rect 526 2776 532 2777
rect 526 2772 527 2776
rect 531 2772 532 2776
rect 526 2771 532 2772
rect 136 2751 138 2771
rect 240 2751 242 2771
rect 376 2751 378 2771
rect 394 2759 400 2760
rect 394 2755 395 2759
rect 399 2755 400 2759
rect 394 2754 400 2755
rect 111 2750 115 2751
rect 111 2745 115 2746
rect 135 2750 139 2751
rect 135 2745 139 2746
rect 231 2750 235 2751
rect 231 2745 235 2746
rect 239 2750 243 2751
rect 239 2745 243 2746
rect 367 2750 371 2751
rect 367 2745 371 2746
rect 375 2750 379 2751
rect 375 2745 379 2746
rect 112 2726 114 2745
rect 136 2729 138 2745
rect 232 2729 234 2745
rect 368 2729 370 2745
rect 134 2728 140 2729
rect 110 2725 116 2726
rect 110 2721 111 2725
rect 115 2721 116 2725
rect 134 2724 135 2728
rect 139 2724 140 2728
rect 134 2723 140 2724
rect 230 2728 236 2729
rect 230 2724 231 2728
rect 235 2724 236 2728
rect 230 2723 236 2724
rect 366 2728 372 2729
rect 366 2724 367 2728
rect 371 2724 372 2728
rect 366 2723 372 2724
rect 110 2720 116 2721
rect 202 2719 208 2720
rect 202 2715 203 2719
rect 207 2715 208 2719
rect 202 2714 208 2715
rect 298 2719 304 2720
rect 298 2715 299 2719
rect 303 2715 304 2719
rect 298 2714 304 2715
rect 194 2711 200 2712
rect 110 2708 116 2709
rect 110 2704 111 2708
rect 115 2704 116 2708
rect 194 2707 195 2711
rect 199 2707 200 2711
rect 194 2706 200 2707
rect 110 2703 116 2704
rect 112 2667 114 2703
rect 142 2690 148 2691
rect 142 2686 143 2690
rect 147 2686 148 2690
rect 142 2685 148 2686
rect 144 2667 146 2685
rect 111 2666 115 2667
rect 111 2661 115 2662
rect 143 2666 147 2667
rect 143 2661 147 2662
rect 112 2633 114 2661
rect 144 2651 146 2661
rect 196 2660 198 2706
rect 204 2680 206 2714
rect 238 2690 244 2691
rect 238 2686 239 2690
rect 243 2686 244 2690
rect 238 2685 244 2686
rect 202 2679 208 2680
rect 202 2675 203 2679
rect 207 2675 208 2679
rect 202 2674 208 2675
rect 240 2667 242 2685
rect 300 2680 302 2714
rect 374 2690 380 2691
rect 374 2686 375 2690
rect 379 2686 380 2690
rect 374 2685 380 2686
rect 298 2679 304 2680
rect 298 2675 299 2679
rect 303 2675 304 2679
rect 298 2674 304 2675
rect 376 2667 378 2685
rect 396 2680 398 2754
rect 528 2751 530 2771
rect 511 2750 515 2751
rect 511 2745 515 2746
rect 527 2750 531 2751
rect 527 2745 531 2746
rect 512 2729 514 2745
rect 510 2728 516 2729
rect 510 2724 511 2728
rect 515 2724 516 2728
rect 510 2723 516 2724
rect 572 2712 574 2818
rect 588 2788 590 2818
rect 688 2815 690 2825
rect 738 2823 744 2824
rect 738 2819 739 2823
rect 743 2819 744 2823
rect 738 2818 744 2819
rect 686 2814 692 2815
rect 686 2810 687 2814
rect 691 2810 692 2814
rect 686 2809 692 2810
rect 740 2788 742 2818
rect 848 2815 850 2825
rect 846 2814 852 2815
rect 846 2810 847 2814
rect 851 2810 852 2814
rect 846 2809 852 2810
rect 856 2788 858 2834
rect 936 2831 938 2845
rect 1016 2840 1018 2874
rect 1062 2850 1068 2851
rect 1062 2846 1063 2850
rect 1067 2846 1068 2850
rect 1062 2845 1068 2846
rect 1006 2839 1012 2840
rect 1006 2835 1007 2839
rect 1011 2835 1012 2839
rect 1006 2834 1012 2835
rect 1014 2839 1020 2840
rect 1014 2835 1015 2839
rect 1019 2835 1020 2839
rect 1014 2834 1020 2835
rect 935 2830 939 2831
rect 935 2825 939 2826
rect 999 2830 1003 2831
rect 999 2825 1003 2826
rect 1000 2815 1002 2825
rect 998 2814 1004 2815
rect 998 2810 999 2814
rect 1003 2810 1004 2814
rect 998 2809 1004 2810
rect 1008 2788 1010 2834
rect 1064 2831 1066 2845
rect 1124 2840 1126 2874
rect 1182 2850 1188 2851
rect 1182 2846 1183 2850
rect 1187 2846 1188 2850
rect 1182 2845 1188 2846
rect 1122 2839 1128 2840
rect 1122 2835 1123 2839
rect 1127 2835 1128 2839
rect 1122 2834 1128 2835
rect 1184 2831 1186 2845
rect 1256 2840 1258 2874
rect 1294 2850 1300 2851
rect 1294 2846 1295 2850
rect 1299 2846 1300 2850
rect 1294 2845 1300 2846
rect 1398 2850 1404 2851
rect 1398 2846 1399 2850
rect 1403 2846 1404 2850
rect 1398 2845 1404 2846
rect 1254 2839 1260 2840
rect 1254 2835 1255 2839
rect 1259 2835 1260 2839
rect 1254 2834 1260 2835
rect 1286 2831 1292 2832
rect 1296 2831 1298 2845
rect 1400 2831 1402 2845
rect 1428 2840 1430 2910
rect 1487 2905 1491 2906
rect 1527 2910 1531 2911
rect 1527 2905 1531 2906
rect 1591 2910 1595 2911
rect 1591 2905 1595 2906
rect 1639 2910 1643 2911
rect 1639 2905 1643 2906
rect 1695 2910 1699 2911
rect 1695 2905 1699 2906
rect 1831 2910 1835 2911
rect 1870 2907 1871 2911
rect 1875 2907 1876 2911
rect 1870 2906 1876 2907
rect 2118 2908 2124 2909
rect 1831 2905 1835 2906
rect 1488 2889 1490 2905
rect 1592 2889 1594 2905
rect 1696 2889 1698 2905
rect 1486 2888 1492 2889
rect 1486 2884 1487 2888
rect 1491 2884 1492 2888
rect 1486 2883 1492 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1590 2883 1596 2884
rect 1694 2888 1700 2889
rect 1694 2884 1695 2888
rect 1699 2884 1700 2888
rect 1832 2886 1834 2905
rect 1872 2887 1874 2906
rect 2118 2904 2119 2908
rect 2123 2904 2124 2908
rect 2118 2903 2124 2904
rect 2198 2908 2204 2909
rect 2198 2904 2199 2908
rect 2203 2904 2204 2908
rect 2198 2903 2204 2904
rect 2278 2908 2284 2909
rect 2278 2904 2279 2908
rect 2283 2904 2284 2908
rect 2278 2903 2284 2904
rect 2082 2891 2088 2892
rect 2082 2887 2083 2891
rect 2087 2887 2088 2891
rect 2120 2887 2122 2903
rect 2200 2887 2202 2903
rect 2280 2887 2282 2903
rect 1871 2886 1875 2887
rect 1694 2883 1700 2884
rect 1830 2885 1836 2886
rect 1830 2881 1831 2885
rect 1835 2881 1836 2885
rect 1871 2881 1875 2882
rect 2047 2886 2051 2887
rect 2082 2886 2088 2887
rect 2119 2886 2123 2887
rect 2047 2881 2051 2882
rect 1830 2880 1836 2881
rect 1462 2879 1468 2880
rect 1462 2875 1463 2879
rect 1467 2875 1468 2879
rect 1462 2874 1468 2875
rect 1562 2879 1568 2880
rect 1562 2875 1563 2879
rect 1567 2875 1568 2879
rect 1562 2874 1568 2875
rect 1666 2879 1672 2880
rect 1666 2875 1667 2879
rect 1671 2875 1672 2879
rect 1666 2874 1672 2875
rect 1674 2879 1680 2880
rect 1674 2875 1675 2879
rect 1679 2875 1680 2879
rect 1674 2874 1680 2875
rect 1435 2852 1439 2853
rect 1435 2847 1439 2848
rect 1426 2839 1432 2840
rect 1426 2835 1427 2839
rect 1431 2835 1432 2839
rect 1426 2834 1432 2835
rect 1063 2830 1067 2831
rect 1063 2825 1067 2826
rect 1143 2830 1147 2831
rect 1143 2825 1147 2826
rect 1183 2830 1187 2831
rect 1183 2825 1187 2826
rect 1279 2830 1283 2831
rect 1286 2827 1287 2831
rect 1291 2827 1292 2831
rect 1286 2826 1292 2827
rect 1295 2830 1299 2831
rect 1279 2825 1283 2826
rect 1144 2815 1146 2825
rect 1202 2823 1208 2824
rect 1202 2819 1203 2823
rect 1207 2819 1208 2823
rect 1202 2818 1208 2819
rect 1230 2823 1236 2824
rect 1230 2819 1231 2823
rect 1235 2819 1236 2823
rect 1230 2818 1236 2819
rect 1142 2814 1148 2815
rect 1142 2810 1143 2814
rect 1147 2810 1148 2814
rect 1142 2809 1148 2810
rect 586 2787 592 2788
rect 586 2783 587 2787
rect 591 2783 592 2787
rect 586 2782 592 2783
rect 738 2787 744 2788
rect 738 2783 739 2787
rect 743 2783 744 2787
rect 738 2782 744 2783
rect 854 2787 860 2788
rect 854 2783 855 2787
rect 859 2783 860 2787
rect 854 2782 860 2783
rect 1006 2787 1012 2788
rect 1006 2783 1007 2787
rect 1011 2783 1012 2787
rect 1006 2782 1012 2783
rect 678 2776 684 2777
rect 678 2772 679 2776
rect 683 2772 684 2776
rect 678 2771 684 2772
rect 838 2776 844 2777
rect 838 2772 839 2776
rect 843 2772 844 2776
rect 838 2771 844 2772
rect 990 2776 996 2777
rect 990 2772 991 2776
rect 995 2772 996 2776
rect 990 2771 996 2772
rect 1134 2776 1140 2777
rect 1134 2772 1135 2776
rect 1139 2772 1140 2776
rect 1134 2771 1140 2772
rect 680 2751 682 2771
rect 840 2751 842 2771
rect 992 2751 994 2771
rect 1136 2751 1138 2771
rect 663 2750 667 2751
rect 663 2745 667 2746
rect 679 2750 683 2751
rect 679 2745 683 2746
rect 815 2750 819 2751
rect 815 2745 819 2746
rect 839 2750 843 2751
rect 839 2745 843 2746
rect 975 2750 979 2751
rect 975 2745 979 2746
rect 991 2750 995 2751
rect 991 2745 995 2746
rect 1135 2750 1139 2751
rect 1135 2745 1139 2746
rect 664 2729 666 2745
rect 816 2729 818 2745
rect 976 2729 978 2745
rect 1136 2729 1138 2745
rect 662 2728 668 2729
rect 662 2724 663 2728
rect 667 2724 668 2728
rect 662 2723 668 2724
rect 814 2728 820 2729
rect 814 2724 815 2728
rect 819 2724 820 2728
rect 814 2723 820 2724
rect 974 2728 980 2729
rect 974 2724 975 2728
rect 979 2724 980 2728
rect 974 2723 980 2724
rect 1134 2728 1140 2729
rect 1134 2724 1135 2728
rect 1139 2724 1140 2728
rect 1134 2723 1140 2724
rect 1204 2720 1206 2818
rect 1232 2788 1234 2818
rect 1280 2815 1282 2825
rect 1278 2814 1284 2815
rect 1278 2810 1279 2814
rect 1283 2810 1284 2814
rect 1278 2809 1284 2810
rect 1288 2788 1290 2826
rect 1295 2825 1299 2826
rect 1399 2830 1403 2831
rect 1399 2825 1403 2826
rect 1407 2830 1411 2831
rect 1407 2825 1411 2826
rect 1408 2815 1410 2825
rect 1436 2824 1438 2847
rect 1464 2840 1466 2874
rect 1494 2850 1500 2851
rect 1494 2846 1495 2850
rect 1499 2846 1500 2850
rect 1494 2845 1500 2846
rect 1462 2839 1468 2840
rect 1462 2835 1463 2839
rect 1467 2835 1468 2839
rect 1462 2834 1468 2835
rect 1496 2831 1498 2845
rect 1564 2840 1566 2874
rect 1598 2850 1604 2851
rect 1598 2846 1599 2850
rect 1603 2846 1604 2850
rect 1598 2845 1604 2846
rect 1562 2839 1568 2840
rect 1562 2835 1563 2839
rect 1567 2835 1568 2839
rect 1562 2834 1568 2835
rect 1600 2831 1602 2845
rect 1668 2840 1670 2874
rect 1676 2853 1678 2874
rect 1830 2868 1836 2869
rect 1830 2864 1831 2868
rect 1835 2864 1836 2868
rect 1830 2863 1836 2864
rect 1675 2852 1679 2853
rect 1675 2847 1679 2848
rect 1702 2850 1708 2851
rect 1702 2846 1703 2850
rect 1707 2846 1708 2850
rect 1702 2845 1708 2846
rect 1666 2839 1672 2840
rect 1666 2835 1667 2839
rect 1671 2835 1672 2839
rect 1666 2834 1672 2835
rect 1704 2831 1706 2845
rect 1832 2831 1834 2863
rect 1872 2862 1874 2881
rect 2048 2865 2050 2881
rect 2046 2864 2052 2865
rect 1870 2861 1876 2862
rect 1870 2857 1871 2861
rect 1875 2857 1876 2861
rect 2046 2860 2047 2864
rect 2051 2860 2052 2864
rect 2046 2859 2052 2860
rect 1870 2856 1876 2857
rect 1870 2844 1876 2845
rect 1870 2840 1871 2844
rect 1875 2840 1876 2844
rect 1870 2839 1876 2840
rect 1495 2830 1499 2831
rect 1495 2825 1499 2826
rect 1527 2830 1531 2831
rect 1527 2825 1531 2826
rect 1599 2830 1603 2831
rect 1599 2825 1603 2826
rect 1647 2830 1651 2831
rect 1647 2825 1651 2826
rect 1703 2830 1707 2831
rect 1703 2825 1707 2826
rect 1751 2830 1755 2831
rect 1751 2825 1755 2826
rect 1831 2830 1835 2831
rect 1831 2825 1835 2826
rect 1434 2823 1440 2824
rect 1434 2819 1435 2823
rect 1439 2819 1440 2823
rect 1434 2818 1440 2819
rect 1458 2823 1464 2824
rect 1458 2819 1459 2823
rect 1463 2819 1464 2823
rect 1458 2818 1464 2819
rect 1406 2814 1412 2815
rect 1406 2810 1407 2814
rect 1411 2810 1412 2814
rect 1406 2809 1412 2810
rect 1460 2788 1462 2818
rect 1528 2815 1530 2825
rect 1578 2823 1584 2824
rect 1578 2819 1579 2823
rect 1583 2819 1584 2823
rect 1578 2818 1584 2819
rect 1526 2814 1532 2815
rect 1526 2810 1527 2814
rect 1531 2810 1532 2814
rect 1526 2809 1532 2810
rect 1580 2788 1582 2818
rect 1648 2815 1650 2825
rect 1714 2823 1720 2824
rect 1714 2819 1715 2823
rect 1719 2819 1720 2823
rect 1714 2818 1720 2819
rect 1646 2814 1652 2815
rect 1646 2810 1647 2814
rect 1651 2810 1652 2814
rect 1646 2809 1652 2810
rect 1716 2788 1718 2818
rect 1752 2815 1754 2825
rect 1750 2814 1756 2815
rect 1750 2810 1751 2814
rect 1755 2810 1756 2814
rect 1750 2809 1756 2810
rect 1832 2797 1834 2825
rect 1872 2799 1874 2839
rect 2054 2826 2060 2827
rect 2054 2822 2055 2826
rect 2059 2822 2060 2826
rect 2054 2821 2060 2822
rect 2022 2799 2028 2800
rect 2056 2799 2058 2821
rect 2084 2816 2086 2886
rect 2119 2881 2123 2882
rect 2135 2886 2139 2887
rect 2135 2881 2139 2882
rect 2199 2886 2203 2887
rect 2199 2881 2203 2882
rect 2239 2886 2243 2887
rect 2239 2881 2243 2882
rect 2279 2886 2283 2887
rect 2279 2881 2283 2882
rect 2136 2865 2138 2881
rect 2240 2865 2242 2881
rect 2134 2864 2140 2865
rect 2134 2860 2135 2864
rect 2139 2860 2140 2864
rect 2134 2859 2140 2860
rect 2238 2864 2244 2865
rect 2238 2860 2239 2864
rect 2243 2860 2244 2864
rect 2238 2859 2244 2860
rect 2114 2855 2120 2856
rect 2114 2851 2115 2855
rect 2119 2851 2120 2855
rect 2114 2850 2120 2851
rect 2306 2855 2312 2856
rect 2306 2851 2307 2855
rect 2311 2851 2312 2855
rect 2306 2850 2312 2851
rect 2116 2816 2118 2850
rect 2194 2847 2200 2848
rect 2194 2843 2195 2847
rect 2199 2843 2200 2847
rect 2194 2842 2200 2843
rect 2142 2826 2148 2827
rect 2142 2822 2143 2826
rect 2147 2822 2148 2826
rect 2142 2821 2148 2822
rect 2082 2815 2088 2816
rect 2082 2811 2083 2815
rect 2087 2811 2088 2815
rect 2082 2810 2088 2811
rect 2114 2815 2120 2816
rect 2114 2811 2115 2815
rect 2119 2811 2120 2815
rect 2114 2810 2120 2811
rect 2144 2799 2146 2821
rect 1871 2798 1875 2799
rect 1830 2796 1836 2797
rect 1830 2792 1831 2796
rect 1835 2792 1836 2796
rect 1871 2793 1875 2794
rect 1903 2798 1907 2799
rect 1903 2793 1907 2794
rect 2015 2798 2019 2799
rect 2022 2795 2023 2799
rect 2027 2795 2028 2799
rect 2022 2794 2028 2795
rect 2055 2798 2059 2799
rect 2015 2793 2019 2794
rect 1830 2791 1836 2792
rect 1230 2787 1236 2788
rect 1230 2783 1231 2787
rect 1235 2783 1236 2787
rect 1230 2782 1236 2783
rect 1286 2787 1292 2788
rect 1286 2783 1287 2787
rect 1291 2783 1292 2787
rect 1286 2782 1292 2783
rect 1458 2787 1464 2788
rect 1458 2783 1459 2787
rect 1463 2783 1464 2787
rect 1458 2782 1464 2783
rect 1578 2787 1584 2788
rect 1578 2783 1579 2787
rect 1583 2783 1584 2787
rect 1578 2782 1584 2783
rect 1714 2787 1720 2788
rect 1714 2783 1715 2787
rect 1719 2783 1720 2787
rect 1714 2782 1720 2783
rect 1830 2779 1836 2780
rect 1270 2776 1276 2777
rect 1270 2772 1271 2776
rect 1275 2772 1276 2776
rect 1270 2771 1276 2772
rect 1398 2776 1404 2777
rect 1398 2772 1399 2776
rect 1403 2772 1404 2776
rect 1398 2771 1404 2772
rect 1518 2776 1524 2777
rect 1518 2772 1519 2776
rect 1523 2772 1524 2776
rect 1518 2771 1524 2772
rect 1638 2776 1644 2777
rect 1638 2772 1639 2776
rect 1643 2772 1644 2776
rect 1638 2771 1644 2772
rect 1742 2776 1748 2777
rect 1742 2772 1743 2776
rect 1747 2772 1748 2776
rect 1830 2775 1831 2779
rect 1835 2775 1836 2779
rect 1830 2774 1836 2775
rect 1742 2771 1748 2772
rect 1272 2751 1274 2771
rect 1400 2751 1402 2771
rect 1520 2751 1522 2771
rect 1640 2751 1642 2771
rect 1730 2759 1736 2760
rect 1730 2755 1731 2759
rect 1735 2755 1736 2759
rect 1730 2754 1736 2755
rect 1271 2750 1275 2751
rect 1271 2745 1275 2746
rect 1287 2750 1291 2751
rect 1287 2745 1291 2746
rect 1399 2750 1403 2751
rect 1399 2745 1403 2746
rect 1447 2750 1451 2751
rect 1447 2745 1451 2746
rect 1519 2750 1523 2751
rect 1519 2745 1523 2746
rect 1607 2750 1611 2751
rect 1607 2745 1611 2746
rect 1639 2750 1643 2751
rect 1639 2745 1643 2746
rect 1288 2729 1290 2745
rect 1448 2729 1450 2745
rect 1608 2729 1610 2745
rect 1286 2728 1292 2729
rect 1286 2724 1287 2728
rect 1291 2724 1292 2728
rect 1286 2723 1292 2724
rect 1446 2728 1452 2729
rect 1446 2724 1447 2728
rect 1451 2724 1452 2728
rect 1446 2723 1452 2724
rect 1606 2728 1612 2729
rect 1606 2724 1607 2728
rect 1611 2724 1612 2728
rect 1606 2723 1612 2724
rect 578 2719 584 2720
rect 578 2715 579 2719
rect 583 2715 584 2719
rect 578 2714 584 2715
rect 730 2719 736 2720
rect 730 2715 731 2719
rect 735 2715 736 2719
rect 730 2714 736 2715
rect 1070 2719 1076 2720
rect 1070 2715 1071 2719
rect 1075 2715 1076 2719
rect 1070 2714 1076 2715
rect 1202 2719 1208 2720
rect 1202 2715 1203 2719
rect 1207 2715 1208 2719
rect 1202 2714 1208 2715
rect 1222 2719 1228 2720
rect 1222 2715 1223 2719
rect 1227 2715 1228 2719
rect 1222 2714 1228 2715
rect 1354 2719 1360 2720
rect 1354 2715 1355 2719
rect 1359 2715 1360 2719
rect 1354 2714 1360 2715
rect 570 2711 576 2712
rect 570 2707 571 2711
rect 575 2707 576 2711
rect 570 2706 576 2707
rect 518 2690 524 2691
rect 518 2686 519 2690
rect 523 2686 524 2690
rect 518 2685 524 2686
rect 394 2679 400 2680
rect 394 2675 395 2679
rect 399 2675 400 2679
rect 394 2674 400 2675
rect 520 2667 522 2685
rect 580 2680 582 2714
rect 670 2690 676 2691
rect 670 2686 671 2690
rect 675 2686 676 2690
rect 670 2685 676 2686
rect 578 2679 584 2680
rect 578 2675 579 2679
rect 583 2675 584 2679
rect 578 2674 584 2675
rect 672 2667 674 2685
rect 732 2680 734 2714
rect 822 2690 828 2691
rect 822 2686 823 2690
rect 827 2686 828 2690
rect 822 2685 828 2686
rect 982 2690 988 2691
rect 982 2686 983 2690
rect 987 2686 988 2690
rect 982 2685 988 2686
rect 730 2679 736 2680
rect 730 2675 731 2679
rect 735 2675 736 2679
rect 730 2674 736 2675
rect 824 2667 826 2685
rect 842 2679 848 2680
rect 842 2675 843 2679
rect 847 2675 848 2679
rect 842 2674 848 2675
rect 239 2666 243 2667
rect 239 2661 243 2662
rect 279 2666 283 2667
rect 279 2661 283 2662
rect 375 2666 379 2667
rect 375 2661 379 2662
rect 447 2666 451 2667
rect 447 2661 451 2662
rect 519 2666 523 2667
rect 519 2661 523 2662
rect 623 2666 627 2667
rect 623 2661 627 2662
rect 671 2666 675 2667
rect 671 2661 675 2662
rect 791 2666 795 2667
rect 791 2661 795 2662
rect 823 2666 827 2667
rect 823 2661 827 2662
rect 194 2659 200 2660
rect 194 2655 195 2659
rect 199 2655 200 2659
rect 194 2654 200 2655
rect 280 2651 282 2661
rect 330 2659 336 2660
rect 330 2655 331 2659
rect 335 2655 336 2659
rect 330 2654 336 2655
rect 142 2650 148 2651
rect 142 2646 143 2650
rect 147 2646 148 2650
rect 142 2645 148 2646
rect 278 2650 284 2651
rect 278 2646 279 2650
rect 283 2646 284 2650
rect 278 2645 284 2646
rect 110 2632 116 2633
rect 110 2628 111 2632
rect 115 2628 116 2632
rect 110 2627 116 2628
rect 332 2624 334 2654
rect 448 2651 450 2661
rect 586 2659 592 2660
rect 586 2655 587 2659
rect 591 2655 592 2659
rect 586 2654 592 2655
rect 446 2650 452 2651
rect 446 2646 447 2650
rect 451 2646 452 2650
rect 446 2645 452 2646
rect 330 2623 336 2624
rect 330 2619 331 2623
rect 335 2619 336 2623
rect 330 2618 336 2619
rect 110 2615 116 2616
rect 110 2611 111 2615
rect 115 2611 116 2615
rect 110 2610 116 2611
rect 134 2612 140 2613
rect 112 2587 114 2610
rect 134 2608 135 2612
rect 139 2608 140 2612
rect 134 2607 140 2608
rect 270 2612 276 2613
rect 270 2608 271 2612
rect 275 2608 276 2612
rect 270 2607 276 2608
rect 438 2612 444 2613
rect 438 2608 439 2612
rect 443 2608 444 2612
rect 438 2607 444 2608
rect 136 2587 138 2607
rect 272 2587 274 2607
rect 402 2595 408 2596
rect 402 2591 403 2595
rect 407 2591 408 2595
rect 402 2590 408 2591
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 135 2586 139 2587
rect 135 2581 139 2582
rect 223 2586 227 2587
rect 223 2581 227 2582
rect 271 2586 275 2587
rect 271 2581 275 2582
rect 367 2586 371 2587
rect 367 2581 371 2582
rect 112 2562 114 2581
rect 136 2565 138 2581
rect 224 2565 226 2581
rect 368 2565 370 2581
rect 134 2564 140 2565
rect 110 2561 116 2562
rect 110 2557 111 2561
rect 115 2557 116 2561
rect 134 2560 135 2564
rect 139 2560 140 2564
rect 134 2559 140 2560
rect 222 2564 228 2565
rect 222 2560 223 2564
rect 227 2560 228 2564
rect 222 2559 228 2560
rect 366 2564 372 2565
rect 366 2560 367 2564
rect 371 2560 372 2564
rect 366 2559 372 2560
rect 110 2556 116 2557
rect 202 2555 208 2556
rect 202 2551 203 2555
rect 207 2551 208 2555
rect 202 2550 208 2551
rect 290 2555 296 2556
rect 290 2551 291 2555
rect 295 2551 296 2555
rect 290 2550 296 2551
rect 194 2547 200 2548
rect 110 2544 116 2545
rect 110 2540 111 2544
rect 115 2540 116 2544
rect 194 2543 195 2547
rect 199 2543 200 2547
rect 194 2542 200 2543
rect 110 2539 116 2540
rect 112 2507 114 2539
rect 142 2526 148 2527
rect 142 2522 143 2526
rect 147 2522 148 2526
rect 142 2521 148 2522
rect 144 2507 146 2521
rect 111 2506 115 2507
rect 111 2501 115 2502
rect 143 2506 147 2507
rect 143 2501 147 2502
rect 112 2473 114 2501
rect 144 2491 146 2501
rect 196 2500 198 2542
rect 204 2516 206 2550
rect 230 2526 236 2527
rect 230 2522 231 2526
rect 235 2522 236 2526
rect 230 2521 236 2522
rect 202 2515 208 2516
rect 202 2511 203 2515
rect 207 2511 208 2515
rect 202 2510 208 2511
rect 232 2507 234 2521
rect 292 2516 294 2550
rect 374 2526 380 2527
rect 374 2522 375 2526
rect 379 2522 380 2526
rect 374 2521 380 2522
rect 290 2515 296 2516
rect 290 2511 291 2515
rect 295 2511 296 2515
rect 290 2510 296 2511
rect 376 2507 378 2521
rect 404 2516 406 2590
rect 440 2587 442 2607
rect 439 2586 443 2587
rect 439 2581 443 2582
rect 527 2586 531 2587
rect 527 2581 531 2582
rect 528 2565 530 2581
rect 526 2564 532 2565
rect 526 2560 527 2564
rect 531 2560 532 2564
rect 526 2559 532 2560
rect 588 2548 590 2654
rect 624 2651 626 2661
rect 792 2651 794 2661
rect 622 2650 628 2651
rect 622 2646 623 2650
rect 627 2646 628 2650
rect 622 2645 628 2646
rect 790 2650 796 2651
rect 790 2646 791 2650
rect 795 2646 796 2650
rect 790 2645 796 2646
rect 844 2624 846 2674
rect 984 2667 986 2685
rect 1007 2684 1011 2685
rect 1072 2680 1074 2714
rect 1142 2690 1148 2691
rect 1142 2686 1143 2690
rect 1147 2686 1148 2690
rect 1142 2685 1148 2686
rect 1224 2685 1226 2714
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1006 2679 1012 2680
rect 1006 2675 1007 2679
rect 1011 2675 1012 2679
rect 1006 2674 1012 2675
rect 1070 2679 1076 2680
rect 1070 2675 1071 2679
rect 1075 2675 1076 2679
rect 1070 2674 1076 2675
rect 1144 2667 1146 2685
rect 1223 2684 1227 2685
rect 1223 2679 1227 2680
rect 1296 2667 1298 2685
rect 1356 2680 1358 2714
rect 1454 2690 1460 2691
rect 1454 2686 1455 2690
rect 1459 2686 1460 2690
rect 1454 2685 1460 2686
rect 1614 2690 1620 2691
rect 1614 2686 1615 2690
rect 1619 2686 1620 2690
rect 1614 2685 1620 2686
rect 1354 2679 1360 2680
rect 1354 2675 1355 2679
rect 1359 2675 1360 2679
rect 1354 2674 1360 2675
rect 1456 2667 1458 2685
rect 1558 2679 1564 2680
rect 1558 2675 1559 2679
rect 1563 2675 1564 2679
rect 1558 2674 1564 2675
rect 951 2666 955 2667
rect 951 2661 955 2662
rect 983 2666 987 2667
rect 983 2661 987 2662
rect 1103 2666 1107 2667
rect 1103 2661 1107 2662
rect 1143 2666 1147 2667
rect 1143 2661 1147 2662
rect 1247 2666 1251 2667
rect 1247 2661 1251 2662
rect 1295 2666 1299 2667
rect 1295 2661 1299 2662
rect 1399 2666 1403 2667
rect 1399 2661 1403 2662
rect 1455 2666 1459 2667
rect 1455 2661 1459 2662
rect 1551 2666 1555 2667
rect 1551 2661 1555 2662
rect 952 2651 954 2661
rect 990 2659 996 2660
rect 990 2655 991 2659
rect 995 2655 996 2659
rect 990 2654 996 2655
rect 1002 2659 1008 2660
rect 1002 2655 1003 2659
rect 1007 2655 1008 2659
rect 1002 2654 1008 2655
rect 950 2650 956 2651
rect 950 2646 951 2650
rect 955 2646 956 2650
rect 950 2645 956 2646
rect 842 2623 848 2624
rect 842 2619 843 2623
rect 847 2619 848 2623
rect 842 2618 848 2619
rect 614 2612 620 2613
rect 614 2608 615 2612
rect 619 2608 620 2612
rect 614 2607 620 2608
rect 782 2612 788 2613
rect 782 2608 783 2612
rect 787 2608 788 2612
rect 782 2607 788 2608
rect 942 2612 948 2613
rect 942 2608 943 2612
rect 947 2608 948 2612
rect 942 2607 948 2608
rect 616 2587 618 2607
rect 784 2587 786 2607
rect 944 2587 946 2607
rect 615 2586 619 2587
rect 615 2581 619 2582
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 783 2586 787 2587
rect 783 2581 787 2582
rect 879 2586 883 2587
rect 879 2581 883 2582
rect 943 2586 947 2587
rect 943 2581 947 2582
rect 704 2565 706 2581
rect 880 2565 882 2581
rect 702 2564 708 2565
rect 702 2560 703 2564
rect 707 2560 708 2564
rect 702 2559 708 2560
rect 878 2564 884 2565
rect 878 2560 879 2564
rect 883 2560 884 2564
rect 878 2559 884 2560
rect 992 2556 994 2654
rect 1004 2624 1006 2654
rect 1104 2651 1106 2661
rect 1154 2659 1160 2660
rect 1154 2655 1155 2659
rect 1159 2655 1160 2659
rect 1154 2654 1160 2655
rect 1102 2650 1108 2651
rect 1102 2646 1103 2650
rect 1107 2646 1108 2650
rect 1102 2645 1108 2646
rect 1156 2624 1158 2654
rect 1248 2651 1250 2661
rect 1390 2659 1396 2660
rect 1390 2655 1391 2659
rect 1395 2655 1396 2659
rect 1390 2654 1396 2655
rect 1246 2650 1252 2651
rect 1246 2646 1247 2650
rect 1251 2646 1252 2650
rect 1246 2645 1252 2646
rect 1392 2624 1394 2654
rect 1400 2651 1402 2661
rect 1542 2659 1548 2660
rect 1542 2655 1543 2659
rect 1547 2655 1548 2659
rect 1542 2654 1548 2655
rect 1398 2650 1404 2651
rect 1398 2646 1399 2650
rect 1403 2646 1404 2650
rect 1398 2645 1404 2646
rect 1544 2624 1546 2654
rect 1552 2651 1554 2661
rect 1550 2650 1556 2651
rect 1550 2646 1551 2650
rect 1555 2646 1556 2650
rect 1550 2645 1556 2646
rect 1560 2624 1562 2674
rect 1616 2667 1618 2685
rect 1732 2680 1734 2754
rect 1744 2751 1746 2771
rect 1832 2751 1834 2774
rect 1872 2765 1874 2793
rect 1904 2783 1906 2793
rect 1954 2791 1960 2792
rect 1954 2787 1955 2791
rect 1959 2787 1960 2791
rect 1954 2786 1960 2787
rect 1902 2782 1908 2783
rect 1902 2778 1903 2782
rect 1907 2778 1908 2782
rect 1902 2777 1908 2778
rect 1870 2764 1876 2765
rect 1870 2760 1871 2764
rect 1875 2760 1876 2764
rect 1870 2759 1876 2760
rect 1956 2756 1958 2786
rect 2016 2783 2018 2793
rect 2014 2782 2020 2783
rect 2014 2778 2015 2782
rect 2019 2778 2020 2782
rect 2014 2777 2020 2778
rect 1954 2755 1960 2756
rect 1954 2751 1955 2755
rect 1959 2751 1960 2755
rect 1743 2750 1747 2751
rect 1743 2745 1747 2746
rect 1831 2750 1835 2751
rect 1954 2750 1960 2751
rect 1831 2745 1835 2746
rect 1870 2747 1876 2748
rect 1744 2729 1746 2745
rect 1742 2728 1748 2729
rect 1742 2724 1743 2728
rect 1747 2724 1748 2728
rect 1832 2726 1834 2745
rect 1870 2743 1871 2747
rect 1875 2743 1876 2747
rect 1870 2742 1876 2743
rect 1894 2744 1900 2745
rect 1742 2723 1748 2724
rect 1830 2725 1836 2726
rect 1830 2721 1831 2725
rect 1835 2721 1836 2725
rect 1872 2723 1874 2742
rect 1894 2740 1895 2744
rect 1899 2740 1900 2744
rect 1894 2739 1900 2740
rect 2006 2744 2012 2745
rect 2006 2740 2007 2744
rect 2011 2740 2012 2744
rect 2006 2739 2012 2740
rect 1896 2723 1898 2739
rect 2008 2723 2010 2739
rect 1830 2720 1836 2721
rect 1871 2722 1875 2723
rect 1842 2719 1848 2720
rect 1738 2715 1744 2716
rect 1738 2711 1739 2715
rect 1743 2711 1744 2715
rect 1842 2715 1843 2719
rect 1847 2715 1848 2719
rect 1871 2717 1875 2718
rect 1895 2722 1899 2723
rect 1895 2717 1899 2718
rect 2007 2722 2011 2723
rect 2007 2717 2011 2718
rect 1842 2714 1848 2715
rect 1738 2710 1744 2711
rect 1740 2680 1742 2710
rect 1830 2708 1836 2709
rect 1830 2704 1831 2708
rect 1835 2704 1836 2708
rect 1830 2703 1836 2704
rect 1750 2690 1756 2691
rect 1750 2686 1751 2690
rect 1755 2686 1756 2690
rect 1750 2685 1756 2686
rect 1730 2679 1736 2680
rect 1730 2675 1731 2679
rect 1735 2675 1736 2679
rect 1730 2674 1736 2675
rect 1738 2679 1744 2680
rect 1738 2675 1739 2679
rect 1743 2675 1744 2679
rect 1738 2674 1744 2675
rect 1752 2667 1754 2685
rect 1832 2667 1834 2703
rect 1615 2666 1619 2667
rect 1615 2661 1619 2662
rect 1751 2666 1755 2667
rect 1751 2661 1755 2662
rect 1831 2666 1835 2667
rect 1831 2661 1835 2662
rect 1832 2633 1834 2661
rect 1844 2652 1846 2714
rect 1872 2698 1874 2717
rect 1896 2701 1898 2717
rect 1894 2700 1900 2701
rect 1870 2697 1876 2698
rect 1870 2693 1871 2697
rect 1875 2693 1876 2697
rect 1894 2696 1895 2700
rect 1899 2696 1900 2700
rect 1894 2695 1900 2696
rect 1870 2692 1876 2693
rect 2024 2684 2026 2794
rect 2055 2793 2059 2794
rect 2143 2798 2147 2799
rect 2143 2793 2147 2794
rect 2167 2798 2171 2799
rect 2167 2793 2171 2794
rect 2168 2783 2170 2793
rect 2196 2792 2198 2842
rect 2246 2826 2252 2827
rect 2246 2822 2247 2826
rect 2251 2822 2252 2826
rect 2246 2821 2252 2822
rect 2248 2799 2250 2821
rect 2308 2816 2310 2850
rect 2316 2848 2318 2950
rect 2352 2920 2354 2950
rect 2368 2947 2370 2957
rect 2418 2955 2424 2956
rect 2418 2951 2419 2955
rect 2423 2951 2424 2955
rect 2418 2950 2424 2951
rect 2366 2946 2372 2947
rect 2366 2942 2367 2946
rect 2371 2942 2372 2946
rect 2366 2941 2372 2942
rect 2420 2920 2422 2950
rect 2448 2947 2450 2957
rect 2498 2955 2504 2956
rect 2498 2951 2499 2955
rect 2503 2951 2504 2955
rect 2498 2950 2504 2951
rect 2446 2946 2452 2947
rect 2446 2942 2447 2946
rect 2451 2942 2452 2946
rect 2446 2941 2452 2942
rect 2500 2920 2502 2950
rect 2528 2947 2530 2957
rect 2578 2955 2584 2956
rect 2578 2951 2579 2955
rect 2583 2951 2584 2955
rect 2578 2950 2584 2951
rect 2526 2946 2532 2947
rect 2526 2942 2527 2946
rect 2531 2942 2532 2946
rect 2526 2941 2532 2942
rect 2580 2920 2582 2950
rect 2608 2947 2610 2957
rect 2658 2955 2664 2956
rect 2658 2951 2659 2955
rect 2663 2951 2664 2955
rect 2658 2950 2664 2951
rect 2606 2946 2612 2947
rect 2606 2942 2607 2946
rect 2611 2942 2612 2946
rect 2606 2941 2612 2942
rect 2660 2920 2662 2950
rect 2696 2947 2698 2957
rect 2746 2955 2752 2956
rect 2746 2951 2747 2955
rect 2751 2951 2752 2955
rect 2746 2950 2752 2951
rect 2694 2946 2700 2947
rect 2694 2942 2695 2946
rect 2699 2942 2700 2946
rect 2694 2941 2700 2942
rect 2748 2920 2750 2950
rect 2792 2947 2794 2957
rect 2912 2947 2914 2957
rect 2946 2955 2952 2956
rect 2946 2951 2947 2955
rect 2951 2951 2952 2955
rect 2946 2950 2952 2951
rect 2962 2955 2968 2956
rect 2962 2951 2963 2955
rect 2967 2951 2968 2955
rect 2962 2950 2968 2951
rect 2790 2946 2796 2947
rect 2790 2942 2791 2946
rect 2795 2942 2796 2946
rect 2790 2941 2796 2942
rect 2910 2946 2916 2947
rect 2910 2942 2911 2946
rect 2915 2942 2916 2946
rect 2910 2941 2916 2942
rect 2350 2919 2356 2920
rect 2350 2915 2351 2919
rect 2355 2915 2356 2919
rect 2350 2914 2356 2915
rect 2418 2919 2424 2920
rect 2418 2915 2419 2919
rect 2423 2915 2424 2919
rect 2418 2914 2424 2915
rect 2498 2919 2504 2920
rect 2498 2915 2499 2919
rect 2503 2915 2504 2919
rect 2498 2914 2504 2915
rect 2578 2919 2584 2920
rect 2578 2915 2579 2919
rect 2583 2915 2584 2919
rect 2578 2914 2584 2915
rect 2658 2919 2664 2920
rect 2658 2915 2659 2919
rect 2663 2915 2664 2919
rect 2658 2914 2664 2915
rect 2746 2919 2752 2920
rect 2746 2915 2747 2919
rect 2751 2915 2752 2919
rect 2746 2914 2752 2915
rect 2358 2908 2364 2909
rect 2358 2904 2359 2908
rect 2363 2904 2364 2908
rect 2358 2903 2364 2904
rect 2438 2908 2444 2909
rect 2438 2904 2439 2908
rect 2443 2904 2444 2908
rect 2438 2903 2444 2904
rect 2518 2908 2524 2909
rect 2518 2904 2519 2908
rect 2523 2904 2524 2908
rect 2518 2903 2524 2904
rect 2598 2908 2604 2909
rect 2598 2904 2599 2908
rect 2603 2904 2604 2908
rect 2598 2903 2604 2904
rect 2686 2908 2692 2909
rect 2686 2904 2687 2908
rect 2691 2904 2692 2908
rect 2686 2903 2692 2904
rect 2782 2908 2788 2909
rect 2782 2904 2783 2908
rect 2787 2904 2788 2908
rect 2782 2903 2788 2904
rect 2902 2908 2908 2909
rect 2902 2904 2903 2908
rect 2907 2904 2908 2908
rect 2902 2903 2908 2904
rect 2360 2887 2362 2903
rect 2440 2887 2442 2903
rect 2520 2887 2522 2903
rect 2600 2887 2602 2903
rect 2626 2891 2632 2892
rect 2626 2887 2627 2891
rect 2631 2887 2632 2891
rect 2688 2887 2690 2903
rect 2784 2887 2786 2903
rect 2904 2887 2906 2903
rect 2343 2886 2347 2887
rect 2343 2881 2347 2882
rect 2359 2886 2363 2887
rect 2359 2881 2363 2882
rect 2439 2886 2443 2887
rect 2439 2881 2443 2882
rect 2463 2886 2467 2887
rect 2463 2881 2467 2882
rect 2519 2886 2523 2887
rect 2519 2881 2523 2882
rect 2591 2886 2595 2887
rect 2591 2881 2595 2882
rect 2599 2886 2603 2887
rect 2626 2886 2632 2887
rect 2687 2886 2691 2887
rect 2599 2881 2603 2882
rect 2344 2865 2346 2881
rect 2464 2865 2466 2881
rect 2592 2865 2594 2881
rect 2342 2864 2348 2865
rect 2342 2860 2343 2864
rect 2347 2860 2348 2864
rect 2342 2859 2348 2860
rect 2462 2864 2468 2865
rect 2462 2860 2463 2864
rect 2467 2860 2468 2864
rect 2462 2859 2468 2860
rect 2590 2864 2596 2865
rect 2590 2860 2591 2864
rect 2595 2860 2596 2864
rect 2590 2859 2596 2860
rect 2410 2855 2416 2856
rect 2410 2851 2411 2855
rect 2415 2851 2416 2855
rect 2410 2850 2416 2851
rect 2314 2847 2320 2848
rect 2314 2843 2315 2847
rect 2319 2843 2320 2847
rect 2314 2842 2320 2843
rect 2350 2826 2356 2827
rect 2350 2822 2351 2826
rect 2355 2822 2356 2826
rect 2350 2821 2356 2822
rect 2306 2815 2312 2816
rect 2306 2811 2307 2815
rect 2311 2811 2312 2815
rect 2306 2810 2312 2811
rect 2352 2799 2354 2821
rect 2412 2816 2414 2850
rect 2470 2826 2476 2827
rect 2470 2822 2471 2826
rect 2475 2822 2476 2826
rect 2470 2821 2476 2822
rect 2598 2826 2604 2827
rect 2598 2822 2599 2826
rect 2603 2822 2604 2826
rect 2598 2821 2604 2822
rect 2410 2815 2416 2816
rect 2410 2811 2411 2815
rect 2415 2811 2416 2815
rect 2410 2810 2416 2811
rect 2472 2799 2474 2821
rect 2494 2815 2500 2816
rect 2494 2811 2495 2815
rect 2499 2811 2500 2815
rect 2494 2810 2500 2811
rect 2247 2798 2251 2799
rect 2247 2793 2251 2794
rect 2327 2798 2331 2799
rect 2327 2793 2331 2794
rect 2351 2798 2355 2799
rect 2351 2793 2355 2794
rect 2471 2798 2475 2799
rect 2471 2793 2475 2794
rect 2487 2798 2491 2799
rect 2487 2793 2491 2794
rect 2194 2791 2200 2792
rect 2194 2787 2195 2791
rect 2199 2787 2200 2791
rect 2194 2786 2200 2787
rect 2218 2791 2224 2792
rect 2218 2787 2219 2791
rect 2223 2787 2224 2791
rect 2218 2786 2224 2787
rect 2166 2782 2172 2783
rect 2067 2780 2071 2781
rect 2166 2778 2167 2782
rect 2171 2778 2172 2782
rect 2166 2777 2172 2778
rect 2067 2775 2071 2776
rect 2068 2756 2070 2775
rect 2220 2756 2222 2786
rect 2328 2783 2330 2793
rect 2418 2791 2424 2792
rect 2418 2787 2419 2791
rect 2423 2787 2424 2791
rect 2418 2786 2424 2787
rect 2326 2782 2332 2783
rect 2326 2778 2327 2782
rect 2331 2778 2332 2782
rect 2420 2781 2422 2786
rect 2488 2783 2490 2793
rect 2486 2782 2492 2783
rect 2326 2777 2332 2778
rect 2419 2780 2423 2781
rect 2486 2778 2487 2782
rect 2491 2778 2492 2782
rect 2486 2777 2492 2778
rect 2419 2775 2423 2776
rect 2496 2756 2498 2810
rect 2600 2799 2602 2821
rect 2628 2816 2630 2886
rect 2687 2881 2691 2882
rect 2727 2886 2731 2887
rect 2727 2881 2731 2882
rect 2783 2886 2787 2887
rect 2783 2881 2787 2882
rect 2879 2886 2883 2887
rect 2879 2881 2883 2882
rect 2903 2886 2907 2887
rect 2903 2881 2907 2882
rect 2728 2865 2730 2881
rect 2880 2865 2882 2881
rect 2726 2864 2732 2865
rect 2726 2860 2727 2864
rect 2731 2860 2732 2864
rect 2726 2859 2732 2860
rect 2878 2864 2884 2865
rect 2878 2860 2879 2864
rect 2883 2860 2884 2864
rect 2878 2859 2884 2860
rect 2948 2856 2950 2950
rect 2964 2920 2966 2950
rect 3040 2947 3042 2957
rect 3100 2956 3102 3006
rect 3108 2980 3110 3014
rect 3190 2990 3196 2991
rect 3190 2986 3191 2990
rect 3195 2986 3196 2990
rect 3190 2985 3196 2986
rect 3106 2979 3112 2980
rect 3106 2975 3107 2979
rect 3111 2975 3112 2979
rect 3106 2974 3112 2975
rect 3192 2963 3194 2985
rect 3252 2980 3254 3014
rect 3284 2980 3286 3090
rect 3590 3087 3596 3088
rect 3382 3084 3388 3085
rect 3382 3080 3383 3084
rect 3387 3080 3388 3084
rect 3590 3083 3591 3087
rect 3595 3083 3596 3087
rect 3590 3082 3596 3083
rect 3382 3079 3388 3080
rect 3384 3051 3386 3079
rect 3592 3051 3594 3082
rect 3327 3050 3331 3051
rect 3327 3045 3331 3046
rect 3383 3050 3387 3051
rect 3383 3045 3387 3046
rect 3591 3050 3595 3051
rect 3591 3045 3595 3046
rect 3328 3029 3330 3045
rect 3326 3028 3332 3029
rect 3326 3024 3327 3028
rect 3331 3024 3332 3028
rect 3592 3026 3594 3045
rect 3326 3023 3332 3024
rect 3590 3025 3596 3026
rect 3590 3021 3591 3025
rect 3595 3021 3596 3025
rect 3590 3020 3596 3021
rect 3590 3008 3596 3009
rect 3590 3004 3591 3008
rect 3595 3004 3596 3008
rect 3590 3003 3596 3004
rect 3334 2990 3340 2991
rect 3334 2986 3335 2990
rect 3339 2986 3340 2990
rect 3334 2985 3340 2986
rect 3250 2979 3256 2980
rect 3250 2975 3251 2979
rect 3255 2975 3256 2979
rect 3250 2974 3256 2975
rect 3282 2979 3288 2980
rect 3282 2975 3283 2979
rect 3287 2975 3288 2979
rect 3282 2974 3288 2975
rect 3336 2963 3338 2985
rect 3592 2963 3594 3003
rect 3183 2962 3187 2963
rect 3183 2957 3187 2958
rect 3191 2962 3195 2963
rect 3191 2957 3195 2958
rect 3335 2962 3339 2963
rect 3335 2957 3339 2958
rect 3495 2962 3499 2963
rect 3495 2957 3499 2958
rect 3591 2962 3595 2963
rect 3591 2957 3595 2958
rect 3098 2955 3104 2956
rect 3098 2951 3099 2955
rect 3103 2951 3104 2955
rect 3098 2950 3104 2951
rect 3184 2947 3186 2957
rect 3234 2955 3240 2956
rect 3234 2951 3235 2955
rect 3239 2951 3240 2955
rect 3234 2950 3240 2951
rect 3038 2946 3044 2947
rect 3038 2942 3039 2946
rect 3043 2942 3044 2946
rect 3038 2941 3044 2942
rect 3182 2946 3188 2947
rect 3182 2942 3183 2946
rect 3187 2942 3188 2946
rect 3182 2941 3188 2942
rect 3236 2920 3238 2950
rect 3336 2947 3338 2957
rect 3438 2955 3444 2956
rect 3438 2951 3439 2955
rect 3443 2951 3444 2955
rect 3438 2950 3444 2951
rect 3334 2946 3340 2947
rect 3334 2942 3335 2946
rect 3339 2942 3340 2946
rect 3334 2941 3340 2942
rect 2962 2919 2968 2920
rect 2962 2915 2963 2919
rect 2967 2915 2968 2919
rect 2962 2914 2968 2915
rect 3234 2919 3240 2920
rect 3234 2915 3235 2919
rect 3239 2915 3240 2919
rect 3234 2914 3240 2915
rect 3030 2908 3036 2909
rect 3030 2904 3031 2908
rect 3035 2904 3036 2908
rect 3030 2903 3036 2904
rect 3174 2908 3180 2909
rect 3174 2904 3175 2908
rect 3179 2904 3180 2908
rect 3174 2903 3180 2904
rect 3326 2908 3332 2909
rect 3326 2904 3327 2908
rect 3331 2904 3332 2908
rect 3326 2903 3332 2904
rect 3032 2887 3034 2903
rect 3176 2887 3178 2903
rect 3226 2891 3232 2892
rect 3226 2887 3227 2891
rect 3231 2887 3232 2891
rect 3328 2887 3330 2903
rect 3031 2886 3035 2887
rect 3031 2881 3035 2882
rect 3175 2886 3179 2887
rect 3175 2881 3179 2882
rect 3191 2886 3195 2887
rect 3226 2886 3232 2887
rect 3327 2886 3331 2887
rect 3191 2881 3195 2882
rect 3032 2865 3034 2881
rect 3192 2865 3194 2881
rect 3030 2864 3036 2865
rect 3030 2860 3031 2864
rect 3035 2860 3036 2864
rect 3030 2859 3036 2860
rect 3190 2864 3196 2865
rect 3190 2860 3191 2864
rect 3195 2860 3196 2864
rect 3190 2859 3196 2860
rect 2682 2855 2688 2856
rect 2682 2851 2683 2855
rect 2687 2851 2688 2855
rect 2682 2850 2688 2851
rect 2794 2855 2800 2856
rect 2794 2851 2795 2855
rect 2799 2851 2800 2855
rect 2794 2850 2800 2851
rect 2946 2855 2952 2856
rect 2946 2851 2947 2855
rect 2951 2851 2952 2855
rect 2946 2850 2952 2851
rect 2958 2855 2964 2856
rect 2958 2851 2959 2855
rect 2963 2851 2964 2855
rect 2958 2850 2964 2851
rect 3098 2855 3104 2856
rect 3098 2851 3099 2855
rect 3103 2851 3104 2855
rect 3098 2850 3104 2851
rect 2667 2820 2671 2821
rect 2684 2816 2686 2850
rect 2734 2826 2740 2827
rect 2734 2822 2735 2826
rect 2739 2822 2740 2826
rect 2734 2821 2740 2822
rect 2626 2815 2632 2816
rect 2667 2815 2671 2816
rect 2682 2815 2688 2816
rect 2626 2811 2627 2815
rect 2631 2811 2632 2815
rect 2626 2810 2632 2811
rect 2599 2798 2603 2799
rect 2599 2793 2603 2794
rect 2639 2798 2643 2799
rect 2639 2793 2643 2794
rect 2640 2783 2642 2793
rect 2668 2792 2670 2815
rect 2682 2811 2683 2815
rect 2687 2811 2688 2815
rect 2682 2810 2688 2811
rect 2736 2799 2738 2821
rect 2796 2816 2798 2850
rect 2886 2826 2892 2827
rect 2886 2822 2887 2826
rect 2891 2822 2892 2826
rect 2886 2821 2892 2822
rect 2960 2821 2962 2850
rect 3038 2826 3044 2827
rect 3038 2822 3039 2826
rect 3043 2822 3044 2826
rect 3038 2821 3044 2822
rect 2794 2815 2800 2816
rect 2794 2811 2795 2815
rect 2799 2811 2800 2815
rect 2794 2810 2800 2811
rect 2888 2799 2890 2821
rect 2959 2820 2963 2821
rect 2959 2815 2963 2816
rect 3040 2799 3042 2821
rect 3100 2816 3102 2850
rect 3198 2826 3204 2827
rect 3198 2822 3199 2826
rect 3203 2822 3204 2826
rect 3198 2821 3204 2822
rect 3098 2815 3104 2816
rect 3098 2811 3099 2815
rect 3103 2811 3104 2815
rect 3098 2810 3104 2811
rect 3200 2799 3202 2821
rect 3228 2816 3230 2886
rect 3327 2881 3331 2882
rect 3359 2886 3363 2887
rect 3359 2881 3363 2882
rect 3360 2865 3362 2881
rect 3358 2864 3364 2865
rect 3358 2860 3359 2864
rect 3363 2860 3364 2864
rect 3358 2859 3364 2860
rect 3440 2856 3442 2950
rect 3496 2947 3498 2957
rect 3494 2946 3500 2947
rect 3494 2942 3495 2946
rect 3499 2942 3500 2946
rect 3494 2941 3500 2942
rect 3592 2929 3594 2957
rect 3590 2928 3596 2929
rect 3590 2924 3591 2928
rect 3595 2924 3596 2928
rect 3590 2923 3596 2924
rect 3534 2919 3540 2920
rect 3534 2915 3535 2919
rect 3539 2915 3540 2919
rect 3534 2914 3540 2915
rect 3486 2908 3492 2909
rect 3486 2904 3487 2908
rect 3491 2904 3492 2908
rect 3486 2903 3492 2904
rect 3488 2887 3490 2903
rect 3487 2886 3491 2887
rect 3487 2881 3491 2882
rect 3503 2886 3507 2887
rect 3503 2881 3507 2882
rect 3504 2865 3506 2881
rect 3502 2864 3508 2865
rect 3502 2860 3503 2864
rect 3507 2860 3508 2864
rect 3502 2859 3508 2860
rect 3438 2855 3444 2856
rect 3438 2851 3439 2855
rect 3443 2851 3444 2855
rect 3438 2850 3444 2851
rect 3366 2826 3372 2827
rect 3366 2822 3367 2826
rect 3371 2822 3372 2826
rect 3366 2821 3372 2822
rect 3510 2826 3516 2827
rect 3510 2822 3511 2826
rect 3515 2822 3516 2826
rect 3510 2821 3516 2822
rect 3226 2815 3232 2816
rect 3226 2811 3227 2815
rect 3231 2811 3232 2815
rect 3226 2810 3232 2811
rect 3368 2799 3370 2821
rect 3390 2815 3396 2816
rect 3390 2811 3391 2815
rect 3395 2811 3396 2815
rect 3390 2810 3396 2811
rect 2735 2798 2739 2799
rect 2735 2793 2739 2794
rect 2791 2798 2795 2799
rect 2791 2793 2795 2794
rect 2887 2798 2891 2799
rect 2887 2793 2891 2794
rect 2943 2798 2947 2799
rect 2943 2793 2947 2794
rect 3039 2798 3043 2799
rect 3039 2793 3043 2794
rect 3087 2798 3091 2799
rect 3087 2793 3091 2794
rect 3199 2798 3203 2799
rect 3199 2793 3203 2794
rect 3231 2798 3235 2799
rect 3231 2793 3235 2794
rect 3367 2798 3371 2799
rect 3367 2793 3371 2794
rect 3383 2798 3387 2799
rect 3383 2793 3387 2794
rect 2666 2791 2672 2792
rect 2666 2787 2667 2791
rect 2671 2787 2672 2791
rect 2666 2786 2672 2787
rect 2690 2791 2696 2792
rect 2690 2787 2691 2791
rect 2695 2787 2696 2791
rect 2690 2786 2696 2787
rect 2638 2782 2644 2783
rect 2638 2778 2639 2782
rect 2643 2778 2644 2782
rect 2638 2777 2644 2778
rect 2692 2756 2694 2786
rect 2792 2783 2794 2793
rect 2842 2791 2848 2792
rect 2842 2787 2843 2791
rect 2847 2787 2848 2791
rect 2842 2786 2848 2787
rect 2790 2782 2796 2783
rect 2790 2778 2791 2782
rect 2795 2778 2796 2782
rect 2790 2777 2796 2778
rect 2844 2756 2846 2786
rect 2944 2783 2946 2793
rect 2994 2791 3000 2792
rect 2994 2787 2995 2791
rect 2999 2787 3000 2791
rect 2994 2786 3000 2787
rect 2942 2782 2948 2783
rect 2942 2778 2943 2782
rect 2947 2778 2948 2782
rect 2942 2777 2948 2778
rect 2996 2756 2998 2786
rect 3088 2783 3090 2793
rect 3138 2791 3144 2792
rect 3138 2787 3139 2791
rect 3143 2787 3144 2791
rect 3138 2786 3144 2787
rect 3086 2782 3092 2783
rect 3086 2778 3087 2782
rect 3091 2778 3092 2782
rect 3086 2777 3092 2778
rect 3140 2756 3142 2786
rect 3232 2783 3234 2793
rect 3384 2783 3386 2793
rect 3230 2782 3236 2783
rect 3230 2778 3231 2782
rect 3235 2778 3236 2782
rect 3230 2777 3236 2778
rect 3382 2782 3388 2783
rect 3382 2778 3383 2782
rect 3387 2778 3388 2782
rect 3382 2777 3388 2778
rect 3392 2756 3394 2810
rect 3512 2799 3514 2821
rect 3536 2816 3538 2914
rect 3590 2911 3596 2912
rect 3590 2907 3591 2911
rect 3595 2907 3596 2911
rect 3590 2906 3596 2907
rect 3592 2887 3594 2906
rect 3591 2886 3595 2887
rect 3591 2881 3595 2882
rect 3592 2862 3594 2881
rect 3590 2861 3596 2862
rect 3590 2857 3591 2861
rect 3595 2857 3596 2861
rect 3590 2856 3596 2857
rect 3562 2847 3568 2848
rect 3562 2843 3563 2847
rect 3567 2843 3568 2847
rect 3562 2842 3568 2843
rect 3590 2844 3596 2845
rect 3534 2815 3540 2816
rect 3534 2811 3535 2815
rect 3539 2811 3540 2815
rect 3534 2810 3540 2811
rect 3511 2798 3515 2799
rect 3511 2793 3515 2794
rect 3442 2791 3448 2792
rect 3442 2787 3443 2791
rect 3447 2787 3448 2791
rect 3442 2786 3448 2787
rect 2066 2755 2072 2756
rect 2066 2751 2067 2755
rect 2071 2751 2072 2755
rect 2066 2750 2072 2751
rect 2218 2755 2224 2756
rect 2218 2751 2219 2755
rect 2223 2751 2224 2755
rect 2218 2750 2224 2751
rect 2358 2755 2364 2756
rect 2358 2751 2359 2755
rect 2363 2751 2364 2755
rect 2358 2750 2364 2751
rect 2494 2755 2500 2756
rect 2494 2751 2495 2755
rect 2499 2751 2500 2755
rect 2494 2750 2500 2751
rect 2690 2755 2696 2756
rect 2690 2751 2691 2755
rect 2695 2751 2696 2755
rect 2690 2750 2696 2751
rect 2842 2755 2848 2756
rect 2842 2751 2843 2755
rect 2847 2751 2848 2755
rect 2842 2750 2848 2751
rect 2994 2755 3000 2756
rect 2994 2751 2995 2755
rect 2999 2751 3000 2755
rect 2994 2750 3000 2751
rect 3138 2755 3144 2756
rect 3138 2751 3139 2755
rect 3143 2751 3144 2755
rect 3138 2750 3144 2751
rect 3390 2755 3396 2756
rect 3390 2751 3391 2755
rect 3395 2751 3396 2755
rect 3390 2750 3396 2751
rect 2158 2744 2164 2745
rect 2158 2740 2159 2744
rect 2163 2740 2164 2744
rect 2158 2739 2164 2740
rect 2318 2744 2324 2745
rect 2318 2740 2319 2744
rect 2323 2740 2324 2744
rect 2318 2739 2324 2740
rect 2160 2723 2162 2739
rect 2320 2723 2322 2739
rect 2103 2722 2107 2723
rect 2103 2717 2107 2718
rect 2159 2722 2163 2723
rect 2159 2717 2163 2718
rect 2319 2722 2323 2723
rect 2319 2717 2323 2718
rect 2327 2722 2331 2723
rect 2327 2717 2331 2718
rect 2104 2701 2106 2717
rect 2328 2701 2330 2717
rect 2102 2700 2108 2701
rect 2102 2696 2103 2700
rect 2107 2696 2108 2700
rect 2102 2695 2108 2696
rect 2326 2700 2332 2701
rect 2326 2696 2327 2700
rect 2331 2696 2332 2700
rect 2326 2695 2332 2696
rect 2022 2683 2028 2684
rect 1870 2680 1876 2681
rect 1870 2676 1871 2680
rect 1875 2676 1876 2680
rect 2022 2679 2023 2683
rect 2027 2679 2028 2683
rect 2022 2678 2028 2679
rect 1870 2675 1876 2676
rect 1842 2651 1848 2652
rect 1842 2647 1843 2651
rect 1847 2647 1848 2651
rect 1842 2646 1848 2647
rect 1872 2639 1874 2675
rect 1902 2662 1908 2663
rect 1902 2658 1903 2662
rect 1907 2658 1908 2662
rect 2110 2662 2116 2663
rect 1902 2657 1908 2658
rect 1931 2660 1935 2661
rect 1904 2639 1906 2657
rect 2110 2658 2111 2662
rect 2115 2658 2116 2662
rect 2110 2657 2116 2658
rect 2334 2662 2340 2663
rect 2334 2658 2335 2662
rect 2339 2658 2340 2662
rect 2334 2657 2340 2658
rect 1931 2655 1935 2656
rect 1871 2638 1875 2639
rect 1871 2633 1875 2634
rect 1903 2638 1907 2639
rect 1903 2633 1907 2634
rect 1830 2632 1836 2633
rect 1830 2628 1831 2632
rect 1835 2628 1836 2632
rect 1830 2627 1836 2628
rect 1002 2623 1008 2624
rect 1002 2619 1003 2623
rect 1007 2619 1008 2623
rect 1002 2618 1008 2619
rect 1154 2623 1160 2624
rect 1154 2619 1155 2623
rect 1159 2619 1160 2623
rect 1154 2618 1160 2619
rect 1390 2623 1396 2624
rect 1390 2619 1391 2623
rect 1395 2619 1396 2623
rect 1390 2618 1396 2619
rect 1542 2623 1548 2624
rect 1542 2619 1543 2623
rect 1547 2619 1548 2623
rect 1542 2618 1548 2619
rect 1558 2623 1564 2624
rect 1558 2619 1559 2623
rect 1563 2619 1564 2623
rect 1558 2618 1564 2619
rect 1830 2615 1836 2616
rect 1094 2612 1100 2613
rect 1094 2608 1095 2612
rect 1099 2608 1100 2612
rect 1094 2607 1100 2608
rect 1238 2612 1244 2613
rect 1238 2608 1239 2612
rect 1243 2608 1244 2612
rect 1238 2607 1244 2608
rect 1390 2612 1396 2613
rect 1390 2608 1391 2612
rect 1395 2608 1396 2612
rect 1390 2607 1396 2608
rect 1542 2612 1548 2613
rect 1542 2608 1543 2612
rect 1547 2608 1548 2612
rect 1830 2611 1831 2615
rect 1835 2611 1836 2615
rect 1830 2610 1836 2611
rect 1542 2607 1548 2608
rect 1096 2587 1098 2607
rect 1240 2587 1242 2607
rect 1392 2587 1394 2607
rect 1544 2587 1546 2607
rect 1832 2587 1834 2610
rect 1872 2605 1874 2633
rect 1904 2623 1906 2633
rect 1932 2632 1934 2655
rect 2112 2639 2114 2657
rect 2336 2639 2338 2657
rect 2360 2652 2362 2750
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2630 2744 2636 2745
rect 2630 2740 2631 2744
rect 2635 2740 2636 2744
rect 2630 2739 2636 2740
rect 2782 2744 2788 2745
rect 2782 2740 2783 2744
rect 2787 2740 2788 2744
rect 2782 2739 2788 2740
rect 2934 2744 2940 2745
rect 2934 2740 2935 2744
rect 2939 2740 2940 2744
rect 2934 2739 2940 2740
rect 3078 2744 3084 2745
rect 3078 2740 3079 2744
rect 3083 2740 3084 2744
rect 3078 2739 3084 2740
rect 3222 2744 3228 2745
rect 3222 2740 3223 2744
rect 3227 2740 3228 2744
rect 3222 2739 3228 2740
rect 3374 2744 3380 2745
rect 3374 2740 3375 2744
rect 3379 2740 3380 2744
rect 3374 2739 3380 2740
rect 2480 2723 2482 2739
rect 2632 2723 2634 2739
rect 2784 2723 2786 2739
rect 2936 2723 2938 2739
rect 3080 2723 3082 2739
rect 3138 2727 3144 2728
rect 3138 2723 3139 2727
rect 3143 2723 3144 2727
rect 3224 2723 3226 2739
rect 3376 2723 3378 2739
rect 2479 2722 2483 2723
rect 2479 2717 2483 2718
rect 2535 2722 2539 2723
rect 2535 2717 2539 2718
rect 2631 2722 2635 2723
rect 2631 2717 2635 2718
rect 2735 2722 2739 2723
rect 2735 2717 2739 2718
rect 2783 2722 2787 2723
rect 2783 2717 2787 2718
rect 2911 2722 2915 2723
rect 2911 2717 2915 2718
rect 2935 2722 2939 2723
rect 2935 2717 2939 2718
rect 3071 2722 3075 2723
rect 3071 2717 3075 2718
rect 3079 2722 3083 2723
rect 3138 2722 3144 2723
rect 3223 2722 3227 2723
rect 3079 2717 3083 2718
rect 2536 2701 2538 2717
rect 2736 2701 2738 2717
rect 2912 2701 2914 2717
rect 3072 2701 3074 2717
rect 2534 2700 2540 2701
rect 2534 2696 2535 2700
rect 2539 2696 2540 2700
rect 2534 2695 2540 2696
rect 2734 2700 2740 2701
rect 2734 2696 2735 2700
rect 2739 2696 2740 2700
rect 2734 2695 2740 2696
rect 2910 2700 2916 2701
rect 2910 2696 2911 2700
rect 2915 2696 2916 2700
rect 2910 2695 2916 2696
rect 3070 2700 3076 2701
rect 3070 2696 3071 2700
rect 3075 2696 3076 2700
rect 3070 2695 3076 2696
rect 2454 2691 2460 2692
rect 2454 2687 2455 2691
rect 2459 2687 2460 2691
rect 2454 2686 2460 2687
rect 2478 2691 2484 2692
rect 2478 2687 2479 2691
rect 2483 2687 2484 2691
rect 2478 2686 2484 2687
rect 3014 2691 3020 2692
rect 3014 2687 3015 2691
rect 3019 2687 3020 2691
rect 3014 2686 3020 2687
rect 2456 2652 2458 2686
rect 2480 2661 2482 2686
rect 2542 2662 2548 2663
rect 2479 2660 2483 2661
rect 2542 2658 2543 2662
rect 2547 2658 2548 2662
rect 2542 2657 2548 2658
rect 2742 2662 2748 2663
rect 2742 2658 2743 2662
rect 2747 2658 2748 2662
rect 2918 2662 2924 2663
rect 2742 2657 2748 2658
rect 2771 2660 2775 2661
rect 2479 2655 2483 2656
rect 2358 2651 2364 2652
rect 2358 2647 2359 2651
rect 2363 2647 2364 2651
rect 2358 2646 2364 2647
rect 2454 2651 2460 2652
rect 2454 2647 2455 2651
rect 2459 2647 2460 2651
rect 2454 2646 2460 2647
rect 2544 2639 2546 2657
rect 2744 2639 2746 2657
rect 2918 2658 2919 2662
rect 2923 2658 2924 2662
rect 2918 2657 2924 2658
rect 2771 2655 2775 2656
rect 2772 2652 2774 2655
rect 2770 2651 2776 2652
rect 2770 2647 2771 2651
rect 2775 2647 2776 2651
rect 2770 2646 2776 2647
rect 2920 2639 2922 2657
rect 3016 2652 3018 2686
rect 3078 2662 3084 2663
rect 3078 2658 3079 2662
rect 3083 2658 3084 2662
rect 3140 2661 3142 2722
rect 3223 2717 3227 2718
rect 3375 2722 3379 2723
rect 3375 2717 3379 2718
rect 3224 2701 3226 2717
rect 3376 2701 3378 2717
rect 3222 2700 3228 2701
rect 3222 2696 3223 2700
rect 3227 2696 3228 2700
rect 3222 2695 3228 2696
rect 3374 2700 3380 2701
rect 3374 2696 3375 2700
rect 3379 2696 3380 2700
rect 3374 2695 3380 2696
rect 3444 2692 3446 2786
rect 3512 2783 3514 2793
rect 3564 2792 3566 2842
rect 3590 2840 3591 2844
rect 3595 2840 3596 2844
rect 3590 2839 3596 2840
rect 3592 2799 3594 2839
rect 3591 2798 3595 2799
rect 3591 2793 3595 2794
rect 3562 2791 3568 2792
rect 3562 2787 3563 2791
rect 3567 2787 3568 2791
rect 3562 2786 3568 2787
rect 3510 2782 3516 2783
rect 3510 2778 3511 2782
rect 3515 2778 3516 2782
rect 3510 2777 3516 2778
rect 3592 2765 3594 2793
rect 3590 2764 3596 2765
rect 3590 2760 3591 2764
rect 3595 2760 3596 2764
rect 3590 2759 3596 2760
rect 3534 2755 3540 2756
rect 3534 2751 3535 2755
rect 3539 2751 3540 2755
rect 3534 2750 3540 2751
rect 3502 2744 3508 2745
rect 3502 2740 3503 2744
rect 3507 2740 3508 2744
rect 3502 2739 3508 2740
rect 3504 2723 3506 2739
rect 3503 2722 3507 2723
rect 3503 2717 3507 2718
rect 3504 2701 3506 2717
rect 3502 2700 3508 2701
rect 3502 2696 3503 2700
rect 3507 2696 3508 2700
rect 3502 2695 3508 2696
rect 3170 2691 3176 2692
rect 3170 2687 3171 2691
rect 3175 2687 3176 2691
rect 3170 2686 3176 2687
rect 3322 2691 3328 2692
rect 3322 2687 3323 2691
rect 3327 2687 3328 2691
rect 3322 2686 3328 2687
rect 3442 2691 3448 2692
rect 3442 2687 3443 2691
rect 3447 2687 3448 2691
rect 3442 2686 3448 2687
rect 3078 2657 3084 2658
rect 3139 2660 3143 2661
rect 3014 2651 3020 2652
rect 3014 2647 3015 2651
rect 3019 2647 3020 2651
rect 3014 2646 3020 2647
rect 3080 2639 3082 2657
rect 3139 2655 3143 2656
rect 3172 2652 3174 2686
rect 3230 2662 3236 2663
rect 3230 2658 3231 2662
rect 3235 2658 3236 2662
rect 3230 2657 3236 2658
rect 3170 2651 3176 2652
rect 3170 2647 3171 2651
rect 3175 2647 3176 2651
rect 3170 2646 3176 2647
rect 3232 2639 3234 2657
rect 3324 2652 3326 2686
rect 3382 2662 3388 2663
rect 3382 2658 3383 2662
rect 3387 2658 3388 2662
rect 3382 2657 3388 2658
rect 3510 2662 3516 2663
rect 3510 2658 3511 2662
rect 3515 2658 3516 2662
rect 3510 2657 3516 2658
rect 3322 2651 3328 2652
rect 3322 2647 3323 2651
rect 3327 2647 3328 2651
rect 3322 2646 3328 2647
rect 3384 2639 3386 2657
rect 3512 2639 3514 2657
rect 3536 2652 3538 2750
rect 3590 2747 3596 2748
rect 3590 2743 3591 2747
rect 3595 2743 3596 2747
rect 3590 2742 3596 2743
rect 3592 2723 3594 2742
rect 3591 2722 3595 2723
rect 3591 2717 3595 2718
rect 3592 2698 3594 2717
rect 3590 2697 3596 2698
rect 3590 2693 3591 2697
rect 3595 2693 3596 2697
rect 3590 2692 3596 2693
rect 3570 2691 3576 2692
rect 3570 2687 3571 2691
rect 3575 2687 3576 2691
rect 3570 2686 3576 2687
rect 3534 2651 3540 2652
rect 3534 2647 3535 2651
rect 3539 2647 3540 2651
rect 3534 2646 3540 2647
rect 2055 2638 2059 2639
rect 2055 2633 2059 2634
rect 2111 2638 2115 2639
rect 2111 2633 2115 2634
rect 2263 2638 2267 2639
rect 2263 2633 2267 2634
rect 2335 2638 2339 2639
rect 2335 2633 2339 2634
rect 2495 2638 2499 2639
rect 2495 2633 2499 2634
rect 2543 2638 2547 2639
rect 2543 2633 2547 2634
rect 2743 2638 2747 2639
rect 2743 2633 2747 2634
rect 2751 2638 2755 2639
rect 2751 2633 2755 2634
rect 2919 2638 2923 2639
rect 2919 2633 2923 2634
rect 3015 2638 3019 2639
rect 3015 2633 3019 2634
rect 3079 2638 3083 2639
rect 3079 2633 3083 2634
rect 3231 2638 3235 2639
rect 3231 2633 3235 2634
rect 3287 2638 3291 2639
rect 3287 2633 3291 2634
rect 3383 2638 3387 2639
rect 3383 2633 3387 2634
rect 3511 2638 3515 2639
rect 3511 2633 3515 2634
rect 1930 2631 1936 2632
rect 1930 2627 1931 2631
rect 1935 2627 1936 2631
rect 1930 2626 1936 2627
rect 1954 2631 1960 2632
rect 1954 2627 1955 2631
rect 1959 2627 1960 2631
rect 1954 2626 1960 2627
rect 1902 2622 1908 2623
rect 1902 2618 1903 2622
rect 1907 2618 1908 2622
rect 1902 2617 1908 2618
rect 1870 2604 1876 2605
rect 1870 2600 1871 2604
rect 1875 2600 1876 2604
rect 1870 2599 1876 2600
rect 1956 2596 1958 2626
rect 2056 2623 2058 2633
rect 2254 2631 2260 2632
rect 2254 2627 2255 2631
rect 2259 2627 2260 2631
rect 2254 2626 2260 2627
rect 2054 2622 2060 2623
rect 2054 2618 2055 2622
rect 2059 2618 2060 2622
rect 2054 2617 2060 2618
rect 2256 2596 2258 2626
rect 2264 2623 2266 2633
rect 2314 2631 2320 2632
rect 2314 2627 2315 2631
rect 2319 2627 2320 2631
rect 2314 2626 2320 2627
rect 2262 2622 2268 2623
rect 2262 2618 2263 2622
rect 2267 2618 2268 2622
rect 2262 2617 2268 2618
rect 2316 2596 2318 2626
rect 2496 2623 2498 2633
rect 2752 2623 2754 2633
rect 3016 2623 3018 2633
rect 3288 2623 3290 2633
rect 3294 2631 3300 2632
rect 3294 2627 3295 2631
rect 3299 2627 3300 2631
rect 3294 2626 3300 2627
rect 3302 2631 3308 2632
rect 3302 2627 3303 2631
rect 3307 2627 3308 2631
rect 3302 2626 3308 2627
rect 2494 2622 2500 2623
rect 2494 2618 2495 2622
rect 2499 2618 2500 2622
rect 2494 2617 2500 2618
rect 2750 2622 2756 2623
rect 2750 2618 2751 2622
rect 2755 2618 2756 2622
rect 2750 2617 2756 2618
rect 3014 2622 3020 2623
rect 3014 2618 3015 2622
rect 3019 2618 3020 2622
rect 3014 2617 3020 2618
rect 3286 2622 3292 2623
rect 3286 2618 3287 2622
rect 3291 2618 3292 2622
rect 3286 2617 3292 2618
rect 3296 2596 3298 2626
rect 1954 2595 1960 2596
rect 1954 2591 1955 2595
rect 1959 2591 1960 2595
rect 1954 2590 1960 2591
rect 2254 2595 2260 2596
rect 2254 2591 2255 2595
rect 2259 2591 2260 2595
rect 2254 2590 2260 2591
rect 2314 2595 2320 2596
rect 2314 2591 2315 2595
rect 2319 2591 2320 2595
rect 2314 2590 2320 2591
rect 3038 2595 3044 2596
rect 3038 2591 3039 2595
rect 3043 2591 3044 2595
rect 3038 2590 3044 2591
rect 3294 2595 3300 2596
rect 3294 2591 3295 2595
rect 3299 2591 3300 2595
rect 3294 2590 3300 2591
rect 1870 2587 1876 2588
rect 1047 2586 1051 2587
rect 1047 2581 1051 2582
rect 1095 2586 1099 2587
rect 1095 2581 1099 2582
rect 1207 2586 1211 2587
rect 1207 2581 1211 2582
rect 1239 2586 1243 2587
rect 1239 2581 1243 2582
rect 1359 2586 1363 2587
rect 1359 2581 1363 2582
rect 1391 2586 1395 2587
rect 1391 2581 1395 2582
rect 1511 2586 1515 2587
rect 1511 2581 1515 2582
rect 1543 2586 1547 2587
rect 1543 2581 1547 2582
rect 1671 2586 1675 2587
rect 1671 2581 1675 2582
rect 1831 2586 1835 2587
rect 1870 2583 1871 2587
rect 1875 2583 1876 2587
rect 1870 2582 1876 2583
rect 1894 2584 1900 2585
rect 1831 2581 1835 2582
rect 1048 2565 1050 2581
rect 1208 2565 1210 2581
rect 1360 2565 1362 2581
rect 1512 2565 1514 2581
rect 1672 2565 1674 2581
rect 1046 2564 1052 2565
rect 1046 2560 1047 2564
rect 1051 2560 1052 2564
rect 1046 2559 1052 2560
rect 1206 2564 1212 2565
rect 1206 2560 1207 2564
rect 1211 2560 1212 2564
rect 1206 2559 1212 2560
rect 1358 2564 1364 2565
rect 1358 2560 1359 2564
rect 1363 2560 1364 2564
rect 1358 2559 1364 2560
rect 1510 2564 1516 2565
rect 1510 2560 1511 2564
rect 1515 2560 1516 2564
rect 1510 2559 1516 2560
rect 1670 2564 1676 2565
rect 1670 2560 1671 2564
rect 1675 2560 1676 2564
rect 1832 2562 1834 2581
rect 1872 2563 1874 2582
rect 1894 2580 1895 2584
rect 1899 2580 1900 2584
rect 1894 2579 1900 2580
rect 2046 2584 2052 2585
rect 2046 2580 2047 2584
rect 2051 2580 2052 2584
rect 2046 2579 2052 2580
rect 2254 2584 2260 2585
rect 2254 2580 2255 2584
rect 2259 2580 2260 2584
rect 2254 2579 2260 2580
rect 2486 2584 2492 2585
rect 2486 2580 2487 2584
rect 2491 2580 2492 2584
rect 2486 2579 2492 2580
rect 2742 2584 2748 2585
rect 2742 2580 2743 2584
rect 2747 2580 2748 2584
rect 2742 2579 2748 2580
rect 3006 2584 3012 2585
rect 3006 2580 3007 2584
rect 3011 2580 3012 2584
rect 3006 2579 3012 2580
rect 1896 2563 1898 2579
rect 2048 2563 2050 2579
rect 2256 2563 2258 2579
rect 2488 2563 2490 2579
rect 2658 2567 2664 2568
rect 2658 2563 2659 2567
rect 2663 2563 2664 2567
rect 2744 2563 2746 2579
rect 3008 2563 3010 2579
rect 1871 2562 1875 2563
rect 1670 2559 1676 2560
rect 1830 2561 1836 2562
rect 1830 2557 1831 2561
rect 1835 2557 1836 2561
rect 1871 2557 1875 2558
rect 1895 2562 1899 2563
rect 1895 2557 1899 2558
rect 2007 2562 2011 2563
rect 2007 2557 2011 2558
rect 2047 2562 2051 2563
rect 2047 2557 2051 2558
rect 2159 2562 2163 2563
rect 2159 2557 2163 2558
rect 2255 2562 2259 2563
rect 2255 2557 2259 2558
rect 2319 2562 2323 2563
rect 2319 2557 2323 2558
rect 2471 2562 2475 2563
rect 2471 2557 2475 2558
rect 2487 2562 2491 2563
rect 2487 2557 2491 2558
rect 2623 2562 2627 2563
rect 2658 2562 2664 2563
rect 2743 2562 2747 2563
rect 2623 2557 2627 2558
rect 1830 2556 1836 2557
rect 594 2555 600 2556
rect 594 2551 595 2555
rect 599 2551 600 2555
rect 594 2550 600 2551
rect 770 2555 776 2556
rect 770 2551 771 2555
rect 775 2551 776 2555
rect 770 2550 776 2551
rect 990 2555 996 2556
rect 990 2551 991 2555
rect 995 2551 996 2555
rect 990 2550 996 2551
rect 1114 2555 1120 2556
rect 1114 2551 1115 2555
rect 1119 2551 1120 2555
rect 1114 2550 1120 2551
rect 1274 2555 1280 2556
rect 1274 2551 1275 2555
rect 1279 2551 1280 2555
rect 1274 2550 1280 2551
rect 1426 2555 1432 2556
rect 1426 2551 1427 2555
rect 1431 2551 1432 2555
rect 1426 2550 1432 2551
rect 1578 2555 1584 2556
rect 1578 2551 1579 2555
rect 1583 2551 1584 2555
rect 1578 2550 1584 2551
rect 586 2547 592 2548
rect 586 2543 587 2547
rect 591 2543 592 2547
rect 586 2542 592 2543
rect 534 2526 540 2527
rect 534 2522 535 2526
rect 539 2522 540 2526
rect 534 2521 540 2522
rect 402 2515 408 2516
rect 402 2511 403 2515
rect 407 2511 408 2515
rect 402 2510 408 2511
rect 536 2507 538 2521
rect 596 2516 598 2550
rect 710 2526 716 2527
rect 710 2522 711 2526
rect 715 2522 716 2526
rect 710 2521 716 2522
rect 594 2515 600 2516
rect 594 2511 595 2515
rect 599 2511 600 2515
rect 594 2510 600 2511
rect 712 2507 714 2521
rect 772 2516 774 2550
rect 886 2526 892 2527
rect 886 2522 887 2526
rect 891 2522 892 2526
rect 886 2521 892 2522
rect 1054 2526 1060 2527
rect 1054 2522 1055 2526
rect 1059 2522 1060 2526
rect 1054 2521 1060 2522
rect 770 2515 776 2516
rect 770 2511 771 2515
rect 775 2511 776 2515
rect 770 2510 776 2511
rect 888 2507 890 2521
rect 934 2515 940 2516
rect 934 2511 935 2515
rect 939 2511 940 2515
rect 934 2510 940 2511
rect 223 2506 227 2507
rect 223 2501 227 2502
rect 231 2506 235 2507
rect 231 2501 235 2502
rect 303 2506 307 2507
rect 303 2501 307 2502
rect 375 2506 379 2507
rect 375 2501 379 2502
rect 391 2506 395 2507
rect 391 2501 395 2502
rect 511 2506 515 2507
rect 511 2501 515 2502
rect 535 2506 539 2507
rect 535 2501 539 2502
rect 647 2506 651 2507
rect 647 2501 651 2502
rect 711 2506 715 2507
rect 711 2501 715 2502
rect 783 2506 787 2507
rect 783 2501 787 2502
rect 887 2506 891 2507
rect 887 2501 891 2502
rect 927 2506 931 2507
rect 927 2501 931 2502
rect 194 2499 200 2500
rect 194 2495 195 2499
rect 199 2495 200 2499
rect 194 2494 200 2495
rect 214 2499 220 2500
rect 214 2495 215 2499
rect 219 2495 220 2499
rect 214 2494 220 2495
rect 142 2490 148 2491
rect 142 2486 143 2490
rect 147 2486 148 2490
rect 142 2485 148 2486
rect 110 2472 116 2473
rect 110 2468 111 2472
rect 115 2468 116 2472
rect 110 2467 116 2468
rect 216 2464 218 2494
rect 224 2491 226 2501
rect 274 2499 280 2500
rect 274 2495 275 2499
rect 279 2495 280 2499
rect 274 2494 280 2495
rect 222 2490 228 2491
rect 222 2486 223 2490
rect 227 2486 228 2490
rect 222 2485 228 2486
rect 276 2464 278 2494
rect 304 2491 306 2501
rect 354 2499 360 2500
rect 354 2495 355 2499
rect 359 2495 360 2499
rect 354 2494 360 2495
rect 302 2490 308 2491
rect 302 2486 303 2490
rect 307 2486 308 2490
rect 302 2485 308 2486
rect 356 2464 358 2494
rect 392 2491 394 2501
rect 442 2499 448 2500
rect 442 2495 443 2499
rect 447 2495 448 2499
rect 442 2494 448 2495
rect 390 2490 396 2491
rect 390 2486 391 2490
rect 395 2486 396 2490
rect 390 2485 396 2486
rect 444 2464 446 2494
rect 512 2491 514 2501
rect 562 2499 568 2500
rect 562 2495 563 2499
rect 567 2495 568 2499
rect 562 2494 568 2495
rect 510 2490 516 2491
rect 510 2486 511 2490
rect 515 2486 516 2490
rect 510 2485 516 2486
rect 564 2464 566 2494
rect 648 2491 650 2501
rect 698 2499 704 2500
rect 698 2495 699 2499
rect 703 2495 704 2499
rect 698 2494 704 2495
rect 646 2490 652 2491
rect 646 2486 647 2490
rect 651 2486 652 2490
rect 646 2485 652 2486
rect 700 2464 702 2494
rect 784 2491 786 2501
rect 834 2499 840 2500
rect 834 2495 835 2499
rect 839 2495 840 2499
rect 834 2494 840 2495
rect 782 2490 788 2491
rect 782 2486 783 2490
rect 787 2486 788 2490
rect 782 2485 788 2486
rect 836 2464 838 2494
rect 928 2491 930 2501
rect 926 2490 932 2491
rect 926 2486 927 2490
rect 931 2486 932 2490
rect 926 2485 932 2486
rect 936 2464 938 2510
rect 1056 2507 1058 2521
rect 1116 2516 1118 2550
rect 1214 2526 1220 2527
rect 1214 2522 1215 2526
rect 1219 2522 1220 2526
rect 1214 2521 1220 2522
rect 1114 2515 1120 2516
rect 1114 2511 1115 2515
rect 1119 2511 1120 2515
rect 1114 2510 1120 2511
rect 1216 2507 1218 2521
rect 1276 2516 1278 2550
rect 1366 2526 1372 2527
rect 1366 2522 1367 2526
rect 1371 2522 1372 2526
rect 1366 2521 1372 2522
rect 1274 2515 1280 2516
rect 1274 2511 1275 2515
rect 1279 2511 1280 2515
rect 1274 2510 1280 2511
rect 1368 2507 1370 2521
rect 1428 2516 1430 2550
rect 1518 2526 1524 2527
rect 1518 2522 1519 2526
rect 1523 2522 1524 2526
rect 1518 2521 1524 2522
rect 1426 2515 1432 2516
rect 1426 2511 1427 2515
rect 1431 2511 1432 2515
rect 1426 2510 1432 2511
rect 1520 2507 1522 2521
rect 1580 2516 1582 2550
rect 1830 2544 1836 2545
rect 1830 2540 1831 2544
rect 1835 2540 1836 2544
rect 1830 2539 1836 2540
rect 1678 2526 1684 2527
rect 1678 2522 1679 2526
rect 1683 2522 1684 2526
rect 1678 2521 1684 2522
rect 1578 2515 1584 2516
rect 1578 2511 1579 2515
rect 1583 2511 1584 2515
rect 1578 2510 1584 2511
rect 1680 2507 1682 2521
rect 1702 2515 1708 2516
rect 1702 2511 1703 2515
rect 1707 2511 1708 2515
rect 1702 2510 1708 2511
rect 1055 2506 1059 2507
rect 1055 2501 1059 2502
rect 1063 2506 1067 2507
rect 1063 2501 1067 2502
rect 1191 2506 1195 2507
rect 1191 2501 1195 2502
rect 1215 2506 1219 2507
rect 1215 2501 1219 2502
rect 1311 2506 1315 2507
rect 1311 2501 1315 2502
rect 1367 2506 1371 2507
rect 1367 2501 1371 2502
rect 1431 2506 1435 2507
rect 1431 2501 1435 2502
rect 1519 2506 1523 2507
rect 1519 2501 1523 2502
rect 1551 2506 1555 2507
rect 1551 2501 1555 2502
rect 1671 2506 1675 2507
rect 1671 2501 1675 2502
rect 1679 2506 1683 2507
rect 1679 2501 1683 2502
rect 1064 2491 1066 2501
rect 1134 2499 1140 2500
rect 1134 2495 1135 2499
rect 1139 2495 1140 2499
rect 1134 2494 1140 2495
rect 1142 2499 1148 2500
rect 1142 2495 1143 2499
rect 1147 2495 1148 2499
rect 1142 2494 1148 2495
rect 1062 2490 1068 2491
rect 1062 2486 1063 2490
rect 1067 2486 1068 2490
rect 1062 2485 1068 2486
rect 214 2463 220 2464
rect 214 2459 215 2463
rect 219 2459 220 2463
rect 214 2458 220 2459
rect 274 2463 280 2464
rect 274 2459 275 2463
rect 279 2459 280 2463
rect 274 2458 280 2459
rect 354 2463 360 2464
rect 354 2459 355 2463
rect 359 2459 360 2463
rect 354 2458 360 2459
rect 442 2463 448 2464
rect 442 2459 443 2463
rect 447 2459 448 2463
rect 442 2458 448 2459
rect 562 2463 568 2464
rect 562 2459 563 2463
rect 567 2459 568 2463
rect 562 2458 568 2459
rect 698 2463 704 2464
rect 698 2459 699 2463
rect 703 2459 704 2463
rect 698 2458 704 2459
rect 834 2463 840 2464
rect 834 2459 835 2463
rect 839 2459 840 2463
rect 834 2458 840 2459
rect 934 2463 940 2464
rect 934 2459 935 2463
rect 939 2459 940 2463
rect 1136 2461 1138 2494
rect 1144 2464 1146 2494
rect 1192 2491 1194 2501
rect 1242 2499 1248 2500
rect 1242 2495 1243 2499
rect 1247 2495 1248 2499
rect 1242 2494 1248 2495
rect 1190 2490 1196 2491
rect 1190 2486 1191 2490
rect 1195 2486 1196 2490
rect 1190 2485 1196 2486
rect 1244 2464 1246 2494
rect 1312 2491 1314 2501
rect 1422 2499 1428 2500
rect 1422 2495 1423 2499
rect 1427 2495 1428 2499
rect 1422 2494 1428 2495
rect 1310 2490 1316 2491
rect 1310 2486 1311 2490
rect 1315 2486 1316 2490
rect 1310 2485 1316 2486
rect 1424 2464 1426 2494
rect 1432 2491 1434 2501
rect 1482 2499 1488 2500
rect 1482 2495 1483 2499
rect 1487 2495 1488 2499
rect 1482 2494 1488 2495
rect 1430 2490 1436 2491
rect 1430 2486 1431 2490
rect 1435 2486 1436 2490
rect 1430 2485 1436 2486
rect 1484 2464 1486 2494
rect 1552 2491 1554 2501
rect 1602 2499 1608 2500
rect 1602 2495 1603 2499
rect 1607 2495 1608 2499
rect 1602 2494 1608 2495
rect 1550 2490 1556 2491
rect 1550 2486 1551 2490
rect 1555 2486 1556 2490
rect 1550 2485 1556 2486
rect 1604 2464 1606 2494
rect 1672 2491 1674 2501
rect 1670 2490 1676 2491
rect 1670 2486 1671 2490
rect 1675 2486 1676 2490
rect 1670 2485 1676 2486
rect 1704 2464 1706 2510
rect 1832 2507 1834 2539
rect 1872 2538 1874 2557
rect 1896 2541 1898 2557
rect 2008 2541 2010 2557
rect 2160 2541 2162 2557
rect 2320 2541 2322 2557
rect 2472 2541 2474 2557
rect 2624 2541 2626 2557
rect 1894 2540 1900 2541
rect 1870 2537 1876 2538
rect 1870 2533 1871 2537
rect 1875 2533 1876 2537
rect 1894 2536 1895 2540
rect 1899 2536 1900 2540
rect 1894 2535 1900 2536
rect 2006 2540 2012 2541
rect 2006 2536 2007 2540
rect 2011 2536 2012 2540
rect 2006 2535 2012 2536
rect 2158 2540 2164 2541
rect 2158 2536 2159 2540
rect 2163 2536 2164 2540
rect 2158 2535 2164 2536
rect 2318 2540 2324 2541
rect 2318 2536 2319 2540
rect 2323 2536 2324 2540
rect 2318 2535 2324 2536
rect 2470 2540 2476 2541
rect 2470 2536 2471 2540
rect 2475 2536 2476 2540
rect 2470 2535 2476 2536
rect 2622 2540 2628 2541
rect 2622 2536 2623 2540
rect 2627 2536 2628 2540
rect 2622 2535 2628 2536
rect 2660 2533 2662 2562
rect 2743 2557 2747 2558
rect 2759 2562 2763 2563
rect 2759 2557 2763 2558
rect 2887 2562 2891 2563
rect 2887 2557 2891 2558
rect 3007 2562 3011 2563
rect 3007 2557 3011 2558
rect 2760 2541 2762 2557
rect 2888 2541 2890 2557
rect 3008 2541 3010 2557
rect 2758 2540 2764 2541
rect 2758 2536 2759 2540
rect 2763 2536 2764 2540
rect 2758 2535 2764 2536
rect 2886 2540 2892 2541
rect 2886 2536 2887 2540
rect 2891 2536 2892 2540
rect 2886 2535 2892 2536
rect 3006 2540 3012 2541
rect 3006 2536 3007 2540
rect 3011 2536 3012 2540
rect 3006 2535 3012 2536
rect 1870 2532 1876 2533
rect 1931 2532 1935 2533
rect 2659 2532 2663 2533
rect 1931 2527 1935 2528
rect 1962 2531 1968 2532
rect 1962 2527 1963 2531
rect 1967 2527 1968 2531
rect 1870 2520 1876 2521
rect 1870 2516 1871 2520
rect 1875 2516 1876 2520
rect 1870 2515 1876 2516
rect 1831 2506 1835 2507
rect 1831 2501 1835 2502
rect 1832 2473 1834 2501
rect 1872 2479 1874 2515
rect 1902 2502 1908 2503
rect 1902 2498 1903 2502
rect 1907 2498 1908 2502
rect 1902 2497 1908 2498
rect 1904 2479 1906 2497
rect 1932 2492 1934 2527
rect 1962 2526 1968 2527
rect 2106 2531 2112 2532
rect 2106 2527 2107 2531
rect 2111 2527 2112 2531
rect 2106 2526 2112 2527
rect 2262 2531 2268 2532
rect 2262 2527 2263 2531
rect 2267 2527 2268 2531
rect 2262 2526 2268 2527
rect 2418 2531 2424 2532
rect 2418 2527 2419 2531
rect 2423 2527 2424 2531
rect 2418 2526 2424 2527
rect 2426 2531 2432 2532
rect 2426 2527 2427 2531
rect 2431 2527 2432 2531
rect 2659 2527 2663 2528
rect 2714 2531 2720 2532
rect 2714 2527 2715 2531
rect 2719 2527 2720 2531
rect 2426 2526 2432 2527
rect 2714 2526 2720 2527
rect 2954 2531 2960 2532
rect 2954 2527 2955 2531
rect 2959 2527 2960 2531
rect 2954 2526 2960 2527
rect 1964 2492 1966 2526
rect 2014 2502 2020 2503
rect 2014 2498 2015 2502
rect 2019 2498 2020 2502
rect 2014 2497 2020 2498
rect 1930 2491 1936 2492
rect 1930 2487 1931 2491
rect 1935 2487 1936 2491
rect 1930 2486 1936 2487
rect 1962 2491 1968 2492
rect 1962 2487 1963 2491
rect 1967 2487 1968 2491
rect 1962 2486 1968 2487
rect 2016 2479 2018 2497
rect 2108 2492 2110 2526
rect 2166 2502 2172 2503
rect 2166 2498 2167 2502
rect 2171 2498 2172 2502
rect 2166 2497 2172 2498
rect 2106 2491 2112 2492
rect 2106 2487 2107 2491
rect 2111 2487 2112 2491
rect 2106 2486 2112 2487
rect 2168 2479 2170 2497
rect 2264 2492 2266 2526
rect 2326 2502 2332 2503
rect 2326 2498 2327 2502
rect 2331 2498 2332 2502
rect 2326 2497 2332 2498
rect 2262 2491 2268 2492
rect 2262 2487 2263 2491
rect 2267 2487 2268 2491
rect 2262 2486 2268 2487
rect 2328 2479 2330 2497
rect 2420 2492 2422 2526
rect 2418 2491 2424 2492
rect 2418 2487 2419 2491
rect 2423 2487 2424 2491
rect 2418 2486 2424 2487
rect 2428 2480 2430 2526
rect 2682 2523 2688 2524
rect 2682 2519 2683 2523
rect 2687 2519 2688 2523
rect 2682 2518 2688 2519
rect 2478 2502 2484 2503
rect 2478 2498 2479 2502
rect 2483 2498 2484 2502
rect 2478 2497 2484 2498
rect 2630 2502 2636 2503
rect 2630 2498 2631 2502
rect 2635 2498 2636 2502
rect 2630 2497 2636 2498
rect 2426 2479 2432 2480
rect 2480 2479 2482 2497
rect 2632 2479 2634 2497
rect 2684 2492 2686 2518
rect 2716 2492 2718 2526
rect 2766 2502 2772 2503
rect 2766 2498 2767 2502
rect 2771 2498 2772 2502
rect 2766 2497 2772 2498
rect 2894 2502 2900 2503
rect 2894 2498 2895 2502
rect 2899 2498 2900 2502
rect 2894 2497 2900 2498
rect 2682 2491 2688 2492
rect 2682 2487 2683 2491
rect 2687 2487 2688 2491
rect 2682 2486 2688 2487
rect 2714 2491 2720 2492
rect 2714 2487 2715 2491
rect 2719 2487 2720 2491
rect 2714 2486 2720 2487
rect 2768 2479 2770 2497
rect 2896 2479 2898 2497
rect 2956 2492 2958 2526
rect 3014 2502 3020 2503
rect 3014 2498 3015 2502
rect 3019 2498 3020 2502
rect 3014 2497 3020 2498
rect 2954 2491 2960 2492
rect 2954 2487 2955 2491
rect 2959 2487 2960 2491
rect 2954 2486 2960 2487
rect 3016 2479 3018 2497
rect 3040 2492 3042 2590
rect 3278 2584 3284 2585
rect 3278 2580 3279 2584
rect 3283 2580 3284 2584
rect 3278 2579 3284 2580
rect 3280 2563 3282 2579
rect 3119 2562 3123 2563
rect 3119 2557 3123 2558
rect 3223 2562 3227 2563
rect 3223 2557 3227 2558
rect 3279 2562 3283 2563
rect 3279 2557 3283 2558
rect 3120 2541 3122 2557
rect 3224 2541 3226 2557
rect 3118 2540 3124 2541
rect 3118 2536 3119 2540
rect 3123 2536 3124 2540
rect 3118 2535 3124 2536
rect 3222 2540 3228 2541
rect 3222 2536 3223 2540
rect 3227 2536 3228 2540
rect 3222 2535 3228 2536
rect 3074 2531 3080 2532
rect 3074 2527 3075 2531
rect 3079 2527 3080 2531
rect 3074 2526 3080 2527
rect 3290 2531 3296 2532
rect 3290 2527 3291 2531
rect 3295 2527 3296 2531
rect 3290 2526 3296 2527
rect 3038 2491 3044 2492
rect 3038 2487 3039 2491
rect 3043 2487 3044 2491
rect 3038 2486 3044 2487
rect 1871 2478 1875 2479
rect 1871 2473 1875 2474
rect 1903 2478 1907 2479
rect 1903 2473 1907 2474
rect 1999 2478 2003 2479
rect 1999 2473 2003 2474
rect 2015 2478 2019 2479
rect 2015 2473 2019 2474
rect 2127 2478 2131 2479
rect 2127 2473 2131 2474
rect 2167 2478 2171 2479
rect 2167 2473 2171 2474
rect 2263 2478 2267 2479
rect 2263 2473 2267 2474
rect 2327 2478 2331 2479
rect 2327 2473 2331 2474
rect 2407 2478 2411 2479
rect 2426 2475 2427 2479
rect 2431 2475 2432 2479
rect 2426 2474 2432 2475
rect 2479 2478 2483 2479
rect 2407 2473 2411 2474
rect 2479 2473 2483 2474
rect 2551 2478 2555 2479
rect 2551 2473 2555 2474
rect 2631 2478 2635 2479
rect 2631 2473 2635 2474
rect 2703 2478 2707 2479
rect 2703 2473 2707 2474
rect 2767 2478 2771 2479
rect 2767 2473 2771 2474
rect 2863 2478 2867 2479
rect 2863 2473 2867 2474
rect 2895 2478 2899 2479
rect 2895 2473 2899 2474
rect 3015 2478 3019 2479
rect 3015 2473 3019 2474
rect 3023 2478 3027 2479
rect 3023 2473 3027 2474
rect 1830 2472 1836 2473
rect 1830 2468 1831 2472
rect 1835 2468 1836 2472
rect 1830 2467 1836 2468
rect 1142 2463 1148 2464
rect 934 2458 940 2459
rect 1135 2460 1139 2461
rect 1142 2459 1143 2463
rect 1147 2459 1148 2463
rect 1142 2458 1148 2459
rect 1242 2463 1248 2464
rect 1242 2459 1243 2463
rect 1247 2459 1248 2463
rect 1242 2458 1248 2459
rect 1422 2463 1428 2464
rect 1422 2459 1423 2463
rect 1427 2459 1428 2463
rect 1482 2463 1488 2464
rect 1422 2458 1428 2459
rect 1471 2460 1475 2461
rect 110 2455 116 2456
rect 1135 2455 1139 2456
rect 1482 2459 1483 2463
rect 1487 2459 1488 2463
rect 1482 2458 1488 2459
rect 1602 2463 1608 2464
rect 1602 2459 1603 2463
rect 1607 2459 1608 2463
rect 1602 2458 1608 2459
rect 1702 2463 1708 2464
rect 1702 2459 1703 2463
rect 1707 2459 1708 2463
rect 1702 2458 1708 2459
rect 1471 2455 1475 2456
rect 1830 2455 1836 2456
rect 110 2451 111 2455
rect 115 2451 116 2455
rect 110 2450 116 2451
rect 134 2452 140 2453
rect 112 2419 114 2450
rect 134 2448 135 2452
rect 139 2448 140 2452
rect 134 2447 140 2448
rect 214 2452 220 2453
rect 214 2448 215 2452
rect 219 2448 220 2452
rect 214 2447 220 2448
rect 294 2452 300 2453
rect 294 2448 295 2452
rect 299 2448 300 2452
rect 294 2447 300 2448
rect 382 2452 388 2453
rect 382 2448 383 2452
rect 387 2448 388 2452
rect 382 2447 388 2448
rect 502 2452 508 2453
rect 502 2448 503 2452
rect 507 2448 508 2452
rect 502 2447 508 2448
rect 638 2452 644 2453
rect 638 2448 639 2452
rect 643 2448 644 2452
rect 638 2447 644 2448
rect 774 2452 780 2453
rect 774 2448 775 2452
rect 779 2448 780 2452
rect 774 2447 780 2448
rect 918 2452 924 2453
rect 918 2448 919 2452
rect 923 2448 924 2452
rect 918 2447 924 2448
rect 1054 2452 1060 2453
rect 1054 2448 1055 2452
rect 1059 2448 1060 2452
rect 1054 2447 1060 2448
rect 1182 2452 1188 2453
rect 1182 2448 1183 2452
rect 1187 2448 1188 2452
rect 1182 2447 1188 2448
rect 1302 2452 1308 2453
rect 1302 2448 1303 2452
rect 1307 2448 1308 2452
rect 1302 2447 1308 2448
rect 1422 2452 1428 2453
rect 1422 2448 1423 2452
rect 1427 2448 1428 2452
rect 1422 2447 1428 2448
rect 136 2419 138 2447
rect 216 2419 218 2447
rect 296 2419 298 2447
rect 384 2419 386 2447
rect 504 2419 506 2447
rect 640 2419 642 2447
rect 776 2419 778 2447
rect 920 2419 922 2447
rect 1056 2419 1058 2447
rect 1184 2419 1186 2447
rect 1304 2419 1306 2447
rect 1424 2419 1426 2447
rect 111 2418 115 2419
rect 111 2413 115 2414
rect 135 2418 139 2419
rect 135 2413 139 2414
rect 215 2418 219 2419
rect 215 2413 219 2414
rect 295 2418 299 2419
rect 295 2413 299 2414
rect 383 2418 387 2419
rect 383 2413 387 2414
rect 503 2418 507 2419
rect 503 2413 507 2414
rect 639 2418 643 2419
rect 639 2413 643 2414
rect 775 2418 779 2419
rect 775 2413 779 2414
rect 919 2418 923 2419
rect 919 2413 923 2414
rect 1055 2418 1059 2419
rect 1055 2413 1059 2414
rect 1063 2418 1067 2419
rect 1063 2413 1067 2414
rect 1143 2418 1147 2419
rect 1143 2413 1147 2414
rect 1183 2418 1187 2419
rect 1183 2413 1187 2414
rect 1223 2418 1227 2419
rect 1223 2413 1227 2414
rect 1303 2418 1307 2419
rect 1303 2413 1307 2414
rect 1383 2418 1387 2419
rect 1383 2413 1387 2414
rect 1423 2418 1427 2419
rect 1423 2413 1427 2414
rect 1463 2418 1467 2419
rect 1463 2413 1467 2414
rect 112 2394 114 2413
rect 1064 2397 1066 2413
rect 1144 2397 1146 2413
rect 1224 2397 1226 2413
rect 1304 2397 1306 2413
rect 1384 2397 1386 2413
rect 1464 2397 1466 2413
rect 1062 2396 1068 2397
rect 110 2393 116 2394
rect 110 2389 111 2393
rect 115 2389 116 2393
rect 1062 2392 1063 2396
rect 1067 2392 1068 2396
rect 1062 2391 1068 2392
rect 1142 2396 1148 2397
rect 1142 2392 1143 2396
rect 1147 2392 1148 2396
rect 1142 2391 1148 2392
rect 1222 2396 1228 2397
rect 1222 2392 1223 2396
rect 1227 2392 1228 2396
rect 1222 2391 1228 2392
rect 1302 2396 1308 2397
rect 1302 2392 1303 2396
rect 1307 2392 1308 2396
rect 1302 2391 1308 2392
rect 1382 2396 1388 2397
rect 1382 2392 1383 2396
rect 1387 2392 1388 2396
rect 1382 2391 1388 2392
rect 1462 2396 1468 2397
rect 1462 2392 1463 2396
rect 1467 2392 1468 2396
rect 1462 2391 1468 2392
rect 110 2388 116 2389
rect 1134 2387 1140 2388
rect 1134 2383 1135 2387
rect 1139 2383 1140 2387
rect 1134 2382 1140 2383
rect 1210 2387 1216 2388
rect 1210 2383 1211 2387
rect 1215 2383 1216 2387
rect 1210 2382 1216 2383
rect 1290 2387 1296 2388
rect 1290 2383 1291 2387
rect 1295 2383 1296 2387
rect 1290 2382 1296 2383
rect 1370 2387 1376 2388
rect 1370 2383 1371 2387
rect 1375 2383 1376 2387
rect 1370 2382 1376 2383
rect 1450 2387 1456 2388
rect 1450 2383 1451 2387
rect 1455 2383 1456 2387
rect 1472 2384 1474 2455
rect 1542 2452 1548 2453
rect 1542 2448 1543 2452
rect 1547 2448 1548 2452
rect 1542 2447 1548 2448
rect 1662 2452 1668 2453
rect 1662 2448 1663 2452
rect 1667 2448 1668 2452
rect 1830 2451 1831 2455
rect 1835 2451 1836 2455
rect 1830 2450 1836 2451
rect 1662 2447 1668 2448
rect 1544 2419 1546 2447
rect 1664 2419 1666 2447
rect 1832 2419 1834 2450
rect 1872 2445 1874 2473
rect 2000 2463 2002 2473
rect 2050 2471 2056 2472
rect 2050 2467 2051 2471
rect 2055 2467 2056 2471
rect 2050 2466 2056 2467
rect 1998 2462 2004 2463
rect 1998 2458 1999 2462
rect 2003 2458 2004 2462
rect 1998 2457 2004 2458
rect 1870 2444 1876 2445
rect 1870 2440 1871 2444
rect 1875 2440 1876 2444
rect 1870 2439 1876 2440
rect 2052 2436 2054 2466
rect 2128 2463 2130 2473
rect 2178 2471 2184 2472
rect 2178 2467 2179 2471
rect 2183 2467 2184 2471
rect 2178 2466 2184 2467
rect 2126 2462 2132 2463
rect 2126 2458 2127 2462
rect 2131 2458 2132 2462
rect 2126 2457 2132 2458
rect 2180 2436 2182 2466
rect 2264 2463 2266 2473
rect 2314 2471 2320 2472
rect 2314 2467 2315 2471
rect 2319 2467 2320 2471
rect 2314 2466 2320 2467
rect 2262 2462 2268 2463
rect 2262 2458 2263 2462
rect 2267 2458 2268 2462
rect 2262 2457 2268 2458
rect 2316 2436 2318 2466
rect 2408 2463 2410 2473
rect 2458 2471 2464 2472
rect 2458 2467 2459 2471
rect 2463 2467 2464 2471
rect 2458 2466 2464 2467
rect 2406 2462 2412 2463
rect 2406 2458 2407 2462
rect 2411 2458 2412 2462
rect 2406 2457 2412 2458
rect 2460 2436 2462 2466
rect 2552 2463 2554 2473
rect 2704 2463 2706 2473
rect 2802 2471 2808 2472
rect 2802 2467 2803 2471
rect 2807 2467 2808 2471
rect 2802 2466 2808 2467
rect 2810 2471 2816 2472
rect 2810 2467 2811 2471
rect 2815 2467 2816 2471
rect 2810 2466 2816 2467
rect 2550 2462 2556 2463
rect 2550 2458 2551 2462
rect 2555 2458 2556 2462
rect 2550 2457 2556 2458
rect 2702 2462 2708 2463
rect 2702 2458 2703 2462
rect 2707 2458 2708 2462
rect 2804 2461 2806 2466
rect 2702 2457 2708 2458
rect 2803 2460 2807 2461
rect 2803 2455 2807 2456
rect 2812 2436 2814 2466
rect 2864 2463 2866 2473
rect 3024 2463 3026 2473
rect 3076 2472 3078 2526
rect 3126 2502 3132 2503
rect 3126 2498 3127 2502
rect 3131 2498 3132 2502
rect 3126 2497 3132 2498
rect 3230 2502 3236 2503
rect 3230 2498 3231 2502
rect 3235 2498 3236 2502
rect 3230 2497 3236 2498
rect 3128 2479 3130 2497
rect 3232 2479 3234 2497
rect 3292 2492 3294 2526
rect 3304 2524 3306 2626
rect 3319 2562 3323 2563
rect 3319 2557 3323 2558
rect 3423 2562 3427 2563
rect 3423 2557 3427 2558
rect 3503 2562 3507 2563
rect 3503 2557 3507 2558
rect 3320 2541 3322 2557
rect 3424 2541 3426 2557
rect 3504 2541 3506 2557
rect 3318 2540 3324 2541
rect 3318 2536 3319 2540
rect 3323 2536 3324 2540
rect 3318 2535 3324 2536
rect 3422 2540 3428 2541
rect 3422 2536 3423 2540
rect 3427 2536 3428 2540
rect 3422 2535 3428 2536
rect 3502 2540 3508 2541
rect 3502 2536 3503 2540
rect 3507 2536 3508 2540
rect 3502 2535 3508 2536
rect 3386 2531 3392 2532
rect 3386 2527 3387 2531
rect 3391 2527 3392 2531
rect 3386 2526 3392 2527
rect 3302 2523 3308 2524
rect 3302 2519 3303 2523
rect 3307 2519 3308 2523
rect 3302 2518 3308 2519
rect 3326 2502 3332 2503
rect 3326 2498 3327 2502
rect 3331 2498 3332 2502
rect 3326 2497 3332 2498
rect 3290 2491 3296 2492
rect 3290 2487 3291 2491
rect 3295 2487 3296 2491
rect 3290 2486 3296 2487
rect 3328 2479 3330 2497
rect 3388 2492 3390 2526
rect 3562 2523 3568 2524
rect 3562 2519 3563 2523
rect 3567 2519 3568 2523
rect 3562 2518 3568 2519
rect 3430 2502 3436 2503
rect 3430 2498 3431 2502
rect 3435 2498 3436 2502
rect 3430 2497 3436 2498
rect 3510 2502 3516 2503
rect 3510 2498 3511 2502
rect 3515 2498 3516 2502
rect 3510 2497 3516 2498
rect 3386 2491 3392 2492
rect 3386 2487 3387 2491
rect 3391 2487 3392 2491
rect 3386 2486 3392 2487
rect 3410 2491 3416 2492
rect 3410 2487 3411 2491
rect 3415 2487 3416 2491
rect 3410 2486 3416 2487
rect 3127 2478 3131 2479
rect 3127 2473 3131 2474
rect 3191 2478 3195 2479
rect 3191 2473 3195 2474
rect 3231 2478 3235 2479
rect 3231 2473 3235 2474
rect 3327 2478 3331 2479
rect 3327 2473 3331 2474
rect 3359 2478 3363 2479
rect 3359 2473 3363 2474
rect 3074 2471 3080 2472
rect 3074 2467 3075 2471
rect 3079 2467 3080 2471
rect 3074 2466 3080 2467
rect 3192 2463 3194 2473
rect 3360 2463 3362 2473
rect 2862 2462 2868 2463
rect 2862 2458 2863 2462
rect 2867 2458 2868 2462
rect 2862 2457 2868 2458
rect 3022 2462 3028 2463
rect 3022 2458 3023 2462
rect 3027 2458 3028 2462
rect 3022 2457 3028 2458
rect 3190 2462 3196 2463
rect 3190 2458 3191 2462
rect 3195 2458 3196 2462
rect 3358 2462 3364 2463
rect 3190 2457 3196 2458
rect 3199 2460 3203 2461
rect 3358 2458 3359 2462
rect 3363 2458 3364 2462
rect 3358 2457 3364 2458
rect 3199 2455 3203 2456
rect 3200 2436 3202 2455
rect 3412 2436 3414 2486
rect 3432 2479 3434 2497
rect 3512 2479 3514 2497
rect 3431 2478 3435 2479
rect 3431 2473 3435 2474
rect 3511 2478 3515 2479
rect 3511 2473 3515 2474
rect 3418 2471 3424 2472
rect 3418 2467 3419 2471
rect 3423 2467 3424 2471
rect 3418 2466 3424 2467
rect 2050 2435 2056 2436
rect 2050 2431 2051 2435
rect 2055 2431 2056 2435
rect 2050 2430 2056 2431
rect 2178 2435 2184 2436
rect 2178 2431 2179 2435
rect 2183 2431 2184 2435
rect 2178 2430 2184 2431
rect 2314 2435 2320 2436
rect 2314 2431 2315 2435
rect 2319 2431 2320 2435
rect 2314 2430 2320 2431
rect 2458 2435 2464 2436
rect 2458 2431 2459 2435
rect 2463 2431 2464 2435
rect 2458 2430 2464 2431
rect 2810 2435 2816 2436
rect 2810 2431 2811 2435
rect 2815 2431 2816 2435
rect 2810 2430 2816 2431
rect 2914 2435 2920 2436
rect 2914 2431 2915 2435
rect 2919 2431 2920 2435
rect 2914 2430 2920 2431
rect 3198 2435 3204 2436
rect 3198 2431 3199 2435
rect 3203 2431 3204 2435
rect 3198 2430 3204 2431
rect 3410 2435 3416 2436
rect 3410 2431 3411 2435
rect 3415 2431 3416 2435
rect 3410 2430 3416 2431
rect 1870 2427 1876 2428
rect 1870 2423 1871 2427
rect 1875 2423 1876 2427
rect 1870 2422 1876 2423
rect 1990 2424 1996 2425
rect 1543 2418 1547 2419
rect 1543 2413 1547 2414
rect 1663 2418 1667 2419
rect 1663 2413 1667 2414
rect 1831 2418 1835 2419
rect 1831 2413 1835 2414
rect 1832 2394 1834 2413
rect 1872 2399 1874 2422
rect 1990 2420 1991 2424
rect 1995 2420 1996 2424
rect 1990 2419 1996 2420
rect 2118 2424 2124 2425
rect 2118 2420 2119 2424
rect 2123 2420 2124 2424
rect 2118 2419 2124 2420
rect 2254 2424 2260 2425
rect 2254 2420 2255 2424
rect 2259 2420 2260 2424
rect 2254 2419 2260 2420
rect 2398 2424 2404 2425
rect 2398 2420 2399 2424
rect 2403 2420 2404 2424
rect 2398 2419 2404 2420
rect 2542 2424 2548 2425
rect 2542 2420 2543 2424
rect 2547 2420 2548 2424
rect 2542 2419 2548 2420
rect 2694 2424 2700 2425
rect 2694 2420 2695 2424
rect 2699 2420 2700 2424
rect 2694 2419 2700 2420
rect 2854 2424 2860 2425
rect 2854 2420 2855 2424
rect 2859 2420 2860 2424
rect 2854 2419 2860 2420
rect 1992 2399 1994 2419
rect 2120 2399 2122 2419
rect 2256 2399 2258 2419
rect 2400 2399 2402 2419
rect 2478 2407 2484 2408
rect 2478 2403 2479 2407
rect 2483 2403 2484 2407
rect 2478 2402 2484 2403
rect 1871 2398 1875 2399
rect 1830 2393 1836 2394
rect 1871 2393 1875 2394
rect 1991 2398 1995 2399
rect 1991 2393 1995 2394
rect 2119 2398 2123 2399
rect 2119 2393 2123 2394
rect 2143 2398 2147 2399
rect 2143 2393 2147 2394
rect 2239 2398 2243 2399
rect 2239 2393 2243 2394
rect 2255 2398 2259 2399
rect 2255 2393 2259 2394
rect 2343 2398 2347 2399
rect 2343 2393 2347 2394
rect 2399 2398 2403 2399
rect 2399 2393 2403 2394
rect 2455 2398 2459 2399
rect 2455 2393 2459 2394
rect 1830 2389 1831 2393
rect 1835 2389 1836 2393
rect 1830 2388 1836 2389
rect 1450 2382 1456 2383
rect 1470 2383 1476 2384
rect 110 2376 116 2377
rect 110 2372 111 2376
rect 115 2372 116 2376
rect 110 2371 116 2372
rect 112 2335 114 2371
rect 1070 2358 1076 2359
rect 1070 2354 1071 2358
rect 1075 2354 1076 2358
rect 1070 2353 1076 2354
rect 926 2335 932 2336
rect 1072 2335 1074 2353
rect 1136 2348 1138 2382
rect 1150 2358 1156 2359
rect 1150 2354 1151 2358
rect 1155 2354 1156 2358
rect 1150 2353 1156 2354
rect 1134 2347 1140 2348
rect 1134 2343 1135 2347
rect 1139 2343 1140 2347
rect 1134 2342 1140 2343
rect 1152 2335 1154 2353
rect 1212 2348 1214 2382
rect 1230 2358 1236 2359
rect 1230 2354 1231 2358
rect 1235 2354 1236 2358
rect 1230 2353 1236 2354
rect 1210 2347 1216 2348
rect 1210 2343 1211 2347
rect 1215 2343 1216 2347
rect 1210 2342 1216 2343
rect 1232 2335 1234 2353
rect 1292 2348 1294 2382
rect 1310 2358 1316 2359
rect 1310 2354 1311 2358
rect 1315 2354 1316 2358
rect 1310 2353 1316 2354
rect 1290 2347 1296 2348
rect 1290 2343 1291 2347
rect 1295 2343 1296 2347
rect 1290 2342 1296 2343
rect 1312 2335 1314 2353
rect 1372 2348 1374 2382
rect 1390 2358 1396 2359
rect 1390 2354 1391 2358
rect 1395 2354 1396 2358
rect 1390 2353 1396 2354
rect 1370 2347 1376 2348
rect 1370 2343 1371 2347
rect 1375 2343 1376 2347
rect 1370 2342 1376 2343
rect 1326 2339 1332 2340
rect 1326 2335 1327 2339
rect 1331 2335 1332 2339
rect 1392 2335 1394 2353
rect 1452 2348 1454 2382
rect 1470 2379 1471 2383
rect 1475 2379 1476 2383
rect 1470 2378 1476 2379
rect 1830 2376 1836 2377
rect 1830 2372 1831 2376
rect 1835 2372 1836 2376
rect 1872 2374 1874 2393
rect 2144 2377 2146 2393
rect 2240 2377 2242 2393
rect 2344 2377 2346 2393
rect 2456 2377 2458 2393
rect 2142 2376 2148 2377
rect 1830 2371 1836 2372
rect 1870 2373 1876 2374
rect 1470 2358 1476 2359
rect 1470 2354 1471 2358
rect 1475 2354 1476 2358
rect 1470 2353 1476 2354
rect 1450 2347 1456 2348
rect 1450 2343 1451 2347
rect 1455 2343 1456 2347
rect 1450 2342 1456 2343
rect 1472 2335 1474 2353
rect 1832 2335 1834 2371
rect 1870 2369 1871 2373
rect 1875 2369 1876 2373
rect 2142 2372 2143 2376
rect 2147 2372 2148 2376
rect 2142 2371 2148 2372
rect 2238 2376 2244 2377
rect 2238 2372 2239 2376
rect 2243 2372 2244 2376
rect 2238 2371 2244 2372
rect 2342 2376 2348 2377
rect 2342 2372 2343 2376
rect 2347 2372 2348 2376
rect 2342 2371 2348 2372
rect 2454 2376 2460 2377
rect 2454 2372 2455 2376
rect 2459 2372 2460 2376
rect 2454 2371 2460 2372
rect 1870 2368 1876 2369
rect 2214 2367 2220 2368
rect 2214 2363 2215 2367
rect 2219 2363 2220 2367
rect 2214 2362 2220 2363
rect 1870 2356 1876 2357
rect 1870 2352 1871 2356
rect 1875 2352 1876 2356
rect 1870 2351 1876 2352
rect 111 2334 115 2335
rect 111 2329 115 2330
rect 359 2334 363 2335
rect 359 2329 363 2330
rect 439 2334 443 2335
rect 439 2329 443 2330
rect 519 2334 523 2335
rect 519 2329 523 2330
rect 599 2334 603 2335
rect 599 2329 603 2330
rect 679 2334 683 2335
rect 679 2329 683 2330
rect 759 2334 763 2335
rect 759 2329 763 2330
rect 839 2334 843 2335
rect 839 2329 843 2330
rect 919 2334 923 2335
rect 926 2331 927 2335
rect 931 2331 932 2335
rect 926 2330 932 2331
rect 999 2334 1003 2335
rect 919 2329 923 2330
rect 112 2301 114 2329
rect 360 2319 362 2329
rect 440 2319 442 2329
rect 446 2327 452 2328
rect 446 2323 447 2327
rect 451 2323 452 2327
rect 446 2322 452 2323
rect 358 2318 364 2319
rect 358 2314 359 2318
rect 363 2314 364 2318
rect 358 2313 364 2314
rect 438 2318 444 2319
rect 438 2314 439 2318
rect 443 2314 444 2318
rect 438 2313 444 2314
rect 110 2300 116 2301
rect 110 2296 111 2300
rect 115 2296 116 2300
rect 110 2295 116 2296
rect 448 2292 450 2322
rect 520 2319 522 2329
rect 526 2327 532 2328
rect 526 2323 527 2327
rect 531 2323 532 2327
rect 526 2322 532 2323
rect 518 2318 524 2319
rect 518 2314 519 2318
rect 523 2314 524 2318
rect 518 2313 524 2314
rect 528 2292 530 2322
rect 600 2319 602 2329
rect 606 2327 612 2328
rect 606 2323 607 2327
rect 611 2323 612 2327
rect 606 2322 612 2323
rect 598 2318 604 2319
rect 598 2314 599 2318
rect 603 2314 604 2318
rect 598 2313 604 2314
rect 608 2292 610 2322
rect 680 2319 682 2329
rect 686 2327 692 2328
rect 686 2323 687 2327
rect 691 2323 692 2327
rect 686 2322 692 2323
rect 678 2318 684 2319
rect 678 2314 679 2318
rect 683 2314 684 2318
rect 678 2313 684 2314
rect 688 2292 690 2322
rect 760 2319 762 2329
rect 766 2327 772 2328
rect 766 2323 767 2327
rect 771 2323 772 2327
rect 766 2322 772 2323
rect 758 2318 764 2319
rect 758 2314 759 2318
rect 763 2314 764 2318
rect 758 2313 764 2314
rect 768 2292 770 2322
rect 840 2319 842 2329
rect 862 2327 868 2328
rect 862 2323 863 2327
rect 867 2323 868 2327
rect 862 2322 868 2323
rect 890 2327 896 2328
rect 890 2323 891 2327
rect 895 2323 896 2327
rect 890 2322 896 2323
rect 838 2318 844 2319
rect 838 2314 839 2318
rect 843 2314 844 2318
rect 838 2313 844 2314
rect 406 2291 412 2292
rect 406 2287 407 2291
rect 411 2287 412 2291
rect 406 2286 412 2287
rect 446 2291 452 2292
rect 446 2287 447 2291
rect 451 2287 452 2291
rect 446 2286 452 2287
rect 526 2291 532 2292
rect 526 2287 527 2291
rect 531 2287 532 2291
rect 526 2286 532 2287
rect 606 2291 612 2292
rect 606 2287 607 2291
rect 611 2287 612 2291
rect 606 2286 612 2287
rect 686 2291 692 2292
rect 686 2287 687 2291
rect 691 2287 692 2291
rect 686 2286 692 2287
rect 766 2291 772 2292
rect 766 2287 767 2291
rect 771 2287 772 2291
rect 766 2286 772 2287
rect 110 2283 116 2284
rect 110 2279 111 2283
rect 115 2279 116 2283
rect 110 2278 116 2279
rect 350 2280 356 2281
rect 112 2259 114 2278
rect 350 2276 351 2280
rect 355 2276 356 2280
rect 350 2275 356 2276
rect 352 2259 354 2275
rect 111 2258 115 2259
rect 111 2253 115 2254
rect 351 2258 355 2259
rect 351 2253 355 2254
rect 375 2258 379 2259
rect 375 2253 379 2254
rect 112 2234 114 2253
rect 376 2237 378 2253
rect 374 2236 380 2237
rect 110 2233 116 2234
rect 110 2229 111 2233
rect 115 2229 116 2233
rect 374 2232 375 2236
rect 379 2232 380 2236
rect 374 2231 380 2232
rect 110 2228 116 2229
rect 110 2216 116 2217
rect 110 2212 111 2216
rect 115 2212 116 2216
rect 110 2211 116 2212
rect 112 2171 114 2211
rect 382 2198 388 2199
rect 382 2194 383 2198
rect 387 2194 388 2198
rect 382 2193 388 2194
rect 384 2171 386 2193
rect 408 2188 410 2286
rect 430 2280 436 2281
rect 430 2276 431 2280
rect 435 2276 436 2280
rect 430 2275 436 2276
rect 510 2280 516 2281
rect 510 2276 511 2280
rect 515 2276 516 2280
rect 510 2275 516 2276
rect 590 2280 596 2281
rect 590 2276 591 2280
rect 595 2276 596 2280
rect 590 2275 596 2276
rect 670 2280 676 2281
rect 670 2276 671 2280
rect 675 2276 676 2280
rect 670 2275 676 2276
rect 750 2280 756 2281
rect 750 2276 751 2280
rect 755 2276 756 2280
rect 750 2275 756 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 432 2259 434 2275
rect 512 2259 514 2275
rect 592 2259 594 2275
rect 672 2259 674 2275
rect 752 2259 754 2275
rect 832 2259 834 2275
rect 431 2258 435 2259
rect 431 2253 435 2254
rect 455 2258 459 2259
rect 455 2253 459 2254
rect 511 2258 515 2259
rect 511 2253 515 2254
rect 535 2258 539 2259
rect 535 2253 539 2254
rect 591 2258 595 2259
rect 591 2253 595 2254
rect 615 2258 619 2259
rect 615 2253 619 2254
rect 671 2258 675 2259
rect 671 2253 675 2254
rect 695 2258 699 2259
rect 695 2253 699 2254
rect 751 2258 755 2259
rect 751 2253 755 2254
rect 775 2258 779 2259
rect 775 2253 779 2254
rect 831 2258 835 2259
rect 831 2253 835 2254
rect 855 2258 859 2259
rect 855 2253 859 2254
rect 456 2237 458 2253
rect 536 2237 538 2253
rect 616 2237 618 2253
rect 696 2237 698 2253
rect 776 2237 778 2253
rect 856 2237 858 2253
rect 454 2236 460 2237
rect 454 2232 455 2236
rect 459 2232 460 2236
rect 454 2231 460 2232
rect 534 2236 540 2237
rect 534 2232 535 2236
rect 539 2232 540 2236
rect 534 2231 540 2232
rect 614 2236 620 2237
rect 614 2232 615 2236
rect 619 2232 620 2236
rect 614 2231 620 2232
rect 694 2236 700 2237
rect 694 2232 695 2236
rect 699 2232 700 2236
rect 694 2231 700 2232
rect 774 2236 780 2237
rect 774 2232 775 2236
rect 779 2232 780 2236
rect 774 2231 780 2232
rect 854 2236 860 2237
rect 854 2232 855 2236
rect 859 2232 860 2236
rect 854 2231 860 2232
rect 442 2227 448 2228
rect 442 2223 443 2227
rect 447 2223 448 2227
rect 442 2222 448 2223
rect 526 2227 532 2228
rect 526 2223 527 2227
rect 531 2223 532 2227
rect 526 2222 532 2223
rect 682 2227 688 2228
rect 682 2223 683 2227
rect 687 2223 688 2227
rect 682 2222 688 2223
rect 762 2227 768 2228
rect 762 2223 763 2227
rect 767 2223 768 2227
rect 864 2224 866 2322
rect 892 2292 894 2322
rect 920 2319 922 2329
rect 918 2318 924 2319
rect 918 2314 919 2318
rect 923 2314 924 2318
rect 918 2313 924 2314
rect 928 2292 930 2330
rect 999 2329 1003 2330
rect 1071 2334 1075 2335
rect 1071 2329 1075 2330
rect 1079 2334 1083 2335
rect 1079 2329 1083 2330
rect 1151 2334 1155 2335
rect 1151 2329 1155 2330
rect 1159 2334 1163 2335
rect 1159 2329 1163 2330
rect 1231 2334 1235 2335
rect 1231 2329 1235 2330
rect 1239 2334 1243 2335
rect 1239 2329 1243 2330
rect 1311 2334 1315 2335
rect 1311 2329 1315 2330
rect 1319 2334 1323 2335
rect 1326 2334 1332 2335
rect 1391 2334 1395 2335
rect 1319 2329 1323 2330
rect 1000 2319 1002 2329
rect 1042 2327 1048 2328
rect 1042 2323 1043 2327
rect 1047 2323 1048 2327
rect 1042 2322 1048 2323
rect 1050 2327 1056 2328
rect 1050 2323 1051 2327
rect 1055 2323 1056 2327
rect 1050 2322 1056 2323
rect 998 2318 1004 2319
rect 998 2314 999 2318
rect 1003 2314 1004 2318
rect 998 2313 1004 2314
rect 890 2291 896 2292
rect 890 2287 891 2291
rect 895 2287 896 2291
rect 890 2286 896 2287
rect 926 2291 932 2292
rect 926 2287 927 2291
rect 931 2287 932 2291
rect 926 2286 932 2287
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 912 2259 914 2275
rect 992 2259 994 2275
rect 1044 2260 1046 2322
rect 1052 2292 1054 2322
rect 1080 2319 1082 2329
rect 1130 2327 1136 2328
rect 1130 2323 1131 2327
rect 1135 2323 1136 2327
rect 1130 2322 1136 2323
rect 1078 2318 1084 2319
rect 1078 2314 1079 2318
rect 1083 2314 1084 2318
rect 1078 2313 1084 2314
rect 1132 2292 1134 2322
rect 1160 2319 1162 2329
rect 1210 2327 1216 2328
rect 1210 2323 1211 2327
rect 1215 2323 1216 2327
rect 1210 2322 1216 2323
rect 1158 2318 1164 2319
rect 1158 2314 1159 2318
rect 1163 2314 1164 2318
rect 1158 2313 1164 2314
rect 1212 2292 1214 2322
rect 1240 2319 1242 2329
rect 1290 2327 1296 2328
rect 1290 2323 1291 2327
rect 1295 2323 1296 2327
rect 1290 2322 1296 2323
rect 1238 2318 1244 2319
rect 1238 2314 1239 2318
rect 1243 2314 1244 2318
rect 1238 2313 1244 2314
rect 1292 2292 1294 2322
rect 1320 2319 1322 2329
rect 1318 2318 1324 2319
rect 1318 2314 1319 2318
rect 1323 2314 1324 2318
rect 1318 2313 1324 2314
rect 1328 2292 1330 2334
rect 1391 2329 1395 2330
rect 1471 2334 1475 2335
rect 1471 2329 1475 2330
rect 1831 2334 1835 2335
rect 1831 2329 1835 2330
rect 1832 2301 1834 2329
rect 1872 2319 1874 2351
rect 2150 2338 2156 2339
rect 2150 2334 2151 2338
rect 2155 2334 2156 2338
rect 2150 2333 2156 2334
rect 2152 2319 2154 2333
rect 2179 2332 2183 2333
rect 2216 2328 2218 2362
rect 2306 2359 2312 2360
rect 2306 2355 2307 2359
rect 2311 2355 2312 2359
rect 2306 2354 2312 2355
rect 2246 2338 2252 2339
rect 2246 2334 2247 2338
rect 2251 2334 2252 2338
rect 2246 2333 2252 2334
rect 2178 2327 2184 2328
rect 2178 2323 2179 2327
rect 2183 2323 2184 2327
rect 2178 2322 2184 2323
rect 2214 2327 2220 2328
rect 2214 2323 2215 2327
rect 2219 2323 2220 2327
rect 2214 2322 2220 2323
rect 2248 2319 2250 2333
rect 1871 2318 1875 2319
rect 1871 2313 1875 2314
rect 2151 2318 2155 2319
rect 2151 2313 2155 2314
rect 2247 2318 2251 2319
rect 2247 2313 2251 2314
rect 2279 2318 2283 2319
rect 2279 2313 2283 2314
rect 1830 2300 1836 2301
rect 1830 2296 1831 2300
rect 1835 2296 1836 2300
rect 1830 2295 1836 2296
rect 1050 2291 1056 2292
rect 1050 2287 1051 2291
rect 1055 2287 1056 2291
rect 1050 2286 1056 2287
rect 1130 2291 1136 2292
rect 1130 2287 1131 2291
rect 1135 2287 1136 2291
rect 1130 2286 1136 2287
rect 1210 2291 1216 2292
rect 1210 2287 1211 2291
rect 1215 2287 1216 2291
rect 1210 2286 1216 2287
rect 1290 2291 1296 2292
rect 1290 2287 1291 2291
rect 1295 2287 1296 2291
rect 1290 2286 1296 2287
rect 1326 2291 1332 2292
rect 1326 2287 1327 2291
rect 1331 2287 1332 2291
rect 1326 2286 1332 2287
rect 1872 2285 1874 2313
rect 2280 2303 2282 2313
rect 2308 2312 2310 2354
rect 2350 2338 2356 2339
rect 2350 2334 2351 2338
rect 2355 2334 2356 2338
rect 2350 2333 2356 2334
rect 2462 2338 2468 2339
rect 2462 2334 2463 2338
rect 2467 2334 2468 2338
rect 2462 2333 2468 2334
rect 2480 2333 2482 2402
rect 2544 2399 2546 2419
rect 2696 2399 2698 2419
rect 2856 2399 2858 2419
rect 2543 2398 2547 2399
rect 2543 2393 2547 2394
rect 2575 2398 2579 2399
rect 2575 2393 2579 2394
rect 2695 2398 2699 2399
rect 2695 2393 2699 2394
rect 2703 2398 2707 2399
rect 2703 2393 2707 2394
rect 2847 2398 2851 2399
rect 2847 2393 2851 2394
rect 2855 2398 2859 2399
rect 2855 2393 2859 2394
rect 2576 2377 2578 2393
rect 2704 2377 2706 2393
rect 2848 2377 2850 2393
rect 2574 2376 2580 2377
rect 2574 2372 2575 2376
rect 2579 2372 2580 2376
rect 2574 2371 2580 2372
rect 2702 2376 2708 2377
rect 2702 2372 2703 2376
rect 2707 2372 2708 2376
rect 2702 2371 2708 2372
rect 2846 2376 2852 2377
rect 2846 2372 2847 2376
rect 2851 2372 2852 2376
rect 2846 2371 2852 2372
rect 2538 2367 2544 2368
rect 2538 2363 2539 2367
rect 2543 2363 2544 2367
rect 2538 2362 2544 2363
rect 2770 2367 2776 2368
rect 2770 2363 2771 2367
rect 2775 2363 2776 2367
rect 2770 2362 2776 2363
rect 2352 2319 2354 2333
rect 2464 2319 2466 2333
rect 2479 2332 2483 2333
rect 2540 2328 2542 2362
rect 2582 2338 2588 2339
rect 2582 2334 2583 2338
rect 2587 2334 2588 2338
rect 2582 2333 2588 2334
rect 2710 2338 2716 2339
rect 2710 2334 2711 2338
rect 2715 2334 2716 2338
rect 2710 2333 2716 2334
rect 2479 2327 2483 2328
rect 2538 2327 2544 2328
rect 2538 2323 2539 2327
rect 2543 2323 2544 2327
rect 2538 2322 2544 2323
rect 2584 2319 2586 2333
rect 2712 2319 2714 2333
rect 2772 2328 2774 2362
rect 2854 2338 2860 2339
rect 2854 2334 2855 2338
rect 2859 2334 2860 2338
rect 2854 2333 2860 2334
rect 2770 2327 2776 2328
rect 2770 2323 2771 2327
rect 2775 2323 2776 2327
rect 2770 2322 2776 2323
rect 2856 2319 2858 2333
rect 2883 2332 2887 2333
rect 2916 2328 2918 2430
rect 3014 2424 3020 2425
rect 3014 2420 3015 2424
rect 3019 2420 3020 2424
rect 3014 2419 3020 2420
rect 3182 2424 3188 2425
rect 3182 2420 3183 2424
rect 3187 2420 3188 2424
rect 3182 2419 3188 2420
rect 3350 2424 3356 2425
rect 3350 2420 3351 2424
rect 3355 2420 3356 2424
rect 3350 2419 3356 2420
rect 3016 2399 3018 2419
rect 3184 2399 3186 2419
rect 3352 2399 3354 2419
rect 3007 2398 3011 2399
rect 3007 2393 3011 2394
rect 3015 2398 3019 2399
rect 3015 2393 3019 2394
rect 3175 2398 3179 2399
rect 3175 2393 3179 2394
rect 3183 2398 3187 2399
rect 3183 2393 3187 2394
rect 3351 2398 3355 2399
rect 3351 2393 3355 2394
rect 3008 2377 3010 2393
rect 3176 2377 3178 2393
rect 3352 2377 3354 2393
rect 3006 2376 3012 2377
rect 3006 2372 3007 2376
rect 3011 2372 3012 2376
rect 3006 2371 3012 2372
rect 3174 2376 3180 2377
rect 3174 2372 3175 2376
rect 3179 2372 3180 2376
rect 3174 2371 3180 2372
rect 3350 2376 3356 2377
rect 3350 2372 3351 2376
rect 3355 2372 3356 2376
rect 3350 2371 3356 2372
rect 3420 2368 3422 2466
rect 3512 2463 3514 2473
rect 3564 2472 3566 2518
rect 3572 2492 3574 2686
rect 3590 2680 3596 2681
rect 3590 2676 3591 2680
rect 3595 2676 3596 2680
rect 3590 2675 3596 2676
rect 3592 2639 3594 2675
rect 3591 2638 3595 2639
rect 3591 2633 3595 2634
rect 3592 2605 3594 2633
rect 3590 2604 3596 2605
rect 3590 2600 3591 2604
rect 3595 2600 3596 2604
rect 3590 2599 3596 2600
rect 3590 2587 3596 2588
rect 3590 2583 3591 2587
rect 3595 2583 3596 2587
rect 3590 2582 3596 2583
rect 3592 2563 3594 2582
rect 3591 2562 3595 2563
rect 3591 2557 3595 2558
rect 3592 2538 3594 2557
rect 3590 2537 3596 2538
rect 3590 2533 3591 2537
rect 3595 2533 3596 2537
rect 3590 2532 3596 2533
rect 3590 2520 3596 2521
rect 3590 2516 3591 2520
rect 3595 2516 3596 2520
rect 3590 2515 3596 2516
rect 3570 2491 3576 2492
rect 3570 2487 3571 2491
rect 3575 2487 3576 2491
rect 3570 2486 3576 2487
rect 3592 2479 3594 2515
rect 3591 2478 3595 2479
rect 3591 2473 3595 2474
rect 3562 2471 3568 2472
rect 3562 2467 3563 2471
rect 3567 2467 3568 2471
rect 3562 2466 3568 2467
rect 3510 2462 3516 2463
rect 3510 2458 3511 2462
rect 3515 2458 3516 2462
rect 3510 2457 3516 2458
rect 3592 2445 3594 2473
rect 3590 2444 3596 2445
rect 3590 2440 3591 2444
rect 3595 2440 3596 2444
rect 3590 2439 3596 2440
rect 3534 2435 3540 2436
rect 3534 2431 3535 2435
rect 3539 2431 3540 2435
rect 3534 2430 3540 2431
rect 3502 2424 3508 2425
rect 3502 2420 3503 2424
rect 3507 2420 3508 2424
rect 3502 2419 3508 2420
rect 3504 2399 3506 2419
rect 3503 2398 3507 2399
rect 3503 2393 3507 2394
rect 3504 2377 3506 2393
rect 3502 2376 3508 2377
rect 3502 2372 3503 2376
rect 3507 2372 3508 2376
rect 3502 2371 3508 2372
rect 3114 2367 3120 2368
rect 3114 2363 3115 2367
rect 3119 2363 3120 2367
rect 3114 2362 3120 2363
rect 3122 2367 3128 2368
rect 3122 2363 3123 2367
rect 3127 2363 3128 2367
rect 3122 2362 3128 2363
rect 3418 2367 3424 2368
rect 3418 2363 3419 2367
rect 3423 2363 3424 2367
rect 3418 2362 3424 2363
rect 3014 2338 3020 2339
rect 3014 2334 3015 2338
rect 3019 2334 3020 2338
rect 3014 2333 3020 2334
rect 2882 2327 2888 2328
rect 2882 2323 2883 2327
rect 2887 2323 2888 2327
rect 2882 2322 2888 2323
rect 2914 2327 2920 2328
rect 2914 2323 2915 2327
rect 2919 2323 2920 2327
rect 2914 2322 2920 2323
rect 2942 2319 2948 2320
rect 3016 2319 3018 2333
rect 3116 2328 3118 2362
rect 3124 2333 3126 2362
rect 3182 2338 3188 2339
rect 3182 2334 3183 2338
rect 3187 2334 3188 2338
rect 3182 2333 3188 2334
rect 3358 2338 3364 2339
rect 3358 2334 3359 2338
rect 3363 2334 3364 2338
rect 3358 2333 3364 2334
rect 3510 2338 3516 2339
rect 3510 2334 3511 2338
rect 3515 2334 3516 2338
rect 3510 2333 3516 2334
rect 3123 2332 3127 2333
rect 3114 2327 3120 2328
rect 3123 2327 3127 2328
rect 3114 2323 3115 2327
rect 3119 2323 3120 2327
rect 3114 2322 3120 2323
rect 3184 2319 3186 2333
rect 3360 2319 3362 2333
rect 3418 2327 3424 2328
rect 3418 2323 3419 2327
rect 3423 2323 3424 2327
rect 3418 2322 3424 2323
rect 2351 2318 2355 2319
rect 2351 2313 2355 2314
rect 2359 2318 2363 2319
rect 2359 2313 2363 2314
rect 2439 2318 2443 2319
rect 2439 2313 2443 2314
rect 2463 2318 2467 2319
rect 2463 2313 2467 2314
rect 2519 2318 2523 2319
rect 2519 2313 2523 2314
rect 2583 2318 2587 2319
rect 2583 2313 2587 2314
rect 2599 2318 2603 2319
rect 2599 2313 2603 2314
rect 2679 2318 2683 2319
rect 2679 2313 2683 2314
rect 2711 2318 2715 2319
rect 2711 2313 2715 2314
rect 2759 2318 2763 2319
rect 2759 2313 2763 2314
rect 2847 2318 2851 2319
rect 2847 2313 2851 2314
rect 2855 2318 2859 2319
rect 2855 2313 2859 2314
rect 2935 2318 2939 2319
rect 2942 2315 2943 2319
rect 2947 2315 2948 2319
rect 2942 2314 2948 2315
rect 3015 2318 3019 2319
rect 2935 2313 2939 2314
rect 2306 2311 2312 2312
rect 2306 2307 2307 2311
rect 2311 2307 2312 2311
rect 2306 2306 2312 2307
rect 2330 2311 2336 2312
rect 2330 2307 2331 2311
rect 2335 2307 2336 2311
rect 2330 2306 2336 2307
rect 2278 2302 2284 2303
rect 2278 2298 2279 2302
rect 2283 2298 2284 2302
rect 2278 2297 2284 2298
rect 1870 2284 1876 2285
rect 1830 2283 1836 2284
rect 1070 2280 1076 2281
rect 1070 2276 1071 2280
rect 1075 2276 1076 2280
rect 1070 2275 1076 2276
rect 1150 2280 1156 2281
rect 1150 2276 1151 2280
rect 1155 2276 1156 2280
rect 1150 2275 1156 2276
rect 1230 2280 1236 2281
rect 1230 2276 1231 2280
rect 1235 2276 1236 2280
rect 1230 2275 1236 2276
rect 1310 2280 1316 2281
rect 1310 2276 1311 2280
rect 1315 2276 1316 2280
rect 1830 2279 1831 2283
rect 1835 2279 1836 2283
rect 1870 2280 1871 2284
rect 1875 2280 1876 2284
rect 1870 2279 1876 2280
rect 1830 2278 1836 2279
rect 1310 2275 1316 2276
rect 1042 2259 1048 2260
rect 1072 2259 1074 2275
rect 1152 2259 1154 2275
rect 1232 2259 1234 2275
rect 1242 2259 1248 2260
rect 1312 2259 1314 2275
rect 1832 2259 1834 2278
rect 2332 2276 2334 2306
rect 2360 2303 2362 2313
rect 2410 2311 2416 2312
rect 2410 2307 2411 2311
rect 2415 2307 2416 2311
rect 2410 2306 2416 2307
rect 2358 2302 2364 2303
rect 2358 2298 2359 2302
rect 2363 2298 2364 2302
rect 2358 2297 2364 2298
rect 2412 2276 2414 2306
rect 2440 2303 2442 2313
rect 2490 2311 2496 2312
rect 2490 2307 2491 2311
rect 2495 2307 2496 2311
rect 2490 2306 2496 2307
rect 2438 2302 2444 2303
rect 2438 2298 2439 2302
rect 2443 2298 2444 2302
rect 2438 2297 2444 2298
rect 2492 2276 2494 2306
rect 2520 2303 2522 2313
rect 2600 2303 2602 2313
rect 2680 2303 2682 2313
rect 2686 2311 2692 2312
rect 2686 2307 2687 2311
rect 2691 2307 2692 2311
rect 2686 2306 2692 2307
rect 2518 2302 2524 2303
rect 2518 2298 2519 2302
rect 2523 2298 2524 2302
rect 2518 2297 2524 2298
rect 2598 2302 2604 2303
rect 2598 2298 2599 2302
rect 2603 2298 2604 2302
rect 2598 2297 2604 2298
rect 2678 2302 2684 2303
rect 2678 2298 2679 2302
rect 2683 2298 2684 2302
rect 2678 2297 2684 2298
rect 2688 2276 2690 2306
rect 2760 2303 2762 2313
rect 2810 2311 2816 2312
rect 2810 2307 2811 2311
rect 2815 2307 2816 2311
rect 2810 2306 2816 2307
rect 2758 2302 2764 2303
rect 2758 2298 2759 2302
rect 2763 2298 2764 2302
rect 2758 2297 2764 2298
rect 2812 2276 2814 2306
rect 2848 2303 2850 2313
rect 2898 2311 2904 2312
rect 2898 2307 2899 2311
rect 2903 2307 2904 2311
rect 2898 2306 2904 2307
rect 2846 2302 2852 2303
rect 2846 2298 2847 2302
rect 2851 2298 2852 2302
rect 2846 2297 2852 2298
rect 2900 2276 2902 2306
rect 2936 2303 2938 2313
rect 2934 2302 2940 2303
rect 2934 2298 2935 2302
rect 2939 2298 2940 2302
rect 2934 2297 2940 2298
rect 2944 2276 2946 2314
rect 3015 2313 3019 2314
rect 3183 2318 3187 2319
rect 3183 2313 3187 2314
rect 3359 2318 3363 2319
rect 3359 2313 3363 2314
rect 2330 2275 2336 2276
rect 2330 2271 2331 2275
rect 2335 2271 2336 2275
rect 2330 2270 2336 2271
rect 2410 2275 2416 2276
rect 2410 2271 2411 2275
rect 2415 2271 2416 2275
rect 2410 2270 2416 2271
rect 2490 2275 2496 2276
rect 2490 2271 2491 2275
rect 2495 2271 2496 2275
rect 2490 2270 2496 2271
rect 2630 2275 2636 2276
rect 2630 2271 2631 2275
rect 2635 2271 2636 2275
rect 2630 2270 2636 2271
rect 2686 2275 2692 2276
rect 2686 2271 2687 2275
rect 2691 2271 2692 2275
rect 2686 2270 2692 2271
rect 2810 2275 2816 2276
rect 2810 2271 2811 2275
rect 2815 2271 2816 2275
rect 2810 2270 2816 2271
rect 2898 2275 2904 2276
rect 2898 2271 2899 2275
rect 2903 2271 2904 2275
rect 2898 2270 2904 2271
rect 2942 2275 2948 2276
rect 2942 2271 2943 2275
rect 2947 2271 2948 2275
rect 2942 2270 2948 2271
rect 1870 2267 1876 2268
rect 1870 2263 1871 2267
rect 1875 2263 1876 2267
rect 1870 2262 1876 2263
rect 2270 2264 2276 2265
rect 911 2258 915 2259
rect 911 2253 915 2254
rect 935 2258 939 2259
rect 935 2253 939 2254
rect 991 2258 995 2259
rect 991 2253 995 2254
rect 1015 2258 1019 2259
rect 1042 2255 1043 2259
rect 1047 2255 1048 2259
rect 1042 2254 1048 2255
rect 1071 2258 1075 2259
rect 1015 2253 1019 2254
rect 1071 2253 1075 2254
rect 1095 2258 1099 2259
rect 1095 2253 1099 2254
rect 1151 2258 1155 2259
rect 1151 2253 1155 2254
rect 1175 2258 1179 2259
rect 1175 2253 1179 2254
rect 1231 2258 1235 2259
rect 1242 2255 1243 2259
rect 1247 2255 1248 2259
rect 1242 2254 1248 2255
rect 1255 2258 1259 2259
rect 1231 2253 1235 2254
rect 936 2237 938 2253
rect 1016 2237 1018 2253
rect 1096 2237 1098 2253
rect 1176 2237 1178 2253
rect 934 2236 940 2237
rect 934 2232 935 2236
rect 939 2232 940 2236
rect 934 2231 940 2232
rect 1014 2236 1020 2237
rect 1014 2232 1015 2236
rect 1019 2232 1020 2236
rect 1014 2231 1020 2232
rect 1094 2236 1100 2237
rect 1094 2232 1095 2236
rect 1099 2232 1100 2236
rect 1094 2231 1100 2232
rect 1174 2236 1180 2237
rect 1174 2232 1175 2236
rect 1179 2232 1180 2236
rect 1174 2231 1180 2232
rect 1244 2228 1246 2254
rect 1255 2253 1259 2254
rect 1311 2258 1315 2259
rect 1311 2253 1315 2254
rect 1831 2258 1835 2259
rect 1831 2253 1835 2254
rect 1256 2237 1258 2253
rect 1254 2236 1260 2237
rect 1254 2232 1255 2236
rect 1259 2232 1260 2236
rect 1832 2234 1834 2253
rect 1872 2243 1874 2262
rect 2270 2260 2271 2264
rect 2275 2260 2276 2264
rect 2270 2259 2276 2260
rect 2350 2264 2356 2265
rect 2350 2260 2351 2264
rect 2355 2260 2356 2264
rect 2350 2259 2356 2260
rect 2430 2264 2436 2265
rect 2430 2260 2431 2264
rect 2435 2260 2436 2264
rect 2430 2259 2436 2260
rect 2510 2264 2516 2265
rect 2510 2260 2511 2264
rect 2515 2260 2516 2264
rect 2510 2259 2516 2260
rect 2590 2264 2596 2265
rect 2590 2260 2591 2264
rect 2595 2260 2596 2264
rect 2590 2259 2596 2260
rect 2272 2243 2274 2259
rect 2352 2243 2354 2259
rect 2358 2247 2364 2248
rect 2358 2243 2359 2247
rect 2363 2243 2364 2247
rect 2432 2243 2434 2259
rect 2512 2243 2514 2259
rect 2592 2243 2594 2259
rect 1871 2242 1875 2243
rect 1871 2237 1875 2238
rect 2271 2242 2275 2243
rect 2271 2237 2275 2238
rect 2311 2242 2315 2243
rect 2311 2237 2315 2238
rect 2351 2242 2355 2243
rect 2358 2242 2364 2243
rect 2399 2242 2403 2243
rect 2351 2237 2355 2238
rect 1254 2231 1260 2232
rect 1830 2233 1836 2234
rect 1830 2229 1831 2233
rect 1835 2229 1836 2233
rect 1830 2228 1836 2229
rect 922 2227 928 2228
rect 762 2222 768 2223
rect 862 2223 868 2224
rect 444 2188 446 2222
rect 514 2219 520 2220
rect 514 2215 515 2219
rect 519 2215 520 2219
rect 514 2214 520 2215
rect 462 2198 468 2199
rect 462 2194 463 2198
rect 467 2194 468 2198
rect 462 2193 468 2194
rect 406 2187 412 2188
rect 406 2183 407 2187
rect 411 2183 412 2187
rect 406 2182 412 2183
rect 442 2187 448 2188
rect 442 2183 443 2187
rect 447 2183 448 2187
rect 442 2182 448 2183
rect 464 2171 466 2193
rect 516 2188 518 2214
rect 514 2187 520 2188
rect 514 2183 515 2187
rect 519 2183 520 2187
rect 514 2182 520 2183
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 311 2170 315 2171
rect 311 2165 315 2166
rect 383 2170 387 2171
rect 383 2165 387 2166
rect 407 2170 411 2171
rect 407 2165 411 2166
rect 463 2170 467 2171
rect 463 2165 467 2166
rect 503 2170 507 2171
rect 503 2165 507 2166
rect 112 2137 114 2165
rect 312 2155 314 2165
rect 408 2155 410 2165
rect 414 2163 420 2164
rect 414 2159 415 2163
rect 419 2159 420 2163
rect 414 2158 420 2159
rect 310 2154 316 2155
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 406 2154 412 2155
rect 406 2150 407 2154
rect 411 2150 412 2154
rect 406 2149 412 2150
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 416 2128 418 2158
rect 504 2155 506 2165
rect 528 2164 530 2222
rect 542 2198 548 2199
rect 542 2194 543 2198
rect 547 2194 548 2198
rect 542 2193 548 2194
rect 622 2198 628 2199
rect 622 2194 623 2198
rect 627 2194 628 2198
rect 622 2193 628 2194
rect 544 2171 546 2193
rect 624 2171 626 2193
rect 684 2188 686 2222
rect 702 2198 708 2199
rect 702 2194 703 2198
rect 707 2194 708 2198
rect 702 2193 708 2194
rect 682 2187 688 2188
rect 682 2183 683 2187
rect 687 2183 688 2187
rect 682 2182 688 2183
rect 704 2171 706 2193
rect 764 2188 766 2222
rect 862 2219 863 2223
rect 867 2219 868 2223
rect 922 2223 923 2227
rect 927 2223 928 2227
rect 922 2222 928 2223
rect 1002 2227 1008 2228
rect 1002 2223 1003 2227
rect 1007 2223 1008 2227
rect 1002 2222 1008 2223
rect 1082 2227 1088 2228
rect 1082 2223 1083 2227
rect 1087 2223 1088 2227
rect 1082 2222 1088 2223
rect 1242 2227 1248 2228
rect 1242 2223 1243 2227
rect 1247 2223 1248 2227
rect 1242 2222 1248 2223
rect 862 2218 868 2219
rect 782 2198 788 2199
rect 782 2194 783 2198
rect 787 2194 788 2198
rect 782 2193 788 2194
rect 862 2198 868 2199
rect 862 2194 863 2198
rect 867 2194 868 2198
rect 862 2193 868 2194
rect 762 2187 768 2188
rect 762 2183 763 2187
rect 767 2183 768 2187
rect 762 2182 768 2183
rect 746 2179 752 2180
rect 746 2175 747 2179
rect 751 2175 752 2179
rect 746 2174 752 2175
rect 543 2170 547 2171
rect 543 2165 547 2166
rect 599 2170 603 2171
rect 599 2165 603 2166
rect 623 2170 627 2171
rect 623 2165 627 2166
rect 687 2170 691 2171
rect 687 2165 691 2166
rect 703 2170 707 2171
rect 703 2165 707 2166
rect 510 2163 516 2164
rect 510 2159 511 2163
rect 515 2159 516 2163
rect 510 2158 516 2159
rect 526 2163 532 2164
rect 526 2159 527 2163
rect 531 2159 532 2163
rect 526 2158 532 2159
rect 502 2154 508 2155
rect 502 2150 503 2154
rect 507 2150 508 2154
rect 502 2149 508 2150
rect 512 2128 514 2158
rect 600 2155 602 2165
rect 634 2163 640 2164
rect 634 2159 635 2163
rect 639 2159 640 2163
rect 634 2158 640 2159
rect 650 2163 656 2164
rect 650 2159 651 2163
rect 655 2159 656 2163
rect 650 2158 656 2159
rect 598 2154 604 2155
rect 598 2150 599 2154
rect 603 2150 604 2154
rect 598 2149 604 2150
rect 414 2127 420 2128
rect 414 2123 415 2127
rect 419 2123 420 2127
rect 414 2122 420 2123
rect 510 2127 516 2128
rect 510 2123 511 2127
rect 515 2123 516 2127
rect 510 2122 516 2123
rect 110 2119 116 2120
rect 110 2115 111 2119
rect 115 2115 116 2119
rect 110 2114 116 2115
rect 302 2116 308 2117
rect 112 2083 114 2114
rect 302 2112 303 2116
rect 307 2112 308 2116
rect 302 2111 308 2112
rect 398 2116 404 2117
rect 398 2112 399 2116
rect 403 2112 404 2116
rect 398 2111 404 2112
rect 494 2116 500 2117
rect 494 2112 495 2116
rect 499 2112 500 2116
rect 494 2111 500 2112
rect 590 2116 596 2117
rect 590 2112 591 2116
rect 595 2112 596 2116
rect 590 2111 596 2112
rect 242 2099 248 2100
rect 242 2095 243 2099
rect 247 2095 248 2099
rect 242 2094 248 2095
rect 111 2082 115 2083
rect 111 2077 115 2078
rect 207 2082 211 2083
rect 207 2077 211 2078
rect 112 2058 114 2077
rect 208 2061 210 2077
rect 206 2060 212 2061
rect 110 2057 116 2058
rect 110 2053 111 2057
rect 115 2053 116 2057
rect 206 2056 207 2060
rect 211 2056 212 2060
rect 206 2055 212 2056
rect 110 2052 116 2053
rect 110 2040 116 2041
rect 110 2036 111 2040
rect 115 2036 116 2040
rect 110 2035 116 2036
rect 112 2003 114 2035
rect 214 2022 220 2023
rect 214 2018 215 2022
rect 219 2018 220 2022
rect 214 2017 220 2018
rect 216 2003 218 2017
rect 244 2012 246 2094
rect 304 2083 306 2111
rect 400 2083 402 2111
rect 496 2083 498 2111
rect 592 2083 594 2111
rect 303 2082 307 2083
rect 303 2077 307 2078
rect 327 2082 331 2083
rect 327 2077 331 2078
rect 399 2082 403 2083
rect 399 2077 403 2078
rect 447 2082 451 2083
rect 447 2077 451 2078
rect 495 2082 499 2083
rect 495 2077 499 2078
rect 575 2082 579 2083
rect 575 2077 579 2078
rect 591 2082 595 2083
rect 591 2077 595 2078
rect 328 2061 330 2077
rect 448 2061 450 2077
rect 576 2061 578 2077
rect 326 2060 332 2061
rect 326 2056 327 2060
rect 331 2056 332 2060
rect 326 2055 332 2056
rect 446 2060 452 2061
rect 446 2056 447 2060
rect 451 2056 452 2060
rect 446 2055 452 2056
rect 574 2060 580 2061
rect 574 2056 575 2060
rect 579 2056 580 2060
rect 574 2055 580 2056
rect 274 2051 280 2052
rect 274 2047 275 2051
rect 279 2047 280 2051
rect 274 2046 280 2047
rect 394 2051 400 2052
rect 394 2047 395 2051
rect 399 2047 400 2051
rect 394 2046 400 2047
rect 276 2012 278 2046
rect 386 2043 392 2044
rect 386 2039 387 2043
rect 391 2039 392 2043
rect 386 2038 392 2039
rect 334 2022 340 2023
rect 334 2018 335 2022
rect 339 2018 340 2022
rect 334 2017 340 2018
rect 242 2011 248 2012
rect 242 2007 243 2011
rect 247 2007 248 2011
rect 242 2006 248 2007
rect 274 2011 280 2012
rect 274 2007 275 2011
rect 279 2007 280 2011
rect 274 2006 280 2007
rect 336 2003 338 2017
rect 388 2012 390 2038
rect 386 2011 392 2012
rect 386 2007 387 2011
rect 391 2007 392 2011
rect 386 2006 392 2007
rect 111 2002 115 2003
rect 111 1997 115 1998
rect 191 2002 195 2003
rect 191 1997 195 1998
rect 215 2002 219 2003
rect 215 1997 219 1998
rect 335 2002 339 2003
rect 335 1997 339 1998
rect 351 2002 355 2003
rect 351 1997 355 1998
rect 112 1969 114 1997
rect 192 1987 194 1997
rect 352 1987 354 1997
rect 396 1996 398 2046
rect 636 2044 638 2158
rect 652 2128 654 2158
rect 688 2155 690 2165
rect 738 2163 744 2164
rect 738 2159 739 2163
rect 743 2159 744 2163
rect 738 2158 744 2159
rect 686 2154 692 2155
rect 686 2150 687 2154
rect 691 2150 692 2154
rect 686 2149 692 2150
rect 740 2128 742 2158
rect 748 2128 750 2174
rect 784 2171 786 2193
rect 864 2171 866 2193
rect 924 2188 926 2222
rect 942 2198 948 2199
rect 942 2194 943 2198
rect 947 2194 948 2198
rect 942 2193 948 2194
rect 886 2187 892 2188
rect 886 2183 887 2187
rect 891 2183 892 2187
rect 886 2182 892 2183
rect 922 2187 928 2188
rect 922 2183 923 2187
rect 927 2183 928 2187
rect 922 2182 928 2183
rect 775 2170 779 2171
rect 775 2165 779 2166
rect 783 2170 787 2171
rect 783 2165 787 2166
rect 863 2170 867 2171
rect 863 2165 867 2166
rect 776 2155 778 2165
rect 864 2155 866 2165
rect 774 2154 780 2155
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 862 2154 868 2155
rect 862 2150 863 2154
rect 867 2150 868 2154
rect 862 2149 868 2150
rect 888 2128 890 2182
rect 944 2171 946 2193
rect 1004 2188 1006 2222
rect 1022 2198 1028 2199
rect 1022 2194 1023 2198
rect 1027 2194 1028 2198
rect 1022 2193 1028 2194
rect 1002 2187 1008 2188
rect 1002 2183 1003 2187
rect 1007 2183 1008 2187
rect 1002 2182 1008 2183
rect 1024 2171 1026 2193
rect 1084 2188 1086 2222
rect 1234 2219 1240 2220
rect 1234 2215 1235 2219
rect 1239 2215 1240 2219
rect 1872 2218 1874 2237
rect 2312 2221 2314 2237
rect 2310 2220 2316 2221
rect 1870 2217 1876 2218
rect 1234 2214 1240 2215
rect 1830 2216 1836 2217
rect 1102 2198 1108 2199
rect 1102 2194 1103 2198
rect 1107 2194 1108 2198
rect 1102 2193 1108 2194
rect 1182 2198 1188 2199
rect 1182 2194 1183 2198
rect 1187 2194 1188 2198
rect 1182 2193 1188 2194
rect 1082 2187 1088 2188
rect 1082 2183 1083 2187
rect 1087 2183 1088 2187
rect 1082 2182 1088 2183
rect 1104 2171 1106 2193
rect 1184 2171 1186 2193
rect 1236 2188 1238 2214
rect 1830 2212 1831 2216
rect 1835 2212 1836 2216
rect 1870 2213 1871 2217
rect 1875 2213 1876 2217
rect 2310 2216 2311 2220
rect 2315 2216 2316 2220
rect 2310 2215 2316 2216
rect 1870 2212 1876 2213
rect 1830 2211 1836 2212
rect 1262 2198 1268 2199
rect 1262 2194 1263 2198
rect 1267 2194 1268 2198
rect 1262 2193 1268 2194
rect 1234 2187 1240 2188
rect 1234 2183 1235 2187
rect 1239 2183 1240 2187
rect 1234 2182 1240 2183
rect 1264 2171 1266 2193
rect 1832 2171 1834 2211
rect 1870 2200 1876 2201
rect 1870 2196 1871 2200
rect 1875 2196 1876 2200
rect 1870 2195 1876 2196
rect 943 2170 947 2171
rect 943 2165 947 2166
rect 951 2170 955 2171
rect 951 2165 955 2166
rect 1023 2170 1027 2171
rect 1023 2165 1027 2166
rect 1039 2170 1043 2171
rect 1039 2165 1043 2166
rect 1103 2170 1107 2171
rect 1103 2165 1107 2166
rect 1127 2170 1131 2171
rect 1127 2165 1131 2166
rect 1183 2170 1187 2171
rect 1183 2165 1187 2166
rect 1223 2170 1227 2171
rect 1223 2165 1227 2166
rect 1263 2170 1267 2171
rect 1263 2165 1267 2166
rect 1831 2170 1835 2171
rect 1831 2165 1835 2166
rect 952 2155 954 2165
rect 958 2163 964 2164
rect 958 2159 959 2163
rect 963 2159 964 2163
rect 958 2158 964 2159
rect 950 2154 956 2155
rect 950 2150 951 2154
rect 955 2150 956 2154
rect 950 2149 956 2150
rect 960 2128 962 2158
rect 1040 2155 1042 2165
rect 1046 2163 1052 2164
rect 1046 2159 1047 2163
rect 1051 2159 1052 2163
rect 1046 2158 1052 2159
rect 1038 2154 1044 2155
rect 1038 2150 1039 2154
rect 1043 2150 1044 2154
rect 1038 2149 1044 2150
rect 1048 2128 1050 2158
rect 1128 2155 1130 2165
rect 1134 2163 1140 2164
rect 1134 2159 1135 2163
rect 1139 2159 1140 2163
rect 1134 2158 1140 2159
rect 1126 2154 1132 2155
rect 1126 2150 1127 2154
rect 1131 2150 1132 2154
rect 1126 2149 1132 2150
rect 1136 2128 1138 2158
rect 1224 2155 1226 2165
rect 1230 2163 1236 2164
rect 1230 2159 1231 2163
rect 1235 2159 1236 2163
rect 1230 2158 1236 2159
rect 1242 2163 1248 2164
rect 1242 2159 1243 2163
rect 1247 2159 1248 2163
rect 1242 2158 1248 2159
rect 1222 2154 1228 2155
rect 1222 2150 1223 2154
rect 1227 2150 1228 2154
rect 1222 2149 1228 2150
rect 1232 2128 1234 2158
rect 650 2127 656 2128
rect 650 2123 651 2127
rect 655 2123 656 2127
rect 650 2122 656 2123
rect 738 2127 744 2128
rect 738 2123 739 2127
rect 743 2123 744 2127
rect 738 2122 744 2123
rect 746 2127 752 2128
rect 746 2123 747 2127
rect 751 2123 752 2127
rect 746 2122 752 2123
rect 886 2127 892 2128
rect 886 2123 887 2127
rect 891 2123 892 2127
rect 886 2122 892 2123
rect 958 2127 964 2128
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 958 2122 964 2123
rect 1046 2127 1052 2128
rect 1046 2123 1047 2127
rect 1051 2123 1052 2127
rect 1046 2122 1052 2123
rect 1134 2127 1140 2128
rect 1134 2123 1135 2127
rect 1139 2123 1140 2127
rect 1134 2122 1140 2123
rect 1230 2127 1236 2128
rect 1230 2123 1231 2127
rect 1235 2123 1236 2127
rect 1230 2122 1236 2123
rect 678 2116 684 2117
rect 678 2112 679 2116
rect 683 2112 684 2116
rect 678 2111 684 2112
rect 766 2116 772 2117
rect 766 2112 767 2116
rect 771 2112 772 2116
rect 766 2111 772 2112
rect 854 2116 860 2117
rect 854 2112 855 2116
rect 859 2112 860 2116
rect 854 2111 860 2112
rect 942 2116 948 2117
rect 942 2112 943 2116
rect 947 2112 948 2116
rect 942 2111 948 2112
rect 1030 2116 1036 2117
rect 1030 2112 1031 2116
rect 1035 2112 1036 2116
rect 1030 2111 1036 2112
rect 1118 2116 1124 2117
rect 1118 2112 1119 2116
rect 1123 2112 1124 2116
rect 1118 2111 1124 2112
rect 1214 2116 1220 2117
rect 1214 2112 1215 2116
rect 1219 2112 1220 2116
rect 1214 2111 1220 2112
rect 680 2083 682 2111
rect 768 2083 770 2111
rect 856 2083 858 2111
rect 944 2083 946 2111
rect 1032 2083 1034 2111
rect 1120 2083 1122 2111
rect 1216 2083 1218 2111
rect 679 2082 683 2083
rect 679 2077 683 2078
rect 703 2082 707 2083
rect 703 2077 707 2078
rect 767 2082 771 2083
rect 767 2077 771 2078
rect 823 2082 827 2083
rect 823 2077 827 2078
rect 855 2082 859 2083
rect 855 2077 859 2078
rect 943 2082 947 2083
rect 943 2077 947 2078
rect 1031 2082 1035 2083
rect 1031 2077 1035 2078
rect 1063 2082 1067 2083
rect 1063 2077 1067 2078
rect 1119 2082 1123 2083
rect 1119 2077 1123 2078
rect 1175 2082 1179 2083
rect 1175 2077 1179 2078
rect 1215 2082 1219 2083
rect 1215 2077 1219 2078
rect 704 2061 706 2077
rect 824 2061 826 2077
rect 944 2061 946 2077
rect 1064 2061 1066 2077
rect 1176 2061 1178 2077
rect 702 2060 708 2061
rect 702 2056 703 2060
rect 707 2056 708 2060
rect 702 2055 708 2056
rect 822 2060 828 2061
rect 822 2056 823 2060
rect 827 2056 828 2060
rect 822 2055 828 2056
rect 942 2060 948 2061
rect 942 2056 943 2060
rect 947 2056 948 2060
rect 942 2055 948 2056
rect 1062 2060 1068 2061
rect 1062 2056 1063 2060
rect 1067 2056 1068 2060
rect 1062 2055 1068 2056
rect 1174 2060 1180 2061
rect 1174 2056 1175 2060
rect 1179 2056 1180 2060
rect 1174 2055 1180 2056
rect 1244 2052 1246 2158
rect 1832 2137 1834 2165
rect 1872 2163 1874 2195
rect 2318 2182 2324 2183
rect 2318 2178 2319 2182
rect 2323 2178 2324 2182
rect 2318 2177 2324 2178
rect 2320 2163 2322 2177
rect 2360 2172 2362 2242
rect 2399 2237 2403 2238
rect 2431 2242 2435 2243
rect 2431 2237 2435 2238
rect 2495 2242 2499 2243
rect 2495 2237 2499 2238
rect 2511 2242 2515 2243
rect 2511 2237 2515 2238
rect 2591 2242 2595 2243
rect 2591 2237 2595 2238
rect 2599 2242 2603 2243
rect 2599 2237 2603 2238
rect 2400 2221 2402 2237
rect 2496 2221 2498 2237
rect 2600 2221 2602 2237
rect 2398 2220 2404 2221
rect 2398 2216 2399 2220
rect 2403 2216 2404 2220
rect 2398 2215 2404 2216
rect 2494 2220 2500 2221
rect 2494 2216 2495 2220
rect 2499 2216 2500 2220
rect 2494 2215 2500 2216
rect 2598 2220 2604 2221
rect 2598 2216 2599 2220
rect 2603 2216 2604 2220
rect 2598 2215 2604 2216
rect 2378 2211 2384 2212
rect 2378 2207 2379 2211
rect 2383 2207 2384 2211
rect 2378 2206 2384 2207
rect 2470 2211 2476 2212
rect 2470 2207 2471 2211
rect 2475 2207 2476 2211
rect 2470 2206 2476 2207
rect 2562 2211 2568 2212
rect 2562 2207 2563 2211
rect 2567 2207 2568 2211
rect 2562 2206 2568 2207
rect 2380 2172 2382 2206
rect 2406 2182 2412 2183
rect 2406 2178 2407 2182
rect 2411 2178 2412 2182
rect 2406 2177 2412 2178
rect 2358 2171 2364 2172
rect 2358 2167 2359 2171
rect 2363 2167 2364 2171
rect 2358 2166 2364 2167
rect 2378 2171 2384 2172
rect 2378 2167 2379 2171
rect 2383 2167 2384 2171
rect 2378 2166 2384 2167
rect 2398 2163 2404 2164
rect 2408 2163 2410 2177
rect 2472 2172 2474 2206
rect 2502 2182 2508 2183
rect 2502 2178 2503 2182
rect 2507 2178 2508 2182
rect 2502 2177 2508 2178
rect 2470 2171 2476 2172
rect 2470 2167 2471 2171
rect 2475 2167 2476 2171
rect 2470 2166 2476 2167
rect 2504 2163 2506 2177
rect 1871 2162 1875 2163
rect 1871 2157 1875 2158
rect 1903 2162 1907 2163
rect 1903 2157 1907 2158
rect 1983 2162 1987 2163
rect 1983 2157 1987 2158
rect 2111 2162 2115 2163
rect 2111 2157 2115 2158
rect 2247 2162 2251 2163
rect 2247 2157 2251 2158
rect 2319 2162 2323 2163
rect 2319 2157 2323 2158
rect 2391 2162 2395 2163
rect 2398 2159 2399 2163
rect 2403 2159 2404 2163
rect 2398 2158 2404 2159
rect 2407 2162 2411 2163
rect 2391 2157 2395 2158
rect 1830 2136 1836 2137
rect 1830 2132 1831 2136
rect 1835 2132 1836 2136
rect 1830 2131 1836 2132
rect 1872 2129 1874 2157
rect 1904 2147 1906 2157
rect 1984 2147 1986 2157
rect 1990 2155 1996 2156
rect 1990 2151 1991 2155
rect 1995 2151 1996 2155
rect 1990 2150 1996 2151
rect 2050 2155 2056 2156
rect 2050 2151 2051 2155
rect 2055 2151 2056 2155
rect 2050 2150 2056 2151
rect 1902 2146 1908 2147
rect 1902 2142 1903 2146
rect 1907 2142 1908 2146
rect 1902 2141 1908 2142
rect 1982 2146 1988 2147
rect 1982 2142 1983 2146
rect 1987 2142 1988 2146
rect 1982 2141 1988 2142
rect 1870 2128 1876 2129
rect 1870 2124 1871 2128
rect 1875 2124 1876 2128
rect 1870 2123 1876 2124
rect 1992 2120 1994 2150
rect 1830 2119 1836 2120
rect 1830 2115 1831 2119
rect 1835 2115 1836 2119
rect 1830 2114 1836 2115
rect 1990 2119 1996 2120
rect 1990 2115 1991 2119
rect 1995 2115 1996 2119
rect 1990 2114 1996 2115
rect 1778 2091 1784 2092
rect 1778 2087 1779 2091
rect 1783 2087 1784 2091
rect 1778 2086 1784 2087
rect 1279 2082 1283 2083
rect 1279 2077 1283 2078
rect 1375 2082 1379 2083
rect 1375 2077 1379 2078
rect 1471 2082 1475 2083
rect 1471 2077 1475 2078
rect 1567 2082 1571 2083
rect 1567 2077 1571 2078
rect 1663 2082 1667 2083
rect 1663 2077 1667 2078
rect 1743 2082 1747 2083
rect 1743 2077 1747 2078
rect 1280 2061 1282 2077
rect 1376 2061 1378 2077
rect 1472 2061 1474 2077
rect 1568 2061 1570 2077
rect 1664 2061 1666 2077
rect 1744 2061 1746 2077
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 1374 2060 1380 2061
rect 1374 2056 1375 2060
rect 1379 2056 1380 2060
rect 1374 2055 1380 2056
rect 1470 2060 1476 2061
rect 1470 2056 1471 2060
rect 1475 2056 1476 2060
rect 1470 2055 1476 2056
rect 1566 2060 1572 2061
rect 1566 2056 1567 2060
rect 1571 2056 1572 2060
rect 1566 2055 1572 2056
rect 1662 2060 1668 2061
rect 1662 2056 1663 2060
rect 1667 2056 1668 2060
rect 1662 2055 1668 2056
rect 1742 2060 1748 2061
rect 1742 2056 1743 2060
rect 1747 2056 1748 2060
rect 1742 2055 1748 2056
rect 642 2051 648 2052
rect 642 2047 643 2051
rect 647 2047 648 2051
rect 642 2046 648 2047
rect 770 2051 776 2052
rect 770 2047 771 2051
rect 775 2047 776 2051
rect 770 2046 776 2047
rect 1030 2051 1036 2052
rect 1030 2047 1031 2051
rect 1035 2047 1036 2051
rect 1030 2046 1036 2047
rect 1130 2051 1136 2052
rect 1130 2047 1131 2051
rect 1135 2047 1136 2051
rect 1130 2046 1136 2047
rect 1242 2051 1248 2052
rect 1242 2047 1243 2051
rect 1247 2047 1248 2051
rect 1242 2046 1248 2047
rect 1346 2051 1352 2052
rect 1346 2047 1347 2051
rect 1351 2047 1352 2051
rect 1346 2046 1352 2047
rect 1442 2051 1448 2052
rect 1442 2047 1443 2051
rect 1447 2047 1448 2051
rect 1442 2046 1448 2047
rect 1538 2051 1544 2052
rect 1538 2047 1539 2051
rect 1543 2047 1544 2051
rect 1538 2046 1544 2047
rect 1634 2051 1640 2052
rect 1634 2047 1635 2051
rect 1639 2047 1640 2051
rect 1634 2046 1640 2047
rect 1730 2051 1736 2052
rect 1730 2047 1731 2051
rect 1735 2047 1736 2051
rect 1730 2046 1736 2047
rect 634 2043 640 2044
rect 634 2039 635 2043
rect 639 2039 640 2043
rect 634 2038 640 2039
rect 454 2022 460 2023
rect 454 2018 455 2022
rect 459 2018 460 2022
rect 454 2017 460 2018
rect 582 2022 588 2023
rect 582 2018 583 2022
rect 587 2018 588 2022
rect 582 2017 588 2018
rect 456 2003 458 2017
rect 584 2003 586 2017
rect 644 2012 646 2046
rect 710 2022 716 2023
rect 710 2018 711 2022
rect 715 2018 716 2022
rect 710 2017 716 2018
rect 642 2011 648 2012
rect 642 2007 643 2011
rect 647 2007 648 2011
rect 642 2006 648 2007
rect 712 2003 714 2017
rect 772 2012 774 2046
rect 830 2022 836 2023
rect 830 2018 831 2022
rect 835 2018 836 2022
rect 830 2017 836 2018
rect 950 2022 956 2023
rect 950 2018 951 2022
rect 955 2018 956 2022
rect 950 2017 956 2018
rect 770 2011 776 2012
rect 770 2007 771 2011
rect 775 2007 776 2011
rect 770 2006 776 2007
rect 832 2003 834 2017
rect 854 2011 860 2012
rect 854 2007 855 2011
rect 859 2009 866 2011
rect 859 2007 860 2009
rect 854 2006 860 2007
rect 455 2002 459 2003
rect 455 1997 459 1998
rect 519 2002 523 2003
rect 519 1997 523 1998
rect 583 2002 587 2003
rect 583 1997 587 1998
rect 687 2002 691 2003
rect 687 1997 691 1998
rect 711 2002 715 2003
rect 711 1997 715 1998
rect 831 2002 835 2003
rect 831 1997 835 1998
rect 855 2002 859 2003
rect 855 1997 859 1998
rect 358 1995 364 1996
rect 358 1991 359 1995
rect 363 1991 364 1995
rect 358 1990 364 1991
rect 394 1995 400 1996
rect 394 1991 395 1995
rect 399 1991 400 1995
rect 394 1990 400 1991
rect 190 1986 196 1987
rect 190 1982 191 1986
rect 195 1982 196 1986
rect 190 1981 196 1982
rect 350 1986 356 1987
rect 350 1982 351 1986
rect 355 1982 356 1986
rect 350 1981 356 1982
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 360 1960 362 1990
rect 520 1987 522 1997
rect 534 1995 540 1996
rect 534 1991 535 1995
rect 539 1991 540 1995
rect 534 1990 540 1991
rect 570 1995 576 1996
rect 570 1991 571 1995
rect 575 1991 576 1995
rect 570 1990 576 1991
rect 518 1986 524 1987
rect 518 1982 519 1986
rect 523 1982 524 1986
rect 518 1981 524 1982
rect 358 1959 364 1960
rect 358 1955 359 1959
rect 363 1955 364 1959
rect 358 1954 364 1955
rect 110 1951 116 1952
rect 110 1947 111 1951
rect 115 1947 116 1951
rect 110 1946 116 1947
rect 182 1948 188 1949
rect 112 1923 114 1946
rect 182 1944 183 1948
rect 187 1944 188 1948
rect 182 1943 188 1944
rect 342 1948 348 1949
rect 342 1944 343 1948
rect 347 1944 348 1948
rect 342 1943 348 1944
rect 510 1948 516 1949
rect 510 1944 511 1948
rect 515 1944 516 1948
rect 510 1943 516 1944
rect 184 1923 186 1943
rect 198 1931 204 1932
rect 198 1927 199 1931
rect 203 1927 204 1931
rect 198 1926 204 1927
rect 111 1922 115 1923
rect 111 1917 115 1918
rect 135 1922 139 1923
rect 135 1917 139 1918
rect 183 1922 187 1923
rect 183 1917 187 1918
rect 112 1898 114 1917
rect 136 1901 138 1917
rect 134 1900 140 1901
rect 110 1897 116 1898
rect 110 1893 111 1897
rect 115 1893 116 1897
rect 134 1896 135 1900
rect 139 1896 140 1900
rect 134 1895 140 1896
rect 110 1892 116 1893
rect 110 1880 116 1881
rect 110 1876 111 1880
rect 115 1876 116 1880
rect 110 1875 116 1876
rect 112 1843 114 1875
rect 142 1862 148 1863
rect 142 1858 143 1862
rect 147 1858 148 1862
rect 142 1857 148 1858
rect 144 1843 146 1857
rect 200 1852 202 1926
rect 344 1923 346 1943
rect 512 1923 514 1943
rect 239 1922 243 1923
rect 239 1917 243 1918
rect 343 1922 347 1923
rect 343 1917 347 1918
rect 375 1922 379 1923
rect 375 1917 379 1918
rect 511 1922 515 1923
rect 511 1917 515 1918
rect 527 1922 531 1923
rect 527 1917 531 1918
rect 240 1901 242 1917
rect 376 1901 378 1917
rect 528 1901 530 1917
rect 238 1900 244 1901
rect 238 1896 239 1900
rect 243 1896 244 1900
rect 238 1895 244 1896
rect 374 1900 380 1901
rect 374 1896 375 1900
rect 379 1896 380 1900
rect 374 1895 380 1896
rect 526 1900 532 1901
rect 526 1896 527 1900
rect 531 1896 532 1900
rect 526 1895 532 1896
rect 210 1891 216 1892
rect 210 1887 211 1891
rect 215 1887 216 1891
rect 210 1886 216 1887
rect 306 1891 312 1892
rect 306 1887 307 1891
rect 311 1887 312 1891
rect 306 1886 312 1887
rect 354 1891 360 1892
rect 354 1887 355 1891
rect 359 1887 360 1891
rect 536 1888 538 1990
rect 572 1960 574 1990
rect 688 1987 690 1997
rect 738 1995 744 1996
rect 738 1991 739 1995
rect 743 1991 744 1995
rect 738 1990 744 1991
rect 686 1986 692 1987
rect 686 1982 687 1986
rect 691 1982 692 1986
rect 686 1981 692 1982
rect 740 1960 742 1990
rect 856 1987 858 1997
rect 854 1986 860 1987
rect 854 1982 855 1986
rect 859 1982 860 1986
rect 854 1981 860 1982
rect 864 1960 866 2009
rect 952 2003 954 2017
rect 1032 2012 1034 2046
rect 1070 2022 1076 2023
rect 1070 2018 1071 2022
rect 1075 2018 1076 2022
rect 1070 2017 1076 2018
rect 1022 2011 1028 2012
rect 1022 2007 1023 2011
rect 1027 2007 1028 2011
rect 1022 2006 1028 2007
rect 1030 2011 1036 2012
rect 1030 2007 1031 2011
rect 1035 2007 1036 2011
rect 1030 2006 1036 2007
rect 951 2002 955 2003
rect 951 1997 955 1998
rect 1015 2002 1019 2003
rect 1015 1997 1019 1998
rect 1016 1987 1018 1997
rect 1014 1986 1020 1987
rect 1014 1982 1015 1986
rect 1019 1982 1020 1986
rect 1014 1981 1020 1982
rect 1024 1960 1026 2006
rect 1072 2003 1074 2017
rect 1132 2012 1134 2046
rect 1338 2043 1344 2044
rect 1338 2039 1339 2043
rect 1343 2039 1344 2043
rect 1338 2038 1344 2039
rect 1182 2022 1188 2023
rect 1182 2018 1183 2022
rect 1187 2018 1188 2022
rect 1182 2017 1188 2018
rect 1286 2022 1292 2023
rect 1286 2018 1287 2022
rect 1291 2018 1292 2022
rect 1286 2017 1292 2018
rect 1130 2011 1136 2012
rect 1130 2007 1131 2011
rect 1135 2007 1136 2011
rect 1130 2006 1136 2007
rect 1184 2003 1186 2017
rect 1288 2003 1290 2017
rect 1071 2002 1075 2003
rect 1071 1997 1075 1998
rect 1167 2002 1171 2003
rect 1167 1997 1171 1998
rect 1183 2002 1187 2003
rect 1183 1997 1187 1998
rect 1287 2002 1291 2003
rect 1287 1997 1291 1998
rect 1311 2002 1315 2003
rect 1311 1997 1315 1998
rect 1168 1987 1170 1997
rect 1174 1995 1180 1996
rect 1174 1991 1175 1995
rect 1179 1991 1180 1995
rect 1174 1990 1180 1991
rect 1218 1995 1224 1996
rect 1218 1991 1219 1995
rect 1223 1991 1224 1995
rect 1218 1990 1224 1991
rect 1166 1986 1172 1987
rect 1166 1982 1167 1986
rect 1171 1982 1172 1986
rect 1166 1981 1172 1982
rect 1176 1960 1178 1990
rect 570 1959 576 1960
rect 570 1955 571 1959
rect 575 1955 576 1959
rect 570 1954 576 1955
rect 738 1959 744 1960
rect 738 1955 739 1959
rect 743 1955 744 1959
rect 738 1954 744 1955
rect 862 1959 868 1960
rect 862 1955 863 1959
rect 867 1955 868 1959
rect 862 1954 868 1955
rect 1022 1959 1028 1960
rect 1022 1955 1023 1959
rect 1027 1955 1028 1959
rect 1022 1954 1028 1955
rect 1174 1959 1180 1960
rect 1174 1955 1175 1959
rect 1179 1955 1180 1959
rect 1174 1954 1180 1955
rect 678 1948 684 1949
rect 678 1944 679 1948
rect 683 1944 684 1948
rect 678 1943 684 1944
rect 846 1948 852 1949
rect 846 1944 847 1948
rect 851 1944 852 1948
rect 846 1943 852 1944
rect 1006 1948 1012 1949
rect 1006 1944 1007 1948
rect 1011 1944 1012 1948
rect 1006 1943 1012 1944
rect 1158 1948 1164 1949
rect 1158 1944 1159 1948
rect 1163 1944 1164 1948
rect 1158 1943 1164 1944
rect 680 1923 682 1943
rect 848 1923 850 1943
rect 1008 1923 1010 1943
rect 1160 1923 1162 1943
rect 679 1922 683 1923
rect 679 1917 683 1918
rect 687 1922 691 1923
rect 687 1917 691 1918
rect 847 1922 851 1923
rect 847 1917 851 1918
rect 1007 1922 1011 1923
rect 1007 1917 1011 1918
rect 1159 1922 1163 1923
rect 1159 1917 1163 1918
rect 688 1901 690 1917
rect 848 1901 850 1917
rect 1008 1901 1010 1917
rect 1160 1901 1162 1917
rect 686 1900 692 1901
rect 686 1896 687 1900
rect 691 1896 692 1900
rect 686 1895 692 1896
rect 846 1900 852 1901
rect 846 1896 847 1900
rect 851 1896 852 1900
rect 846 1895 852 1896
rect 1006 1900 1012 1901
rect 1006 1896 1007 1900
rect 1011 1896 1012 1900
rect 1006 1895 1012 1896
rect 1158 1900 1164 1901
rect 1158 1896 1159 1900
rect 1163 1896 1164 1900
rect 1158 1895 1164 1896
rect 594 1891 600 1892
rect 354 1886 360 1887
rect 534 1887 540 1888
rect 212 1852 214 1886
rect 246 1862 252 1863
rect 246 1858 247 1862
rect 251 1858 252 1862
rect 246 1857 252 1858
rect 198 1851 204 1852
rect 198 1847 199 1851
rect 203 1847 204 1851
rect 198 1846 204 1847
rect 210 1851 216 1852
rect 210 1847 211 1851
rect 215 1847 216 1851
rect 210 1846 216 1847
rect 248 1843 250 1857
rect 308 1852 310 1886
rect 306 1851 312 1852
rect 306 1847 307 1851
rect 311 1847 312 1851
rect 306 1846 312 1847
rect 111 1842 115 1843
rect 111 1837 115 1838
rect 143 1842 147 1843
rect 143 1837 147 1838
rect 247 1842 251 1843
rect 247 1837 251 1838
rect 287 1842 291 1843
rect 287 1837 291 1838
rect 112 1809 114 1837
rect 144 1827 146 1837
rect 288 1827 290 1837
rect 356 1836 358 1886
rect 534 1883 535 1887
rect 539 1883 540 1887
rect 594 1887 595 1891
rect 599 1887 600 1891
rect 594 1886 600 1887
rect 754 1891 760 1892
rect 754 1887 755 1891
rect 759 1887 760 1891
rect 754 1886 760 1887
rect 1078 1891 1084 1892
rect 1078 1887 1079 1891
rect 1083 1887 1084 1891
rect 1078 1886 1084 1887
rect 534 1882 540 1883
rect 382 1862 388 1863
rect 382 1858 383 1862
rect 387 1858 388 1862
rect 382 1857 388 1858
rect 534 1862 540 1863
rect 534 1858 535 1862
rect 539 1858 540 1862
rect 534 1857 540 1858
rect 384 1843 386 1857
rect 536 1843 538 1857
rect 596 1852 598 1886
rect 694 1862 700 1863
rect 694 1858 695 1862
rect 699 1858 700 1862
rect 694 1857 700 1858
rect 594 1851 600 1852
rect 594 1847 595 1851
rect 599 1847 600 1851
rect 594 1846 600 1847
rect 696 1843 698 1857
rect 756 1852 758 1886
rect 854 1862 860 1863
rect 854 1858 855 1862
rect 859 1858 860 1862
rect 854 1857 860 1858
rect 1014 1862 1020 1863
rect 1014 1858 1015 1862
rect 1019 1858 1020 1862
rect 1014 1857 1020 1858
rect 754 1851 760 1852
rect 754 1847 755 1851
rect 759 1847 760 1851
rect 754 1846 760 1847
rect 856 1843 858 1857
rect 878 1851 884 1852
rect 878 1847 879 1851
rect 883 1847 884 1851
rect 878 1846 884 1847
rect 383 1842 387 1843
rect 383 1837 387 1838
rect 471 1842 475 1843
rect 471 1837 475 1838
rect 535 1842 539 1843
rect 535 1837 539 1838
rect 663 1842 667 1843
rect 663 1837 667 1838
rect 695 1842 699 1843
rect 695 1837 699 1838
rect 847 1842 851 1843
rect 847 1837 851 1838
rect 855 1842 859 1843
rect 855 1837 859 1838
rect 294 1835 300 1836
rect 294 1831 295 1835
rect 299 1831 300 1835
rect 294 1830 300 1831
rect 354 1835 360 1836
rect 354 1831 355 1835
rect 359 1831 360 1835
rect 354 1830 360 1831
rect 142 1826 148 1827
rect 142 1822 143 1826
rect 147 1822 148 1826
rect 142 1821 148 1822
rect 286 1826 292 1827
rect 286 1822 287 1826
rect 291 1822 292 1826
rect 286 1821 292 1822
rect 110 1808 116 1809
rect 110 1804 111 1808
rect 115 1804 116 1808
rect 110 1803 116 1804
rect 296 1800 298 1830
rect 472 1827 474 1837
rect 486 1835 492 1836
rect 486 1831 487 1835
rect 491 1831 492 1835
rect 486 1830 492 1831
rect 522 1835 528 1836
rect 522 1831 523 1835
rect 527 1831 528 1835
rect 522 1830 528 1831
rect 470 1826 476 1827
rect 470 1822 471 1826
rect 475 1822 476 1826
rect 470 1821 476 1822
rect 166 1799 172 1800
rect 166 1795 167 1799
rect 171 1795 172 1799
rect 166 1794 172 1795
rect 294 1799 300 1800
rect 294 1795 295 1799
rect 299 1795 300 1799
rect 294 1794 300 1795
rect 110 1791 116 1792
rect 110 1787 111 1791
rect 115 1787 116 1791
rect 110 1786 116 1787
rect 134 1788 140 1789
rect 112 1759 114 1786
rect 134 1784 135 1788
rect 139 1784 140 1788
rect 134 1783 140 1784
rect 136 1759 138 1783
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 135 1758 139 1759
rect 135 1753 139 1754
rect 112 1734 114 1753
rect 136 1737 138 1753
rect 134 1736 140 1737
rect 110 1733 116 1734
rect 110 1729 111 1733
rect 115 1729 116 1733
rect 134 1732 135 1736
rect 139 1732 140 1736
rect 134 1731 140 1732
rect 110 1728 116 1729
rect 110 1716 116 1717
rect 110 1712 111 1716
rect 115 1712 116 1716
rect 110 1711 116 1712
rect 112 1679 114 1711
rect 142 1698 148 1699
rect 142 1694 143 1698
rect 147 1694 148 1698
rect 142 1693 148 1694
rect 144 1679 146 1693
rect 168 1688 170 1794
rect 278 1788 284 1789
rect 278 1784 279 1788
rect 283 1784 284 1788
rect 278 1783 284 1784
rect 462 1788 468 1789
rect 462 1784 463 1788
rect 467 1784 468 1788
rect 462 1783 468 1784
rect 280 1759 282 1783
rect 464 1759 466 1783
rect 215 1758 219 1759
rect 215 1753 219 1754
rect 279 1758 283 1759
rect 279 1753 283 1754
rect 343 1758 347 1759
rect 343 1753 347 1754
rect 463 1758 467 1759
rect 463 1753 467 1754
rect 216 1737 218 1753
rect 344 1737 346 1753
rect 214 1736 220 1737
rect 214 1732 215 1736
rect 219 1732 220 1736
rect 214 1731 220 1732
rect 342 1736 348 1737
rect 342 1732 343 1736
rect 347 1732 348 1736
rect 342 1731 348 1732
rect 488 1728 490 1830
rect 524 1800 526 1830
rect 664 1827 666 1837
rect 714 1835 720 1836
rect 714 1831 715 1835
rect 719 1831 720 1835
rect 714 1830 720 1831
rect 662 1826 668 1827
rect 662 1822 663 1826
rect 667 1822 668 1826
rect 662 1821 668 1822
rect 716 1800 718 1830
rect 848 1827 850 1837
rect 846 1826 852 1827
rect 846 1822 847 1826
rect 851 1822 852 1826
rect 846 1821 852 1822
rect 880 1800 882 1846
rect 1016 1843 1018 1857
rect 1080 1852 1082 1886
rect 1220 1884 1222 1990
rect 1312 1987 1314 1997
rect 1340 1996 1342 2038
rect 1348 2012 1350 2046
rect 1382 2022 1388 2023
rect 1382 2018 1383 2022
rect 1387 2018 1388 2022
rect 1382 2017 1388 2018
rect 1346 2011 1352 2012
rect 1346 2007 1347 2011
rect 1351 2007 1352 2011
rect 1346 2006 1352 2007
rect 1384 2003 1386 2017
rect 1444 2012 1446 2046
rect 1478 2022 1484 2023
rect 1478 2018 1479 2022
rect 1483 2018 1484 2022
rect 1478 2017 1484 2018
rect 1442 2011 1448 2012
rect 1442 2007 1443 2011
rect 1447 2007 1448 2011
rect 1442 2006 1448 2007
rect 1480 2003 1482 2017
rect 1540 2012 1542 2046
rect 1574 2022 1580 2023
rect 1574 2018 1575 2022
rect 1579 2018 1580 2022
rect 1574 2017 1580 2018
rect 1538 2011 1544 2012
rect 1538 2007 1539 2011
rect 1543 2007 1544 2011
rect 1538 2006 1544 2007
rect 1576 2003 1578 2017
rect 1636 2012 1638 2046
rect 1670 2022 1676 2023
rect 1670 2018 1671 2022
rect 1675 2018 1676 2022
rect 1670 2017 1676 2018
rect 1634 2011 1640 2012
rect 1634 2007 1635 2011
rect 1639 2007 1640 2011
rect 1634 2006 1640 2007
rect 1672 2003 1674 2017
rect 1732 2012 1734 2046
rect 1750 2022 1756 2023
rect 1750 2018 1751 2022
rect 1755 2018 1756 2022
rect 1750 2017 1756 2018
rect 1730 2011 1736 2012
rect 1730 2007 1731 2011
rect 1735 2007 1736 2011
rect 1730 2006 1736 2007
rect 1752 2003 1754 2017
rect 1780 2012 1782 2086
rect 1832 2083 1834 2114
rect 1870 2111 1876 2112
rect 1870 2107 1871 2111
rect 1875 2107 1876 2111
rect 1870 2106 1876 2107
rect 1894 2108 1900 2109
rect 1831 2082 1835 2083
rect 1872 2079 1874 2106
rect 1894 2104 1895 2108
rect 1899 2104 1900 2108
rect 1894 2103 1900 2104
rect 1974 2108 1980 2109
rect 1974 2104 1975 2108
rect 1979 2104 1980 2108
rect 1974 2103 1980 2104
rect 1896 2079 1898 2103
rect 1976 2079 1978 2103
rect 1831 2077 1835 2078
rect 1871 2078 1875 2079
rect 1832 2058 1834 2077
rect 1871 2073 1875 2074
rect 1895 2078 1899 2079
rect 1895 2073 1899 2074
rect 1967 2078 1971 2079
rect 1967 2073 1971 2074
rect 1975 2078 1979 2079
rect 1975 2073 1979 2074
rect 1830 2057 1836 2058
rect 1830 2053 1831 2057
rect 1835 2053 1836 2057
rect 1872 2054 1874 2073
rect 1968 2057 1970 2073
rect 1966 2056 1972 2057
rect 1830 2052 1836 2053
rect 1870 2053 1876 2054
rect 1870 2049 1871 2053
rect 1875 2049 1876 2053
rect 1966 2052 1967 2056
rect 1971 2052 1972 2056
rect 1966 2051 1972 2052
rect 1870 2048 1876 2049
rect 2052 2048 2054 2150
rect 2112 2147 2114 2157
rect 2162 2155 2168 2156
rect 2162 2151 2163 2155
rect 2167 2151 2168 2155
rect 2162 2150 2168 2151
rect 2110 2146 2116 2147
rect 2110 2142 2111 2146
rect 2115 2142 2116 2146
rect 2110 2141 2116 2142
rect 2164 2120 2166 2150
rect 2248 2147 2250 2157
rect 2298 2155 2304 2156
rect 2298 2151 2299 2155
rect 2303 2151 2304 2155
rect 2298 2150 2304 2151
rect 2246 2146 2252 2147
rect 2246 2142 2247 2146
rect 2251 2142 2252 2146
rect 2246 2141 2252 2142
rect 2300 2120 2302 2150
rect 2392 2147 2394 2157
rect 2390 2146 2396 2147
rect 2390 2142 2391 2146
rect 2395 2142 2396 2146
rect 2390 2141 2396 2142
rect 2400 2120 2402 2158
rect 2407 2157 2411 2158
rect 2503 2162 2507 2163
rect 2503 2157 2507 2158
rect 2543 2162 2547 2163
rect 2543 2157 2547 2158
rect 2544 2147 2546 2157
rect 2564 2156 2566 2206
rect 2606 2182 2612 2183
rect 2606 2178 2607 2182
rect 2611 2178 2612 2182
rect 2606 2177 2612 2178
rect 2608 2163 2610 2177
rect 2632 2172 2634 2270
rect 2670 2264 2676 2265
rect 2670 2260 2671 2264
rect 2675 2260 2676 2264
rect 2670 2259 2676 2260
rect 2750 2264 2756 2265
rect 2750 2260 2751 2264
rect 2755 2260 2756 2264
rect 2750 2259 2756 2260
rect 2838 2264 2844 2265
rect 2838 2260 2839 2264
rect 2843 2260 2844 2264
rect 2838 2259 2844 2260
rect 2926 2264 2932 2265
rect 2926 2260 2927 2264
rect 2931 2260 2932 2264
rect 2926 2259 2932 2260
rect 2672 2243 2674 2259
rect 2752 2243 2754 2259
rect 2840 2243 2842 2259
rect 2928 2243 2930 2259
rect 2671 2242 2675 2243
rect 2671 2237 2675 2238
rect 2719 2242 2723 2243
rect 2719 2237 2723 2238
rect 2751 2242 2755 2243
rect 2751 2237 2755 2238
rect 2839 2242 2843 2243
rect 2839 2237 2843 2238
rect 2855 2242 2859 2243
rect 2855 2237 2859 2238
rect 2927 2242 2931 2243
rect 2927 2237 2931 2238
rect 3007 2242 3011 2243
rect 3007 2237 3011 2238
rect 3175 2242 3179 2243
rect 3175 2237 3179 2238
rect 3351 2242 3355 2243
rect 3351 2237 3355 2238
rect 2720 2221 2722 2237
rect 2856 2221 2858 2237
rect 3008 2221 3010 2237
rect 3176 2221 3178 2237
rect 3352 2221 3354 2237
rect 2718 2220 2724 2221
rect 2718 2216 2719 2220
rect 2723 2216 2724 2220
rect 2718 2215 2724 2216
rect 2854 2220 2860 2221
rect 2854 2216 2855 2220
rect 2859 2216 2860 2220
rect 2854 2215 2860 2216
rect 3006 2220 3012 2221
rect 3006 2216 3007 2220
rect 3011 2216 3012 2220
rect 3006 2215 3012 2216
rect 3174 2220 3180 2221
rect 3174 2216 3175 2220
rect 3179 2216 3180 2220
rect 3174 2215 3180 2216
rect 3350 2220 3356 2221
rect 3350 2216 3351 2220
rect 3355 2216 3356 2220
rect 3350 2215 3356 2216
rect 3420 2212 3422 2322
rect 3512 2319 3514 2333
rect 3536 2328 3538 2430
rect 3590 2427 3596 2428
rect 3590 2423 3591 2427
rect 3595 2423 3596 2427
rect 3590 2422 3596 2423
rect 3592 2399 3594 2422
rect 3591 2398 3595 2399
rect 3591 2393 3595 2394
rect 3592 2374 3594 2393
rect 3590 2373 3596 2374
rect 3590 2369 3591 2373
rect 3595 2369 3596 2373
rect 3590 2368 3596 2369
rect 3570 2367 3576 2368
rect 3570 2363 3571 2367
rect 3575 2363 3576 2367
rect 3570 2362 3576 2363
rect 3534 2327 3540 2328
rect 3534 2323 3535 2327
rect 3539 2323 3540 2327
rect 3534 2322 3540 2323
rect 3511 2318 3515 2319
rect 3511 2313 3515 2314
rect 3503 2242 3507 2243
rect 3503 2237 3507 2238
rect 3504 2221 3506 2237
rect 3502 2220 3508 2221
rect 3502 2216 3503 2220
rect 3507 2216 3508 2220
rect 3502 2215 3508 2216
rect 2678 2211 2684 2212
rect 2678 2207 2679 2211
rect 2683 2207 2684 2211
rect 2678 2206 2684 2207
rect 2786 2211 2792 2212
rect 2786 2207 2787 2211
rect 2791 2207 2792 2211
rect 2786 2206 2792 2207
rect 3074 2211 3080 2212
rect 3074 2207 3075 2211
rect 3079 2207 3080 2211
rect 3074 2206 3080 2207
rect 3082 2211 3088 2212
rect 3082 2207 3083 2211
rect 3087 2207 3088 2211
rect 3082 2206 3088 2207
rect 3418 2211 3424 2212
rect 3418 2207 3419 2211
rect 3423 2207 3424 2211
rect 3418 2206 3424 2207
rect 2680 2172 2682 2206
rect 2726 2182 2732 2183
rect 2726 2178 2727 2182
rect 2731 2178 2732 2182
rect 2726 2177 2732 2178
rect 2735 2180 2739 2181
rect 2630 2171 2636 2172
rect 2630 2167 2631 2171
rect 2635 2167 2636 2171
rect 2630 2166 2636 2167
rect 2678 2171 2684 2172
rect 2678 2167 2679 2171
rect 2683 2167 2684 2171
rect 2678 2166 2684 2167
rect 2728 2163 2730 2177
rect 2735 2175 2739 2176
rect 2607 2162 2611 2163
rect 2607 2157 2611 2158
rect 2695 2162 2699 2163
rect 2695 2157 2699 2158
rect 2727 2162 2731 2163
rect 2727 2157 2731 2158
rect 2562 2155 2568 2156
rect 2562 2151 2563 2155
rect 2567 2151 2568 2155
rect 2562 2150 2568 2151
rect 2696 2147 2698 2157
rect 2736 2156 2738 2175
rect 2788 2172 2790 2206
rect 2862 2182 2868 2183
rect 2862 2178 2863 2182
rect 2867 2178 2868 2182
rect 2862 2177 2868 2178
rect 3014 2182 3020 2183
rect 3014 2178 3015 2182
rect 3019 2178 3020 2182
rect 3014 2177 3020 2178
rect 2786 2171 2792 2172
rect 2786 2167 2787 2171
rect 2791 2167 2792 2171
rect 2786 2166 2792 2167
rect 2864 2163 2866 2177
rect 3016 2163 3018 2177
rect 3076 2172 3078 2206
rect 3084 2181 3086 2206
rect 3562 2203 3568 2204
rect 3562 2199 3563 2203
rect 3567 2199 3568 2203
rect 3562 2198 3568 2199
rect 3182 2182 3188 2183
rect 3083 2180 3087 2181
rect 3182 2178 3183 2182
rect 3187 2178 3188 2182
rect 3182 2177 3188 2178
rect 3358 2182 3364 2183
rect 3358 2178 3359 2182
rect 3363 2178 3364 2182
rect 3358 2177 3364 2178
rect 3510 2182 3516 2183
rect 3510 2178 3511 2182
rect 3515 2178 3516 2182
rect 3510 2177 3516 2178
rect 3083 2175 3087 2176
rect 3074 2171 3080 2172
rect 3074 2167 3075 2171
rect 3079 2167 3080 2171
rect 3074 2166 3080 2167
rect 3184 2163 3186 2177
rect 3360 2163 3362 2177
rect 3386 2171 3392 2172
rect 3386 2167 3387 2171
rect 3391 2167 3392 2171
rect 3386 2166 3392 2167
rect 2847 2162 2851 2163
rect 2847 2157 2851 2158
rect 2863 2162 2867 2163
rect 2863 2157 2867 2158
rect 3007 2162 3011 2163
rect 3007 2157 3011 2158
rect 3015 2162 3019 2163
rect 3015 2157 3019 2158
rect 3175 2162 3179 2163
rect 3175 2157 3179 2158
rect 3183 2162 3187 2163
rect 3183 2157 3187 2158
rect 3351 2162 3355 2163
rect 3351 2157 3355 2158
rect 3359 2162 3363 2163
rect 3359 2157 3363 2158
rect 2734 2155 2740 2156
rect 2734 2151 2735 2155
rect 2739 2151 2740 2155
rect 2734 2150 2740 2151
rect 2746 2155 2752 2156
rect 2746 2151 2747 2155
rect 2751 2151 2752 2155
rect 2746 2150 2752 2151
rect 2542 2146 2548 2147
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2694 2146 2700 2147
rect 2694 2142 2695 2146
rect 2699 2142 2700 2146
rect 2694 2141 2700 2142
rect 2748 2120 2750 2150
rect 2848 2147 2850 2157
rect 2898 2155 2904 2156
rect 2898 2151 2899 2155
rect 2903 2151 2904 2155
rect 2898 2150 2904 2151
rect 2846 2146 2852 2147
rect 2846 2142 2847 2146
rect 2851 2142 2852 2146
rect 2846 2141 2852 2142
rect 2900 2120 2902 2150
rect 3008 2147 3010 2157
rect 3058 2155 3064 2156
rect 3058 2151 3059 2155
rect 3063 2151 3064 2155
rect 3058 2150 3064 2151
rect 3006 2146 3012 2147
rect 3006 2142 3007 2146
rect 3011 2142 3012 2146
rect 3006 2141 3012 2142
rect 3060 2120 3062 2150
rect 3176 2147 3178 2157
rect 3226 2155 3232 2156
rect 3226 2151 3227 2155
rect 3231 2151 3232 2155
rect 3226 2150 3232 2151
rect 3174 2146 3180 2147
rect 3174 2142 3175 2146
rect 3179 2142 3180 2146
rect 3174 2141 3180 2142
rect 3228 2120 3230 2150
rect 3352 2147 3354 2157
rect 3350 2146 3356 2147
rect 3350 2142 3351 2146
rect 3355 2142 3356 2146
rect 3350 2141 3356 2142
rect 2162 2119 2168 2120
rect 2162 2115 2163 2119
rect 2167 2115 2168 2119
rect 2162 2114 2168 2115
rect 2298 2119 2304 2120
rect 2298 2115 2299 2119
rect 2303 2115 2304 2119
rect 2298 2114 2304 2115
rect 2398 2119 2404 2120
rect 2398 2115 2399 2119
rect 2403 2115 2404 2119
rect 2398 2114 2404 2115
rect 2746 2119 2752 2120
rect 2746 2115 2747 2119
rect 2751 2115 2752 2119
rect 2746 2114 2752 2115
rect 2898 2119 2904 2120
rect 2898 2115 2899 2119
rect 2903 2115 2904 2119
rect 2898 2114 2904 2115
rect 3058 2119 3064 2120
rect 3058 2115 3059 2119
rect 3063 2115 3064 2119
rect 3058 2114 3064 2115
rect 3226 2119 3232 2120
rect 3226 2115 3227 2119
rect 3231 2115 3232 2119
rect 3226 2114 3232 2115
rect 2102 2108 2108 2109
rect 2102 2104 2103 2108
rect 2107 2104 2108 2108
rect 2102 2103 2108 2104
rect 2238 2108 2244 2109
rect 2238 2104 2239 2108
rect 2243 2104 2244 2108
rect 2238 2103 2244 2104
rect 2382 2108 2388 2109
rect 2382 2104 2383 2108
rect 2387 2104 2388 2108
rect 2382 2103 2388 2104
rect 2534 2108 2540 2109
rect 2534 2104 2535 2108
rect 2539 2104 2540 2108
rect 2534 2103 2540 2104
rect 2686 2108 2692 2109
rect 2686 2104 2687 2108
rect 2691 2104 2692 2108
rect 2686 2103 2692 2104
rect 2838 2108 2844 2109
rect 2838 2104 2839 2108
rect 2843 2104 2844 2108
rect 2838 2103 2844 2104
rect 2998 2108 3004 2109
rect 2998 2104 2999 2108
rect 3003 2104 3004 2108
rect 2998 2103 3004 2104
rect 3166 2108 3172 2109
rect 3166 2104 3167 2108
rect 3171 2104 3172 2108
rect 3166 2103 3172 2104
rect 3342 2108 3348 2109
rect 3342 2104 3343 2108
rect 3347 2104 3348 2108
rect 3342 2103 3348 2104
rect 2104 2079 2106 2103
rect 2240 2079 2242 2103
rect 2384 2079 2386 2103
rect 2482 2091 2488 2092
rect 2482 2087 2483 2091
rect 2487 2087 2488 2091
rect 2482 2086 2488 2087
rect 2103 2078 2107 2079
rect 2103 2073 2107 2074
rect 2215 2078 2219 2079
rect 2215 2073 2219 2074
rect 2239 2078 2243 2079
rect 2239 2073 2243 2074
rect 2383 2078 2387 2079
rect 2383 2073 2387 2074
rect 2447 2078 2451 2079
rect 2447 2073 2451 2074
rect 2216 2057 2218 2073
rect 2448 2057 2450 2073
rect 2214 2056 2220 2057
rect 2214 2052 2215 2056
rect 2219 2052 2220 2056
rect 2214 2051 2220 2052
rect 2446 2056 2452 2057
rect 2446 2052 2447 2056
rect 2451 2052 2452 2056
rect 2446 2051 2452 2052
rect 2050 2047 2056 2048
rect 2050 2043 2051 2047
rect 2055 2043 2056 2047
rect 2050 2042 2056 2043
rect 2282 2047 2288 2048
rect 2282 2043 2283 2047
rect 2287 2043 2288 2047
rect 2282 2042 2288 2043
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 2274 2039 2280 2040
rect 1830 2035 1836 2036
rect 1870 2036 1876 2037
rect 1778 2011 1784 2012
rect 1778 2007 1779 2011
rect 1783 2007 1784 2011
rect 1778 2006 1784 2007
rect 1832 2003 1834 2035
rect 1870 2032 1871 2036
rect 1875 2032 1876 2036
rect 2274 2035 2275 2039
rect 2279 2035 2280 2039
rect 2274 2034 2280 2035
rect 1870 2031 1876 2032
rect 1872 2003 1874 2031
rect 1974 2018 1980 2019
rect 1974 2014 1975 2018
rect 1979 2014 1980 2018
rect 1974 2013 1980 2014
rect 2222 2018 2228 2019
rect 2222 2014 2223 2018
rect 2227 2014 2228 2018
rect 2222 2013 2228 2014
rect 1976 2003 1978 2013
rect 1998 2007 2004 2008
rect 1998 2003 1999 2007
rect 2003 2003 2004 2007
rect 2224 2003 2226 2013
rect 1383 2002 1387 2003
rect 1383 1997 1387 1998
rect 1447 2002 1451 2003
rect 1447 1997 1451 1998
rect 1479 2002 1483 2003
rect 1479 1997 1483 1998
rect 1575 2002 1579 2003
rect 1575 1997 1579 1998
rect 1583 2002 1587 2003
rect 1583 1997 1587 1998
rect 1671 2002 1675 2003
rect 1671 1997 1675 1998
rect 1719 2002 1723 2003
rect 1719 1997 1723 1998
rect 1751 2002 1755 2003
rect 1751 1997 1755 1998
rect 1831 2002 1835 2003
rect 1831 1997 1835 1998
rect 1871 2002 1875 2003
rect 1871 1997 1875 1998
rect 1959 2002 1963 2003
rect 1959 1997 1963 1998
rect 1975 2002 1979 2003
rect 1998 2002 2004 2003
rect 2079 2002 2083 2003
rect 1975 1997 1979 1998
rect 1338 1995 1344 1996
rect 1338 1991 1339 1995
rect 1343 1991 1344 1995
rect 1338 1990 1344 1991
rect 1362 1995 1368 1996
rect 1362 1991 1363 1995
rect 1367 1991 1368 1995
rect 1362 1990 1368 1991
rect 1310 1986 1316 1987
rect 1310 1982 1311 1986
rect 1315 1982 1316 1986
rect 1310 1981 1316 1982
rect 1364 1960 1366 1990
rect 1448 1987 1450 1997
rect 1498 1995 1504 1996
rect 1498 1991 1499 1995
rect 1503 1991 1504 1995
rect 1498 1990 1504 1991
rect 1446 1986 1452 1987
rect 1446 1982 1447 1986
rect 1451 1982 1452 1986
rect 1446 1981 1452 1982
rect 1500 1960 1502 1990
rect 1584 1987 1586 1997
rect 1634 1995 1640 1996
rect 1634 1991 1635 1995
rect 1639 1991 1640 1995
rect 1634 1990 1640 1991
rect 1582 1986 1588 1987
rect 1582 1982 1583 1986
rect 1587 1982 1588 1986
rect 1582 1981 1588 1982
rect 1636 1960 1638 1990
rect 1720 1987 1722 1997
rect 1718 1986 1724 1987
rect 1718 1982 1719 1986
rect 1723 1982 1724 1986
rect 1718 1981 1724 1982
rect 1832 1969 1834 1997
rect 1872 1969 1874 1997
rect 1960 1987 1962 1997
rect 1958 1986 1964 1987
rect 1958 1982 1959 1986
rect 1963 1982 1964 1986
rect 1958 1981 1964 1982
rect 1830 1968 1836 1969
rect 1830 1964 1831 1968
rect 1835 1964 1836 1968
rect 1830 1963 1836 1964
rect 1870 1968 1876 1969
rect 1870 1964 1871 1968
rect 1875 1964 1876 1968
rect 1870 1963 1876 1964
rect 2000 1960 2002 2002
rect 2079 1997 2083 1998
rect 2199 2002 2203 2003
rect 2199 1997 2203 1998
rect 2223 2002 2227 2003
rect 2223 1997 2227 1998
rect 2080 1987 2082 1997
rect 2086 1995 2092 1996
rect 2086 1991 2087 1995
rect 2091 1991 2092 1995
rect 2086 1990 2092 1991
rect 2078 1986 2084 1987
rect 2078 1982 2079 1986
rect 2083 1982 2084 1986
rect 2078 1981 2084 1982
rect 2088 1960 2090 1990
rect 2200 1987 2202 1997
rect 2276 1996 2278 2034
rect 2284 2008 2286 2042
rect 2454 2018 2460 2019
rect 2454 2014 2455 2018
rect 2459 2014 2460 2018
rect 2454 2013 2460 2014
rect 2282 2007 2288 2008
rect 2282 2003 2283 2007
rect 2287 2003 2288 2007
rect 2456 2003 2458 2013
rect 2484 2008 2486 2086
rect 2536 2079 2538 2103
rect 2688 2079 2690 2103
rect 2840 2079 2842 2103
rect 3000 2079 3002 2103
rect 3168 2079 3170 2103
rect 3306 2091 3312 2092
rect 3306 2087 3307 2091
rect 3311 2087 3312 2091
rect 3306 2086 3312 2087
rect 2535 2078 2539 2079
rect 2535 2073 2539 2074
rect 2655 2078 2659 2079
rect 2655 2073 2659 2074
rect 2687 2078 2691 2079
rect 2687 2073 2691 2074
rect 2839 2078 2843 2079
rect 2839 2073 2843 2074
rect 2999 2078 3003 2079
rect 2999 2073 3003 2074
rect 3143 2078 3147 2079
rect 3143 2073 3147 2074
rect 3167 2078 3171 2079
rect 3167 2073 3171 2074
rect 3271 2078 3275 2079
rect 3271 2073 3275 2074
rect 2656 2057 2658 2073
rect 2840 2057 2842 2073
rect 3000 2057 3002 2073
rect 3144 2057 3146 2073
rect 3272 2057 3274 2073
rect 2654 2056 2660 2057
rect 2654 2052 2655 2056
rect 2659 2052 2660 2056
rect 2654 2051 2660 2052
rect 2838 2056 2844 2057
rect 2838 2052 2839 2056
rect 2843 2052 2844 2056
rect 2838 2051 2844 2052
rect 2998 2056 3004 2057
rect 2998 2052 2999 2056
rect 3003 2052 3004 2056
rect 2998 2051 3004 2052
rect 3142 2056 3148 2057
rect 3142 2052 3143 2056
rect 3147 2052 3148 2056
rect 3142 2051 3148 2052
rect 3270 2056 3276 2057
rect 3270 2052 3271 2056
rect 3275 2052 3276 2056
rect 3270 2051 3276 2052
rect 2754 2047 2760 2048
rect 2754 2043 2755 2047
rect 2759 2043 2760 2047
rect 2754 2042 2760 2043
rect 2942 2047 2948 2048
rect 2942 2043 2943 2047
rect 2947 2043 2948 2047
rect 2942 2042 2948 2043
rect 3078 2047 3084 2048
rect 3078 2043 3079 2047
rect 3083 2043 3084 2047
rect 3078 2042 3084 2043
rect 3086 2047 3092 2048
rect 3086 2043 3087 2047
rect 3091 2043 3092 2047
rect 3086 2042 3092 2043
rect 3210 2047 3216 2048
rect 3210 2043 3211 2047
rect 3215 2043 3216 2047
rect 3210 2042 3216 2043
rect 2662 2018 2668 2019
rect 2662 2014 2663 2018
rect 2667 2014 2668 2018
rect 2662 2013 2668 2014
rect 2482 2007 2488 2008
rect 2482 2003 2483 2007
rect 2487 2003 2488 2007
rect 2664 2003 2666 2013
rect 2687 2012 2691 2013
rect 2756 2008 2758 2042
rect 2846 2018 2852 2019
rect 2846 2014 2847 2018
rect 2851 2014 2852 2018
rect 2846 2013 2852 2014
rect 2686 2007 2692 2008
rect 2686 2003 2687 2007
rect 2691 2003 2692 2007
rect 2754 2007 2760 2008
rect 2754 2003 2755 2007
rect 2759 2003 2760 2007
rect 2848 2003 2850 2013
rect 2944 2008 2946 2042
rect 3006 2018 3012 2019
rect 3006 2014 3007 2018
rect 3011 2014 3012 2018
rect 3006 2013 3012 2014
rect 2942 2007 2948 2008
rect 2942 2003 2943 2007
rect 2947 2003 2948 2007
rect 3008 2003 3010 2013
rect 2282 2002 2288 2003
rect 2319 2002 2323 2003
rect 2319 1997 2323 1998
rect 2447 2002 2451 2003
rect 2447 1997 2451 1998
rect 2455 2002 2459 2003
rect 2482 2002 2488 2003
rect 2583 2002 2587 2003
rect 2455 1997 2459 1998
rect 2583 1997 2587 1998
rect 2663 2002 2667 2003
rect 2686 2002 2692 2003
rect 2743 2002 2747 2003
rect 2754 2002 2760 2003
rect 2847 2002 2851 2003
rect 2663 1997 2667 1998
rect 2743 1997 2747 1998
rect 2847 1997 2851 1998
rect 2919 2002 2923 2003
rect 2942 2002 2948 2003
rect 3007 2002 3011 2003
rect 2919 1997 2923 1998
rect 3007 1997 3011 1998
rect 2206 1995 2212 1996
rect 2206 1991 2207 1995
rect 2211 1991 2212 1995
rect 2274 1995 2280 1996
rect 2206 1990 2212 1991
rect 2222 1991 2228 1992
rect 2198 1986 2204 1987
rect 2198 1982 2199 1986
rect 2203 1982 2204 1986
rect 2198 1981 2204 1982
rect 2208 1960 2210 1990
rect 2222 1987 2223 1991
rect 2227 1987 2228 1991
rect 2274 1991 2275 1995
rect 2279 1991 2280 1995
rect 2274 1990 2280 1991
rect 2320 1987 2322 1997
rect 2448 1987 2450 1997
rect 2584 1987 2586 1997
rect 2590 1995 2596 1996
rect 2590 1991 2591 1995
rect 2595 1991 2596 1995
rect 2590 1990 2596 1991
rect 2222 1986 2228 1987
rect 2318 1986 2324 1987
rect 1362 1959 1368 1960
rect 1362 1955 1363 1959
rect 1367 1955 1368 1959
rect 1362 1954 1368 1955
rect 1498 1959 1504 1960
rect 1498 1955 1499 1959
rect 1503 1955 1504 1959
rect 1498 1954 1504 1955
rect 1634 1959 1640 1960
rect 1634 1955 1635 1959
rect 1639 1955 1640 1959
rect 1634 1954 1640 1955
rect 1998 1959 2004 1960
rect 1998 1955 1999 1959
rect 2003 1955 2004 1959
rect 1998 1954 2004 1955
rect 2086 1959 2092 1960
rect 2086 1955 2087 1959
rect 2091 1955 2092 1959
rect 2086 1954 2092 1955
rect 2206 1959 2212 1960
rect 2206 1955 2207 1959
rect 2211 1955 2212 1959
rect 2206 1954 2212 1955
rect 1830 1951 1836 1952
rect 1302 1948 1308 1949
rect 1302 1944 1303 1948
rect 1307 1944 1308 1948
rect 1302 1943 1308 1944
rect 1438 1948 1444 1949
rect 1438 1944 1439 1948
rect 1443 1944 1444 1948
rect 1438 1943 1444 1944
rect 1574 1948 1580 1949
rect 1574 1944 1575 1948
rect 1579 1944 1580 1948
rect 1574 1943 1580 1944
rect 1710 1948 1716 1949
rect 1710 1944 1711 1948
rect 1715 1944 1716 1948
rect 1830 1947 1831 1951
rect 1835 1947 1836 1951
rect 1830 1946 1836 1947
rect 1870 1951 1876 1952
rect 1870 1947 1871 1951
rect 1875 1947 1876 1951
rect 1870 1946 1876 1947
rect 1950 1948 1956 1949
rect 1710 1943 1716 1944
rect 1304 1923 1306 1943
rect 1440 1923 1442 1943
rect 1576 1923 1578 1943
rect 1712 1923 1714 1943
rect 1726 1931 1732 1932
rect 1726 1927 1727 1931
rect 1731 1927 1732 1931
rect 1726 1926 1732 1927
rect 1303 1922 1307 1923
rect 1303 1917 1307 1918
rect 1439 1922 1443 1923
rect 1439 1917 1443 1918
rect 1455 1922 1459 1923
rect 1455 1917 1459 1918
rect 1575 1922 1579 1923
rect 1575 1917 1579 1918
rect 1607 1922 1611 1923
rect 1607 1917 1611 1918
rect 1711 1922 1715 1923
rect 1711 1917 1715 1918
rect 1304 1901 1306 1917
rect 1456 1901 1458 1917
rect 1608 1901 1610 1917
rect 1302 1900 1308 1901
rect 1302 1896 1303 1900
rect 1307 1896 1308 1900
rect 1302 1895 1308 1896
rect 1454 1900 1460 1901
rect 1454 1896 1455 1900
rect 1459 1896 1460 1900
rect 1454 1895 1460 1896
rect 1606 1900 1612 1901
rect 1606 1896 1607 1900
rect 1611 1896 1612 1900
rect 1606 1895 1612 1896
rect 1226 1891 1232 1892
rect 1226 1887 1227 1891
rect 1231 1887 1232 1891
rect 1226 1886 1232 1887
rect 1370 1891 1376 1892
rect 1370 1887 1371 1891
rect 1375 1887 1376 1891
rect 1370 1886 1376 1887
rect 1522 1891 1528 1892
rect 1522 1887 1523 1891
rect 1527 1887 1528 1891
rect 1522 1886 1528 1887
rect 1218 1883 1224 1884
rect 1218 1879 1219 1883
rect 1223 1879 1224 1883
rect 1218 1878 1224 1879
rect 1166 1862 1172 1863
rect 1166 1858 1167 1862
rect 1171 1858 1172 1862
rect 1166 1857 1172 1858
rect 1038 1851 1044 1852
rect 1038 1847 1039 1851
rect 1043 1847 1044 1851
rect 1038 1846 1044 1847
rect 1078 1851 1084 1852
rect 1078 1847 1079 1851
rect 1083 1847 1084 1851
rect 1078 1846 1084 1847
rect 1015 1842 1019 1843
rect 1015 1837 1019 1838
rect 1023 1842 1027 1843
rect 1023 1837 1027 1838
rect 1024 1827 1026 1837
rect 1022 1826 1028 1827
rect 1022 1822 1023 1826
rect 1027 1822 1028 1826
rect 1022 1821 1028 1822
rect 1040 1800 1042 1846
rect 1168 1843 1170 1857
rect 1167 1842 1171 1843
rect 1167 1837 1171 1838
rect 1191 1842 1195 1843
rect 1191 1837 1195 1838
rect 1102 1835 1108 1836
rect 1102 1831 1103 1835
rect 1107 1831 1108 1835
rect 1102 1830 1108 1831
rect 522 1799 528 1800
rect 522 1795 523 1799
rect 527 1795 528 1799
rect 522 1794 528 1795
rect 714 1799 720 1800
rect 714 1795 715 1799
rect 719 1795 720 1799
rect 714 1794 720 1795
rect 878 1799 884 1800
rect 878 1795 879 1799
rect 883 1795 884 1799
rect 878 1794 884 1795
rect 1038 1799 1044 1800
rect 1038 1795 1039 1799
rect 1043 1795 1044 1799
rect 1038 1794 1044 1795
rect 654 1788 660 1789
rect 654 1784 655 1788
rect 659 1784 660 1788
rect 654 1783 660 1784
rect 838 1788 844 1789
rect 838 1784 839 1788
rect 843 1784 844 1788
rect 838 1783 844 1784
rect 1014 1788 1020 1789
rect 1014 1784 1015 1788
rect 1019 1784 1020 1788
rect 1014 1783 1020 1784
rect 656 1759 658 1783
rect 840 1759 842 1783
rect 1016 1759 1018 1783
rect 495 1758 499 1759
rect 495 1753 499 1754
rect 655 1758 659 1759
rect 655 1753 659 1754
rect 663 1758 667 1759
rect 663 1753 667 1754
rect 839 1758 843 1759
rect 839 1753 843 1754
rect 1007 1758 1011 1759
rect 1007 1753 1011 1754
rect 1015 1758 1019 1759
rect 1015 1753 1019 1754
rect 496 1737 498 1753
rect 664 1737 666 1753
rect 840 1737 842 1753
rect 1008 1737 1010 1753
rect 494 1736 500 1737
rect 494 1732 495 1736
rect 499 1732 500 1736
rect 494 1731 500 1732
rect 662 1736 668 1737
rect 662 1732 663 1736
rect 667 1732 668 1736
rect 662 1731 668 1732
rect 838 1736 844 1737
rect 838 1732 839 1736
rect 843 1732 844 1736
rect 838 1731 844 1732
rect 1006 1736 1012 1737
rect 1006 1732 1007 1736
rect 1011 1732 1012 1736
rect 1006 1731 1012 1732
rect 1104 1728 1106 1830
rect 1192 1827 1194 1837
rect 1228 1836 1230 1886
rect 1310 1862 1316 1863
rect 1310 1858 1311 1862
rect 1315 1858 1316 1862
rect 1310 1857 1316 1858
rect 1312 1843 1314 1857
rect 1372 1852 1374 1886
rect 1462 1862 1468 1863
rect 1462 1858 1463 1862
rect 1467 1858 1468 1862
rect 1462 1857 1468 1858
rect 1370 1851 1376 1852
rect 1370 1847 1371 1851
rect 1375 1847 1376 1851
rect 1370 1846 1376 1847
rect 1464 1843 1466 1857
rect 1524 1852 1526 1886
rect 1614 1862 1620 1863
rect 1614 1858 1615 1862
rect 1619 1858 1620 1862
rect 1614 1857 1620 1858
rect 1522 1851 1528 1852
rect 1522 1847 1523 1851
rect 1527 1847 1528 1851
rect 1522 1846 1528 1847
rect 1616 1843 1618 1857
rect 1728 1852 1730 1926
rect 1832 1923 1834 1946
rect 1831 1922 1835 1923
rect 1872 1919 1874 1946
rect 1950 1944 1951 1948
rect 1955 1944 1956 1948
rect 1950 1943 1956 1944
rect 2070 1948 2076 1949
rect 2070 1944 2071 1948
rect 2075 1944 2076 1948
rect 2070 1943 2076 1944
rect 2190 1948 2196 1949
rect 2190 1944 2191 1948
rect 2195 1944 2196 1948
rect 2190 1943 2196 1944
rect 1952 1919 1954 1943
rect 2072 1919 2074 1943
rect 2192 1919 2194 1943
rect 1831 1917 1835 1918
rect 1871 1918 1875 1919
rect 1832 1898 1834 1917
rect 1871 1913 1875 1914
rect 1951 1918 1955 1919
rect 1951 1913 1955 1914
rect 2063 1918 2067 1919
rect 2063 1913 2067 1914
rect 2071 1918 2075 1919
rect 2071 1913 2075 1914
rect 2151 1918 2155 1919
rect 2151 1913 2155 1914
rect 2191 1918 2195 1919
rect 2191 1913 2195 1914
rect 1830 1897 1836 1898
rect 1830 1893 1831 1897
rect 1835 1893 1836 1897
rect 1872 1894 1874 1913
rect 2064 1897 2066 1913
rect 2152 1897 2154 1913
rect 2062 1896 2068 1897
rect 1830 1892 1836 1893
rect 1870 1893 1876 1894
rect 1870 1889 1871 1893
rect 1875 1889 1876 1893
rect 2062 1892 2063 1896
rect 2067 1892 2068 1896
rect 2062 1891 2068 1892
rect 2150 1896 2156 1897
rect 2150 1892 2151 1896
rect 2155 1892 2156 1896
rect 2150 1891 2156 1892
rect 1870 1888 1876 1889
rect 2224 1888 2226 1986
rect 2318 1982 2319 1986
rect 2323 1982 2324 1986
rect 2318 1981 2324 1982
rect 2446 1986 2452 1987
rect 2446 1982 2447 1986
rect 2451 1982 2452 1986
rect 2446 1981 2452 1982
rect 2582 1986 2588 1987
rect 2582 1982 2583 1986
rect 2587 1982 2588 1986
rect 2582 1981 2588 1982
rect 2592 1960 2594 1990
rect 2744 1987 2746 1997
rect 2750 1995 2756 1996
rect 2750 1991 2751 1995
rect 2755 1991 2756 1995
rect 2750 1990 2756 1991
rect 2742 1986 2748 1987
rect 2742 1982 2743 1986
rect 2747 1982 2748 1986
rect 2742 1981 2748 1982
rect 2752 1960 2754 1990
rect 2920 1987 2922 1997
rect 3080 1996 3082 2042
rect 3088 2013 3090 2042
rect 3150 2018 3156 2019
rect 3150 2014 3151 2018
rect 3155 2014 3156 2018
rect 3150 2013 3156 2014
rect 3087 2012 3091 2013
rect 3087 2007 3091 2008
rect 3152 2003 3154 2013
rect 3212 2008 3214 2042
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3210 2007 3216 2008
rect 3166 2003 3172 2004
rect 3210 2003 3211 2007
rect 3215 2003 3216 2007
rect 3280 2003 3282 2013
rect 3308 2008 3310 2086
rect 3344 2079 3346 2103
rect 3343 2078 3347 2079
rect 3343 2073 3347 2074
rect 3388 2048 3390 2166
rect 3512 2163 3514 2177
rect 3511 2162 3515 2163
rect 3511 2157 3515 2158
rect 3512 2147 3514 2157
rect 3564 2156 3566 2198
rect 3572 2172 3574 2362
rect 3590 2356 3596 2357
rect 3590 2352 3591 2356
rect 3595 2352 3596 2356
rect 3590 2351 3596 2352
rect 3592 2319 3594 2351
rect 3591 2318 3595 2319
rect 3591 2313 3595 2314
rect 3592 2285 3594 2313
rect 3590 2284 3596 2285
rect 3590 2280 3591 2284
rect 3595 2280 3596 2284
rect 3590 2279 3596 2280
rect 3590 2267 3596 2268
rect 3590 2263 3591 2267
rect 3595 2263 3596 2267
rect 3590 2262 3596 2263
rect 3592 2243 3594 2262
rect 3591 2242 3595 2243
rect 3591 2237 3595 2238
rect 3592 2218 3594 2237
rect 3590 2217 3596 2218
rect 3590 2213 3591 2217
rect 3595 2213 3596 2217
rect 3590 2212 3596 2213
rect 3590 2200 3596 2201
rect 3590 2196 3591 2200
rect 3595 2196 3596 2200
rect 3590 2195 3596 2196
rect 3570 2171 3576 2172
rect 3570 2167 3571 2171
rect 3575 2167 3576 2171
rect 3570 2166 3576 2167
rect 3592 2163 3594 2195
rect 3591 2162 3595 2163
rect 3591 2157 3595 2158
rect 3562 2155 3568 2156
rect 3562 2151 3563 2155
rect 3567 2151 3568 2155
rect 3562 2150 3568 2151
rect 3510 2146 3516 2147
rect 3510 2142 3511 2146
rect 3515 2142 3516 2146
rect 3510 2141 3516 2142
rect 3592 2129 3594 2157
rect 3590 2128 3596 2129
rect 3590 2124 3591 2128
rect 3595 2124 3596 2128
rect 3590 2123 3596 2124
rect 3534 2119 3540 2120
rect 3534 2115 3535 2119
rect 3539 2115 3540 2119
rect 3534 2114 3540 2115
rect 3502 2108 3508 2109
rect 3502 2104 3503 2108
rect 3507 2104 3508 2108
rect 3502 2103 3508 2104
rect 3504 2079 3506 2103
rect 3399 2078 3403 2079
rect 3399 2073 3403 2074
rect 3503 2078 3507 2079
rect 3503 2073 3507 2074
rect 3400 2057 3402 2073
rect 3504 2057 3506 2073
rect 3398 2056 3404 2057
rect 3398 2052 3399 2056
rect 3403 2052 3404 2056
rect 3398 2051 3404 2052
rect 3502 2056 3508 2057
rect 3502 2052 3503 2056
rect 3507 2052 3508 2056
rect 3502 2051 3508 2052
rect 3386 2047 3392 2048
rect 3386 2043 3387 2047
rect 3391 2043 3392 2047
rect 3386 2042 3392 2043
rect 3406 2018 3412 2019
rect 3406 2014 3407 2018
rect 3411 2014 3412 2018
rect 3406 2013 3412 2014
rect 3510 2018 3516 2019
rect 3510 2014 3511 2018
rect 3515 2014 3516 2018
rect 3510 2013 3516 2014
rect 3306 2007 3312 2008
rect 3306 2003 3307 2007
rect 3311 2003 3312 2007
rect 3408 2003 3410 2013
rect 3450 2007 3456 2008
rect 3450 2003 3451 2007
rect 3455 2003 3456 2007
rect 3512 2003 3514 2013
rect 3536 2008 3538 2114
rect 3590 2111 3596 2112
rect 3590 2107 3591 2111
rect 3595 2107 3596 2111
rect 3590 2106 3596 2107
rect 3592 2079 3594 2106
rect 3591 2078 3595 2079
rect 3591 2073 3595 2074
rect 3592 2054 3594 2073
rect 3590 2053 3596 2054
rect 3590 2049 3591 2053
rect 3595 2049 3596 2053
rect 3590 2048 3596 2049
rect 3562 2039 3568 2040
rect 3562 2035 3563 2039
rect 3567 2035 3568 2039
rect 3562 2034 3568 2035
rect 3590 2036 3596 2037
rect 3534 2007 3540 2008
rect 3534 2003 3535 2007
rect 3539 2003 3540 2007
rect 3119 2002 3123 2003
rect 3119 1997 3123 1998
rect 3151 2002 3155 2003
rect 3166 1999 3167 2003
rect 3171 2001 3182 2003
rect 3210 2002 3216 2003
rect 3279 2002 3283 2003
rect 3306 2002 3312 2003
rect 3327 2002 3331 2003
rect 3171 1999 3172 2001
rect 3166 1998 3172 1999
rect 3151 1997 3155 1998
rect 2926 1995 2932 1996
rect 2926 1991 2927 1995
rect 2931 1991 2932 1995
rect 2926 1990 2932 1991
rect 3078 1995 3084 1996
rect 3078 1991 3079 1995
rect 3083 1991 3084 1995
rect 3078 1990 3084 1991
rect 2918 1986 2924 1987
rect 2918 1982 2919 1986
rect 2923 1982 2924 1986
rect 2918 1981 2924 1982
rect 2928 1960 2930 1990
rect 3120 1987 3122 1997
rect 3170 1995 3176 1996
rect 3170 1991 3171 1995
rect 3175 1991 3176 1995
rect 3170 1990 3176 1991
rect 3118 1986 3124 1987
rect 3118 1982 3119 1986
rect 3123 1982 3124 1986
rect 3118 1981 3124 1982
rect 3172 1960 3174 1990
rect 3180 1960 3182 2001
rect 3279 1997 3283 1998
rect 3327 1997 3331 1998
rect 3407 2002 3411 2003
rect 3450 2002 3456 2003
rect 3511 2002 3515 2003
rect 3534 2002 3540 2003
rect 3407 1997 3411 1998
rect 3328 1987 3330 1997
rect 3326 1986 3332 1987
rect 3326 1982 3327 1986
rect 3331 1982 3332 1986
rect 3326 1981 3332 1982
rect 2590 1959 2596 1960
rect 2590 1955 2591 1959
rect 2595 1955 2596 1959
rect 2590 1954 2596 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2926 1959 2932 1960
rect 2926 1955 2927 1959
rect 2931 1955 2932 1959
rect 2926 1954 2932 1955
rect 3170 1959 3176 1960
rect 3170 1955 3171 1959
rect 3175 1955 3176 1959
rect 3170 1954 3176 1955
rect 3178 1959 3184 1960
rect 3178 1955 3179 1959
rect 3183 1955 3184 1959
rect 3178 1954 3184 1955
rect 2310 1948 2316 1949
rect 2310 1944 2311 1948
rect 2315 1944 2316 1948
rect 2310 1943 2316 1944
rect 2438 1948 2444 1949
rect 2438 1944 2439 1948
rect 2443 1944 2444 1948
rect 2438 1943 2444 1944
rect 2574 1948 2580 1949
rect 2574 1944 2575 1948
rect 2579 1944 2580 1948
rect 2574 1943 2580 1944
rect 2734 1948 2740 1949
rect 2734 1944 2735 1948
rect 2739 1944 2740 1948
rect 2734 1943 2740 1944
rect 2910 1948 2916 1949
rect 2910 1944 2911 1948
rect 2915 1944 2916 1948
rect 2910 1943 2916 1944
rect 3110 1948 3116 1949
rect 3110 1944 3111 1948
rect 3115 1944 3116 1948
rect 3110 1943 3116 1944
rect 3318 1948 3324 1949
rect 3318 1944 3319 1948
rect 3323 1944 3324 1948
rect 3318 1943 3324 1944
rect 2302 1931 2308 1932
rect 2302 1927 2303 1931
rect 2307 1927 2308 1931
rect 2302 1926 2308 1927
rect 2239 1918 2243 1919
rect 2239 1913 2243 1914
rect 2240 1897 2242 1913
rect 2238 1896 2244 1897
rect 2238 1892 2239 1896
rect 2243 1892 2244 1896
rect 2238 1891 2244 1892
rect 2130 1887 2136 1888
rect 2130 1883 2131 1887
rect 2135 1883 2136 1887
rect 2130 1882 2136 1883
rect 2222 1887 2228 1888
rect 2222 1883 2223 1887
rect 2227 1883 2228 1887
rect 2222 1882 2228 1883
rect 1830 1880 1836 1881
rect 1830 1876 1831 1880
rect 1835 1876 1836 1880
rect 1830 1875 1836 1876
rect 1870 1876 1876 1877
rect 1726 1851 1732 1852
rect 1726 1847 1727 1851
rect 1731 1847 1732 1851
rect 1726 1846 1732 1847
rect 1832 1843 1834 1875
rect 1870 1872 1871 1876
rect 1875 1872 1876 1876
rect 1870 1871 1876 1872
rect 1311 1842 1315 1843
rect 1311 1837 1315 1838
rect 1351 1842 1355 1843
rect 1351 1837 1355 1838
rect 1463 1842 1467 1843
rect 1463 1837 1467 1838
rect 1511 1842 1515 1843
rect 1511 1837 1515 1838
rect 1615 1842 1619 1843
rect 1615 1837 1619 1838
rect 1679 1842 1683 1843
rect 1679 1837 1683 1838
rect 1831 1842 1835 1843
rect 1831 1837 1835 1838
rect 1226 1835 1232 1836
rect 1226 1831 1227 1835
rect 1231 1831 1232 1835
rect 1226 1830 1232 1831
rect 1242 1835 1248 1836
rect 1242 1831 1243 1835
rect 1247 1831 1248 1835
rect 1242 1830 1248 1831
rect 1190 1826 1196 1827
rect 1190 1822 1191 1826
rect 1195 1822 1196 1826
rect 1190 1821 1196 1822
rect 1244 1800 1246 1830
rect 1352 1827 1354 1837
rect 1402 1835 1408 1836
rect 1402 1831 1403 1835
rect 1407 1831 1408 1835
rect 1402 1830 1408 1831
rect 1350 1826 1356 1827
rect 1350 1822 1351 1826
rect 1355 1822 1356 1826
rect 1350 1821 1356 1822
rect 1404 1800 1406 1830
rect 1512 1827 1514 1837
rect 1562 1835 1568 1836
rect 1562 1831 1563 1835
rect 1567 1831 1568 1835
rect 1562 1830 1568 1831
rect 1510 1826 1516 1827
rect 1510 1822 1511 1826
rect 1515 1822 1516 1826
rect 1510 1821 1516 1822
rect 1564 1800 1566 1830
rect 1680 1827 1682 1837
rect 1678 1826 1684 1827
rect 1678 1822 1679 1826
rect 1683 1822 1684 1826
rect 1678 1821 1684 1822
rect 1832 1809 1834 1837
rect 1872 1827 1874 1871
rect 2070 1858 2076 1859
rect 2070 1854 2071 1858
rect 2075 1854 2076 1858
rect 2070 1853 2076 1854
rect 2072 1827 2074 1853
rect 2132 1848 2134 1882
rect 2158 1858 2164 1859
rect 2158 1854 2159 1858
rect 2163 1854 2164 1858
rect 2158 1853 2164 1854
rect 2246 1858 2252 1859
rect 2246 1854 2247 1858
rect 2251 1854 2252 1858
rect 2246 1853 2252 1854
rect 2094 1847 2100 1848
rect 2094 1843 2095 1847
rect 2099 1843 2100 1847
rect 2130 1847 2136 1848
rect 2130 1843 2131 1847
rect 2135 1843 2136 1847
rect 2094 1842 2106 1843
rect 2130 1842 2136 1843
rect 2096 1841 2106 1842
rect 1871 1826 1875 1827
rect 1871 1821 1875 1822
rect 2071 1826 2075 1827
rect 2071 1821 2075 1822
rect 2095 1826 2099 1827
rect 2095 1821 2099 1822
rect 1830 1808 1836 1809
rect 1830 1804 1831 1808
rect 1835 1804 1836 1808
rect 1830 1803 1836 1804
rect 1242 1799 1248 1800
rect 1242 1795 1243 1799
rect 1247 1795 1248 1799
rect 1242 1794 1248 1795
rect 1402 1799 1408 1800
rect 1402 1795 1403 1799
rect 1407 1795 1408 1799
rect 1402 1794 1408 1795
rect 1562 1799 1568 1800
rect 1562 1795 1563 1799
rect 1567 1795 1568 1799
rect 1562 1794 1568 1795
rect 1872 1793 1874 1821
rect 2096 1811 2098 1821
rect 2094 1810 2100 1811
rect 2094 1806 2095 1810
rect 2099 1806 2100 1810
rect 2094 1805 2100 1806
rect 1870 1792 1876 1793
rect 1830 1791 1836 1792
rect 1182 1788 1188 1789
rect 1182 1784 1183 1788
rect 1187 1784 1188 1788
rect 1182 1783 1188 1784
rect 1342 1788 1348 1789
rect 1342 1784 1343 1788
rect 1347 1784 1348 1788
rect 1342 1783 1348 1784
rect 1502 1788 1508 1789
rect 1502 1784 1503 1788
rect 1507 1784 1508 1788
rect 1502 1783 1508 1784
rect 1670 1788 1676 1789
rect 1670 1784 1671 1788
rect 1675 1784 1676 1788
rect 1830 1787 1831 1791
rect 1835 1787 1836 1791
rect 1870 1788 1871 1792
rect 1875 1788 1876 1792
rect 1870 1787 1876 1788
rect 1830 1786 1836 1787
rect 1670 1783 1676 1784
rect 1184 1759 1186 1783
rect 1344 1759 1346 1783
rect 1354 1771 1360 1772
rect 1354 1767 1355 1771
rect 1359 1767 1360 1771
rect 1354 1766 1360 1767
rect 1167 1758 1171 1759
rect 1167 1753 1171 1754
rect 1183 1758 1187 1759
rect 1183 1753 1187 1754
rect 1319 1758 1323 1759
rect 1319 1753 1323 1754
rect 1343 1758 1347 1759
rect 1343 1753 1347 1754
rect 1168 1737 1170 1753
rect 1320 1737 1322 1753
rect 1166 1736 1172 1737
rect 1166 1732 1167 1736
rect 1171 1732 1172 1736
rect 1166 1731 1172 1732
rect 1318 1736 1324 1737
rect 1318 1732 1319 1736
rect 1323 1732 1324 1736
rect 1318 1731 1324 1732
rect 202 1727 208 1728
rect 202 1723 203 1727
rect 207 1723 208 1727
rect 202 1722 208 1723
rect 282 1727 288 1728
rect 282 1723 283 1727
rect 287 1723 288 1727
rect 282 1722 288 1723
rect 486 1727 492 1728
rect 486 1723 487 1727
rect 491 1723 492 1727
rect 486 1722 492 1723
rect 562 1727 568 1728
rect 562 1723 563 1727
rect 567 1723 568 1727
rect 562 1722 568 1723
rect 730 1727 736 1728
rect 730 1723 731 1727
rect 735 1723 736 1727
rect 730 1722 736 1723
rect 1090 1727 1096 1728
rect 1090 1723 1091 1727
rect 1095 1723 1096 1727
rect 1090 1722 1096 1723
rect 1102 1727 1108 1728
rect 1102 1723 1103 1727
rect 1107 1723 1108 1727
rect 1102 1722 1108 1723
rect 204 1688 206 1722
rect 222 1698 228 1699
rect 222 1694 223 1698
rect 227 1694 228 1698
rect 222 1693 228 1694
rect 166 1687 172 1688
rect 166 1683 167 1687
rect 171 1683 172 1687
rect 166 1682 172 1683
rect 202 1687 208 1688
rect 202 1683 203 1687
rect 207 1683 208 1687
rect 202 1682 208 1683
rect 224 1679 226 1693
rect 284 1688 286 1722
rect 350 1698 356 1699
rect 350 1694 351 1698
rect 355 1694 356 1698
rect 350 1693 356 1694
rect 502 1698 508 1699
rect 502 1694 503 1698
rect 507 1694 508 1698
rect 502 1693 508 1694
rect 282 1687 288 1688
rect 282 1683 283 1687
rect 287 1683 288 1687
rect 282 1682 288 1683
rect 352 1679 354 1693
rect 504 1679 506 1693
rect 564 1688 566 1722
rect 670 1698 676 1699
rect 670 1694 671 1698
rect 675 1694 676 1698
rect 670 1693 676 1694
rect 562 1687 568 1688
rect 562 1683 563 1687
rect 567 1683 568 1687
rect 562 1682 568 1683
rect 672 1679 674 1693
rect 732 1688 734 1722
rect 846 1698 852 1699
rect 846 1694 847 1698
rect 851 1694 852 1698
rect 846 1693 852 1694
rect 1014 1698 1020 1699
rect 1014 1694 1015 1698
rect 1019 1694 1020 1698
rect 1014 1693 1020 1694
rect 730 1687 736 1688
rect 730 1683 731 1687
rect 735 1683 736 1687
rect 730 1682 736 1683
rect 814 1687 820 1688
rect 814 1683 815 1687
rect 819 1683 820 1687
rect 814 1682 820 1683
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 143 1678 147 1679
rect 143 1673 147 1674
rect 223 1678 227 1679
rect 223 1673 227 1674
rect 295 1678 299 1679
rect 295 1673 299 1674
rect 351 1678 355 1679
rect 351 1673 355 1674
rect 479 1678 483 1679
rect 479 1673 483 1674
rect 503 1678 507 1679
rect 503 1673 507 1674
rect 671 1678 675 1679
rect 671 1673 675 1674
rect 112 1645 114 1673
rect 144 1663 146 1673
rect 296 1663 298 1673
rect 302 1671 308 1672
rect 302 1667 303 1671
rect 307 1667 308 1671
rect 302 1666 308 1667
rect 142 1662 148 1663
rect 142 1658 143 1662
rect 147 1658 148 1662
rect 142 1657 148 1658
rect 294 1662 300 1663
rect 294 1658 295 1662
rect 299 1658 300 1662
rect 294 1657 300 1658
rect 110 1644 116 1645
rect 110 1640 111 1644
rect 115 1640 116 1644
rect 110 1639 116 1640
rect 304 1636 306 1666
rect 480 1663 482 1673
rect 530 1671 536 1672
rect 530 1667 531 1671
rect 535 1667 536 1671
rect 530 1666 536 1667
rect 478 1662 484 1663
rect 478 1658 479 1662
rect 483 1658 484 1662
rect 478 1657 484 1658
rect 532 1636 534 1666
rect 672 1663 674 1673
rect 670 1662 676 1663
rect 670 1658 671 1662
rect 675 1658 676 1662
rect 670 1657 676 1658
rect 816 1636 818 1682
rect 848 1679 850 1693
rect 862 1679 868 1680
rect 1016 1679 1018 1693
rect 1092 1688 1094 1722
rect 1174 1698 1180 1699
rect 1174 1694 1175 1698
rect 1179 1694 1180 1698
rect 1174 1693 1180 1694
rect 1326 1698 1332 1699
rect 1326 1694 1327 1698
rect 1331 1694 1332 1698
rect 1326 1693 1332 1694
rect 1038 1687 1044 1688
rect 1038 1683 1039 1687
rect 1043 1683 1044 1687
rect 1038 1682 1044 1683
rect 1090 1687 1096 1688
rect 1090 1683 1091 1687
rect 1095 1683 1096 1687
rect 1090 1682 1096 1683
rect 847 1678 851 1679
rect 847 1673 851 1674
rect 855 1678 859 1679
rect 862 1675 863 1679
rect 867 1675 868 1679
rect 862 1674 868 1675
rect 1015 1678 1019 1679
rect 855 1673 859 1674
rect 856 1663 858 1673
rect 854 1662 860 1663
rect 854 1658 855 1662
rect 859 1658 860 1662
rect 854 1657 860 1658
rect 864 1636 866 1674
rect 1015 1673 1019 1674
rect 1031 1678 1035 1679
rect 1031 1673 1035 1674
rect 914 1671 920 1672
rect 914 1667 915 1671
rect 919 1667 920 1671
rect 914 1666 920 1667
rect 190 1635 196 1636
rect 190 1631 191 1635
rect 195 1631 196 1635
rect 190 1630 196 1631
rect 302 1635 308 1636
rect 302 1631 303 1635
rect 307 1631 308 1635
rect 302 1630 308 1631
rect 530 1635 536 1636
rect 530 1631 531 1635
rect 535 1631 536 1635
rect 530 1630 536 1631
rect 814 1635 820 1636
rect 814 1631 815 1635
rect 819 1631 820 1635
rect 814 1630 820 1631
rect 862 1635 868 1636
rect 862 1631 863 1635
rect 867 1631 868 1635
rect 862 1630 868 1631
rect 110 1627 116 1628
rect 110 1623 111 1627
rect 115 1623 116 1627
rect 110 1622 116 1623
rect 134 1624 140 1625
rect 112 1603 114 1622
rect 134 1620 135 1624
rect 139 1620 140 1624
rect 134 1619 140 1620
rect 136 1603 138 1619
rect 111 1602 115 1603
rect 111 1597 115 1598
rect 135 1602 139 1603
rect 135 1597 139 1598
rect 159 1602 163 1603
rect 159 1597 163 1598
rect 112 1578 114 1597
rect 160 1581 162 1597
rect 158 1580 164 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 158 1576 159 1580
rect 163 1576 164 1580
rect 158 1575 164 1576
rect 110 1572 116 1573
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 110 1555 116 1556
rect 112 1523 114 1555
rect 166 1542 172 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 168 1523 170 1537
rect 192 1532 194 1630
rect 286 1624 292 1625
rect 286 1620 287 1624
rect 291 1620 292 1624
rect 286 1619 292 1620
rect 470 1624 476 1625
rect 470 1620 471 1624
rect 475 1620 476 1624
rect 470 1619 476 1620
rect 662 1624 668 1625
rect 662 1620 663 1624
rect 667 1620 668 1624
rect 662 1619 668 1620
rect 846 1624 852 1625
rect 846 1620 847 1624
rect 851 1620 852 1624
rect 846 1619 852 1620
rect 288 1603 290 1619
rect 472 1603 474 1619
rect 664 1603 666 1619
rect 848 1603 850 1619
rect 287 1602 291 1603
rect 287 1597 291 1598
rect 423 1602 427 1603
rect 423 1597 427 1598
rect 471 1602 475 1603
rect 471 1597 475 1598
rect 567 1602 571 1603
rect 567 1597 571 1598
rect 663 1602 667 1603
rect 663 1597 667 1598
rect 711 1602 715 1603
rect 711 1597 715 1598
rect 847 1602 851 1603
rect 847 1597 851 1598
rect 288 1581 290 1597
rect 424 1581 426 1597
rect 568 1581 570 1597
rect 712 1581 714 1597
rect 848 1581 850 1597
rect 286 1580 292 1581
rect 286 1576 287 1580
rect 291 1576 292 1580
rect 286 1575 292 1576
rect 422 1580 428 1581
rect 422 1576 423 1580
rect 427 1576 428 1580
rect 422 1575 428 1576
rect 566 1580 572 1581
rect 566 1576 567 1580
rect 571 1576 572 1580
rect 566 1575 572 1576
rect 710 1580 716 1581
rect 710 1576 711 1580
rect 715 1576 716 1580
rect 710 1575 716 1576
rect 846 1580 852 1581
rect 846 1576 847 1580
rect 851 1576 852 1580
rect 846 1575 852 1576
rect 916 1572 918 1666
rect 1032 1663 1034 1673
rect 1030 1662 1036 1663
rect 1030 1658 1031 1662
rect 1035 1658 1036 1662
rect 1030 1657 1036 1658
rect 1040 1636 1042 1682
rect 1176 1679 1178 1693
rect 1328 1679 1330 1693
rect 1356 1688 1358 1766
rect 1504 1759 1506 1783
rect 1672 1759 1674 1783
rect 1832 1759 1834 1786
rect 2104 1784 2106 1841
rect 2160 1827 2162 1853
rect 2248 1827 2250 1853
rect 2304 1848 2306 1926
rect 2312 1919 2314 1943
rect 2378 1931 2384 1932
rect 2378 1927 2379 1931
rect 2383 1927 2384 1931
rect 2378 1926 2384 1927
rect 2311 1918 2315 1919
rect 2311 1913 2315 1914
rect 2319 1918 2323 1919
rect 2319 1913 2323 1914
rect 2320 1897 2322 1913
rect 2318 1896 2324 1897
rect 2318 1892 2319 1896
rect 2323 1892 2324 1896
rect 2318 1891 2324 1892
rect 2326 1858 2332 1859
rect 2326 1854 2327 1858
rect 2331 1854 2332 1858
rect 2326 1853 2332 1854
rect 2302 1847 2308 1848
rect 2302 1843 2303 1847
rect 2307 1843 2308 1847
rect 2302 1842 2308 1843
rect 2328 1827 2330 1853
rect 2380 1848 2382 1926
rect 2440 1919 2442 1943
rect 2576 1919 2578 1943
rect 2736 1919 2738 1943
rect 2912 1919 2914 1943
rect 3112 1919 3114 1943
rect 3320 1919 3322 1943
rect 2399 1918 2403 1919
rect 2399 1913 2403 1914
rect 2439 1918 2443 1919
rect 2439 1913 2443 1914
rect 2487 1918 2491 1919
rect 2487 1913 2491 1914
rect 2575 1918 2579 1919
rect 2575 1913 2579 1914
rect 2663 1918 2667 1919
rect 2663 1913 2667 1914
rect 2735 1918 2739 1919
rect 2735 1913 2739 1914
rect 2759 1918 2763 1919
rect 2759 1913 2763 1914
rect 2871 1918 2875 1919
rect 2871 1913 2875 1914
rect 2911 1918 2915 1919
rect 2911 1913 2915 1914
rect 2991 1918 2995 1919
rect 2991 1913 2995 1914
rect 3111 1918 3115 1919
rect 3111 1913 3115 1914
rect 3119 1918 3123 1919
rect 3119 1913 3123 1914
rect 3247 1918 3251 1919
rect 3247 1913 3251 1914
rect 3319 1918 3323 1919
rect 3319 1913 3323 1914
rect 3383 1918 3387 1919
rect 3383 1913 3387 1914
rect 2400 1897 2402 1913
rect 2488 1897 2490 1913
rect 2576 1897 2578 1913
rect 2664 1897 2666 1913
rect 2760 1897 2762 1913
rect 2872 1897 2874 1913
rect 2992 1897 2994 1913
rect 3120 1897 3122 1913
rect 3248 1897 3250 1913
rect 3384 1897 3386 1913
rect 2398 1896 2404 1897
rect 2398 1892 2399 1896
rect 2403 1892 2404 1896
rect 2398 1891 2404 1892
rect 2486 1896 2492 1897
rect 2486 1892 2487 1896
rect 2491 1892 2492 1896
rect 2486 1891 2492 1892
rect 2574 1896 2580 1897
rect 2574 1892 2575 1896
rect 2579 1892 2580 1896
rect 2574 1891 2580 1892
rect 2662 1896 2668 1897
rect 2662 1892 2663 1896
rect 2667 1892 2668 1896
rect 2662 1891 2668 1892
rect 2758 1896 2764 1897
rect 2758 1892 2759 1896
rect 2763 1892 2764 1896
rect 2758 1891 2764 1892
rect 2870 1896 2876 1897
rect 2870 1892 2871 1896
rect 2875 1892 2876 1896
rect 2870 1891 2876 1892
rect 2990 1896 2996 1897
rect 2990 1892 2991 1896
rect 2995 1892 2996 1896
rect 2990 1891 2996 1892
rect 3118 1896 3124 1897
rect 3118 1892 3119 1896
rect 3123 1892 3124 1896
rect 3118 1891 3124 1892
rect 3246 1896 3252 1897
rect 3246 1892 3247 1896
rect 3251 1892 3252 1896
rect 3246 1891 3252 1892
rect 3382 1896 3388 1897
rect 3382 1892 3383 1896
rect 3387 1892 3388 1896
rect 3382 1891 3388 1892
rect 3452 1888 3454 2002
rect 3511 1997 3515 1998
rect 3512 1987 3514 1997
rect 3564 1996 3566 2034
rect 3590 2032 3591 2036
rect 3595 2032 3596 2036
rect 3590 2031 3596 2032
rect 3592 2003 3594 2031
rect 3591 2002 3595 2003
rect 3591 1997 3595 1998
rect 3562 1995 3568 1996
rect 3562 1991 3563 1995
rect 3567 1991 3568 1995
rect 3562 1990 3568 1991
rect 3510 1986 3516 1987
rect 3510 1982 3511 1986
rect 3515 1982 3516 1986
rect 3510 1981 3516 1982
rect 3592 1969 3594 1997
rect 3590 1968 3596 1969
rect 3590 1964 3591 1968
rect 3595 1964 3596 1968
rect 3590 1963 3596 1964
rect 3534 1959 3540 1960
rect 3534 1955 3535 1959
rect 3539 1955 3540 1959
rect 3534 1954 3540 1955
rect 3502 1948 3508 1949
rect 3502 1944 3503 1948
rect 3507 1944 3508 1948
rect 3502 1943 3508 1944
rect 3504 1919 3506 1943
rect 3503 1918 3507 1919
rect 3503 1913 3507 1914
rect 3504 1897 3506 1913
rect 3502 1896 3508 1897
rect 3502 1892 3503 1896
rect 3507 1892 3508 1896
rect 3502 1891 3508 1892
rect 2386 1887 2392 1888
rect 2386 1883 2387 1887
rect 2391 1883 2392 1887
rect 2386 1882 2392 1883
rect 2466 1887 2472 1888
rect 2466 1883 2467 1887
rect 2471 1883 2472 1887
rect 2466 1882 2472 1883
rect 2554 1887 2560 1888
rect 2554 1883 2555 1887
rect 2559 1883 2560 1887
rect 2554 1882 2560 1883
rect 2642 1887 2648 1888
rect 2642 1883 2643 1887
rect 2647 1883 2648 1887
rect 2642 1882 2648 1883
rect 2734 1887 2740 1888
rect 2734 1883 2735 1887
rect 2739 1883 2740 1887
rect 2734 1882 2740 1883
rect 2954 1887 2960 1888
rect 2954 1883 2955 1887
rect 2959 1883 2960 1887
rect 2954 1882 2960 1883
rect 3078 1887 3084 1888
rect 3078 1883 3079 1887
rect 3083 1883 3084 1887
rect 3078 1882 3084 1883
rect 3194 1887 3200 1888
rect 3194 1883 3195 1887
rect 3199 1883 3200 1887
rect 3194 1882 3200 1883
rect 3202 1887 3208 1888
rect 3202 1883 3203 1887
rect 3207 1883 3208 1887
rect 3202 1882 3208 1883
rect 3450 1887 3456 1888
rect 3450 1883 3451 1887
rect 3455 1883 3456 1887
rect 3450 1882 3456 1883
rect 3458 1887 3464 1888
rect 3458 1883 3459 1887
rect 3463 1883 3464 1887
rect 3458 1882 3464 1883
rect 2388 1848 2390 1882
rect 2458 1879 2464 1880
rect 2458 1875 2459 1879
rect 2463 1875 2464 1879
rect 2458 1874 2464 1875
rect 2406 1858 2412 1859
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2378 1847 2384 1848
rect 2378 1843 2379 1847
rect 2383 1843 2384 1847
rect 2378 1842 2384 1843
rect 2386 1847 2392 1848
rect 2386 1843 2387 1847
rect 2391 1843 2392 1847
rect 2386 1842 2392 1843
rect 2408 1827 2410 1853
rect 2159 1826 2163 1827
rect 2159 1821 2163 1822
rect 2239 1826 2243 1827
rect 2239 1821 2243 1822
rect 2247 1826 2251 1827
rect 2247 1821 2251 1822
rect 2327 1826 2331 1827
rect 2327 1821 2331 1822
rect 2399 1826 2403 1827
rect 2399 1821 2403 1822
rect 2407 1826 2411 1827
rect 2407 1821 2411 1822
rect 2240 1811 2242 1821
rect 2334 1819 2340 1820
rect 2334 1815 2335 1819
rect 2339 1815 2340 1819
rect 2334 1814 2340 1815
rect 2238 1810 2244 1811
rect 2238 1806 2239 1810
rect 2243 1806 2244 1810
rect 2238 1805 2244 1806
rect 2336 1784 2338 1814
rect 2400 1811 2402 1821
rect 2460 1820 2462 1874
rect 2468 1848 2470 1882
rect 2494 1858 2500 1859
rect 2494 1854 2495 1858
rect 2499 1854 2500 1858
rect 2494 1853 2500 1854
rect 2466 1847 2472 1848
rect 2466 1843 2467 1847
rect 2471 1843 2472 1847
rect 2466 1842 2472 1843
rect 2496 1827 2498 1853
rect 2556 1848 2558 1882
rect 2582 1858 2588 1859
rect 2582 1854 2583 1858
rect 2587 1854 2588 1858
rect 2582 1853 2588 1854
rect 2554 1847 2560 1848
rect 2554 1843 2555 1847
rect 2559 1843 2560 1847
rect 2554 1842 2560 1843
rect 2584 1827 2586 1853
rect 2644 1848 2646 1882
rect 2670 1858 2676 1859
rect 2670 1854 2671 1858
rect 2675 1854 2676 1858
rect 2670 1853 2676 1854
rect 2642 1847 2648 1848
rect 2642 1843 2643 1847
rect 2647 1843 2648 1847
rect 2642 1842 2648 1843
rect 2672 1827 2674 1853
rect 2736 1848 2738 1882
rect 2766 1858 2772 1859
rect 2766 1854 2767 1858
rect 2771 1854 2772 1858
rect 2766 1853 2772 1854
rect 2878 1858 2884 1859
rect 2878 1854 2879 1858
rect 2883 1854 2884 1858
rect 2878 1853 2884 1854
rect 2734 1847 2740 1848
rect 2734 1843 2735 1847
rect 2739 1843 2740 1847
rect 2734 1842 2740 1843
rect 2768 1827 2770 1853
rect 2880 1827 2882 1853
rect 2956 1848 2958 1882
rect 2998 1858 3004 1859
rect 2998 1854 2999 1858
rect 3003 1854 3004 1858
rect 2998 1853 3004 1854
rect 2954 1847 2960 1848
rect 2954 1843 2955 1847
rect 2959 1843 2960 1847
rect 2954 1842 2960 1843
rect 3000 1827 3002 1853
rect 3080 1848 3082 1882
rect 3126 1858 3132 1859
rect 3126 1854 3127 1858
rect 3131 1854 3132 1858
rect 3126 1853 3132 1854
rect 3078 1847 3084 1848
rect 3078 1843 3079 1847
rect 3083 1843 3084 1847
rect 3078 1842 3084 1843
rect 3128 1827 3130 1853
rect 3196 1848 3198 1882
rect 3194 1847 3200 1848
rect 3194 1843 3195 1847
rect 3199 1843 3200 1847
rect 3194 1842 3200 1843
rect 2495 1826 2499 1827
rect 2495 1821 2499 1822
rect 2559 1826 2563 1827
rect 2559 1821 2563 1822
rect 2583 1826 2587 1827
rect 2583 1821 2587 1822
rect 2671 1826 2675 1827
rect 2671 1821 2675 1822
rect 2719 1826 2723 1827
rect 2719 1821 2723 1822
rect 2767 1826 2771 1827
rect 2767 1821 2771 1822
rect 2879 1826 2883 1827
rect 2879 1821 2883 1822
rect 2999 1826 3003 1827
rect 2999 1821 3003 1822
rect 3031 1826 3035 1827
rect 3031 1821 3035 1822
rect 3127 1826 3131 1827
rect 3127 1821 3131 1822
rect 3175 1826 3179 1827
rect 3175 1821 3179 1822
rect 2450 1819 2456 1820
rect 2450 1815 2451 1819
rect 2455 1815 2456 1819
rect 2450 1814 2456 1815
rect 2458 1819 2464 1820
rect 2458 1815 2459 1819
rect 2463 1815 2464 1819
rect 2458 1814 2464 1815
rect 2398 1810 2404 1811
rect 2398 1806 2399 1810
rect 2403 1806 2404 1810
rect 2398 1805 2404 1806
rect 2102 1783 2108 1784
rect 2102 1779 2103 1783
rect 2107 1779 2108 1783
rect 2102 1778 2108 1779
rect 2334 1783 2340 1784
rect 2334 1779 2335 1783
rect 2339 1779 2340 1783
rect 2334 1778 2340 1779
rect 1870 1775 1876 1776
rect 1870 1771 1871 1775
rect 1875 1771 1876 1775
rect 1870 1770 1876 1771
rect 2086 1772 2092 1773
rect 1463 1758 1467 1759
rect 1463 1753 1467 1754
rect 1503 1758 1507 1759
rect 1503 1753 1507 1754
rect 1607 1758 1611 1759
rect 1607 1753 1611 1754
rect 1671 1758 1675 1759
rect 1671 1753 1675 1754
rect 1743 1758 1747 1759
rect 1743 1753 1747 1754
rect 1831 1758 1835 1759
rect 1831 1753 1835 1754
rect 1464 1737 1466 1753
rect 1608 1737 1610 1753
rect 1744 1737 1746 1753
rect 1462 1736 1468 1737
rect 1462 1732 1463 1736
rect 1467 1732 1468 1736
rect 1462 1731 1468 1732
rect 1606 1736 1612 1737
rect 1606 1732 1607 1736
rect 1611 1732 1612 1736
rect 1606 1731 1612 1732
rect 1742 1736 1748 1737
rect 1742 1732 1743 1736
rect 1747 1732 1748 1736
rect 1832 1734 1834 1753
rect 1872 1747 1874 1770
rect 2086 1768 2087 1772
rect 2091 1768 2092 1772
rect 2086 1767 2092 1768
rect 2230 1772 2236 1773
rect 2230 1768 2231 1772
rect 2235 1768 2236 1772
rect 2230 1767 2236 1768
rect 2390 1772 2396 1773
rect 2390 1768 2391 1772
rect 2395 1768 2396 1772
rect 2390 1767 2396 1768
rect 2088 1747 2090 1767
rect 2232 1747 2234 1767
rect 2392 1747 2394 1767
rect 1871 1746 1875 1747
rect 1871 1741 1875 1742
rect 2087 1746 2091 1747
rect 2087 1741 2091 1742
rect 2103 1746 2107 1747
rect 2103 1741 2107 1742
rect 2231 1746 2235 1747
rect 2231 1741 2235 1742
rect 2239 1746 2243 1747
rect 2239 1741 2243 1742
rect 2383 1746 2387 1747
rect 2383 1741 2387 1742
rect 2391 1746 2395 1747
rect 2391 1741 2395 1742
rect 1742 1731 1748 1732
rect 1830 1733 1836 1734
rect 1830 1729 1831 1733
rect 1835 1729 1836 1733
rect 1830 1728 1836 1729
rect 1410 1727 1416 1728
rect 1410 1723 1411 1727
rect 1415 1723 1416 1727
rect 1410 1722 1416 1723
rect 1554 1727 1560 1728
rect 1554 1723 1555 1727
rect 1559 1723 1560 1727
rect 1554 1722 1560 1723
rect 1690 1727 1696 1728
rect 1690 1723 1691 1727
rect 1695 1723 1696 1727
rect 1690 1722 1696 1723
rect 1706 1727 1712 1728
rect 1706 1723 1707 1727
rect 1711 1723 1712 1727
rect 1706 1722 1712 1723
rect 1872 1722 1874 1741
rect 2104 1725 2106 1741
rect 2240 1725 2242 1741
rect 2384 1725 2386 1741
rect 2102 1724 2108 1725
rect 1412 1688 1414 1722
rect 1470 1698 1476 1699
rect 1470 1694 1471 1698
rect 1475 1694 1476 1698
rect 1470 1693 1476 1694
rect 1354 1687 1360 1688
rect 1354 1683 1355 1687
rect 1359 1683 1360 1687
rect 1354 1682 1360 1683
rect 1410 1687 1416 1688
rect 1410 1683 1411 1687
rect 1415 1683 1416 1687
rect 1410 1682 1416 1683
rect 1472 1679 1474 1693
rect 1556 1688 1558 1722
rect 1614 1698 1620 1699
rect 1614 1694 1615 1698
rect 1619 1694 1620 1698
rect 1614 1693 1620 1694
rect 1554 1687 1560 1688
rect 1554 1683 1555 1687
rect 1559 1683 1560 1687
rect 1554 1682 1560 1683
rect 1616 1679 1618 1693
rect 1692 1688 1694 1722
rect 1690 1687 1696 1688
rect 1690 1683 1691 1687
rect 1695 1683 1696 1687
rect 1690 1682 1696 1683
rect 1175 1678 1179 1679
rect 1175 1673 1179 1674
rect 1199 1678 1203 1679
rect 1199 1673 1203 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 1359 1678 1363 1679
rect 1359 1673 1363 1674
rect 1471 1678 1475 1679
rect 1471 1673 1475 1674
rect 1519 1678 1523 1679
rect 1519 1673 1523 1674
rect 1615 1678 1619 1679
rect 1615 1673 1619 1674
rect 1679 1678 1683 1679
rect 1679 1673 1683 1674
rect 1058 1671 1064 1672
rect 1058 1667 1059 1671
rect 1063 1667 1064 1671
rect 1058 1666 1064 1667
rect 1038 1635 1044 1636
rect 1038 1631 1039 1635
rect 1043 1631 1044 1635
rect 1038 1630 1044 1631
rect 1022 1624 1028 1625
rect 1022 1620 1023 1624
rect 1027 1620 1028 1624
rect 1022 1619 1028 1620
rect 1024 1603 1026 1619
rect 983 1602 987 1603
rect 983 1597 987 1598
rect 1023 1602 1027 1603
rect 1023 1597 1027 1598
rect 984 1581 986 1597
rect 982 1580 988 1581
rect 982 1576 983 1580
rect 987 1576 988 1580
rect 982 1575 988 1576
rect 1060 1572 1062 1666
rect 1200 1663 1202 1673
rect 1360 1663 1362 1673
rect 1366 1671 1372 1672
rect 1366 1667 1367 1671
rect 1371 1667 1372 1671
rect 1366 1666 1372 1667
rect 1198 1662 1204 1663
rect 1198 1658 1199 1662
rect 1203 1658 1204 1662
rect 1198 1657 1204 1658
rect 1358 1662 1364 1663
rect 1358 1658 1359 1662
rect 1363 1658 1364 1662
rect 1358 1657 1364 1658
rect 1368 1636 1370 1666
rect 1520 1663 1522 1673
rect 1526 1671 1532 1672
rect 1526 1667 1527 1671
rect 1531 1667 1532 1671
rect 1526 1666 1532 1667
rect 1518 1662 1524 1663
rect 1518 1658 1519 1662
rect 1523 1658 1524 1662
rect 1518 1657 1524 1658
rect 1528 1636 1530 1666
rect 1680 1663 1682 1673
rect 1708 1672 1710 1722
rect 1870 1721 1876 1722
rect 1870 1717 1871 1721
rect 1875 1717 1876 1721
rect 2102 1720 2103 1724
rect 2107 1720 2108 1724
rect 2102 1719 2108 1720
rect 2238 1724 2244 1725
rect 2238 1720 2239 1724
rect 2243 1720 2244 1724
rect 2238 1719 2244 1720
rect 2382 1724 2388 1725
rect 2382 1720 2383 1724
rect 2387 1720 2388 1724
rect 2382 1719 2388 1720
rect 1830 1716 1836 1717
rect 1870 1716 1876 1717
rect 2452 1716 2454 1814
rect 2560 1811 2562 1821
rect 2610 1819 2616 1820
rect 2610 1815 2611 1819
rect 2615 1815 2616 1819
rect 2610 1814 2616 1815
rect 2558 1810 2564 1811
rect 2558 1806 2559 1810
rect 2563 1806 2564 1810
rect 2558 1805 2564 1806
rect 2612 1784 2614 1814
rect 2720 1811 2722 1821
rect 2880 1811 2882 1821
rect 3032 1811 3034 1821
rect 3038 1819 3044 1820
rect 3038 1815 3039 1819
rect 3043 1815 3044 1819
rect 3038 1814 3044 1815
rect 3118 1819 3124 1820
rect 3118 1815 3119 1819
rect 3123 1815 3124 1819
rect 3118 1814 3124 1815
rect 2718 1810 2724 1811
rect 2718 1806 2719 1810
rect 2723 1806 2724 1810
rect 2718 1805 2724 1806
rect 2878 1810 2884 1811
rect 2878 1806 2879 1810
rect 2883 1806 2884 1810
rect 2878 1805 2884 1806
rect 3030 1810 3036 1811
rect 3030 1806 3031 1810
rect 3035 1806 3036 1810
rect 3030 1805 3036 1806
rect 3040 1784 3042 1814
rect 2610 1783 2616 1784
rect 2610 1779 2611 1783
rect 2615 1779 2616 1783
rect 2610 1778 2616 1779
rect 3038 1783 3044 1784
rect 3038 1779 3039 1783
rect 3043 1779 3044 1783
rect 3038 1778 3044 1779
rect 2550 1772 2556 1773
rect 2550 1768 2551 1772
rect 2555 1768 2556 1772
rect 2550 1767 2556 1768
rect 2710 1772 2716 1773
rect 2710 1768 2711 1772
rect 2715 1768 2716 1772
rect 2710 1767 2716 1768
rect 2870 1772 2876 1773
rect 2870 1768 2871 1772
rect 2875 1768 2876 1772
rect 2870 1767 2876 1768
rect 3022 1772 3028 1773
rect 3022 1768 3023 1772
rect 3027 1768 3028 1772
rect 3022 1767 3028 1768
rect 2552 1747 2554 1767
rect 2698 1755 2704 1756
rect 2698 1751 2699 1755
rect 2703 1751 2704 1755
rect 2698 1750 2704 1751
rect 2527 1746 2531 1747
rect 2527 1741 2531 1742
rect 2551 1746 2555 1747
rect 2551 1741 2555 1742
rect 2663 1746 2667 1747
rect 2663 1741 2667 1742
rect 2528 1725 2530 1741
rect 2664 1725 2666 1741
rect 2526 1724 2532 1725
rect 2526 1720 2527 1724
rect 2531 1720 2532 1724
rect 2526 1719 2532 1720
rect 2662 1724 2668 1725
rect 2662 1720 2663 1724
rect 2667 1720 2668 1724
rect 2662 1719 2668 1720
rect 1830 1712 1831 1716
rect 1835 1712 1836 1716
rect 1830 1711 1836 1712
rect 2186 1715 2192 1716
rect 2186 1711 2187 1715
rect 2191 1711 2192 1715
rect 1750 1698 1756 1699
rect 1750 1694 1751 1698
rect 1755 1694 1756 1698
rect 1750 1693 1756 1694
rect 1752 1679 1754 1693
rect 1832 1679 1834 1711
rect 2186 1710 2192 1711
rect 2330 1715 2336 1716
rect 2330 1711 2331 1715
rect 2335 1711 2336 1715
rect 2330 1710 2336 1711
rect 2450 1715 2456 1716
rect 2450 1711 2451 1715
rect 2455 1711 2456 1715
rect 2450 1710 2456 1711
rect 2594 1715 2600 1716
rect 2594 1711 2595 1715
rect 2599 1711 2600 1715
rect 2594 1710 2600 1711
rect 1870 1704 1876 1705
rect 1870 1700 1871 1704
rect 1875 1700 1876 1704
rect 1870 1699 1876 1700
rect 1751 1678 1755 1679
rect 1751 1673 1755 1674
rect 1831 1678 1835 1679
rect 1831 1673 1835 1674
rect 1686 1671 1692 1672
rect 1686 1667 1687 1671
rect 1691 1667 1692 1671
rect 1686 1666 1692 1667
rect 1706 1671 1712 1672
rect 1706 1667 1707 1671
rect 1711 1667 1712 1671
rect 1706 1666 1712 1667
rect 1678 1662 1684 1663
rect 1678 1658 1679 1662
rect 1683 1658 1684 1662
rect 1678 1657 1684 1658
rect 1688 1636 1690 1666
rect 1832 1645 1834 1673
rect 1872 1667 1874 1699
rect 2110 1686 2116 1687
rect 2110 1682 2111 1686
rect 2115 1682 2116 1686
rect 2110 1681 2116 1682
rect 2112 1667 2114 1681
rect 2188 1676 2190 1710
rect 2246 1686 2252 1687
rect 2246 1682 2247 1686
rect 2251 1682 2252 1686
rect 2246 1681 2252 1682
rect 2186 1675 2192 1676
rect 2186 1671 2187 1675
rect 2191 1671 2192 1675
rect 2186 1670 2192 1671
rect 2248 1667 2250 1681
rect 2332 1676 2334 1710
rect 2390 1686 2396 1687
rect 2390 1682 2391 1686
rect 2395 1682 2396 1686
rect 2390 1681 2396 1682
rect 2534 1686 2540 1687
rect 2534 1682 2535 1686
rect 2539 1682 2540 1686
rect 2534 1681 2540 1682
rect 2330 1675 2336 1676
rect 2330 1671 2331 1675
rect 2335 1671 2336 1675
rect 2330 1670 2336 1671
rect 2358 1667 2364 1668
rect 2392 1667 2394 1681
rect 2536 1667 2538 1681
rect 2596 1676 2598 1710
rect 2654 1707 2660 1708
rect 2654 1703 2655 1707
rect 2659 1703 2660 1707
rect 2654 1702 2660 1703
rect 2594 1675 2600 1676
rect 2594 1671 2595 1675
rect 2599 1671 2600 1675
rect 2594 1670 2600 1671
rect 1871 1666 1875 1667
rect 1871 1661 1875 1662
rect 1967 1666 1971 1667
rect 1967 1661 1971 1662
rect 2087 1666 2091 1667
rect 2087 1661 2091 1662
rect 2111 1666 2115 1667
rect 2111 1661 2115 1662
rect 2215 1666 2219 1667
rect 2215 1661 2219 1662
rect 2247 1666 2251 1667
rect 2247 1661 2251 1662
rect 2351 1666 2355 1667
rect 2358 1663 2359 1667
rect 2363 1663 2364 1667
rect 2358 1662 2364 1663
rect 2391 1666 2395 1667
rect 2351 1661 2355 1662
rect 1830 1644 1836 1645
rect 1830 1640 1831 1644
rect 1835 1640 1836 1644
rect 1830 1639 1836 1640
rect 1262 1635 1268 1636
rect 1262 1631 1263 1635
rect 1267 1631 1268 1635
rect 1262 1630 1268 1631
rect 1366 1635 1372 1636
rect 1366 1631 1367 1635
rect 1371 1631 1372 1635
rect 1366 1630 1372 1631
rect 1526 1635 1532 1636
rect 1526 1631 1527 1635
rect 1531 1631 1532 1635
rect 1526 1630 1532 1631
rect 1686 1635 1692 1636
rect 1686 1631 1687 1635
rect 1691 1631 1692 1635
rect 1872 1633 1874 1661
rect 1968 1651 1970 1661
rect 1974 1659 1980 1660
rect 1974 1655 1975 1659
rect 1979 1655 1980 1659
rect 1974 1654 1980 1655
rect 2018 1659 2024 1660
rect 2018 1655 2019 1659
rect 2023 1655 2024 1659
rect 2018 1654 2024 1655
rect 1966 1650 1972 1651
rect 1966 1646 1967 1650
rect 1971 1646 1972 1650
rect 1966 1645 1972 1646
rect 1686 1630 1692 1631
rect 1870 1632 1876 1633
rect 1190 1624 1196 1625
rect 1190 1620 1191 1624
rect 1195 1620 1196 1624
rect 1190 1619 1196 1620
rect 1192 1603 1194 1619
rect 1119 1602 1123 1603
rect 1119 1597 1123 1598
rect 1191 1602 1195 1603
rect 1191 1597 1195 1598
rect 1247 1602 1251 1603
rect 1247 1597 1251 1598
rect 1120 1581 1122 1597
rect 1248 1581 1250 1597
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1246 1580 1252 1581
rect 1246 1576 1247 1580
rect 1251 1576 1252 1580
rect 1246 1575 1252 1576
rect 230 1571 236 1572
rect 230 1567 231 1571
rect 235 1567 236 1571
rect 230 1566 236 1567
rect 258 1571 264 1572
rect 258 1567 259 1571
rect 263 1567 264 1571
rect 258 1566 264 1567
rect 534 1571 540 1572
rect 534 1567 535 1571
rect 539 1567 540 1571
rect 534 1566 540 1567
rect 658 1571 664 1572
rect 658 1567 659 1571
rect 663 1567 664 1571
rect 658 1566 664 1567
rect 802 1571 808 1572
rect 802 1567 803 1571
rect 807 1567 808 1571
rect 802 1566 808 1567
rect 914 1571 920 1572
rect 914 1567 915 1571
rect 919 1567 920 1571
rect 914 1566 920 1567
rect 1050 1571 1056 1572
rect 1050 1567 1051 1571
rect 1055 1567 1056 1571
rect 1050 1566 1056 1567
rect 1058 1571 1064 1572
rect 1058 1567 1059 1571
rect 1063 1567 1064 1571
rect 1058 1566 1064 1567
rect 232 1532 234 1566
rect 190 1531 196 1532
rect 190 1527 191 1531
rect 195 1527 196 1531
rect 190 1526 196 1527
rect 230 1531 236 1532
rect 230 1527 231 1531
rect 235 1527 236 1531
rect 230 1526 236 1527
rect 111 1522 115 1523
rect 111 1517 115 1518
rect 167 1522 171 1523
rect 167 1517 171 1518
rect 231 1522 235 1523
rect 231 1517 235 1518
rect 112 1489 114 1517
rect 232 1507 234 1517
rect 260 1516 262 1566
rect 294 1542 300 1543
rect 294 1538 295 1542
rect 299 1538 300 1542
rect 294 1537 300 1538
rect 430 1542 436 1543
rect 430 1538 431 1542
rect 435 1538 436 1542
rect 430 1537 436 1538
rect 296 1523 298 1537
rect 432 1523 434 1537
rect 536 1532 538 1566
rect 574 1542 580 1543
rect 574 1538 575 1542
rect 579 1538 580 1542
rect 574 1537 580 1538
rect 526 1531 532 1532
rect 526 1527 527 1531
rect 531 1527 532 1531
rect 526 1526 532 1527
rect 534 1531 540 1532
rect 534 1527 535 1531
rect 539 1527 540 1531
rect 534 1526 540 1527
rect 295 1522 299 1523
rect 295 1517 299 1518
rect 375 1522 379 1523
rect 375 1517 379 1518
rect 431 1522 435 1523
rect 431 1517 435 1518
rect 519 1522 523 1523
rect 519 1517 523 1518
rect 258 1515 264 1516
rect 258 1511 259 1515
rect 263 1511 264 1515
rect 258 1510 264 1511
rect 282 1515 288 1516
rect 282 1511 283 1515
rect 287 1511 288 1515
rect 282 1510 288 1511
rect 230 1506 236 1507
rect 230 1502 231 1506
rect 235 1502 236 1506
rect 230 1501 236 1502
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 110 1483 116 1484
rect 284 1480 286 1510
rect 376 1507 378 1517
rect 520 1507 522 1517
rect 374 1506 380 1507
rect 374 1502 375 1506
rect 379 1502 380 1506
rect 374 1501 380 1502
rect 518 1506 524 1507
rect 518 1502 519 1506
rect 523 1502 524 1506
rect 518 1501 524 1502
rect 528 1480 530 1526
rect 576 1523 578 1537
rect 660 1532 662 1566
rect 718 1542 724 1543
rect 718 1538 719 1542
rect 723 1538 724 1542
rect 718 1537 724 1538
rect 658 1531 664 1532
rect 658 1527 659 1531
rect 663 1527 664 1531
rect 658 1526 664 1527
rect 720 1523 722 1537
rect 804 1532 806 1566
rect 854 1542 860 1543
rect 854 1538 855 1542
rect 859 1538 860 1542
rect 854 1537 860 1538
rect 990 1542 996 1543
rect 990 1538 991 1542
rect 995 1538 996 1542
rect 990 1537 996 1538
rect 802 1531 808 1532
rect 802 1527 803 1531
rect 807 1527 808 1531
rect 802 1526 808 1527
rect 790 1523 796 1524
rect 856 1523 858 1537
rect 992 1523 994 1537
rect 1052 1532 1054 1566
rect 1126 1542 1132 1543
rect 1126 1538 1127 1542
rect 1131 1538 1132 1542
rect 1126 1537 1132 1538
rect 1254 1542 1260 1543
rect 1254 1538 1255 1542
rect 1259 1538 1260 1542
rect 1254 1537 1260 1538
rect 1014 1531 1020 1532
rect 1050 1531 1056 1532
rect 1014 1527 1015 1531
rect 1019 1529 1026 1531
rect 1019 1527 1020 1529
rect 1014 1526 1020 1527
rect 575 1522 579 1523
rect 575 1517 579 1518
rect 655 1522 659 1523
rect 655 1517 659 1518
rect 719 1522 723 1523
rect 719 1517 723 1518
rect 783 1522 787 1523
rect 790 1519 791 1523
rect 795 1519 796 1523
rect 790 1518 796 1519
rect 855 1522 859 1523
rect 783 1517 787 1518
rect 656 1507 658 1517
rect 698 1515 704 1516
rect 698 1511 699 1515
rect 703 1511 704 1515
rect 698 1510 704 1511
rect 706 1515 712 1516
rect 706 1511 707 1515
rect 711 1511 712 1515
rect 706 1510 712 1511
rect 654 1506 660 1507
rect 654 1502 655 1506
rect 659 1502 660 1506
rect 654 1501 660 1502
rect 282 1479 288 1480
rect 282 1475 283 1479
rect 287 1475 288 1479
rect 282 1474 288 1475
rect 426 1479 432 1480
rect 426 1475 427 1479
rect 431 1475 432 1479
rect 426 1474 432 1475
rect 526 1479 532 1480
rect 526 1475 527 1479
rect 531 1475 532 1479
rect 526 1474 532 1475
rect 110 1471 116 1472
rect 110 1467 111 1471
rect 115 1467 116 1471
rect 110 1466 116 1467
rect 222 1468 228 1469
rect 112 1439 114 1466
rect 222 1464 223 1468
rect 227 1464 228 1468
rect 222 1463 228 1464
rect 366 1468 372 1469
rect 366 1464 367 1468
rect 371 1464 372 1468
rect 366 1463 372 1464
rect 224 1439 226 1463
rect 368 1439 370 1463
rect 111 1438 115 1439
rect 111 1433 115 1434
rect 223 1438 227 1439
rect 223 1433 227 1434
rect 255 1438 259 1439
rect 255 1433 259 1434
rect 351 1438 355 1439
rect 351 1433 355 1434
rect 367 1438 371 1439
rect 367 1433 371 1434
rect 112 1414 114 1433
rect 256 1417 258 1433
rect 352 1417 354 1433
rect 254 1416 260 1417
rect 110 1413 116 1414
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 254 1412 255 1416
rect 259 1412 260 1416
rect 254 1411 260 1412
rect 350 1416 356 1417
rect 350 1412 351 1416
rect 355 1412 356 1416
rect 350 1411 356 1412
rect 110 1408 116 1409
rect 342 1407 348 1408
rect 342 1403 343 1407
rect 347 1403 348 1407
rect 342 1402 348 1403
rect 418 1407 424 1408
rect 418 1403 419 1407
rect 423 1403 424 1407
rect 418 1402 424 1403
rect 314 1399 320 1400
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 314 1395 315 1399
rect 319 1395 320 1399
rect 314 1394 320 1395
rect 110 1391 116 1392
rect 112 1363 114 1391
rect 262 1378 268 1379
rect 262 1374 263 1378
rect 267 1374 268 1378
rect 262 1373 268 1374
rect 264 1363 266 1373
rect 111 1362 115 1363
rect 111 1357 115 1358
rect 263 1362 267 1363
rect 263 1357 267 1358
rect 112 1329 114 1357
rect 316 1356 318 1394
rect 344 1368 346 1402
rect 358 1378 364 1379
rect 358 1374 359 1378
rect 363 1374 364 1378
rect 358 1373 364 1374
rect 342 1367 348 1368
rect 342 1363 343 1367
rect 347 1363 348 1367
rect 360 1363 362 1373
rect 420 1368 422 1402
rect 428 1368 430 1474
rect 510 1468 516 1469
rect 510 1464 511 1468
rect 515 1464 516 1468
rect 510 1463 516 1464
rect 646 1468 652 1469
rect 646 1464 647 1468
rect 651 1464 652 1468
rect 646 1463 652 1464
rect 512 1439 514 1463
rect 648 1439 650 1463
rect 447 1438 451 1439
rect 447 1433 451 1434
rect 511 1438 515 1439
rect 511 1433 515 1434
rect 543 1438 547 1439
rect 543 1433 547 1434
rect 631 1438 635 1439
rect 631 1433 635 1434
rect 647 1438 651 1439
rect 647 1433 651 1434
rect 448 1417 450 1433
rect 544 1417 546 1433
rect 632 1417 634 1433
rect 446 1416 452 1417
rect 446 1412 447 1416
rect 451 1412 452 1416
rect 446 1411 452 1412
rect 542 1416 548 1417
rect 542 1412 543 1416
rect 547 1412 548 1416
rect 542 1411 548 1412
rect 630 1416 636 1417
rect 630 1412 631 1416
rect 635 1412 636 1416
rect 630 1411 636 1412
rect 700 1408 702 1510
rect 708 1480 710 1510
rect 784 1507 786 1517
rect 782 1506 788 1507
rect 782 1502 783 1506
rect 787 1502 788 1506
rect 782 1501 788 1502
rect 792 1480 794 1518
rect 855 1517 859 1518
rect 903 1522 907 1523
rect 903 1517 907 1518
rect 991 1522 995 1523
rect 991 1517 995 1518
rect 1015 1522 1019 1523
rect 1015 1517 1019 1518
rect 904 1507 906 1517
rect 926 1515 932 1516
rect 926 1511 927 1515
rect 931 1511 932 1515
rect 926 1510 932 1511
rect 954 1515 960 1516
rect 954 1511 955 1515
rect 959 1511 960 1515
rect 954 1510 960 1511
rect 902 1506 908 1507
rect 902 1502 903 1506
rect 907 1502 908 1506
rect 902 1501 908 1502
rect 706 1479 712 1480
rect 706 1475 707 1479
rect 711 1475 712 1479
rect 706 1474 712 1475
rect 790 1479 796 1480
rect 790 1475 791 1479
rect 795 1475 796 1479
rect 790 1474 796 1475
rect 774 1468 780 1469
rect 774 1464 775 1468
rect 779 1464 780 1468
rect 774 1463 780 1464
rect 894 1468 900 1469
rect 894 1464 895 1468
rect 899 1464 900 1468
rect 894 1463 900 1464
rect 776 1439 778 1463
rect 896 1439 898 1463
rect 719 1438 723 1439
rect 719 1433 723 1434
rect 775 1438 779 1439
rect 775 1433 779 1434
rect 807 1438 811 1439
rect 807 1433 811 1434
rect 895 1438 899 1439
rect 895 1433 899 1434
rect 919 1438 923 1439
rect 919 1433 923 1434
rect 720 1417 722 1433
rect 808 1417 810 1433
rect 920 1417 922 1433
rect 718 1416 724 1417
rect 718 1412 719 1416
rect 723 1412 724 1416
rect 718 1411 724 1412
rect 806 1416 812 1417
rect 806 1412 807 1416
rect 811 1412 812 1416
rect 806 1411 812 1412
rect 918 1416 924 1417
rect 918 1412 919 1416
rect 923 1412 924 1416
rect 918 1411 924 1412
rect 610 1407 616 1408
rect 610 1403 611 1407
rect 615 1403 616 1407
rect 610 1402 616 1403
rect 698 1407 704 1408
rect 698 1403 699 1407
rect 703 1403 704 1407
rect 698 1402 704 1403
rect 786 1407 792 1408
rect 786 1403 787 1407
rect 791 1403 792 1407
rect 928 1404 930 1510
rect 956 1480 958 1510
rect 1016 1507 1018 1517
rect 1014 1506 1020 1507
rect 1014 1502 1015 1506
rect 1019 1502 1020 1506
rect 1014 1501 1020 1502
rect 1024 1480 1026 1529
rect 1050 1527 1051 1531
rect 1055 1527 1056 1531
rect 1050 1526 1056 1527
rect 1128 1523 1130 1537
rect 1256 1523 1258 1537
rect 1264 1532 1266 1630
rect 1870 1628 1871 1632
rect 1875 1628 1876 1632
rect 1830 1627 1836 1628
rect 1870 1627 1876 1628
rect 1350 1624 1356 1625
rect 1350 1620 1351 1624
rect 1355 1620 1356 1624
rect 1350 1619 1356 1620
rect 1510 1624 1516 1625
rect 1510 1620 1511 1624
rect 1515 1620 1516 1624
rect 1510 1619 1516 1620
rect 1670 1624 1676 1625
rect 1670 1620 1671 1624
rect 1675 1620 1676 1624
rect 1830 1623 1831 1627
rect 1835 1623 1836 1627
rect 1830 1622 1836 1623
rect 1670 1619 1676 1620
rect 1352 1603 1354 1619
rect 1512 1603 1514 1619
rect 1672 1603 1674 1619
rect 1832 1603 1834 1622
rect 1870 1615 1876 1616
rect 1870 1611 1871 1615
rect 1875 1611 1876 1615
rect 1870 1610 1876 1611
rect 1958 1612 1964 1613
rect 1351 1602 1355 1603
rect 1351 1597 1355 1598
rect 1375 1602 1379 1603
rect 1375 1597 1379 1598
rect 1511 1602 1515 1603
rect 1511 1597 1515 1598
rect 1671 1602 1675 1603
rect 1671 1597 1675 1598
rect 1831 1602 1835 1603
rect 1831 1597 1835 1598
rect 1376 1581 1378 1597
rect 1512 1581 1514 1597
rect 1374 1580 1380 1581
rect 1374 1576 1375 1580
rect 1379 1576 1380 1580
rect 1374 1575 1380 1576
rect 1510 1580 1516 1581
rect 1510 1576 1511 1580
rect 1515 1576 1516 1580
rect 1832 1578 1834 1597
rect 1872 1583 1874 1610
rect 1958 1608 1959 1612
rect 1963 1608 1964 1612
rect 1958 1607 1964 1608
rect 1960 1583 1962 1607
rect 1871 1582 1875 1583
rect 1510 1575 1516 1576
rect 1830 1577 1836 1578
rect 1871 1577 1875 1578
rect 1895 1582 1899 1583
rect 1895 1577 1899 1578
rect 1959 1582 1963 1583
rect 1959 1577 1963 1578
rect 1830 1573 1831 1577
rect 1835 1573 1836 1577
rect 1830 1572 1836 1573
rect 1330 1571 1336 1572
rect 1330 1567 1331 1571
rect 1335 1567 1336 1571
rect 1330 1566 1336 1567
rect 1442 1571 1448 1572
rect 1442 1567 1443 1571
rect 1447 1567 1448 1571
rect 1442 1566 1448 1567
rect 1450 1571 1456 1572
rect 1450 1567 1451 1571
rect 1455 1567 1456 1571
rect 1450 1566 1456 1567
rect 1332 1532 1334 1566
rect 1382 1542 1388 1543
rect 1382 1538 1383 1542
rect 1387 1538 1388 1542
rect 1382 1537 1388 1538
rect 1262 1531 1268 1532
rect 1262 1527 1263 1531
rect 1267 1527 1268 1531
rect 1262 1526 1268 1527
rect 1330 1531 1336 1532
rect 1330 1527 1331 1531
rect 1335 1527 1336 1531
rect 1330 1526 1336 1527
rect 1384 1523 1386 1537
rect 1444 1532 1446 1566
rect 1442 1531 1448 1532
rect 1442 1527 1443 1531
rect 1447 1527 1448 1531
rect 1442 1526 1448 1527
rect 1119 1522 1123 1523
rect 1119 1517 1123 1518
rect 1127 1522 1131 1523
rect 1127 1517 1131 1518
rect 1215 1522 1219 1523
rect 1215 1517 1219 1518
rect 1255 1522 1259 1523
rect 1255 1517 1259 1518
rect 1319 1522 1323 1523
rect 1319 1517 1323 1518
rect 1383 1522 1387 1523
rect 1383 1517 1387 1518
rect 1423 1522 1427 1523
rect 1423 1517 1427 1518
rect 1120 1507 1122 1517
rect 1154 1515 1160 1516
rect 1154 1511 1155 1515
rect 1159 1511 1160 1515
rect 1154 1510 1160 1511
rect 1170 1515 1176 1516
rect 1170 1511 1171 1515
rect 1175 1511 1176 1515
rect 1170 1510 1176 1511
rect 1118 1506 1124 1507
rect 1118 1502 1119 1506
rect 1123 1502 1124 1506
rect 1118 1501 1124 1502
rect 1156 1501 1158 1510
rect 1155 1500 1159 1501
rect 1155 1495 1159 1496
rect 1172 1480 1174 1510
rect 1216 1507 1218 1517
rect 1266 1515 1272 1516
rect 1266 1511 1267 1515
rect 1271 1511 1272 1515
rect 1266 1510 1272 1511
rect 1214 1506 1220 1507
rect 1214 1502 1215 1506
rect 1219 1502 1220 1506
rect 1214 1501 1220 1502
rect 1268 1480 1270 1510
rect 1320 1507 1322 1517
rect 1424 1507 1426 1517
rect 1452 1516 1454 1566
rect 1830 1560 1836 1561
rect 1830 1556 1831 1560
rect 1835 1556 1836 1560
rect 1872 1558 1874 1577
rect 1896 1561 1898 1577
rect 1894 1560 1900 1561
rect 1830 1555 1836 1556
rect 1870 1557 1876 1558
rect 1518 1542 1524 1543
rect 1518 1538 1519 1542
rect 1523 1538 1524 1542
rect 1518 1537 1524 1538
rect 1520 1523 1522 1537
rect 1832 1523 1834 1555
rect 1870 1553 1871 1557
rect 1875 1553 1876 1557
rect 1894 1556 1895 1560
rect 1899 1556 1900 1560
rect 1894 1555 1900 1556
rect 1870 1552 1876 1553
rect 1962 1551 1968 1552
rect 1962 1547 1963 1551
rect 1967 1547 1968 1551
rect 1962 1546 1968 1547
rect 1870 1540 1876 1541
rect 1870 1536 1871 1540
rect 1875 1536 1876 1540
rect 1870 1535 1876 1536
rect 1519 1522 1523 1523
rect 1519 1517 1523 1518
rect 1831 1522 1835 1523
rect 1831 1517 1835 1518
rect 1450 1515 1456 1516
rect 1450 1511 1451 1515
rect 1455 1511 1456 1515
rect 1450 1510 1456 1511
rect 1431 1508 1435 1509
rect 1318 1506 1324 1507
rect 1318 1502 1319 1506
rect 1323 1502 1324 1506
rect 1318 1501 1324 1502
rect 1422 1506 1428 1507
rect 1422 1502 1423 1506
rect 1427 1502 1428 1506
rect 1431 1503 1435 1504
rect 1422 1501 1428 1502
rect 1432 1480 1434 1503
rect 1832 1489 1834 1517
rect 1872 1499 1874 1535
rect 1902 1522 1908 1523
rect 1902 1518 1903 1522
rect 1907 1518 1908 1522
rect 1902 1517 1908 1518
rect 1904 1499 1906 1517
rect 1964 1512 1966 1546
rect 1976 1544 1978 1654
rect 2020 1624 2022 1654
rect 2088 1651 2090 1661
rect 2138 1659 2144 1660
rect 2138 1655 2139 1659
rect 2143 1655 2144 1659
rect 2138 1654 2144 1655
rect 2086 1650 2092 1651
rect 2086 1646 2087 1650
rect 2091 1646 2092 1650
rect 2086 1645 2092 1646
rect 2140 1624 2142 1654
rect 2216 1651 2218 1661
rect 2266 1659 2272 1660
rect 2266 1655 2267 1659
rect 2271 1655 2272 1659
rect 2266 1654 2272 1655
rect 2214 1650 2220 1651
rect 2214 1646 2215 1650
rect 2219 1646 2220 1650
rect 2214 1645 2220 1646
rect 2268 1624 2270 1654
rect 2352 1651 2354 1661
rect 2350 1650 2356 1651
rect 2350 1646 2351 1650
rect 2355 1646 2356 1650
rect 2350 1645 2356 1646
rect 2360 1624 2362 1662
rect 2391 1661 2395 1662
rect 2495 1666 2499 1667
rect 2495 1661 2499 1662
rect 2535 1666 2539 1667
rect 2535 1661 2539 1662
rect 2639 1666 2643 1667
rect 2639 1661 2643 1662
rect 2496 1651 2498 1661
rect 2640 1651 2642 1661
rect 2656 1660 2658 1702
rect 2670 1686 2676 1687
rect 2670 1682 2671 1686
rect 2675 1682 2676 1686
rect 2670 1681 2676 1682
rect 2672 1667 2674 1681
rect 2700 1676 2702 1750
rect 2712 1747 2714 1767
rect 2834 1755 2840 1756
rect 2834 1751 2835 1755
rect 2839 1751 2840 1755
rect 2834 1750 2840 1751
rect 2711 1746 2715 1747
rect 2711 1741 2715 1742
rect 2799 1746 2803 1747
rect 2799 1741 2803 1742
rect 2800 1725 2802 1741
rect 2798 1724 2804 1725
rect 2798 1720 2799 1724
rect 2803 1720 2804 1724
rect 2798 1719 2804 1720
rect 2806 1686 2812 1687
rect 2806 1682 2807 1686
rect 2811 1682 2812 1686
rect 2806 1681 2812 1682
rect 2698 1675 2704 1676
rect 2698 1671 2699 1675
rect 2703 1671 2704 1675
rect 2698 1670 2704 1671
rect 2808 1667 2810 1681
rect 2836 1676 2838 1750
rect 2872 1747 2874 1767
rect 3024 1747 3026 1767
rect 2871 1746 2875 1747
rect 2871 1741 2875 1742
rect 2927 1746 2931 1747
rect 2927 1741 2931 1742
rect 3023 1746 3027 1747
rect 3023 1741 3027 1742
rect 3047 1746 3051 1747
rect 3047 1741 3051 1742
rect 2928 1725 2930 1741
rect 3048 1725 3050 1741
rect 2926 1724 2932 1725
rect 2926 1720 2927 1724
rect 2931 1720 2932 1724
rect 2926 1719 2932 1720
rect 3046 1724 3052 1725
rect 3046 1720 3047 1724
rect 3051 1720 3052 1724
rect 3046 1719 3052 1720
rect 3120 1716 3122 1814
rect 3176 1811 3178 1821
rect 3204 1820 3206 1882
rect 3254 1858 3260 1859
rect 3254 1854 3255 1858
rect 3259 1854 3260 1858
rect 3254 1853 3260 1854
rect 3390 1858 3396 1859
rect 3390 1854 3391 1858
rect 3395 1854 3396 1858
rect 3390 1853 3396 1854
rect 3256 1827 3258 1853
rect 3392 1827 3394 1853
rect 3460 1848 3462 1882
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 3458 1847 3464 1848
rect 3458 1843 3459 1847
rect 3463 1843 3464 1847
rect 3458 1842 3464 1843
rect 3512 1827 3514 1853
rect 3536 1848 3538 1954
rect 3590 1951 3596 1952
rect 3590 1947 3591 1951
rect 3595 1947 3596 1951
rect 3590 1946 3596 1947
rect 3592 1919 3594 1946
rect 3591 1918 3595 1919
rect 3591 1913 3595 1914
rect 3592 1894 3594 1913
rect 3590 1893 3596 1894
rect 3590 1889 3591 1893
rect 3595 1889 3596 1893
rect 3590 1888 3596 1889
rect 3590 1876 3596 1877
rect 3590 1872 3591 1876
rect 3595 1872 3596 1876
rect 3590 1871 3596 1872
rect 3534 1847 3540 1848
rect 3534 1843 3535 1847
rect 3539 1843 3540 1847
rect 3534 1842 3540 1843
rect 3592 1827 3594 1871
rect 3255 1826 3259 1827
rect 3255 1821 3259 1822
rect 3319 1826 3323 1827
rect 3319 1821 3323 1822
rect 3391 1826 3395 1827
rect 3391 1821 3395 1822
rect 3471 1826 3475 1827
rect 3471 1821 3475 1822
rect 3511 1826 3515 1827
rect 3511 1821 3515 1822
rect 3591 1826 3595 1827
rect 3591 1821 3595 1822
rect 3202 1819 3208 1820
rect 3202 1815 3203 1819
rect 3207 1815 3208 1819
rect 3202 1814 3208 1815
rect 3226 1819 3232 1820
rect 3226 1815 3227 1819
rect 3231 1815 3232 1819
rect 3226 1814 3232 1815
rect 3174 1810 3180 1811
rect 3174 1806 3175 1810
rect 3179 1806 3180 1810
rect 3174 1805 3180 1806
rect 3228 1784 3230 1814
rect 3320 1811 3322 1821
rect 3370 1819 3376 1820
rect 3370 1815 3371 1819
rect 3375 1815 3376 1819
rect 3370 1814 3376 1815
rect 3318 1810 3324 1811
rect 3318 1806 3319 1810
rect 3323 1806 3324 1810
rect 3318 1805 3324 1806
rect 3372 1784 3374 1814
rect 3472 1811 3474 1821
rect 3470 1810 3476 1811
rect 3470 1806 3471 1810
rect 3475 1806 3476 1810
rect 3470 1805 3476 1806
rect 3592 1793 3594 1821
rect 3590 1792 3596 1793
rect 3590 1788 3591 1792
rect 3595 1788 3596 1792
rect 3590 1787 3596 1788
rect 3226 1783 3232 1784
rect 3226 1779 3227 1783
rect 3231 1779 3232 1783
rect 3226 1778 3232 1779
rect 3370 1783 3376 1784
rect 3370 1779 3371 1783
rect 3375 1779 3376 1783
rect 3370 1778 3376 1779
rect 3590 1775 3596 1776
rect 3166 1772 3172 1773
rect 3166 1768 3167 1772
rect 3171 1768 3172 1772
rect 3166 1767 3172 1768
rect 3310 1772 3316 1773
rect 3310 1768 3311 1772
rect 3315 1768 3316 1772
rect 3310 1767 3316 1768
rect 3462 1772 3468 1773
rect 3462 1768 3463 1772
rect 3467 1768 3468 1772
rect 3590 1771 3591 1775
rect 3595 1771 3596 1775
rect 3590 1770 3596 1771
rect 3462 1767 3468 1768
rect 3168 1747 3170 1767
rect 3312 1747 3314 1767
rect 3426 1755 3432 1756
rect 3426 1751 3427 1755
rect 3431 1751 3432 1755
rect 3426 1750 3432 1751
rect 3159 1746 3163 1747
rect 3159 1741 3163 1742
rect 3167 1746 3171 1747
rect 3167 1741 3171 1742
rect 3271 1746 3275 1747
rect 3271 1741 3275 1742
rect 3311 1746 3315 1747
rect 3311 1741 3315 1742
rect 3391 1746 3395 1747
rect 3391 1741 3395 1742
rect 3160 1725 3162 1741
rect 3272 1725 3274 1741
rect 3392 1725 3394 1741
rect 3158 1724 3164 1725
rect 3158 1720 3159 1724
rect 3163 1720 3164 1724
rect 3158 1719 3164 1720
rect 3270 1724 3276 1725
rect 3270 1720 3271 1724
rect 3275 1720 3276 1724
rect 3270 1719 3276 1720
rect 3390 1724 3396 1725
rect 3390 1720 3391 1724
rect 3395 1720 3396 1724
rect 3390 1719 3396 1720
rect 2898 1715 2904 1716
rect 2898 1711 2899 1715
rect 2903 1711 2904 1715
rect 2898 1710 2904 1711
rect 3002 1715 3008 1716
rect 3002 1711 3003 1715
rect 3007 1711 3008 1715
rect 3002 1710 3008 1711
rect 3118 1715 3124 1716
rect 3118 1711 3119 1715
rect 3123 1711 3124 1715
rect 3118 1710 3124 1711
rect 3226 1715 3232 1716
rect 3226 1711 3227 1715
rect 3231 1711 3232 1715
rect 3226 1710 3232 1711
rect 2900 1676 2902 1710
rect 2934 1686 2940 1687
rect 2934 1682 2935 1686
rect 2939 1682 2940 1686
rect 2934 1681 2940 1682
rect 2834 1675 2840 1676
rect 2834 1671 2835 1675
rect 2839 1671 2840 1675
rect 2834 1670 2840 1671
rect 2898 1675 2904 1676
rect 2898 1671 2899 1675
rect 2903 1671 2904 1675
rect 2898 1670 2904 1671
rect 2936 1667 2938 1681
rect 3004 1676 3006 1710
rect 3106 1707 3112 1708
rect 3106 1703 3107 1707
rect 3111 1703 3112 1707
rect 3106 1702 3112 1703
rect 3054 1686 3060 1687
rect 3054 1682 3055 1686
rect 3059 1682 3060 1686
rect 3054 1681 3060 1682
rect 3002 1675 3008 1676
rect 3002 1671 3003 1675
rect 3007 1671 3008 1675
rect 3002 1670 3008 1671
rect 3056 1667 3058 1681
rect 2671 1666 2675 1667
rect 2671 1661 2675 1662
rect 2783 1666 2787 1667
rect 2783 1661 2787 1662
rect 2807 1666 2811 1667
rect 2807 1661 2811 1662
rect 2927 1666 2931 1667
rect 2927 1661 2931 1662
rect 2935 1666 2939 1667
rect 2935 1661 2939 1662
rect 3055 1666 3059 1667
rect 3055 1661 3059 1662
rect 3071 1666 3075 1667
rect 3071 1661 3075 1662
rect 2646 1659 2652 1660
rect 2646 1655 2647 1659
rect 2651 1655 2652 1659
rect 2646 1654 2652 1655
rect 2654 1659 2660 1660
rect 2654 1655 2655 1659
rect 2659 1655 2660 1659
rect 2654 1654 2660 1655
rect 2494 1650 2500 1651
rect 2494 1646 2495 1650
rect 2499 1646 2500 1650
rect 2494 1645 2500 1646
rect 2638 1650 2644 1651
rect 2638 1646 2639 1650
rect 2643 1646 2644 1650
rect 2638 1645 2644 1646
rect 2648 1624 2650 1654
rect 2784 1651 2786 1661
rect 2928 1651 2930 1661
rect 3072 1651 3074 1661
rect 3108 1660 3110 1702
rect 3166 1686 3172 1687
rect 3166 1682 3167 1686
rect 3171 1682 3172 1686
rect 3166 1681 3172 1682
rect 3168 1667 3170 1681
rect 3228 1676 3230 1710
rect 3278 1686 3284 1687
rect 3278 1682 3279 1686
rect 3283 1682 3284 1686
rect 3278 1681 3284 1682
rect 3398 1686 3404 1687
rect 3398 1682 3399 1686
rect 3403 1682 3404 1686
rect 3398 1681 3404 1682
rect 3226 1675 3232 1676
rect 3226 1671 3227 1675
rect 3231 1671 3232 1675
rect 3226 1670 3232 1671
rect 3280 1667 3282 1681
rect 3382 1675 3388 1676
rect 3382 1671 3383 1675
rect 3387 1671 3388 1675
rect 3382 1670 3388 1671
rect 3167 1666 3171 1667
rect 3167 1661 3171 1662
rect 3223 1666 3227 1667
rect 3223 1661 3227 1662
rect 3279 1666 3283 1667
rect 3279 1661 3283 1662
rect 3375 1666 3379 1667
rect 3375 1661 3379 1662
rect 3078 1659 3084 1660
rect 3078 1655 3079 1659
rect 3083 1655 3084 1659
rect 3078 1654 3084 1655
rect 3106 1659 3112 1660
rect 3106 1655 3107 1659
rect 3111 1655 3112 1659
rect 3106 1654 3112 1655
rect 3178 1659 3184 1660
rect 3178 1655 3179 1659
rect 3183 1655 3184 1659
rect 3178 1654 3184 1655
rect 2782 1650 2788 1651
rect 2782 1646 2783 1650
rect 2787 1646 2788 1650
rect 2782 1645 2788 1646
rect 2926 1650 2932 1651
rect 2926 1646 2927 1650
rect 2931 1646 2932 1650
rect 2926 1645 2932 1646
rect 3070 1650 3076 1651
rect 3070 1646 3071 1650
rect 3075 1646 3076 1650
rect 3070 1645 3076 1646
rect 3080 1624 3082 1654
rect 2018 1623 2024 1624
rect 2018 1619 2019 1623
rect 2023 1619 2024 1623
rect 2018 1618 2024 1619
rect 2138 1623 2144 1624
rect 2138 1619 2139 1623
rect 2143 1619 2144 1623
rect 2138 1618 2144 1619
rect 2266 1623 2272 1624
rect 2266 1619 2267 1623
rect 2271 1619 2272 1623
rect 2266 1618 2272 1619
rect 2358 1623 2364 1624
rect 2358 1619 2359 1623
rect 2363 1619 2364 1623
rect 2358 1618 2364 1619
rect 2546 1623 2552 1624
rect 2546 1619 2547 1623
rect 2551 1619 2552 1623
rect 2546 1618 2552 1619
rect 2646 1623 2652 1624
rect 2646 1619 2647 1623
rect 2651 1619 2652 1623
rect 2646 1618 2652 1619
rect 3078 1623 3084 1624
rect 3078 1619 3079 1623
rect 3083 1619 3084 1623
rect 3078 1618 3084 1619
rect 2078 1612 2084 1613
rect 2078 1608 2079 1612
rect 2083 1608 2084 1612
rect 2078 1607 2084 1608
rect 2206 1612 2212 1613
rect 2206 1608 2207 1612
rect 2211 1608 2212 1612
rect 2206 1607 2212 1608
rect 2342 1612 2348 1613
rect 2342 1608 2343 1612
rect 2347 1608 2348 1612
rect 2342 1607 2348 1608
rect 2486 1612 2492 1613
rect 2486 1608 2487 1612
rect 2491 1608 2492 1612
rect 2486 1607 2492 1608
rect 2080 1583 2082 1607
rect 2208 1583 2210 1607
rect 2344 1583 2346 1607
rect 2488 1583 2490 1607
rect 2047 1582 2051 1583
rect 2047 1577 2051 1578
rect 2079 1582 2083 1583
rect 2079 1577 2083 1578
rect 2207 1582 2211 1583
rect 2207 1577 2211 1578
rect 2343 1582 2347 1583
rect 2343 1577 2347 1578
rect 2367 1582 2371 1583
rect 2367 1577 2371 1578
rect 2487 1582 2491 1583
rect 2487 1577 2491 1578
rect 2527 1582 2531 1583
rect 2527 1577 2531 1578
rect 2048 1561 2050 1577
rect 2208 1561 2210 1577
rect 2368 1561 2370 1577
rect 2528 1561 2530 1577
rect 2046 1560 2052 1561
rect 2046 1556 2047 1560
rect 2051 1556 2052 1560
rect 2046 1555 2052 1556
rect 2206 1560 2212 1561
rect 2206 1556 2207 1560
rect 2211 1556 2212 1560
rect 2206 1555 2212 1556
rect 2366 1560 2372 1561
rect 2366 1556 2367 1560
rect 2371 1556 2372 1560
rect 2366 1555 2372 1556
rect 2526 1560 2532 1561
rect 2526 1556 2527 1560
rect 2531 1556 2532 1560
rect 2526 1555 2532 1556
rect 2114 1551 2120 1552
rect 2114 1547 2115 1551
rect 2119 1547 2120 1551
rect 2114 1546 2120 1547
rect 2434 1551 2440 1552
rect 2434 1547 2435 1551
rect 2439 1547 2440 1551
rect 2434 1546 2440 1547
rect 1974 1543 1980 1544
rect 1974 1539 1975 1543
rect 1979 1539 1980 1543
rect 1974 1538 1980 1539
rect 2054 1522 2060 1523
rect 2054 1518 2055 1522
rect 2059 1518 2060 1522
rect 2054 1517 2060 1518
rect 1962 1511 1968 1512
rect 1962 1507 1963 1511
rect 1967 1507 1968 1511
rect 1962 1506 1968 1507
rect 2056 1499 2058 1517
rect 2116 1512 2118 1546
rect 2214 1522 2220 1523
rect 2214 1518 2215 1522
rect 2219 1518 2220 1522
rect 2214 1517 2220 1518
rect 2374 1522 2380 1523
rect 2374 1518 2375 1522
rect 2379 1518 2380 1522
rect 2374 1517 2380 1518
rect 2114 1511 2120 1512
rect 2114 1507 2115 1511
rect 2119 1507 2120 1511
rect 2114 1506 2120 1507
rect 2186 1511 2192 1512
rect 2186 1507 2187 1511
rect 2191 1507 2192 1511
rect 2186 1506 2192 1507
rect 1871 1498 1875 1499
rect 1871 1493 1875 1494
rect 1903 1498 1907 1499
rect 1903 1493 1907 1494
rect 2007 1498 2011 1499
rect 2007 1493 2011 1494
rect 2055 1498 2059 1499
rect 2055 1493 2059 1494
rect 2135 1498 2139 1499
rect 2135 1493 2139 1494
rect 1830 1488 1836 1489
rect 1830 1484 1831 1488
rect 1835 1484 1836 1488
rect 1830 1483 1836 1484
rect 954 1479 960 1480
rect 954 1475 955 1479
rect 959 1475 960 1479
rect 954 1474 960 1475
rect 1022 1479 1028 1480
rect 1022 1475 1023 1479
rect 1027 1475 1028 1479
rect 1022 1474 1028 1475
rect 1170 1479 1176 1480
rect 1170 1475 1171 1479
rect 1175 1475 1176 1479
rect 1170 1474 1176 1475
rect 1266 1479 1272 1480
rect 1266 1475 1267 1479
rect 1271 1475 1272 1479
rect 1266 1474 1272 1475
rect 1370 1479 1376 1480
rect 1370 1475 1371 1479
rect 1375 1475 1376 1479
rect 1370 1474 1376 1475
rect 1430 1479 1436 1480
rect 1430 1475 1431 1479
rect 1435 1475 1436 1479
rect 1430 1474 1436 1475
rect 1006 1468 1012 1469
rect 1006 1464 1007 1468
rect 1011 1464 1012 1468
rect 1006 1463 1012 1464
rect 1110 1468 1116 1469
rect 1110 1464 1111 1468
rect 1115 1464 1116 1468
rect 1110 1463 1116 1464
rect 1206 1468 1212 1469
rect 1206 1464 1207 1468
rect 1211 1464 1212 1468
rect 1206 1463 1212 1464
rect 1310 1468 1316 1469
rect 1310 1464 1311 1468
rect 1315 1464 1316 1468
rect 1310 1463 1316 1464
rect 1008 1439 1010 1463
rect 1112 1439 1114 1463
rect 1208 1439 1210 1463
rect 1312 1439 1314 1463
rect 1007 1438 1011 1439
rect 1007 1433 1011 1434
rect 1047 1438 1051 1439
rect 1047 1433 1051 1434
rect 1111 1438 1115 1439
rect 1111 1433 1115 1434
rect 1207 1438 1211 1439
rect 1207 1433 1211 1434
rect 1311 1438 1315 1439
rect 1311 1433 1315 1434
rect 1048 1417 1050 1433
rect 1208 1417 1210 1433
rect 1046 1416 1052 1417
rect 1046 1412 1047 1416
rect 1051 1412 1052 1416
rect 1046 1411 1052 1412
rect 1206 1416 1212 1417
rect 1206 1412 1207 1416
rect 1211 1412 1212 1416
rect 1206 1411 1212 1412
rect 986 1407 992 1408
rect 786 1402 792 1403
rect 926 1403 932 1404
rect 602 1399 608 1400
rect 602 1395 603 1399
rect 607 1395 608 1399
rect 602 1394 608 1395
rect 454 1378 460 1379
rect 454 1374 455 1378
rect 459 1374 460 1378
rect 454 1373 460 1374
rect 550 1378 556 1379
rect 550 1374 551 1378
rect 555 1374 556 1378
rect 550 1373 556 1374
rect 418 1367 424 1368
rect 418 1363 419 1367
rect 423 1363 424 1367
rect 342 1362 348 1363
rect 359 1362 363 1363
rect 418 1362 424 1363
rect 426 1367 432 1368
rect 426 1363 427 1367
rect 431 1363 432 1367
rect 456 1363 458 1373
rect 552 1363 554 1373
rect 604 1368 606 1394
rect 612 1368 614 1402
rect 638 1378 644 1379
rect 638 1374 639 1378
rect 643 1374 644 1378
rect 638 1373 644 1374
rect 726 1378 732 1379
rect 726 1374 727 1378
rect 731 1374 732 1378
rect 726 1373 732 1374
rect 602 1367 608 1368
rect 602 1363 603 1367
rect 607 1363 608 1367
rect 426 1362 432 1363
rect 455 1362 459 1363
rect 359 1357 363 1358
rect 455 1357 459 1358
rect 471 1362 475 1363
rect 471 1357 475 1358
rect 551 1362 555 1363
rect 551 1357 555 1358
rect 591 1362 595 1363
rect 602 1362 608 1363
rect 610 1367 616 1368
rect 610 1363 611 1367
rect 615 1363 616 1367
rect 640 1363 642 1373
rect 728 1363 730 1373
rect 788 1368 790 1402
rect 926 1399 927 1403
rect 931 1399 932 1403
rect 986 1403 987 1407
rect 991 1403 992 1407
rect 986 1402 992 1403
rect 1114 1407 1120 1408
rect 1114 1403 1115 1407
rect 1119 1403 1120 1407
rect 1114 1402 1120 1403
rect 926 1398 932 1399
rect 988 1388 990 1402
rect 870 1387 876 1388
rect 870 1383 871 1387
rect 875 1383 876 1387
rect 870 1382 876 1383
rect 986 1387 992 1388
rect 986 1383 987 1387
rect 991 1383 992 1387
rect 986 1382 992 1383
rect 814 1378 820 1379
rect 814 1374 815 1378
rect 819 1374 820 1378
rect 814 1373 820 1374
rect 786 1367 792 1368
rect 786 1363 787 1367
rect 791 1363 792 1367
rect 816 1363 818 1373
rect 872 1368 874 1382
rect 926 1378 932 1379
rect 926 1374 927 1378
rect 931 1374 932 1378
rect 926 1373 932 1374
rect 1054 1378 1060 1379
rect 1054 1374 1055 1378
rect 1059 1374 1060 1378
rect 1054 1373 1060 1374
rect 870 1367 876 1368
rect 870 1363 871 1367
rect 875 1363 876 1367
rect 610 1362 616 1363
rect 639 1362 643 1363
rect 591 1357 595 1358
rect 639 1357 643 1358
rect 727 1362 731 1363
rect 786 1362 792 1363
rect 815 1362 819 1363
rect 727 1357 731 1358
rect 815 1357 819 1358
rect 863 1362 867 1363
rect 870 1362 876 1363
rect 914 1367 920 1368
rect 914 1363 915 1367
rect 919 1363 920 1367
rect 928 1363 930 1373
rect 1056 1363 1058 1373
rect 1116 1368 1118 1402
rect 1214 1378 1220 1379
rect 1214 1374 1215 1378
rect 1219 1374 1220 1378
rect 1214 1373 1220 1374
rect 1114 1367 1120 1368
rect 1114 1363 1115 1367
rect 1119 1363 1120 1367
rect 1216 1363 1218 1373
rect 1243 1372 1247 1373
rect 1372 1368 1374 1474
rect 1830 1471 1836 1472
rect 1414 1468 1420 1469
rect 1414 1464 1415 1468
rect 1419 1464 1420 1468
rect 1830 1467 1831 1471
rect 1835 1467 1836 1471
rect 1830 1466 1836 1467
rect 1414 1463 1420 1464
rect 1416 1439 1418 1463
rect 1832 1439 1834 1466
rect 1872 1465 1874 1493
rect 1904 1483 1906 1493
rect 1962 1491 1968 1492
rect 1962 1487 1963 1491
rect 1967 1487 1968 1491
rect 1962 1486 1968 1487
rect 1970 1491 1976 1492
rect 1970 1487 1971 1491
rect 1975 1487 1976 1491
rect 1970 1486 1976 1487
rect 1902 1482 1908 1483
rect 1902 1478 1903 1482
rect 1907 1478 1908 1482
rect 1902 1477 1908 1478
rect 1870 1464 1876 1465
rect 1870 1460 1871 1464
rect 1875 1460 1876 1464
rect 1870 1459 1876 1460
rect 1870 1447 1876 1448
rect 1870 1443 1871 1447
rect 1875 1443 1876 1447
rect 1870 1442 1876 1443
rect 1894 1444 1900 1445
rect 1383 1438 1387 1439
rect 1383 1433 1387 1434
rect 1415 1438 1419 1439
rect 1415 1433 1419 1434
rect 1575 1438 1579 1439
rect 1575 1433 1579 1434
rect 1743 1438 1747 1439
rect 1743 1433 1747 1434
rect 1831 1438 1835 1439
rect 1831 1433 1835 1434
rect 1384 1417 1386 1433
rect 1576 1417 1578 1433
rect 1744 1417 1746 1433
rect 1382 1416 1388 1417
rect 1382 1412 1383 1416
rect 1387 1412 1388 1416
rect 1382 1411 1388 1412
rect 1574 1416 1580 1417
rect 1574 1412 1575 1416
rect 1579 1412 1580 1416
rect 1574 1411 1580 1412
rect 1742 1416 1748 1417
rect 1742 1412 1743 1416
rect 1747 1412 1748 1416
rect 1832 1414 1834 1433
rect 1872 1423 1874 1442
rect 1894 1440 1895 1444
rect 1899 1440 1900 1444
rect 1894 1439 1900 1440
rect 1896 1423 1898 1439
rect 1871 1422 1875 1423
rect 1871 1417 1875 1418
rect 1895 1422 1899 1423
rect 1895 1417 1899 1418
rect 1742 1411 1748 1412
rect 1830 1413 1836 1414
rect 1830 1409 1831 1413
rect 1835 1409 1836 1413
rect 1830 1408 1836 1409
rect 1502 1407 1508 1408
rect 1502 1403 1503 1407
rect 1507 1403 1508 1407
rect 1502 1402 1508 1403
rect 1518 1407 1524 1408
rect 1518 1403 1519 1407
rect 1523 1403 1524 1407
rect 1518 1402 1524 1403
rect 1810 1407 1816 1408
rect 1810 1403 1811 1407
rect 1815 1403 1816 1407
rect 1810 1402 1816 1403
rect 1390 1378 1396 1379
rect 1390 1374 1391 1378
rect 1395 1374 1396 1378
rect 1390 1373 1396 1374
rect 1242 1367 1248 1368
rect 1242 1363 1243 1367
rect 1247 1363 1248 1367
rect 1370 1367 1376 1368
rect 1370 1363 1371 1367
rect 1375 1363 1376 1367
rect 1392 1363 1394 1373
rect 1504 1368 1506 1402
rect 1520 1373 1522 1402
rect 1582 1378 1588 1379
rect 1582 1374 1583 1378
rect 1587 1374 1588 1378
rect 1582 1373 1588 1374
rect 1750 1378 1756 1379
rect 1750 1374 1751 1378
rect 1755 1374 1756 1378
rect 1750 1373 1756 1374
rect 1519 1372 1523 1373
rect 1502 1367 1508 1368
rect 1519 1367 1523 1368
rect 1502 1363 1503 1367
rect 1507 1363 1508 1367
rect 1584 1363 1586 1373
rect 1752 1363 1754 1373
rect 1774 1367 1780 1368
rect 1774 1363 1775 1367
rect 1779 1363 1780 1367
rect 914 1362 920 1363
rect 927 1362 931 1363
rect 863 1357 867 1358
rect 314 1355 320 1356
rect 314 1351 315 1355
rect 319 1351 320 1355
rect 314 1350 320 1351
rect 360 1347 362 1357
rect 410 1355 416 1356
rect 410 1351 411 1355
rect 415 1351 416 1355
rect 410 1350 416 1351
rect 358 1346 364 1347
rect 358 1342 359 1346
rect 363 1342 364 1346
rect 358 1341 364 1342
rect 110 1328 116 1329
rect 110 1324 111 1328
rect 115 1324 116 1328
rect 110 1323 116 1324
rect 412 1320 414 1350
rect 472 1347 474 1357
rect 522 1355 528 1356
rect 522 1351 523 1355
rect 527 1351 528 1355
rect 522 1350 528 1351
rect 470 1346 476 1347
rect 470 1342 471 1346
rect 475 1342 476 1346
rect 470 1341 476 1342
rect 524 1320 526 1350
rect 592 1347 594 1357
rect 718 1355 724 1356
rect 718 1351 719 1355
rect 723 1351 724 1355
rect 718 1350 724 1351
rect 590 1346 596 1347
rect 590 1342 591 1346
rect 595 1342 596 1346
rect 590 1341 596 1342
rect 720 1320 722 1350
rect 728 1347 730 1357
rect 864 1347 866 1357
rect 726 1346 732 1347
rect 726 1342 727 1346
rect 731 1342 732 1346
rect 726 1341 732 1342
rect 862 1346 868 1347
rect 862 1342 863 1346
rect 867 1342 868 1346
rect 862 1341 868 1342
rect 916 1320 918 1362
rect 927 1357 931 1358
rect 1007 1362 1011 1363
rect 1007 1357 1011 1358
rect 1055 1362 1059 1363
rect 1114 1362 1120 1363
rect 1143 1362 1147 1363
rect 1055 1357 1059 1358
rect 1143 1357 1147 1358
rect 1215 1362 1219 1363
rect 1242 1362 1248 1363
rect 1279 1362 1283 1363
rect 1370 1362 1376 1363
rect 1391 1362 1395 1363
rect 1215 1357 1219 1358
rect 1279 1357 1283 1358
rect 1391 1357 1395 1358
rect 1407 1362 1411 1363
rect 1502 1362 1508 1363
rect 1527 1362 1531 1363
rect 1407 1357 1411 1358
rect 1527 1357 1531 1358
rect 1583 1362 1587 1363
rect 1583 1357 1587 1358
rect 1647 1362 1651 1363
rect 1647 1357 1651 1358
rect 1751 1362 1755 1363
rect 1774 1362 1780 1363
rect 1751 1357 1755 1358
rect 1008 1347 1010 1357
rect 1014 1355 1020 1356
rect 1014 1351 1015 1355
rect 1019 1351 1020 1355
rect 1014 1350 1020 1351
rect 1006 1346 1012 1347
rect 1006 1342 1007 1346
rect 1011 1342 1012 1346
rect 1006 1341 1012 1342
rect 1016 1320 1018 1350
rect 1144 1347 1146 1357
rect 1150 1355 1156 1356
rect 1150 1351 1151 1355
rect 1155 1351 1156 1355
rect 1150 1350 1156 1351
rect 1170 1355 1176 1356
rect 1170 1351 1171 1355
rect 1175 1351 1176 1355
rect 1170 1350 1176 1351
rect 1142 1346 1148 1347
rect 1142 1342 1143 1346
rect 1147 1342 1148 1346
rect 1142 1341 1148 1342
rect 1152 1320 1154 1350
rect 410 1319 416 1320
rect 410 1315 411 1319
rect 415 1315 416 1319
rect 410 1314 416 1315
rect 522 1319 528 1320
rect 522 1315 523 1319
rect 527 1315 528 1319
rect 522 1314 528 1315
rect 718 1319 724 1320
rect 718 1315 719 1319
rect 723 1315 724 1319
rect 718 1314 724 1315
rect 914 1319 920 1320
rect 914 1315 915 1319
rect 919 1315 920 1319
rect 914 1314 920 1315
rect 1014 1319 1020 1320
rect 1014 1315 1015 1319
rect 1019 1315 1020 1319
rect 1014 1314 1020 1315
rect 1150 1319 1156 1320
rect 1150 1315 1151 1319
rect 1155 1315 1156 1319
rect 1150 1314 1156 1315
rect 110 1311 116 1312
rect 110 1307 111 1311
rect 115 1307 116 1311
rect 110 1306 116 1307
rect 350 1308 356 1309
rect 112 1283 114 1306
rect 350 1304 351 1308
rect 355 1304 356 1308
rect 350 1303 356 1304
rect 462 1308 468 1309
rect 462 1304 463 1308
rect 467 1304 468 1308
rect 462 1303 468 1304
rect 582 1308 588 1309
rect 582 1304 583 1308
rect 587 1304 588 1308
rect 582 1303 588 1304
rect 718 1308 724 1309
rect 718 1304 719 1308
rect 723 1304 724 1308
rect 718 1303 724 1304
rect 854 1308 860 1309
rect 854 1304 855 1308
rect 859 1304 860 1308
rect 854 1303 860 1304
rect 998 1308 1004 1309
rect 998 1304 999 1308
rect 1003 1304 1004 1308
rect 998 1303 1004 1304
rect 1134 1308 1140 1309
rect 1134 1304 1135 1308
rect 1139 1304 1140 1308
rect 1134 1303 1140 1304
rect 352 1283 354 1303
rect 464 1283 466 1303
rect 584 1283 586 1303
rect 706 1291 712 1292
rect 706 1287 707 1291
rect 711 1287 712 1291
rect 706 1286 712 1287
rect 111 1282 115 1283
rect 111 1277 115 1278
rect 311 1282 315 1283
rect 311 1277 315 1278
rect 351 1282 355 1283
rect 351 1277 355 1278
rect 415 1282 419 1283
rect 415 1277 419 1278
rect 463 1282 467 1283
rect 463 1277 467 1278
rect 535 1282 539 1283
rect 535 1277 539 1278
rect 583 1282 587 1283
rect 583 1277 587 1278
rect 671 1282 675 1283
rect 671 1277 675 1278
rect 112 1258 114 1277
rect 312 1261 314 1277
rect 416 1261 418 1277
rect 536 1261 538 1277
rect 672 1261 674 1277
rect 310 1260 316 1261
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 310 1256 311 1260
rect 315 1256 316 1260
rect 310 1255 316 1256
rect 414 1260 420 1261
rect 414 1256 415 1260
rect 419 1256 420 1260
rect 414 1255 420 1256
rect 534 1260 540 1261
rect 534 1256 535 1260
rect 539 1256 540 1260
rect 534 1255 540 1256
rect 670 1260 676 1261
rect 670 1256 671 1260
rect 675 1256 676 1260
rect 670 1255 676 1256
rect 110 1252 116 1253
rect 266 1251 272 1252
rect 266 1247 267 1251
rect 271 1247 272 1251
rect 266 1246 272 1247
rect 378 1251 384 1252
rect 378 1247 379 1251
rect 383 1247 384 1251
rect 378 1246 384 1247
rect 482 1251 488 1252
rect 482 1247 483 1251
rect 487 1247 488 1251
rect 482 1246 488 1247
rect 602 1251 608 1252
rect 602 1247 603 1251
rect 607 1247 608 1251
rect 602 1246 608 1247
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 112 1207 114 1235
rect 111 1206 115 1207
rect 111 1201 115 1202
rect 239 1206 243 1207
rect 239 1201 243 1202
rect 112 1173 114 1201
rect 240 1191 242 1201
rect 268 1200 270 1246
rect 318 1222 324 1223
rect 318 1218 319 1222
rect 323 1218 324 1222
rect 318 1217 324 1218
rect 320 1207 322 1217
rect 380 1212 382 1246
rect 422 1222 428 1223
rect 422 1218 423 1222
rect 427 1218 428 1222
rect 422 1217 428 1218
rect 378 1211 384 1212
rect 378 1207 379 1211
rect 383 1207 384 1211
rect 424 1207 426 1217
rect 484 1212 486 1246
rect 542 1222 548 1223
rect 542 1218 543 1222
rect 547 1218 548 1222
rect 542 1217 548 1218
rect 482 1211 488 1212
rect 482 1207 483 1211
rect 487 1207 488 1211
rect 544 1207 546 1217
rect 604 1212 606 1246
rect 678 1222 684 1223
rect 678 1218 679 1222
rect 683 1218 684 1222
rect 678 1217 684 1218
rect 602 1211 608 1212
rect 602 1207 603 1211
rect 607 1207 608 1211
rect 680 1207 682 1217
rect 708 1212 710 1286
rect 720 1283 722 1303
rect 856 1283 858 1303
rect 1000 1283 1002 1303
rect 1136 1283 1138 1303
rect 719 1282 723 1283
rect 719 1277 723 1278
rect 815 1282 819 1283
rect 815 1277 819 1278
rect 855 1282 859 1283
rect 855 1277 859 1278
rect 959 1282 963 1283
rect 959 1277 963 1278
rect 999 1282 1003 1283
rect 999 1277 1003 1278
rect 1103 1282 1107 1283
rect 1103 1277 1107 1278
rect 1135 1282 1139 1283
rect 1135 1277 1139 1278
rect 816 1261 818 1277
rect 960 1261 962 1277
rect 1104 1261 1106 1277
rect 814 1260 820 1261
rect 814 1256 815 1260
rect 819 1256 820 1260
rect 814 1255 820 1256
rect 958 1260 964 1261
rect 958 1256 959 1260
rect 963 1256 964 1260
rect 958 1255 964 1256
rect 1102 1260 1108 1261
rect 1102 1256 1103 1260
rect 1107 1256 1108 1260
rect 1102 1255 1108 1256
rect 1172 1252 1174 1350
rect 1280 1347 1282 1357
rect 1306 1355 1312 1356
rect 1306 1351 1307 1355
rect 1311 1351 1312 1355
rect 1306 1350 1312 1351
rect 1330 1355 1336 1356
rect 1330 1351 1331 1355
rect 1335 1351 1336 1355
rect 1330 1350 1336 1351
rect 1278 1346 1284 1347
rect 1278 1342 1279 1346
rect 1283 1342 1284 1346
rect 1278 1341 1284 1342
rect 1270 1308 1276 1309
rect 1270 1304 1271 1308
rect 1275 1304 1276 1308
rect 1270 1303 1276 1304
rect 1272 1283 1274 1303
rect 1308 1301 1310 1350
rect 1332 1320 1334 1350
rect 1408 1347 1410 1357
rect 1458 1355 1464 1356
rect 1458 1351 1459 1355
rect 1463 1351 1464 1355
rect 1458 1350 1464 1351
rect 1406 1346 1412 1347
rect 1406 1342 1407 1346
rect 1411 1342 1412 1346
rect 1406 1341 1412 1342
rect 1460 1320 1462 1350
rect 1528 1347 1530 1357
rect 1648 1347 1650 1357
rect 1698 1355 1704 1356
rect 1698 1351 1699 1355
rect 1703 1351 1704 1355
rect 1698 1350 1704 1351
rect 1526 1346 1532 1347
rect 1526 1342 1527 1346
rect 1531 1342 1532 1346
rect 1526 1341 1532 1342
rect 1646 1346 1652 1347
rect 1646 1342 1647 1346
rect 1651 1342 1652 1346
rect 1646 1341 1652 1342
rect 1700 1320 1702 1350
rect 1752 1347 1754 1357
rect 1750 1346 1756 1347
rect 1750 1342 1751 1346
rect 1755 1342 1756 1346
rect 1750 1341 1756 1342
rect 1776 1320 1778 1362
rect 1812 1352 1814 1402
rect 1872 1398 1874 1417
rect 1896 1401 1898 1417
rect 1894 1400 1900 1401
rect 1870 1397 1876 1398
rect 1830 1396 1836 1397
rect 1830 1392 1831 1396
rect 1835 1392 1836 1396
rect 1870 1393 1871 1397
rect 1875 1393 1876 1397
rect 1894 1396 1895 1400
rect 1899 1396 1900 1400
rect 1894 1395 1900 1396
rect 1870 1392 1876 1393
rect 1964 1392 1966 1486
rect 1972 1456 1974 1486
rect 2008 1483 2010 1493
rect 2126 1491 2132 1492
rect 2126 1487 2127 1491
rect 2131 1487 2132 1491
rect 2126 1486 2132 1487
rect 2006 1482 2012 1483
rect 2006 1478 2007 1482
rect 2011 1478 2012 1482
rect 2006 1477 2012 1478
rect 2128 1456 2130 1486
rect 2136 1483 2138 1493
rect 2134 1482 2140 1483
rect 2134 1478 2135 1482
rect 2139 1478 2140 1482
rect 2134 1477 2140 1478
rect 2188 1456 2190 1506
rect 2216 1499 2218 1517
rect 2376 1499 2378 1517
rect 2436 1512 2438 1546
rect 2442 1543 2448 1544
rect 2442 1539 2443 1543
rect 2447 1539 2448 1543
rect 2442 1538 2448 1539
rect 2434 1511 2440 1512
rect 2434 1507 2435 1511
rect 2439 1507 2440 1511
rect 2434 1506 2440 1507
rect 2215 1498 2219 1499
rect 2215 1493 2219 1494
rect 2271 1498 2275 1499
rect 2271 1493 2275 1494
rect 2375 1498 2379 1499
rect 2375 1493 2379 1494
rect 2415 1498 2419 1499
rect 2415 1493 2419 1494
rect 2272 1483 2274 1493
rect 2416 1483 2418 1493
rect 2444 1492 2446 1538
rect 2534 1522 2540 1523
rect 2534 1518 2535 1522
rect 2539 1518 2540 1522
rect 2534 1517 2540 1518
rect 2536 1499 2538 1517
rect 2548 1512 2550 1618
rect 2630 1612 2636 1613
rect 2630 1608 2631 1612
rect 2635 1608 2636 1612
rect 2630 1607 2636 1608
rect 2774 1612 2780 1613
rect 2774 1608 2775 1612
rect 2779 1608 2780 1612
rect 2774 1607 2780 1608
rect 2918 1612 2924 1613
rect 2918 1608 2919 1612
rect 2923 1608 2924 1612
rect 2918 1607 2924 1608
rect 3062 1612 3068 1613
rect 3062 1608 3063 1612
rect 3067 1608 3068 1612
rect 3062 1607 3068 1608
rect 2632 1583 2634 1607
rect 2722 1595 2728 1596
rect 2722 1591 2723 1595
rect 2727 1591 2728 1595
rect 2722 1590 2728 1591
rect 2631 1582 2635 1583
rect 2631 1577 2635 1578
rect 2687 1582 2691 1583
rect 2687 1577 2691 1578
rect 2688 1561 2690 1577
rect 2686 1560 2692 1561
rect 2686 1556 2687 1560
rect 2691 1556 2692 1560
rect 2686 1555 2692 1556
rect 2694 1522 2700 1523
rect 2694 1518 2695 1522
rect 2699 1518 2700 1522
rect 2694 1517 2700 1518
rect 2546 1511 2552 1512
rect 2546 1507 2547 1511
rect 2551 1507 2552 1511
rect 2546 1506 2552 1507
rect 2696 1499 2698 1517
rect 2724 1512 2726 1590
rect 2776 1583 2778 1607
rect 2920 1583 2922 1607
rect 3064 1583 3066 1607
rect 2775 1582 2779 1583
rect 2775 1577 2779 1578
rect 2839 1582 2843 1583
rect 2839 1577 2843 1578
rect 2919 1582 2923 1583
rect 2919 1577 2923 1578
rect 2983 1582 2987 1583
rect 2983 1577 2987 1578
rect 3063 1582 3067 1583
rect 3063 1577 3067 1578
rect 3119 1582 3123 1583
rect 3119 1577 3123 1578
rect 2840 1561 2842 1577
rect 2984 1561 2986 1577
rect 3120 1561 3122 1577
rect 2838 1560 2844 1561
rect 2838 1556 2839 1560
rect 2843 1556 2844 1560
rect 2838 1555 2844 1556
rect 2982 1560 2988 1561
rect 2982 1556 2983 1560
rect 2987 1556 2988 1560
rect 2982 1555 2988 1556
rect 3118 1560 3124 1561
rect 3118 1556 3119 1560
rect 3123 1556 3124 1560
rect 3118 1555 3124 1556
rect 2754 1551 2760 1552
rect 2754 1547 2755 1551
rect 2759 1547 2760 1551
rect 2754 1546 2760 1547
rect 2930 1551 2936 1552
rect 2930 1547 2931 1551
rect 2935 1547 2936 1551
rect 2930 1546 2936 1547
rect 3054 1551 3060 1552
rect 3054 1547 3055 1551
rect 3059 1547 3060 1551
rect 3054 1546 3060 1547
rect 2756 1512 2758 1546
rect 2846 1522 2852 1523
rect 2846 1518 2847 1522
rect 2851 1518 2852 1522
rect 2846 1517 2852 1518
rect 2722 1511 2728 1512
rect 2722 1507 2723 1511
rect 2727 1507 2728 1511
rect 2722 1506 2728 1507
rect 2754 1511 2760 1512
rect 2754 1507 2755 1511
rect 2759 1507 2760 1511
rect 2754 1506 2760 1507
rect 2848 1499 2850 1517
rect 2932 1512 2934 1546
rect 2990 1522 2996 1523
rect 2990 1518 2991 1522
rect 2995 1518 2996 1522
rect 2990 1517 2996 1518
rect 2930 1511 2936 1512
rect 2930 1507 2931 1511
rect 2935 1507 2936 1511
rect 2930 1506 2936 1507
rect 2992 1499 2994 1517
rect 2535 1498 2539 1499
rect 2535 1493 2539 1494
rect 2567 1498 2571 1499
rect 2567 1493 2571 1494
rect 2695 1498 2699 1499
rect 2695 1493 2699 1494
rect 2719 1498 2723 1499
rect 2719 1493 2723 1494
rect 2847 1498 2851 1499
rect 2847 1493 2851 1494
rect 2879 1498 2883 1499
rect 2879 1493 2883 1494
rect 2991 1498 2995 1499
rect 2991 1493 2995 1494
rect 3039 1498 3043 1499
rect 3039 1493 3043 1494
rect 2422 1491 2428 1492
rect 2422 1487 2423 1491
rect 2427 1487 2428 1491
rect 2422 1486 2428 1487
rect 2442 1491 2448 1492
rect 2442 1487 2443 1491
rect 2447 1487 2448 1491
rect 2442 1486 2448 1487
rect 2270 1482 2276 1483
rect 2270 1478 2271 1482
rect 2275 1478 2276 1482
rect 2270 1477 2276 1478
rect 2414 1482 2420 1483
rect 2414 1478 2415 1482
rect 2419 1478 2420 1482
rect 2414 1477 2420 1478
rect 2424 1456 2426 1486
rect 2568 1483 2570 1493
rect 2720 1483 2722 1493
rect 2726 1491 2732 1492
rect 2726 1487 2727 1491
rect 2731 1487 2732 1491
rect 2726 1486 2732 1487
rect 2566 1482 2572 1483
rect 2566 1478 2567 1482
rect 2571 1478 2572 1482
rect 2566 1477 2572 1478
rect 2718 1482 2724 1483
rect 2718 1478 2719 1482
rect 2723 1478 2724 1482
rect 2718 1477 2724 1478
rect 2728 1456 2730 1486
rect 2880 1483 2882 1493
rect 2886 1491 2892 1492
rect 2886 1487 2887 1491
rect 2891 1487 2892 1491
rect 2886 1486 2892 1487
rect 2878 1482 2884 1483
rect 2878 1478 2879 1482
rect 2883 1478 2884 1482
rect 2878 1477 2884 1478
rect 2888 1456 2890 1486
rect 3040 1483 3042 1493
rect 3056 1492 3058 1546
rect 3180 1544 3182 1654
rect 3224 1651 3226 1661
rect 3330 1659 3336 1660
rect 3330 1655 3331 1659
rect 3335 1655 3336 1659
rect 3330 1654 3336 1655
rect 3222 1650 3228 1651
rect 3222 1646 3223 1650
rect 3227 1646 3228 1650
rect 3222 1645 3228 1646
rect 3332 1624 3334 1654
rect 3376 1651 3378 1661
rect 3374 1650 3380 1651
rect 3374 1646 3375 1650
rect 3379 1646 3380 1650
rect 3374 1645 3380 1646
rect 3384 1624 3386 1670
rect 3400 1667 3402 1681
rect 3428 1676 3430 1750
rect 3464 1747 3466 1767
rect 3592 1747 3594 1770
rect 3463 1746 3467 1747
rect 3463 1741 3467 1742
rect 3503 1746 3507 1747
rect 3503 1741 3507 1742
rect 3591 1746 3595 1747
rect 3591 1741 3595 1742
rect 3504 1725 3506 1741
rect 3502 1724 3508 1725
rect 3502 1720 3503 1724
rect 3507 1720 3508 1724
rect 3592 1722 3594 1741
rect 3502 1719 3508 1720
rect 3590 1721 3596 1722
rect 3590 1717 3591 1721
rect 3595 1717 3596 1721
rect 3590 1716 3596 1717
rect 3458 1715 3464 1716
rect 3458 1711 3459 1715
rect 3463 1711 3464 1715
rect 3458 1710 3464 1711
rect 3460 1676 3462 1710
rect 3562 1707 3568 1708
rect 3562 1703 3563 1707
rect 3567 1703 3568 1707
rect 3562 1702 3568 1703
rect 3590 1704 3596 1705
rect 3510 1686 3516 1687
rect 3510 1682 3511 1686
rect 3515 1682 3516 1686
rect 3510 1681 3516 1682
rect 3426 1675 3432 1676
rect 3426 1671 3427 1675
rect 3431 1671 3432 1675
rect 3426 1670 3432 1671
rect 3458 1675 3464 1676
rect 3458 1671 3459 1675
rect 3463 1671 3464 1675
rect 3458 1670 3464 1671
rect 3512 1667 3514 1681
rect 3399 1666 3403 1667
rect 3399 1661 3403 1662
rect 3511 1666 3515 1667
rect 3511 1661 3515 1662
rect 3512 1651 3514 1661
rect 3564 1660 3566 1702
rect 3590 1700 3591 1704
rect 3595 1700 3596 1704
rect 3590 1699 3596 1700
rect 3592 1667 3594 1699
rect 3591 1666 3595 1667
rect 3591 1661 3595 1662
rect 3562 1659 3568 1660
rect 3562 1655 3563 1659
rect 3567 1655 3568 1659
rect 3562 1654 3568 1655
rect 3510 1650 3516 1651
rect 3510 1646 3511 1650
rect 3515 1646 3516 1650
rect 3510 1645 3516 1646
rect 3592 1633 3594 1661
rect 3590 1632 3596 1633
rect 3590 1628 3591 1632
rect 3595 1628 3596 1632
rect 3590 1627 3596 1628
rect 3330 1623 3336 1624
rect 3330 1619 3331 1623
rect 3335 1619 3336 1623
rect 3330 1618 3336 1619
rect 3382 1623 3388 1624
rect 3382 1619 3383 1623
rect 3387 1619 3388 1623
rect 3382 1618 3388 1619
rect 3534 1623 3540 1624
rect 3534 1619 3535 1623
rect 3539 1619 3540 1623
rect 3534 1618 3540 1619
rect 3214 1612 3220 1613
rect 3214 1608 3215 1612
rect 3219 1608 3220 1612
rect 3214 1607 3220 1608
rect 3366 1612 3372 1613
rect 3366 1608 3367 1612
rect 3371 1608 3372 1612
rect 3366 1607 3372 1608
rect 3502 1612 3508 1613
rect 3502 1608 3503 1612
rect 3507 1608 3508 1612
rect 3502 1607 3508 1608
rect 3216 1583 3218 1607
rect 3368 1583 3370 1607
rect 3504 1583 3506 1607
rect 3215 1582 3219 1583
rect 3215 1577 3219 1578
rect 3255 1582 3259 1583
rect 3255 1577 3259 1578
rect 3367 1582 3371 1583
rect 3367 1577 3371 1578
rect 3391 1582 3395 1583
rect 3391 1577 3395 1578
rect 3503 1582 3507 1583
rect 3503 1577 3507 1578
rect 3256 1561 3258 1577
rect 3392 1561 3394 1577
rect 3504 1561 3506 1577
rect 3254 1560 3260 1561
rect 3254 1556 3255 1560
rect 3259 1556 3260 1560
rect 3254 1555 3260 1556
rect 3390 1560 3396 1561
rect 3390 1556 3391 1560
rect 3395 1556 3396 1560
rect 3390 1555 3396 1556
rect 3502 1560 3508 1561
rect 3502 1556 3503 1560
rect 3507 1556 3508 1560
rect 3502 1555 3508 1556
rect 3186 1551 3192 1552
rect 3186 1547 3187 1551
rect 3191 1547 3192 1551
rect 3186 1546 3192 1547
rect 3322 1551 3328 1552
rect 3322 1547 3323 1551
rect 3327 1547 3328 1551
rect 3322 1546 3328 1547
rect 3178 1543 3184 1544
rect 3178 1539 3179 1543
rect 3183 1539 3184 1543
rect 3178 1538 3184 1539
rect 3126 1522 3132 1523
rect 3126 1518 3127 1522
rect 3131 1518 3132 1522
rect 3126 1517 3132 1518
rect 3128 1499 3130 1517
rect 3188 1512 3190 1546
rect 3262 1522 3268 1523
rect 3262 1518 3263 1522
rect 3267 1518 3268 1522
rect 3262 1517 3268 1518
rect 3186 1511 3192 1512
rect 3186 1507 3187 1511
rect 3191 1507 3192 1511
rect 3186 1506 3192 1507
rect 3264 1499 3266 1517
rect 3324 1512 3326 1546
rect 3398 1522 3404 1523
rect 3398 1518 3399 1522
rect 3403 1518 3404 1522
rect 3398 1517 3404 1518
rect 3510 1522 3516 1523
rect 3510 1518 3511 1522
rect 3515 1518 3516 1522
rect 3510 1517 3516 1518
rect 3322 1511 3328 1512
rect 3322 1507 3323 1511
rect 3327 1507 3328 1511
rect 3322 1506 3328 1507
rect 3400 1499 3402 1517
rect 3418 1511 3424 1512
rect 3418 1507 3419 1511
rect 3423 1507 3424 1511
rect 3418 1506 3424 1507
rect 3127 1498 3131 1499
rect 3127 1493 3131 1494
rect 3199 1498 3203 1499
rect 3199 1493 3203 1494
rect 3263 1498 3267 1499
rect 3263 1493 3267 1494
rect 3367 1498 3371 1499
rect 3367 1493 3371 1494
rect 3399 1498 3403 1499
rect 3399 1493 3403 1494
rect 3046 1491 3052 1492
rect 3046 1487 3047 1491
rect 3051 1487 3052 1491
rect 3046 1486 3052 1487
rect 3054 1491 3060 1492
rect 3054 1487 3055 1491
rect 3059 1487 3060 1491
rect 3054 1486 3060 1487
rect 3038 1482 3044 1483
rect 3038 1478 3039 1482
rect 3043 1478 3044 1482
rect 3038 1477 3044 1478
rect 3048 1456 3050 1486
rect 3200 1483 3202 1493
rect 3250 1491 3256 1492
rect 3250 1487 3251 1491
rect 3255 1487 3256 1491
rect 3250 1486 3256 1487
rect 3198 1482 3204 1483
rect 3198 1478 3199 1482
rect 3203 1478 3204 1482
rect 3198 1477 3204 1478
rect 3252 1456 3254 1486
rect 3368 1483 3370 1493
rect 3366 1482 3372 1483
rect 3366 1478 3367 1482
rect 3371 1478 3372 1482
rect 3366 1477 3372 1478
rect 3420 1456 3422 1506
rect 3512 1499 3514 1517
rect 3536 1512 3538 1618
rect 3590 1615 3596 1616
rect 3590 1611 3591 1615
rect 3595 1611 3596 1615
rect 3590 1610 3596 1611
rect 3592 1583 3594 1610
rect 3591 1582 3595 1583
rect 3591 1577 3595 1578
rect 3592 1558 3594 1577
rect 3590 1557 3596 1558
rect 3590 1553 3591 1557
rect 3595 1553 3596 1557
rect 3590 1552 3596 1553
rect 3562 1543 3568 1544
rect 3562 1539 3563 1543
rect 3567 1539 3568 1543
rect 3562 1538 3568 1539
rect 3590 1540 3596 1541
rect 3534 1511 3540 1512
rect 3534 1507 3535 1511
rect 3539 1507 3540 1511
rect 3534 1506 3540 1507
rect 3518 1499 3524 1500
rect 3511 1498 3515 1499
rect 3518 1495 3519 1499
rect 3523 1495 3524 1499
rect 3518 1494 3524 1495
rect 3511 1493 3515 1494
rect 3512 1483 3514 1493
rect 3510 1482 3516 1483
rect 3510 1478 3511 1482
rect 3515 1478 3516 1482
rect 3510 1477 3516 1478
rect 3520 1456 3522 1494
rect 3564 1492 3566 1538
rect 3590 1536 3591 1540
rect 3595 1536 3596 1540
rect 3590 1535 3596 1536
rect 3592 1499 3594 1535
rect 3591 1498 3595 1499
rect 3591 1493 3595 1494
rect 3562 1491 3568 1492
rect 3562 1487 3563 1491
rect 3567 1487 3568 1491
rect 3562 1486 3568 1487
rect 3592 1465 3594 1493
rect 3590 1464 3596 1465
rect 3590 1460 3591 1464
rect 3595 1460 3596 1464
rect 3590 1459 3596 1460
rect 1970 1455 1976 1456
rect 1970 1451 1971 1455
rect 1975 1451 1976 1455
rect 1970 1450 1976 1451
rect 2126 1455 2132 1456
rect 2126 1451 2127 1455
rect 2131 1451 2132 1455
rect 2126 1450 2132 1451
rect 2186 1455 2192 1456
rect 2186 1451 2187 1455
rect 2191 1451 2192 1455
rect 2186 1450 2192 1451
rect 2422 1455 2428 1456
rect 2422 1451 2423 1455
rect 2427 1451 2428 1455
rect 2422 1450 2428 1451
rect 2726 1455 2732 1456
rect 2726 1451 2727 1455
rect 2731 1451 2732 1455
rect 2726 1450 2732 1451
rect 2886 1455 2892 1456
rect 2886 1451 2887 1455
rect 2891 1451 2892 1455
rect 2886 1450 2892 1451
rect 3046 1455 3052 1456
rect 3046 1451 3047 1455
rect 3051 1451 3052 1455
rect 3046 1450 3052 1451
rect 3250 1455 3256 1456
rect 3250 1451 3251 1455
rect 3255 1451 3256 1455
rect 3250 1450 3256 1451
rect 3418 1455 3424 1456
rect 3418 1451 3419 1455
rect 3423 1451 3424 1455
rect 3418 1450 3424 1451
rect 3518 1455 3524 1456
rect 3518 1451 3519 1455
rect 3523 1451 3524 1455
rect 3518 1450 3524 1451
rect 3590 1447 3596 1448
rect 1998 1444 2004 1445
rect 1998 1440 1999 1444
rect 2003 1440 2004 1444
rect 1998 1439 2004 1440
rect 2126 1444 2132 1445
rect 2126 1440 2127 1444
rect 2131 1440 2132 1444
rect 2126 1439 2132 1440
rect 2262 1444 2268 1445
rect 2262 1440 2263 1444
rect 2267 1440 2268 1444
rect 2262 1439 2268 1440
rect 2406 1444 2412 1445
rect 2406 1440 2407 1444
rect 2411 1440 2412 1444
rect 2406 1439 2412 1440
rect 2558 1444 2564 1445
rect 2558 1440 2559 1444
rect 2563 1440 2564 1444
rect 2558 1439 2564 1440
rect 2710 1444 2716 1445
rect 2710 1440 2711 1444
rect 2715 1440 2716 1444
rect 2710 1439 2716 1440
rect 2870 1444 2876 1445
rect 2870 1440 2871 1444
rect 2875 1440 2876 1444
rect 2870 1439 2876 1440
rect 3030 1444 3036 1445
rect 3030 1440 3031 1444
rect 3035 1440 3036 1444
rect 3030 1439 3036 1440
rect 3190 1444 3196 1445
rect 3190 1440 3191 1444
rect 3195 1440 3196 1444
rect 3190 1439 3196 1440
rect 3358 1444 3364 1445
rect 3358 1440 3359 1444
rect 3363 1440 3364 1444
rect 3358 1439 3364 1440
rect 3502 1444 3508 1445
rect 3502 1440 3503 1444
rect 3507 1440 3508 1444
rect 3590 1443 3591 1447
rect 3595 1443 3596 1447
rect 3590 1442 3596 1443
rect 3502 1439 3508 1440
rect 2000 1423 2002 1439
rect 2058 1427 2064 1428
rect 2058 1423 2059 1427
rect 2063 1423 2064 1427
rect 2128 1423 2130 1439
rect 2264 1423 2266 1439
rect 2408 1423 2410 1439
rect 2466 1427 2472 1428
rect 2466 1423 2467 1427
rect 2471 1423 2472 1427
rect 2560 1423 2562 1439
rect 2712 1423 2714 1439
rect 2872 1423 2874 1439
rect 3032 1423 3034 1439
rect 3192 1423 3194 1439
rect 3360 1423 3362 1439
rect 3504 1423 3506 1439
rect 3592 1423 3594 1442
rect 1999 1422 2003 1423
rect 1999 1417 2003 1418
rect 2023 1422 2027 1423
rect 2058 1422 2064 1423
rect 2127 1422 2131 1423
rect 2023 1417 2027 1418
rect 2024 1401 2026 1417
rect 2022 1400 2028 1401
rect 2022 1396 2023 1400
rect 2027 1396 2028 1400
rect 2022 1395 2028 1396
rect 1830 1391 1836 1392
rect 1962 1391 1968 1392
rect 1832 1363 1834 1391
rect 1962 1387 1963 1391
rect 1967 1387 1968 1391
rect 1962 1386 1968 1387
rect 1870 1380 1876 1381
rect 1870 1376 1871 1380
rect 1875 1376 1876 1380
rect 1870 1375 1876 1376
rect 1831 1362 1835 1363
rect 1831 1357 1835 1358
rect 1810 1351 1816 1352
rect 1810 1347 1811 1351
rect 1815 1347 1816 1351
rect 1810 1346 1816 1347
rect 1832 1329 1834 1357
rect 1872 1339 1874 1375
rect 1902 1362 1908 1363
rect 1902 1358 1903 1362
rect 1907 1358 1908 1362
rect 1902 1357 1908 1358
rect 2030 1362 2036 1363
rect 2030 1358 2031 1362
rect 2035 1358 2036 1362
rect 2030 1357 2036 1358
rect 1904 1339 1906 1357
rect 2032 1339 2034 1357
rect 2060 1352 2062 1422
rect 2127 1417 2131 1418
rect 2167 1422 2171 1423
rect 2167 1417 2171 1418
rect 2263 1422 2267 1423
rect 2263 1417 2267 1418
rect 2303 1422 2307 1423
rect 2303 1417 2307 1418
rect 2407 1422 2411 1423
rect 2407 1417 2411 1418
rect 2431 1422 2435 1423
rect 2466 1422 2472 1423
rect 2551 1422 2555 1423
rect 2431 1417 2435 1418
rect 2168 1401 2170 1417
rect 2304 1401 2306 1417
rect 2432 1401 2434 1417
rect 2166 1400 2172 1401
rect 2166 1396 2167 1400
rect 2171 1396 2172 1400
rect 2166 1395 2172 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2430 1400 2436 1401
rect 2430 1396 2431 1400
rect 2435 1396 2436 1400
rect 2430 1395 2436 1396
rect 2114 1391 2120 1392
rect 2114 1387 2115 1391
rect 2119 1387 2120 1391
rect 2114 1386 2120 1387
rect 2258 1391 2264 1392
rect 2258 1387 2259 1391
rect 2263 1387 2264 1391
rect 2258 1386 2264 1387
rect 2378 1391 2384 1392
rect 2378 1387 2379 1391
rect 2383 1387 2384 1391
rect 2378 1386 2384 1387
rect 2116 1352 2118 1386
rect 2174 1362 2180 1363
rect 2174 1358 2175 1362
rect 2179 1358 2180 1362
rect 2174 1357 2180 1358
rect 2058 1351 2064 1352
rect 2058 1347 2059 1351
rect 2063 1347 2064 1351
rect 2058 1346 2064 1347
rect 2114 1351 2120 1352
rect 2114 1347 2115 1351
rect 2119 1347 2120 1351
rect 2114 1346 2120 1347
rect 2176 1339 2178 1357
rect 2260 1352 2262 1386
rect 2310 1362 2316 1363
rect 2310 1358 2311 1362
rect 2315 1358 2316 1362
rect 2310 1357 2316 1358
rect 2258 1351 2264 1352
rect 2258 1347 2259 1351
rect 2263 1347 2264 1351
rect 2258 1346 2264 1347
rect 2312 1339 2314 1357
rect 2380 1340 2382 1386
rect 2438 1362 2444 1363
rect 2438 1358 2439 1362
rect 2443 1358 2444 1362
rect 2438 1357 2444 1358
rect 2378 1339 2384 1340
rect 2440 1339 2442 1357
rect 2468 1352 2470 1422
rect 2551 1417 2555 1418
rect 2559 1422 2563 1423
rect 2559 1417 2563 1418
rect 2671 1422 2675 1423
rect 2671 1417 2675 1418
rect 2711 1422 2715 1423
rect 2711 1417 2715 1418
rect 2791 1422 2795 1423
rect 2791 1417 2795 1418
rect 2871 1422 2875 1423
rect 2871 1417 2875 1418
rect 2911 1422 2915 1423
rect 2911 1417 2915 1418
rect 3031 1422 3035 1423
rect 3031 1417 3035 1418
rect 3191 1422 3195 1423
rect 3191 1417 3195 1418
rect 3359 1422 3363 1423
rect 3359 1417 3363 1418
rect 3503 1422 3507 1423
rect 3503 1417 3507 1418
rect 3591 1422 3595 1423
rect 3591 1417 3595 1418
rect 2552 1401 2554 1417
rect 2672 1401 2674 1417
rect 2792 1401 2794 1417
rect 2912 1401 2914 1417
rect 2550 1400 2556 1401
rect 2550 1396 2551 1400
rect 2555 1396 2556 1400
rect 2550 1395 2556 1396
rect 2670 1400 2676 1401
rect 2670 1396 2671 1400
rect 2675 1396 2676 1400
rect 2670 1395 2676 1396
rect 2790 1400 2796 1401
rect 2790 1396 2791 1400
rect 2795 1396 2796 1400
rect 2790 1395 2796 1396
rect 2910 1400 2916 1401
rect 2910 1396 2911 1400
rect 2915 1396 2916 1400
rect 3592 1398 3594 1417
rect 2910 1395 2916 1396
rect 3590 1397 3596 1398
rect 3590 1393 3591 1397
rect 3595 1393 3596 1397
rect 3590 1392 3596 1393
rect 2514 1391 2520 1392
rect 2514 1387 2515 1391
rect 2519 1387 2520 1391
rect 2514 1386 2520 1387
rect 2634 1391 2640 1392
rect 2634 1387 2635 1391
rect 2639 1387 2640 1391
rect 2634 1386 2640 1387
rect 2754 1391 2760 1392
rect 2754 1387 2755 1391
rect 2759 1387 2760 1391
rect 2754 1386 2760 1387
rect 2866 1391 2872 1392
rect 2866 1387 2867 1391
rect 2871 1387 2872 1391
rect 2866 1386 2872 1387
rect 2874 1391 2880 1392
rect 2874 1387 2875 1391
rect 2879 1387 2880 1391
rect 2874 1386 2880 1387
rect 2516 1352 2518 1386
rect 2558 1362 2564 1363
rect 2558 1358 2559 1362
rect 2563 1358 2564 1362
rect 2558 1357 2564 1358
rect 2466 1351 2472 1352
rect 2466 1347 2467 1351
rect 2471 1347 2472 1351
rect 2466 1346 2472 1347
rect 2514 1351 2520 1352
rect 2514 1347 2515 1351
rect 2519 1347 2520 1351
rect 2514 1346 2520 1347
rect 2560 1339 2562 1357
rect 2636 1352 2638 1386
rect 2678 1362 2684 1363
rect 2678 1358 2679 1362
rect 2683 1358 2684 1362
rect 2678 1357 2684 1358
rect 2634 1351 2640 1352
rect 2619 1348 2623 1349
rect 2634 1347 2635 1351
rect 2639 1347 2640 1351
rect 2634 1346 2640 1347
rect 2619 1343 2623 1344
rect 1871 1338 1875 1339
rect 1871 1333 1875 1334
rect 1903 1338 1907 1339
rect 1903 1333 1907 1334
rect 1927 1338 1931 1339
rect 1927 1333 1931 1334
rect 2031 1338 2035 1339
rect 2031 1333 2035 1334
rect 2047 1338 2051 1339
rect 2047 1333 2051 1334
rect 2175 1338 2179 1339
rect 2175 1333 2179 1334
rect 2183 1338 2187 1339
rect 2183 1333 2187 1334
rect 2311 1338 2315 1339
rect 2311 1333 2315 1334
rect 2319 1338 2323 1339
rect 2378 1335 2379 1339
rect 2383 1335 2384 1339
rect 2378 1334 2384 1335
rect 2439 1338 2443 1339
rect 2319 1333 2323 1334
rect 2439 1333 2443 1334
rect 2455 1338 2459 1339
rect 2455 1333 2459 1334
rect 2559 1338 2563 1339
rect 2559 1333 2563 1334
rect 2591 1338 2595 1339
rect 2591 1333 2595 1334
rect 1830 1328 1836 1329
rect 1830 1324 1831 1328
rect 1835 1324 1836 1328
rect 1830 1323 1836 1324
rect 1330 1319 1336 1320
rect 1330 1315 1331 1319
rect 1335 1315 1336 1319
rect 1330 1314 1336 1315
rect 1458 1319 1464 1320
rect 1458 1315 1459 1319
rect 1463 1315 1464 1319
rect 1458 1314 1464 1315
rect 1698 1319 1704 1320
rect 1698 1315 1699 1319
rect 1703 1315 1704 1319
rect 1698 1314 1704 1315
rect 1774 1319 1780 1320
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1774 1314 1780 1315
rect 1830 1311 1836 1312
rect 1398 1308 1404 1309
rect 1398 1304 1399 1308
rect 1403 1304 1404 1308
rect 1398 1303 1404 1304
rect 1518 1308 1524 1309
rect 1518 1304 1519 1308
rect 1523 1304 1524 1308
rect 1518 1303 1524 1304
rect 1638 1308 1644 1309
rect 1638 1304 1639 1308
rect 1643 1304 1644 1308
rect 1638 1303 1644 1304
rect 1742 1308 1748 1309
rect 1742 1304 1743 1308
rect 1747 1304 1748 1308
rect 1830 1307 1831 1311
rect 1835 1307 1836 1311
rect 1830 1306 1836 1307
rect 1742 1303 1748 1304
rect 1307 1300 1311 1301
rect 1307 1295 1311 1296
rect 1400 1283 1402 1303
rect 1520 1283 1522 1303
rect 1599 1300 1603 1301
rect 1599 1295 1603 1296
rect 1239 1282 1243 1283
rect 1239 1277 1243 1278
rect 1271 1282 1275 1283
rect 1271 1277 1275 1278
rect 1375 1282 1379 1283
rect 1375 1277 1379 1278
rect 1399 1282 1403 1283
rect 1399 1277 1403 1278
rect 1503 1282 1507 1283
rect 1503 1277 1507 1278
rect 1519 1282 1523 1283
rect 1519 1277 1523 1278
rect 1240 1261 1242 1277
rect 1376 1261 1378 1277
rect 1504 1261 1506 1277
rect 1238 1260 1244 1261
rect 1238 1256 1239 1260
rect 1243 1256 1244 1260
rect 1238 1255 1244 1256
rect 1374 1260 1380 1261
rect 1374 1256 1375 1260
rect 1379 1256 1380 1260
rect 1374 1255 1380 1256
rect 1502 1260 1508 1261
rect 1502 1256 1503 1260
rect 1507 1256 1508 1260
rect 1502 1255 1508 1256
rect 1600 1252 1602 1295
rect 1640 1283 1642 1303
rect 1744 1283 1746 1303
rect 1832 1283 1834 1306
rect 1872 1305 1874 1333
rect 1928 1323 1930 1333
rect 1978 1331 1984 1332
rect 1978 1327 1979 1331
rect 1983 1327 1984 1331
rect 1978 1326 1984 1327
rect 1926 1322 1932 1323
rect 1926 1318 1927 1322
rect 1931 1318 1932 1322
rect 1926 1317 1932 1318
rect 1870 1304 1876 1305
rect 1870 1300 1871 1304
rect 1875 1300 1876 1304
rect 1870 1299 1876 1300
rect 1980 1296 1982 1326
rect 1987 1324 1991 1325
rect 1986 1319 1987 1324
rect 1991 1319 1992 1324
rect 2048 1323 2050 1333
rect 2098 1331 2104 1332
rect 2098 1327 2099 1331
rect 2103 1327 2104 1331
rect 2098 1326 2104 1327
rect 1986 1318 1992 1319
rect 2046 1322 2052 1323
rect 2046 1318 2047 1322
rect 2051 1318 2052 1322
rect 2046 1317 2052 1318
rect 2100 1296 2102 1326
rect 2184 1323 2186 1333
rect 2320 1323 2322 1333
rect 2327 1324 2331 1325
rect 2182 1322 2188 1323
rect 2182 1318 2183 1322
rect 2187 1318 2188 1322
rect 2182 1317 2188 1318
rect 2318 1322 2324 1323
rect 2318 1318 2319 1322
rect 2323 1318 2324 1322
rect 2456 1323 2458 1333
rect 2462 1331 2468 1332
rect 2462 1327 2463 1331
rect 2467 1327 2468 1331
rect 2462 1326 2468 1327
rect 2327 1319 2331 1320
rect 2454 1322 2460 1323
rect 2318 1317 2324 1318
rect 2328 1296 2330 1319
rect 2454 1318 2455 1322
rect 2459 1318 2460 1322
rect 2454 1317 2460 1318
rect 2464 1296 2466 1326
rect 2592 1323 2594 1333
rect 2620 1332 2622 1343
rect 2680 1339 2682 1357
rect 2756 1352 2758 1386
rect 2798 1362 2804 1363
rect 2798 1358 2799 1362
rect 2803 1358 2804 1362
rect 2798 1357 2804 1358
rect 2754 1351 2760 1352
rect 2754 1347 2755 1351
rect 2759 1347 2760 1351
rect 2754 1346 2760 1347
rect 2800 1339 2802 1357
rect 2868 1352 2870 1386
rect 2866 1351 2872 1352
rect 2866 1347 2867 1351
rect 2871 1347 2872 1351
rect 2876 1349 2878 1386
rect 3590 1380 3596 1381
rect 3590 1376 3591 1380
rect 3595 1376 3596 1380
rect 3590 1375 3596 1376
rect 2918 1362 2924 1363
rect 2918 1358 2919 1362
rect 2923 1358 2924 1362
rect 2918 1357 2924 1358
rect 2866 1346 2872 1347
rect 2875 1348 2879 1349
rect 2875 1343 2879 1344
rect 2920 1339 2922 1357
rect 3592 1339 3594 1375
rect 2679 1338 2683 1339
rect 2679 1333 2683 1334
rect 2719 1338 2723 1339
rect 2719 1333 2723 1334
rect 2799 1338 2803 1339
rect 2799 1333 2803 1334
rect 2839 1338 2843 1339
rect 2839 1333 2843 1334
rect 2919 1338 2923 1339
rect 2919 1333 2923 1334
rect 2951 1338 2955 1339
rect 2951 1333 2955 1334
rect 3063 1338 3067 1339
rect 3063 1333 3067 1334
rect 3183 1338 3187 1339
rect 3183 1333 3187 1334
rect 3591 1338 3595 1339
rect 3591 1333 3595 1334
rect 2618 1331 2624 1332
rect 2618 1327 2619 1331
rect 2623 1327 2624 1331
rect 2618 1326 2624 1327
rect 2642 1331 2648 1332
rect 2642 1327 2643 1331
rect 2647 1327 2648 1331
rect 2642 1326 2648 1327
rect 2590 1322 2596 1323
rect 2590 1318 2591 1322
rect 2595 1318 2596 1322
rect 2590 1317 2596 1318
rect 2644 1296 2646 1326
rect 2720 1323 2722 1333
rect 2770 1331 2776 1332
rect 2770 1327 2771 1331
rect 2775 1327 2776 1331
rect 2770 1326 2776 1327
rect 2718 1322 2724 1323
rect 2718 1318 2719 1322
rect 2723 1318 2724 1322
rect 2718 1317 2724 1318
rect 2772 1296 2774 1326
rect 2840 1323 2842 1333
rect 2890 1331 2896 1332
rect 2890 1327 2891 1331
rect 2895 1327 2896 1331
rect 2890 1326 2896 1327
rect 2838 1322 2844 1323
rect 2838 1318 2839 1322
rect 2843 1318 2844 1322
rect 2838 1317 2844 1318
rect 2892 1296 2894 1326
rect 2952 1323 2954 1333
rect 3002 1331 3008 1332
rect 3002 1327 3003 1331
rect 3007 1327 3008 1331
rect 3002 1326 3008 1327
rect 2950 1322 2956 1323
rect 2950 1318 2951 1322
rect 2955 1318 2956 1322
rect 2950 1317 2956 1318
rect 3004 1296 3006 1326
rect 3064 1323 3066 1333
rect 3114 1331 3120 1332
rect 3114 1327 3115 1331
rect 3119 1327 3120 1331
rect 3114 1326 3120 1327
rect 3062 1322 3068 1323
rect 3062 1318 3063 1322
rect 3067 1318 3068 1322
rect 3062 1317 3068 1318
rect 3116 1296 3118 1326
rect 3184 1323 3186 1333
rect 3182 1322 3188 1323
rect 3182 1318 3183 1322
rect 3187 1318 3188 1322
rect 3182 1317 3188 1318
rect 3592 1305 3594 1333
rect 3590 1304 3596 1305
rect 3590 1300 3591 1304
rect 3595 1300 3596 1304
rect 3590 1299 3596 1300
rect 1978 1295 1984 1296
rect 1978 1291 1979 1295
rect 1983 1291 1984 1295
rect 1978 1290 1984 1291
rect 2098 1295 2104 1296
rect 2098 1291 2099 1295
rect 2103 1291 2104 1295
rect 2098 1290 2104 1291
rect 2234 1295 2240 1296
rect 2234 1291 2235 1295
rect 2239 1291 2240 1295
rect 2234 1290 2240 1291
rect 2326 1295 2332 1296
rect 2326 1291 2327 1295
rect 2331 1291 2332 1295
rect 2326 1290 2332 1291
rect 2462 1295 2468 1296
rect 2462 1291 2463 1295
rect 2467 1291 2468 1295
rect 2462 1290 2468 1291
rect 2642 1295 2648 1296
rect 2642 1291 2643 1295
rect 2647 1291 2648 1295
rect 2642 1290 2648 1291
rect 2770 1295 2776 1296
rect 2770 1291 2771 1295
rect 2775 1291 2776 1295
rect 2770 1290 2776 1291
rect 2890 1295 2896 1296
rect 2890 1291 2891 1295
rect 2895 1291 2896 1295
rect 2890 1290 2896 1291
rect 3002 1295 3008 1296
rect 3002 1291 3003 1295
rect 3007 1291 3008 1295
rect 3002 1290 3008 1291
rect 3114 1295 3120 1296
rect 3114 1291 3115 1295
rect 3119 1291 3120 1295
rect 3114 1290 3120 1291
rect 1870 1287 1876 1288
rect 1870 1283 1871 1287
rect 1875 1283 1876 1287
rect 1631 1282 1635 1283
rect 1631 1277 1635 1278
rect 1639 1282 1643 1283
rect 1639 1277 1643 1278
rect 1743 1282 1747 1283
rect 1743 1277 1747 1278
rect 1831 1282 1835 1283
rect 1870 1282 1876 1283
rect 1918 1284 1924 1285
rect 1831 1277 1835 1278
rect 1632 1261 1634 1277
rect 1744 1261 1746 1277
rect 1630 1260 1636 1261
rect 1630 1256 1631 1260
rect 1635 1256 1636 1260
rect 1630 1255 1636 1256
rect 1742 1260 1748 1261
rect 1742 1256 1743 1260
rect 1747 1256 1748 1260
rect 1832 1258 1834 1277
rect 1742 1255 1748 1256
rect 1830 1257 1836 1258
rect 1830 1253 1831 1257
rect 1835 1253 1836 1257
rect 1872 1255 1874 1282
rect 1918 1280 1919 1284
rect 1923 1280 1924 1284
rect 1918 1279 1924 1280
rect 2038 1284 2044 1285
rect 2038 1280 2039 1284
rect 2043 1280 2044 1284
rect 2038 1279 2044 1280
rect 2174 1284 2180 1285
rect 2174 1280 2175 1284
rect 2179 1280 2180 1284
rect 2174 1279 2180 1280
rect 1920 1255 1922 1279
rect 2040 1255 2042 1279
rect 2176 1255 2178 1279
rect 1830 1252 1836 1253
rect 1871 1254 1875 1255
rect 906 1251 912 1252
rect 906 1247 907 1251
rect 911 1247 912 1251
rect 906 1246 912 1247
rect 1050 1251 1056 1252
rect 1050 1247 1051 1251
rect 1055 1247 1056 1251
rect 1050 1246 1056 1247
rect 1170 1251 1176 1252
rect 1170 1247 1171 1251
rect 1175 1247 1176 1251
rect 1170 1246 1176 1247
rect 1330 1251 1336 1252
rect 1330 1247 1331 1251
rect 1335 1247 1336 1251
rect 1330 1246 1336 1247
rect 1462 1251 1468 1252
rect 1462 1247 1463 1251
rect 1467 1247 1468 1251
rect 1462 1246 1468 1247
rect 1590 1251 1596 1252
rect 1590 1247 1591 1251
rect 1595 1247 1596 1251
rect 1590 1246 1596 1247
rect 1598 1251 1604 1252
rect 1598 1247 1599 1251
rect 1603 1247 1604 1251
rect 1871 1249 1875 1250
rect 1895 1254 1899 1255
rect 1895 1249 1899 1250
rect 1919 1254 1923 1255
rect 1919 1249 1923 1250
rect 2039 1254 2043 1255
rect 2039 1249 2043 1250
rect 2071 1254 2075 1255
rect 2071 1249 2075 1250
rect 2175 1254 2179 1255
rect 2175 1249 2179 1250
rect 1598 1246 1604 1247
rect 822 1222 828 1223
rect 822 1218 823 1222
rect 827 1218 828 1222
rect 822 1217 828 1218
rect 706 1211 712 1212
rect 706 1207 707 1211
rect 711 1207 712 1211
rect 810 1211 816 1212
rect 810 1207 811 1211
rect 815 1207 816 1211
rect 824 1207 826 1217
rect 908 1212 910 1246
rect 966 1222 972 1223
rect 966 1218 967 1222
rect 971 1218 972 1222
rect 966 1217 972 1218
rect 906 1211 912 1212
rect 906 1207 907 1211
rect 911 1207 912 1211
rect 968 1207 970 1217
rect 1052 1212 1054 1246
rect 1110 1222 1116 1223
rect 1110 1218 1111 1222
rect 1115 1218 1116 1222
rect 1110 1217 1116 1218
rect 1246 1222 1252 1223
rect 1246 1218 1247 1222
rect 1251 1218 1252 1222
rect 1246 1217 1252 1218
rect 1050 1211 1056 1212
rect 1050 1207 1051 1211
rect 1055 1207 1056 1211
rect 1112 1207 1114 1217
rect 1248 1207 1250 1217
rect 1332 1212 1334 1246
rect 1382 1222 1388 1223
rect 1382 1218 1383 1222
rect 1387 1218 1388 1222
rect 1382 1217 1388 1218
rect 1330 1211 1336 1212
rect 1330 1207 1331 1211
rect 1335 1207 1336 1211
rect 1384 1207 1386 1217
rect 1464 1212 1466 1246
rect 1510 1222 1516 1223
rect 1510 1218 1511 1222
rect 1515 1218 1516 1222
rect 1510 1217 1516 1218
rect 1462 1211 1468 1212
rect 1462 1207 1463 1211
rect 1467 1207 1468 1211
rect 1512 1207 1514 1217
rect 1592 1212 1594 1246
rect 1802 1243 1808 1244
rect 1802 1239 1803 1243
rect 1807 1239 1808 1243
rect 1802 1238 1808 1239
rect 1830 1240 1836 1241
rect 1638 1222 1644 1223
rect 1638 1218 1639 1222
rect 1643 1218 1644 1222
rect 1638 1217 1644 1218
rect 1750 1222 1756 1223
rect 1750 1218 1751 1222
rect 1755 1218 1756 1222
rect 1750 1217 1756 1218
rect 1590 1211 1596 1212
rect 1590 1207 1591 1211
rect 1595 1207 1596 1211
rect 1640 1207 1642 1217
rect 1752 1207 1754 1217
rect 319 1206 323 1207
rect 378 1206 384 1207
rect 415 1206 419 1207
rect 319 1201 323 1202
rect 415 1201 419 1202
rect 423 1206 427 1207
rect 482 1206 488 1207
rect 543 1206 547 1207
rect 423 1201 427 1202
rect 543 1201 547 1202
rect 591 1206 595 1207
rect 602 1206 608 1207
rect 679 1206 683 1207
rect 706 1206 712 1207
rect 759 1206 763 1207
rect 810 1206 816 1207
rect 823 1206 827 1207
rect 906 1206 912 1207
rect 927 1206 931 1207
rect 591 1201 595 1202
rect 679 1201 683 1202
rect 759 1201 763 1202
rect 266 1199 272 1200
rect 266 1195 267 1199
rect 271 1195 272 1199
rect 266 1194 272 1195
rect 290 1199 296 1200
rect 290 1195 291 1199
rect 295 1195 296 1199
rect 290 1194 296 1195
rect 238 1190 244 1191
rect 238 1186 239 1190
rect 243 1186 244 1190
rect 238 1185 244 1186
rect 110 1172 116 1173
rect 110 1168 111 1172
rect 115 1168 116 1172
rect 110 1167 116 1168
rect 292 1164 294 1194
rect 416 1191 418 1201
rect 466 1199 472 1200
rect 466 1195 467 1199
rect 471 1195 472 1199
rect 466 1194 472 1195
rect 414 1190 420 1191
rect 414 1186 415 1190
rect 419 1186 420 1190
rect 414 1185 420 1186
rect 468 1164 470 1194
rect 592 1191 594 1201
rect 760 1191 762 1201
rect 590 1190 596 1191
rect 590 1186 591 1190
rect 595 1186 596 1190
rect 590 1185 596 1186
rect 758 1190 764 1191
rect 758 1186 759 1190
rect 763 1186 764 1190
rect 758 1185 764 1186
rect 812 1164 814 1206
rect 823 1201 827 1202
rect 927 1201 931 1202
rect 967 1206 971 1207
rect 1050 1206 1056 1207
rect 1079 1206 1083 1207
rect 967 1201 971 1202
rect 1079 1201 1083 1202
rect 1111 1206 1115 1207
rect 1111 1201 1115 1202
rect 1223 1206 1227 1207
rect 1223 1201 1227 1202
rect 1247 1206 1251 1207
rect 1330 1206 1336 1207
rect 1367 1206 1371 1207
rect 1247 1201 1251 1202
rect 1367 1201 1371 1202
rect 1383 1206 1387 1207
rect 1462 1206 1468 1207
rect 1503 1206 1507 1207
rect 1383 1201 1387 1202
rect 1503 1201 1507 1202
rect 1511 1206 1515 1207
rect 1590 1206 1596 1207
rect 1639 1206 1643 1207
rect 1511 1201 1515 1202
rect 1639 1201 1643 1202
rect 1751 1206 1755 1207
rect 1751 1201 1755 1202
rect 928 1191 930 1201
rect 934 1199 940 1200
rect 934 1195 935 1199
rect 939 1195 940 1199
rect 934 1194 940 1195
rect 942 1199 948 1200
rect 942 1195 943 1199
rect 947 1195 948 1199
rect 942 1194 948 1195
rect 926 1190 932 1191
rect 926 1186 927 1190
rect 931 1186 932 1190
rect 926 1185 932 1186
rect 936 1164 938 1194
rect 290 1163 296 1164
rect 290 1159 291 1163
rect 295 1159 296 1163
rect 290 1158 296 1159
rect 466 1163 472 1164
rect 466 1159 467 1163
rect 471 1159 472 1163
rect 466 1158 472 1159
rect 810 1163 816 1164
rect 810 1159 811 1163
rect 815 1159 816 1163
rect 810 1158 816 1159
rect 934 1163 940 1164
rect 934 1159 935 1163
rect 939 1159 940 1163
rect 934 1158 940 1159
rect 110 1155 116 1156
rect 110 1151 111 1155
rect 115 1151 116 1155
rect 110 1150 116 1151
rect 230 1152 236 1153
rect 112 1127 114 1150
rect 230 1148 231 1152
rect 235 1148 236 1152
rect 230 1147 236 1148
rect 406 1152 412 1153
rect 406 1148 407 1152
rect 411 1148 412 1152
rect 406 1147 412 1148
rect 582 1152 588 1153
rect 582 1148 583 1152
rect 587 1148 588 1152
rect 582 1147 588 1148
rect 750 1152 756 1153
rect 750 1148 751 1152
rect 755 1148 756 1152
rect 750 1147 756 1148
rect 918 1152 924 1153
rect 918 1148 919 1152
rect 923 1148 924 1152
rect 918 1147 924 1148
rect 232 1127 234 1147
rect 408 1127 410 1147
rect 458 1135 464 1136
rect 458 1131 459 1135
rect 463 1131 464 1135
rect 458 1130 464 1131
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 143 1126 147 1127
rect 143 1121 147 1122
rect 231 1126 235 1127
rect 231 1121 235 1122
rect 279 1126 283 1127
rect 279 1121 283 1122
rect 407 1126 411 1127
rect 407 1121 411 1122
rect 423 1126 427 1127
rect 423 1121 427 1122
rect 112 1102 114 1121
rect 144 1105 146 1121
rect 280 1105 282 1121
rect 424 1105 426 1121
rect 142 1104 148 1105
rect 110 1101 116 1102
rect 110 1097 111 1101
rect 115 1097 116 1101
rect 142 1100 143 1104
rect 147 1100 148 1104
rect 142 1099 148 1100
rect 278 1104 284 1105
rect 278 1100 279 1104
rect 283 1100 284 1104
rect 278 1099 284 1100
rect 422 1104 428 1105
rect 422 1100 423 1104
rect 427 1100 428 1104
rect 422 1099 428 1100
rect 110 1096 116 1097
rect 210 1095 216 1096
rect 210 1091 211 1095
rect 215 1091 216 1095
rect 210 1090 216 1091
rect 346 1095 352 1096
rect 346 1091 347 1095
rect 351 1091 352 1095
rect 346 1090 352 1091
rect 202 1087 208 1088
rect 110 1084 116 1085
rect 110 1080 111 1084
rect 115 1080 116 1084
rect 202 1083 203 1087
rect 207 1083 208 1087
rect 202 1082 208 1083
rect 110 1079 116 1080
rect 112 1043 114 1079
rect 150 1066 156 1067
rect 150 1062 151 1066
rect 155 1062 156 1066
rect 150 1061 156 1062
rect 152 1043 154 1061
rect 111 1042 115 1043
rect 111 1037 115 1038
rect 143 1042 147 1043
rect 143 1037 147 1038
rect 151 1042 155 1043
rect 151 1037 155 1038
rect 112 1009 114 1037
rect 144 1027 146 1037
rect 204 1036 206 1082
rect 212 1056 214 1090
rect 286 1066 292 1067
rect 286 1062 287 1066
rect 291 1062 292 1066
rect 286 1061 292 1062
rect 210 1055 216 1056
rect 210 1051 211 1055
rect 215 1051 216 1055
rect 210 1050 216 1051
rect 288 1043 290 1061
rect 348 1056 350 1090
rect 430 1066 436 1067
rect 430 1062 431 1066
rect 435 1062 436 1066
rect 430 1061 436 1062
rect 346 1055 352 1056
rect 346 1051 347 1055
rect 351 1051 352 1055
rect 346 1050 352 1051
rect 414 1043 420 1044
rect 432 1043 434 1061
rect 460 1056 462 1130
rect 584 1127 586 1147
rect 752 1127 754 1147
rect 920 1127 922 1147
rect 567 1126 571 1127
rect 567 1121 571 1122
rect 583 1126 587 1127
rect 583 1121 587 1122
rect 711 1126 715 1127
rect 711 1121 715 1122
rect 751 1126 755 1127
rect 751 1121 755 1122
rect 847 1126 851 1127
rect 847 1121 851 1122
rect 919 1126 923 1127
rect 919 1121 923 1122
rect 568 1105 570 1121
rect 712 1105 714 1121
rect 848 1105 850 1121
rect 566 1104 572 1105
rect 566 1100 567 1104
rect 571 1100 572 1104
rect 566 1099 572 1100
rect 710 1104 716 1105
rect 710 1100 711 1104
rect 715 1100 716 1104
rect 710 1099 716 1100
rect 846 1104 852 1105
rect 846 1100 847 1104
rect 851 1100 852 1104
rect 846 1099 852 1100
rect 944 1096 946 1194
rect 1080 1191 1082 1201
rect 1122 1199 1128 1200
rect 1122 1195 1123 1199
rect 1127 1195 1128 1199
rect 1122 1194 1128 1195
rect 1130 1199 1136 1200
rect 1130 1195 1131 1199
rect 1135 1195 1136 1199
rect 1130 1194 1136 1195
rect 1078 1190 1084 1191
rect 1078 1186 1079 1190
rect 1083 1186 1084 1190
rect 1078 1185 1084 1186
rect 1070 1152 1076 1153
rect 1070 1148 1071 1152
rect 1075 1148 1076 1152
rect 1070 1147 1076 1148
rect 1072 1127 1074 1147
rect 1124 1128 1126 1194
rect 1132 1164 1134 1194
rect 1224 1191 1226 1201
rect 1274 1199 1280 1200
rect 1274 1195 1275 1199
rect 1279 1195 1280 1199
rect 1274 1194 1280 1195
rect 1222 1190 1228 1191
rect 1222 1186 1223 1190
rect 1227 1186 1228 1190
rect 1222 1185 1228 1186
rect 1276 1164 1278 1194
rect 1368 1191 1370 1201
rect 1418 1199 1424 1200
rect 1418 1195 1419 1199
rect 1423 1195 1424 1199
rect 1418 1194 1424 1195
rect 1366 1190 1372 1191
rect 1366 1186 1367 1190
rect 1371 1186 1372 1190
rect 1366 1185 1372 1186
rect 1420 1164 1422 1194
rect 1504 1191 1506 1201
rect 1554 1199 1560 1200
rect 1554 1195 1555 1199
rect 1559 1195 1560 1199
rect 1554 1194 1560 1195
rect 1502 1190 1508 1191
rect 1502 1186 1503 1190
rect 1507 1186 1508 1190
rect 1502 1185 1508 1186
rect 1556 1164 1558 1194
rect 1640 1191 1642 1201
rect 1752 1191 1754 1201
rect 1804 1200 1806 1238
rect 1830 1236 1831 1240
rect 1835 1236 1836 1240
rect 1830 1235 1836 1236
rect 1832 1207 1834 1235
rect 1872 1230 1874 1249
rect 1896 1233 1898 1249
rect 2072 1233 2074 1249
rect 1894 1232 1900 1233
rect 1870 1229 1876 1230
rect 1870 1225 1871 1229
rect 1875 1225 1876 1229
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 1894 1227 1900 1228
rect 2070 1232 2076 1233
rect 2070 1228 2071 1232
rect 2075 1228 2076 1232
rect 2070 1227 2076 1228
rect 1870 1224 1876 1225
rect 2138 1223 2144 1224
rect 2138 1219 2139 1223
rect 2143 1219 2144 1223
rect 2138 1218 2144 1219
rect 1954 1215 1960 1216
rect 1870 1212 1876 1213
rect 1870 1208 1871 1212
rect 1875 1208 1876 1212
rect 1954 1211 1955 1215
rect 1959 1211 1960 1215
rect 1954 1210 1960 1211
rect 1870 1207 1876 1208
rect 1831 1206 1835 1207
rect 1831 1201 1835 1202
rect 1802 1199 1808 1200
rect 1802 1195 1803 1199
rect 1807 1195 1808 1199
rect 1802 1194 1808 1195
rect 1638 1190 1644 1191
rect 1638 1186 1639 1190
rect 1643 1186 1644 1190
rect 1638 1185 1644 1186
rect 1750 1190 1756 1191
rect 1750 1186 1751 1190
rect 1755 1186 1756 1190
rect 1750 1185 1756 1186
rect 1802 1183 1808 1184
rect 1802 1179 1803 1183
rect 1807 1179 1808 1183
rect 1802 1178 1808 1179
rect 1804 1164 1806 1178
rect 1832 1173 1834 1201
rect 1872 1175 1874 1207
rect 1902 1194 1908 1195
rect 1902 1190 1903 1194
rect 1907 1190 1908 1194
rect 1902 1189 1908 1190
rect 1904 1175 1906 1189
rect 1871 1174 1875 1175
rect 1830 1172 1836 1173
rect 1830 1168 1831 1172
rect 1835 1168 1836 1172
rect 1871 1169 1875 1170
rect 1903 1174 1907 1175
rect 1903 1169 1907 1170
rect 1830 1167 1836 1168
rect 1130 1163 1136 1164
rect 1130 1159 1131 1163
rect 1135 1159 1136 1163
rect 1130 1158 1136 1159
rect 1274 1163 1280 1164
rect 1274 1159 1275 1163
rect 1279 1159 1280 1163
rect 1274 1158 1280 1159
rect 1418 1163 1424 1164
rect 1418 1159 1419 1163
rect 1423 1159 1424 1163
rect 1418 1158 1424 1159
rect 1554 1163 1560 1164
rect 1554 1159 1555 1163
rect 1559 1159 1560 1163
rect 1554 1158 1560 1159
rect 1802 1163 1808 1164
rect 1802 1159 1803 1163
rect 1807 1159 1808 1163
rect 1802 1158 1808 1159
rect 1830 1155 1836 1156
rect 1214 1152 1220 1153
rect 1214 1148 1215 1152
rect 1219 1148 1220 1152
rect 1214 1147 1220 1148
rect 1358 1152 1364 1153
rect 1358 1148 1359 1152
rect 1363 1148 1364 1152
rect 1358 1147 1364 1148
rect 1494 1152 1500 1153
rect 1494 1148 1495 1152
rect 1499 1148 1500 1152
rect 1494 1147 1500 1148
rect 1630 1152 1636 1153
rect 1630 1148 1631 1152
rect 1635 1148 1636 1152
rect 1630 1147 1636 1148
rect 1742 1152 1748 1153
rect 1742 1148 1743 1152
rect 1747 1148 1748 1152
rect 1830 1151 1831 1155
rect 1835 1151 1836 1155
rect 1830 1150 1836 1151
rect 1742 1147 1748 1148
rect 1122 1127 1128 1128
rect 1216 1127 1218 1147
rect 1360 1127 1362 1147
rect 1438 1127 1444 1128
rect 1496 1127 1498 1147
rect 1632 1127 1634 1147
rect 1744 1127 1746 1147
rect 1832 1127 1834 1150
rect 1872 1141 1874 1169
rect 1904 1159 1906 1169
rect 1956 1168 1958 1210
rect 2078 1194 2084 1195
rect 2078 1190 2079 1194
rect 2083 1190 2084 1194
rect 2078 1189 2084 1190
rect 2080 1175 2082 1189
rect 2140 1184 2142 1218
rect 2236 1184 2238 1290
rect 3590 1287 3596 1288
rect 2310 1284 2316 1285
rect 2310 1280 2311 1284
rect 2315 1280 2316 1284
rect 2310 1279 2316 1280
rect 2446 1284 2452 1285
rect 2446 1280 2447 1284
rect 2451 1280 2452 1284
rect 2446 1279 2452 1280
rect 2582 1284 2588 1285
rect 2582 1280 2583 1284
rect 2587 1280 2588 1284
rect 2582 1279 2588 1280
rect 2710 1284 2716 1285
rect 2710 1280 2711 1284
rect 2715 1280 2716 1284
rect 2710 1279 2716 1280
rect 2830 1284 2836 1285
rect 2830 1280 2831 1284
rect 2835 1280 2836 1284
rect 2830 1279 2836 1280
rect 2942 1284 2948 1285
rect 2942 1280 2943 1284
rect 2947 1280 2948 1284
rect 2942 1279 2948 1280
rect 3054 1284 3060 1285
rect 3054 1280 3055 1284
rect 3059 1280 3060 1284
rect 3054 1279 3060 1280
rect 3174 1284 3180 1285
rect 3174 1280 3175 1284
rect 3179 1280 3180 1284
rect 3590 1283 3591 1287
rect 3595 1283 3596 1287
rect 3590 1282 3596 1283
rect 3174 1279 3180 1280
rect 2312 1255 2314 1279
rect 2448 1255 2450 1279
rect 2584 1255 2586 1279
rect 2712 1255 2714 1279
rect 2832 1255 2834 1279
rect 2944 1255 2946 1279
rect 3056 1255 3058 1279
rect 3062 1267 3068 1268
rect 3062 1263 3063 1267
rect 3067 1263 3068 1267
rect 3062 1262 3068 1263
rect 2271 1254 2275 1255
rect 2271 1249 2275 1250
rect 2311 1254 2315 1255
rect 2311 1249 2315 1250
rect 2447 1254 2451 1255
rect 2447 1249 2451 1250
rect 2471 1254 2475 1255
rect 2471 1249 2475 1250
rect 2583 1254 2587 1255
rect 2583 1249 2587 1250
rect 2663 1254 2667 1255
rect 2663 1249 2667 1250
rect 2711 1254 2715 1255
rect 2711 1249 2715 1250
rect 2831 1254 2835 1255
rect 2831 1249 2835 1250
rect 2847 1254 2851 1255
rect 2847 1249 2851 1250
rect 2943 1254 2947 1255
rect 2943 1249 2947 1250
rect 3023 1254 3027 1255
rect 3023 1249 3027 1250
rect 3055 1254 3059 1255
rect 3055 1249 3059 1250
rect 2272 1233 2274 1249
rect 2472 1233 2474 1249
rect 2664 1233 2666 1249
rect 2848 1233 2850 1249
rect 3024 1233 3026 1249
rect 2270 1232 2276 1233
rect 2270 1228 2271 1232
rect 2275 1228 2276 1232
rect 2270 1227 2276 1228
rect 2470 1232 2476 1233
rect 2470 1228 2471 1232
rect 2475 1228 2476 1232
rect 2470 1227 2476 1228
rect 2662 1232 2668 1233
rect 2662 1228 2663 1232
rect 2667 1228 2668 1232
rect 2662 1227 2668 1228
rect 2846 1232 2852 1233
rect 2846 1228 2847 1232
rect 2851 1228 2852 1232
rect 2846 1227 2852 1228
rect 3022 1232 3028 1233
rect 3022 1228 3023 1232
rect 3027 1228 3028 1232
rect 3022 1227 3028 1228
rect 2590 1223 2596 1224
rect 2590 1219 2591 1223
rect 2595 1219 2596 1223
rect 2590 1218 2596 1219
rect 2778 1223 2784 1224
rect 2778 1219 2779 1223
rect 2783 1219 2784 1223
rect 2778 1218 2784 1219
rect 2914 1223 2920 1224
rect 2914 1219 2915 1223
rect 2919 1219 2920 1223
rect 2914 1218 2920 1219
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2478 1194 2484 1195
rect 2478 1190 2479 1194
rect 2483 1190 2484 1194
rect 2478 1189 2484 1190
rect 2138 1183 2144 1184
rect 2138 1179 2139 1183
rect 2143 1179 2144 1183
rect 2138 1178 2144 1179
rect 2234 1183 2240 1184
rect 2234 1179 2235 1183
rect 2239 1179 2240 1183
rect 2234 1178 2240 1179
rect 2280 1175 2282 1189
rect 2480 1175 2482 1189
rect 2507 1188 2511 1189
rect 2592 1184 2594 1218
rect 2722 1215 2728 1216
rect 2722 1211 2723 1215
rect 2727 1211 2728 1215
rect 2722 1210 2728 1211
rect 2670 1194 2676 1195
rect 2670 1190 2671 1194
rect 2675 1190 2676 1194
rect 2670 1189 2676 1190
rect 2506 1183 2512 1184
rect 2506 1179 2507 1183
rect 2511 1179 2512 1183
rect 2506 1178 2512 1179
rect 2590 1183 2596 1184
rect 2590 1179 2591 1183
rect 2595 1179 2596 1183
rect 2590 1178 2596 1179
rect 2672 1175 2674 1189
rect 1983 1174 1987 1175
rect 1983 1169 1987 1170
rect 2079 1174 2083 1175
rect 2079 1169 2083 1170
rect 2087 1174 2091 1175
rect 2087 1169 2091 1170
rect 2215 1174 2219 1175
rect 2215 1169 2219 1170
rect 2279 1174 2283 1175
rect 2279 1169 2283 1170
rect 2367 1174 2371 1175
rect 2367 1169 2371 1170
rect 2479 1174 2483 1175
rect 2479 1169 2483 1170
rect 2527 1174 2531 1175
rect 2527 1169 2531 1170
rect 2671 1174 2675 1175
rect 2671 1169 2675 1170
rect 2687 1174 2691 1175
rect 2687 1169 2691 1170
rect 1954 1167 1960 1168
rect 1954 1163 1955 1167
rect 1959 1163 1960 1167
rect 1954 1162 1960 1163
rect 1962 1167 1968 1168
rect 1962 1163 1963 1167
rect 1967 1163 1968 1167
rect 1962 1162 1968 1163
rect 1902 1158 1908 1159
rect 1902 1154 1903 1158
rect 1907 1154 1908 1158
rect 1902 1153 1908 1154
rect 1870 1140 1876 1141
rect 1870 1136 1871 1140
rect 1875 1136 1876 1140
rect 1870 1135 1876 1136
rect 1964 1132 1966 1162
rect 1984 1159 1986 1169
rect 2034 1167 2040 1168
rect 2034 1163 2035 1167
rect 2039 1163 2040 1167
rect 2034 1162 2040 1163
rect 1982 1158 1988 1159
rect 1982 1154 1983 1158
rect 1987 1154 1988 1158
rect 1982 1153 1988 1154
rect 2036 1132 2038 1162
rect 2088 1159 2090 1169
rect 2138 1167 2144 1168
rect 2138 1163 2139 1167
rect 2143 1163 2144 1167
rect 2138 1162 2144 1163
rect 2086 1158 2092 1159
rect 2086 1154 2087 1158
rect 2091 1154 2092 1158
rect 2086 1153 2092 1154
rect 2140 1132 2142 1162
rect 2216 1159 2218 1169
rect 2266 1167 2272 1168
rect 2266 1163 2267 1167
rect 2271 1163 2272 1167
rect 2266 1162 2272 1163
rect 2214 1158 2220 1159
rect 2214 1154 2215 1158
rect 2219 1154 2220 1158
rect 2214 1153 2220 1154
rect 2268 1132 2270 1162
rect 2368 1159 2370 1169
rect 2418 1167 2424 1168
rect 2418 1163 2419 1167
rect 2423 1163 2424 1167
rect 2418 1162 2424 1163
rect 2366 1158 2372 1159
rect 2366 1154 2367 1158
rect 2371 1154 2372 1158
rect 2366 1153 2372 1154
rect 2420 1132 2422 1162
rect 2528 1159 2530 1169
rect 2688 1159 2690 1169
rect 2724 1168 2726 1210
rect 2780 1189 2782 1218
rect 2854 1194 2860 1195
rect 2854 1190 2855 1194
rect 2859 1190 2860 1194
rect 2854 1189 2860 1190
rect 2779 1188 2783 1189
rect 2779 1183 2783 1184
rect 2856 1175 2858 1189
rect 2916 1184 2918 1218
rect 3030 1194 3036 1195
rect 3030 1190 3031 1194
rect 3035 1190 3036 1194
rect 3030 1189 3036 1190
rect 2914 1183 2920 1184
rect 2914 1179 2915 1183
rect 2919 1179 2920 1183
rect 2914 1178 2920 1179
rect 3032 1175 3034 1189
rect 3055 1183 3061 1184
rect 3055 1179 3056 1183
rect 3060 1182 3061 1183
rect 3064 1182 3066 1262
rect 3176 1255 3178 1279
rect 3592 1255 3594 1282
rect 3175 1254 3179 1255
rect 3175 1249 3179 1250
rect 3191 1254 3195 1255
rect 3191 1249 3195 1250
rect 3359 1254 3363 1255
rect 3359 1249 3363 1250
rect 3503 1254 3507 1255
rect 3503 1249 3507 1250
rect 3591 1254 3595 1255
rect 3591 1249 3595 1250
rect 3192 1233 3194 1249
rect 3360 1233 3362 1249
rect 3504 1233 3506 1249
rect 3190 1232 3196 1233
rect 3190 1228 3191 1232
rect 3195 1228 3196 1232
rect 3190 1227 3196 1228
rect 3358 1232 3364 1233
rect 3358 1228 3359 1232
rect 3363 1228 3364 1232
rect 3358 1227 3364 1228
rect 3502 1232 3508 1233
rect 3502 1228 3503 1232
rect 3507 1228 3508 1232
rect 3592 1230 3594 1249
rect 3502 1227 3508 1228
rect 3590 1229 3596 1230
rect 3590 1225 3591 1229
rect 3595 1225 3596 1229
rect 3590 1224 3596 1225
rect 3262 1223 3268 1224
rect 3262 1219 3263 1223
rect 3267 1219 3268 1223
rect 3262 1218 3268 1219
rect 3450 1223 3456 1224
rect 3450 1219 3451 1223
rect 3455 1219 3456 1223
rect 3450 1218 3456 1219
rect 3198 1194 3204 1195
rect 3198 1190 3199 1194
rect 3203 1190 3204 1194
rect 3198 1189 3204 1190
rect 3060 1180 3066 1182
rect 3060 1179 3061 1180
rect 3055 1178 3061 1179
rect 3200 1175 3202 1189
rect 3264 1184 3266 1218
rect 3366 1194 3372 1195
rect 3366 1190 3367 1194
rect 3371 1190 3372 1194
rect 3366 1189 3372 1190
rect 3262 1183 3268 1184
rect 3262 1179 3263 1183
rect 3267 1179 3268 1183
rect 3262 1178 3268 1179
rect 3368 1175 3370 1189
rect 3452 1184 3454 1218
rect 3562 1215 3568 1216
rect 3562 1211 3563 1215
rect 3567 1211 3568 1215
rect 3562 1210 3568 1211
rect 3590 1212 3596 1213
rect 3510 1194 3516 1195
rect 3510 1190 3511 1194
rect 3515 1190 3516 1194
rect 3510 1189 3516 1190
rect 3450 1183 3456 1184
rect 3450 1179 3451 1183
rect 3455 1179 3456 1183
rect 3450 1178 3456 1179
rect 3406 1175 3412 1176
rect 3512 1175 3514 1189
rect 2839 1174 2843 1175
rect 2839 1169 2843 1170
rect 2855 1174 2859 1175
rect 2855 1169 2859 1170
rect 2983 1174 2987 1175
rect 2983 1169 2987 1170
rect 3031 1174 3035 1175
rect 3031 1169 3035 1170
rect 3127 1174 3131 1175
rect 3127 1169 3131 1170
rect 3199 1174 3203 1175
rect 3199 1169 3203 1170
rect 3263 1174 3267 1175
rect 3263 1169 3267 1170
rect 3367 1174 3371 1175
rect 3367 1169 3371 1170
rect 3399 1174 3403 1175
rect 3406 1171 3407 1175
rect 3411 1171 3412 1175
rect 3406 1170 3412 1171
rect 3511 1174 3515 1175
rect 3399 1169 3403 1170
rect 2722 1167 2728 1168
rect 2722 1163 2723 1167
rect 2727 1163 2728 1167
rect 2722 1162 2728 1163
rect 2738 1167 2744 1168
rect 2738 1163 2739 1167
rect 2743 1163 2744 1167
rect 2738 1162 2744 1163
rect 2526 1158 2532 1159
rect 2526 1154 2527 1158
rect 2531 1154 2532 1158
rect 2526 1153 2532 1154
rect 2686 1158 2692 1159
rect 2686 1154 2687 1158
rect 2691 1154 2692 1158
rect 2686 1153 2692 1154
rect 2740 1132 2742 1162
rect 2840 1159 2842 1169
rect 2984 1159 2986 1169
rect 3010 1167 3016 1168
rect 3010 1163 3011 1167
rect 3015 1163 3016 1167
rect 3010 1162 3016 1163
rect 2838 1158 2844 1159
rect 2838 1154 2839 1158
rect 2843 1154 2844 1158
rect 2838 1153 2844 1154
rect 2982 1158 2988 1159
rect 2982 1154 2983 1158
rect 2987 1154 2988 1158
rect 2982 1153 2988 1154
rect 1962 1131 1968 1132
rect 1962 1127 1963 1131
rect 1967 1127 1968 1131
rect 975 1126 979 1127
rect 975 1121 979 1122
rect 1071 1126 1075 1127
rect 1071 1121 1075 1122
rect 1103 1126 1107 1127
rect 1122 1123 1123 1127
rect 1127 1123 1128 1127
rect 1122 1122 1128 1123
rect 1215 1126 1219 1127
rect 1103 1121 1107 1122
rect 1215 1121 1219 1122
rect 1223 1126 1227 1127
rect 1223 1121 1227 1122
rect 1343 1126 1347 1127
rect 1343 1121 1347 1122
rect 1359 1126 1363 1127
rect 1438 1123 1439 1127
rect 1443 1123 1444 1127
rect 1438 1122 1444 1123
rect 1471 1126 1475 1127
rect 1359 1121 1363 1122
rect 976 1105 978 1121
rect 1104 1105 1106 1121
rect 1224 1105 1226 1121
rect 1344 1105 1346 1121
rect 974 1104 980 1105
rect 974 1100 975 1104
rect 979 1100 980 1104
rect 974 1099 980 1100
rect 1102 1104 1108 1105
rect 1102 1100 1103 1104
rect 1107 1100 1108 1104
rect 1102 1099 1108 1100
rect 1222 1104 1228 1105
rect 1222 1100 1223 1104
rect 1227 1100 1228 1104
rect 1222 1099 1228 1100
rect 1342 1104 1348 1105
rect 1342 1100 1343 1104
rect 1347 1100 1348 1104
rect 1342 1099 1348 1100
rect 1440 1096 1442 1122
rect 1471 1121 1475 1122
rect 1495 1126 1499 1127
rect 1495 1121 1499 1122
rect 1631 1126 1635 1127
rect 1631 1121 1635 1122
rect 1743 1126 1747 1127
rect 1743 1121 1747 1122
rect 1831 1126 1835 1127
rect 1962 1126 1968 1127
rect 2034 1131 2040 1132
rect 2034 1127 2035 1131
rect 2039 1127 2040 1131
rect 2034 1126 2040 1127
rect 2138 1131 2144 1132
rect 2138 1127 2139 1131
rect 2143 1127 2144 1131
rect 2138 1126 2144 1127
rect 2266 1131 2272 1132
rect 2266 1127 2267 1131
rect 2271 1127 2272 1131
rect 2266 1126 2272 1127
rect 2418 1131 2424 1132
rect 2418 1127 2419 1131
rect 2423 1127 2424 1131
rect 2418 1126 2424 1127
rect 2738 1131 2744 1132
rect 2738 1127 2739 1131
rect 2743 1127 2744 1131
rect 2738 1126 2744 1127
rect 2918 1131 2924 1132
rect 2918 1127 2919 1131
rect 2923 1127 2924 1131
rect 2918 1126 2924 1127
rect 1831 1121 1835 1122
rect 1870 1123 1876 1124
rect 1472 1105 1474 1121
rect 1470 1104 1476 1105
rect 1470 1100 1471 1104
rect 1475 1100 1476 1104
rect 1832 1102 1834 1121
rect 1870 1119 1871 1123
rect 1875 1119 1876 1123
rect 1870 1118 1876 1119
rect 1894 1120 1900 1121
rect 1470 1099 1476 1100
rect 1830 1101 1836 1102
rect 1830 1097 1831 1101
rect 1835 1097 1836 1101
rect 1830 1096 1836 1097
rect 634 1095 640 1096
rect 634 1091 635 1095
rect 639 1091 640 1095
rect 634 1090 640 1091
rect 802 1095 808 1096
rect 802 1091 803 1095
rect 807 1091 808 1095
rect 802 1090 808 1091
rect 942 1095 948 1096
rect 942 1091 943 1095
rect 947 1091 948 1095
rect 942 1090 948 1091
rect 1062 1095 1068 1096
rect 1062 1091 1063 1095
rect 1067 1091 1068 1095
rect 1062 1090 1068 1091
rect 1186 1095 1192 1096
rect 1186 1091 1187 1095
rect 1191 1091 1192 1095
rect 1186 1090 1192 1091
rect 1306 1095 1312 1096
rect 1306 1091 1307 1095
rect 1311 1091 1312 1095
rect 1306 1090 1312 1091
rect 1430 1095 1436 1096
rect 1430 1091 1431 1095
rect 1435 1091 1436 1095
rect 1430 1090 1436 1091
rect 1438 1095 1444 1096
rect 1438 1091 1439 1095
rect 1443 1091 1444 1095
rect 1872 1091 1874 1118
rect 1894 1116 1895 1120
rect 1899 1116 1900 1120
rect 1894 1115 1900 1116
rect 1974 1120 1980 1121
rect 1974 1116 1975 1120
rect 1979 1116 1980 1120
rect 1974 1115 1980 1116
rect 2078 1120 2084 1121
rect 2078 1116 2079 1120
rect 2083 1116 2084 1120
rect 2078 1115 2084 1116
rect 2206 1120 2212 1121
rect 2206 1116 2207 1120
rect 2211 1116 2212 1120
rect 2206 1115 2212 1116
rect 2358 1120 2364 1121
rect 2358 1116 2359 1120
rect 2363 1116 2364 1120
rect 2358 1115 2364 1116
rect 2518 1120 2524 1121
rect 2518 1116 2519 1120
rect 2523 1116 2524 1120
rect 2518 1115 2524 1116
rect 2678 1120 2684 1121
rect 2678 1116 2679 1120
rect 2683 1116 2684 1120
rect 2678 1115 2684 1116
rect 2830 1120 2836 1121
rect 2830 1116 2831 1120
rect 2835 1116 2836 1120
rect 2830 1115 2836 1116
rect 1896 1091 1898 1115
rect 1976 1091 1978 1115
rect 2080 1091 2082 1115
rect 2208 1091 2210 1115
rect 2214 1103 2220 1104
rect 2214 1099 2215 1103
rect 2219 1099 2220 1103
rect 2214 1098 2220 1099
rect 1438 1090 1444 1091
rect 1871 1090 1875 1091
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 458 1055 464 1056
rect 458 1051 459 1055
rect 463 1051 464 1055
rect 458 1050 464 1051
rect 576 1043 578 1061
rect 636 1056 638 1090
rect 718 1066 724 1067
rect 718 1062 719 1066
rect 723 1062 724 1066
rect 718 1061 724 1062
rect 598 1055 604 1056
rect 598 1051 599 1055
rect 603 1051 604 1055
rect 598 1050 604 1051
rect 634 1055 640 1056
rect 634 1051 635 1055
rect 639 1051 640 1055
rect 634 1050 640 1051
rect 263 1042 267 1043
rect 263 1037 267 1038
rect 287 1042 291 1043
rect 287 1037 291 1038
rect 407 1042 411 1043
rect 414 1039 415 1043
rect 419 1039 420 1043
rect 414 1038 420 1039
rect 431 1042 435 1043
rect 407 1037 411 1038
rect 202 1035 208 1036
rect 202 1031 203 1035
rect 207 1031 208 1035
rect 202 1030 208 1031
rect 264 1027 266 1037
rect 314 1035 320 1036
rect 314 1031 315 1035
rect 319 1031 320 1035
rect 314 1030 320 1031
rect 142 1026 148 1027
rect 142 1022 143 1026
rect 147 1022 148 1026
rect 142 1021 148 1022
rect 262 1026 268 1027
rect 262 1022 263 1026
rect 267 1022 268 1026
rect 262 1021 268 1022
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 316 1000 318 1030
rect 408 1027 410 1037
rect 406 1026 412 1027
rect 406 1022 407 1026
rect 411 1022 412 1026
rect 406 1021 412 1022
rect 416 1000 418 1038
rect 431 1037 435 1038
rect 551 1042 555 1043
rect 551 1037 555 1038
rect 575 1042 579 1043
rect 575 1037 579 1038
rect 552 1027 554 1037
rect 550 1026 556 1027
rect 550 1022 551 1026
rect 555 1022 556 1026
rect 550 1021 556 1022
rect 600 1000 602 1050
rect 720 1043 722 1061
rect 804 1056 806 1090
rect 854 1066 860 1067
rect 854 1062 855 1066
rect 859 1062 860 1066
rect 854 1061 860 1062
rect 982 1066 988 1067
rect 982 1062 983 1066
rect 987 1062 988 1066
rect 982 1061 988 1062
rect 802 1055 808 1056
rect 802 1051 803 1055
rect 807 1051 808 1055
rect 802 1050 808 1051
rect 856 1043 858 1061
rect 984 1043 986 1061
rect 1064 1056 1066 1090
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1054 1055 1060 1056
rect 1054 1050 1055 1055
rect 1059 1050 1060 1055
rect 1062 1055 1068 1056
rect 1062 1051 1063 1055
rect 1067 1051 1068 1055
rect 1062 1050 1068 1051
rect 1055 1047 1059 1048
rect 1112 1043 1114 1061
rect 1188 1056 1190 1090
rect 1230 1066 1236 1067
rect 1230 1062 1231 1066
rect 1235 1062 1236 1066
rect 1230 1061 1236 1062
rect 1186 1055 1192 1056
rect 1186 1051 1187 1055
rect 1191 1051 1192 1055
rect 1186 1050 1192 1051
rect 1232 1043 1234 1061
rect 1308 1056 1310 1090
rect 1350 1066 1356 1067
rect 1350 1062 1351 1066
rect 1355 1062 1356 1066
rect 1350 1061 1356 1062
rect 1306 1055 1312 1056
rect 1306 1051 1307 1055
rect 1311 1051 1312 1055
rect 1306 1050 1312 1051
rect 1352 1043 1354 1061
rect 1432 1056 1434 1090
rect 1871 1085 1875 1086
rect 1895 1090 1899 1091
rect 1895 1085 1899 1086
rect 1975 1090 1979 1091
rect 1975 1085 1979 1086
rect 2079 1090 2083 1091
rect 2079 1085 2083 1086
rect 2167 1090 2171 1091
rect 2167 1085 2171 1086
rect 2207 1090 2211 1091
rect 2207 1085 2211 1086
rect 1830 1084 1836 1085
rect 1830 1080 1831 1084
rect 1835 1080 1836 1084
rect 1830 1079 1836 1080
rect 1478 1066 1484 1067
rect 1478 1062 1479 1066
rect 1483 1062 1484 1066
rect 1478 1061 1484 1062
rect 1430 1055 1436 1056
rect 1367 1052 1371 1053
rect 1430 1051 1431 1055
rect 1435 1051 1436 1055
rect 1430 1050 1436 1051
rect 1367 1047 1371 1048
rect 687 1042 691 1043
rect 687 1037 691 1038
rect 719 1042 723 1043
rect 719 1037 723 1038
rect 807 1042 811 1043
rect 807 1037 811 1038
rect 855 1042 859 1043
rect 855 1037 859 1038
rect 927 1042 931 1043
rect 927 1037 931 1038
rect 983 1042 987 1043
rect 983 1037 987 1038
rect 1039 1042 1043 1043
rect 1039 1037 1043 1038
rect 1111 1042 1115 1043
rect 1111 1037 1115 1038
rect 1143 1042 1147 1043
rect 1143 1037 1147 1038
rect 1231 1042 1235 1043
rect 1231 1037 1235 1038
rect 1247 1042 1251 1043
rect 1247 1037 1251 1038
rect 1351 1042 1355 1043
rect 1351 1037 1355 1038
rect 1359 1042 1363 1043
rect 1359 1037 1363 1038
rect 688 1027 690 1037
rect 694 1035 700 1036
rect 694 1031 695 1035
rect 699 1031 700 1035
rect 694 1030 700 1031
rect 754 1035 760 1036
rect 754 1031 755 1035
rect 759 1031 760 1035
rect 754 1030 760 1031
rect 686 1026 692 1027
rect 686 1022 687 1026
rect 691 1022 692 1026
rect 686 1021 692 1022
rect 696 1000 698 1030
rect 166 999 172 1000
rect 166 995 167 999
rect 171 995 172 999
rect 166 994 172 995
rect 314 999 320 1000
rect 314 995 315 999
rect 319 995 320 999
rect 314 994 320 995
rect 414 999 420 1000
rect 414 995 415 999
rect 419 995 420 999
rect 414 994 420 995
rect 598 999 604 1000
rect 598 995 599 999
rect 603 995 604 999
rect 598 994 604 995
rect 694 999 700 1000
rect 694 995 695 999
rect 699 995 700 999
rect 694 994 700 995
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 110 986 116 987
rect 134 988 140 989
rect 112 959 114 986
rect 134 984 135 988
rect 139 984 140 988
rect 134 983 140 984
rect 136 959 138 983
rect 111 958 115 959
rect 111 953 115 954
rect 135 958 139 959
rect 135 953 139 954
rect 112 934 114 953
rect 136 937 138 953
rect 134 936 140 937
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 134 932 135 936
rect 139 932 140 936
rect 134 931 140 932
rect 110 928 116 929
rect 110 916 116 917
rect 110 912 111 916
rect 115 912 116 916
rect 110 911 116 912
rect 112 875 114 911
rect 142 898 148 899
rect 142 894 143 898
rect 147 894 148 898
rect 142 893 148 894
rect 144 875 146 893
rect 168 888 170 994
rect 254 988 260 989
rect 254 984 255 988
rect 259 984 260 988
rect 254 983 260 984
rect 398 988 404 989
rect 398 984 399 988
rect 403 984 404 988
rect 398 983 404 984
rect 542 988 548 989
rect 542 984 543 988
rect 547 984 548 988
rect 542 983 548 984
rect 678 988 684 989
rect 678 984 679 988
rect 683 984 684 988
rect 678 983 684 984
rect 256 959 258 983
rect 400 959 402 983
rect 544 959 546 983
rect 680 959 682 983
rect 215 958 219 959
rect 215 953 219 954
rect 255 958 259 959
rect 255 953 259 954
rect 327 958 331 959
rect 327 953 331 954
rect 399 958 403 959
rect 399 953 403 954
rect 447 958 451 959
rect 447 953 451 954
rect 543 958 547 959
rect 543 953 547 954
rect 567 958 571 959
rect 567 953 571 954
rect 679 958 683 959
rect 679 953 683 954
rect 687 958 691 959
rect 687 953 691 954
rect 216 937 218 953
rect 328 937 330 953
rect 448 937 450 953
rect 568 937 570 953
rect 688 937 690 953
rect 214 936 220 937
rect 214 932 215 936
rect 219 932 220 936
rect 214 931 220 932
rect 326 936 332 937
rect 326 932 327 936
rect 331 932 332 936
rect 326 931 332 932
rect 446 936 452 937
rect 446 932 447 936
rect 451 932 452 936
rect 446 931 452 932
rect 566 936 572 937
rect 566 932 567 936
rect 571 932 572 936
rect 566 931 572 932
rect 686 936 692 937
rect 686 932 687 936
rect 691 932 692 936
rect 686 931 692 932
rect 756 928 758 1030
rect 808 1027 810 1037
rect 918 1035 924 1036
rect 918 1031 919 1035
rect 923 1031 924 1035
rect 918 1030 924 1031
rect 806 1026 812 1027
rect 806 1022 807 1026
rect 811 1022 812 1026
rect 806 1021 812 1022
rect 920 1000 922 1030
rect 928 1027 930 1037
rect 1030 1035 1036 1036
rect 1030 1031 1031 1035
rect 1035 1031 1036 1035
rect 1030 1030 1036 1031
rect 926 1026 932 1027
rect 926 1022 927 1026
rect 931 1022 932 1026
rect 926 1021 932 1022
rect 1032 1000 1034 1030
rect 1040 1027 1042 1037
rect 1090 1035 1096 1036
rect 1090 1031 1091 1035
rect 1095 1031 1096 1035
rect 1090 1030 1096 1031
rect 1038 1026 1044 1027
rect 1038 1022 1039 1026
rect 1043 1022 1044 1026
rect 1038 1021 1044 1022
rect 1092 1000 1094 1030
rect 1144 1027 1146 1037
rect 1194 1035 1200 1036
rect 1194 1031 1195 1035
rect 1199 1031 1200 1035
rect 1194 1030 1200 1031
rect 1142 1026 1148 1027
rect 1142 1022 1143 1026
rect 1147 1022 1148 1026
rect 1142 1021 1148 1022
rect 1196 1000 1198 1030
rect 1248 1027 1250 1037
rect 1298 1035 1304 1036
rect 1298 1031 1299 1035
rect 1303 1031 1304 1035
rect 1298 1030 1304 1031
rect 1246 1026 1252 1027
rect 1246 1022 1247 1026
rect 1251 1022 1252 1026
rect 1246 1021 1252 1022
rect 1300 1000 1302 1030
rect 1360 1027 1362 1037
rect 1358 1026 1364 1027
rect 1358 1022 1359 1026
rect 1363 1022 1364 1026
rect 1358 1021 1364 1022
rect 1368 1000 1370 1047
rect 1480 1043 1482 1061
rect 1832 1043 1834 1079
rect 1872 1066 1874 1085
rect 2168 1069 2170 1085
rect 2166 1068 2172 1069
rect 1870 1065 1876 1066
rect 1870 1061 1871 1065
rect 1875 1061 1876 1065
rect 2166 1064 2167 1068
rect 2171 1064 2172 1068
rect 2166 1063 2172 1064
rect 1870 1060 1876 1061
rect 1870 1048 1876 1049
rect 1870 1044 1871 1048
rect 1875 1044 1876 1048
rect 1870 1043 1876 1044
rect 1479 1042 1483 1043
rect 1479 1037 1483 1038
rect 1831 1042 1835 1043
rect 1831 1037 1835 1038
rect 1832 1009 1834 1037
rect 1872 1015 1874 1043
rect 2174 1030 2180 1031
rect 2174 1026 2175 1030
rect 2179 1026 2180 1030
rect 2174 1025 2180 1026
rect 2176 1015 2178 1025
rect 2216 1020 2218 1098
rect 2360 1091 2362 1115
rect 2520 1091 2522 1115
rect 2680 1091 2682 1115
rect 2832 1091 2834 1115
rect 2255 1090 2259 1091
rect 2255 1085 2259 1086
rect 2359 1090 2363 1091
rect 2359 1085 2363 1086
rect 2479 1090 2483 1091
rect 2479 1085 2483 1086
rect 2519 1090 2523 1091
rect 2519 1085 2523 1086
rect 2607 1090 2611 1091
rect 2607 1085 2611 1086
rect 2679 1090 2683 1091
rect 2679 1085 2683 1086
rect 2751 1090 2755 1091
rect 2751 1085 2755 1086
rect 2831 1090 2835 1091
rect 2831 1085 2835 1086
rect 2895 1090 2899 1091
rect 2895 1085 2899 1086
rect 2256 1069 2258 1085
rect 2360 1069 2362 1085
rect 2480 1069 2482 1085
rect 2608 1069 2610 1085
rect 2752 1069 2754 1085
rect 2896 1069 2898 1085
rect 2254 1068 2260 1069
rect 2254 1064 2255 1068
rect 2259 1064 2260 1068
rect 2254 1063 2260 1064
rect 2358 1068 2364 1069
rect 2358 1064 2359 1068
rect 2363 1064 2364 1068
rect 2358 1063 2364 1064
rect 2478 1068 2484 1069
rect 2478 1064 2479 1068
rect 2483 1064 2484 1068
rect 2478 1063 2484 1064
rect 2606 1068 2612 1069
rect 2606 1064 2607 1068
rect 2611 1064 2612 1068
rect 2606 1063 2612 1064
rect 2750 1068 2756 1069
rect 2750 1064 2751 1068
rect 2755 1064 2756 1068
rect 2750 1063 2756 1064
rect 2894 1068 2900 1069
rect 2894 1064 2895 1068
rect 2899 1064 2900 1068
rect 2894 1063 2900 1064
rect 2234 1059 2240 1060
rect 2234 1055 2235 1059
rect 2239 1055 2240 1059
rect 2234 1054 2240 1055
rect 2330 1059 2336 1060
rect 2330 1055 2331 1059
rect 2335 1055 2336 1059
rect 2330 1054 2336 1055
rect 2434 1059 2440 1060
rect 2434 1055 2435 1059
rect 2439 1055 2440 1059
rect 2434 1054 2440 1055
rect 2554 1059 2560 1060
rect 2554 1055 2555 1059
rect 2559 1055 2560 1059
rect 2554 1054 2560 1055
rect 2562 1059 2568 1060
rect 2562 1055 2563 1059
rect 2567 1055 2568 1059
rect 2562 1054 2568 1055
rect 2818 1059 2824 1060
rect 2818 1055 2819 1059
rect 2823 1055 2824 1059
rect 2818 1054 2824 1055
rect 2236 1020 2238 1054
rect 2262 1030 2268 1031
rect 2262 1026 2263 1030
rect 2267 1026 2268 1030
rect 2262 1025 2268 1026
rect 2214 1019 2220 1020
rect 2214 1015 2215 1019
rect 2219 1015 2220 1019
rect 1871 1014 1875 1015
rect 1871 1009 1875 1010
rect 2175 1014 2179 1015
rect 2214 1014 2220 1015
rect 2234 1019 2240 1020
rect 2234 1015 2235 1019
rect 2239 1015 2240 1019
rect 2264 1015 2266 1025
rect 2332 1020 2334 1054
rect 2366 1030 2372 1031
rect 2347 1028 2351 1029
rect 2366 1026 2367 1030
rect 2371 1026 2372 1030
rect 2366 1025 2372 1026
rect 2347 1023 2351 1024
rect 2330 1019 2336 1020
rect 2330 1015 2331 1019
rect 2335 1015 2336 1019
rect 2234 1014 2240 1015
rect 2263 1014 2267 1015
rect 2175 1009 2179 1010
rect 2263 1009 2267 1010
rect 2303 1014 2307 1015
rect 2330 1014 2336 1015
rect 2303 1009 2307 1010
rect 1830 1008 1836 1009
rect 1830 1004 1831 1008
rect 1835 1004 1836 1008
rect 1830 1003 1836 1004
rect 918 999 924 1000
rect 918 995 919 999
rect 923 995 924 999
rect 918 994 924 995
rect 1030 999 1036 1000
rect 1030 995 1031 999
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1090 999 1096 1000
rect 1090 995 1091 999
rect 1095 995 1096 999
rect 1090 994 1096 995
rect 1194 999 1200 1000
rect 1194 995 1195 999
rect 1199 995 1200 999
rect 1194 994 1200 995
rect 1298 999 1304 1000
rect 1298 995 1299 999
rect 1303 995 1304 999
rect 1298 994 1304 995
rect 1366 999 1372 1000
rect 1366 995 1367 999
rect 1371 995 1372 999
rect 1366 994 1372 995
rect 1830 991 1836 992
rect 798 988 804 989
rect 798 984 799 988
rect 803 984 804 988
rect 798 983 804 984
rect 918 988 924 989
rect 918 984 919 988
rect 923 984 924 988
rect 918 983 924 984
rect 1030 988 1036 989
rect 1030 984 1031 988
rect 1035 984 1036 988
rect 1030 983 1036 984
rect 1134 988 1140 989
rect 1134 984 1135 988
rect 1139 984 1140 988
rect 1134 983 1140 984
rect 1238 988 1244 989
rect 1238 984 1239 988
rect 1243 984 1244 988
rect 1238 983 1244 984
rect 1350 988 1356 989
rect 1350 984 1351 988
rect 1355 984 1356 988
rect 1830 987 1831 991
rect 1835 987 1836 991
rect 1830 986 1836 987
rect 1350 983 1356 984
rect 800 959 802 983
rect 920 959 922 983
rect 1032 959 1034 983
rect 1136 959 1138 983
rect 1240 959 1242 983
rect 1352 959 1354 983
rect 1832 959 1834 986
rect 1872 981 1874 1009
rect 2304 999 2306 1009
rect 2348 1008 2350 1023
rect 2368 1015 2370 1025
rect 2436 1020 2438 1054
rect 2486 1030 2492 1031
rect 2486 1026 2487 1030
rect 2491 1026 2492 1030
rect 2486 1025 2492 1026
rect 2434 1019 2440 1020
rect 2434 1015 2435 1019
rect 2439 1015 2440 1019
rect 2488 1015 2490 1025
rect 2556 1020 2558 1054
rect 2564 1029 2566 1054
rect 2810 1051 2816 1052
rect 2810 1047 2811 1051
rect 2815 1047 2816 1051
rect 2810 1046 2816 1047
rect 2614 1030 2620 1031
rect 2563 1028 2567 1029
rect 2614 1026 2615 1030
rect 2619 1026 2620 1030
rect 2614 1025 2620 1026
rect 2758 1030 2764 1031
rect 2758 1026 2759 1030
rect 2763 1026 2764 1030
rect 2758 1025 2764 1026
rect 2563 1023 2567 1024
rect 2554 1019 2560 1020
rect 2554 1015 2555 1019
rect 2559 1015 2560 1019
rect 2616 1015 2618 1025
rect 2760 1015 2762 1025
rect 2367 1014 2371 1015
rect 2367 1009 2371 1010
rect 2383 1014 2387 1015
rect 2434 1014 2440 1015
rect 2471 1014 2475 1015
rect 2383 1009 2387 1010
rect 2471 1009 2475 1010
rect 2487 1014 2491 1015
rect 2554 1014 2560 1015
rect 2567 1014 2571 1015
rect 2487 1009 2491 1010
rect 2567 1009 2571 1010
rect 2615 1014 2619 1015
rect 2615 1009 2619 1010
rect 2671 1014 2675 1015
rect 2671 1009 2675 1010
rect 2759 1014 2763 1015
rect 2759 1009 2763 1010
rect 2783 1014 2787 1015
rect 2783 1009 2787 1010
rect 2346 1007 2352 1008
rect 2346 1003 2347 1007
rect 2351 1003 2352 1007
rect 2346 1002 2352 1003
rect 2354 1007 2360 1008
rect 2354 1003 2355 1007
rect 2359 1003 2360 1007
rect 2354 1002 2360 1003
rect 2302 998 2308 999
rect 2302 994 2303 998
rect 2307 994 2308 998
rect 2302 993 2308 994
rect 1870 980 1876 981
rect 1870 976 1871 980
rect 1875 976 1876 980
rect 1870 975 1876 976
rect 2356 972 2358 1002
rect 2384 999 2386 1009
rect 2434 1007 2440 1008
rect 2434 1003 2435 1007
rect 2439 1003 2440 1007
rect 2434 1002 2440 1003
rect 2382 998 2388 999
rect 2382 994 2383 998
rect 2387 994 2388 998
rect 2382 993 2388 994
rect 2436 972 2438 1002
rect 2472 999 2474 1009
rect 2522 1007 2528 1008
rect 2522 1003 2523 1007
rect 2527 1003 2528 1007
rect 2522 1002 2528 1003
rect 2470 998 2476 999
rect 2470 994 2471 998
rect 2475 994 2476 998
rect 2470 993 2476 994
rect 2524 972 2526 1002
rect 2568 999 2570 1009
rect 2672 999 2674 1009
rect 2784 999 2786 1009
rect 2812 1008 2814 1046
rect 2820 1020 2822 1054
rect 2902 1030 2908 1031
rect 2902 1026 2903 1030
rect 2907 1026 2908 1030
rect 2902 1025 2908 1026
rect 2818 1019 2824 1020
rect 2818 1015 2819 1019
rect 2823 1015 2824 1019
rect 2904 1015 2906 1025
rect 2920 1020 2922 1126
rect 2974 1120 2980 1121
rect 2974 1116 2975 1120
rect 2979 1116 2980 1120
rect 2974 1115 2980 1116
rect 2976 1091 2978 1115
rect 2975 1090 2979 1091
rect 2975 1085 2979 1086
rect 3012 1060 3014 1162
rect 3128 1159 3130 1169
rect 3178 1167 3184 1168
rect 3178 1163 3179 1167
rect 3183 1163 3184 1167
rect 3178 1162 3184 1163
rect 3126 1158 3132 1159
rect 3126 1154 3127 1158
rect 3131 1154 3132 1158
rect 3126 1153 3132 1154
rect 3180 1132 3182 1162
rect 3264 1159 3266 1169
rect 3314 1167 3320 1168
rect 3314 1163 3315 1167
rect 3319 1163 3320 1167
rect 3314 1162 3320 1163
rect 3262 1158 3268 1159
rect 3262 1154 3263 1158
rect 3267 1154 3268 1158
rect 3262 1153 3268 1154
rect 3316 1132 3318 1162
rect 3400 1159 3402 1169
rect 3398 1158 3404 1159
rect 3398 1154 3399 1158
rect 3403 1154 3404 1158
rect 3398 1153 3404 1154
rect 3408 1132 3410 1170
rect 3511 1169 3515 1170
rect 3512 1159 3514 1169
rect 3564 1168 3566 1210
rect 3590 1208 3591 1212
rect 3595 1208 3596 1212
rect 3590 1207 3596 1208
rect 3592 1175 3594 1207
rect 3591 1174 3595 1175
rect 3591 1169 3595 1170
rect 3562 1167 3568 1168
rect 3562 1163 3563 1167
rect 3567 1163 3568 1167
rect 3562 1162 3568 1163
rect 3510 1158 3516 1159
rect 3510 1154 3511 1158
rect 3515 1154 3516 1158
rect 3510 1153 3516 1154
rect 3592 1141 3594 1169
rect 3590 1140 3596 1141
rect 3590 1136 3591 1140
rect 3595 1136 3596 1140
rect 3590 1135 3596 1136
rect 3178 1131 3184 1132
rect 3178 1127 3179 1131
rect 3183 1127 3184 1131
rect 3178 1126 3184 1127
rect 3314 1131 3320 1132
rect 3314 1127 3315 1131
rect 3319 1127 3320 1131
rect 3314 1126 3320 1127
rect 3406 1131 3412 1132
rect 3406 1127 3407 1131
rect 3411 1127 3412 1131
rect 3406 1126 3412 1127
rect 3534 1131 3540 1132
rect 3534 1127 3535 1131
rect 3539 1127 3540 1131
rect 3534 1126 3540 1127
rect 3118 1120 3124 1121
rect 3118 1116 3119 1120
rect 3123 1116 3124 1120
rect 3118 1115 3124 1116
rect 3254 1120 3260 1121
rect 3254 1116 3255 1120
rect 3259 1116 3260 1120
rect 3254 1115 3260 1116
rect 3390 1120 3396 1121
rect 3390 1116 3391 1120
rect 3395 1116 3396 1120
rect 3390 1115 3396 1116
rect 3502 1120 3508 1121
rect 3502 1116 3503 1120
rect 3507 1116 3508 1120
rect 3502 1115 3508 1116
rect 3120 1091 3122 1115
rect 3256 1091 3258 1115
rect 3392 1091 3394 1115
rect 3504 1091 3506 1115
rect 3047 1090 3051 1091
rect 3047 1085 3051 1086
rect 3119 1090 3123 1091
rect 3119 1085 3123 1086
rect 3207 1090 3211 1091
rect 3207 1085 3211 1086
rect 3255 1090 3259 1091
rect 3255 1085 3259 1086
rect 3367 1090 3371 1091
rect 3367 1085 3371 1086
rect 3391 1090 3395 1091
rect 3391 1085 3395 1086
rect 3503 1090 3507 1091
rect 3503 1085 3507 1086
rect 3048 1069 3050 1085
rect 3208 1069 3210 1085
rect 3368 1069 3370 1085
rect 3504 1069 3506 1085
rect 3046 1068 3052 1069
rect 3046 1064 3047 1068
rect 3051 1064 3052 1068
rect 3046 1063 3052 1064
rect 3206 1068 3212 1069
rect 3206 1064 3207 1068
rect 3211 1064 3212 1068
rect 3206 1063 3212 1064
rect 3366 1068 3372 1069
rect 3366 1064 3367 1068
rect 3371 1064 3372 1068
rect 3366 1063 3372 1064
rect 3502 1068 3508 1069
rect 3502 1064 3503 1068
rect 3507 1064 3508 1068
rect 3502 1063 3508 1064
rect 3010 1059 3016 1060
rect 3010 1055 3011 1059
rect 3015 1055 3016 1059
rect 3010 1054 3016 1055
rect 3114 1059 3120 1060
rect 3114 1055 3115 1059
rect 3119 1055 3120 1059
rect 3114 1054 3120 1055
rect 3274 1059 3280 1060
rect 3274 1055 3275 1059
rect 3279 1055 3280 1059
rect 3274 1054 3280 1055
rect 3054 1030 3060 1031
rect 3054 1026 3055 1030
rect 3059 1026 3060 1030
rect 3054 1025 3060 1026
rect 2918 1019 2924 1020
rect 2918 1015 2919 1019
rect 2923 1015 2924 1019
rect 3056 1015 3058 1025
rect 3116 1020 3118 1054
rect 3214 1030 3220 1031
rect 3214 1026 3215 1030
rect 3219 1026 3220 1030
rect 3214 1025 3220 1026
rect 3114 1019 3120 1020
rect 3114 1015 3115 1019
rect 3119 1015 3120 1019
rect 3216 1015 3218 1025
rect 3276 1020 3278 1054
rect 3374 1030 3380 1031
rect 3374 1026 3375 1030
rect 3379 1026 3380 1030
rect 3374 1025 3380 1026
rect 3510 1030 3516 1031
rect 3510 1026 3511 1030
rect 3515 1026 3516 1030
rect 3510 1025 3516 1026
rect 3274 1019 3280 1020
rect 3274 1015 3275 1019
rect 3279 1015 3280 1019
rect 3376 1015 3378 1025
rect 3398 1019 3404 1020
rect 3398 1015 3399 1019
rect 3403 1015 3404 1019
rect 3512 1015 3514 1025
rect 3536 1020 3538 1126
rect 3590 1123 3596 1124
rect 3590 1119 3591 1123
rect 3595 1119 3596 1123
rect 3590 1118 3596 1119
rect 3592 1091 3594 1118
rect 3591 1090 3595 1091
rect 3591 1085 3595 1086
rect 3592 1066 3594 1085
rect 3590 1065 3596 1066
rect 3590 1061 3591 1065
rect 3595 1061 3596 1065
rect 3590 1060 3596 1061
rect 3562 1051 3568 1052
rect 3562 1047 3563 1051
rect 3567 1047 3568 1051
rect 3562 1046 3568 1047
rect 3590 1048 3596 1049
rect 3534 1019 3540 1020
rect 3534 1015 3535 1019
rect 3539 1015 3540 1019
rect 2818 1014 2824 1015
rect 2903 1014 2907 1015
rect 2903 1009 2907 1010
rect 2911 1014 2915 1015
rect 2918 1014 2924 1015
rect 3055 1014 3059 1015
rect 3114 1014 3120 1015
rect 3207 1014 3211 1015
rect 2911 1009 2915 1010
rect 3055 1009 3059 1010
rect 3207 1009 3211 1010
rect 3215 1014 3219 1015
rect 3274 1014 3280 1015
rect 3367 1014 3371 1015
rect 3215 1009 3219 1010
rect 3367 1009 3371 1010
rect 3375 1014 3379 1015
rect 3398 1014 3404 1015
rect 3511 1014 3515 1015
rect 3534 1014 3540 1015
rect 3375 1009 3379 1010
rect 2810 1007 2816 1008
rect 2810 1003 2811 1007
rect 2815 1003 2816 1007
rect 2810 1002 2816 1003
rect 2834 1007 2840 1008
rect 2834 1003 2835 1007
rect 2839 1003 2840 1007
rect 2834 1002 2840 1003
rect 2566 998 2572 999
rect 2566 994 2567 998
rect 2571 994 2572 998
rect 2566 993 2572 994
rect 2670 998 2676 999
rect 2670 994 2671 998
rect 2675 994 2676 998
rect 2670 993 2676 994
rect 2782 998 2788 999
rect 2782 994 2783 998
rect 2787 994 2788 998
rect 2782 993 2788 994
rect 2836 972 2838 1002
rect 2912 999 2914 1009
rect 3056 999 3058 1009
rect 3074 1007 3080 1008
rect 3074 1003 3075 1007
rect 3079 1003 3080 1007
rect 3074 1002 3080 1003
rect 3106 1007 3112 1008
rect 3106 1003 3107 1007
rect 3111 1003 3112 1007
rect 3106 1002 3112 1003
rect 2910 998 2916 999
rect 2910 994 2911 998
rect 2915 994 2916 998
rect 2910 993 2916 994
rect 3054 998 3060 999
rect 3054 994 3055 998
rect 3059 994 3060 998
rect 3054 993 3060 994
rect 2354 971 2360 972
rect 2354 967 2355 971
rect 2359 967 2360 971
rect 2354 966 2360 967
rect 2434 971 2440 972
rect 2434 967 2435 971
rect 2439 967 2440 971
rect 2434 966 2440 967
rect 2522 971 2528 972
rect 2522 967 2523 971
rect 2527 967 2528 971
rect 2522 966 2528 967
rect 2722 971 2728 972
rect 2722 967 2723 971
rect 2727 967 2728 971
rect 2722 966 2728 967
rect 2834 971 2840 972
rect 2834 967 2835 971
rect 2839 967 2840 971
rect 2834 966 2840 967
rect 1870 963 1876 964
rect 1870 959 1871 963
rect 1875 959 1876 963
rect 799 958 803 959
rect 799 953 803 954
rect 911 958 915 959
rect 911 953 915 954
rect 919 958 923 959
rect 919 953 923 954
rect 1015 958 1019 959
rect 1015 953 1019 954
rect 1031 958 1035 959
rect 1031 953 1035 954
rect 1119 958 1123 959
rect 1119 953 1123 954
rect 1135 958 1139 959
rect 1135 953 1139 954
rect 1223 958 1227 959
rect 1223 953 1227 954
rect 1239 958 1243 959
rect 1239 953 1243 954
rect 1327 958 1331 959
rect 1327 953 1331 954
rect 1351 958 1355 959
rect 1351 953 1355 954
rect 1831 958 1835 959
rect 1870 958 1876 959
rect 2294 960 2300 961
rect 1831 953 1835 954
rect 800 937 802 953
rect 912 937 914 953
rect 1016 937 1018 953
rect 1120 937 1122 953
rect 1224 937 1226 953
rect 1328 937 1330 953
rect 798 936 804 937
rect 798 932 799 936
rect 803 932 804 936
rect 798 931 804 932
rect 910 936 916 937
rect 910 932 911 936
rect 915 932 916 936
rect 910 931 916 932
rect 1014 936 1020 937
rect 1014 932 1015 936
rect 1019 932 1020 936
rect 1014 931 1020 932
rect 1118 936 1124 937
rect 1118 932 1119 936
rect 1123 932 1124 936
rect 1118 931 1124 932
rect 1222 936 1228 937
rect 1222 932 1223 936
rect 1227 932 1228 936
rect 1222 931 1228 932
rect 1326 936 1332 937
rect 1326 932 1327 936
rect 1331 932 1332 936
rect 1832 934 1834 953
rect 1326 931 1332 932
rect 1830 933 1836 934
rect 1830 929 1831 933
rect 1835 929 1836 933
rect 1872 931 1874 958
rect 2294 956 2295 960
rect 2299 956 2300 960
rect 2294 955 2300 956
rect 2374 960 2380 961
rect 2374 956 2375 960
rect 2379 956 2380 960
rect 2374 955 2380 956
rect 2462 960 2468 961
rect 2462 956 2463 960
rect 2467 956 2468 960
rect 2462 955 2468 956
rect 2558 960 2564 961
rect 2558 956 2559 960
rect 2563 956 2564 960
rect 2558 955 2564 956
rect 2662 960 2668 961
rect 2662 956 2663 960
rect 2667 956 2668 960
rect 2662 955 2668 956
rect 2296 931 2298 955
rect 2376 931 2378 955
rect 2464 931 2466 955
rect 2560 931 2562 955
rect 2664 931 2666 955
rect 1830 928 1836 929
rect 1871 930 1875 931
rect 202 927 208 928
rect 202 923 203 927
rect 207 923 208 927
rect 202 922 208 923
rect 282 927 288 928
rect 282 923 283 927
rect 287 923 288 927
rect 282 922 288 923
rect 398 927 404 928
rect 398 923 399 927
rect 403 923 404 927
rect 398 922 404 923
rect 426 927 432 928
rect 426 923 427 927
rect 431 923 432 927
rect 426 922 432 923
rect 650 927 656 928
rect 650 923 651 927
rect 655 923 656 927
rect 650 922 656 923
rect 754 927 760 928
rect 754 923 755 927
rect 759 923 760 927
rect 754 922 760 923
rect 866 927 872 928
rect 866 923 867 927
rect 871 923 872 927
rect 866 922 872 923
rect 978 927 984 928
rect 978 923 979 927
rect 983 923 984 927
rect 978 922 984 923
rect 1082 927 1088 928
rect 1082 923 1083 927
rect 1087 923 1088 927
rect 1082 922 1088 923
rect 1298 927 1304 928
rect 1298 923 1299 927
rect 1303 923 1304 927
rect 1871 925 1875 926
rect 2279 930 2283 931
rect 2279 925 2283 926
rect 2295 930 2299 931
rect 2295 925 2299 926
rect 2359 930 2363 931
rect 2359 925 2363 926
rect 2375 930 2379 931
rect 2375 925 2379 926
rect 2439 930 2443 931
rect 2439 925 2443 926
rect 2463 930 2467 931
rect 2463 925 2467 926
rect 2519 930 2523 931
rect 2519 925 2523 926
rect 2559 930 2563 931
rect 2559 925 2563 926
rect 2607 930 2611 931
rect 2607 925 2611 926
rect 2663 930 2667 931
rect 2663 925 2667 926
rect 2703 930 2707 931
rect 2703 925 2707 926
rect 1298 922 1304 923
rect 204 888 206 922
rect 222 898 228 899
rect 222 894 223 898
rect 227 894 228 898
rect 222 893 228 894
rect 166 887 172 888
rect 166 883 167 887
rect 171 883 172 887
rect 166 882 172 883
rect 202 887 208 888
rect 202 883 203 887
rect 207 883 208 887
rect 202 882 208 883
rect 224 875 226 893
rect 284 888 286 922
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 282 887 288 888
rect 282 883 283 887
rect 287 883 288 887
rect 282 882 288 883
rect 336 875 338 893
rect 400 888 402 922
rect 398 887 404 888
rect 398 883 399 887
rect 403 883 404 887
rect 398 882 404 883
rect 111 874 115 875
rect 111 869 115 870
rect 143 874 147 875
rect 143 869 147 870
rect 223 874 227 875
rect 223 869 227 870
rect 255 874 259 875
rect 255 869 259 870
rect 335 874 339 875
rect 335 869 339 870
rect 399 874 403 875
rect 399 869 403 870
rect 112 841 114 869
rect 144 859 146 869
rect 256 859 258 869
rect 262 867 268 868
rect 262 863 263 867
rect 267 863 268 867
rect 262 862 268 863
rect 142 858 148 859
rect 142 854 143 858
rect 147 854 148 858
rect 142 853 148 854
rect 254 858 260 859
rect 254 854 255 858
rect 259 854 260 858
rect 254 853 260 854
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 110 835 116 836
rect 264 832 266 862
rect 400 859 402 869
rect 428 868 430 922
rect 454 898 460 899
rect 454 894 455 898
rect 459 894 460 898
rect 454 893 460 894
rect 574 898 580 899
rect 574 894 575 898
rect 579 894 580 898
rect 574 893 580 894
rect 456 875 458 893
rect 576 875 578 893
rect 652 888 654 922
rect 694 898 700 899
rect 694 894 695 898
rect 699 894 700 898
rect 694 893 700 894
rect 806 898 812 899
rect 806 894 807 898
rect 811 894 812 898
rect 806 893 812 894
rect 598 887 604 888
rect 598 883 599 887
rect 603 883 604 887
rect 598 882 604 883
rect 650 887 656 888
rect 650 883 651 887
rect 655 883 656 887
rect 650 882 656 883
rect 455 874 459 875
rect 455 869 459 870
rect 559 874 563 875
rect 559 869 563 870
rect 575 874 579 875
rect 575 869 579 870
rect 406 867 412 868
rect 406 863 407 867
rect 411 863 412 867
rect 406 862 412 863
rect 426 867 432 868
rect 426 863 427 867
rect 431 863 432 867
rect 426 862 432 863
rect 398 858 404 859
rect 398 854 399 858
rect 403 854 404 858
rect 398 853 404 854
rect 408 832 410 862
rect 560 859 562 869
rect 558 858 564 859
rect 558 854 559 858
rect 563 854 564 858
rect 558 853 564 854
rect 600 832 602 882
rect 696 875 698 893
rect 808 875 810 893
rect 868 888 870 922
rect 918 898 924 899
rect 918 894 919 898
rect 923 894 924 898
rect 918 893 924 894
rect 866 887 872 888
rect 866 883 867 887
rect 871 883 872 887
rect 866 882 872 883
rect 920 875 922 893
rect 980 888 982 922
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 978 887 984 888
rect 978 883 979 887
rect 983 883 984 887
rect 978 882 984 883
rect 1024 875 1026 893
rect 1084 888 1086 922
rect 1194 919 1200 920
rect 1194 915 1195 919
rect 1199 915 1200 919
rect 1194 914 1200 915
rect 1126 898 1132 899
rect 1126 894 1127 898
rect 1131 894 1132 898
rect 1126 893 1132 894
rect 1082 887 1088 888
rect 1082 883 1083 887
rect 1087 883 1088 887
rect 1082 882 1088 883
rect 1128 875 1130 893
rect 1196 888 1198 914
rect 1230 898 1236 899
rect 1230 894 1231 898
rect 1235 894 1236 898
rect 1230 893 1236 894
rect 1194 887 1200 888
rect 1194 883 1195 887
rect 1199 883 1200 887
rect 1194 882 1200 883
rect 1202 887 1208 888
rect 1202 883 1203 887
rect 1207 883 1208 887
rect 1202 882 1208 883
rect 695 874 699 875
rect 695 869 699 870
rect 719 874 723 875
rect 719 869 723 870
rect 807 874 811 875
rect 807 869 811 870
rect 871 874 875 875
rect 871 869 875 870
rect 919 874 923 875
rect 919 869 923 870
rect 1015 874 1019 875
rect 1015 869 1019 870
rect 1023 874 1027 875
rect 1023 869 1027 870
rect 1127 874 1131 875
rect 1127 869 1131 870
rect 1151 874 1155 875
rect 1151 869 1155 870
rect 720 859 722 869
rect 726 867 732 868
rect 726 863 727 867
rect 731 863 732 867
rect 726 862 732 863
rect 718 858 724 859
rect 718 854 719 858
rect 723 854 724 858
rect 718 853 724 854
rect 728 832 730 862
rect 872 859 874 869
rect 878 867 884 868
rect 878 863 879 867
rect 883 863 884 867
rect 878 862 884 863
rect 886 867 892 868
rect 886 863 887 867
rect 891 863 892 867
rect 886 862 892 863
rect 870 858 876 859
rect 870 854 871 858
rect 875 854 876 858
rect 870 853 876 854
rect 880 832 882 862
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 262 831 268 832
rect 262 827 263 831
rect 267 827 268 831
rect 262 826 268 827
rect 406 831 412 832
rect 406 827 407 831
rect 411 827 412 831
rect 406 826 412 827
rect 598 831 604 832
rect 598 827 599 831
rect 603 827 604 831
rect 598 826 604 827
rect 726 831 732 832
rect 726 827 727 831
rect 731 827 732 831
rect 726 826 732 827
rect 878 831 884 832
rect 878 827 879 831
rect 883 827 884 831
rect 878 826 884 827
rect 110 823 116 824
rect 110 819 111 823
rect 115 819 116 823
rect 110 818 116 819
rect 134 820 140 821
rect 112 787 114 818
rect 134 816 135 820
rect 139 816 140 820
rect 134 815 140 816
rect 136 787 138 815
rect 111 786 115 787
rect 111 781 115 782
rect 135 786 139 787
rect 135 781 139 782
rect 112 762 114 781
rect 136 765 138 781
rect 134 764 140 765
rect 110 761 116 762
rect 110 757 111 761
rect 115 757 116 761
rect 134 760 135 764
rect 139 760 140 764
rect 134 759 140 760
rect 110 756 116 757
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 110 739 116 740
rect 112 699 114 739
rect 142 726 148 727
rect 142 722 143 726
rect 147 722 148 726
rect 142 721 148 722
rect 144 699 146 721
rect 168 716 170 826
rect 246 820 252 821
rect 246 816 247 820
rect 251 816 252 820
rect 246 815 252 816
rect 390 820 396 821
rect 390 816 391 820
rect 395 816 396 820
rect 390 815 396 816
rect 550 820 556 821
rect 550 816 551 820
rect 555 816 556 820
rect 550 815 556 816
rect 710 820 716 821
rect 710 816 711 820
rect 715 816 716 820
rect 710 815 716 816
rect 862 820 868 821
rect 862 816 863 820
rect 867 816 868 820
rect 862 815 868 816
rect 248 787 250 815
rect 392 787 394 815
rect 552 787 554 815
rect 712 787 714 815
rect 864 787 866 815
rect 247 786 251 787
rect 247 781 251 782
rect 263 786 267 787
rect 263 781 267 782
rect 391 786 395 787
rect 391 781 395 782
rect 431 786 435 787
rect 431 781 435 782
rect 551 786 555 787
rect 551 781 555 782
rect 607 786 611 787
rect 607 781 611 782
rect 711 786 715 787
rect 711 781 715 782
rect 783 786 787 787
rect 783 781 787 782
rect 863 786 867 787
rect 863 781 867 782
rect 264 765 266 781
rect 432 765 434 781
rect 608 765 610 781
rect 784 765 786 781
rect 262 764 268 765
rect 262 760 263 764
rect 267 760 268 764
rect 262 759 268 760
rect 430 764 436 765
rect 430 760 431 764
rect 435 760 436 764
rect 430 759 436 760
rect 606 764 612 765
rect 606 760 607 764
rect 611 760 612 764
rect 606 759 612 760
rect 782 764 788 765
rect 782 760 783 764
rect 787 760 788 764
rect 782 759 788 760
rect 218 755 224 756
rect 218 751 219 755
rect 223 751 224 755
rect 218 750 224 751
rect 330 755 336 756
rect 330 751 331 755
rect 335 751 336 755
rect 330 750 336 751
rect 850 755 856 756
rect 850 751 851 755
rect 855 751 856 755
rect 850 750 856 751
rect 220 716 222 750
rect 322 747 328 748
rect 322 743 323 747
rect 327 743 328 747
rect 322 742 328 743
rect 270 726 276 727
rect 270 722 271 726
rect 275 722 276 726
rect 270 721 276 722
rect 166 715 172 716
rect 166 711 167 715
rect 171 711 172 715
rect 166 710 172 711
rect 218 715 224 716
rect 218 711 219 715
rect 223 711 224 715
rect 218 710 224 711
rect 272 699 274 721
rect 111 698 115 699
rect 111 693 115 694
rect 143 698 147 699
rect 143 693 147 694
rect 271 698 275 699
rect 271 693 275 694
rect 295 698 299 699
rect 295 693 299 694
rect 112 665 114 693
rect 296 683 298 693
rect 324 692 326 742
rect 332 716 334 750
rect 438 726 444 727
rect 438 722 439 726
rect 443 722 444 726
rect 438 721 444 722
rect 614 726 620 727
rect 614 722 615 726
rect 619 722 620 726
rect 614 721 620 722
rect 790 726 796 727
rect 790 722 791 726
rect 795 722 796 726
rect 790 721 796 722
rect 330 715 336 716
rect 330 711 331 715
rect 335 711 336 715
rect 330 710 336 711
rect 440 699 442 721
rect 616 699 618 721
rect 792 699 794 721
rect 852 716 854 750
rect 888 748 890 862
rect 1016 859 1018 869
rect 1106 863 1112 864
rect 1106 859 1107 863
rect 1111 859 1112 863
rect 1152 859 1154 869
rect 1014 858 1020 859
rect 1106 858 1112 859
rect 1150 858 1156 859
rect 1014 854 1015 858
rect 1019 854 1020 858
rect 1014 853 1020 854
rect 1108 832 1110 858
rect 1150 854 1151 858
rect 1155 854 1156 858
rect 1150 853 1156 854
rect 1204 832 1206 882
rect 1232 875 1234 893
rect 1300 888 1302 922
rect 1830 916 1836 917
rect 1830 912 1831 916
rect 1835 912 1836 916
rect 1830 911 1836 912
rect 1334 898 1340 899
rect 1334 894 1335 898
rect 1339 894 1340 898
rect 1334 893 1340 894
rect 1298 887 1304 888
rect 1298 883 1299 887
rect 1303 883 1304 887
rect 1298 882 1304 883
rect 1286 875 1292 876
rect 1336 875 1338 893
rect 1832 875 1834 911
rect 1872 906 1874 925
rect 2280 909 2282 925
rect 2360 909 2362 925
rect 2440 909 2442 925
rect 2520 909 2522 925
rect 2608 909 2610 925
rect 2704 909 2706 925
rect 2278 908 2284 909
rect 1870 905 1876 906
rect 1870 901 1871 905
rect 1875 901 1876 905
rect 2278 904 2279 908
rect 2283 904 2284 908
rect 2278 903 2284 904
rect 2358 908 2364 909
rect 2358 904 2359 908
rect 2363 904 2364 908
rect 2358 903 2364 904
rect 2438 908 2444 909
rect 2438 904 2439 908
rect 2443 904 2444 908
rect 2438 903 2444 904
rect 2518 908 2524 909
rect 2518 904 2519 908
rect 2523 904 2524 908
rect 2518 903 2524 904
rect 2606 908 2612 909
rect 2606 904 2607 908
rect 2611 904 2612 908
rect 2606 903 2612 904
rect 2702 908 2708 909
rect 2702 904 2703 908
rect 2707 904 2708 908
rect 2702 903 2708 904
rect 1870 900 1876 901
rect 2346 899 2352 900
rect 2346 895 2347 899
rect 2351 895 2352 899
rect 2346 894 2352 895
rect 2430 899 2436 900
rect 2430 895 2431 899
rect 2435 895 2436 899
rect 2430 894 2436 895
rect 2506 899 2512 900
rect 2506 895 2507 899
rect 2511 895 2512 899
rect 2506 894 2512 895
rect 2586 899 2592 900
rect 2586 895 2587 899
rect 2591 895 2592 899
rect 2586 894 2592 895
rect 2674 899 2680 900
rect 2674 895 2675 899
rect 2679 895 2680 899
rect 2674 894 2680 895
rect 2338 891 2344 892
rect 1870 888 1876 889
rect 1870 884 1871 888
rect 1875 884 1876 888
rect 2338 887 2339 891
rect 2343 887 2344 891
rect 2338 886 2344 887
rect 1870 883 1876 884
rect 1231 874 1235 875
rect 1231 869 1235 870
rect 1279 874 1283 875
rect 1286 871 1287 875
rect 1291 871 1292 875
rect 1286 870 1292 871
rect 1335 874 1339 875
rect 1279 869 1283 870
rect 1280 859 1282 869
rect 1278 858 1284 859
rect 1278 854 1279 858
rect 1283 854 1284 858
rect 1278 853 1284 854
rect 1288 832 1290 870
rect 1335 869 1339 870
rect 1399 874 1403 875
rect 1399 869 1403 870
rect 1519 874 1523 875
rect 1519 869 1523 870
rect 1647 874 1651 875
rect 1647 869 1651 870
rect 1831 874 1835 875
rect 1831 869 1835 870
rect 1400 859 1402 869
rect 1406 867 1412 868
rect 1406 863 1407 867
rect 1411 863 1412 867
rect 1406 862 1412 863
rect 1398 858 1404 859
rect 1398 854 1399 858
rect 1403 854 1404 858
rect 1398 853 1404 854
rect 1408 832 1410 862
rect 1520 859 1522 869
rect 1526 867 1532 868
rect 1526 863 1527 867
rect 1531 863 1532 867
rect 1526 862 1532 863
rect 1518 858 1524 859
rect 1518 854 1519 858
rect 1523 854 1524 858
rect 1518 853 1524 854
rect 1528 832 1530 862
rect 1648 859 1650 869
rect 1654 867 1660 868
rect 1654 863 1655 867
rect 1659 863 1660 867
rect 1654 862 1660 863
rect 1710 867 1716 868
rect 1710 863 1711 867
rect 1715 863 1716 867
rect 1710 862 1716 863
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 1646 853 1652 854
rect 1656 832 1658 862
rect 1106 831 1112 832
rect 1106 827 1107 831
rect 1111 827 1112 831
rect 1106 826 1112 827
rect 1202 831 1208 832
rect 1202 827 1203 831
rect 1207 827 1208 831
rect 1202 826 1208 827
rect 1286 831 1292 832
rect 1286 827 1287 831
rect 1291 827 1292 831
rect 1286 826 1292 827
rect 1406 831 1412 832
rect 1406 827 1407 831
rect 1411 827 1412 831
rect 1406 826 1412 827
rect 1526 831 1532 832
rect 1526 827 1527 831
rect 1531 827 1532 831
rect 1526 826 1532 827
rect 1654 831 1660 832
rect 1654 827 1655 831
rect 1659 827 1660 831
rect 1654 826 1660 827
rect 1006 820 1012 821
rect 1006 816 1007 820
rect 1011 816 1012 820
rect 1006 815 1012 816
rect 1142 820 1148 821
rect 1142 816 1143 820
rect 1147 816 1148 820
rect 1142 815 1148 816
rect 1270 820 1276 821
rect 1270 816 1271 820
rect 1275 816 1276 820
rect 1270 815 1276 816
rect 1390 820 1396 821
rect 1390 816 1391 820
rect 1395 816 1396 820
rect 1390 815 1396 816
rect 1510 820 1516 821
rect 1510 816 1511 820
rect 1515 816 1516 820
rect 1510 815 1516 816
rect 1638 820 1644 821
rect 1638 816 1639 820
rect 1643 816 1644 820
rect 1638 815 1644 816
rect 1008 787 1010 815
rect 1144 787 1146 815
rect 1272 787 1274 815
rect 1392 787 1394 815
rect 1512 787 1514 815
rect 1640 787 1642 815
rect 951 786 955 787
rect 951 781 955 782
rect 1007 786 1011 787
rect 1007 781 1011 782
rect 1103 786 1107 787
rect 1103 781 1107 782
rect 1143 786 1147 787
rect 1143 781 1147 782
rect 1247 786 1251 787
rect 1247 781 1251 782
rect 1271 786 1275 787
rect 1271 781 1275 782
rect 1383 786 1387 787
rect 1383 781 1387 782
rect 1391 786 1395 787
rect 1391 781 1395 782
rect 1511 786 1515 787
rect 1511 781 1515 782
rect 1639 786 1643 787
rect 1639 781 1643 782
rect 952 765 954 781
rect 1104 765 1106 781
rect 1248 765 1250 781
rect 1384 765 1386 781
rect 1512 765 1514 781
rect 1640 765 1642 781
rect 950 764 956 765
rect 950 760 951 764
rect 955 760 956 764
rect 950 759 956 760
rect 1102 764 1108 765
rect 1102 760 1103 764
rect 1107 760 1108 764
rect 1102 759 1108 760
rect 1246 764 1252 765
rect 1246 760 1247 764
rect 1251 760 1252 764
rect 1246 759 1252 760
rect 1382 764 1388 765
rect 1382 760 1383 764
rect 1387 760 1388 764
rect 1382 759 1388 760
rect 1510 764 1516 765
rect 1510 760 1511 764
rect 1515 760 1516 764
rect 1510 759 1516 760
rect 1638 764 1644 765
rect 1638 760 1639 764
rect 1643 760 1644 764
rect 1638 759 1644 760
rect 1712 756 1714 862
rect 1832 841 1834 869
rect 1872 843 1874 883
rect 2286 870 2292 871
rect 2286 866 2287 870
rect 2291 866 2292 870
rect 2286 865 2292 866
rect 2288 843 2290 865
rect 2340 860 2342 886
rect 2348 860 2350 894
rect 2366 870 2372 871
rect 2366 866 2367 870
rect 2371 866 2372 870
rect 2366 865 2372 866
rect 2338 859 2344 860
rect 2338 855 2339 859
rect 2343 855 2344 859
rect 2338 854 2344 855
rect 2346 859 2352 860
rect 2346 855 2347 859
rect 2351 855 2352 859
rect 2346 854 2352 855
rect 2334 843 2340 844
rect 2368 843 2370 865
rect 1871 842 1875 843
rect 1830 840 1836 841
rect 1830 836 1831 840
rect 1835 836 1836 840
rect 1871 837 1875 838
rect 2167 842 2171 843
rect 2167 837 2171 838
rect 2247 842 2251 843
rect 2247 837 2251 838
rect 2287 842 2291 843
rect 2287 837 2291 838
rect 2327 842 2331 843
rect 2334 839 2335 843
rect 2339 839 2340 843
rect 2334 838 2340 839
rect 2367 842 2371 843
rect 2327 837 2331 838
rect 1830 835 1836 836
rect 1830 823 1836 824
rect 1830 819 1831 823
rect 1835 819 1836 823
rect 1830 818 1836 819
rect 1832 787 1834 818
rect 1872 809 1874 837
rect 2168 827 2170 837
rect 2218 835 2224 836
rect 2218 831 2219 835
rect 2223 831 2224 835
rect 2218 830 2224 831
rect 2166 826 2172 827
rect 2166 822 2167 826
rect 2171 822 2172 826
rect 2166 821 2172 822
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 2220 800 2222 830
rect 2248 827 2250 837
rect 2328 827 2330 837
rect 2246 826 2252 827
rect 2246 822 2247 826
rect 2251 822 2252 826
rect 2246 821 2252 822
rect 2326 826 2332 827
rect 2326 822 2327 826
rect 2331 822 2332 826
rect 2326 821 2332 822
rect 2336 800 2338 838
rect 2367 837 2371 838
rect 2423 842 2427 843
rect 2423 837 2427 838
rect 2424 827 2426 837
rect 2432 836 2434 894
rect 2446 870 2452 871
rect 2446 866 2447 870
rect 2451 866 2452 870
rect 2446 865 2452 866
rect 2448 843 2450 865
rect 2508 860 2510 894
rect 2526 870 2532 871
rect 2526 866 2527 870
rect 2531 866 2532 870
rect 2526 865 2532 866
rect 2506 859 2512 860
rect 2506 855 2507 859
rect 2511 855 2512 859
rect 2506 854 2512 855
rect 2528 843 2530 865
rect 2588 860 2590 894
rect 2614 870 2620 871
rect 2614 866 2615 870
rect 2619 866 2620 870
rect 2614 865 2620 866
rect 2586 859 2592 860
rect 2586 855 2587 859
rect 2591 855 2592 859
rect 2586 854 2592 855
rect 2616 843 2618 865
rect 2676 860 2678 894
rect 2710 870 2716 871
rect 2710 866 2711 870
rect 2715 866 2716 870
rect 2710 865 2716 866
rect 2674 859 2680 860
rect 2674 855 2675 859
rect 2679 855 2680 859
rect 2674 854 2680 855
rect 2662 843 2668 844
rect 2712 843 2714 865
rect 2724 860 2726 966
rect 2774 960 2780 961
rect 2774 956 2775 960
rect 2779 956 2780 960
rect 2774 955 2780 956
rect 2902 960 2908 961
rect 2902 956 2903 960
rect 2907 956 2908 960
rect 2902 955 2908 956
rect 3046 960 3052 961
rect 3046 956 3047 960
rect 3051 956 3052 960
rect 3046 955 3052 956
rect 2776 931 2778 955
rect 2842 943 2848 944
rect 2842 939 2843 943
rect 2847 939 2848 943
rect 2842 938 2848 939
rect 2775 930 2779 931
rect 2775 925 2779 926
rect 2807 930 2811 931
rect 2807 925 2811 926
rect 2808 909 2810 925
rect 2806 908 2812 909
rect 2806 904 2807 908
rect 2811 904 2812 908
rect 2806 903 2812 904
rect 2814 870 2820 871
rect 2814 866 2815 870
rect 2819 866 2820 870
rect 2814 865 2820 866
rect 2722 859 2728 860
rect 2722 855 2723 859
rect 2727 855 2728 859
rect 2722 854 2728 855
rect 2816 843 2818 865
rect 2844 860 2846 938
rect 2904 931 2906 955
rect 3048 931 3050 955
rect 2903 930 2907 931
rect 2903 925 2907 926
rect 2911 930 2915 931
rect 2911 925 2915 926
rect 3015 930 3019 931
rect 3015 925 3019 926
rect 3047 930 3051 931
rect 3047 925 3051 926
rect 2912 909 2914 925
rect 3016 909 3018 925
rect 2910 908 2916 909
rect 2910 904 2911 908
rect 2915 904 2916 908
rect 2910 903 2916 904
rect 3014 908 3020 909
rect 3014 904 3015 908
rect 3019 904 3020 908
rect 3014 903 3020 904
rect 2890 899 2896 900
rect 2890 895 2891 899
rect 2895 895 2896 899
rect 2890 894 2896 895
rect 2918 895 2924 896
rect 2892 860 2894 894
rect 2918 891 2919 895
rect 2923 891 2924 895
rect 3076 892 3078 1002
rect 3108 972 3110 1002
rect 3208 999 3210 1009
rect 3258 1007 3264 1008
rect 3258 1003 3259 1007
rect 3263 1003 3264 1007
rect 3258 1002 3264 1003
rect 3206 998 3212 999
rect 3206 994 3207 998
rect 3211 994 3212 998
rect 3206 993 3212 994
rect 3260 972 3262 1002
rect 3368 999 3370 1009
rect 3366 998 3372 999
rect 3366 994 3367 998
rect 3371 994 3372 998
rect 3366 993 3372 994
rect 3400 972 3402 1014
rect 3511 1009 3515 1010
rect 3512 999 3514 1009
rect 3564 1008 3566 1046
rect 3590 1044 3591 1048
rect 3595 1044 3596 1048
rect 3590 1043 3596 1044
rect 3592 1015 3594 1043
rect 3591 1014 3595 1015
rect 3591 1009 3595 1010
rect 3562 1007 3568 1008
rect 3562 1003 3563 1007
rect 3567 1003 3568 1007
rect 3562 1002 3568 1003
rect 3510 998 3516 999
rect 3510 994 3511 998
rect 3515 994 3516 998
rect 3510 993 3516 994
rect 3592 981 3594 1009
rect 3590 980 3596 981
rect 3590 976 3591 980
rect 3595 976 3596 980
rect 3590 975 3596 976
rect 3106 971 3112 972
rect 3106 967 3107 971
rect 3111 967 3112 971
rect 3106 966 3112 967
rect 3258 971 3264 972
rect 3258 967 3259 971
rect 3263 967 3264 971
rect 3258 966 3264 967
rect 3398 971 3404 972
rect 3398 967 3399 971
rect 3403 967 3404 971
rect 3398 966 3404 967
rect 3534 971 3540 972
rect 3534 967 3535 971
rect 3539 967 3540 971
rect 3534 966 3540 967
rect 3198 960 3204 961
rect 3198 956 3199 960
rect 3203 956 3204 960
rect 3198 955 3204 956
rect 3358 960 3364 961
rect 3358 956 3359 960
rect 3363 956 3364 960
rect 3358 955 3364 956
rect 3502 960 3508 961
rect 3502 956 3503 960
rect 3507 956 3508 960
rect 3502 955 3508 956
rect 3200 931 3202 955
rect 3360 931 3362 955
rect 3504 931 3506 955
rect 3111 930 3115 931
rect 3111 925 3115 926
rect 3199 930 3203 931
rect 3199 925 3203 926
rect 3215 930 3219 931
rect 3215 925 3219 926
rect 3319 930 3323 931
rect 3319 925 3323 926
rect 3359 930 3363 931
rect 3359 925 3363 926
rect 3423 930 3427 931
rect 3423 925 3427 926
rect 3503 930 3507 931
rect 3503 925 3507 926
rect 3112 909 3114 925
rect 3216 909 3218 925
rect 3320 909 3322 925
rect 3424 909 3426 925
rect 3504 909 3506 925
rect 3110 908 3116 909
rect 3110 904 3111 908
rect 3115 904 3116 908
rect 3110 903 3116 904
rect 3214 908 3220 909
rect 3214 904 3215 908
rect 3219 904 3220 908
rect 3214 903 3220 904
rect 3318 908 3324 909
rect 3318 904 3319 908
rect 3323 904 3324 908
rect 3318 903 3324 904
rect 3422 908 3428 909
rect 3422 904 3423 908
rect 3427 904 3428 908
rect 3422 903 3428 904
rect 3502 908 3508 909
rect 3502 904 3503 908
rect 3507 904 3508 908
rect 3502 903 3508 904
rect 3082 899 3088 900
rect 3082 895 3083 899
rect 3087 895 3088 899
rect 3082 894 3088 895
rect 3178 899 3184 900
rect 3178 895 3179 899
rect 3183 895 3184 899
rect 3178 894 3184 895
rect 3282 899 3288 900
rect 3282 895 3283 899
rect 3287 895 3288 899
rect 3282 894 3288 895
rect 3490 899 3496 900
rect 3490 895 3491 899
rect 3495 895 3496 899
rect 3490 894 3496 895
rect 2918 890 2924 891
rect 3074 891 3080 892
rect 2920 875 2922 890
rect 3074 887 3075 891
rect 3079 887 3080 891
rect 3074 886 3080 887
rect 2920 873 2930 875
rect 2918 870 2924 871
rect 2918 866 2919 870
rect 2923 866 2924 870
rect 2918 865 2924 866
rect 2842 859 2848 860
rect 2842 855 2843 859
rect 2847 855 2848 859
rect 2842 854 2848 855
rect 2890 859 2896 860
rect 2890 855 2891 859
rect 2895 855 2896 859
rect 2890 854 2896 855
rect 2920 843 2922 865
rect 2447 842 2451 843
rect 2447 837 2451 838
rect 2527 842 2531 843
rect 2527 837 2531 838
rect 2535 842 2539 843
rect 2535 837 2539 838
rect 2615 842 2619 843
rect 2615 837 2619 838
rect 2655 842 2659 843
rect 2662 839 2663 843
rect 2667 839 2668 843
rect 2662 838 2668 839
rect 2711 842 2715 843
rect 2655 837 2659 838
rect 2430 835 2436 836
rect 2430 831 2431 835
rect 2435 831 2436 835
rect 2430 830 2436 831
rect 2474 835 2480 836
rect 2474 831 2475 835
rect 2479 831 2480 835
rect 2474 830 2480 831
rect 2422 826 2428 827
rect 2422 822 2423 826
rect 2427 822 2428 826
rect 2422 821 2428 822
rect 2476 800 2478 830
rect 2536 827 2538 837
rect 2586 835 2592 836
rect 2586 831 2587 835
rect 2591 831 2592 835
rect 2586 830 2592 831
rect 2534 826 2540 827
rect 2534 822 2535 826
rect 2539 822 2540 826
rect 2534 821 2540 822
rect 2588 800 2590 830
rect 2656 827 2658 837
rect 2654 826 2660 827
rect 2654 822 2655 826
rect 2659 822 2660 826
rect 2654 821 2660 822
rect 2664 800 2666 838
rect 2711 837 2715 838
rect 2783 842 2787 843
rect 2783 837 2787 838
rect 2815 842 2819 843
rect 2815 837 2819 838
rect 2911 842 2915 843
rect 2911 837 2915 838
rect 2919 842 2923 843
rect 2919 837 2923 838
rect 2784 827 2786 837
rect 2858 835 2864 836
rect 2858 831 2859 835
rect 2863 831 2864 835
rect 2858 830 2864 831
rect 2782 826 2788 827
rect 2782 822 2783 826
rect 2787 822 2788 826
rect 2782 821 2788 822
rect 2860 800 2862 830
rect 2912 827 2914 837
rect 2928 836 2930 873
rect 3022 870 3028 871
rect 3022 866 3023 870
rect 3027 866 3028 870
rect 3022 865 3028 866
rect 3024 843 3026 865
rect 3084 860 3086 894
rect 3118 870 3124 871
rect 3118 866 3119 870
rect 3123 866 3124 870
rect 3118 865 3124 866
rect 3082 859 3088 860
rect 3082 855 3083 859
rect 3087 855 3088 859
rect 3082 854 3088 855
rect 3120 843 3122 865
rect 3180 860 3182 894
rect 3222 870 3228 871
rect 3222 866 3223 870
rect 3227 866 3228 870
rect 3222 865 3228 866
rect 3178 859 3184 860
rect 3178 855 3179 859
rect 3183 855 3184 859
rect 3178 854 3184 855
rect 3224 843 3226 865
rect 3284 860 3286 894
rect 3482 891 3488 892
rect 3482 887 3483 891
rect 3487 887 3488 891
rect 3482 886 3488 887
rect 3326 870 3332 871
rect 3326 866 3327 870
rect 3331 866 3332 870
rect 3326 865 3332 866
rect 3430 870 3436 871
rect 3430 866 3431 870
rect 3435 866 3436 870
rect 3430 865 3436 866
rect 3282 859 3288 860
rect 3282 855 3283 859
rect 3287 855 3288 859
rect 3282 854 3288 855
rect 3328 843 3330 865
rect 3414 859 3420 860
rect 3414 855 3415 859
rect 3419 855 3420 859
rect 3414 854 3420 855
rect 3023 842 3027 843
rect 3023 837 3027 838
rect 3039 842 3043 843
rect 3039 837 3043 838
rect 3119 842 3123 843
rect 3119 837 3123 838
rect 3159 842 3163 843
rect 3159 837 3163 838
rect 3223 842 3227 843
rect 3223 837 3227 838
rect 3279 842 3283 843
rect 3279 837 3283 838
rect 3327 842 3331 843
rect 3327 837 3331 838
rect 3407 842 3411 843
rect 3407 837 3411 838
rect 2926 835 2932 836
rect 2926 831 2927 835
rect 2931 831 2932 835
rect 2926 830 2932 831
rect 3040 827 3042 837
rect 3054 835 3060 836
rect 3054 831 3055 835
rect 3059 831 3060 835
rect 3054 830 3060 831
rect 3090 835 3096 836
rect 3090 831 3091 835
rect 3095 831 3096 835
rect 3090 830 3096 831
rect 2910 826 2916 827
rect 2910 822 2911 826
rect 2915 822 2916 826
rect 2910 821 2916 822
rect 3038 826 3044 827
rect 3038 822 3039 826
rect 3043 822 3044 826
rect 3038 821 3044 822
rect 2218 799 2224 800
rect 2218 795 2219 799
rect 2223 795 2224 799
rect 2218 794 2224 795
rect 2298 799 2304 800
rect 2298 795 2299 799
rect 2303 795 2304 799
rect 2298 794 2304 795
rect 2334 799 2340 800
rect 2334 795 2335 799
rect 2339 795 2340 799
rect 2334 794 2340 795
rect 2474 799 2480 800
rect 2474 795 2475 799
rect 2479 795 2480 799
rect 2474 794 2480 795
rect 2586 799 2592 800
rect 2586 795 2587 799
rect 2591 795 2592 799
rect 2586 794 2592 795
rect 2662 799 2668 800
rect 2662 795 2663 799
rect 2667 795 2668 799
rect 2662 794 2668 795
rect 2834 799 2840 800
rect 2834 795 2835 799
rect 2839 795 2840 799
rect 2834 794 2840 795
rect 2858 799 2864 800
rect 2858 795 2859 799
rect 2863 795 2864 799
rect 2858 794 2864 795
rect 1870 791 1876 792
rect 1870 787 1871 791
rect 1875 787 1876 791
rect 1743 786 1747 787
rect 1743 781 1747 782
rect 1831 786 1835 787
rect 1870 786 1876 787
rect 2158 788 2164 789
rect 1831 781 1835 782
rect 1744 765 1746 781
rect 1742 764 1748 765
rect 1742 760 1743 764
rect 1747 760 1748 764
rect 1832 762 1834 781
rect 1742 759 1748 760
rect 1830 761 1836 762
rect 1830 757 1831 761
rect 1835 757 1836 761
rect 1872 759 1874 786
rect 2158 784 2159 788
rect 2163 784 2164 788
rect 2158 783 2164 784
rect 2238 788 2244 789
rect 2238 784 2239 788
rect 2243 784 2244 788
rect 2238 783 2244 784
rect 2160 759 2162 783
rect 2240 759 2242 783
rect 1830 756 1836 757
rect 1871 758 1875 759
rect 1210 755 1216 756
rect 1210 751 1211 755
rect 1215 751 1216 755
rect 1210 750 1216 751
rect 1338 755 1344 756
rect 1338 751 1339 755
rect 1343 751 1344 755
rect 1338 750 1344 751
rect 1470 755 1476 756
rect 1470 751 1471 755
rect 1475 751 1476 755
rect 1470 750 1476 751
rect 1598 755 1604 756
rect 1598 751 1599 755
rect 1603 751 1604 755
rect 1598 750 1604 751
rect 1710 755 1716 756
rect 1710 751 1711 755
rect 1715 751 1716 755
rect 1871 753 1875 754
rect 1895 758 1899 759
rect 1895 753 1899 754
rect 1975 758 1979 759
rect 1975 753 1979 754
rect 2071 758 2075 759
rect 2071 753 2075 754
rect 2159 758 2163 759
rect 2159 753 2163 754
rect 2183 758 2187 759
rect 2183 753 2187 754
rect 2239 758 2243 759
rect 2239 753 2243 754
rect 1710 750 1716 751
rect 886 747 892 748
rect 886 743 887 747
rect 891 743 892 747
rect 886 742 892 743
rect 958 726 964 727
rect 958 722 959 726
rect 963 722 964 726
rect 958 721 964 722
rect 1110 726 1116 727
rect 1110 722 1111 726
rect 1115 722 1116 726
rect 1110 721 1116 722
rect 850 715 856 716
rect 850 711 851 715
rect 855 711 856 715
rect 850 710 856 711
rect 960 699 962 721
rect 966 715 972 716
rect 966 711 967 715
rect 971 711 972 715
rect 966 710 972 711
rect 407 698 411 699
rect 407 693 411 694
rect 439 698 443 699
rect 439 693 443 694
rect 527 698 531 699
rect 527 693 531 694
rect 615 698 619 699
rect 615 693 619 694
rect 655 698 659 699
rect 655 693 659 694
rect 783 698 787 699
rect 783 693 787 694
rect 791 698 795 699
rect 791 693 795 694
rect 903 698 907 699
rect 903 693 907 694
rect 959 698 963 699
rect 959 693 963 694
rect 322 691 328 692
rect 322 687 323 691
rect 327 687 328 691
rect 322 686 328 687
rect 346 691 352 692
rect 346 687 347 691
rect 351 687 352 691
rect 346 686 352 687
rect 294 682 300 683
rect 294 678 295 682
rect 299 678 300 682
rect 294 677 300 678
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 348 656 350 686
rect 408 683 410 693
rect 458 691 464 692
rect 458 687 459 691
rect 463 687 464 691
rect 458 686 464 687
rect 406 682 412 683
rect 406 678 407 682
rect 411 678 412 682
rect 406 677 412 678
rect 460 656 462 686
rect 528 683 530 693
rect 656 683 658 693
rect 714 691 720 692
rect 714 687 715 691
rect 719 687 720 691
rect 714 686 720 687
rect 774 691 780 692
rect 774 687 775 691
rect 779 687 780 691
rect 774 686 780 687
rect 526 682 532 683
rect 526 678 527 682
rect 531 678 532 682
rect 526 677 532 678
rect 654 682 660 683
rect 654 678 655 682
rect 659 678 660 682
rect 654 677 660 678
rect 346 655 352 656
rect 346 651 347 655
rect 351 651 352 655
rect 346 650 352 651
rect 458 655 464 656
rect 458 651 459 655
rect 463 651 464 655
rect 458 650 464 651
rect 578 655 584 656
rect 578 651 579 655
rect 583 651 584 655
rect 578 650 584 651
rect 110 647 116 648
rect 110 643 111 647
rect 115 643 116 647
rect 110 642 116 643
rect 286 644 292 645
rect 112 619 114 642
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 398 644 404 645
rect 398 640 399 644
rect 403 640 404 644
rect 398 639 404 640
rect 518 644 524 645
rect 518 640 519 644
rect 523 640 524 644
rect 518 639 524 640
rect 288 619 290 639
rect 400 619 402 639
rect 520 619 522 639
rect 111 618 115 619
rect 111 613 115 614
rect 287 618 291 619
rect 287 613 291 614
rect 311 618 315 619
rect 311 613 315 614
rect 391 618 395 619
rect 391 613 395 614
rect 399 618 403 619
rect 399 613 403 614
rect 471 618 475 619
rect 471 613 475 614
rect 519 618 523 619
rect 519 613 523 614
rect 559 618 563 619
rect 559 613 563 614
rect 112 594 114 613
rect 312 597 314 613
rect 392 597 394 613
rect 472 597 474 613
rect 560 597 562 613
rect 310 596 316 597
rect 110 593 116 594
rect 110 589 111 593
rect 115 589 116 593
rect 310 592 311 596
rect 315 592 316 596
rect 310 591 316 592
rect 390 596 396 597
rect 390 592 391 596
rect 395 592 396 596
rect 390 591 396 592
rect 470 596 476 597
rect 470 592 471 596
rect 475 592 476 596
rect 470 591 476 592
rect 558 596 564 597
rect 558 592 559 596
rect 563 592 564 596
rect 558 591 564 592
rect 110 588 116 589
rect 266 587 272 588
rect 266 583 267 587
rect 271 583 272 587
rect 266 582 272 583
rect 378 587 384 588
rect 378 583 379 587
rect 383 583 384 587
rect 378 582 384 583
rect 458 587 464 588
rect 458 583 459 587
rect 463 583 464 587
rect 458 582 464 583
rect 538 587 544 588
rect 538 583 539 587
rect 543 583 544 587
rect 538 582 544 583
rect 110 576 116 577
rect 110 572 111 576
rect 115 572 116 576
rect 110 571 116 572
rect 112 531 114 571
rect 111 530 115 531
rect 111 525 115 526
rect 239 530 243 531
rect 239 525 243 526
rect 112 497 114 525
rect 240 515 242 525
rect 268 524 270 582
rect 318 558 324 559
rect 318 554 319 558
rect 323 554 324 558
rect 318 553 324 554
rect 320 531 322 553
rect 380 548 382 582
rect 398 558 404 559
rect 398 554 399 558
rect 403 554 404 558
rect 398 553 404 554
rect 378 547 384 548
rect 378 543 379 547
rect 383 543 384 547
rect 378 542 384 543
rect 400 531 402 553
rect 460 548 462 582
rect 478 558 484 559
rect 478 554 479 558
rect 483 554 484 558
rect 478 553 484 554
rect 458 547 464 548
rect 458 543 459 547
rect 463 543 464 547
rect 458 542 464 543
rect 480 531 482 553
rect 540 548 542 582
rect 566 558 572 559
rect 566 554 567 558
rect 571 554 572 558
rect 566 553 572 554
rect 538 547 544 548
rect 538 543 539 547
rect 543 543 544 547
rect 538 542 544 543
rect 568 531 570 553
rect 580 548 582 650
rect 646 644 652 645
rect 646 640 647 644
rect 651 640 652 644
rect 646 639 652 640
rect 648 619 650 639
rect 647 618 651 619
rect 647 613 651 614
rect 648 597 650 613
rect 646 596 652 597
rect 646 592 647 596
rect 651 592 652 596
rect 646 591 652 592
rect 716 588 718 686
rect 776 656 778 686
rect 784 683 786 693
rect 834 691 840 692
rect 834 687 835 691
rect 839 687 840 691
rect 834 686 840 687
rect 782 682 788 683
rect 782 678 783 682
rect 787 678 788 682
rect 782 677 788 678
rect 836 656 838 686
rect 904 683 906 693
rect 902 682 908 683
rect 902 678 903 682
rect 907 678 908 682
rect 902 677 908 678
rect 968 656 970 710
rect 1112 699 1114 721
rect 1212 716 1214 750
rect 1254 726 1260 727
rect 1254 722 1255 726
rect 1259 722 1260 726
rect 1254 721 1260 722
rect 1198 715 1204 716
rect 1198 711 1199 715
rect 1203 711 1204 715
rect 1198 710 1204 711
rect 1210 715 1216 716
rect 1210 711 1211 715
rect 1215 711 1216 715
rect 1210 710 1216 711
rect 1023 698 1027 699
rect 1023 693 1027 694
rect 1111 698 1115 699
rect 1111 693 1115 694
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1024 683 1026 693
rect 1058 691 1064 692
rect 1058 687 1059 691
rect 1063 687 1064 691
rect 1058 686 1064 687
rect 1074 691 1080 692
rect 1074 687 1075 691
rect 1079 687 1080 691
rect 1074 686 1080 687
rect 1022 682 1028 683
rect 1022 678 1023 682
rect 1027 678 1028 682
rect 1022 677 1028 678
rect 774 655 780 656
rect 774 651 775 655
rect 779 651 780 655
rect 774 650 780 651
rect 834 655 840 656
rect 834 651 835 655
rect 839 651 840 655
rect 834 650 840 651
rect 966 655 972 656
rect 966 651 967 655
rect 971 651 972 655
rect 966 650 972 651
rect 774 644 780 645
rect 774 640 775 644
rect 779 640 780 644
rect 774 639 780 640
rect 894 644 900 645
rect 894 640 895 644
rect 899 640 900 644
rect 894 639 900 640
rect 1014 644 1020 645
rect 1014 640 1015 644
rect 1019 640 1020 644
rect 1014 639 1020 640
rect 776 619 778 639
rect 896 619 898 639
rect 1016 619 1018 639
rect 735 618 739 619
rect 735 613 739 614
rect 775 618 779 619
rect 775 613 779 614
rect 823 618 827 619
rect 823 613 827 614
rect 895 618 899 619
rect 895 613 899 614
rect 911 618 915 619
rect 911 613 915 614
rect 999 618 1003 619
rect 999 613 1003 614
rect 1015 618 1019 619
rect 1015 613 1019 614
rect 736 597 738 613
rect 824 597 826 613
rect 912 597 914 613
rect 1000 597 1002 613
rect 734 596 740 597
rect 734 592 735 596
rect 739 592 740 596
rect 734 591 740 592
rect 822 596 828 597
rect 822 592 823 596
rect 827 592 828 596
rect 822 591 828 592
rect 910 596 916 597
rect 910 592 911 596
rect 915 592 916 596
rect 910 591 916 592
rect 998 596 1004 597
rect 998 592 999 596
rect 1003 592 1004 596
rect 998 591 1004 592
rect 714 587 720 588
rect 714 583 715 587
rect 719 583 720 587
rect 714 582 720 583
rect 890 587 896 588
rect 890 583 891 587
rect 895 583 896 587
rect 890 582 896 583
rect 978 587 984 588
rect 978 583 979 587
rect 983 583 984 587
rect 978 582 984 583
rect 706 579 712 580
rect 706 575 707 579
rect 711 575 712 579
rect 706 574 712 575
rect 654 558 660 559
rect 654 554 655 558
rect 659 554 660 558
rect 654 553 660 554
rect 578 547 584 548
rect 578 543 579 547
rect 583 543 584 547
rect 578 542 584 543
rect 622 547 628 548
rect 622 543 623 547
rect 627 543 628 547
rect 622 542 628 543
rect 319 530 323 531
rect 319 525 323 526
rect 343 530 347 531
rect 343 525 347 526
rect 399 530 403 531
rect 399 525 403 526
rect 439 530 443 531
rect 439 525 443 526
rect 479 530 483 531
rect 479 525 483 526
rect 535 530 539 531
rect 535 525 539 526
rect 567 530 571 531
rect 567 525 571 526
rect 266 523 272 524
rect 266 519 267 523
rect 271 519 272 523
rect 266 518 272 519
rect 290 523 296 524
rect 290 519 291 523
rect 295 519 296 523
rect 290 518 296 519
rect 238 514 244 515
rect 238 510 239 514
rect 243 510 244 514
rect 238 509 244 510
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 292 488 294 518
rect 344 515 346 525
rect 440 515 442 525
rect 466 523 472 524
rect 466 519 467 523
rect 471 519 472 523
rect 466 518 472 519
rect 490 523 496 524
rect 490 519 491 523
rect 495 519 496 523
rect 490 518 496 519
rect 342 514 348 515
rect 342 510 343 514
rect 347 510 348 514
rect 342 509 348 510
rect 438 514 444 515
rect 438 510 439 514
rect 443 510 444 514
rect 438 509 444 510
rect 290 487 296 488
rect 290 483 291 487
rect 295 483 296 487
rect 290 482 296 483
rect 394 487 400 488
rect 394 483 395 487
rect 399 483 400 487
rect 394 482 400 483
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 230 476 236 477
rect 112 447 114 474
rect 230 472 231 476
rect 235 472 236 476
rect 230 471 236 472
rect 334 476 340 477
rect 334 472 335 476
rect 339 472 340 476
rect 334 471 340 472
rect 232 447 234 471
rect 336 447 338 471
rect 111 446 115 447
rect 111 441 115 442
rect 135 446 139 447
rect 135 441 139 442
rect 231 446 235 447
rect 231 441 235 442
rect 247 446 251 447
rect 247 441 251 442
rect 335 446 339 447
rect 335 441 339 442
rect 375 446 379 447
rect 375 441 379 442
rect 112 422 114 441
rect 136 425 138 441
rect 248 425 250 441
rect 376 425 378 441
rect 134 424 140 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 134 420 135 424
rect 139 420 140 424
rect 134 419 140 420
rect 246 424 252 425
rect 246 420 247 424
rect 251 420 252 424
rect 246 419 252 420
rect 374 424 380 425
rect 374 420 375 424
rect 379 420 380 424
rect 374 419 380 420
rect 110 416 116 417
rect 202 415 208 416
rect 202 411 203 415
rect 207 411 208 415
rect 202 410 208 411
rect 314 415 320 416
rect 314 411 315 415
rect 319 411 320 415
rect 314 410 320 411
rect 194 407 200 408
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 194 403 195 407
rect 199 403 200 407
rect 194 402 200 403
rect 110 399 116 400
rect 112 359 114 399
rect 142 386 148 387
rect 142 382 143 386
rect 147 382 148 386
rect 142 381 148 382
rect 144 359 146 381
rect 111 358 115 359
rect 111 353 115 354
rect 143 358 147 359
rect 143 353 147 354
rect 112 325 114 353
rect 144 343 146 353
rect 196 352 198 402
rect 204 376 206 410
rect 254 386 260 387
rect 254 382 255 386
rect 259 382 260 386
rect 254 381 260 382
rect 202 375 208 376
rect 202 371 203 375
rect 207 371 208 375
rect 202 370 208 371
rect 256 359 258 381
rect 316 376 318 410
rect 382 386 388 387
rect 382 382 383 386
rect 387 382 388 386
rect 382 381 388 382
rect 314 375 320 376
rect 314 371 315 375
rect 319 371 320 375
rect 314 370 320 371
rect 384 359 386 381
rect 396 376 398 482
rect 430 476 436 477
rect 430 472 431 476
rect 435 472 436 476
rect 430 471 436 472
rect 432 447 434 471
rect 431 446 435 447
rect 431 441 435 442
rect 468 416 470 518
rect 492 488 494 518
rect 536 515 538 525
rect 534 514 540 515
rect 534 510 535 514
rect 539 510 540 514
rect 534 509 540 510
rect 624 488 626 542
rect 656 531 658 553
rect 708 548 710 574
rect 742 558 748 559
rect 742 554 743 558
rect 747 554 748 558
rect 742 553 748 554
rect 830 558 836 559
rect 830 554 831 558
rect 835 554 836 558
rect 830 553 836 554
rect 706 547 712 548
rect 706 543 707 547
rect 711 543 712 547
rect 706 542 712 543
rect 744 531 746 553
rect 786 531 792 532
rect 832 531 834 553
rect 892 548 894 582
rect 918 558 924 559
rect 918 554 919 558
rect 923 554 924 558
rect 918 553 924 554
rect 882 547 888 548
rect 882 543 883 547
rect 887 543 888 547
rect 882 542 888 543
rect 890 547 896 548
rect 890 543 891 547
rect 895 543 896 547
rect 890 542 896 543
rect 631 530 635 531
rect 631 525 635 526
rect 655 530 659 531
rect 655 525 659 526
rect 719 530 723 531
rect 719 525 723 526
rect 743 530 747 531
rect 786 527 787 531
rect 791 527 792 531
rect 786 526 792 527
rect 807 530 811 531
rect 743 525 747 526
rect 632 515 634 525
rect 682 523 688 524
rect 682 519 683 523
rect 687 519 688 523
rect 682 518 688 519
rect 630 514 636 515
rect 630 510 631 514
rect 635 510 636 514
rect 630 509 636 510
rect 684 488 686 518
rect 720 515 722 525
rect 770 523 776 524
rect 770 519 771 523
rect 775 519 776 523
rect 770 518 776 519
rect 718 514 724 515
rect 718 510 719 514
rect 723 510 724 514
rect 718 509 724 510
rect 772 488 774 518
rect 490 487 496 488
rect 490 483 491 487
rect 495 483 496 487
rect 490 482 496 483
rect 622 487 628 488
rect 622 483 623 487
rect 627 483 628 487
rect 622 482 628 483
rect 682 487 688 488
rect 682 483 683 487
rect 687 483 688 487
rect 682 482 688 483
rect 770 487 776 488
rect 770 483 771 487
rect 775 483 776 487
rect 770 482 776 483
rect 526 476 532 477
rect 526 472 527 476
rect 531 472 532 476
rect 526 471 532 472
rect 622 476 628 477
rect 622 472 623 476
rect 627 472 628 476
rect 622 471 628 472
rect 710 476 716 477
rect 710 472 711 476
rect 715 472 716 476
rect 710 471 716 472
rect 528 447 530 471
rect 624 447 626 471
rect 712 447 714 471
rect 495 446 499 447
rect 495 441 499 442
rect 527 446 531 447
rect 527 441 531 442
rect 607 446 611 447
rect 607 441 611 442
rect 623 446 627 447
rect 623 441 627 442
rect 711 446 715 447
rect 711 441 715 442
rect 719 446 723 447
rect 719 441 723 442
rect 496 425 498 441
rect 608 425 610 441
rect 720 425 722 441
rect 494 424 500 425
rect 494 420 495 424
rect 499 420 500 424
rect 494 419 500 420
rect 606 424 612 425
rect 606 420 607 424
rect 611 420 612 424
rect 606 419 612 420
rect 718 424 724 425
rect 718 420 719 424
rect 723 420 724 424
rect 718 419 724 420
rect 788 416 790 526
rect 807 525 811 526
rect 831 530 835 531
rect 831 525 835 526
rect 808 515 810 525
rect 858 523 864 524
rect 858 519 859 523
rect 863 519 864 523
rect 858 518 864 519
rect 806 514 812 515
rect 806 510 807 514
rect 811 510 812 514
rect 806 509 812 510
rect 860 488 862 518
rect 884 517 886 542
rect 920 531 922 553
rect 980 548 982 582
rect 1060 580 1062 686
rect 1076 656 1078 686
rect 1136 683 1138 693
rect 1186 691 1192 692
rect 1186 687 1187 691
rect 1191 687 1192 691
rect 1186 686 1192 687
rect 1134 682 1140 683
rect 1134 678 1135 682
rect 1139 678 1140 682
rect 1134 677 1140 678
rect 1188 656 1190 686
rect 1200 685 1202 710
rect 1256 699 1258 721
rect 1340 716 1342 750
rect 1390 726 1396 727
rect 1390 722 1391 726
rect 1395 722 1396 726
rect 1390 721 1396 722
rect 1338 715 1344 716
rect 1338 711 1339 715
rect 1343 711 1344 715
rect 1338 710 1344 711
rect 1392 699 1394 721
rect 1472 716 1474 750
rect 1518 726 1524 727
rect 1518 722 1519 726
rect 1523 722 1524 726
rect 1518 721 1524 722
rect 1470 715 1476 716
rect 1470 711 1471 715
rect 1475 711 1476 715
rect 1470 710 1476 711
rect 1520 699 1522 721
rect 1600 716 1602 750
rect 1698 747 1704 748
rect 1698 743 1699 747
rect 1703 743 1704 747
rect 1698 742 1704 743
rect 1830 744 1836 745
rect 1646 726 1652 727
rect 1646 722 1647 726
rect 1651 722 1652 726
rect 1646 721 1652 722
rect 1598 715 1604 716
rect 1598 711 1599 715
rect 1603 711 1604 715
rect 1598 710 1604 711
rect 1648 699 1650 721
rect 1700 716 1702 742
rect 1830 740 1831 744
rect 1835 740 1836 744
rect 1830 739 1836 740
rect 1750 726 1756 727
rect 1750 722 1751 726
rect 1755 722 1756 726
rect 1750 721 1756 722
rect 1698 715 1704 716
rect 1698 711 1699 715
rect 1703 711 1704 715
rect 1698 710 1704 711
rect 1752 699 1754 721
rect 1832 699 1834 739
rect 1872 734 1874 753
rect 1896 737 1898 753
rect 1976 737 1978 753
rect 2072 737 2074 753
rect 2184 737 2186 753
rect 1894 736 1900 737
rect 1870 733 1876 734
rect 1870 729 1871 733
rect 1875 729 1876 733
rect 1894 732 1895 736
rect 1899 732 1900 736
rect 1894 731 1900 732
rect 1974 736 1980 737
rect 1974 732 1975 736
rect 1979 732 1980 736
rect 1974 731 1980 732
rect 2070 736 2076 737
rect 2070 732 2071 736
rect 2075 732 2076 736
rect 2070 731 2076 732
rect 2182 736 2188 737
rect 2182 732 2183 736
rect 2187 732 2188 736
rect 2182 731 2188 732
rect 1870 728 1876 729
rect 2050 727 2056 728
rect 1970 723 1976 724
rect 1970 719 1971 723
rect 1975 719 1976 723
rect 2050 723 2051 727
rect 2055 723 2056 727
rect 2050 722 2056 723
rect 2138 727 2144 728
rect 2138 723 2139 727
rect 2143 723 2144 727
rect 2138 722 2144 723
rect 1970 718 1976 719
rect 1870 716 1876 717
rect 1870 712 1871 716
rect 1875 712 1876 716
rect 1870 711 1876 712
rect 1247 698 1251 699
rect 1247 693 1251 694
rect 1255 698 1259 699
rect 1255 693 1259 694
rect 1351 698 1355 699
rect 1351 693 1355 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1455 698 1459 699
rect 1455 693 1459 694
rect 1519 698 1523 699
rect 1519 693 1523 694
rect 1559 698 1563 699
rect 1559 693 1563 694
rect 1647 698 1651 699
rect 1647 693 1651 694
rect 1663 698 1667 699
rect 1663 693 1667 694
rect 1751 698 1755 699
rect 1751 693 1755 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 1199 684 1203 685
rect 1248 683 1250 693
rect 1298 691 1304 692
rect 1298 687 1299 691
rect 1303 687 1304 691
rect 1298 686 1304 687
rect 1199 679 1203 680
rect 1246 682 1252 683
rect 1246 678 1247 682
rect 1251 678 1252 682
rect 1246 677 1252 678
rect 1300 656 1302 686
rect 1352 683 1354 693
rect 1402 691 1408 692
rect 1402 687 1403 691
rect 1407 687 1408 691
rect 1402 686 1408 687
rect 1350 682 1356 683
rect 1350 678 1351 682
rect 1355 678 1356 682
rect 1350 677 1356 678
rect 1404 656 1406 686
rect 1456 683 1458 693
rect 1506 691 1512 692
rect 1506 687 1507 691
rect 1511 687 1512 691
rect 1506 686 1512 687
rect 1454 682 1460 683
rect 1454 678 1455 682
rect 1459 678 1460 682
rect 1454 677 1460 678
rect 1508 656 1510 686
rect 1560 683 1562 693
rect 1567 684 1571 685
rect 1558 682 1564 683
rect 1558 678 1559 682
rect 1563 678 1564 682
rect 1664 683 1666 693
rect 1706 691 1712 692
rect 1706 687 1707 691
rect 1711 687 1712 691
rect 1706 686 1712 687
rect 1714 691 1720 692
rect 1714 687 1715 691
rect 1719 687 1720 691
rect 1714 686 1720 687
rect 1567 679 1571 680
rect 1662 682 1668 683
rect 1558 677 1564 678
rect 1568 656 1570 679
rect 1662 678 1663 682
rect 1667 678 1668 682
rect 1662 677 1668 678
rect 1708 661 1710 686
rect 1707 660 1711 661
rect 1716 656 1718 686
rect 1752 683 1754 693
rect 1750 682 1756 683
rect 1750 678 1751 682
rect 1755 678 1756 682
rect 1750 677 1756 678
rect 1832 665 1834 693
rect 1872 679 1874 711
rect 1902 698 1908 699
rect 1902 694 1903 698
rect 1907 694 1908 698
rect 1902 693 1908 694
rect 1904 679 1906 693
rect 1972 688 1974 718
rect 1982 698 1988 699
rect 1982 694 1983 698
rect 1987 694 1988 698
rect 1982 693 1988 694
rect 1970 687 1976 688
rect 1970 683 1971 687
rect 1975 683 1976 687
rect 1970 682 1976 683
rect 1984 679 1986 693
rect 2052 688 2054 722
rect 2130 719 2136 720
rect 2130 715 2131 719
rect 2135 715 2136 719
rect 2130 714 2136 715
rect 2078 698 2084 699
rect 2078 694 2079 698
rect 2083 694 2084 698
rect 2078 693 2084 694
rect 2050 687 2056 688
rect 2050 683 2051 687
rect 2055 683 2056 687
rect 2050 682 2056 683
rect 2080 679 2082 693
rect 1871 678 1875 679
rect 1871 673 1875 674
rect 1903 678 1907 679
rect 1903 673 1907 674
rect 1983 678 1987 679
rect 1983 673 1987 674
rect 2079 678 2083 679
rect 2079 673 2083 674
rect 2095 678 2099 679
rect 2095 673 2099 674
rect 1830 664 1836 665
rect 1830 660 1831 664
rect 1835 660 1836 664
rect 1830 659 1836 660
rect 1074 655 1080 656
rect 1074 651 1075 655
rect 1079 651 1080 655
rect 1074 650 1080 651
rect 1186 655 1192 656
rect 1186 651 1187 655
rect 1191 651 1192 655
rect 1186 650 1192 651
rect 1298 655 1304 656
rect 1298 651 1299 655
rect 1303 651 1304 655
rect 1298 650 1304 651
rect 1402 655 1408 656
rect 1402 651 1403 655
rect 1407 651 1408 655
rect 1402 650 1408 651
rect 1506 655 1512 656
rect 1506 651 1507 655
rect 1511 651 1512 655
rect 1506 650 1512 651
rect 1566 655 1572 656
rect 1707 655 1711 656
rect 1714 655 1720 656
rect 1566 651 1567 655
rect 1571 651 1572 655
rect 1566 650 1572 651
rect 1714 651 1715 655
rect 1719 651 1720 655
rect 1714 650 1720 651
rect 1830 647 1836 648
rect 1126 644 1132 645
rect 1126 640 1127 644
rect 1131 640 1132 644
rect 1126 639 1132 640
rect 1238 644 1244 645
rect 1238 640 1239 644
rect 1243 640 1244 644
rect 1238 639 1244 640
rect 1342 644 1348 645
rect 1342 640 1343 644
rect 1347 640 1348 644
rect 1342 639 1348 640
rect 1446 644 1452 645
rect 1446 640 1447 644
rect 1451 640 1452 644
rect 1446 639 1452 640
rect 1550 644 1556 645
rect 1550 640 1551 644
rect 1555 640 1556 644
rect 1550 639 1556 640
rect 1654 644 1660 645
rect 1654 640 1655 644
rect 1659 640 1660 644
rect 1654 639 1660 640
rect 1742 644 1748 645
rect 1742 640 1743 644
rect 1747 640 1748 644
rect 1830 643 1831 647
rect 1835 643 1836 647
rect 1872 645 1874 673
rect 1904 663 1906 673
rect 2096 663 2098 673
rect 2132 672 2134 714
rect 2140 680 2142 722
rect 2262 719 2268 720
rect 2262 715 2263 719
rect 2267 715 2268 719
rect 2262 714 2268 715
rect 2190 698 2196 699
rect 2190 694 2191 698
rect 2195 694 2196 698
rect 2190 693 2196 694
rect 2138 679 2144 680
rect 2192 679 2194 693
rect 2264 688 2266 714
rect 2300 688 2302 794
rect 2318 788 2324 789
rect 2318 784 2319 788
rect 2323 784 2324 788
rect 2318 783 2324 784
rect 2414 788 2420 789
rect 2414 784 2415 788
rect 2419 784 2420 788
rect 2414 783 2420 784
rect 2526 788 2532 789
rect 2526 784 2527 788
rect 2531 784 2532 788
rect 2526 783 2532 784
rect 2646 788 2652 789
rect 2646 784 2647 788
rect 2651 784 2652 788
rect 2646 783 2652 784
rect 2774 788 2780 789
rect 2774 784 2775 788
rect 2779 784 2780 788
rect 2774 783 2780 784
rect 2320 759 2322 783
rect 2416 759 2418 783
rect 2528 759 2530 783
rect 2648 759 2650 783
rect 2776 759 2778 783
rect 2311 758 2315 759
rect 2311 753 2315 754
rect 2319 758 2323 759
rect 2319 753 2323 754
rect 2415 758 2419 759
rect 2415 753 2419 754
rect 2447 758 2451 759
rect 2447 753 2451 754
rect 2527 758 2531 759
rect 2527 753 2531 754
rect 2591 758 2595 759
rect 2591 753 2595 754
rect 2647 758 2651 759
rect 2647 753 2651 754
rect 2743 758 2747 759
rect 2743 753 2747 754
rect 2775 758 2779 759
rect 2775 753 2779 754
rect 2312 737 2314 753
rect 2448 737 2450 753
rect 2592 737 2594 753
rect 2744 737 2746 753
rect 2310 736 2316 737
rect 2310 732 2311 736
rect 2315 732 2316 736
rect 2310 731 2316 732
rect 2446 736 2452 737
rect 2446 732 2447 736
rect 2451 732 2452 736
rect 2446 731 2452 732
rect 2590 736 2596 737
rect 2590 732 2591 736
rect 2595 732 2596 736
rect 2590 731 2596 732
rect 2742 736 2748 737
rect 2742 732 2743 736
rect 2747 732 2748 736
rect 2742 731 2748 732
rect 2402 727 2408 728
rect 2402 723 2403 727
rect 2407 723 2408 727
rect 2402 722 2408 723
rect 2514 727 2520 728
rect 2514 723 2515 727
rect 2519 723 2520 727
rect 2514 722 2520 723
rect 2658 727 2664 728
rect 2658 723 2659 727
rect 2663 723 2664 727
rect 2658 722 2664 723
rect 2810 727 2816 728
rect 2810 723 2811 727
rect 2815 723 2816 727
rect 2810 722 2816 723
rect 2318 698 2324 699
rect 2318 694 2319 698
rect 2323 694 2324 698
rect 2318 693 2324 694
rect 2262 687 2268 688
rect 2262 683 2263 687
rect 2267 683 2268 687
rect 2262 682 2268 683
rect 2298 687 2304 688
rect 2298 683 2299 687
rect 2303 683 2304 687
rect 2298 682 2304 683
rect 2320 679 2322 693
rect 2404 688 2406 722
rect 2454 698 2460 699
rect 2454 694 2455 698
rect 2459 694 2460 698
rect 2454 693 2460 694
rect 2402 687 2408 688
rect 2402 683 2403 687
rect 2407 683 2408 687
rect 2402 682 2408 683
rect 2456 679 2458 693
rect 2138 675 2139 679
rect 2143 675 2144 679
rect 2138 674 2144 675
rect 2191 678 2195 679
rect 2191 673 2195 674
rect 2295 678 2299 679
rect 2295 673 2299 674
rect 2319 678 2323 679
rect 2319 673 2323 674
rect 2455 678 2459 679
rect 2455 673 2459 674
rect 2479 678 2483 679
rect 2479 673 2483 674
rect 2130 671 2136 672
rect 2130 667 2131 671
rect 2135 667 2136 671
rect 2130 666 2136 667
rect 2146 671 2152 672
rect 2146 667 2147 671
rect 2151 667 2152 671
rect 2146 666 2152 667
rect 1902 662 1908 663
rect 1902 658 1903 662
rect 1907 658 1908 662
rect 1902 657 1908 658
rect 2094 662 2100 663
rect 2094 658 2095 662
rect 2099 658 2100 662
rect 2094 657 2100 658
rect 1830 642 1836 643
rect 1870 644 1876 645
rect 1742 639 1748 640
rect 1128 619 1130 639
rect 1240 619 1242 639
rect 1344 619 1346 639
rect 1448 619 1450 639
rect 1552 619 1554 639
rect 1656 619 1658 639
rect 1744 619 1746 639
rect 1832 619 1834 642
rect 1870 640 1871 644
rect 1875 640 1876 644
rect 1870 639 1876 640
rect 2148 636 2150 666
rect 2296 663 2298 673
rect 2480 663 2482 673
rect 2516 672 2518 722
rect 2598 698 2604 699
rect 2598 694 2599 698
rect 2603 694 2604 698
rect 2598 693 2604 694
rect 2600 679 2602 693
rect 2660 688 2662 722
rect 2750 698 2756 699
rect 2750 694 2751 698
rect 2755 694 2756 698
rect 2750 693 2756 694
rect 2658 687 2664 688
rect 2658 683 2659 687
rect 2663 683 2664 687
rect 2658 682 2664 683
rect 2752 679 2754 693
rect 2812 688 2814 722
rect 2836 688 2838 794
rect 2902 788 2908 789
rect 2902 784 2903 788
rect 2907 784 2908 788
rect 2902 783 2908 784
rect 3030 788 3036 789
rect 3030 784 3031 788
rect 3035 784 3036 788
rect 3030 783 3036 784
rect 2904 759 2906 783
rect 3032 759 3034 783
rect 2895 758 2899 759
rect 2895 753 2899 754
rect 2903 758 2907 759
rect 2903 753 2907 754
rect 3031 758 3035 759
rect 3031 753 3035 754
rect 3047 758 3051 759
rect 3047 753 3051 754
rect 2896 737 2898 753
rect 3048 737 3050 753
rect 2894 736 2900 737
rect 2894 732 2895 736
rect 2899 732 2900 736
rect 2894 731 2900 732
rect 3046 736 3052 737
rect 3046 732 3047 736
rect 3051 732 3052 736
rect 3046 731 3052 732
rect 3056 724 3058 830
rect 3092 800 3094 830
rect 3160 827 3162 837
rect 3210 835 3216 836
rect 3210 831 3211 835
rect 3215 831 3216 835
rect 3210 830 3216 831
rect 3158 826 3164 827
rect 3158 822 3159 826
rect 3163 822 3164 826
rect 3158 821 3164 822
rect 3212 800 3214 830
rect 3280 827 3282 837
rect 3394 835 3400 836
rect 3394 831 3395 835
rect 3399 831 3400 835
rect 3394 830 3400 831
rect 3278 826 3284 827
rect 3278 822 3279 826
rect 3283 822 3284 826
rect 3278 821 3284 822
rect 3396 800 3398 830
rect 3408 827 3410 837
rect 3406 826 3412 827
rect 3406 822 3407 826
rect 3411 822 3412 826
rect 3406 821 3412 822
rect 3416 800 3418 854
rect 3432 843 3434 865
rect 3431 842 3435 843
rect 3431 837 3435 838
rect 3484 836 3486 886
rect 3492 860 3494 894
rect 3510 870 3516 871
rect 3510 866 3511 870
rect 3515 866 3516 870
rect 3510 865 3516 866
rect 3490 859 3496 860
rect 3490 855 3491 859
rect 3495 855 3496 859
rect 3490 854 3496 855
rect 3512 843 3514 865
rect 3536 860 3538 966
rect 3590 963 3596 964
rect 3590 959 3591 963
rect 3595 959 3596 963
rect 3590 958 3596 959
rect 3592 931 3594 958
rect 3591 930 3595 931
rect 3591 925 3595 926
rect 3592 906 3594 925
rect 3590 905 3596 906
rect 3590 901 3591 905
rect 3595 901 3596 905
rect 3590 900 3596 901
rect 3590 888 3596 889
rect 3590 884 3591 888
rect 3595 884 3596 888
rect 3590 883 3596 884
rect 3534 859 3540 860
rect 3534 855 3535 859
rect 3539 855 3540 859
rect 3534 854 3540 855
rect 3592 843 3594 883
rect 3511 842 3515 843
rect 3511 837 3515 838
rect 3591 842 3595 843
rect 3591 837 3595 838
rect 3482 835 3488 836
rect 3482 831 3483 835
rect 3487 831 3488 835
rect 3482 830 3488 831
rect 3512 827 3514 837
rect 3510 826 3516 827
rect 3510 822 3511 826
rect 3515 822 3516 826
rect 3510 821 3516 822
rect 3592 809 3594 837
rect 3590 808 3596 809
rect 3590 804 3591 808
rect 3595 804 3596 808
rect 3590 803 3596 804
rect 3090 799 3096 800
rect 3090 795 3091 799
rect 3095 795 3096 799
rect 3090 794 3096 795
rect 3210 799 3216 800
rect 3210 795 3211 799
rect 3215 795 3216 799
rect 3210 794 3216 795
rect 3394 799 3400 800
rect 3394 795 3395 799
rect 3399 795 3400 799
rect 3394 794 3400 795
rect 3414 799 3420 800
rect 3414 795 3415 799
rect 3419 795 3420 799
rect 3414 794 3420 795
rect 3534 799 3540 800
rect 3534 795 3535 799
rect 3539 795 3540 799
rect 3534 794 3540 795
rect 3150 788 3156 789
rect 3150 784 3151 788
rect 3155 784 3156 788
rect 3150 783 3156 784
rect 3270 788 3276 789
rect 3270 784 3271 788
rect 3275 784 3276 788
rect 3270 783 3276 784
rect 3398 788 3404 789
rect 3398 784 3399 788
rect 3403 784 3404 788
rect 3398 783 3404 784
rect 3502 788 3508 789
rect 3502 784 3503 788
rect 3507 784 3508 788
rect 3502 783 3508 784
rect 3152 759 3154 783
rect 3272 759 3274 783
rect 3400 759 3402 783
rect 3504 759 3506 783
rect 3151 758 3155 759
rect 3151 753 3155 754
rect 3199 758 3203 759
rect 3199 753 3203 754
rect 3271 758 3275 759
rect 3271 753 3275 754
rect 3359 758 3363 759
rect 3359 753 3363 754
rect 3399 758 3403 759
rect 3399 753 3403 754
rect 3503 758 3507 759
rect 3503 753 3507 754
rect 3200 737 3202 753
rect 3360 737 3362 753
rect 3504 737 3506 753
rect 3198 736 3204 737
rect 3198 732 3199 736
rect 3203 732 3204 736
rect 3198 731 3204 732
rect 3358 736 3364 737
rect 3358 732 3359 736
rect 3363 732 3364 736
rect 3358 731 3364 732
rect 3502 736 3508 737
rect 3502 732 3503 736
rect 3507 732 3508 736
rect 3502 731 3508 732
rect 3114 727 3120 728
rect 3054 723 3060 724
rect 3054 719 3055 723
rect 3059 719 3060 723
rect 3114 723 3115 727
rect 3119 723 3120 727
rect 3114 722 3120 723
rect 3266 727 3272 728
rect 3266 723 3267 727
rect 3271 723 3272 727
rect 3266 722 3272 723
rect 3054 718 3060 719
rect 2902 698 2908 699
rect 2902 694 2903 698
rect 2907 694 2908 698
rect 2902 693 2908 694
rect 3054 698 3060 699
rect 3054 694 3055 698
rect 3059 694 3060 698
rect 3054 693 3060 694
rect 2810 687 2816 688
rect 2810 683 2811 687
rect 2815 683 2816 687
rect 2810 682 2816 683
rect 2834 687 2840 688
rect 2834 683 2835 687
rect 2839 683 2840 687
rect 2834 682 2840 683
rect 2904 679 2906 693
rect 3056 679 3058 693
rect 3116 688 3118 722
rect 3206 698 3212 699
rect 3206 694 3207 698
rect 3211 694 3212 698
rect 3206 693 3212 694
rect 3114 687 3120 688
rect 3114 683 3115 687
rect 3119 683 3120 687
rect 3114 682 3120 683
rect 3208 679 3210 693
rect 3268 688 3270 722
rect 3366 698 3372 699
rect 3366 694 3367 698
rect 3371 694 3372 698
rect 3366 693 3372 694
rect 3510 698 3516 699
rect 3510 694 3511 698
rect 3515 694 3516 698
rect 3510 693 3516 694
rect 3266 687 3272 688
rect 3266 683 3267 687
rect 3271 683 3272 687
rect 3266 682 3272 683
rect 3368 679 3370 693
rect 3390 687 3396 688
rect 3390 683 3391 687
rect 3395 683 3396 687
rect 3390 682 3396 683
rect 2599 678 2603 679
rect 2599 673 2603 674
rect 2655 678 2659 679
rect 2655 673 2659 674
rect 2751 678 2755 679
rect 2751 673 2755 674
rect 2831 678 2835 679
rect 2831 673 2835 674
rect 2903 678 2907 679
rect 2903 673 2907 674
rect 3007 678 3011 679
rect 3007 673 3011 674
rect 3055 678 3059 679
rect 3055 673 3059 674
rect 3183 678 3187 679
rect 3183 673 3187 674
rect 3207 678 3211 679
rect 3207 673 3211 674
rect 3359 678 3363 679
rect 3359 673 3363 674
rect 3367 678 3371 679
rect 3367 673 3371 674
rect 2514 671 2520 672
rect 2514 667 2515 671
rect 2519 667 2520 671
rect 2514 666 2520 667
rect 2530 671 2536 672
rect 2530 667 2531 671
rect 2535 667 2536 671
rect 2530 666 2536 667
rect 2294 662 2300 663
rect 2294 658 2295 662
rect 2299 658 2300 662
rect 2478 662 2484 663
rect 2294 657 2300 658
rect 2303 660 2307 661
rect 2478 658 2479 662
rect 2483 658 2484 662
rect 2478 657 2484 658
rect 2303 655 2307 656
rect 2304 636 2306 655
rect 2532 636 2534 666
rect 2656 663 2658 673
rect 2832 663 2834 673
rect 2874 671 2880 672
rect 2874 667 2875 671
rect 2879 667 2880 671
rect 2874 666 2880 667
rect 2882 671 2888 672
rect 2882 667 2883 671
rect 2887 667 2888 671
rect 2882 666 2888 667
rect 2654 662 2660 663
rect 2654 658 2655 662
rect 2659 658 2660 662
rect 2654 657 2660 658
rect 2830 662 2836 663
rect 2830 658 2831 662
rect 2835 658 2836 662
rect 2830 657 2836 658
rect 1926 635 1932 636
rect 1926 631 1927 635
rect 1931 631 1932 635
rect 1926 630 1932 631
rect 2146 635 2152 636
rect 2146 631 2147 635
rect 2151 631 2152 635
rect 2146 630 2152 631
rect 2302 635 2308 636
rect 2302 631 2303 635
rect 2307 631 2308 635
rect 2302 630 2308 631
rect 2530 635 2536 636
rect 2530 631 2531 635
rect 2535 631 2536 635
rect 2530 630 2536 631
rect 2678 635 2684 636
rect 2678 631 2679 635
rect 2683 631 2684 635
rect 2678 630 2684 631
rect 1870 627 1876 628
rect 1870 623 1871 627
rect 1875 623 1876 627
rect 1870 622 1876 623
rect 1894 624 1900 625
rect 1087 618 1091 619
rect 1087 613 1091 614
rect 1127 618 1131 619
rect 1127 613 1131 614
rect 1175 618 1179 619
rect 1175 613 1179 614
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 1263 618 1267 619
rect 1263 613 1267 614
rect 1343 618 1347 619
rect 1343 613 1347 614
rect 1447 618 1451 619
rect 1447 613 1451 614
rect 1551 618 1555 619
rect 1551 613 1555 614
rect 1655 618 1659 619
rect 1655 613 1659 614
rect 1743 618 1747 619
rect 1743 613 1747 614
rect 1831 618 1835 619
rect 1831 613 1835 614
rect 1088 597 1090 613
rect 1176 597 1178 613
rect 1264 597 1266 613
rect 1086 596 1092 597
rect 1086 592 1087 596
rect 1091 592 1092 596
rect 1086 591 1092 592
rect 1174 596 1180 597
rect 1174 592 1175 596
rect 1179 592 1180 596
rect 1174 591 1180 592
rect 1262 596 1268 597
rect 1262 592 1263 596
rect 1267 592 1268 596
rect 1832 594 1834 613
rect 1872 599 1874 622
rect 1894 620 1895 624
rect 1899 620 1900 624
rect 1894 619 1900 620
rect 1896 599 1898 619
rect 1871 598 1875 599
rect 1262 591 1268 592
rect 1830 593 1836 594
rect 1871 593 1875 594
rect 1895 598 1899 599
rect 1895 593 1899 594
rect 1830 589 1831 593
rect 1835 589 1836 593
rect 1830 588 1836 589
rect 1066 587 1072 588
rect 1066 583 1067 587
rect 1071 583 1072 587
rect 1066 582 1072 583
rect 1154 587 1160 588
rect 1154 583 1155 587
rect 1159 583 1160 587
rect 1154 582 1160 583
rect 1242 587 1248 588
rect 1242 583 1243 587
rect 1247 583 1248 587
rect 1242 582 1248 583
rect 1058 579 1064 580
rect 1058 575 1059 579
rect 1063 575 1064 579
rect 1058 574 1064 575
rect 1006 558 1012 559
rect 1006 554 1007 558
rect 1011 554 1012 558
rect 1006 553 1012 554
rect 978 547 984 548
rect 978 543 979 547
rect 983 543 984 547
rect 978 542 984 543
rect 1008 531 1010 553
rect 1068 548 1070 582
rect 1094 558 1100 559
rect 1094 554 1095 558
rect 1099 554 1100 558
rect 1094 553 1100 554
rect 1066 547 1072 548
rect 1066 543 1067 547
rect 1071 543 1072 547
rect 1066 542 1072 543
rect 1096 531 1098 553
rect 1156 548 1158 582
rect 1182 558 1188 559
rect 1182 554 1183 558
rect 1187 554 1188 558
rect 1182 553 1188 554
rect 1154 547 1160 548
rect 1154 543 1155 547
rect 1159 543 1160 547
rect 1154 542 1160 543
rect 1184 531 1186 553
rect 1244 548 1246 582
rect 1830 576 1836 577
rect 1830 572 1831 576
rect 1835 572 1836 576
rect 1872 574 1874 593
rect 1896 577 1898 593
rect 1894 576 1900 577
rect 1830 571 1836 572
rect 1870 573 1876 574
rect 1270 558 1276 559
rect 1270 554 1271 558
rect 1275 554 1276 558
rect 1270 553 1276 554
rect 1242 547 1248 548
rect 1242 543 1243 547
rect 1247 543 1248 547
rect 1242 542 1248 543
rect 1272 531 1274 553
rect 1832 531 1834 571
rect 1870 569 1871 573
rect 1875 569 1876 573
rect 1894 572 1895 576
rect 1899 572 1900 576
rect 1894 571 1900 572
rect 1870 568 1876 569
rect 1870 556 1876 557
rect 1870 552 1871 556
rect 1875 552 1876 556
rect 1870 551 1876 552
rect 895 530 899 531
rect 895 525 899 526
rect 919 530 923 531
rect 919 525 923 526
rect 983 530 987 531
rect 983 525 987 526
rect 1007 530 1011 531
rect 1007 525 1011 526
rect 1071 530 1075 531
rect 1071 525 1075 526
rect 1095 530 1099 531
rect 1095 525 1099 526
rect 1159 530 1163 531
rect 1159 525 1163 526
rect 1183 530 1187 531
rect 1183 525 1187 526
rect 1247 530 1251 531
rect 1247 525 1251 526
rect 1271 530 1275 531
rect 1271 525 1275 526
rect 1831 530 1835 531
rect 1831 525 1835 526
rect 883 516 887 517
rect 896 515 898 525
rect 946 523 952 524
rect 946 519 947 523
rect 951 519 952 523
rect 946 518 952 519
rect 883 511 887 512
rect 894 514 900 515
rect 894 510 895 514
rect 899 510 900 514
rect 894 509 900 510
rect 948 488 950 518
rect 984 515 986 525
rect 1034 523 1040 524
rect 1034 519 1035 523
rect 1039 519 1040 523
rect 1034 518 1040 519
rect 982 514 988 515
rect 982 510 983 514
rect 987 510 988 514
rect 982 509 988 510
rect 1036 488 1038 518
rect 1072 515 1074 525
rect 1122 523 1128 524
rect 1122 519 1123 523
rect 1127 519 1128 523
rect 1122 518 1128 519
rect 1070 514 1076 515
rect 1070 510 1071 514
rect 1075 510 1076 514
rect 1070 509 1076 510
rect 1124 488 1126 518
rect 1160 515 1162 525
rect 1210 523 1216 524
rect 1210 519 1211 523
rect 1215 519 1216 523
rect 1210 518 1216 519
rect 1158 514 1164 515
rect 1158 510 1159 514
rect 1163 510 1164 514
rect 1158 509 1164 510
rect 1212 488 1214 518
rect 1248 515 1250 525
rect 1255 516 1259 517
rect 1246 514 1252 515
rect 1246 510 1247 514
rect 1251 510 1252 514
rect 1255 511 1259 512
rect 1246 509 1252 510
rect 1256 488 1258 511
rect 1832 497 1834 525
rect 1872 523 1874 551
rect 1902 538 1908 539
rect 1902 534 1903 538
rect 1907 534 1908 538
rect 1902 533 1908 534
rect 1904 523 1906 533
rect 1928 528 1930 630
rect 2086 624 2092 625
rect 2086 620 2087 624
rect 2091 620 2092 624
rect 2086 619 2092 620
rect 2286 624 2292 625
rect 2286 620 2287 624
rect 2291 620 2292 624
rect 2286 619 2292 620
rect 2470 624 2476 625
rect 2470 620 2471 624
rect 2475 620 2476 624
rect 2470 619 2476 620
rect 2646 624 2652 625
rect 2646 620 2647 624
rect 2651 620 2652 624
rect 2646 619 2652 620
rect 2088 599 2090 619
rect 2288 599 2290 619
rect 2472 599 2474 619
rect 2648 599 2650 619
rect 1975 598 1979 599
rect 1975 593 1979 594
rect 2087 598 2091 599
rect 2087 593 2091 594
rect 2215 598 2219 599
rect 2215 593 2219 594
rect 2287 598 2291 599
rect 2287 593 2291 594
rect 2351 598 2355 599
rect 2351 593 2355 594
rect 2471 598 2475 599
rect 2471 593 2475 594
rect 2495 598 2499 599
rect 2495 593 2499 594
rect 2647 598 2651 599
rect 2647 593 2651 594
rect 1976 577 1978 593
rect 2088 577 2090 593
rect 2216 577 2218 593
rect 2352 577 2354 593
rect 2496 577 2498 593
rect 2648 577 2650 593
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2086 576 2092 577
rect 2086 572 2087 576
rect 2091 572 2092 576
rect 2086 571 2092 572
rect 2214 576 2220 577
rect 2214 572 2215 576
rect 2219 572 2220 576
rect 2214 571 2220 572
rect 2350 576 2356 577
rect 2350 572 2351 576
rect 2355 572 2356 576
rect 2350 571 2356 572
rect 2494 576 2500 577
rect 2494 572 2495 576
rect 2499 572 2500 576
rect 2494 571 2500 572
rect 2646 576 2652 577
rect 2646 572 2647 576
rect 2651 572 2652 576
rect 2646 571 2652 572
rect 1962 567 1968 568
rect 1962 563 1963 567
rect 1967 563 1968 567
rect 1962 562 1968 563
rect 2058 567 2064 568
rect 2058 563 2059 567
rect 2063 563 2064 567
rect 2058 562 2064 563
rect 2162 567 2168 568
rect 2162 563 2163 567
rect 2167 563 2168 567
rect 2162 562 2168 563
rect 2298 567 2304 568
rect 2298 563 2299 567
rect 2303 563 2304 567
rect 2298 562 2304 563
rect 2442 567 2448 568
rect 2442 563 2443 567
rect 2447 563 2448 567
rect 2442 562 2448 563
rect 2450 567 2456 568
rect 2450 563 2451 567
rect 2455 563 2456 567
rect 2450 562 2456 563
rect 1964 528 1966 562
rect 1982 538 1988 539
rect 1982 534 1983 538
rect 1987 534 1988 538
rect 1982 533 1988 534
rect 1926 527 1932 528
rect 1926 523 1927 527
rect 1931 523 1932 527
rect 1871 522 1875 523
rect 1871 517 1875 518
rect 1903 522 1907 523
rect 1926 522 1932 523
rect 1962 527 1968 528
rect 1962 523 1963 527
rect 1967 523 1968 527
rect 1984 523 1986 533
rect 2060 528 2062 562
rect 2094 538 2100 539
rect 2094 534 2095 538
rect 2099 534 2100 538
rect 2094 533 2100 534
rect 2058 527 2064 528
rect 2058 523 2059 527
rect 2063 523 2064 527
rect 2096 523 2098 533
rect 2164 528 2166 562
rect 2179 540 2183 541
rect 2179 535 2183 536
rect 2222 538 2228 539
rect 2162 527 2168 528
rect 2162 523 2163 527
rect 2167 523 2168 527
rect 1962 522 1968 523
rect 1983 522 1987 523
rect 2058 522 2064 523
rect 2095 522 2099 523
rect 1903 517 1907 518
rect 1983 517 1987 518
rect 2095 517 2099 518
rect 2151 522 2155 523
rect 2162 522 2168 523
rect 2151 517 2155 518
rect 1830 496 1836 497
rect 1830 492 1831 496
rect 1835 492 1836 496
rect 1830 491 1836 492
rect 1872 489 1874 517
rect 2152 507 2154 517
rect 2180 516 2182 535
rect 2222 534 2223 538
rect 2227 534 2228 538
rect 2222 533 2228 534
rect 2224 523 2226 533
rect 2300 528 2302 562
rect 2358 538 2364 539
rect 2358 534 2359 538
rect 2363 534 2364 538
rect 2358 533 2364 534
rect 2298 527 2304 528
rect 2298 523 2299 527
rect 2303 523 2304 527
rect 2360 523 2362 533
rect 2444 528 2446 562
rect 2452 541 2454 562
rect 2451 540 2455 541
rect 2451 535 2455 536
rect 2502 538 2508 539
rect 2502 534 2503 538
rect 2507 534 2508 538
rect 2502 533 2508 534
rect 2654 538 2660 539
rect 2654 534 2655 538
rect 2659 534 2660 538
rect 2654 533 2660 534
rect 2442 527 2448 528
rect 2442 523 2443 527
rect 2447 523 2448 527
rect 2504 523 2506 533
rect 2656 523 2658 533
rect 2680 528 2682 630
rect 2822 624 2828 625
rect 2822 620 2823 624
rect 2827 620 2828 624
rect 2822 619 2828 620
rect 2824 599 2826 619
rect 2807 598 2811 599
rect 2807 593 2811 594
rect 2823 598 2827 599
rect 2823 593 2827 594
rect 2808 577 2810 593
rect 2806 576 2812 577
rect 2806 572 2807 576
rect 2811 572 2812 576
rect 2806 571 2812 572
rect 2876 568 2878 666
rect 2884 636 2886 666
rect 3008 663 3010 673
rect 3174 671 3180 672
rect 3174 667 3175 671
rect 3179 667 3180 671
rect 3174 666 3180 667
rect 3006 662 3012 663
rect 3006 658 3007 662
rect 3011 658 3012 662
rect 3006 657 3012 658
rect 3176 636 3178 666
rect 3184 663 3186 673
rect 3234 671 3240 672
rect 3234 667 3235 671
rect 3239 667 3240 671
rect 3234 666 3240 667
rect 3182 662 3188 663
rect 3182 658 3183 662
rect 3187 658 3188 662
rect 3182 657 3188 658
rect 3236 636 3238 666
rect 3360 663 3362 673
rect 3358 662 3364 663
rect 3358 658 3359 662
rect 3363 658 3364 662
rect 3358 657 3364 658
rect 3392 636 3394 682
rect 3512 679 3514 693
rect 3536 688 3538 794
rect 3590 791 3596 792
rect 3590 787 3591 791
rect 3595 787 3596 791
rect 3590 786 3596 787
rect 3592 759 3594 786
rect 3591 758 3595 759
rect 3591 753 3595 754
rect 3592 734 3594 753
rect 3590 733 3596 734
rect 3590 729 3591 733
rect 3595 729 3596 733
rect 3590 728 3596 729
rect 3562 719 3568 720
rect 3562 715 3563 719
rect 3567 715 3568 719
rect 3562 714 3568 715
rect 3590 716 3596 717
rect 3534 687 3540 688
rect 3534 683 3535 687
rect 3539 683 3540 687
rect 3534 682 3540 683
rect 3511 678 3515 679
rect 3511 673 3515 674
rect 3512 663 3514 673
rect 3564 672 3566 714
rect 3590 712 3591 716
rect 3595 712 3596 716
rect 3590 711 3596 712
rect 3592 679 3594 711
rect 3591 678 3595 679
rect 3591 673 3595 674
rect 3562 671 3568 672
rect 3562 667 3563 671
rect 3567 667 3568 671
rect 3562 666 3568 667
rect 3510 662 3516 663
rect 3510 658 3511 662
rect 3515 658 3516 662
rect 3510 657 3516 658
rect 3592 645 3594 673
rect 3590 644 3596 645
rect 3590 640 3591 644
rect 3595 640 3596 644
rect 3590 639 3596 640
rect 2882 635 2888 636
rect 2882 631 2883 635
rect 2887 631 2888 635
rect 2882 630 2888 631
rect 3174 635 3180 636
rect 3174 631 3175 635
rect 3179 631 3180 635
rect 3174 630 3180 631
rect 3234 635 3240 636
rect 3234 631 3235 635
rect 3239 631 3240 635
rect 3234 630 3240 631
rect 3390 635 3396 636
rect 3390 631 3391 635
rect 3395 631 3396 635
rect 3390 630 3396 631
rect 3534 635 3540 636
rect 3534 631 3535 635
rect 3539 631 3540 635
rect 3534 630 3540 631
rect 2998 624 3004 625
rect 2998 620 2999 624
rect 3003 620 3004 624
rect 2998 619 3004 620
rect 3174 624 3180 625
rect 3174 620 3175 624
rect 3179 620 3180 624
rect 3174 619 3180 620
rect 3350 624 3356 625
rect 3350 620 3351 624
rect 3355 620 3356 624
rect 3350 619 3356 620
rect 3502 624 3508 625
rect 3502 620 3503 624
rect 3507 620 3508 624
rect 3502 619 3508 620
rect 3000 599 3002 619
rect 3176 599 3178 619
rect 3352 599 3354 619
rect 3504 599 3506 619
rect 2975 598 2979 599
rect 2975 593 2979 594
rect 2999 598 3003 599
rect 2999 593 3003 594
rect 3151 598 3155 599
rect 3151 593 3155 594
rect 3175 598 3179 599
rect 3175 593 3179 594
rect 3335 598 3339 599
rect 3335 593 3339 594
rect 3351 598 3355 599
rect 3351 593 3355 594
rect 3503 598 3507 599
rect 3503 593 3507 594
rect 2976 577 2978 593
rect 3152 577 3154 593
rect 3336 577 3338 593
rect 3504 577 3506 593
rect 2974 576 2980 577
rect 2974 572 2975 576
rect 2979 572 2980 576
rect 2974 571 2980 572
rect 3150 576 3156 577
rect 3150 572 3151 576
rect 3155 572 3156 576
rect 3150 571 3156 572
rect 3334 576 3340 577
rect 3334 572 3335 576
rect 3339 572 3340 576
rect 3334 571 3340 572
rect 3502 576 3508 577
rect 3502 572 3503 576
rect 3507 572 3508 576
rect 3502 571 3508 572
rect 2746 567 2752 568
rect 2746 563 2747 567
rect 2751 563 2752 567
rect 2746 562 2752 563
rect 2874 567 2880 568
rect 2874 563 2875 567
rect 2879 563 2880 567
rect 2874 562 2880 563
rect 3042 567 3048 568
rect 3042 563 3043 567
rect 3047 563 3048 567
rect 3042 562 3048 563
rect 3218 567 3224 568
rect 3218 563 3219 567
rect 3223 563 3224 567
rect 3218 562 3224 563
rect 2748 528 2750 562
rect 2866 559 2872 560
rect 2866 555 2867 559
rect 2871 555 2872 559
rect 2866 554 2872 555
rect 2814 538 2820 539
rect 2814 534 2815 538
rect 2819 534 2820 538
rect 2814 533 2820 534
rect 2678 527 2684 528
rect 2678 523 2679 527
rect 2683 523 2684 527
rect 2746 527 2752 528
rect 2746 523 2747 527
rect 2751 523 2752 527
rect 2816 523 2818 533
rect 2223 522 2227 523
rect 2223 517 2227 518
rect 2231 522 2235 523
rect 2298 522 2304 523
rect 2327 522 2331 523
rect 2231 517 2235 518
rect 2327 517 2331 518
rect 2359 522 2363 523
rect 2359 517 2363 518
rect 2431 522 2435 523
rect 2442 522 2448 523
rect 2503 522 2507 523
rect 2431 517 2435 518
rect 2503 517 2507 518
rect 2551 522 2555 523
rect 2551 517 2555 518
rect 2655 522 2659 523
rect 2678 522 2684 523
rect 2687 522 2691 523
rect 2746 522 2752 523
rect 2815 522 2819 523
rect 2655 517 2659 518
rect 2687 517 2691 518
rect 2815 517 2819 518
rect 2839 522 2843 523
rect 2839 517 2843 518
rect 2178 515 2184 516
rect 2178 511 2179 515
rect 2183 511 2184 515
rect 2178 510 2184 511
rect 2202 515 2208 516
rect 2202 511 2203 515
rect 2207 511 2208 515
rect 2202 510 2208 511
rect 2150 506 2156 507
rect 2150 502 2151 506
rect 2155 502 2156 506
rect 2150 501 2156 502
rect 1870 488 1876 489
rect 858 487 864 488
rect 858 483 859 487
rect 863 483 864 487
rect 858 482 864 483
rect 946 487 952 488
rect 946 483 947 487
rect 951 483 952 487
rect 946 482 952 483
rect 1034 487 1040 488
rect 1034 483 1035 487
rect 1039 483 1040 487
rect 1034 482 1040 483
rect 1122 487 1128 488
rect 1122 483 1123 487
rect 1127 483 1128 487
rect 1122 482 1128 483
rect 1210 487 1216 488
rect 1210 483 1211 487
rect 1215 483 1216 487
rect 1210 482 1216 483
rect 1254 487 1260 488
rect 1254 483 1255 487
rect 1259 483 1260 487
rect 1870 484 1871 488
rect 1875 484 1876 488
rect 1870 483 1876 484
rect 1254 482 1260 483
rect 2204 480 2206 510
rect 2232 507 2234 517
rect 2282 515 2288 516
rect 2282 511 2283 515
rect 2287 511 2288 515
rect 2282 510 2288 511
rect 2230 506 2236 507
rect 2230 502 2231 506
rect 2235 502 2236 506
rect 2230 501 2236 502
rect 2284 480 2286 510
rect 2328 507 2330 517
rect 2378 515 2384 516
rect 2378 511 2379 515
rect 2383 511 2384 515
rect 2378 510 2384 511
rect 2326 506 2332 507
rect 2326 502 2327 506
rect 2331 502 2332 506
rect 2326 501 2332 502
rect 2380 480 2382 510
rect 2432 507 2434 517
rect 2482 515 2488 516
rect 2482 511 2483 515
rect 2487 511 2488 515
rect 2482 510 2488 511
rect 2430 506 2436 507
rect 2430 502 2431 506
rect 2435 502 2436 506
rect 2430 501 2436 502
rect 2484 480 2486 510
rect 2552 507 2554 517
rect 2602 515 2608 516
rect 2602 511 2603 515
rect 2607 511 2608 515
rect 2602 510 2608 511
rect 2550 506 2556 507
rect 2550 502 2551 506
rect 2555 502 2556 506
rect 2550 501 2556 502
rect 2604 480 2606 510
rect 2688 507 2690 517
rect 2840 507 2842 517
rect 2868 516 2870 554
rect 2982 538 2988 539
rect 2982 534 2983 538
rect 2987 534 2988 538
rect 2982 533 2988 534
rect 2984 523 2986 533
rect 3044 528 3046 562
rect 3158 538 3164 539
rect 3158 534 3159 538
rect 3163 534 3164 538
rect 3158 533 3164 534
rect 3042 527 3048 528
rect 3042 523 3043 527
rect 3047 523 3048 527
rect 3160 523 3162 533
rect 3220 528 3222 562
rect 3342 538 3348 539
rect 3342 534 3343 538
rect 3347 534 3348 538
rect 3342 533 3348 534
rect 3510 538 3516 539
rect 3510 534 3511 538
rect 3515 534 3516 538
rect 3510 533 3516 534
rect 3218 527 3224 528
rect 3218 523 3219 527
rect 3223 523 3224 527
rect 3344 523 3346 533
rect 3366 527 3372 528
rect 3366 523 3367 527
rect 3371 523 3372 527
rect 3512 523 3514 533
rect 3536 528 3538 630
rect 3590 627 3596 628
rect 3590 623 3591 627
rect 3595 623 3596 627
rect 3590 622 3596 623
rect 3592 599 3594 622
rect 3591 598 3595 599
rect 3591 593 3595 594
rect 3592 574 3594 593
rect 3590 573 3596 574
rect 3590 569 3591 573
rect 3595 569 3596 573
rect 3590 568 3596 569
rect 3562 559 3568 560
rect 3562 555 3563 559
rect 3567 555 3568 559
rect 3562 554 3568 555
rect 3590 556 3596 557
rect 3534 527 3540 528
rect 3534 523 3535 527
rect 3539 523 3540 527
rect 2983 522 2987 523
rect 2983 517 2987 518
rect 2999 522 3003 523
rect 3042 522 3048 523
rect 3159 522 3163 523
rect 2999 517 3003 518
rect 3159 517 3163 518
rect 3175 522 3179 523
rect 3218 522 3224 523
rect 3343 522 3347 523
rect 3175 517 3179 518
rect 3343 517 3347 518
rect 3351 522 3355 523
rect 3366 522 3372 523
rect 3511 522 3515 523
rect 3534 522 3540 523
rect 3351 517 3355 518
rect 2866 515 2872 516
rect 2866 511 2867 515
rect 2871 511 2872 515
rect 2866 510 2872 511
rect 2890 515 2896 516
rect 2890 511 2891 515
rect 2895 511 2896 515
rect 2890 510 2896 511
rect 2686 506 2692 507
rect 2686 502 2687 506
rect 2691 502 2692 506
rect 2686 501 2692 502
rect 2838 506 2844 507
rect 2838 502 2839 506
rect 2843 502 2844 506
rect 2838 501 2844 502
rect 2892 480 2894 510
rect 3000 507 3002 517
rect 3176 507 3178 517
rect 3202 515 3208 516
rect 3202 511 3203 515
rect 3207 511 3208 515
rect 3202 510 3208 511
rect 3226 515 3232 516
rect 3226 511 3227 515
rect 3231 511 3232 515
rect 3226 510 3232 511
rect 2998 506 3004 507
rect 2998 502 2999 506
rect 3003 502 3004 506
rect 2998 501 3004 502
rect 3174 506 3180 507
rect 3174 502 3175 506
rect 3179 502 3180 506
rect 3174 501 3180 502
rect 1830 479 1836 480
rect 798 476 804 477
rect 798 472 799 476
rect 803 472 804 476
rect 798 471 804 472
rect 886 476 892 477
rect 886 472 887 476
rect 891 472 892 476
rect 886 471 892 472
rect 974 476 980 477
rect 974 472 975 476
rect 979 472 980 476
rect 974 471 980 472
rect 1062 476 1068 477
rect 1062 472 1063 476
rect 1067 472 1068 476
rect 1062 471 1068 472
rect 1150 476 1156 477
rect 1150 472 1151 476
rect 1155 472 1156 476
rect 1150 471 1156 472
rect 1238 476 1244 477
rect 1238 472 1239 476
rect 1243 472 1244 476
rect 1830 475 1831 479
rect 1835 475 1836 479
rect 1830 474 1836 475
rect 2202 479 2208 480
rect 2202 475 2203 479
rect 2207 475 2208 479
rect 2202 474 2208 475
rect 2282 479 2288 480
rect 2282 475 2283 479
rect 2287 475 2288 479
rect 2282 474 2288 475
rect 2378 479 2384 480
rect 2378 475 2379 479
rect 2383 475 2384 479
rect 2378 474 2384 475
rect 2482 479 2488 480
rect 2482 475 2483 479
rect 2487 475 2488 479
rect 2482 474 2488 475
rect 2602 479 2608 480
rect 2602 475 2603 479
rect 2607 475 2608 479
rect 2602 474 2608 475
rect 2718 479 2724 480
rect 2718 475 2719 479
rect 2723 475 2724 479
rect 2718 474 2724 475
rect 2890 479 2896 480
rect 2890 475 2891 479
rect 2895 475 2896 479
rect 2890 474 2896 475
rect 3050 479 3056 480
rect 3050 475 3051 479
rect 3055 475 3056 479
rect 3050 474 3056 475
rect 1238 471 1244 472
rect 800 447 802 471
rect 888 447 890 471
rect 976 447 978 471
rect 1064 447 1066 471
rect 1152 447 1154 471
rect 1240 447 1242 471
rect 1832 447 1834 474
rect 1870 471 1876 472
rect 1870 467 1871 471
rect 1875 467 1876 471
rect 1870 466 1876 467
rect 2142 468 2148 469
rect 799 446 803 447
rect 799 441 803 442
rect 823 446 827 447
rect 823 441 827 442
rect 887 446 891 447
rect 887 441 891 442
rect 919 446 923 447
rect 919 441 923 442
rect 975 446 979 447
rect 975 441 979 442
rect 1007 446 1011 447
rect 1007 441 1011 442
rect 1063 446 1067 447
rect 1063 441 1067 442
rect 1103 446 1107 447
rect 1103 441 1107 442
rect 1151 446 1155 447
rect 1151 441 1155 442
rect 1199 446 1203 447
rect 1199 441 1203 442
rect 1239 446 1243 447
rect 1239 441 1243 442
rect 1295 446 1299 447
rect 1295 441 1299 442
rect 1831 446 1835 447
rect 1872 443 1874 466
rect 2142 464 2143 468
rect 2147 464 2148 468
rect 2142 463 2148 464
rect 2222 468 2228 469
rect 2222 464 2223 468
rect 2227 464 2228 468
rect 2222 463 2228 464
rect 2318 468 2324 469
rect 2318 464 2319 468
rect 2323 464 2324 468
rect 2318 463 2324 464
rect 2422 468 2428 469
rect 2422 464 2423 468
rect 2427 464 2428 468
rect 2422 463 2428 464
rect 2542 468 2548 469
rect 2542 464 2543 468
rect 2547 464 2548 468
rect 2542 463 2548 464
rect 2678 468 2684 469
rect 2678 464 2679 468
rect 2683 464 2684 468
rect 2678 463 2684 464
rect 2144 443 2146 463
rect 2224 443 2226 463
rect 2320 443 2322 463
rect 2424 443 2426 463
rect 2544 443 2546 463
rect 2680 443 2682 463
rect 1831 441 1835 442
rect 1871 442 1875 443
rect 824 425 826 441
rect 920 425 922 441
rect 1008 425 1010 441
rect 1104 425 1106 441
rect 1200 425 1202 441
rect 1296 425 1298 441
rect 822 424 828 425
rect 822 420 823 424
rect 827 420 828 424
rect 822 419 828 420
rect 918 424 924 425
rect 918 420 919 424
rect 923 420 924 424
rect 918 419 924 420
rect 1006 424 1012 425
rect 1006 420 1007 424
rect 1011 420 1012 424
rect 1006 419 1012 420
rect 1102 424 1108 425
rect 1102 420 1103 424
rect 1107 420 1108 424
rect 1102 419 1108 420
rect 1198 424 1204 425
rect 1198 420 1199 424
rect 1203 420 1204 424
rect 1198 419 1204 420
rect 1294 424 1300 425
rect 1294 420 1295 424
rect 1299 420 1300 424
rect 1832 422 1834 441
rect 1871 437 1875 438
rect 2143 442 2147 443
rect 2143 437 2147 438
rect 2223 442 2227 443
rect 2223 437 2227 438
rect 2319 442 2323 443
rect 2319 437 2323 438
rect 2335 442 2339 443
rect 2335 437 2339 438
rect 2415 442 2419 443
rect 2415 437 2419 438
rect 2423 442 2427 443
rect 2423 437 2427 438
rect 2495 442 2499 443
rect 2495 437 2499 438
rect 2543 442 2547 443
rect 2543 437 2547 438
rect 2583 442 2587 443
rect 2583 437 2587 438
rect 2679 442 2683 443
rect 2679 437 2683 438
rect 2687 442 2691 443
rect 2687 437 2691 438
rect 1294 419 1300 420
rect 1830 421 1836 422
rect 1830 417 1831 421
rect 1835 417 1836 421
rect 1872 418 1874 437
rect 2336 421 2338 437
rect 2416 421 2418 437
rect 2496 421 2498 437
rect 2584 421 2586 437
rect 2688 421 2690 437
rect 2334 420 2340 421
rect 1830 416 1836 417
rect 1870 417 1876 418
rect 466 415 472 416
rect 466 411 467 415
rect 471 411 472 415
rect 466 410 472 411
rect 562 415 568 416
rect 562 411 563 415
rect 567 411 568 415
rect 562 410 568 411
rect 674 415 680 416
rect 674 411 675 415
rect 679 411 680 415
rect 674 410 680 411
rect 786 415 792 416
rect 786 411 787 415
rect 791 411 792 415
rect 786 410 792 411
rect 890 415 896 416
rect 890 411 891 415
rect 895 411 896 415
rect 890 410 896 411
rect 986 415 992 416
rect 986 411 987 415
rect 991 411 992 415
rect 986 410 992 411
rect 1074 415 1080 416
rect 1074 411 1075 415
rect 1079 411 1080 415
rect 1074 410 1080 411
rect 1270 415 1276 416
rect 1270 411 1271 415
rect 1275 411 1276 415
rect 1870 413 1871 417
rect 1875 413 1876 417
rect 2334 416 2335 420
rect 2339 416 2340 420
rect 2334 415 2340 416
rect 2414 420 2420 421
rect 2414 416 2415 420
rect 2419 416 2420 420
rect 2414 415 2420 416
rect 2494 420 2500 421
rect 2494 416 2495 420
rect 2499 416 2500 420
rect 2494 415 2500 416
rect 2582 420 2588 421
rect 2582 416 2583 420
rect 2587 416 2588 420
rect 2582 415 2588 416
rect 2686 420 2692 421
rect 2686 416 2687 420
rect 2691 416 2692 420
rect 2686 415 2692 416
rect 1870 412 1876 413
rect 1270 410 1276 411
rect 2402 411 2408 412
rect 502 386 508 387
rect 502 382 503 386
rect 507 382 508 386
rect 502 381 508 382
rect 394 375 400 376
rect 394 371 395 375
rect 399 371 400 375
rect 394 370 400 371
rect 504 359 506 381
rect 564 376 566 410
rect 614 386 620 387
rect 614 382 615 386
rect 619 382 620 386
rect 614 381 620 382
rect 562 375 568 376
rect 562 371 563 375
rect 567 371 568 375
rect 562 370 568 371
rect 616 359 618 381
rect 676 376 678 410
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 674 375 680 376
rect 674 371 675 375
rect 679 371 680 375
rect 674 370 680 371
rect 728 359 730 381
rect 782 375 788 376
rect 782 371 783 375
rect 787 371 788 375
rect 782 370 788 371
rect 247 358 251 359
rect 247 353 251 354
rect 255 358 259 359
rect 255 353 259 354
rect 375 358 379 359
rect 375 353 379 354
rect 383 358 387 359
rect 383 353 387 354
rect 503 358 507 359
rect 503 353 507 354
rect 511 358 515 359
rect 511 353 515 354
rect 615 358 619 359
rect 615 353 619 354
rect 647 358 651 359
rect 647 353 651 354
rect 727 358 731 359
rect 727 353 731 354
rect 775 358 779 359
rect 775 353 779 354
rect 194 351 200 352
rect 194 347 195 351
rect 199 347 200 351
rect 194 346 200 347
rect 248 343 250 353
rect 298 351 304 352
rect 298 347 299 351
rect 303 347 304 351
rect 298 346 304 347
rect 142 342 148 343
rect 142 338 143 342
rect 147 338 148 342
rect 142 337 148 338
rect 246 342 252 343
rect 246 338 247 342
rect 251 338 252 342
rect 246 337 252 338
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 110 319 116 320
rect 300 316 302 346
rect 376 343 378 353
rect 426 351 432 352
rect 426 347 427 351
rect 431 347 432 351
rect 426 346 432 347
rect 374 342 380 343
rect 374 338 375 342
rect 379 338 380 342
rect 374 337 380 338
rect 428 316 430 346
rect 512 343 514 353
rect 648 343 650 353
rect 662 351 668 352
rect 662 347 663 351
rect 667 347 668 351
rect 662 346 668 347
rect 698 351 704 352
rect 698 347 699 351
rect 703 347 704 351
rect 698 346 704 347
rect 510 342 516 343
rect 510 338 511 342
rect 515 338 516 342
rect 510 337 516 338
rect 646 342 652 343
rect 646 338 647 342
rect 651 338 652 342
rect 646 337 652 338
rect 298 315 304 316
rect 298 311 299 315
rect 303 311 304 315
rect 298 310 304 311
rect 426 315 432 316
rect 426 311 427 315
rect 431 311 432 315
rect 426 310 432 311
rect 110 307 116 308
rect 110 303 111 307
rect 115 303 116 307
rect 110 302 116 303
rect 134 304 140 305
rect 112 275 114 302
rect 134 300 135 304
rect 139 300 140 304
rect 134 299 140 300
rect 238 304 244 305
rect 238 300 239 304
rect 243 300 244 304
rect 238 299 244 300
rect 366 304 372 305
rect 366 300 367 304
rect 371 300 372 304
rect 366 299 372 300
rect 502 304 508 305
rect 502 300 503 304
rect 507 300 508 304
rect 502 299 508 300
rect 638 304 644 305
rect 638 300 639 304
rect 643 300 644 304
rect 638 299 644 300
rect 136 275 138 299
rect 240 275 242 299
rect 368 275 370 299
rect 504 275 506 299
rect 510 287 516 288
rect 510 283 511 287
rect 515 283 516 287
rect 510 282 516 283
rect 111 274 115 275
rect 111 269 115 270
rect 135 274 139 275
rect 135 269 139 270
rect 223 274 227 275
rect 223 269 227 270
rect 239 274 243 275
rect 239 269 243 270
rect 335 274 339 275
rect 335 269 339 270
rect 367 274 371 275
rect 367 269 371 270
rect 463 274 467 275
rect 463 269 467 270
rect 503 274 507 275
rect 503 269 507 270
rect 112 250 114 269
rect 224 253 226 269
rect 336 253 338 269
rect 464 253 466 269
rect 222 252 228 253
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 222 248 223 252
rect 227 248 228 252
rect 222 247 228 248
rect 334 252 340 253
rect 334 248 335 252
rect 339 248 340 252
rect 334 247 340 248
rect 462 252 468 253
rect 462 248 463 252
rect 467 248 468 252
rect 462 247 468 248
rect 110 244 116 245
rect 186 243 192 244
rect 186 239 187 243
rect 191 239 192 243
rect 186 238 192 239
rect 290 243 296 244
rect 290 239 291 243
rect 295 239 296 243
rect 290 238 296 239
rect 402 243 408 244
rect 402 239 403 243
rect 407 239 408 243
rect 402 238 408 239
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 110 227 116 228
rect 112 167 114 227
rect 111 166 115 167
rect 111 161 115 162
rect 159 166 163 167
rect 159 161 163 162
rect 112 133 114 161
rect 160 151 162 161
rect 188 160 190 238
rect 230 214 236 215
rect 230 210 231 214
rect 235 210 236 214
rect 230 209 236 210
rect 232 167 234 209
rect 292 204 294 238
rect 342 214 348 215
rect 342 210 343 214
rect 347 210 348 214
rect 342 209 348 210
rect 290 203 296 204
rect 290 199 291 203
rect 295 199 296 203
rect 290 198 296 199
rect 344 167 346 209
rect 404 204 406 238
rect 470 214 476 215
rect 470 210 471 214
rect 475 210 476 214
rect 470 209 476 210
rect 402 203 408 204
rect 402 199 403 203
rect 407 199 408 203
rect 402 198 408 199
rect 472 167 474 209
rect 512 204 514 282
rect 640 275 642 299
rect 599 274 603 275
rect 599 269 603 270
rect 639 274 643 275
rect 639 269 643 270
rect 600 253 602 269
rect 664 253 666 346
rect 700 316 702 346
rect 776 343 778 353
rect 774 342 780 343
rect 774 338 775 342
rect 779 338 780 342
rect 774 337 780 338
rect 784 316 786 370
rect 832 359 834 381
rect 892 376 894 410
rect 926 386 932 387
rect 926 382 927 386
rect 931 382 932 386
rect 926 381 932 382
rect 890 375 896 376
rect 890 371 891 375
rect 895 371 896 375
rect 890 370 896 371
rect 928 359 930 381
rect 988 376 990 410
rect 1014 386 1020 387
rect 1014 382 1015 386
rect 1019 382 1020 386
rect 1014 381 1020 382
rect 986 375 992 376
rect 986 371 987 375
rect 991 371 992 375
rect 986 370 992 371
rect 1016 359 1018 381
rect 1076 376 1078 410
rect 1162 407 1168 408
rect 1162 403 1163 407
rect 1167 403 1168 407
rect 1162 402 1168 403
rect 1110 386 1116 387
rect 1110 382 1111 386
rect 1115 382 1116 386
rect 1110 381 1116 382
rect 1074 375 1080 376
rect 1074 371 1075 375
rect 1079 371 1080 375
rect 1074 370 1080 371
rect 1112 359 1114 381
rect 1164 376 1166 402
rect 1206 386 1212 387
rect 1206 382 1207 386
rect 1211 382 1212 386
rect 1206 381 1212 382
rect 1162 375 1168 376
rect 1162 371 1163 375
rect 1167 371 1168 375
rect 1162 370 1168 371
rect 1170 375 1176 376
rect 1170 371 1171 375
rect 1175 371 1176 375
rect 1170 370 1176 371
rect 831 358 835 359
rect 831 353 835 354
rect 895 358 899 359
rect 895 353 899 354
rect 927 358 931 359
rect 927 353 931 354
rect 1007 358 1011 359
rect 1007 353 1011 354
rect 1015 358 1019 359
rect 1015 353 1019 354
rect 1111 358 1115 359
rect 1111 353 1115 354
rect 1119 358 1123 359
rect 1119 353 1123 354
rect 896 343 898 353
rect 1008 343 1010 353
rect 1030 351 1036 352
rect 1030 347 1031 351
rect 1035 347 1036 351
rect 1030 346 1036 347
rect 1058 351 1064 352
rect 1058 347 1059 351
rect 1063 347 1064 351
rect 1058 346 1064 347
rect 894 342 900 343
rect 894 338 895 342
rect 899 338 900 342
rect 894 337 900 338
rect 1006 342 1012 343
rect 1006 338 1007 342
rect 1011 338 1012 342
rect 1006 337 1012 338
rect 698 315 704 316
rect 698 311 699 315
rect 703 311 704 315
rect 698 310 704 311
rect 782 315 788 316
rect 782 311 783 315
rect 787 311 788 315
rect 782 310 788 311
rect 1006 315 1012 316
rect 1006 311 1007 315
rect 1011 314 1012 315
rect 1032 314 1034 346
rect 1060 316 1062 346
rect 1120 343 1122 353
rect 1118 342 1124 343
rect 1118 338 1119 342
rect 1123 338 1124 342
rect 1118 337 1124 338
rect 1172 316 1174 370
rect 1208 359 1210 381
rect 1272 376 1274 410
rect 2402 407 2403 411
rect 2407 407 2408 411
rect 2402 406 2408 407
rect 2482 411 2488 412
rect 2482 407 2483 411
rect 2487 407 2488 411
rect 2482 406 2488 407
rect 2562 411 2568 412
rect 2562 407 2563 411
rect 2567 407 2568 411
rect 2562 406 2568 407
rect 2650 411 2656 412
rect 2650 407 2651 411
rect 2655 407 2656 411
rect 2650 406 2656 407
rect 1830 404 1836 405
rect 1830 400 1831 404
rect 1835 400 1836 404
rect 2394 403 2400 404
rect 1830 399 1836 400
rect 1870 400 1876 401
rect 1302 386 1308 387
rect 1302 382 1303 386
rect 1307 382 1308 386
rect 1302 381 1308 382
rect 1270 375 1276 376
rect 1270 371 1271 375
rect 1275 371 1276 375
rect 1270 370 1276 371
rect 1230 359 1236 360
rect 1304 359 1306 381
rect 1446 359 1452 360
rect 1832 359 1834 399
rect 1870 396 1871 400
rect 1875 396 1876 400
rect 2394 399 2395 403
rect 2399 399 2400 403
rect 2394 398 2400 399
rect 1870 395 1876 396
rect 1872 359 1874 395
rect 2342 382 2348 383
rect 2342 378 2343 382
rect 2347 378 2348 382
rect 2342 377 2348 378
rect 2270 359 2276 360
rect 2344 359 2346 377
rect 2396 372 2398 398
rect 2404 372 2406 406
rect 2422 382 2428 383
rect 2422 378 2423 382
rect 2427 378 2428 382
rect 2422 377 2428 378
rect 2394 371 2400 372
rect 2394 367 2395 371
rect 2399 367 2400 371
rect 2394 366 2400 367
rect 2402 371 2408 372
rect 2402 367 2403 371
rect 2407 367 2408 371
rect 2402 366 2408 367
rect 2424 359 2426 377
rect 2484 376 2486 406
rect 2502 382 2508 383
rect 2502 378 2503 382
rect 2507 378 2508 382
rect 2502 377 2508 378
rect 2482 375 2488 376
rect 2482 371 2483 375
rect 2487 371 2488 375
rect 2482 370 2488 371
rect 2504 359 2506 377
rect 2518 375 2524 376
rect 2518 371 2519 375
rect 2523 371 2524 375
rect 2564 372 2566 406
rect 2590 382 2596 383
rect 2590 378 2591 382
rect 2595 378 2596 382
rect 2590 377 2596 378
rect 2562 371 2568 372
rect 2518 370 2530 371
rect 2520 369 2530 370
rect 1207 358 1211 359
rect 1207 353 1211 354
rect 1223 358 1227 359
rect 1230 355 1231 359
rect 1235 355 1236 359
rect 1230 354 1236 355
rect 1303 358 1307 359
rect 1223 353 1227 354
rect 1224 343 1226 353
rect 1222 342 1228 343
rect 1222 338 1223 342
rect 1227 338 1228 342
rect 1222 337 1228 338
rect 1232 316 1234 354
rect 1303 353 1307 354
rect 1327 358 1331 359
rect 1327 353 1331 354
rect 1439 358 1443 359
rect 1446 355 1447 359
rect 1451 355 1452 359
rect 1446 354 1452 355
rect 1831 358 1835 359
rect 1439 353 1443 354
rect 1328 343 1330 353
rect 1342 351 1348 352
rect 1342 347 1343 351
rect 1347 347 1348 351
rect 1342 346 1348 347
rect 1378 351 1384 352
rect 1378 347 1379 351
rect 1383 347 1384 351
rect 1378 346 1384 347
rect 1326 342 1332 343
rect 1326 338 1327 342
rect 1331 338 1332 342
rect 1326 337 1332 338
rect 1011 312 1034 314
rect 1058 315 1064 316
rect 1011 311 1012 312
rect 1006 310 1012 311
rect 1058 311 1059 315
rect 1063 311 1064 315
rect 1058 310 1064 311
rect 1170 315 1176 316
rect 1170 311 1171 315
rect 1175 311 1176 315
rect 1170 310 1176 311
rect 1230 315 1236 316
rect 1230 311 1231 315
rect 1235 311 1236 315
rect 1230 310 1236 311
rect 766 304 772 305
rect 766 300 767 304
rect 771 300 772 304
rect 766 299 772 300
rect 886 304 892 305
rect 886 300 887 304
rect 891 300 892 304
rect 886 299 892 300
rect 998 304 1004 305
rect 998 300 999 304
rect 1003 300 1004 304
rect 998 299 1004 300
rect 1110 304 1116 305
rect 1110 300 1111 304
rect 1115 300 1116 304
rect 1110 299 1116 300
rect 1214 304 1220 305
rect 1214 300 1215 304
rect 1219 300 1220 304
rect 1214 299 1220 300
rect 1318 304 1324 305
rect 1318 300 1319 304
rect 1323 300 1324 304
rect 1318 299 1324 300
rect 768 275 770 299
rect 888 275 890 299
rect 1000 275 1002 299
rect 1112 275 1114 299
rect 1216 275 1218 299
rect 1320 275 1322 299
rect 735 274 739 275
rect 735 269 739 270
rect 767 274 771 275
rect 767 269 771 270
rect 871 274 875 275
rect 871 269 875 270
rect 887 274 891 275
rect 887 269 891 270
rect 999 274 1003 275
rect 999 269 1003 270
rect 1007 274 1011 275
rect 1007 269 1011 270
rect 1111 274 1115 275
rect 1111 269 1115 270
rect 1135 274 1139 275
rect 1135 269 1139 270
rect 1215 274 1219 275
rect 1215 269 1219 270
rect 1255 274 1259 275
rect 1255 269 1259 270
rect 1319 274 1323 275
rect 1319 269 1323 270
rect 736 253 738 269
rect 872 253 874 269
rect 1008 253 1010 269
rect 1136 253 1138 269
rect 1256 253 1258 269
rect 598 252 604 253
rect 598 248 599 252
rect 603 248 604 252
rect 598 247 604 248
rect 660 251 666 253
rect 734 252 740 253
rect 660 236 662 251
rect 734 248 735 252
rect 739 248 740 252
rect 734 247 740 248
rect 870 252 876 253
rect 870 248 871 252
rect 875 248 876 252
rect 870 247 876 248
rect 1006 252 1012 253
rect 1006 248 1007 252
rect 1011 248 1012 252
rect 1006 247 1012 248
rect 1134 252 1140 253
rect 1134 248 1135 252
rect 1139 248 1140 252
rect 1134 247 1140 248
rect 1254 252 1260 253
rect 1254 248 1255 252
rect 1259 248 1260 252
rect 1254 247 1260 248
rect 1344 244 1346 346
rect 1380 316 1382 346
rect 1440 343 1442 353
rect 1438 342 1444 343
rect 1438 338 1439 342
rect 1443 338 1444 342
rect 1438 337 1444 338
rect 1448 316 1450 354
rect 1831 353 1835 354
rect 1871 358 1875 359
rect 1871 353 1875 354
rect 2079 358 2083 359
rect 2079 353 2083 354
rect 2167 358 2171 359
rect 2167 353 2171 354
rect 2263 358 2267 359
rect 2270 355 2271 359
rect 2275 355 2276 359
rect 2270 354 2276 355
rect 2343 358 2347 359
rect 2263 353 2267 354
rect 1832 325 1834 353
rect 1872 325 1874 353
rect 2080 343 2082 353
rect 2130 351 2136 352
rect 2130 347 2131 351
rect 2135 347 2136 351
rect 2130 346 2136 347
rect 2078 342 2084 343
rect 2078 338 2079 342
rect 2083 338 2084 342
rect 2078 337 2084 338
rect 1830 324 1836 325
rect 1830 320 1831 324
rect 1835 320 1836 324
rect 1830 319 1836 320
rect 1870 324 1876 325
rect 1870 320 1871 324
rect 1875 320 1876 324
rect 1870 319 1876 320
rect 2132 316 2134 346
rect 2168 343 2170 353
rect 2264 343 2266 353
rect 2166 342 2172 343
rect 2166 338 2167 342
rect 2171 338 2172 342
rect 2166 337 2172 338
rect 2262 342 2268 343
rect 2262 338 2263 342
rect 2267 338 2268 342
rect 2262 337 2268 338
rect 2272 316 2274 354
rect 2343 353 2347 354
rect 2375 358 2379 359
rect 2375 353 2379 354
rect 2423 358 2427 359
rect 2423 353 2427 354
rect 2503 358 2507 359
rect 2503 353 2507 354
rect 2376 343 2378 353
rect 2382 351 2388 352
rect 2382 347 2383 351
rect 2387 347 2388 351
rect 2382 346 2388 347
rect 2374 342 2380 343
rect 2374 338 2375 342
rect 2379 338 2380 342
rect 2374 337 2380 338
rect 2384 316 2386 346
rect 2504 343 2506 353
rect 2528 352 2530 369
rect 2562 367 2563 371
rect 2567 367 2568 371
rect 2562 366 2568 367
rect 2592 359 2594 377
rect 2652 372 2654 406
rect 2694 382 2700 383
rect 2694 378 2695 382
rect 2699 378 2700 382
rect 2694 377 2700 378
rect 2650 371 2656 372
rect 2650 367 2651 371
rect 2655 367 2656 371
rect 2650 366 2656 367
rect 2646 359 2652 360
rect 2696 359 2698 377
rect 2720 372 2722 474
rect 2830 468 2836 469
rect 2830 464 2831 468
rect 2835 464 2836 468
rect 2830 463 2836 464
rect 2990 468 2996 469
rect 2990 464 2991 468
rect 2995 464 2996 468
rect 2990 463 2996 464
rect 2832 443 2834 463
rect 2992 443 2994 463
rect 2799 442 2803 443
rect 2799 437 2803 438
rect 2831 442 2835 443
rect 2831 437 2835 438
rect 2927 442 2931 443
rect 2927 437 2931 438
rect 2991 442 2995 443
rect 2991 437 2995 438
rect 2800 421 2802 437
rect 2928 421 2930 437
rect 2798 420 2804 421
rect 2798 416 2799 420
rect 2803 416 2804 420
rect 2798 415 2804 416
rect 2926 420 2932 421
rect 2926 416 2927 420
rect 2931 416 2932 420
rect 2926 415 2932 416
rect 2866 411 2872 412
rect 2798 407 2804 408
rect 2798 403 2799 407
rect 2803 403 2804 407
rect 2866 407 2867 411
rect 2871 407 2872 411
rect 2866 406 2872 407
rect 2994 411 3000 412
rect 2994 407 2995 411
rect 2999 407 3000 411
rect 2994 406 3000 407
rect 2798 402 2804 403
rect 2718 371 2724 372
rect 2718 367 2719 371
rect 2723 367 2724 371
rect 2718 366 2724 367
rect 2591 358 2595 359
rect 2591 353 2595 354
rect 2639 358 2643 359
rect 2646 355 2647 359
rect 2651 355 2652 359
rect 2646 354 2652 355
rect 2695 358 2699 359
rect 2639 353 2643 354
rect 2526 351 2532 352
rect 2526 347 2527 351
rect 2531 347 2532 351
rect 2526 346 2532 347
rect 2554 351 2560 352
rect 2554 347 2555 351
rect 2559 347 2560 351
rect 2554 346 2560 347
rect 2502 342 2508 343
rect 2502 338 2503 342
rect 2507 338 2508 342
rect 2502 337 2508 338
rect 2556 316 2558 346
rect 2640 343 2642 353
rect 2638 342 2644 343
rect 2638 338 2639 342
rect 2643 338 2644 342
rect 2638 337 2644 338
rect 2648 316 2650 354
rect 2695 353 2699 354
rect 2775 358 2779 359
rect 2775 353 2779 354
rect 2776 343 2778 353
rect 2800 352 2802 402
rect 2806 382 2812 383
rect 2806 378 2807 382
rect 2811 378 2812 382
rect 2806 377 2812 378
rect 2808 359 2810 377
rect 2868 372 2870 406
rect 2934 382 2940 383
rect 2934 378 2935 382
rect 2939 378 2940 382
rect 2934 377 2940 378
rect 2866 371 2872 372
rect 2866 367 2867 371
rect 2871 367 2872 371
rect 2866 366 2872 367
rect 2936 359 2938 377
rect 2996 372 2998 406
rect 3052 372 3054 474
rect 3166 468 3172 469
rect 3166 464 3167 468
rect 3171 464 3172 468
rect 3166 463 3172 464
rect 3168 443 3170 463
rect 3071 442 3075 443
rect 3071 437 3075 438
rect 3167 442 3171 443
rect 3167 437 3171 438
rect 3072 421 3074 437
rect 3070 420 3076 421
rect 3070 416 3071 420
rect 3075 416 3076 420
rect 3070 415 3076 416
rect 3204 412 3206 510
rect 3228 480 3230 510
rect 3352 507 3354 517
rect 3350 506 3356 507
rect 3350 502 3351 506
rect 3355 502 3356 506
rect 3350 501 3356 502
rect 3368 480 3370 522
rect 3511 517 3515 518
rect 3512 507 3514 517
rect 3564 516 3566 554
rect 3590 552 3591 556
rect 3595 552 3596 556
rect 3590 551 3596 552
rect 3592 523 3594 551
rect 3591 522 3595 523
rect 3591 517 3595 518
rect 3562 515 3568 516
rect 3562 511 3563 515
rect 3567 511 3568 515
rect 3562 510 3568 511
rect 3510 506 3516 507
rect 3510 502 3511 506
rect 3515 502 3516 506
rect 3510 501 3516 502
rect 3592 489 3594 517
rect 3590 488 3596 489
rect 3590 484 3591 488
rect 3595 484 3596 488
rect 3590 483 3596 484
rect 3226 479 3232 480
rect 3226 475 3227 479
rect 3231 475 3232 479
rect 3226 474 3232 475
rect 3366 479 3372 480
rect 3366 475 3367 479
rect 3371 475 3372 479
rect 3366 474 3372 475
rect 3534 479 3540 480
rect 3534 475 3535 479
rect 3539 475 3540 479
rect 3534 474 3540 475
rect 3342 468 3348 469
rect 3342 464 3343 468
rect 3347 464 3348 468
rect 3342 463 3348 464
rect 3502 468 3508 469
rect 3502 464 3503 468
rect 3507 464 3508 468
rect 3502 463 3508 464
rect 3344 443 3346 463
rect 3504 443 3506 463
rect 3215 442 3219 443
rect 3215 437 3219 438
rect 3343 442 3347 443
rect 3343 437 3347 438
rect 3367 442 3371 443
rect 3367 437 3371 438
rect 3503 442 3507 443
rect 3503 437 3507 438
rect 3216 421 3218 437
rect 3368 421 3370 437
rect 3504 421 3506 437
rect 3214 420 3220 421
rect 3214 416 3215 420
rect 3219 416 3220 420
rect 3214 415 3220 416
rect 3366 420 3372 421
rect 3366 416 3367 420
rect 3371 416 3372 420
rect 3366 415 3372 416
rect 3502 420 3508 421
rect 3502 416 3503 420
rect 3507 416 3508 420
rect 3502 415 3508 416
rect 3202 411 3208 412
rect 3202 407 3203 411
rect 3207 407 3208 411
rect 3202 406 3208 407
rect 3282 411 3288 412
rect 3282 407 3283 411
rect 3287 407 3288 411
rect 3282 406 3288 407
rect 3434 411 3440 412
rect 3434 407 3435 411
rect 3439 407 3440 411
rect 3434 406 3440 407
rect 3078 382 3084 383
rect 3078 378 3079 382
rect 3083 378 3084 382
rect 3078 377 3084 378
rect 3222 382 3228 383
rect 3222 378 3223 382
rect 3227 378 3228 382
rect 3222 377 3228 378
rect 2994 371 3000 372
rect 2994 367 2995 371
rect 2999 367 3000 371
rect 2994 366 3000 367
rect 3050 371 3056 372
rect 3050 367 3051 371
rect 3055 367 3056 371
rect 3050 366 3056 367
rect 3080 359 3082 377
rect 3224 359 3226 377
rect 3284 372 3286 406
rect 3374 382 3380 383
rect 3374 378 3375 382
rect 3379 378 3380 382
rect 3374 377 3380 378
rect 3282 371 3288 372
rect 3282 367 3283 371
rect 3287 367 3288 371
rect 3282 366 3288 367
rect 3338 371 3344 372
rect 3338 367 3339 371
rect 3343 367 3344 371
rect 3338 366 3344 367
rect 2807 358 2811 359
rect 2807 353 2811 354
rect 2911 358 2915 359
rect 2911 353 2915 354
rect 2935 358 2939 359
rect 2935 353 2939 354
rect 3039 358 3043 359
rect 3039 353 3043 354
rect 3079 358 3083 359
rect 3079 353 3083 354
rect 3167 358 3171 359
rect 3167 353 3171 354
rect 3223 358 3227 359
rect 3223 353 3227 354
rect 3287 358 3291 359
rect 3287 353 3291 354
rect 2798 351 2804 352
rect 2798 347 2799 351
rect 2803 347 2804 351
rect 2798 346 2804 347
rect 2826 351 2832 352
rect 2826 347 2827 351
rect 2831 347 2832 351
rect 2826 346 2832 347
rect 2774 342 2780 343
rect 2774 338 2775 342
rect 2779 338 2780 342
rect 2774 337 2780 338
rect 2828 316 2830 346
rect 2912 343 2914 353
rect 3040 343 3042 353
rect 3066 351 3072 352
rect 3066 347 3067 351
rect 3071 347 3072 351
rect 3066 346 3072 347
rect 3090 351 3096 352
rect 3090 347 3091 351
rect 3095 347 3096 351
rect 3090 346 3096 347
rect 2910 342 2916 343
rect 2910 338 2911 342
rect 2915 338 2916 342
rect 2910 337 2916 338
rect 3038 342 3044 343
rect 3038 338 3039 342
rect 3043 338 3044 342
rect 3038 337 3044 338
rect 1378 315 1384 316
rect 1378 311 1379 315
rect 1383 311 1384 315
rect 1378 310 1384 311
rect 1446 315 1452 316
rect 1446 311 1447 315
rect 1451 311 1452 315
rect 1446 310 1452 311
rect 2130 315 2136 316
rect 2130 311 2131 315
rect 2135 311 2136 315
rect 2130 310 2136 311
rect 2238 315 2244 316
rect 2238 311 2239 315
rect 2243 311 2244 315
rect 2238 310 2244 311
rect 2270 315 2276 316
rect 2270 311 2271 315
rect 2275 311 2276 315
rect 2270 310 2276 311
rect 2382 315 2388 316
rect 2382 311 2383 315
rect 2387 311 2388 315
rect 2382 310 2388 311
rect 2554 315 2560 316
rect 2554 311 2555 315
rect 2559 311 2560 315
rect 2554 310 2560 311
rect 2646 315 2652 316
rect 2646 311 2647 315
rect 2651 311 2652 315
rect 2646 310 2652 311
rect 2826 315 2832 316
rect 2826 311 2827 315
rect 2831 311 2832 315
rect 2826 310 2832 311
rect 2962 315 2968 316
rect 2962 311 2963 315
rect 2967 311 2968 315
rect 2962 310 2968 311
rect 1830 307 1836 308
rect 1430 304 1436 305
rect 1430 300 1431 304
rect 1435 300 1436 304
rect 1830 303 1831 307
rect 1835 303 1836 307
rect 1830 302 1836 303
rect 1870 307 1876 308
rect 1870 303 1871 307
rect 1875 303 1876 307
rect 1870 302 1876 303
rect 2070 304 2076 305
rect 1430 299 1436 300
rect 1432 275 1434 299
rect 1832 275 1834 302
rect 1872 275 1874 302
rect 2070 300 2071 304
rect 2075 300 2076 304
rect 2070 299 2076 300
rect 2158 304 2164 305
rect 2158 300 2159 304
rect 2163 300 2164 304
rect 2158 299 2164 300
rect 2072 275 2074 299
rect 2160 275 2162 299
rect 1367 274 1371 275
rect 1367 269 1371 270
rect 1431 274 1435 275
rect 1431 269 1435 270
rect 1479 274 1483 275
rect 1479 269 1483 270
rect 1599 274 1603 275
rect 1599 269 1603 270
rect 1831 274 1835 275
rect 1831 269 1835 270
rect 1871 274 1875 275
rect 1871 269 1875 270
rect 1895 274 1899 275
rect 1895 269 1899 270
rect 1983 274 1987 275
rect 1983 269 1987 270
rect 2071 274 2075 275
rect 2071 269 2075 270
rect 2095 274 2099 275
rect 2095 269 2099 270
rect 2159 274 2163 275
rect 2159 269 2163 270
rect 2223 274 2227 275
rect 2223 269 2227 270
rect 1368 253 1370 269
rect 1480 253 1482 269
rect 1600 253 1602 269
rect 1366 252 1372 253
rect 1366 248 1367 252
rect 1371 248 1372 252
rect 1366 247 1372 248
rect 1478 252 1484 253
rect 1478 248 1479 252
rect 1483 248 1484 252
rect 1478 247 1484 248
rect 1598 252 1604 253
rect 1598 248 1599 252
rect 1603 248 1604 252
rect 1832 250 1834 269
rect 1872 250 1874 269
rect 1896 253 1898 269
rect 1984 253 1986 269
rect 2096 253 2098 269
rect 2224 253 2226 269
rect 1894 252 1900 253
rect 1598 247 1604 248
rect 1830 249 1836 250
rect 1830 245 1831 249
rect 1835 245 1836 249
rect 1830 244 1836 245
rect 1870 249 1876 250
rect 1870 245 1871 249
rect 1875 245 1876 249
rect 1894 248 1895 252
rect 1899 248 1900 252
rect 1894 247 1900 248
rect 1982 252 1988 253
rect 1982 248 1983 252
rect 1987 248 1988 252
rect 1982 247 1988 248
rect 2094 252 2100 253
rect 2094 248 2095 252
rect 2099 248 2100 252
rect 2094 247 2100 248
rect 2222 252 2228 253
rect 2222 248 2223 252
rect 2227 248 2228 252
rect 2222 247 2228 248
rect 1870 244 1876 245
rect 666 243 672 244
rect 666 239 667 243
rect 671 239 672 243
rect 666 238 672 239
rect 802 243 808 244
rect 802 239 803 243
rect 807 239 808 243
rect 802 238 808 239
rect 1078 243 1084 244
rect 1078 239 1079 243
rect 1083 239 1084 243
rect 1078 238 1084 239
rect 1210 243 1216 244
rect 1210 239 1211 243
rect 1215 239 1216 243
rect 1210 238 1216 239
rect 1342 243 1348 244
rect 1342 239 1343 243
rect 1347 239 1348 243
rect 1342 238 1348 239
rect 1446 243 1452 244
rect 1446 239 1447 243
rect 1451 239 1452 243
rect 1446 238 1452 239
rect 1562 243 1568 244
rect 1562 239 1563 243
rect 1567 239 1568 243
rect 1562 238 1568 239
rect 1570 243 1576 244
rect 1570 239 1571 243
rect 1575 239 1576 243
rect 1570 238 1576 239
rect 1962 243 1968 244
rect 1962 239 1963 243
rect 1967 239 1968 243
rect 1962 238 1968 239
rect 2062 243 2068 244
rect 2062 239 2063 243
rect 2067 239 2068 243
rect 2062 238 2068 239
rect 2162 243 2168 244
rect 2162 239 2163 243
rect 2167 239 2168 243
rect 2162 238 2168 239
rect 658 235 664 236
rect 658 231 659 235
rect 663 231 664 235
rect 658 230 664 231
rect 606 214 612 215
rect 606 210 607 214
rect 611 210 612 214
rect 606 209 612 210
rect 510 203 516 204
rect 510 199 511 203
rect 515 199 516 203
rect 510 198 516 199
rect 608 167 610 209
rect 668 204 670 238
rect 742 214 748 215
rect 742 210 743 214
rect 747 210 748 214
rect 742 209 748 210
rect 666 203 672 204
rect 666 199 667 203
rect 671 199 672 203
rect 666 198 672 199
rect 744 167 746 209
rect 804 204 806 238
rect 878 214 884 215
rect 878 210 879 214
rect 883 210 884 214
rect 878 209 884 210
rect 1014 214 1020 215
rect 1014 210 1015 214
rect 1019 210 1020 214
rect 1014 209 1020 210
rect 1043 212 1047 213
rect 802 203 808 204
rect 802 199 803 203
rect 807 199 808 203
rect 802 198 808 199
rect 880 167 882 209
rect 902 203 908 204
rect 902 199 903 203
rect 907 199 908 203
rect 902 198 908 199
rect 231 166 235 167
rect 231 161 235 162
rect 239 166 243 167
rect 239 161 243 162
rect 319 166 323 167
rect 319 161 323 162
rect 343 166 347 167
rect 343 161 347 162
rect 399 166 403 167
rect 399 161 403 162
rect 471 166 475 167
rect 471 161 475 162
rect 479 166 483 167
rect 479 161 483 162
rect 559 166 563 167
rect 559 161 563 162
rect 607 166 611 167
rect 607 161 611 162
rect 647 166 651 167
rect 647 161 651 162
rect 735 166 739 167
rect 735 161 739 162
rect 743 166 747 167
rect 743 161 747 162
rect 823 166 827 167
rect 823 161 827 162
rect 879 166 883 167
rect 879 161 883 162
rect 186 159 192 160
rect 186 155 187 159
rect 191 155 192 159
rect 186 154 192 155
rect 210 159 216 160
rect 210 155 211 159
rect 215 155 216 159
rect 210 154 216 155
rect 158 150 164 151
rect 158 146 159 150
rect 163 146 164 150
rect 158 145 164 146
rect 110 132 116 133
rect 110 128 111 132
rect 115 128 116 132
rect 110 127 116 128
rect 212 124 214 154
rect 240 151 242 161
rect 290 159 296 160
rect 290 155 291 159
rect 295 155 296 159
rect 290 154 296 155
rect 238 150 244 151
rect 238 146 239 150
rect 243 146 244 150
rect 238 145 244 146
rect 292 124 294 154
rect 320 151 322 161
rect 370 159 376 160
rect 370 155 371 159
rect 375 155 376 159
rect 370 154 376 155
rect 318 150 324 151
rect 318 146 319 150
rect 323 146 324 150
rect 318 145 324 146
rect 372 124 374 154
rect 400 151 402 161
rect 450 159 456 160
rect 450 155 451 159
rect 455 155 456 159
rect 450 154 456 155
rect 398 150 404 151
rect 398 146 399 150
rect 403 146 404 150
rect 398 145 404 146
rect 452 124 454 154
rect 480 151 482 161
rect 530 159 536 160
rect 530 155 531 159
rect 535 155 536 159
rect 530 154 536 155
rect 478 150 484 151
rect 478 146 479 150
rect 483 146 484 150
rect 478 145 484 146
rect 532 124 534 154
rect 560 151 562 161
rect 638 159 644 160
rect 638 155 639 159
rect 643 155 644 159
rect 638 154 644 155
rect 558 150 564 151
rect 558 146 559 150
rect 563 146 564 150
rect 558 145 564 146
rect 640 124 642 154
rect 648 151 650 161
rect 698 159 704 160
rect 698 155 699 159
rect 703 155 704 159
rect 698 154 704 155
rect 646 150 652 151
rect 646 146 647 150
rect 651 146 652 150
rect 646 145 652 146
rect 700 124 702 154
rect 736 151 738 161
rect 786 159 792 160
rect 786 155 787 159
rect 791 155 792 159
rect 786 154 792 155
rect 734 150 740 151
rect 734 146 735 150
rect 739 146 740 150
rect 734 145 740 146
rect 788 124 790 154
rect 824 151 826 161
rect 822 150 828 151
rect 822 146 823 150
rect 827 146 828 150
rect 822 145 828 146
rect 904 124 906 198
rect 1016 167 1018 209
rect 1043 207 1047 208
rect 1044 204 1046 207
rect 1080 204 1082 238
rect 1142 214 1148 215
rect 1142 210 1143 214
rect 1147 210 1148 214
rect 1142 209 1148 210
rect 1042 203 1048 204
rect 1042 199 1043 203
rect 1047 199 1048 203
rect 1042 198 1048 199
rect 1078 203 1084 204
rect 1078 199 1079 203
rect 1083 199 1084 203
rect 1078 198 1084 199
rect 1144 167 1146 209
rect 1212 204 1214 238
rect 1262 214 1268 215
rect 1262 210 1263 214
rect 1267 210 1268 214
rect 1262 209 1268 210
rect 1374 214 1380 215
rect 1374 210 1375 214
rect 1379 210 1380 214
rect 1374 209 1380 210
rect 1210 203 1216 204
rect 1210 199 1211 203
rect 1215 199 1216 203
rect 1210 198 1216 199
rect 1158 195 1164 196
rect 1158 191 1159 195
rect 1163 191 1164 195
rect 1158 190 1164 191
rect 911 166 915 167
rect 911 161 915 162
rect 999 166 1003 167
rect 999 161 1003 162
rect 1015 166 1019 167
rect 1015 161 1019 162
rect 1087 166 1091 167
rect 1087 161 1091 162
rect 1143 166 1147 167
rect 1143 161 1147 162
rect 912 151 914 161
rect 1000 151 1002 161
rect 1022 159 1028 160
rect 1022 155 1023 159
rect 1027 155 1028 159
rect 1022 154 1028 155
rect 1050 159 1056 160
rect 1050 155 1051 159
rect 1055 155 1056 159
rect 1050 154 1056 155
rect 910 150 916 151
rect 910 146 911 150
rect 915 146 916 150
rect 910 145 916 146
rect 998 150 1004 151
rect 998 146 999 150
rect 1003 146 1004 150
rect 998 145 1004 146
rect 1024 139 1026 154
rect 1000 137 1026 139
rect 1000 124 1002 137
rect 1052 124 1054 154
rect 1088 151 1090 161
rect 1086 150 1092 151
rect 1086 146 1087 150
rect 1091 146 1092 150
rect 1086 145 1092 146
rect 1160 124 1162 190
rect 1174 167 1180 168
rect 1264 167 1266 209
rect 1376 167 1378 209
rect 1448 204 1450 238
rect 1486 214 1492 215
rect 1486 210 1487 214
rect 1491 210 1492 214
rect 1486 209 1492 210
rect 1446 203 1452 204
rect 1446 199 1447 203
rect 1451 199 1452 203
rect 1446 198 1452 199
rect 1488 167 1490 209
rect 1564 204 1566 238
rect 1572 213 1574 238
rect 1830 232 1836 233
rect 1830 228 1831 232
rect 1835 228 1836 232
rect 1830 227 1836 228
rect 1870 232 1876 233
rect 1870 228 1871 232
rect 1875 228 1876 232
rect 1870 227 1876 228
rect 1606 214 1612 215
rect 1571 212 1575 213
rect 1606 210 1607 214
rect 1611 210 1612 214
rect 1606 209 1612 210
rect 1571 207 1575 208
rect 1562 203 1568 204
rect 1562 199 1563 203
rect 1567 199 1568 203
rect 1562 198 1568 199
rect 1608 167 1610 209
rect 1832 167 1834 227
rect 1872 187 1874 227
rect 1902 214 1908 215
rect 1902 210 1903 214
rect 1907 210 1908 214
rect 1902 209 1908 210
rect 1931 212 1935 213
rect 1904 187 1906 209
rect 1931 207 1935 208
rect 1932 204 1934 207
rect 1964 204 1966 238
rect 1990 214 1996 215
rect 1990 210 1991 214
rect 1995 210 1996 214
rect 1990 209 1996 210
rect 1930 203 1936 204
rect 1930 199 1931 203
rect 1935 199 1936 203
rect 1930 198 1936 199
rect 1962 203 1968 204
rect 1962 199 1963 203
rect 1967 199 1968 203
rect 1962 198 1968 199
rect 1992 187 1994 209
rect 2064 204 2066 238
rect 2102 214 2108 215
rect 2102 210 2103 214
rect 2107 210 2108 214
rect 2102 209 2108 210
rect 2062 203 2068 204
rect 2062 199 2063 203
rect 2067 199 2068 203
rect 2062 198 2068 199
rect 2104 187 2106 209
rect 1871 186 1875 187
rect 1871 181 1875 182
rect 1903 186 1907 187
rect 1903 181 1907 182
rect 1983 186 1987 187
rect 1983 181 1987 182
rect 1991 186 1995 187
rect 1991 181 1995 182
rect 2087 186 2091 187
rect 2087 181 2091 182
rect 2103 186 2107 187
rect 2103 181 2107 182
rect 1167 166 1171 167
rect 1174 163 1175 167
rect 1179 163 1180 167
rect 1174 162 1180 163
rect 1247 166 1251 167
rect 1167 161 1171 162
rect 1168 151 1170 161
rect 1166 150 1172 151
rect 1166 146 1167 150
rect 1171 146 1172 150
rect 1166 145 1172 146
rect 1176 124 1178 162
rect 1247 161 1251 162
rect 1263 166 1267 167
rect 1263 161 1267 162
rect 1335 166 1339 167
rect 1335 161 1339 162
rect 1375 166 1379 167
rect 1375 161 1379 162
rect 1423 166 1427 167
rect 1423 161 1427 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1511 166 1515 167
rect 1511 161 1515 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1607 166 1611 167
rect 1607 161 1611 162
rect 1671 166 1675 167
rect 1671 161 1675 162
rect 1751 166 1755 167
rect 1751 161 1755 162
rect 1831 166 1835 167
rect 1831 161 1835 162
rect 1248 151 1250 161
rect 1254 159 1260 160
rect 1254 155 1255 159
rect 1259 155 1260 159
rect 1254 154 1260 155
rect 1246 150 1252 151
rect 1246 146 1247 150
rect 1251 146 1252 150
rect 1246 145 1252 146
rect 1256 124 1258 154
rect 1336 151 1338 161
rect 1342 159 1348 160
rect 1342 155 1343 159
rect 1347 155 1348 159
rect 1342 154 1348 155
rect 1334 150 1340 151
rect 1334 146 1335 150
rect 1339 146 1340 150
rect 1334 145 1340 146
rect 1344 124 1346 154
rect 1424 151 1426 161
rect 1430 159 1436 160
rect 1430 155 1431 159
rect 1435 155 1436 159
rect 1430 154 1436 155
rect 1422 150 1428 151
rect 1422 146 1423 150
rect 1427 146 1428 150
rect 1422 145 1428 146
rect 1432 124 1434 154
rect 1512 151 1514 161
rect 1518 159 1524 160
rect 1518 155 1519 159
rect 1523 155 1524 159
rect 1518 154 1524 155
rect 1510 150 1516 151
rect 1510 146 1511 150
rect 1515 146 1516 150
rect 1510 145 1516 146
rect 1520 124 1522 154
rect 1592 151 1594 161
rect 1598 159 1604 160
rect 1598 155 1599 159
rect 1603 155 1604 159
rect 1598 154 1604 155
rect 1590 150 1596 151
rect 1590 146 1591 150
rect 1595 146 1596 150
rect 1590 145 1596 146
rect 1600 124 1602 154
rect 1672 151 1674 161
rect 1678 159 1684 160
rect 1678 155 1679 159
rect 1683 155 1684 159
rect 1678 154 1684 155
rect 1670 150 1676 151
rect 1670 146 1671 150
rect 1675 146 1676 150
rect 1670 145 1676 146
rect 1680 124 1682 154
rect 1752 151 1754 161
rect 1758 159 1764 160
rect 1758 155 1759 159
rect 1763 155 1764 159
rect 1758 154 1764 155
rect 1750 150 1756 151
rect 1750 146 1751 150
rect 1755 146 1756 150
rect 1750 145 1756 146
rect 1760 124 1762 154
rect 1832 133 1834 161
rect 1872 153 1874 181
rect 1904 171 1906 181
rect 1962 179 1968 180
rect 1962 175 1963 179
rect 1967 175 1968 179
rect 1962 174 1968 175
rect 1902 170 1908 171
rect 1902 166 1903 170
rect 1907 166 1908 170
rect 1902 165 1908 166
rect 1870 152 1876 153
rect 1870 148 1871 152
rect 1875 148 1876 152
rect 1870 147 1876 148
rect 1964 144 1966 174
rect 1984 171 1986 181
rect 2088 171 2090 181
rect 2164 180 2166 238
rect 2230 214 2236 215
rect 2230 210 2231 214
rect 2235 210 2236 214
rect 2230 209 2236 210
rect 2232 187 2234 209
rect 2240 204 2242 310
rect 2254 304 2260 305
rect 2254 300 2255 304
rect 2259 300 2260 304
rect 2254 299 2260 300
rect 2366 304 2372 305
rect 2366 300 2367 304
rect 2371 300 2372 304
rect 2366 299 2372 300
rect 2494 304 2500 305
rect 2494 300 2495 304
rect 2499 300 2500 304
rect 2494 299 2500 300
rect 2630 304 2636 305
rect 2630 300 2631 304
rect 2635 300 2636 304
rect 2630 299 2636 300
rect 2766 304 2772 305
rect 2766 300 2767 304
rect 2771 300 2772 304
rect 2766 299 2772 300
rect 2902 304 2908 305
rect 2902 300 2903 304
rect 2907 300 2908 304
rect 2902 299 2908 300
rect 2256 275 2258 299
rect 2368 275 2370 299
rect 2496 275 2498 299
rect 2632 275 2634 299
rect 2768 275 2770 299
rect 2904 275 2906 299
rect 2255 274 2259 275
rect 2255 269 2259 270
rect 2359 274 2363 275
rect 2359 269 2363 270
rect 2367 274 2371 275
rect 2367 269 2371 270
rect 2495 274 2499 275
rect 2495 269 2499 270
rect 2503 274 2507 275
rect 2503 269 2507 270
rect 2631 274 2635 275
rect 2631 269 2635 270
rect 2647 274 2651 275
rect 2647 269 2651 270
rect 2767 274 2771 275
rect 2767 269 2771 270
rect 2791 274 2795 275
rect 2791 269 2795 270
rect 2903 274 2907 275
rect 2903 269 2907 270
rect 2935 274 2939 275
rect 2935 269 2939 270
rect 2360 253 2362 269
rect 2504 253 2506 269
rect 2648 253 2650 269
rect 2792 253 2794 269
rect 2936 253 2938 269
rect 2358 252 2364 253
rect 2358 248 2359 252
rect 2363 248 2364 252
rect 2358 247 2364 248
rect 2502 252 2508 253
rect 2502 248 2503 252
rect 2507 248 2508 252
rect 2502 247 2508 248
rect 2646 252 2652 253
rect 2646 248 2647 252
rect 2651 248 2652 252
rect 2646 247 2652 248
rect 2790 252 2796 253
rect 2790 248 2791 252
rect 2795 248 2796 252
rect 2790 247 2796 248
rect 2934 252 2940 253
rect 2934 248 2935 252
rect 2939 248 2940 252
rect 2934 247 2940 248
rect 2314 243 2320 244
rect 2314 239 2315 243
rect 2319 239 2320 243
rect 2314 238 2320 239
rect 2450 243 2456 244
rect 2450 239 2451 243
rect 2455 239 2456 243
rect 2450 238 2456 239
rect 2458 243 2464 244
rect 2458 239 2459 243
rect 2463 239 2464 243
rect 2458 238 2464 239
rect 2610 243 2616 244
rect 2610 239 2611 243
rect 2615 239 2616 243
rect 2610 238 2616 239
rect 2714 243 2720 244
rect 2714 239 2715 243
rect 2719 239 2720 243
rect 2714 238 2720 239
rect 2878 243 2884 244
rect 2878 239 2879 243
rect 2883 239 2884 243
rect 2878 238 2884 239
rect 2316 204 2318 238
rect 2366 214 2372 215
rect 2366 210 2367 214
rect 2371 210 2372 214
rect 2366 209 2372 210
rect 2238 203 2244 204
rect 2238 199 2239 203
rect 2243 199 2244 203
rect 2238 198 2244 199
rect 2314 203 2320 204
rect 2314 199 2315 203
rect 2319 199 2320 203
rect 2314 198 2320 199
rect 2368 187 2370 209
rect 2452 204 2454 238
rect 2460 213 2462 238
rect 2510 214 2516 215
rect 2459 212 2463 213
rect 2510 210 2511 214
rect 2515 210 2516 214
rect 2510 209 2516 210
rect 2459 207 2463 208
rect 2450 203 2456 204
rect 2450 199 2451 203
rect 2455 199 2456 203
rect 2450 198 2456 199
rect 2512 187 2514 209
rect 2207 186 2211 187
rect 2207 181 2211 182
rect 2231 186 2235 187
rect 2231 181 2235 182
rect 2335 186 2339 187
rect 2335 181 2339 182
rect 2367 186 2371 187
rect 2367 181 2371 182
rect 2463 186 2467 187
rect 2463 181 2467 182
rect 2511 186 2515 187
rect 2511 181 2515 182
rect 2583 186 2587 187
rect 2583 181 2587 182
rect 2094 179 2100 180
rect 2094 175 2095 179
rect 2099 175 2100 179
rect 2162 179 2168 180
rect 2094 174 2100 175
rect 2154 175 2160 176
rect 1982 170 1988 171
rect 1982 166 1983 170
rect 1987 166 1988 170
rect 1982 165 1988 166
rect 2086 170 2092 171
rect 2086 166 2087 170
rect 2091 166 2092 170
rect 2086 165 2092 166
rect 2096 144 2098 174
rect 2154 170 2155 175
rect 2159 170 2160 175
rect 2162 175 2163 179
rect 2167 175 2168 179
rect 2162 174 2168 175
rect 2208 171 2210 181
rect 2258 179 2264 180
rect 2258 175 2259 179
rect 2263 175 2264 179
rect 2258 174 2264 175
rect 2206 170 2212 171
rect 2155 167 2159 168
rect 2206 166 2207 170
rect 2211 166 2212 170
rect 2206 165 2212 166
rect 2260 144 2262 174
rect 2336 171 2338 181
rect 2386 179 2392 180
rect 2386 175 2387 179
rect 2391 175 2392 179
rect 2386 174 2392 175
rect 2334 170 2340 171
rect 2334 166 2335 170
rect 2339 166 2340 170
rect 2334 165 2340 166
rect 2388 144 2390 174
rect 2464 171 2466 181
rect 2471 172 2475 173
rect 2462 170 2468 171
rect 2462 166 2463 170
rect 2467 166 2468 170
rect 2584 171 2586 181
rect 2612 180 2614 238
rect 2654 214 2660 215
rect 2654 210 2655 214
rect 2659 210 2660 214
rect 2654 209 2660 210
rect 2656 187 2658 209
rect 2716 204 2718 238
rect 2798 214 2804 215
rect 2798 210 2799 214
rect 2803 210 2804 214
rect 2798 209 2804 210
rect 2714 203 2720 204
rect 2714 199 2715 203
rect 2719 199 2720 203
rect 2714 198 2720 199
rect 2800 187 2802 209
rect 2880 204 2882 238
rect 2942 214 2948 215
rect 2942 210 2943 214
rect 2947 210 2948 214
rect 2942 209 2948 210
rect 2878 203 2884 204
rect 2878 199 2879 203
rect 2883 199 2884 203
rect 2878 198 2884 199
rect 2944 187 2946 209
rect 2964 204 2966 310
rect 3030 304 3036 305
rect 3030 300 3031 304
rect 3035 300 3036 304
rect 3030 299 3036 300
rect 3032 275 3034 299
rect 3031 274 3035 275
rect 3031 269 3035 270
rect 3068 244 3070 346
rect 3092 316 3094 346
rect 3168 343 3170 353
rect 3278 351 3284 352
rect 3278 347 3279 351
rect 3283 347 3284 351
rect 3278 346 3284 347
rect 3166 342 3172 343
rect 3166 338 3167 342
rect 3171 338 3172 342
rect 3166 337 3172 338
rect 3280 316 3282 346
rect 3288 343 3290 353
rect 3286 342 3292 343
rect 3286 338 3287 342
rect 3291 338 3292 342
rect 3286 337 3292 338
rect 3340 316 3342 366
rect 3376 359 3378 377
rect 3375 358 3379 359
rect 3375 353 3379 354
rect 3407 358 3411 359
rect 3407 353 3411 354
rect 3408 343 3410 353
rect 3436 352 3438 406
rect 3510 382 3516 383
rect 3510 378 3511 382
rect 3515 378 3516 382
rect 3510 377 3516 378
rect 3512 359 3514 377
rect 3536 372 3538 474
rect 3590 471 3596 472
rect 3590 467 3591 471
rect 3595 467 3596 471
rect 3590 466 3596 467
rect 3592 443 3594 466
rect 3591 442 3595 443
rect 3591 437 3595 438
rect 3592 418 3594 437
rect 3590 417 3596 418
rect 3590 413 3591 417
rect 3595 413 3596 417
rect 3590 412 3596 413
rect 3590 400 3596 401
rect 3590 396 3591 400
rect 3595 396 3596 400
rect 3590 395 3596 396
rect 3534 371 3540 372
rect 3534 367 3535 371
rect 3539 367 3540 371
rect 3534 366 3540 367
rect 3592 359 3594 395
rect 3511 358 3515 359
rect 3511 353 3515 354
rect 3591 358 3595 359
rect 3591 353 3595 354
rect 3434 351 3440 352
rect 3434 347 3435 351
rect 3439 347 3440 351
rect 3434 346 3440 347
rect 3458 351 3464 352
rect 3458 347 3459 351
rect 3463 347 3464 351
rect 3458 346 3464 347
rect 3406 342 3412 343
rect 3406 338 3407 342
rect 3411 338 3412 342
rect 3406 337 3412 338
rect 3460 316 3462 346
rect 3512 343 3514 353
rect 3510 342 3516 343
rect 3510 338 3511 342
rect 3515 338 3516 342
rect 3510 337 3516 338
rect 3592 325 3594 353
rect 3590 324 3596 325
rect 3590 320 3591 324
rect 3595 320 3596 324
rect 3590 319 3596 320
rect 3090 315 3096 316
rect 3090 311 3091 315
rect 3095 311 3096 315
rect 3090 310 3096 311
rect 3278 315 3284 316
rect 3278 311 3279 315
rect 3283 311 3284 315
rect 3278 310 3284 311
rect 3338 315 3344 316
rect 3338 311 3339 315
rect 3343 311 3344 315
rect 3338 310 3344 311
rect 3458 315 3464 316
rect 3458 311 3459 315
rect 3463 311 3464 315
rect 3458 310 3464 311
rect 3534 315 3540 316
rect 3534 311 3535 315
rect 3539 311 3540 315
rect 3534 310 3540 311
rect 3158 304 3164 305
rect 3158 300 3159 304
rect 3163 300 3164 304
rect 3158 299 3164 300
rect 3278 304 3284 305
rect 3278 300 3279 304
rect 3283 300 3284 304
rect 3278 299 3284 300
rect 3398 304 3404 305
rect 3398 300 3399 304
rect 3403 300 3404 304
rect 3398 299 3404 300
rect 3502 304 3508 305
rect 3502 300 3503 304
rect 3507 300 3508 304
rect 3502 299 3508 300
rect 3160 275 3162 299
rect 3280 275 3282 299
rect 3400 275 3402 299
rect 3504 275 3506 299
rect 3079 274 3083 275
rect 3079 269 3083 270
rect 3159 274 3163 275
rect 3159 269 3163 270
rect 3223 274 3227 275
rect 3223 269 3227 270
rect 3279 274 3283 275
rect 3279 269 3283 270
rect 3375 274 3379 275
rect 3375 269 3379 270
rect 3399 274 3403 275
rect 3399 269 3403 270
rect 3503 274 3507 275
rect 3503 269 3507 270
rect 3080 253 3082 269
rect 3224 253 3226 269
rect 3376 253 3378 269
rect 3504 253 3506 269
rect 3078 252 3084 253
rect 3078 248 3079 252
rect 3083 248 3084 252
rect 3078 247 3084 248
rect 3222 252 3228 253
rect 3222 248 3223 252
rect 3227 248 3228 252
rect 3222 247 3228 248
rect 3374 252 3380 253
rect 3374 248 3375 252
rect 3379 248 3380 252
rect 3374 247 3380 248
rect 3502 252 3508 253
rect 3502 248 3503 252
rect 3507 248 3508 252
rect 3502 247 3508 248
rect 3066 243 3072 244
rect 3066 239 3067 243
rect 3071 239 3072 243
rect 3066 238 3072 239
rect 3146 243 3152 244
rect 3146 239 3147 243
rect 3151 239 3152 243
rect 3146 238 3152 239
rect 3290 243 3296 244
rect 3290 239 3291 243
rect 3295 239 3296 243
rect 3290 238 3296 239
rect 3086 214 3092 215
rect 3086 210 3087 214
rect 3091 210 3092 214
rect 3086 209 3092 210
rect 2962 203 2968 204
rect 2962 199 2963 203
rect 2967 199 2968 203
rect 2962 198 2968 199
rect 3088 187 3090 209
rect 3148 204 3150 238
rect 3230 214 3236 215
rect 3230 210 3231 214
rect 3235 210 3236 214
rect 3230 209 3236 210
rect 3146 203 3152 204
rect 3146 199 3147 203
rect 3151 199 3152 203
rect 3146 198 3152 199
rect 3232 187 3234 209
rect 3292 204 3294 238
rect 3382 214 3388 215
rect 3382 210 3383 214
rect 3387 210 3388 214
rect 3382 209 3388 210
rect 3510 214 3516 215
rect 3510 210 3511 214
rect 3515 210 3516 214
rect 3510 209 3516 210
rect 3290 203 3296 204
rect 3290 199 3291 203
rect 3295 199 3296 203
rect 3290 198 3296 199
rect 3384 187 3386 209
rect 3406 203 3412 204
rect 3406 199 3407 203
rect 3411 199 3412 203
rect 3406 198 3412 199
rect 2655 186 2659 187
rect 2655 181 2659 182
rect 2703 186 2707 187
rect 2703 181 2707 182
rect 2799 186 2803 187
rect 2799 181 2803 182
rect 2815 186 2819 187
rect 2815 181 2819 182
rect 2919 186 2923 187
rect 2919 181 2923 182
rect 2943 186 2947 187
rect 2943 181 2947 182
rect 3015 186 3019 187
rect 3015 181 3019 182
rect 3087 186 3091 187
rect 3087 181 3091 182
rect 3111 186 3115 187
rect 3111 181 3115 182
rect 3207 186 3211 187
rect 3207 181 3211 182
rect 3231 186 3235 187
rect 3231 181 3235 182
rect 3303 186 3307 187
rect 3303 181 3307 182
rect 3383 186 3387 187
rect 3383 181 3387 182
rect 3399 186 3403 187
rect 3399 181 3403 182
rect 2610 179 2616 180
rect 2610 175 2611 179
rect 2615 175 2616 179
rect 2610 174 2616 175
rect 2634 179 2640 180
rect 2634 175 2635 179
rect 2639 175 2640 179
rect 2634 174 2640 175
rect 2471 167 2475 168
rect 2582 170 2588 171
rect 2462 165 2468 166
rect 2472 144 2474 167
rect 2582 166 2583 170
rect 2587 166 2588 170
rect 2582 165 2588 166
rect 2636 144 2638 174
rect 2704 171 2706 181
rect 2754 179 2760 180
rect 2754 175 2755 179
rect 2759 175 2760 179
rect 2754 174 2760 175
rect 2702 170 2708 171
rect 2702 166 2703 170
rect 2707 166 2708 170
rect 2702 165 2708 166
rect 2756 144 2758 174
rect 2816 171 2818 181
rect 2866 179 2872 180
rect 2866 175 2867 179
rect 2871 175 2872 179
rect 2866 174 2872 175
rect 2814 170 2820 171
rect 2814 166 2815 170
rect 2819 166 2820 170
rect 2814 165 2820 166
rect 2868 144 2870 174
rect 2920 171 2922 181
rect 2970 179 2976 180
rect 2970 175 2971 179
rect 2975 175 2976 179
rect 2970 174 2976 175
rect 2918 170 2924 171
rect 2918 166 2919 170
rect 2923 166 2924 170
rect 2918 165 2924 166
rect 2972 144 2974 174
rect 3016 171 3018 181
rect 3066 179 3072 180
rect 3066 175 3067 179
rect 3071 175 3072 179
rect 3066 174 3072 175
rect 3014 170 3020 171
rect 3014 166 3015 170
rect 3019 166 3020 170
rect 3014 165 3020 166
rect 3068 144 3070 174
rect 3112 171 3114 181
rect 3162 179 3168 180
rect 3162 175 3163 179
rect 3167 175 3168 179
rect 3162 174 3168 175
rect 3110 170 3116 171
rect 3110 166 3111 170
rect 3115 166 3116 170
rect 3110 165 3116 166
rect 3164 144 3166 174
rect 3208 171 3210 181
rect 3258 179 3264 180
rect 3258 175 3259 179
rect 3263 175 3264 179
rect 3258 174 3264 175
rect 3206 170 3212 171
rect 3206 166 3207 170
rect 3211 166 3212 170
rect 3206 165 3212 166
rect 3260 144 3262 174
rect 3304 171 3306 181
rect 3354 179 3360 180
rect 3354 175 3355 179
rect 3359 175 3360 179
rect 3354 174 3360 175
rect 3302 170 3308 171
rect 3302 166 3303 170
rect 3307 166 3308 170
rect 3302 165 3308 166
rect 3356 144 3358 174
rect 3400 171 3402 181
rect 3398 170 3404 171
rect 3398 166 3399 170
rect 3403 166 3404 170
rect 3398 165 3404 166
rect 3408 144 3410 198
rect 3512 187 3514 209
rect 3536 204 3538 310
rect 3590 307 3596 308
rect 3590 303 3591 307
rect 3595 303 3596 307
rect 3590 302 3596 303
rect 3592 275 3594 302
rect 3591 274 3595 275
rect 3591 269 3595 270
rect 3592 250 3594 269
rect 3590 249 3596 250
rect 3590 245 3591 249
rect 3595 245 3596 249
rect 3590 244 3596 245
rect 3590 232 3596 233
rect 3590 228 3591 232
rect 3595 228 3596 232
rect 3590 227 3596 228
rect 3534 203 3540 204
rect 3534 199 3535 203
rect 3539 199 3540 203
rect 3534 198 3540 199
rect 3592 187 3594 227
rect 3511 186 3515 187
rect 3511 181 3515 182
rect 3591 186 3595 187
rect 3591 181 3595 182
rect 3592 153 3594 181
rect 3590 152 3596 153
rect 3590 148 3591 152
rect 3595 148 3596 152
rect 3590 147 3596 148
rect 1962 143 1968 144
rect 1962 139 1963 143
rect 1967 139 1968 143
rect 1962 138 1968 139
rect 2094 143 2100 144
rect 2094 139 2095 143
rect 2099 139 2100 143
rect 2094 138 2100 139
rect 2258 143 2264 144
rect 2258 139 2259 143
rect 2263 139 2264 143
rect 2258 138 2264 139
rect 2386 143 2392 144
rect 2386 139 2387 143
rect 2391 139 2392 143
rect 2386 138 2392 139
rect 2470 143 2476 144
rect 2470 139 2471 143
rect 2475 139 2476 143
rect 2470 138 2476 139
rect 2634 143 2640 144
rect 2634 139 2635 143
rect 2639 139 2640 143
rect 2634 138 2640 139
rect 2754 143 2760 144
rect 2754 139 2755 143
rect 2759 139 2760 143
rect 2754 138 2760 139
rect 2866 143 2872 144
rect 2866 139 2867 143
rect 2871 139 2872 143
rect 2866 138 2872 139
rect 2970 143 2976 144
rect 2970 139 2971 143
rect 2975 139 2976 143
rect 2970 138 2976 139
rect 3066 143 3072 144
rect 3066 139 3067 143
rect 3071 139 3072 143
rect 3066 138 3072 139
rect 3162 143 3168 144
rect 3162 139 3163 143
rect 3167 139 3168 143
rect 3162 138 3168 139
rect 3258 143 3264 144
rect 3258 139 3259 143
rect 3263 139 3264 143
rect 3258 138 3264 139
rect 3354 143 3360 144
rect 3354 139 3355 143
rect 3359 139 3360 143
rect 3354 138 3360 139
rect 3406 143 3412 144
rect 3406 139 3407 143
rect 3411 139 3412 143
rect 3406 138 3412 139
rect 1870 135 1876 136
rect 1830 132 1836 133
rect 1830 128 1831 132
rect 1835 128 1836 132
rect 1870 131 1871 135
rect 1875 131 1876 135
rect 3590 135 3596 136
rect 1870 130 1876 131
rect 1894 132 1900 133
rect 1830 127 1836 128
rect 210 123 216 124
rect 210 119 211 123
rect 215 119 216 123
rect 210 118 216 119
rect 290 123 296 124
rect 290 119 291 123
rect 295 119 296 123
rect 290 118 296 119
rect 370 123 376 124
rect 370 119 371 123
rect 375 119 376 123
rect 370 118 376 119
rect 450 123 456 124
rect 450 119 451 123
rect 455 119 456 123
rect 450 118 456 119
rect 530 123 536 124
rect 530 119 531 123
rect 535 119 536 123
rect 530 118 536 119
rect 638 123 644 124
rect 638 119 639 123
rect 643 119 644 123
rect 638 118 644 119
rect 698 123 704 124
rect 698 119 699 123
rect 703 119 704 123
rect 698 118 704 119
rect 786 123 792 124
rect 786 119 787 123
rect 791 119 792 123
rect 786 118 792 119
rect 902 123 908 124
rect 902 119 903 123
rect 907 119 908 123
rect 902 118 908 119
rect 998 123 1004 124
rect 998 119 999 123
rect 1003 119 1004 123
rect 998 118 1004 119
rect 1050 123 1056 124
rect 1050 119 1051 123
rect 1055 119 1056 123
rect 1050 118 1056 119
rect 1158 123 1164 124
rect 1158 119 1159 123
rect 1163 119 1164 123
rect 1158 118 1164 119
rect 1174 123 1180 124
rect 1174 119 1175 123
rect 1179 119 1180 123
rect 1174 118 1180 119
rect 1254 123 1260 124
rect 1254 119 1255 123
rect 1259 119 1260 123
rect 1254 118 1260 119
rect 1342 123 1348 124
rect 1342 119 1343 123
rect 1347 119 1348 123
rect 1342 118 1348 119
rect 1430 123 1436 124
rect 1430 119 1431 123
rect 1435 119 1436 123
rect 1430 118 1436 119
rect 1518 123 1524 124
rect 1518 119 1519 123
rect 1523 119 1524 123
rect 1518 118 1524 119
rect 1598 123 1604 124
rect 1598 119 1599 123
rect 1603 119 1604 123
rect 1598 118 1604 119
rect 1678 123 1684 124
rect 1678 119 1679 123
rect 1683 119 1684 123
rect 1678 118 1684 119
rect 1758 123 1764 124
rect 1758 119 1759 123
rect 1763 119 1764 123
rect 1758 118 1764 119
rect 110 115 116 116
rect 110 111 111 115
rect 115 111 116 115
rect 1830 115 1836 116
rect 110 110 116 111
rect 150 112 156 113
rect 112 91 114 110
rect 150 108 151 112
rect 155 108 156 112
rect 150 107 156 108
rect 230 112 236 113
rect 230 108 231 112
rect 235 108 236 112
rect 230 107 236 108
rect 310 112 316 113
rect 310 108 311 112
rect 315 108 316 112
rect 310 107 316 108
rect 390 112 396 113
rect 390 108 391 112
rect 395 108 396 112
rect 390 107 396 108
rect 470 112 476 113
rect 470 108 471 112
rect 475 108 476 112
rect 470 107 476 108
rect 550 112 556 113
rect 550 108 551 112
rect 555 108 556 112
rect 550 107 556 108
rect 638 112 644 113
rect 638 108 639 112
rect 643 108 644 112
rect 638 107 644 108
rect 726 112 732 113
rect 726 108 727 112
rect 731 108 732 112
rect 726 107 732 108
rect 814 112 820 113
rect 814 108 815 112
rect 819 108 820 112
rect 814 107 820 108
rect 902 112 908 113
rect 902 108 903 112
rect 907 108 908 112
rect 902 107 908 108
rect 990 112 996 113
rect 990 108 991 112
rect 995 108 996 112
rect 990 107 996 108
rect 1078 112 1084 113
rect 1078 108 1079 112
rect 1083 108 1084 112
rect 1078 107 1084 108
rect 1158 112 1164 113
rect 1158 108 1159 112
rect 1163 108 1164 112
rect 1158 107 1164 108
rect 1238 112 1244 113
rect 1238 108 1239 112
rect 1243 108 1244 112
rect 1238 107 1244 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1326 107 1332 108
rect 1414 112 1420 113
rect 1414 108 1415 112
rect 1419 108 1420 112
rect 1414 107 1420 108
rect 1502 112 1508 113
rect 1502 108 1503 112
rect 1507 108 1508 112
rect 1502 107 1508 108
rect 1582 112 1588 113
rect 1582 108 1583 112
rect 1587 108 1588 112
rect 1582 107 1588 108
rect 1662 112 1668 113
rect 1662 108 1663 112
rect 1667 108 1668 112
rect 1662 107 1668 108
rect 1742 112 1748 113
rect 1742 108 1743 112
rect 1747 108 1748 112
rect 1830 111 1831 115
rect 1835 111 1836 115
rect 1872 111 1874 130
rect 1894 128 1895 132
rect 1899 128 1900 132
rect 1894 127 1900 128
rect 1974 132 1980 133
rect 1974 128 1975 132
rect 1979 128 1980 132
rect 1974 127 1980 128
rect 2078 132 2084 133
rect 2078 128 2079 132
rect 2083 128 2084 132
rect 2078 127 2084 128
rect 2198 132 2204 133
rect 2198 128 2199 132
rect 2203 128 2204 132
rect 2198 127 2204 128
rect 2326 132 2332 133
rect 2326 128 2327 132
rect 2331 128 2332 132
rect 2326 127 2332 128
rect 2454 132 2460 133
rect 2454 128 2455 132
rect 2459 128 2460 132
rect 2454 127 2460 128
rect 2574 132 2580 133
rect 2574 128 2575 132
rect 2579 128 2580 132
rect 2574 127 2580 128
rect 2694 132 2700 133
rect 2694 128 2695 132
rect 2699 128 2700 132
rect 2694 127 2700 128
rect 2806 132 2812 133
rect 2806 128 2807 132
rect 2811 128 2812 132
rect 2806 127 2812 128
rect 2910 132 2916 133
rect 2910 128 2911 132
rect 2915 128 2916 132
rect 2910 127 2916 128
rect 3006 132 3012 133
rect 3006 128 3007 132
rect 3011 128 3012 132
rect 3006 127 3012 128
rect 3102 132 3108 133
rect 3102 128 3103 132
rect 3107 128 3108 132
rect 3102 127 3108 128
rect 3198 132 3204 133
rect 3198 128 3199 132
rect 3203 128 3204 132
rect 3198 127 3204 128
rect 3294 132 3300 133
rect 3294 128 3295 132
rect 3299 128 3300 132
rect 3294 127 3300 128
rect 3390 132 3396 133
rect 3390 128 3391 132
rect 3395 128 3396 132
rect 3590 131 3591 135
rect 3595 131 3596 135
rect 3590 130 3596 131
rect 3390 127 3396 128
rect 1896 111 1898 127
rect 1976 111 1978 127
rect 2080 111 2082 127
rect 2200 111 2202 127
rect 2328 111 2330 127
rect 2456 111 2458 127
rect 2576 111 2578 127
rect 2696 111 2698 127
rect 2808 111 2810 127
rect 2912 111 2914 127
rect 3008 111 3010 127
rect 3104 111 3106 127
rect 3200 111 3202 127
rect 3296 111 3298 127
rect 3392 111 3394 127
rect 3592 111 3594 130
rect 1830 110 1836 111
rect 1871 110 1875 111
rect 1742 107 1748 108
rect 152 91 154 107
rect 232 91 234 107
rect 312 91 314 107
rect 392 91 394 107
rect 472 91 474 107
rect 552 91 554 107
rect 640 91 642 107
rect 728 91 730 107
rect 816 91 818 107
rect 904 91 906 107
rect 992 91 994 107
rect 1080 91 1082 107
rect 1160 91 1162 107
rect 1240 91 1242 107
rect 1328 91 1330 107
rect 1416 91 1418 107
rect 1504 91 1506 107
rect 1584 91 1586 107
rect 1664 91 1666 107
rect 1744 91 1746 107
rect 1832 91 1834 110
rect 1871 105 1875 106
rect 1895 110 1899 111
rect 1895 105 1899 106
rect 1975 110 1979 111
rect 1975 105 1979 106
rect 2079 110 2083 111
rect 2079 105 2083 106
rect 2199 110 2203 111
rect 2199 105 2203 106
rect 2327 110 2331 111
rect 2327 105 2331 106
rect 2455 110 2459 111
rect 2455 105 2459 106
rect 2575 110 2579 111
rect 2575 105 2579 106
rect 2695 110 2699 111
rect 2695 105 2699 106
rect 2807 110 2811 111
rect 2807 105 2811 106
rect 2911 110 2915 111
rect 2911 105 2915 106
rect 3007 110 3011 111
rect 3007 105 3011 106
rect 3103 110 3107 111
rect 3103 105 3107 106
rect 3199 110 3203 111
rect 3199 105 3203 106
rect 3295 110 3299 111
rect 3295 105 3299 106
rect 3391 110 3395 111
rect 3391 105 3395 106
rect 3591 110 3595 111
rect 3591 105 3595 106
rect 111 90 115 91
rect 111 85 115 86
rect 151 90 155 91
rect 151 85 155 86
rect 231 90 235 91
rect 231 85 235 86
rect 311 90 315 91
rect 311 85 315 86
rect 391 90 395 91
rect 391 85 395 86
rect 471 90 475 91
rect 471 85 475 86
rect 551 90 555 91
rect 551 85 555 86
rect 639 90 643 91
rect 639 85 643 86
rect 727 90 731 91
rect 727 85 731 86
rect 815 90 819 91
rect 815 85 819 86
rect 903 90 907 91
rect 903 85 907 86
rect 991 90 995 91
rect 991 85 995 86
rect 1079 90 1083 91
rect 1079 85 1083 86
rect 1159 90 1163 91
rect 1159 85 1163 86
rect 1239 90 1243 91
rect 1239 85 1243 86
rect 1327 90 1331 91
rect 1327 85 1331 86
rect 1415 90 1419 91
rect 1415 85 1419 86
rect 1503 90 1507 91
rect 1503 85 1507 86
rect 1583 90 1587 91
rect 1583 85 1587 86
rect 1663 90 1667 91
rect 1663 85 1667 86
rect 1743 90 1747 91
rect 1743 85 1747 86
rect 1831 90 1835 91
rect 1831 85 1835 86
<< m4c >>
rect 1871 3666 1875 3670
rect 2151 3666 2155 3670
rect 2439 3666 2443 3670
rect 2727 3666 2731 3670
rect 3015 3666 3019 3670
rect 3591 3666 3595 3670
rect 111 3638 115 3642
rect 143 3638 147 3642
rect 239 3638 243 3642
rect 367 3638 371 3642
rect 503 3638 507 3642
rect 639 3638 643 3642
rect 775 3638 779 3642
rect 911 3638 915 3642
rect 1055 3638 1059 3642
rect 1199 3638 1203 3642
rect 1831 3638 1835 3642
rect 1871 3590 1875 3594
rect 1903 3590 1907 3594
rect 1983 3590 1987 3594
rect 2071 3590 2075 3594
rect 2159 3590 2163 3594
rect 2175 3590 2179 3594
rect 111 3562 115 3566
rect 135 3562 139 3566
rect 183 3562 187 3566
rect 231 3562 235 3566
rect 303 3562 307 3566
rect 359 3562 363 3566
rect 415 3562 419 3566
rect 111 3478 115 3482
rect 191 3478 195 3482
rect 231 3478 235 3482
rect 311 3478 315 3482
rect 367 3478 371 3482
rect 495 3562 499 3566
rect 527 3562 531 3566
rect 631 3562 635 3566
rect 735 3562 739 3566
rect 767 3562 771 3566
rect 831 3562 835 3566
rect 903 3562 907 3566
rect 919 3562 923 3566
rect 1007 3562 1011 3566
rect 1047 3562 1051 3566
rect 987 3504 991 3508
rect 423 3478 427 3482
rect 503 3478 507 3482
rect 535 3478 539 3482
rect 623 3478 627 3482
rect 639 3478 643 3482
rect 735 3478 739 3482
rect 743 3478 747 3482
rect 839 3478 843 3482
rect 111 3398 115 3402
rect 215 3398 219 3402
rect 223 3398 227 3402
rect 359 3398 363 3402
rect 367 3398 371 3402
rect 495 3398 499 3402
rect 511 3398 515 3402
rect 927 3478 931 3482
rect 943 3478 947 3482
rect 1095 3562 1099 3566
rect 1183 3562 1187 3566
rect 1191 3562 1195 3566
rect 1271 3562 1275 3566
rect 1359 3562 1363 3566
rect 1447 3562 1451 3566
rect 1831 3562 1835 3566
rect 1435 3504 1439 3508
rect 1871 3514 1875 3518
rect 1895 3514 1899 3518
rect 2295 3590 2299 3594
rect 2423 3590 2427 3594
rect 2447 3590 2451 3594
rect 2559 3590 2563 3594
rect 2695 3590 2699 3594
rect 2735 3590 2739 3594
rect 2831 3590 2835 3594
rect 2975 3590 2979 3594
rect 3023 3590 3027 3594
rect 2503 3568 2507 3572
rect 1967 3514 1971 3518
rect 1975 3514 1979 3518
rect 2063 3514 2067 3518
rect 2151 3514 2155 3518
rect 2167 3514 2171 3518
rect 2287 3514 2291 3518
rect 2335 3514 2339 3518
rect 2415 3514 2419 3518
rect 2511 3514 2515 3518
rect 2551 3514 2555 3518
rect 1015 3478 1019 3482
rect 1039 3478 1043 3482
rect 1103 3478 1107 3482
rect 1135 3478 1139 3482
rect 1191 3478 1195 3482
rect 1231 3478 1235 3482
rect 1279 3478 1283 3482
rect 1327 3478 1331 3482
rect 1367 3478 1371 3482
rect 1455 3478 1459 3482
rect 1831 3478 1835 3482
rect 2671 3514 2675 3518
rect 2687 3514 2691 3518
rect 3119 3590 3123 3594
rect 3263 3590 3267 3594
rect 3591 3590 3595 3594
rect 2839 3568 2843 3572
rect 2823 3514 2827 3518
rect 2959 3514 2963 3518
rect 2967 3514 2971 3518
rect 3079 3514 3083 3518
rect 3111 3514 3115 3518
rect 3191 3514 3195 3518
rect 3255 3514 3259 3518
rect 3303 3514 3307 3518
rect 3415 3514 3419 3518
rect 3503 3514 3507 3518
rect 3591 3514 3595 3518
rect 1871 3438 1875 3442
rect 1975 3438 1979 3442
rect 2007 3438 2011 3442
rect 2127 3438 2131 3442
rect 2159 3438 2163 3442
rect 615 3398 619 3402
rect 647 3398 651 3402
rect 727 3398 731 3402
rect 775 3398 779 3402
rect 831 3398 835 3402
rect 895 3398 899 3402
rect 935 3398 939 3402
rect 1015 3398 1019 3402
rect 1031 3398 1035 3402
rect 1127 3398 1131 3402
rect 1223 3398 1227 3402
rect 1239 3398 1243 3402
rect 111 3318 115 3322
rect 207 3318 211 3322
rect 223 3318 227 3322
rect 367 3318 371 3322
rect 375 3318 379 3322
rect 927 3352 931 3356
rect 519 3318 523 3322
rect 655 3318 659 3322
rect 671 3318 675 3322
rect 783 3318 787 3322
rect 815 3318 819 3322
rect 111 3242 115 3246
rect 135 3242 139 3246
rect 199 3242 203 3246
rect 111 3158 115 3162
rect 143 3158 147 3162
rect 175 3158 179 3162
rect 271 3242 275 3246
rect 359 3242 363 3246
rect 415 3242 419 3246
rect 511 3242 515 3246
rect 979 3336 983 3340
rect 903 3318 907 3322
rect 951 3318 955 3322
rect 1319 3398 1323 3402
rect 1351 3398 1355 3402
rect 1831 3398 1835 3402
rect 2255 3438 2259 3442
rect 2343 3438 2347 3442
rect 2391 3438 2395 3442
rect 2519 3438 2523 3442
rect 2535 3438 2539 3442
rect 2679 3438 2683 3442
rect 2831 3438 2835 3442
rect 1247 3352 1251 3356
rect 1871 3362 1875 3366
rect 1999 3362 2003 3366
rect 2015 3362 2019 3366
rect 2119 3362 2123 3366
rect 2151 3362 2155 3366
rect 2247 3362 2251 3366
rect 1327 3336 1331 3340
rect 2967 3438 2971 3442
rect 2999 3438 3003 3442
rect 3087 3438 3091 3442
rect 3167 3438 3171 3442
rect 3199 3438 3203 3442
rect 3311 3438 3315 3442
rect 3343 3438 3347 3442
rect 3423 3438 3427 3442
rect 3511 3438 3515 3442
rect 2295 3362 2299 3366
rect 2383 3362 2387 3366
rect 2439 3362 2443 3366
rect 2527 3362 2531 3366
rect 2583 3362 2587 3366
rect 1023 3318 1027 3322
rect 1087 3318 1091 3322
rect 1135 3318 1139 3322
rect 1215 3318 1219 3322
rect 1247 3318 1251 3322
rect 1343 3318 1347 3322
rect 1359 3318 1363 3322
rect 1471 3318 1475 3322
rect 1831 3318 1835 3322
rect 1871 3286 1875 3290
rect 1927 3286 1931 3290
rect 2023 3286 2027 3290
rect 2063 3286 2067 3290
rect 2159 3286 2163 3290
rect 2191 3286 2195 3290
rect 2303 3286 2307 3290
rect 2319 3286 2323 3290
rect 2447 3286 2451 3290
rect 575 3242 579 3246
rect 663 3242 667 3246
rect 735 3242 739 3246
rect 807 3242 811 3246
rect 895 3242 899 3246
rect 943 3242 947 3246
rect 1047 3242 1051 3246
rect 1079 3242 1083 3246
rect 1191 3242 1195 3246
rect 1207 3242 1211 3246
rect 1327 3242 1331 3246
rect 1335 3242 1339 3246
rect 911 3168 915 3172
rect 279 3158 283 3162
rect 319 3158 323 3162
rect 423 3158 427 3162
rect 463 3158 467 3162
rect 583 3158 587 3162
rect 607 3158 611 3162
rect 743 3158 747 3162
rect 871 3158 875 3162
rect 903 3158 907 3162
rect 111 3070 115 3074
rect 135 3070 139 3074
rect 167 3070 171 3074
rect 223 3070 227 3074
rect 311 3070 315 3074
rect 327 3070 331 3074
rect 111 2982 115 2986
rect 143 2982 147 2986
rect 159 2982 163 2986
rect 439 3070 443 3074
rect 455 3070 459 3074
rect 1079 3176 1083 3180
rect 1463 3242 1467 3246
rect 1607 3242 1611 3246
rect 1831 3242 1835 3246
rect 1871 3210 1875 3214
rect 1399 3176 1403 3180
rect 1895 3210 1899 3214
rect 1919 3210 1923 3214
rect 2007 3210 2011 3214
rect 2055 3210 2059 3214
rect 2143 3210 2147 3214
rect 2183 3210 2187 3214
rect 1587 3192 1591 3196
rect 2671 3362 2675 3366
rect 2727 3362 2731 3366
rect 2823 3362 2827 3366
rect 2871 3362 2875 3366
rect 2991 3362 2995 3366
rect 3023 3362 3027 3366
rect 3159 3362 3163 3366
rect 3183 3362 3187 3366
rect 3335 3362 3339 3366
rect 3351 3362 3355 3366
rect 3591 3438 3595 3442
rect 3503 3362 3507 3366
rect 2591 3286 2595 3290
rect 2735 3286 2739 3290
rect 3591 3362 3595 3366
rect 2743 3286 2747 3290
rect 2295 3210 2299 3214
rect 2311 3210 2315 3214
rect 991 3158 995 3162
rect 1055 3158 1059 3162
rect 1103 3158 1107 3162
rect 1199 3158 1203 3162
rect 1207 3158 1211 3162
rect 1311 3158 1315 3162
rect 1335 3158 1339 3162
rect 1407 3158 1411 3162
rect 1471 3158 1475 3162
rect 1495 3158 1499 3162
rect 1583 3158 1587 3162
rect 1615 3158 1619 3162
rect 1671 3158 1675 3162
rect 1751 3158 1755 3162
rect 1831 3158 1835 3162
rect 1871 3134 1875 3138
rect 2439 3210 2443 3214
rect 2455 3210 2459 3214
rect 2583 3210 2587 3214
rect 2879 3286 2883 3290
rect 2919 3286 2923 3290
rect 3031 3286 3035 3290
rect 3111 3286 3115 3290
rect 3191 3286 3195 3290
rect 3311 3286 3315 3290
rect 3359 3286 3363 3290
rect 3511 3286 3515 3290
rect 2787 3264 2791 3268
rect 3591 3286 3595 3290
rect 3319 3264 3323 3268
rect 2623 3210 2627 3214
rect 2735 3210 2739 3214
rect 2799 3210 2803 3214
rect 2911 3210 2915 3214
rect 2975 3210 2979 3214
rect 3103 3210 3107 3214
rect 3151 3210 3155 3214
rect 3303 3210 3307 3214
rect 3327 3210 3331 3214
rect 3503 3210 3507 3214
rect 1903 3134 1907 3138
rect 2015 3134 2019 3138
rect 2071 3134 2075 3138
rect 2151 3134 2155 3138
rect 2263 3134 2267 3138
rect 2303 3134 2307 3138
rect 2455 3134 2459 3138
rect 2463 3134 2467 3138
rect 551 3070 555 3074
rect 599 3070 603 3074
rect 663 3070 667 3074
rect 735 3070 739 3074
rect 863 3070 867 3074
rect 983 3070 987 3074
rect 1095 3070 1099 3074
rect 1199 3070 1203 3074
rect 1303 3070 1307 3074
rect 1399 3070 1403 3074
rect 1487 3070 1491 3074
rect 1575 3070 1579 3074
rect 1663 3070 1667 3074
rect 1743 3070 1747 3074
rect 1831 3070 1835 3074
rect 2631 3134 2635 3138
rect 2647 3134 2651 3138
rect 2807 3134 2811 3138
rect 2831 3134 2835 3138
rect 2983 3134 2987 3138
rect 1871 3046 1875 3050
rect 1895 3046 1899 3050
rect 2063 3046 2067 3050
rect 2199 3046 2203 3050
rect 2255 3046 2259 3050
rect 231 2982 235 2986
rect 319 2982 323 2986
rect 335 2982 339 2986
rect 447 2982 451 2986
rect 487 2982 491 2986
rect 559 2982 563 2986
rect 647 2982 651 2986
rect 671 2982 675 2986
rect 799 2982 803 2986
rect 111 2906 115 2910
rect 151 2906 155 2910
rect 311 2906 315 2910
rect 111 2826 115 2830
rect 143 2826 147 2830
rect 471 2906 475 2910
rect 479 2906 483 2910
rect 943 2982 947 2986
rect 1079 2982 1083 2986
rect 1199 2982 1203 2986
rect 1311 2982 1315 2986
rect 631 2906 635 2910
rect 639 2906 643 2910
rect 783 2906 787 2910
rect 791 2906 795 2910
rect 927 2906 931 2910
rect 935 2906 939 2910
rect 1055 2906 1059 2910
rect 1071 2906 1075 2910
rect 1175 2906 1179 2910
rect 1191 2906 1195 2910
rect 1423 2982 1427 2986
rect 1535 2982 1539 2986
rect 1647 2982 1651 2986
rect 1831 2982 1835 2986
rect 1871 2958 1875 2962
rect 2127 2958 2131 2962
rect 2207 2958 2211 2962
rect 2335 3046 2339 3050
rect 2447 3046 2451 3050
rect 2479 3046 2483 3050
rect 2623 3046 2627 3050
rect 2639 3046 2643 3050
rect 3015 3134 3019 3138
rect 3159 3134 3163 3138
rect 3199 3134 3203 3138
rect 3335 3134 3339 3138
rect 3391 3134 3395 3138
rect 3591 3210 3595 3214
rect 3511 3134 3515 3138
rect 3591 3134 3595 3138
rect 2767 3046 2771 3050
rect 2823 3046 2827 3050
rect 2903 3046 2907 3050
rect 3007 3046 3011 3050
rect 3039 3046 3043 3050
rect 3183 3046 3187 3050
rect 3191 3046 3195 3050
rect 2287 2958 2291 2962
rect 2343 2958 2347 2962
rect 2367 2958 2371 2962
rect 2447 2958 2451 2962
rect 2487 2958 2491 2962
rect 2527 2958 2531 2962
rect 2607 2958 2611 2962
rect 2631 2958 2635 2962
rect 2695 2958 2699 2962
rect 2775 2958 2779 2962
rect 2791 2958 2795 2962
rect 2911 2958 2915 2962
rect 3039 2958 3043 2962
rect 3047 2958 3051 2962
rect 1287 2906 1291 2910
rect 1303 2906 1307 2910
rect 1391 2906 1395 2910
rect 1415 2906 1419 2910
rect 159 2826 163 2830
rect 247 2826 251 2830
rect 319 2826 323 2830
rect 383 2826 387 2830
rect 479 2826 483 2830
rect 535 2826 539 2830
rect 639 2826 643 2830
rect 687 2826 691 2830
rect 791 2826 795 2830
rect 847 2826 851 2830
rect 111 2746 115 2750
rect 135 2746 139 2750
rect 231 2746 235 2750
rect 239 2746 243 2750
rect 367 2746 371 2750
rect 375 2746 379 2750
rect 111 2662 115 2666
rect 143 2662 147 2666
rect 511 2746 515 2750
rect 527 2746 531 2750
rect 935 2826 939 2830
rect 999 2826 1003 2830
rect 1487 2906 1491 2910
rect 1527 2906 1531 2910
rect 1591 2906 1595 2910
rect 1639 2906 1643 2910
rect 1695 2906 1699 2910
rect 1831 2906 1835 2910
rect 1871 2882 1875 2886
rect 2047 2882 2051 2886
rect 1435 2848 1439 2852
rect 1063 2826 1067 2830
rect 1143 2826 1147 2830
rect 1183 2826 1187 2830
rect 1279 2826 1283 2830
rect 1295 2826 1299 2830
rect 663 2746 667 2750
rect 679 2746 683 2750
rect 815 2746 819 2750
rect 839 2746 843 2750
rect 975 2746 979 2750
rect 991 2746 995 2750
rect 1135 2746 1139 2750
rect 1399 2826 1403 2830
rect 1407 2826 1411 2830
rect 1675 2848 1679 2852
rect 1495 2826 1499 2830
rect 1527 2826 1531 2830
rect 1599 2826 1603 2830
rect 1647 2826 1651 2830
rect 1703 2826 1707 2830
rect 1751 2826 1755 2830
rect 1831 2826 1835 2830
rect 2119 2882 2123 2886
rect 2135 2882 2139 2886
rect 2199 2882 2203 2886
rect 2239 2882 2243 2886
rect 2279 2882 2283 2886
rect 1871 2794 1875 2798
rect 1903 2794 1907 2798
rect 2015 2794 2019 2798
rect 2055 2794 2059 2798
rect 1271 2746 1275 2750
rect 1287 2746 1291 2750
rect 1399 2746 1403 2750
rect 1447 2746 1451 2750
rect 1519 2746 1523 2750
rect 1607 2746 1611 2750
rect 1639 2746 1643 2750
rect 239 2662 243 2666
rect 279 2662 283 2666
rect 375 2662 379 2666
rect 447 2662 451 2666
rect 519 2662 523 2666
rect 623 2662 627 2666
rect 671 2662 675 2666
rect 791 2662 795 2666
rect 823 2662 827 2666
rect 111 2582 115 2586
rect 135 2582 139 2586
rect 223 2582 227 2586
rect 271 2582 275 2586
rect 367 2582 371 2586
rect 111 2502 115 2506
rect 143 2502 147 2506
rect 439 2582 443 2586
rect 527 2582 531 2586
rect 1007 2680 1011 2684
rect 1223 2680 1227 2684
rect 951 2662 955 2666
rect 983 2662 987 2666
rect 1103 2662 1107 2666
rect 1143 2662 1147 2666
rect 1247 2662 1251 2666
rect 1295 2662 1299 2666
rect 1399 2662 1403 2666
rect 1455 2662 1459 2666
rect 1551 2662 1555 2666
rect 615 2582 619 2586
rect 703 2582 707 2586
rect 783 2582 787 2586
rect 879 2582 883 2586
rect 943 2582 947 2586
rect 1743 2746 1747 2750
rect 1831 2746 1835 2750
rect 1871 2718 1875 2722
rect 1895 2718 1899 2722
rect 2007 2718 2011 2722
rect 1615 2662 1619 2666
rect 1751 2662 1755 2666
rect 1831 2662 1835 2666
rect 2143 2794 2147 2798
rect 2167 2794 2171 2798
rect 2343 2882 2347 2886
rect 2359 2882 2363 2886
rect 2439 2882 2443 2886
rect 2463 2882 2467 2886
rect 2519 2882 2523 2886
rect 2591 2882 2595 2886
rect 2599 2882 2603 2886
rect 2247 2794 2251 2798
rect 2327 2794 2331 2798
rect 2351 2794 2355 2798
rect 2471 2794 2475 2798
rect 2487 2794 2491 2798
rect 2067 2776 2071 2780
rect 2419 2776 2423 2780
rect 2687 2882 2691 2886
rect 2727 2882 2731 2886
rect 2783 2882 2787 2886
rect 2879 2882 2883 2886
rect 2903 2882 2907 2886
rect 3327 3046 3331 3050
rect 3383 3046 3387 3050
rect 3591 3046 3595 3050
rect 3183 2958 3187 2962
rect 3191 2958 3195 2962
rect 3335 2958 3339 2962
rect 3495 2958 3499 2962
rect 3591 2958 3595 2962
rect 3031 2882 3035 2886
rect 3175 2882 3179 2886
rect 3191 2882 3195 2886
rect 2667 2816 2671 2820
rect 2599 2794 2603 2798
rect 2639 2794 2643 2798
rect 2959 2816 2963 2820
rect 3327 2882 3331 2886
rect 3359 2882 3363 2886
rect 3487 2882 3491 2886
rect 3503 2882 3507 2886
rect 2735 2794 2739 2798
rect 2791 2794 2795 2798
rect 2887 2794 2891 2798
rect 2943 2794 2947 2798
rect 3039 2794 3043 2798
rect 3087 2794 3091 2798
rect 3199 2794 3203 2798
rect 3231 2794 3235 2798
rect 3367 2794 3371 2798
rect 3383 2794 3387 2798
rect 3591 2882 3595 2886
rect 3511 2794 3515 2798
rect 2103 2718 2107 2722
rect 2159 2718 2163 2722
rect 2319 2718 2323 2722
rect 2327 2718 2331 2722
rect 1931 2656 1935 2660
rect 1871 2634 1875 2638
rect 1903 2634 1907 2638
rect 2479 2718 2483 2722
rect 2535 2718 2539 2722
rect 2631 2718 2635 2722
rect 2735 2718 2739 2722
rect 2783 2718 2787 2722
rect 2911 2718 2915 2722
rect 2935 2718 2939 2722
rect 3071 2718 3075 2722
rect 3079 2718 3083 2722
rect 2479 2656 2483 2660
rect 2771 2656 2775 2660
rect 3223 2718 3227 2722
rect 3375 2718 3379 2722
rect 3591 2794 3595 2798
rect 3503 2718 3507 2722
rect 3139 2656 3143 2660
rect 3591 2718 3595 2722
rect 2055 2634 2059 2638
rect 2111 2634 2115 2638
rect 2263 2634 2267 2638
rect 2335 2634 2339 2638
rect 2495 2634 2499 2638
rect 2543 2634 2547 2638
rect 2743 2634 2747 2638
rect 2751 2634 2755 2638
rect 2919 2634 2923 2638
rect 3015 2634 3019 2638
rect 3079 2634 3083 2638
rect 3231 2634 3235 2638
rect 3287 2634 3291 2638
rect 3383 2634 3387 2638
rect 3511 2634 3515 2638
rect 1047 2582 1051 2586
rect 1095 2582 1099 2586
rect 1207 2582 1211 2586
rect 1239 2582 1243 2586
rect 1359 2582 1363 2586
rect 1391 2582 1395 2586
rect 1511 2582 1515 2586
rect 1543 2582 1547 2586
rect 1671 2582 1675 2586
rect 1831 2582 1835 2586
rect 1871 2558 1875 2562
rect 1895 2558 1899 2562
rect 2007 2558 2011 2562
rect 2047 2558 2051 2562
rect 2159 2558 2163 2562
rect 2255 2558 2259 2562
rect 2319 2558 2323 2562
rect 2471 2558 2475 2562
rect 2487 2558 2491 2562
rect 2623 2558 2627 2562
rect 223 2502 227 2506
rect 231 2502 235 2506
rect 303 2502 307 2506
rect 375 2502 379 2506
rect 391 2502 395 2506
rect 511 2502 515 2506
rect 535 2502 539 2506
rect 647 2502 651 2506
rect 711 2502 715 2506
rect 783 2502 787 2506
rect 887 2502 891 2506
rect 927 2502 931 2506
rect 1055 2502 1059 2506
rect 1063 2502 1067 2506
rect 1191 2502 1195 2506
rect 1215 2502 1219 2506
rect 1311 2502 1315 2506
rect 1367 2502 1371 2506
rect 1431 2502 1435 2506
rect 1519 2502 1523 2506
rect 1551 2502 1555 2506
rect 1671 2502 1675 2506
rect 1679 2502 1683 2506
rect 2743 2558 2747 2562
rect 2759 2558 2763 2562
rect 2887 2558 2891 2562
rect 3007 2558 3011 2562
rect 1931 2528 1935 2532
rect 1831 2502 1835 2506
rect 2659 2528 2663 2532
rect 3119 2558 3123 2562
rect 3223 2558 3227 2562
rect 3279 2558 3283 2562
rect 1871 2474 1875 2478
rect 1903 2474 1907 2478
rect 1999 2474 2003 2478
rect 2015 2474 2019 2478
rect 2127 2474 2131 2478
rect 2167 2474 2171 2478
rect 2263 2474 2267 2478
rect 2327 2474 2331 2478
rect 2407 2474 2411 2478
rect 2479 2474 2483 2478
rect 2551 2474 2555 2478
rect 2631 2474 2635 2478
rect 2703 2474 2707 2478
rect 2767 2474 2771 2478
rect 2863 2474 2867 2478
rect 2895 2474 2899 2478
rect 3015 2474 3019 2478
rect 3023 2474 3027 2478
rect 1135 2456 1139 2460
rect 1471 2456 1475 2460
rect 111 2414 115 2418
rect 135 2414 139 2418
rect 215 2414 219 2418
rect 295 2414 299 2418
rect 383 2414 387 2418
rect 503 2414 507 2418
rect 639 2414 643 2418
rect 775 2414 779 2418
rect 919 2414 923 2418
rect 1055 2414 1059 2418
rect 1063 2414 1067 2418
rect 1143 2414 1147 2418
rect 1183 2414 1187 2418
rect 1223 2414 1227 2418
rect 1303 2414 1307 2418
rect 1383 2414 1387 2418
rect 1423 2414 1427 2418
rect 1463 2414 1467 2418
rect 2803 2456 2807 2460
rect 3319 2558 3323 2562
rect 3423 2558 3427 2562
rect 3503 2558 3507 2562
rect 3127 2474 3131 2478
rect 3191 2474 3195 2478
rect 3231 2474 3235 2478
rect 3327 2474 3331 2478
rect 3359 2474 3363 2478
rect 3199 2456 3203 2460
rect 3431 2474 3435 2478
rect 3511 2474 3515 2478
rect 1543 2414 1547 2418
rect 1663 2414 1667 2418
rect 1831 2414 1835 2418
rect 1871 2394 1875 2398
rect 1991 2394 1995 2398
rect 2119 2394 2123 2398
rect 2143 2394 2147 2398
rect 2239 2394 2243 2398
rect 2255 2394 2259 2398
rect 2343 2394 2347 2398
rect 2399 2394 2403 2398
rect 2455 2394 2459 2398
rect 111 2330 115 2334
rect 359 2330 363 2334
rect 439 2330 443 2334
rect 519 2330 523 2334
rect 599 2330 603 2334
rect 679 2330 683 2334
rect 759 2330 763 2334
rect 839 2330 843 2334
rect 919 2330 923 2334
rect 999 2330 1003 2334
rect 111 2254 115 2258
rect 351 2254 355 2258
rect 375 2254 379 2258
rect 431 2254 435 2258
rect 455 2254 459 2258
rect 511 2254 515 2258
rect 535 2254 539 2258
rect 591 2254 595 2258
rect 615 2254 619 2258
rect 671 2254 675 2258
rect 695 2254 699 2258
rect 751 2254 755 2258
rect 775 2254 779 2258
rect 831 2254 835 2258
rect 855 2254 859 2258
rect 1071 2330 1075 2334
rect 1079 2330 1083 2334
rect 1151 2330 1155 2334
rect 1159 2330 1163 2334
rect 1231 2330 1235 2334
rect 1239 2330 1243 2334
rect 1311 2330 1315 2334
rect 1319 2330 1323 2334
rect 1391 2330 1395 2334
rect 1471 2330 1475 2334
rect 1831 2330 1835 2334
rect 2179 2328 2183 2332
rect 1871 2314 1875 2318
rect 2151 2314 2155 2318
rect 2247 2314 2251 2318
rect 2279 2314 2283 2318
rect 2543 2394 2547 2398
rect 2575 2394 2579 2398
rect 2695 2394 2699 2398
rect 2703 2394 2707 2398
rect 2847 2394 2851 2398
rect 2855 2394 2859 2398
rect 2479 2328 2483 2332
rect 2883 2328 2887 2332
rect 3007 2394 3011 2398
rect 3015 2394 3019 2398
rect 3175 2394 3179 2398
rect 3183 2394 3187 2398
rect 3351 2394 3355 2398
rect 3591 2634 3595 2638
rect 3591 2558 3595 2562
rect 3591 2474 3595 2478
rect 3503 2394 3507 2398
rect 3123 2328 3127 2332
rect 2351 2314 2355 2318
rect 2359 2314 2363 2318
rect 2439 2314 2443 2318
rect 2463 2314 2467 2318
rect 2519 2314 2523 2318
rect 2583 2314 2587 2318
rect 2599 2314 2603 2318
rect 2679 2314 2683 2318
rect 2711 2314 2715 2318
rect 2759 2314 2763 2318
rect 2847 2314 2851 2318
rect 2855 2314 2859 2318
rect 2935 2314 2939 2318
rect 3015 2314 3019 2318
rect 3183 2314 3187 2318
rect 3359 2314 3363 2318
rect 911 2254 915 2258
rect 935 2254 939 2258
rect 991 2254 995 2258
rect 1015 2254 1019 2258
rect 1071 2254 1075 2258
rect 1095 2254 1099 2258
rect 1151 2254 1155 2258
rect 1175 2254 1179 2258
rect 1231 2254 1235 2258
rect 1255 2254 1259 2258
rect 1311 2254 1315 2258
rect 1831 2254 1835 2258
rect 1871 2238 1875 2242
rect 2271 2238 2275 2242
rect 2311 2238 2315 2242
rect 2351 2238 2355 2242
rect 111 2166 115 2170
rect 311 2166 315 2170
rect 383 2166 387 2170
rect 407 2166 411 2170
rect 463 2166 467 2170
rect 503 2166 507 2170
rect 543 2166 547 2170
rect 599 2166 603 2170
rect 623 2166 627 2170
rect 687 2166 691 2170
rect 703 2166 707 2170
rect 111 2078 115 2082
rect 207 2078 211 2082
rect 303 2078 307 2082
rect 327 2078 331 2082
rect 399 2078 403 2082
rect 447 2078 451 2082
rect 495 2078 499 2082
rect 575 2078 579 2082
rect 591 2078 595 2082
rect 111 1998 115 2002
rect 191 1998 195 2002
rect 215 1998 219 2002
rect 335 1998 339 2002
rect 351 1998 355 2002
rect 775 2166 779 2170
rect 783 2166 787 2170
rect 863 2166 867 2170
rect 943 2166 947 2170
rect 951 2166 955 2170
rect 1023 2166 1027 2170
rect 1039 2166 1043 2170
rect 1103 2166 1107 2170
rect 1127 2166 1131 2170
rect 1183 2166 1187 2170
rect 1223 2166 1227 2170
rect 1263 2166 1267 2170
rect 1831 2166 1835 2170
rect 679 2078 683 2082
rect 703 2078 707 2082
rect 767 2078 771 2082
rect 823 2078 827 2082
rect 855 2078 859 2082
rect 943 2078 947 2082
rect 1031 2078 1035 2082
rect 1063 2078 1067 2082
rect 1119 2078 1123 2082
rect 1175 2078 1179 2082
rect 1215 2078 1219 2082
rect 2399 2238 2403 2242
rect 2431 2238 2435 2242
rect 2495 2238 2499 2242
rect 2511 2238 2515 2242
rect 2591 2238 2595 2242
rect 2599 2238 2603 2242
rect 1871 2158 1875 2162
rect 1903 2158 1907 2162
rect 1983 2158 1987 2162
rect 2111 2158 2115 2162
rect 2247 2158 2251 2162
rect 2319 2158 2323 2162
rect 2391 2158 2395 2162
rect 2407 2158 2411 2162
rect 1279 2078 1283 2082
rect 1375 2078 1379 2082
rect 1471 2078 1475 2082
rect 1567 2078 1571 2082
rect 1663 2078 1667 2082
rect 1743 2078 1747 2082
rect 455 1998 459 2002
rect 519 1998 523 2002
rect 583 1998 587 2002
rect 687 1998 691 2002
rect 711 1998 715 2002
rect 831 1998 835 2002
rect 855 1998 859 2002
rect 111 1918 115 1922
rect 135 1918 139 1922
rect 183 1918 187 1922
rect 239 1918 243 1922
rect 343 1918 347 1922
rect 375 1918 379 1922
rect 511 1918 515 1922
rect 527 1918 531 1922
rect 951 1998 955 2002
rect 1015 1998 1019 2002
rect 1071 1998 1075 2002
rect 1167 1998 1171 2002
rect 1183 1998 1187 2002
rect 1287 1998 1291 2002
rect 1311 1998 1315 2002
rect 679 1918 683 1922
rect 687 1918 691 1922
rect 847 1918 851 1922
rect 1007 1918 1011 1922
rect 1159 1918 1163 1922
rect 111 1838 115 1842
rect 143 1838 147 1842
rect 247 1838 251 1842
rect 287 1838 291 1842
rect 383 1838 387 1842
rect 471 1838 475 1842
rect 535 1838 539 1842
rect 663 1838 667 1842
rect 695 1838 699 1842
rect 847 1838 851 1842
rect 855 1838 859 1842
rect 111 1754 115 1758
rect 135 1754 139 1758
rect 215 1754 219 1758
rect 279 1754 283 1758
rect 343 1754 347 1758
rect 463 1754 467 1758
rect 1831 2078 1835 2082
rect 1871 2074 1875 2078
rect 1895 2074 1899 2078
rect 1967 2074 1971 2078
rect 1975 2074 1979 2078
rect 2503 2158 2507 2162
rect 2543 2158 2547 2162
rect 2671 2238 2675 2242
rect 2719 2238 2723 2242
rect 2751 2238 2755 2242
rect 2839 2238 2843 2242
rect 2855 2238 2859 2242
rect 2927 2238 2931 2242
rect 3007 2238 3011 2242
rect 3175 2238 3179 2242
rect 3351 2238 3355 2242
rect 3591 2394 3595 2398
rect 3511 2314 3515 2318
rect 3503 2238 3507 2242
rect 2735 2176 2739 2180
rect 2607 2158 2611 2162
rect 2695 2158 2699 2162
rect 2727 2158 2731 2162
rect 3083 2176 3087 2180
rect 2847 2158 2851 2162
rect 2863 2158 2867 2162
rect 3007 2158 3011 2162
rect 3015 2158 3019 2162
rect 3175 2158 3179 2162
rect 3183 2158 3187 2162
rect 3351 2158 3355 2162
rect 3359 2158 3363 2162
rect 2103 2074 2107 2078
rect 2215 2074 2219 2078
rect 2239 2074 2243 2078
rect 2383 2074 2387 2078
rect 2447 2074 2451 2078
rect 1383 1998 1387 2002
rect 1447 1998 1451 2002
rect 1479 1998 1483 2002
rect 1575 1998 1579 2002
rect 1583 1998 1587 2002
rect 1671 1998 1675 2002
rect 1719 1998 1723 2002
rect 1751 1998 1755 2002
rect 1831 1998 1835 2002
rect 1871 1998 1875 2002
rect 1959 1998 1963 2002
rect 1975 1998 1979 2002
rect 2079 1998 2083 2002
rect 2199 1998 2203 2002
rect 2223 1998 2227 2002
rect 2535 2074 2539 2078
rect 2655 2074 2659 2078
rect 2687 2074 2691 2078
rect 2839 2074 2843 2078
rect 2999 2074 3003 2078
rect 3143 2074 3147 2078
rect 3167 2074 3171 2078
rect 3271 2074 3275 2078
rect 2687 2008 2691 2012
rect 2319 1998 2323 2002
rect 2447 1998 2451 2002
rect 2455 1998 2459 2002
rect 2583 1998 2587 2002
rect 2663 1998 2667 2002
rect 2743 1998 2747 2002
rect 2847 1998 2851 2002
rect 2919 1998 2923 2002
rect 3007 1998 3011 2002
rect 1303 1918 1307 1922
rect 1439 1918 1443 1922
rect 1455 1918 1459 1922
rect 1575 1918 1579 1922
rect 1607 1918 1611 1922
rect 1711 1918 1715 1922
rect 1015 1838 1019 1842
rect 1023 1838 1027 1842
rect 1167 1838 1171 1842
rect 1191 1838 1195 1842
rect 495 1754 499 1758
rect 655 1754 659 1758
rect 663 1754 667 1758
rect 839 1754 843 1758
rect 1007 1754 1011 1758
rect 1015 1754 1019 1758
rect 1831 1918 1835 1922
rect 1871 1914 1875 1918
rect 1951 1914 1955 1918
rect 2063 1914 2067 1918
rect 2071 1914 2075 1918
rect 2151 1914 2155 1918
rect 2191 1914 2195 1918
rect 3087 2008 3091 2012
rect 3343 2074 3347 2078
rect 3511 2158 3515 2162
rect 3591 2314 3595 2318
rect 3591 2238 3595 2242
rect 3591 2158 3595 2162
rect 3399 2074 3403 2078
rect 3503 2074 3507 2078
rect 3591 2074 3595 2078
rect 3119 1998 3123 2002
rect 3151 1998 3155 2002
rect 3279 1998 3283 2002
rect 3327 1998 3331 2002
rect 3407 1998 3411 2002
rect 2239 1914 2243 1918
rect 1311 1838 1315 1842
rect 1351 1838 1355 1842
rect 1463 1838 1467 1842
rect 1511 1838 1515 1842
rect 1615 1838 1619 1842
rect 1679 1838 1683 1842
rect 1831 1838 1835 1842
rect 1871 1822 1875 1826
rect 2071 1822 2075 1826
rect 2095 1822 2099 1826
rect 1167 1754 1171 1758
rect 1183 1754 1187 1758
rect 1319 1754 1323 1758
rect 1343 1754 1347 1758
rect 111 1674 115 1678
rect 143 1674 147 1678
rect 223 1674 227 1678
rect 295 1674 299 1678
rect 351 1674 355 1678
rect 479 1674 483 1678
rect 503 1674 507 1678
rect 671 1674 675 1678
rect 847 1674 851 1678
rect 855 1674 859 1678
rect 1015 1674 1019 1678
rect 1031 1674 1035 1678
rect 111 1598 115 1602
rect 135 1598 139 1602
rect 159 1598 163 1602
rect 287 1598 291 1602
rect 423 1598 427 1602
rect 471 1598 475 1602
rect 567 1598 571 1602
rect 663 1598 667 1602
rect 711 1598 715 1602
rect 847 1598 851 1602
rect 2311 1914 2315 1918
rect 2319 1914 2323 1918
rect 2399 1914 2403 1918
rect 2439 1914 2443 1918
rect 2487 1914 2491 1918
rect 2575 1914 2579 1918
rect 2663 1914 2667 1918
rect 2735 1914 2739 1918
rect 2759 1914 2763 1918
rect 2871 1914 2875 1918
rect 2911 1914 2915 1918
rect 2991 1914 2995 1918
rect 3111 1914 3115 1918
rect 3119 1914 3123 1918
rect 3247 1914 3251 1918
rect 3319 1914 3323 1918
rect 3383 1914 3387 1918
rect 3511 1998 3515 2002
rect 3591 1998 3595 2002
rect 3503 1914 3507 1918
rect 2159 1822 2163 1826
rect 2239 1822 2243 1826
rect 2247 1822 2251 1826
rect 2327 1822 2331 1826
rect 2399 1822 2403 1826
rect 2407 1822 2411 1826
rect 2495 1822 2499 1826
rect 2559 1822 2563 1826
rect 2583 1822 2587 1826
rect 2671 1822 2675 1826
rect 2719 1822 2723 1826
rect 2767 1822 2771 1826
rect 2879 1822 2883 1826
rect 2999 1822 3003 1826
rect 3031 1822 3035 1826
rect 3127 1822 3131 1826
rect 3175 1822 3179 1826
rect 1463 1754 1467 1758
rect 1503 1754 1507 1758
rect 1607 1754 1611 1758
rect 1671 1754 1675 1758
rect 1743 1754 1747 1758
rect 1831 1754 1835 1758
rect 1871 1742 1875 1746
rect 2087 1742 2091 1746
rect 2103 1742 2107 1746
rect 2231 1742 2235 1746
rect 2239 1742 2243 1746
rect 2383 1742 2387 1746
rect 2391 1742 2395 1746
rect 1175 1674 1179 1678
rect 1199 1674 1203 1678
rect 1327 1674 1331 1678
rect 1359 1674 1363 1678
rect 1471 1674 1475 1678
rect 1519 1674 1523 1678
rect 1615 1674 1619 1678
rect 1679 1674 1683 1678
rect 983 1598 987 1602
rect 1023 1598 1027 1602
rect 2527 1742 2531 1746
rect 2551 1742 2555 1746
rect 2663 1742 2667 1746
rect 1751 1674 1755 1678
rect 1831 1674 1835 1678
rect 1871 1662 1875 1666
rect 1967 1662 1971 1666
rect 2087 1662 2091 1666
rect 2111 1662 2115 1666
rect 2215 1662 2219 1666
rect 2247 1662 2251 1666
rect 2351 1662 2355 1666
rect 2391 1662 2395 1666
rect 1119 1598 1123 1602
rect 1191 1598 1195 1602
rect 1247 1598 1251 1602
rect 111 1518 115 1522
rect 167 1518 171 1522
rect 231 1518 235 1522
rect 295 1518 299 1522
rect 375 1518 379 1522
rect 431 1518 435 1522
rect 519 1518 523 1522
rect 575 1518 579 1522
rect 655 1518 659 1522
rect 719 1518 723 1522
rect 783 1518 787 1522
rect 855 1518 859 1522
rect 111 1434 115 1438
rect 223 1434 227 1438
rect 255 1434 259 1438
rect 351 1434 355 1438
rect 367 1434 371 1438
rect 111 1358 115 1362
rect 263 1358 267 1362
rect 447 1434 451 1438
rect 511 1434 515 1438
rect 543 1434 547 1438
rect 631 1434 635 1438
rect 647 1434 651 1438
rect 903 1518 907 1522
rect 991 1518 995 1522
rect 1015 1518 1019 1522
rect 719 1434 723 1438
rect 775 1434 779 1438
rect 807 1434 811 1438
rect 895 1434 899 1438
rect 919 1434 923 1438
rect 1351 1598 1355 1602
rect 1375 1598 1379 1602
rect 1511 1598 1515 1602
rect 1671 1598 1675 1602
rect 1831 1598 1835 1602
rect 1871 1578 1875 1582
rect 1895 1578 1899 1582
rect 1959 1578 1963 1582
rect 1119 1518 1123 1522
rect 1127 1518 1131 1522
rect 1215 1518 1219 1522
rect 1255 1518 1259 1522
rect 1319 1518 1323 1522
rect 1383 1518 1387 1522
rect 1423 1518 1427 1522
rect 1155 1496 1159 1500
rect 1519 1518 1523 1522
rect 1831 1518 1835 1522
rect 1431 1504 1435 1508
rect 2495 1662 2499 1666
rect 2535 1662 2539 1666
rect 2639 1662 2643 1666
rect 2711 1742 2715 1746
rect 2799 1742 2803 1746
rect 2871 1742 2875 1746
rect 2927 1742 2931 1746
rect 3023 1742 3027 1746
rect 3047 1742 3051 1746
rect 3591 1914 3595 1918
rect 3255 1822 3259 1826
rect 3319 1822 3323 1826
rect 3391 1822 3395 1826
rect 3471 1822 3475 1826
rect 3511 1822 3515 1826
rect 3591 1822 3595 1826
rect 3159 1742 3163 1746
rect 3167 1742 3171 1746
rect 3271 1742 3275 1746
rect 3311 1742 3315 1746
rect 3391 1742 3395 1746
rect 2671 1662 2675 1666
rect 2783 1662 2787 1666
rect 2807 1662 2811 1666
rect 2927 1662 2931 1666
rect 2935 1662 2939 1666
rect 3055 1662 3059 1666
rect 3071 1662 3075 1666
rect 3167 1662 3171 1666
rect 3223 1662 3227 1666
rect 3279 1662 3283 1666
rect 3375 1662 3379 1666
rect 2047 1578 2051 1582
rect 2079 1578 2083 1582
rect 2207 1578 2211 1582
rect 2343 1578 2347 1582
rect 2367 1578 2371 1582
rect 2487 1578 2491 1582
rect 2527 1578 2531 1582
rect 1871 1494 1875 1498
rect 1903 1494 1907 1498
rect 2007 1494 2011 1498
rect 2055 1494 2059 1498
rect 2135 1494 2139 1498
rect 1007 1434 1011 1438
rect 1047 1434 1051 1438
rect 1111 1434 1115 1438
rect 1207 1434 1211 1438
rect 1311 1434 1315 1438
rect 359 1358 363 1362
rect 455 1358 459 1362
rect 471 1358 475 1362
rect 551 1358 555 1362
rect 591 1358 595 1362
rect 639 1358 643 1362
rect 727 1358 731 1362
rect 815 1358 819 1362
rect 1243 1368 1247 1372
rect 1383 1434 1387 1438
rect 1415 1434 1419 1438
rect 1575 1434 1579 1438
rect 1743 1434 1747 1438
rect 1831 1434 1835 1438
rect 1871 1418 1875 1422
rect 1895 1418 1899 1422
rect 1519 1368 1523 1372
rect 863 1358 867 1362
rect 927 1358 931 1362
rect 1007 1358 1011 1362
rect 1055 1358 1059 1362
rect 1143 1358 1147 1362
rect 1215 1358 1219 1362
rect 1279 1358 1283 1362
rect 1391 1358 1395 1362
rect 1407 1358 1411 1362
rect 1527 1358 1531 1362
rect 1583 1358 1587 1362
rect 1647 1358 1651 1362
rect 1751 1358 1755 1362
rect 111 1278 115 1282
rect 311 1278 315 1282
rect 351 1278 355 1282
rect 415 1278 419 1282
rect 463 1278 467 1282
rect 535 1278 539 1282
rect 583 1278 587 1282
rect 671 1278 675 1282
rect 111 1202 115 1206
rect 239 1202 243 1206
rect 719 1278 723 1282
rect 815 1278 819 1282
rect 855 1278 859 1282
rect 959 1278 963 1282
rect 999 1278 1003 1282
rect 1103 1278 1107 1282
rect 1135 1278 1139 1282
rect 2215 1494 2219 1498
rect 2271 1494 2275 1498
rect 2375 1494 2379 1498
rect 2415 1494 2419 1498
rect 2631 1578 2635 1582
rect 2687 1578 2691 1582
rect 2775 1578 2779 1582
rect 2839 1578 2843 1582
rect 2919 1578 2923 1582
rect 2983 1578 2987 1582
rect 3063 1578 3067 1582
rect 3119 1578 3123 1582
rect 2535 1494 2539 1498
rect 2567 1494 2571 1498
rect 2695 1494 2699 1498
rect 2719 1494 2723 1498
rect 2847 1494 2851 1498
rect 2879 1494 2883 1498
rect 2991 1494 2995 1498
rect 3039 1494 3043 1498
rect 3463 1742 3467 1746
rect 3503 1742 3507 1746
rect 3591 1742 3595 1746
rect 3399 1662 3403 1666
rect 3511 1662 3515 1666
rect 3591 1662 3595 1666
rect 3215 1578 3219 1582
rect 3255 1578 3259 1582
rect 3367 1578 3371 1582
rect 3391 1578 3395 1582
rect 3503 1578 3507 1582
rect 3127 1494 3131 1498
rect 3199 1494 3203 1498
rect 3263 1494 3267 1498
rect 3367 1494 3371 1498
rect 3399 1494 3403 1498
rect 3591 1578 3595 1582
rect 3511 1494 3515 1498
rect 3591 1494 3595 1498
rect 1999 1418 2003 1422
rect 2023 1418 2027 1422
rect 1831 1358 1835 1362
rect 2127 1418 2131 1422
rect 2167 1418 2171 1422
rect 2263 1418 2267 1422
rect 2303 1418 2307 1422
rect 2407 1418 2411 1422
rect 2431 1418 2435 1422
rect 2551 1418 2555 1422
rect 2559 1418 2563 1422
rect 2671 1418 2675 1422
rect 2711 1418 2715 1422
rect 2791 1418 2795 1422
rect 2871 1418 2875 1422
rect 2911 1418 2915 1422
rect 3031 1418 3035 1422
rect 3191 1418 3195 1422
rect 3359 1418 3363 1422
rect 3503 1418 3507 1422
rect 3591 1418 3595 1422
rect 2619 1344 2623 1348
rect 1871 1334 1875 1338
rect 1903 1334 1907 1338
rect 1927 1334 1931 1338
rect 2031 1334 2035 1338
rect 2047 1334 2051 1338
rect 2175 1334 2179 1338
rect 2183 1334 2187 1338
rect 2311 1334 2315 1338
rect 2319 1334 2323 1338
rect 2439 1334 2443 1338
rect 2455 1334 2459 1338
rect 2559 1334 2563 1338
rect 2591 1334 2595 1338
rect 1307 1296 1311 1300
rect 1599 1296 1603 1300
rect 1239 1278 1243 1282
rect 1271 1278 1275 1282
rect 1375 1278 1379 1282
rect 1399 1278 1403 1282
rect 1503 1278 1507 1282
rect 1519 1278 1523 1282
rect 1987 1323 1991 1324
rect 1987 1320 1991 1323
rect 2327 1320 2331 1324
rect 2875 1344 2879 1348
rect 2679 1334 2683 1338
rect 2719 1334 2723 1338
rect 2799 1334 2803 1338
rect 2839 1334 2843 1338
rect 2919 1334 2923 1338
rect 2951 1334 2955 1338
rect 3063 1334 3067 1338
rect 3183 1334 3187 1338
rect 3591 1334 3595 1338
rect 1631 1278 1635 1282
rect 1639 1278 1643 1282
rect 1743 1278 1747 1282
rect 1831 1278 1835 1282
rect 1871 1250 1875 1254
rect 1895 1250 1899 1254
rect 1919 1250 1923 1254
rect 2039 1250 2043 1254
rect 2071 1250 2075 1254
rect 2175 1250 2179 1254
rect 319 1202 323 1206
rect 415 1202 419 1206
rect 423 1202 427 1206
rect 543 1202 547 1206
rect 591 1202 595 1206
rect 679 1202 683 1206
rect 759 1202 763 1206
rect 823 1202 827 1206
rect 927 1202 931 1206
rect 967 1202 971 1206
rect 1079 1202 1083 1206
rect 1111 1202 1115 1206
rect 1223 1202 1227 1206
rect 1247 1202 1251 1206
rect 1367 1202 1371 1206
rect 1383 1202 1387 1206
rect 1503 1202 1507 1206
rect 1511 1202 1515 1206
rect 1639 1202 1643 1206
rect 1751 1202 1755 1206
rect 111 1122 115 1126
rect 143 1122 147 1126
rect 231 1122 235 1126
rect 279 1122 283 1126
rect 407 1122 411 1126
rect 423 1122 427 1126
rect 111 1038 115 1042
rect 143 1038 147 1042
rect 151 1038 155 1042
rect 567 1122 571 1126
rect 583 1122 587 1126
rect 711 1122 715 1126
rect 751 1122 755 1126
rect 847 1122 851 1126
rect 919 1122 923 1126
rect 1831 1202 1835 1206
rect 1871 1170 1875 1174
rect 1903 1170 1907 1174
rect 2271 1250 2275 1254
rect 2311 1250 2315 1254
rect 2447 1250 2451 1254
rect 2471 1250 2475 1254
rect 2583 1250 2587 1254
rect 2663 1250 2667 1254
rect 2711 1250 2715 1254
rect 2831 1250 2835 1254
rect 2847 1250 2851 1254
rect 2943 1250 2947 1254
rect 3023 1250 3027 1254
rect 3055 1250 3059 1254
rect 2507 1184 2511 1188
rect 1983 1170 1987 1174
rect 2079 1170 2083 1174
rect 2087 1170 2091 1174
rect 2215 1170 2219 1174
rect 2279 1170 2283 1174
rect 2367 1170 2371 1174
rect 2479 1170 2483 1174
rect 2527 1170 2531 1174
rect 2671 1170 2675 1174
rect 2687 1170 2691 1174
rect 2779 1184 2783 1188
rect 3175 1250 3179 1254
rect 3191 1250 3195 1254
rect 3359 1250 3363 1254
rect 3503 1250 3507 1254
rect 3591 1250 3595 1254
rect 2839 1170 2843 1174
rect 2855 1170 2859 1174
rect 2983 1170 2987 1174
rect 3031 1170 3035 1174
rect 3127 1170 3131 1174
rect 3199 1170 3203 1174
rect 3263 1170 3267 1174
rect 3367 1170 3371 1174
rect 3399 1170 3403 1174
rect 3511 1170 3515 1174
rect 975 1122 979 1126
rect 1071 1122 1075 1126
rect 1103 1122 1107 1126
rect 1215 1122 1219 1126
rect 1223 1122 1227 1126
rect 1343 1122 1347 1126
rect 1359 1122 1363 1126
rect 1471 1122 1475 1126
rect 1495 1122 1499 1126
rect 1631 1122 1635 1126
rect 1743 1122 1747 1126
rect 1831 1122 1835 1126
rect 263 1038 267 1042
rect 287 1038 291 1042
rect 407 1038 411 1042
rect 431 1038 435 1042
rect 551 1038 555 1042
rect 575 1038 579 1042
rect 1055 1051 1059 1052
rect 1055 1048 1059 1051
rect 1871 1086 1875 1090
rect 1895 1086 1899 1090
rect 1975 1086 1979 1090
rect 2079 1086 2083 1090
rect 2167 1086 2171 1090
rect 2207 1086 2211 1090
rect 1367 1048 1371 1052
rect 687 1038 691 1042
rect 719 1038 723 1042
rect 807 1038 811 1042
rect 855 1038 859 1042
rect 927 1038 931 1042
rect 983 1038 987 1042
rect 1039 1038 1043 1042
rect 1111 1038 1115 1042
rect 1143 1038 1147 1042
rect 1231 1038 1235 1042
rect 1247 1038 1251 1042
rect 1351 1038 1355 1042
rect 1359 1038 1363 1042
rect 111 954 115 958
rect 135 954 139 958
rect 215 954 219 958
rect 255 954 259 958
rect 327 954 331 958
rect 399 954 403 958
rect 447 954 451 958
rect 543 954 547 958
rect 567 954 571 958
rect 679 954 683 958
rect 687 954 691 958
rect 1479 1038 1483 1042
rect 1831 1038 1835 1042
rect 2255 1086 2259 1090
rect 2359 1086 2363 1090
rect 2479 1086 2483 1090
rect 2519 1086 2523 1090
rect 2607 1086 2611 1090
rect 2679 1086 2683 1090
rect 2751 1086 2755 1090
rect 2831 1086 2835 1090
rect 2895 1086 2899 1090
rect 1871 1010 1875 1014
rect 2347 1024 2351 1028
rect 2175 1010 2179 1014
rect 2263 1010 2267 1014
rect 2303 1010 2307 1014
rect 2563 1024 2567 1028
rect 2367 1010 2371 1014
rect 2383 1010 2387 1014
rect 2471 1010 2475 1014
rect 2487 1010 2491 1014
rect 2567 1010 2571 1014
rect 2615 1010 2619 1014
rect 2671 1010 2675 1014
rect 2759 1010 2763 1014
rect 2783 1010 2787 1014
rect 2975 1086 2979 1090
rect 3591 1170 3595 1174
rect 3047 1086 3051 1090
rect 3119 1086 3123 1090
rect 3207 1086 3211 1090
rect 3255 1086 3259 1090
rect 3367 1086 3371 1090
rect 3391 1086 3395 1090
rect 3503 1086 3507 1090
rect 3591 1086 3595 1090
rect 2903 1010 2907 1014
rect 2911 1010 2915 1014
rect 3055 1010 3059 1014
rect 3207 1010 3211 1014
rect 3215 1010 3219 1014
rect 3367 1010 3371 1014
rect 3375 1010 3379 1014
rect 799 954 803 958
rect 911 954 915 958
rect 919 954 923 958
rect 1015 954 1019 958
rect 1031 954 1035 958
rect 1119 954 1123 958
rect 1135 954 1139 958
rect 1223 954 1227 958
rect 1239 954 1243 958
rect 1327 954 1331 958
rect 1351 954 1355 958
rect 1831 954 1835 958
rect 1871 926 1875 930
rect 2279 926 2283 930
rect 2295 926 2299 930
rect 2359 926 2363 930
rect 2375 926 2379 930
rect 2439 926 2443 930
rect 2463 926 2467 930
rect 2519 926 2523 930
rect 2559 926 2563 930
rect 2607 926 2611 930
rect 2663 926 2667 930
rect 2703 926 2707 930
rect 111 870 115 874
rect 143 870 147 874
rect 223 870 227 874
rect 255 870 259 874
rect 335 870 339 874
rect 399 870 403 874
rect 455 870 459 874
rect 559 870 563 874
rect 575 870 579 874
rect 695 870 699 874
rect 719 870 723 874
rect 807 870 811 874
rect 871 870 875 874
rect 919 870 923 874
rect 1015 870 1019 874
rect 1023 870 1027 874
rect 1127 870 1131 874
rect 1151 870 1155 874
rect 111 782 115 786
rect 135 782 139 786
rect 247 782 251 786
rect 263 782 267 786
rect 391 782 395 786
rect 431 782 435 786
rect 551 782 555 786
rect 607 782 611 786
rect 711 782 715 786
rect 783 782 787 786
rect 863 782 867 786
rect 111 694 115 698
rect 143 694 147 698
rect 271 694 275 698
rect 295 694 299 698
rect 1231 870 1235 874
rect 1279 870 1283 874
rect 1335 870 1339 874
rect 1399 870 1403 874
rect 1519 870 1523 874
rect 1647 870 1651 874
rect 1831 870 1835 874
rect 951 782 955 786
rect 1007 782 1011 786
rect 1103 782 1107 786
rect 1143 782 1147 786
rect 1247 782 1251 786
rect 1271 782 1275 786
rect 1383 782 1387 786
rect 1391 782 1395 786
rect 1511 782 1515 786
rect 1639 782 1643 786
rect 1871 838 1875 842
rect 2167 838 2171 842
rect 2247 838 2251 842
rect 2287 838 2291 842
rect 2327 838 2331 842
rect 2367 838 2371 842
rect 2423 838 2427 842
rect 2775 926 2779 930
rect 2807 926 2811 930
rect 2903 926 2907 930
rect 2911 926 2915 930
rect 3015 926 3019 930
rect 3047 926 3051 930
rect 3511 1010 3515 1014
rect 3591 1010 3595 1014
rect 3111 926 3115 930
rect 3199 926 3203 930
rect 3215 926 3219 930
rect 3319 926 3323 930
rect 3359 926 3363 930
rect 3423 926 3427 930
rect 3503 926 3507 930
rect 2447 838 2451 842
rect 2527 838 2531 842
rect 2535 838 2539 842
rect 2615 838 2619 842
rect 2655 838 2659 842
rect 2711 838 2715 842
rect 2783 838 2787 842
rect 2815 838 2819 842
rect 2911 838 2915 842
rect 2919 838 2923 842
rect 3023 838 3027 842
rect 3039 838 3043 842
rect 3119 838 3123 842
rect 3159 838 3163 842
rect 3223 838 3227 842
rect 3279 838 3283 842
rect 3327 838 3331 842
rect 3407 838 3411 842
rect 1743 782 1747 786
rect 1831 782 1835 786
rect 1871 754 1875 758
rect 1895 754 1899 758
rect 1975 754 1979 758
rect 2071 754 2075 758
rect 2159 754 2163 758
rect 2183 754 2187 758
rect 2239 754 2243 758
rect 407 694 411 698
rect 439 694 443 698
rect 527 694 531 698
rect 615 694 619 698
rect 655 694 659 698
rect 783 694 787 698
rect 791 694 795 698
rect 903 694 907 698
rect 959 694 963 698
rect 111 614 115 618
rect 287 614 291 618
rect 311 614 315 618
rect 391 614 395 618
rect 399 614 403 618
rect 471 614 475 618
rect 519 614 523 618
rect 559 614 563 618
rect 111 526 115 530
rect 239 526 243 530
rect 647 614 651 618
rect 1023 694 1027 698
rect 1111 694 1115 698
rect 1135 694 1139 698
rect 735 614 739 618
rect 775 614 779 618
rect 823 614 827 618
rect 895 614 899 618
rect 911 614 915 618
rect 999 614 1003 618
rect 1015 614 1019 618
rect 319 526 323 530
rect 343 526 347 530
rect 399 526 403 530
rect 439 526 443 530
rect 479 526 483 530
rect 535 526 539 530
rect 567 526 571 530
rect 111 442 115 446
rect 135 442 139 446
rect 231 442 235 446
rect 247 442 251 446
rect 335 442 339 446
rect 375 442 379 446
rect 111 354 115 358
rect 143 354 147 358
rect 431 442 435 446
rect 631 526 635 530
rect 655 526 659 530
rect 719 526 723 530
rect 743 526 747 530
rect 807 526 811 530
rect 495 442 499 446
rect 527 442 531 446
rect 607 442 611 446
rect 623 442 627 446
rect 711 442 715 446
rect 719 442 723 446
rect 831 526 835 530
rect 1247 694 1251 698
rect 1255 694 1259 698
rect 1351 694 1355 698
rect 1391 694 1395 698
rect 1455 694 1459 698
rect 1519 694 1523 698
rect 1559 694 1563 698
rect 1647 694 1651 698
rect 1663 694 1667 698
rect 1751 694 1755 698
rect 1831 694 1835 698
rect 1199 680 1203 684
rect 1567 680 1571 684
rect 1707 656 1711 660
rect 1871 674 1875 678
rect 1903 674 1907 678
rect 1983 674 1987 678
rect 2079 674 2083 678
rect 2095 674 2099 678
rect 2311 754 2315 758
rect 2319 754 2323 758
rect 2415 754 2419 758
rect 2447 754 2451 758
rect 2527 754 2531 758
rect 2591 754 2595 758
rect 2647 754 2651 758
rect 2743 754 2747 758
rect 2775 754 2779 758
rect 2191 674 2195 678
rect 2295 674 2299 678
rect 2319 674 2323 678
rect 2455 674 2459 678
rect 2479 674 2483 678
rect 2895 754 2899 758
rect 2903 754 2907 758
rect 3031 754 3035 758
rect 3047 754 3051 758
rect 3431 838 3435 842
rect 3591 926 3595 930
rect 3511 838 3515 842
rect 3591 838 3595 842
rect 3151 754 3155 758
rect 3199 754 3203 758
rect 3271 754 3275 758
rect 3359 754 3363 758
rect 3399 754 3403 758
rect 3503 754 3507 758
rect 2599 674 2603 678
rect 2655 674 2659 678
rect 2751 674 2755 678
rect 2831 674 2835 678
rect 2903 674 2907 678
rect 3007 674 3011 678
rect 3055 674 3059 678
rect 3183 674 3187 678
rect 3207 674 3211 678
rect 3359 674 3363 678
rect 3367 674 3371 678
rect 2303 656 2307 660
rect 1087 614 1091 618
rect 1127 614 1131 618
rect 1175 614 1179 618
rect 1239 614 1243 618
rect 1263 614 1267 618
rect 1343 614 1347 618
rect 1447 614 1451 618
rect 1551 614 1555 618
rect 1655 614 1659 618
rect 1743 614 1747 618
rect 1831 614 1835 618
rect 1871 594 1875 598
rect 1895 594 1899 598
rect 895 526 899 530
rect 919 526 923 530
rect 983 526 987 530
rect 1007 526 1011 530
rect 1071 526 1075 530
rect 1095 526 1099 530
rect 1159 526 1163 530
rect 1183 526 1187 530
rect 1247 526 1251 530
rect 1271 526 1275 530
rect 1831 526 1835 530
rect 883 512 887 516
rect 1255 512 1259 516
rect 1975 594 1979 598
rect 2087 594 2091 598
rect 2215 594 2219 598
rect 2287 594 2291 598
rect 2351 594 2355 598
rect 2471 594 2475 598
rect 2495 594 2499 598
rect 2647 594 2651 598
rect 1871 518 1875 522
rect 2179 536 2183 540
rect 1903 518 1907 522
rect 1983 518 1987 522
rect 2095 518 2099 522
rect 2151 518 2155 522
rect 2451 536 2455 540
rect 2807 594 2811 598
rect 2823 594 2827 598
rect 3591 754 3595 758
rect 3511 674 3515 678
rect 3591 674 3595 678
rect 2975 594 2979 598
rect 2999 594 3003 598
rect 3151 594 3155 598
rect 3175 594 3179 598
rect 3335 594 3339 598
rect 3351 594 3355 598
rect 3503 594 3507 598
rect 2223 518 2227 522
rect 2231 518 2235 522
rect 2327 518 2331 522
rect 2359 518 2363 522
rect 2431 518 2435 522
rect 2503 518 2507 522
rect 2551 518 2555 522
rect 2655 518 2659 522
rect 2687 518 2691 522
rect 2815 518 2819 522
rect 2839 518 2843 522
rect 3591 594 3595 598
rect 2983 518 2987 522
rect 2999 518 3003 522
rect 3159 518 3163 522
rect 3175 518 3179 522
rect 3343 518 3347 522
rect 3351 518 3355 522
rect 799 442 803 446
rect 823 442 827 446
rect 887 442 891 446
rect 919 442 923 446
rect 975 442 979 446
rect 1007 442 1011 446
rect 1063 442 1067 446
rect 1103 442 1107 446
rect 1151 442 1155 446
rect 1199 442 1203 446
rect 1239 442 1243 446
rect 1295 442 1299 446
rect 1831 442 1835 446
rect 1871 438 1875 442
rect 2143 438 2147 442
rect 2223 438 2227 442
rect 2319 438 2323 442
rect 2335 438 2339 442
rect 2415 438 2419 442
rect 2423 438 2427 442
rect 2495 438 2499 442
rect 2543 438 2547 442
rect 2583 438 2587 442
rect 2679 438 2683 442
rect 2687 438 2691 442
rect 247 354 251 358
rect 255 354 259 358
rect 375 354 379 358
rect 383 354 387 358
rect 503 354 507 358
rect 511 354 515 358
rect 615 354 619 358
rect 647 354 651 358
rect 727 354 731 358
rect 775 354 779 358
rect 111 270 115 274
rect 135 270 139 274
rect 223 270 227 274
rect 239 270 243 274
rect 335 270 339 274
rect 367 270 371 274
rect 463 270 467 274
rect 503 270 507 274
rect 111 162 115 166
rect 159 162 163 166
rect 599 270 603 274
rect 639 270 643 274
rect 831 354 835 358
rect 895 354 899 358
rect 927 354 931 358
rect 1007 354 1011 358
rect 1015 354 1019 358
rect 1111 354 1115 358
rect 1119 354 1123 358
rect 1207 354 1211 358
rect 1223 354 1227 358
rect 1303 354 1307 358
rect 1327 354 1331 358
rect 1439 354 1443 358
rect 1831 354 1835 358
rect 735 270 739 274
rect 767 270 771 274
rect 871 270 875 274
rect 887 270 891 274
rect 999 270 1003 274
rect 1007 270 1011 274
rect 1111 270 1115 274
rect 1135 270 1139 274
rect 1215 270 1219 274
rect 1255 270 1259 274
rect 1319 270 1323 274
rect 1871 354 1875 358
rect 2079 354 2083 358
rect 2167 354 2171 358
rect 2263 354 2267 358
rect 2343 354 2347 358
rect 2375 354 2379 358
rect 2423 354 2427 358
rect 2503 354 2507 358
rect 2799 438 2803 442
rect 2831 438 2835 442
rect 2927 438 2931 442
rect 2991 438 2995 442
rect 2591 354 2595 358
rect 2639 354 2643 358
rect 2695 354 2699 358
rect 2775 354 2779 358
rect 3071 438 3075 442
rect 3167 438 3171 442
rect 3511 518 3515 522
rect 3591 518 3595 522
rect 3215 438 3219 442
rect 3343 438 3347 442
rect 3367 438 3371 442
rect 3503 438 3507 442
rect 2807 354 2811 358
rect 2911 354 2915 358
rect 2935 354 2939 358
rect 3039 354 3043 358
rect 3079 354 3083 358
rect 3167 354 3171 358
rect 3223 354 3227 358
rect 3287 354 3291 358
rect 1367 270 1371 274
rect 1431 270 1435 274
rect 1479 270 1483 274
rect 1599 270 1603 274
rect 1831 270 1835 274
rect 1871 270 1875 274
rect 1895 270 1899 274
rect 1983 270 1987 274
rect 2071 270 2075 274
rect 2095 270 2099 274
rect 2159 270 2163 274
rect 2223 270 2227 274
rect 231 162 235 166
rect 239 162 243 166
rect 319 162 323 166
rect 343 162 347 166
rect 399 162 403 166
rect 471 162 475 166
rect 479 162 483 166
rect 559 162 563 166
rect 607 162 611 166
rect 647 162 651 166
rect 735 162 739 166
rect 743 162 747 166
rect 823 162 827 166
rect 879 162 883 166
rect 1043 208 1047 212
rect 911 162 915 166
rect 999 162 1003 166
rect 1015 162 1019 166
rect 1087 162 1091 166
rect 1143 162 1147 166
rect 1571 208 1575 212
rect 1931 208 1935 212
rect 1871 182 1875 186
rect 1903 182 1907 186
rect 1983 182 1987 186
rect 1991 182 1995 186
rect 2087 182 2091 186
rect 2103 182 2107 186
rect 1167 162 1171 166
rect 1247 162 1251 166
rect 1263 162 1267 166
rect 1335 162 1339 166
rect 1375 162 1379 166
rect 1423 162 1427 166
rect 1487 162 1491 166
rect 1511 162 1515 166
rect 1591 162 1595 166
rect 1607 162 1611 166
rect 1671 162 1675 166
rect 1751 162 1755 166
rect 1831 162 1835 166
rect 2255 270 2259 274
rect 2359 270 2363 274
rect 2367 270 2371 274
rect 2495 270 2499 274
rect 2503 270 2507 274
rect 2631 270 2635 274
rect 2647 270 2651 274
rect 2767 270 2771 274
rect 2791 270 2795 274
rect 2903 270 2907 274
rect 2935 270 2939 274
rect 2459 208 2463 212
rect 2207 182 2211 186
rect 2231 182 2235 186
rect 2335 182 2339 186
rect 2367 182 2371 186
rect 2463 182 2467 186
rect 2511 182 2515 186
rect 2583 182 2587 186
rect 2155 171 2159 172
rect 2155 168 2159 171
rect 2471 168 2475 172
rect 3031 270 3035 274
rect 3375 354 3379 358
rect 3407 354 3411 358
rect 3591 438 3595 442
rect 3511 354 3515 358
rect 3591 354 3595 358
rect 3079 270 3083 274
rect 3159 270 3163 274
rect 3223 270 3227 274
rect 3279 270 3283 274
rect 3375 270 3379 274
rect 3399 270 3403 274
rect 3503 270 3507 274
rect 2655 182 2659 186
rect 2703 182 2707 186
rect 2799 182 2803 186
rect 2815 182 2819 186
rect 2919 182 2923 186
rect 2943 182 2947 186
rect 3015 182 3019 186
rect 3087 182 3091 186
rect 3111 182 3115 186
rect 3207 182 3211 186
rect 3231 182 3235 186
rect 3303 182 3307 186
rect 3383 182 3387 186
rect 3399 182 3403 186
rect 3591 270 3595 274
rect 3511 182 3515 186
rect 3591 182 3595 186
rect 1871 106 1875 110
rect 1895 106 1899 110
rect 1975 106 1979 110
rect 2079 106 2083 110
rect 2199 106 2203 110
rect 2327 106 2331 110
rect 2455 106 2459 110
rect 2575 106 2579 110
rect 2695 106 2699 110
rect 2807 106 2811 110
rect 2911 106 2915 110
rect 3007 106 3011 110
rect 3103 106 3107 110
rect 3199 106 3203 110
rect 3295 106 3299 110
rect 3391 106 3395 110
rect 3591 106 3595 110
rect 111 86 115 90
rect 151 86 155 90
rect 231 86 235 90
rect 311 86 315 90
rect 391 86 395 90
rect 471 86 475 90
rect 551 86 555 90
rect 639 86 643 90
rect 727 86 731 90
rect 815 86 819 90
rect 903 86 907 90
rect 991 86 995 90
rect 1079 86 1083 90
rect 1159 86 1163 90
rect 1239 86 1243 90
rect 1327 86 1331 90
rect 1415 86 1419 90
rect 1503 86 1507 90
rect 1583 86 1587 90
rect 1663 86 1667 90
rect 1743 86 1747 90
rect 1831 86 1835 90
<< m4 >>
rect 1842 3665 1843 3671
rect 1849 3670 3619 3671
rect 1849 3666 1871 3670
rect 1875 3666 2151 3670
rect 2155 3666 2439 3670
rect 2443 3666 2727 3670
rect 2731 3666 3015 3670
rect 3019 3666 3591 3670
rect 3595 3666 3619 3670
rect 1849 3665 3619 3666
rect 3625 3665 3626 3671
rect 96 3637 97 3643
rect 103 3642 1855 3643
rect 103 3638 111 3642
rect 115 3638 143 3642
rect 147 3638 239 3642
rect 243 3638 367 3642
rect 371 3638 503 3642
rect 507 3638 639 3642
rect 643 3638 775 3642
rect 779 3638 911 3642
rect 915 3638 1055 3642
rect 1059 3638 1199 3642
rect 1203 3638 1831 3642
rect 1835 3638 1855 3642
rect 103 3637 1855 3638
rect 1861 3637 1862 3643
rect 1854 3589 1855 3595
rect 1861 3594 3631 3595
rect 1861 3590 1871 3594
rect 1875 3590 1903 3594
rect 1907 3590 1983 3594
rect 1987 3590 2071 3594
rect 2075 3590 2159 3594
rect 2163 3590 2175 3594
rect 2179 3590 2295 3594
rect 2299 3590 2423 3594
rect 2427 3590 2447 3594
rect 2451 3590 2559 3594
rect 2563 3590 2695 3594
rect 2699 3590 2735 3594
rect 2739 3590 2831 3594
rect 2835 3590 2975 3594
rect 2979 3590 3023 3594
rect 3027 3590 3119 3594
rect 3123 3590 3263 3594
rect 3267 3590 3591 3594
rect 3595 3590 3631 3594
rect 1861 3589 3631 3590
rect 3637 3589 3638 3595
rect 2502 3572 2508 3573
rect 2838 3572 2844 3573
rect 2502 3568 2503 3572
rect 2507 3568 2839 3572
rect 2843 3568 2844 3572
rect 2502 3567 2508 3568
rect 2838 3567 2844 3568
rect 84 3561 85 3567
rect 91 3566 1843 3567
rect 91 3562 111 3566
rect 115 3562 135 3566
rect 139 3562 183 3566
rect 187 3562 231 3566
rect 235 3562 303 3566
rect 307 3562 359 3566
rect 363 3562 415 3566
rect 419 3562 495 3566
rect 499 3562 527 3566
rect 531 3562 631 3566
rect 635 3562 735 3566
rect 739 3562 767 3566
rect 771 3562 831 3566
rect 835 3562 903 3566
rect 907 3562 919 3566
rect 923 3562 1007 3566
rect 1011 3562 1047 3566
rect 1051 3562 1095 3566
rect 1099 3562 1183 3566
rect 1187 3562 1191 3566
rect 1195 3562 1271 3566
rect 1275 3562 1359 3566
rect 1363 3562 1447 3566
rect 1451 3562 1831 3566
rect 1835 3562 1843 3566
rect 91 3561 1843 3562
rect 1849 3561 1850 3567
rect 1842 3513 1843 3519
rect 1849 3518 3619 3519
rect 1849 3514 1871 3518
rect 1875 3514 1895 3518
rect 1899 3514 1967 3518
rect 1971 3514 1975 3518
rect 1979 3514 2063 3518
rect 2067 3514 2151 3518
rect 2155 3514 2167 3518
rect 2171 3514 2287 3518
rect 2291 3514 2335 3518
rect 2339 3514 2415 3518
rect 2419 3514 2511 3518
rect 2515 3514 2551 3518
rect 2555 3514 2671 3518
rect 2675 3514 2687 3518
rect 2691 3514 2823 3518
rect 2827 3514 2959 3518
rect 2963 3514 2967 3518
rect 2971 3514 3079 3518
rect 3083 3514 3111 3518
rect 3115 3514 3191 3518
rect 3195 3514 3255 3518
rect 3259 3514 3303 3518
rect 3307 3514 3415 3518
rect 3419 3514 3503 3518
rect 3507 3514 3591 3518
rect 3595 3514 3619 3518
rect 1849 3513 3619 3514
rect 3625 3513 3626 3519
rect 986 3508 992 3509
rect 1434 3508 1440 3509
rect 986 3504 987 3508
rect 991 3504 1435 3508
rect 1439 3504 1440 3508
rect 986 3503 992 3504
rect 1434 3503 1440 3504
rect 96 3477 97 3483
rect 103 3482 1855 3483
rect 103 3478 111 3482
rect 115 3478 191 3482
rect 195 3478 231 3482
rect 235 3478 311 3482
rect 315 3478 367 3482
rect 371 3478 423 3482
rect 427 3478 503 3482
rect 507 3478 535 3482
rect 539 3478 623 3482
rect 627 3478 639 3482
rect 643 3478 735 3482
rect 739 3478 743 3482
rect 747 3478 839 3482
rect 843 3478 927 3482
rect 931 3478 943 3482
rect 947 3478 1015 3482
rect 1019 3478 1039 3482
rect 1043 3478 1103 3482
rect 1107 3478 1135 3482
rect 1139 3478 1191 3482
rect 1195 3478 1231 3482
rect 1235 3478 1279 3482
rect 1283 3478 1327 3482
rect 1331 3478 1367 3482
rect 1371 3478 1455 3482
rect 1459 3478 1831 3482
rect 1835 3478 1855 3482
rect 103 3477 1855 3478
rect 1861 3477 1862 3483
rect 1854 3437 1855 3443
rect 1861 3442 3631 3443
rect 1861 3438 1871 3442
rect 1875 3438 1975 3442
rect 1979 3438 2007 3442
rect 2011 3438 2127 3442
rect 2131 3438 2159 3442
rect 2163 3438 2255 3442
rect 2259 3438 2343 3442
rect 2347 3438 2391 3442
rect 2395 3438 2519 3442
rect 2523 3438 2535 3442
rect 2539 3438 2679 3442
rect 2683 3438 2831 3442
rect 2835 3438 2967 3442
rect 2971 3438 2999 3442
rect 3003 3438 3087 3442
rect 3091 3438 3167 3442
rect 3171 3438 3199 3442
rect 3203 3438 3311 3442
rect 3315 3438 3343 3442
rect 3347 3438 3423 3442
rect 3427 3438 3511 3442
rect 3515 3438 3591 3442
rect 3595 3438 3631 3442
rect 1861 3437 3631 3438
rect 3637 3437 3638 3443
rect 84 3397 85 3403
rect 91 3402 1843 3403
rect 91 3398 111 3402
rect 115 3398 215 3402
rect 219 3398 223 3402
rect 227 3398 359 3402
rect 363 3398 367 3402
rect 371 3398 495 3402
rect 499 3398 511 3402
rect 515 3398 615 3402
rect 619 3398 647 3402
rect 651 3398 727 3402
rect 731 3398 775 3402
rect 779 3398 831 3402
rect 835 3398 895 3402
rect 899 3398 935 3402
rect 939 3398 1015 3402
rect 1019 3398 1031 3402
rect 1035 3398 1127 3402
rect 1131 3398 1223 3402
rect 1227 3398 1239 3402
rect 1243 3398 1319 3402
rect 1323 3398 1351 3402
rect 1355 3398 1831 3402
rect 1835 3398 1843 3402
rect 91 3397 1843 3398
rect 1849 3397 1850 3403
rect 1842 3361 1843 3367
rect 1849 3366 3619 3367
rect 1849 3362 1871 3366
rect 1875 3362 1999 3366
rect 2003 3362 2015 3366
rect 2019 3362 2119 3366
rect 2123 3362 2151 3366
rect 2155 3362 2247 3366
rect 2251 3362 2295 3366
rect 2299 3362 2383 3366
rect 2387 3362 2439 3366
rect 2443 3362 2527 3366
rect 2531 3362 2583 3366
rect 2587 3362 2671 3366
rect 2675 3362 2727 3366
rect 2731 3362 2823 3366
rect 2827 3362 2871 3366
rect 2875 3362 2991 3366
rect 2995 3362 3023 3366
rect 3027 3362 3159 3366
rect 3163 3362 3183 3366
rect 3187 3362 3335 3366
rect 3339 3362 3351 3366
rect 3355 3362 3503 3366
rect 3507 3362 3591 3366
rect 3595 3362 3619 3366
rect 1849 3361 3619 3362
rect 3625 3361 3626 3367
rect 926 3356 932 3357
rect 1246 3356 1252 3357
rect 926 3352 927 3356
rect 931 3352 1247 3356
rect 1251 3352 1252 3356
rect 926 3351 932 3352
rect 1246 3351 1252 3352
rect 978 3340 984 3341
rect 1326 3340 1332 3341
rect 978 3336 979 3340
rect 983 3336 1327 3340
rect 1331 3336 1332 3340
rect 978 3335 984 3336
rect 1326 3335 1332 3336
rect 96 3317 97 3323
rect 103 3322 1855 3323
rect 103 3318 111 3322
rect 115 3318 207 3322
rect 211 3318 223 3322
rect 227 3318 367 3322
rect 371 3318 375 3322
rect 379 3318 519 3322
rect 523 3318 655 3322
rect 659 3318 671 3322
rect 675 3318 783 3322
rect 787 3318 815 3322
rect 819 3318 903 3322
rect 907 3318 951 3322
rect 955 3318 1023 3322
rect 1027 3318 1087 3322
rect 1091 3318 1135 3322
rect 1139 3318 1215 3322
rect 1219 3318 1247 3322
rect 1251 3318 1343 3322
rect 1347 3318 1359 3322
rect 1363 3318 1471 3322
rect 1475 3318 1831 3322
rect 1835 3318 1855 3322
rect 103 3317 1855 3318
rect 1861 3317 1862 3323
rect 1854 3285 1855 3291
rect 1861 3290 3631 3291
rect 1861 3286 1871 3290
rect 1875 3286 1927 3290
rect 1931 3286 2023 3290
rect 2027 3286 2063 3290
rect 2067 3286 2159 3290
rect 2163 3286 2191 3290
rect 2195 3286 2303 3290
rect 2307 3286 2319 3290
rect 2323 3286 2447 3290
rect 2451 3286 2591 3290
rect 2595 3286 2735 3290
rect 2739 3286 2743 3290
rect 2747 3286 2879 3290
rect 2883 3286 2919 3290
rect 2923 3286 3031 3290
rect 3035 3286 3111 3290
rect 3115 3286 3191 3290
rect 3195 3286 3311 3290
rect 3315 3286 3359 3290
rect 3363 3286 3511 3290
rect 3515 3286 3591 3290
rect 3595 3286 3631 3290
rect 1861 3285 3631 3286
rect 3637 3285 3638 3291
rect 2786 3268 2792 3269
rect 3318 3268 3324 3269
rect 2786 3264 2787 3268
rect 2791 3264 3319 3268
rect 3323 3264 3324 3268
rect 2786 3263 2792 3264
rect 3318 3263 3324 3264
rect 84 3241 85 3247
rect 91 3246 1843 3247
rect 91 3242 111 3246
rect 115 3242 135 3246
rect 139 3242 199 3246
rect 203 3242 271 3246
rect 275 3242 359 3246
rect 363 3242 415 3246
rect 419 3242 511 3246
rect 515 3242 575 3246
rect 579 3242 663 3246
rect 667 3242 735 3246
rect 739 3242 807 3246
rect 811 3242 895 3246
rect 899 3242 943 3246
rect 947 3242 1047 3246
rect 1051 3242 1079 3246
rect 1083 3242 1191 3246
rect 1195 3242 1207 3246
rect 1211 3242 1327 3246
rect 1331 3242 1335 3246
rect 1339 3242 1463 3246
rect 1467 3242 1607 3246
rect 1611 3242 1831 3246
rect 1835 3242 1843 3246
rect 91 3241 1843 3242
rect 1849 3241 1850 3247
rect 1842 3209 1843 3215
rect 1849 3214 3619 3215
rect 1849 3210 1871 3214
rect 1875 3210 1895 3214
rect 1899 3210 1919 3214
rect 1923 3210 2007 3214
rect 2011 3210 2055 3214
rect 2059 3210 2143 3214
rect 2147 3210 2183 3214
rect 2187 3210 2295 3214
rect 2299 3210 2311 3214
rect 2315 3210 2439 3214
rect 2443 3210 2455 3214
rect 2459 3210 2583 3214
rect 2587 3210 2623 3214
rect 2627 3210 2735 3214
rect 2739 3210 2799 3214
rect 2803 3210 2911 3214
rect 2915 3210 2975 3214
rect 2979 3210 3103 3214
rect 3107 3210 3151 3214
rect 3155 3210 3303 3214
rect 3307 3210 3327 3214
rect 3331 3210 3503 3214
rect 3507 3210 3591 3214
rect 3595 3210 3619 3214
rect 1849 3209 3619 3210
rect 3625 3209 3626 3215
rect 1582 3191 1583 3197
rect 1589 3196 1592 3197
rect 1591 3192 1592 3196
rect 1589 3191 1592 3192
rect 1078 3180 1084 3181
rect 1398 3180 1404 3181
rect 1078 3176 1079 3180
rect 1083 3176 1399 3180
rect 1403 3176 1404 3180
rect 1078 3175 1084 3176
rect 1398 3175 1404 3176
rect 910 3167 911 3173
rect 917 3167 918 3173
rect 96 3157 97 3163
rect 103 3162 1855 3163
rect 103 3158 111 3162
rect 115 3158 143 3162
rect 147 3158 175 3162
rect 179 3158 279 3162
rect 283 3158 319 3162
rect 323 3158 423 3162
rect 427 3158 463 3162
rect 467 3158 583 3162
rect 587 3158 607 3162
rect 611 3158 743 3162
rect 747 3158 871 3162
rect 875 3158 903 3162
rect 907 3158 991 3162
rect 995 3158 1055 3162
rect 1059 3158 1103 3162
rect 1107 3158 1199 3162
rect 1203 3158 1207 3162
rect 1211 3158 1311 3162
rect 1315 3158 1335 3162
rect 1339 3158 1407 3162
rect 1411 3158 1471 3162
rect 1475 3158 1495 3162
rect 1499 3158 1583 3162
rect 1587 3158 1615 3162
rect 1619 3158 1671 3162
rect 1675 3158 1751 3162
rect 1755 3158 1831 3162
rect 1835 3158 1855 3162
rect 103 3157 1855 3158
rect 1861 3157 1862 3163
rect 1854 3133 1855 3139
rect 1861 3138 3631 3139
rect 1861 3134 1871 3138
rect 1875 3134 1903 3138
rect 1907 3134 2015 3138
rect 2019 3134 2071 3138
rect 2075 3134 2151 3138
rect 2155 3134 2263 3138
rect 2267 3134 2303 3138
rect 2307 3134 2455 3138
rect 2459 3134 2463 3138
rect 2467 3134 2631 3138
rect 2635 3134 2647 3138
rect 2651 3134 2807 3138
rect 2811 3134 2831 3138
rect 2835 3134 2983 3138
rect 2987 3134 3015 3138
rect 3019 3134 3159 3138
rect 3163 3134 3199 3138
rect 3203 3134 3335 3138
rect 3339 3134 3391 3138
rect 3395 3134 3511 3138
rect 3515 3134 3591 3138
rect 3595 3134 3631 3138
rect 1861 3133 3631 3134
rect 3637 3133 3638 3139
rect 84 3069 85 3075
rect 91 3074 1843 3075
rect 91 3070 111 3074
rect 115 3070 135 3074
rect 139 3070 167 3074
rect 171 3070 223 3074
rect 227 3070 311 3074
rect 315 3070 327 3074
rect 331 3070 439 3074
rect 443 3070 455 3074
rect 459 3070 551 3074
rect 555 3070 599 3074
rect 603 3070 663 3074
rect 667 3070 735 3074
rect 739 3070 863 3074
rect 867 3070 983 3074
rect 987 3070 1095 3074
rect 1099 3070 1199 3074
rect 1203 3070 1303 3074
rect 1307 3070 1399 3074
rect 1403 3070 1487 3074
rect 1491 3070 1575 3074
rect 1579 3070 1663 3074
rect 1667 3070 1743 3074
rect 1747 3070 1831 3074
rect 1835 3070 1843 3074
rect 91 3069 1843 3070
rect 1849 3069 1850 3075
rect 1842 3045 1843 3051
rect 1849 3050 3619 3051
rect 1849 3046 1871 3050
rect 1875 3046 1895 3050
rect 1899 3046 2063 3050
rect 2067 3046 2199 3050
rect 2203 3046 2255 3050
rect 2259 3046 2335 3050
rect 2339 3046 2447 3050
rect 2451 3046 2479 3050
rect 2483 3046 2623 3050
rect 2627 3046 2639 3050
rect 2643 3046 2767 3050
rect 2771 3046 2823 3050
rect 2827 3046 2903 3050
rect 2907 3046 3007 3050
rect 3011 3046 3039 3050
rect 3043 3046 3183 3050
rect 3187 3046 3191 3050
rect 3195 3046 3327 3050
rect 3331 3046 3383 3050
rect 3387 3046 3591 3050
rect 3595 3046 3619 3050
rect 1849 3045 3619 3046
rect 3625 3045 3626 3051
rect 96 2981 97 2987
rect 103 2986 1855 2987
rect 103 2982 111 2986
rect 115 2982 143 2986
rect 147 2982 159 2986
rect 163 2982 231 2986
rect 235 2982 319 2986
rect 323 2982 335 2986
rect 339 2982 447 2986
rect 451 2982 487 2986
rect 491 2982 559 2986
rect 563 2982 647 2986
rect 651 2982 671 2986
rect 675 2982 799 2986
rect 803 2982 943 2986
rect 947 2982 1079 2986
rect 1083 2982 1199 2986
rect 1203 2982 1311 2986
rect 1315 2982 1423 2986
rect 1427 2982 1535 2986
rect 1539 2982 1647 2986
rect 1651 2982 1831 2986
rect 1835 2982 1855 2986
rect 103 2981 1855 2982
rect 1861 2981 1862 2987
rect 1854 2957 1855 2963
rect 1861 2962 3631 2963
rect 1861 2958 1871 2962
rect 1875 2958 2127 2962
rect 2131 2958 2207 2962
rect 2211 2958 2287 2962
rect 2291 2958 2343 2962
rect 2347 2958 2367 2962
rect 2371 2958 2447 2962
rect 2451 2958 2487 2962
rect 2491 2958 2527 2962
rect 2531 2958 2607 2962
rect 2611 2958 2631 2962
rect 2635 2958 2695 2962
rect 2699 2958 2775 2962
rect 2779 2958 2791 2962
rect 2795 2958 2911 2962
rect 2915 2958 3039 2962
rect 3043 2958 3047 2962
rect 3051 2958 3183 2962
rect 3187 2958 3191 2962
rect 3195 2958 3335 2962
rect 3339 2958 3495 2962
rect 3499 2958 3591 2962
rect 3595 2958 3631 2962
rect 1861 2957 3631 2958
rect 3637 2957 3638 2963
rect 84 2905 85 2911
rect 91 2910 1843 2911
rect 91 2906 111 2910
rect 115 2906 151 2910
rect 155 2906 311 2910
rect 315 2906 471 2910
rect 475 2906 479 2910
rect 483 2906 631 2910
rect 635 2906 639 2910
rect 643 2906 783 2910
rect 787 2906 791 2910
rect 795 2906 927 2910
rect 931 2906 935 2910
rect 939 2906 1055 2910
rect 1059 2906 1071 2910
rect 1075 2906 1175 2910
rect 1179 2906 1191 2910
rect 1195 2906 1287 2910
rect 1291 2906 1303 2910
rect 1307 2906 1391 2910
rect 1395 2906 1415 2910
rect 1419 2906 1487 2910
rect 1491 2906 1527 2910
rect 1531 2906 1591 2910
rect 1595 2906 1639 2910
rect 1643 2906 1695 2910
rect 1699 2906 1831 2910
rect 1835 2906 1843 2910
rect 91 2905 1843 2906
rect 1849 2905 1850 2911
rect 1842 2881 1843 2887
rect 1849 2886 3619 2887
rect 1849 2882 1871 2886
rect 1875 2882 2047 2886
rect 2051 2882 2119 2886
rect 2123 2882 2135 2886
rect 2139 2882 2199 2886
rect 2203 2882 2239 2886
rect 2243 2882 2279 2886
rect 2283 2882 2343 2886
rect 2347 2882 2359 2886
rect 2363 2882 2439 2886
rect 2443 2882 2463 2886
rect 2467 2882 2519 2886
rect 2523 2882 2591 2886
rect 2595 2882 2599 2886
rect 2603 2882 2687 2886
rect 2691 2882 2727 2886
rect 2731 2882 2783 2886
rect 2787 2882 2879 2886
rect 2883 2882 2903 2886
rect 2907 2882 3031 2886
rect 3035 2882 3175 2886
rect 3179 2882 3191 2886
rect 3195 2882 3327 2886
rect 3331 2882 3359 2886
rect 3363 2882 3487 2886
rect 3491 2882 3503 2886
rect 3507 2882 3591 2886
rect 3595 2882 3619 2886
rect 1849 2881 3619 2882
rect 3625 2881 3626 2887
rect 1434 2852 1440 2853
rect 1674 2852 1680 2853
rect 1434 2848 1435 2852
rect 1439 2848 1675 2852
rect 1679 2848 1680 2852
rect 1434 2847 1440 2848
rect 1674 2847 1680 2848
rect 96 2825 97 2831
rect 103 2830 1855 2831
rect 103 2826 111 2830
rect 115 2826 143 2830
rect 147 2826 159 2830
rect 163 2826 247 2830
rect 251 2826 319 2830
rect 323 2826 383 2830
rect 387 2826 479 2830
rect 483 2826 535 2830
rect 539 2826 639 2830
rect 643 2826 687 2830
rect 691 2826 791 2830
rect 795 2826 847 2830
rect 851 2826 935 2830
rect 939 2826 999 2830
rect 1003 2826 1063 2830
rect 1067 2826 1143 2830
rect 1147 2826 1183 2830
rect 1187 2826 1279 2830
rect 1283 2826 1295 2830
rect 1299 2826 1399 2830
rect 1403 2826 1407 2830
rect 1411 2826 1495 2830
rect 1499 2826 1527 2830
rect 1531 2826 1599 2830
rect 1603 2826 1647 2830
rect 1651 2826 1703 2830
rect 1707 2826 1751 2830
rect 1755 2826 1831 2830
rect 1835 2826 1855 2830
rect 103 2825 1855 2826
rect 1861 2825 1862 2831
rect 2666 2820 2672 2821
rect 2958 2820 2964 2821
rect 2666 2816 2667 2820
rect 2671 2816 2959 2820
rect 2963 2816 2964 2820
rect 2666 2815 2672 2816
rect 2958 2815 2964 2816
rect 1854 2793 1855 2799
rect 1861 2798 3631 2799
rect 1861 2794 1871 2798
rect 1875 2794 1903 2798
rect 1907 2794 2015 2798
rect 2019 2794 2055 2798
rect 2059 2794 2143 2798
rect 2147 2794 2167 2798
rect 2171 2794 2247 2798
rect 2251 2794 2327 2798
rect 2331 2794 2351 2798
rect 2355 2794 2471 2798
rect 2475 2794 2487 2798
rect 2491 2794 2599 2798
rect 2603 2794 2639 2798
rect 2643 2794 2735 2798
rect 2739 2794 2791 2798
rect 2795 2794 2887 2798
rect 2891 2794 2943 2798
rect 2947 2794 3039 2798
rect 3043 2794 3087 2798
rect 3091 2794 3199 2798
rect 3203 2794 3231 2798
rect 3235 2794 3367 2798
rect 3371 2794 3383 2798
rect 3387 2794 3511 2798
rect 3515 2794 3591 2798
rect 3595 2794 3631 2798
rect 1861 2793 3631 2794
rect 3637 2793 3638 2799
rect 2066 2780 2072 2781
rect 2418 2780 2424 2781
rect 2066 2776 2067 2780
rect 2071 2776 2419 2780
rect 2423 2776 2424 2780
rect 2066 2775 2072 2776
rect 2418 2775 2424 2776
rect 84 2745 85 2751
rect 91 2750 1843 2751
rect 91 2746 111 2750
rect 115 2746 135 2750
rect 139 2746 231 2750
rect 235 2746 239 2750
rect 243 2746 367 2750
rect 371 2746 375 2750
rect 379 2746 511 2750
rect 515 2746 527 2750
rect 531 2746 663 2750
rect 667 2746 679 2750
rect 683 2746 815 2750
rect 819 2746 839 2750
rect 843 2746 975 2750
rect 979 2746 991 2750
rect 995 2746 1135 2750
rect 1139 2746 1271 2750
rect 1275 2746 1287 2750
rect 1291 2746 1399 2750
rect 1403 2746 1447 2750
rect 1451 2746 1519 2750
rect 1523 2746 1607 2750
rect 1611 2746 1639 2750
rect 1643 2746 1743 2750
rect 1747 2746 1831 2750
rect 1835 2746 1843 2750
rect 91 2745 1843 2746
rect 1849 2745 1850 2751
rect 1842 2717 1843 2723
rect 1849 2722 3619 2723
rect 1849 2718 1871 2722
rect 1875 2718 1895 2722
rect 1899 2718 2007 2722
rect 2011 2718 2103 2722
rect 2107 2718 2159 2722
rect 2163 2718 2319 2722
rect 2323 2718 2327 2722
rect 2331 2718 2479 2722
rect 2483 2718 2535 2722
rect 2539 2718 2631 2722
rect 2635 2718 2735 2722
rect 2739 2718 2783 2722
rect 2787 2718 2911 2722
rect 2915 2718 2935 2722
rect 2939 2718 3071 2722
rect 3075 2718 3079 2722
rect 3083 2718 3223 2722
rect 3227 2718 3375 2722
rect 3379 2718 3503 2722
rect 3507 2718 3591 2722
rect 3595 2718 3619 2722
rect 1849 2717 3619 2718
rect 3625 2717 3626 2723
rect 1006 2684 1012 2685
rect 1222 2684 1228 2685
rect 1006 2680 1007 2684
rect 1011 2680 1223 2684
rect 1227 2680 1228 2684
rect 1006 2679 1012 2680
rect 1222 2679 1228 2680
rect 96 2661 97 2667
rect 103 2666 1855 2667
rect 103 2662 111 2666
rect 115 2662 143 2666
rect 147 2662 239 2666
rect 243 2662 279 2666
rect 283 2662 375 2666
rect 379 2662 447 2666
rect 451 2662 519 2666
rect 523 2662 623 2666
rect 627 2662 671 2666
rect 675 2662 791 2666
rect 795 2662 823 2666
rect 827 2662 951 2666
rect 955 2662 983 2666
rect 987 2662 1103 2666
rect 1107 2662 1143 2666
rect 1147 2662 1247 2666
rect 1251 2662 1295 2666
rect 1299 2662 1399 2666
rect 1403 2662 1455 2666
rect 1459 2662 1551 2666
rect 1555 2662 1615 2666
rect 1619 2662 1751 2666
rect 1755 2662 1831 2666
rect 1835 2662 1855 2666
rect 103 2661 1855 2662
rect 1861 2661 1862 2667
rect 1930 2660 1936 2661
rect 2478 2660 2484 2661
rect 1930 2656 1931 2660
rect 1935 2656 2479 2660
rect 2483 2656 2484 2660
rect 1930 2655 1936 2656
rect 2478 2655 2484 2656
rect 2770 2660 2776 2661
rect 3138 2660 3144 2661
rect 2770 2656 2771 2660
rect 2775 2656 3139 2660
rect 3143 2656 3144 2660
rect 2770 2655 2776 2656
rect 3138 2655 3144 2656
rect 1854 2633 1855 2639
rect 1861 2638 3631 2639
rect 1861 2634 1871 2638
rect 1875 2634 1903 2638
rect 1907 2634 2055 2638
rect 2059 2634 2111 2638
rect 2115 2634 2263 2638
rect 2267 2634 2335 2638
rect 2339 2634 2495 2638
rect 2499 2634 2543 2638
rect 2547 2634 2743 2638
rect 2747 2634 2751 2638
rect 2755 2634 2919 2638
rect 2923 2634 3015 2638
rect 3019 2634 3079 2638
rect 3083 2634 3231 2638
rect 3235 2634 3287 2638
rect 3291 2634 3383 2638
rect 3387 2634 3511 2638
rect 3515 2634 3591 2638
rect 3595 2634 3631 2638
rect 1861 2633 3631 2634
rect 3637 2633 3638 2639
rect 84 2581 85 2587
rect 91 2586 1843 2587
rect 91 2582 111 2586
rect 115 2582 135 2586
rect 139 2582 223 2586
rect 227 2582 271 2586
rect 275 2582 367 2586
rect 371 2582 439 2586
rect 443 2582 527 2586
rect 531 2582 615 2586
rect 619 2582 703 2586
rect 707 2582 783 2586
rect 787 2582 879 2586
rect 883 2582 943 2586
rect 947 2582 1047 2586
rect 1051 2582 1095 2586
rect 1099 2582 1207 2586
rect 1211 2582 1239 2586
rect 1243 2582 1359 2586
rect 1363 2582 1391 2586
rect 1395 2582 1511 2586
rect 1515 2582 1543 2586
rect 1547 2582 1671 2586
rect 1675 2582 1831 2586
rect 1835 2582 1843 2586
rect 91 2581 1843 2582
rect 1849 2581 1850 2587
rect 1842 2557 1843 2563
rect 1849 2562 3619 2563
rect 1849 2558 1871 2562
rect 1875 2558 1895 2562
rect 1899 2558 2007 2562
rect 2011 2558 2047 2562
rect 2051 2558 2159 2562
rect 2163 2558 2255 2562
rect 2259 2558 2319 2562
rect 2323 2558 2471 2562
rect 2475 2558 2487 2562
rect 2491 2558 2623 2562
rect 2627 2558 2743 2562
rect 2747 2558 2759 2562
rect 2763 2558 2887 2562
rect 2891 2558 3007 2562
rect 3011 2558 3119 2562
rect 3123 2558 3223 2562
rect 3227 2558 3279 2562
rect 3283 2558 3319 2562
rect 3323 2558 3423 2562
rect 3427 2558 3503 2562
rect 3507 2558 3591 2562
rect 3595 2558 3619 2562
rect 1849 2557 3619 2558
rect 3625 2557 3626 2563
rect 1930 2532 1936 2533
rect 2658 2532 2664 2533
rect 1930 2528 1931 2532
rect 1935 2528 2659 2532
rect 2663 2528 2664 2532
rect 1930 2527 1936 2528
rect 2658 2527 2664 2528
rect 96 2501 97 2507
rect 103 2506 1855 2507
rect 103 2502 111 2506
rect 115 2502 143 2506
rect 147 2502 223 2506
rect 227 2502 231 2506
rect 235 2502 303 2506
rect 307 2502 375 2506
rect 379 2502 391 2506
rect 395 2502 511 2506
rect 515 2502 535 2506
rect 539 2502 647 2506
rect 651 2502 711 2506
rect 715 2502 783 2506
rect 787 2502 887 2506
rect 891 2502 927 2506
rect 931 2502 1055 2506
rect 1059 2502 1063 2506
rect 1067 2502 1191 2506
rect 1195 2502 1215 2506
rect 1219 2502 1311 2506
rect 1315 2502 1367 2506
rect 1371 2502 1431 2506
rect 1435 2502 1519 2506
rect 1523 2502 1551 2506
rect 1555 2502 1671 2506
rect 1675 2502 1679 2506
rect 1683 2502 1831 2506
rect 1835 2502 1855 2506
rect 103 2501 1855 2502
rect 1861 2501 1862 2507
rect 1854 2473 1855 2479
rect 1861 2478 3631 2479
rect 1861 2474 1871 2478
rect 1875 2474 1903 2478
rect 1907 2474 1999 2478
rect 2003 2474 2015 2478
rect 2019 2474 2127 2478
rect 2131 2474 2167 2478
rect 2171 2474 2263 2478
rect 2267 2474 2327 2478
rect 2331 2474 2407 2478
rect 2411 2474 2479 2478
rect 2483 2474 2551 2478
rect 2555 2474 2631 2478
rect 2635 2474 2703 2478
rect 2707 2474 2767 2478
rect 2771 2474 2863 2478
rect 2867 2474 2895 2478
rect 2899 2474 3015 2478
rect 3019 2474 3023 2478
rect 3027 2474 3127 2478
rect 3131 2474 3191 2478
rect 3195 2474 3231 2478
rect 3235 2474 3327 2478
rect 3331 2474 3359 2478
rect 3363 2474 3431 2478
rect 3435 2474 3511 2478
rect 3515 2474 3591 2478
rect 3595 2474 3631 2478
rect 1861 2473 3631 2474
rect 3637 2473 3638 2479
rect 1134 2460 1140 2461
rect 1470 2460 1476 2461
rect 1134 2456 1135 2460
rect 1139 2456 1471 2460
rect 1475 2456 1476 2460
rect 1134 2455 1140 2456
rect 1470 2455 1476 2456
rect 2802 2460 2808 2461
rect 3198 2460 3204 2461
rect 2802 2456 2803 2460
rect 2807 2456 3199 2460
rect 3203 2456 3204 2460
rect 2802 2455 2808 2456
rect 3198 2455 3204 2456
rect 84 2413 85 2419
rect 91 2418 1843 2419
rect 91 2414 111 2418
rect 115 2414 135 2418
rect 139 2414 215 2418
rect 219 2414 295 2418
rect 299 2414 383 2418
rect 387 2414 503 2418
rect 507 2414 639 2418
rect 643 2414 775 2418
rect 779 2414 919 2418
rect 923 2414 1055 2418
rect 1059 2414 1063 2418
rect 1067 2414 1143 2418
rect 1147 2414 1183 2418
rect 1187 2414 1223 2418
rect 1227 2414 1303 2418
rect 1307 2414 1383 2418
rect 1387 2414 1423 2418
rect 1427 2414 1463 2418
rect 1467 2414 1543 2418
rect 1547 2414 1663 2418
rect 1667 2414 1831 2418
rect 1835 2414 1843 2418
rect 91 2413 1843 2414
rect 1849 2413 1850 2419
rect 1842 2393 1843 2399
rect 1849 2398 3619 2399
rect 1849 2394 1871 2398
rect 1875 2394 1991 2398
rect 1995 2394 2119 2398
rect 2123 2394 2143 2398
rect 2147 2394 2239 2398
rect 2243 2394 2255 2398
rect 2259 2394 2343 2398
rect 2347 2394 2399 2398
rect 2403 2394 2455 2398
rect 2459 2394 2543 2398
rect 2547 2394 2575 2398
rect 2579 2394 2695 2398
rect 2699 2394 2703 2398
rect 2707 2394 2847 2398
rect 2851 2394 2855 2398
rect 2859 2394 3007 2398
rect 3011 2394 3015 2398
rect 3019 2394 3175 2398
rect 3179 2394 3183 2398
rect 3187 2394 3351 2398
rect 3355 2394 3503 2398
rect 3507 2394 3591 2398
rect 3595 2394 3619 2398
rect 1849 2393 3619 2394
rect 3625 2393 3626 2399
rect 96 2329 97 2335
rect 103 2334 1855 2335
rect 103 2330 111 2334
rect 115 2330 359 2334
rect 363 2330 439 2334
rect 443 2330 519 2334
rect 523 2330 599 2334
rect 603 2330 679 2334
rect 683 2330 759 2334
rect 763 2330 839 2334
rect 843 2330 919 2334
rect 923 2330 999 2334
rect 1003 2330 1071 2334
rect 1075 2330 1079 2334
rect 1083 2330 1151 2334
rect 1155 2330 1159 2334
rect 1163 2330 1231 2334
rect 1235 2330 1239 2334
rect 1243 2330 1311 2334
rect 1315 2330 1319 2334
rect 1323 2330 1391 2334
rect 1395 2330 1471 2334
rect 1475 2330 1831 2334
rect 1835 2330 1855 2334
rect 103 2329 1855 2330
rect 1861 2329 1862 2335
rect 2178 2332 2184 2333
rect 2478 2332 2484 2333
rect 2178 2328 2179 2332
rect 2183 2328 2479 2332
rect 2483 2328 2484 2332
rect 2178 2327 2184 2328
rect 2478 2327 2484 2328
rect 2882 2332 2888 2333
rect 3122 2332 3128 2333
rect 2882 2328 2883 2332
rect 2887 2328 3123 2332
rect 3127 2328 3128 2332
rect 2882 2327 2888 2328
rect 3122 2327 3128 2328
rect 1854 2313 1855 2319
rect 1861 2318 3631 2319
rect 1861 2314 1871 2318
rect 1875 2314 2151 2318
rect 2155 2314 2247 2318
rect 2251 2314 2279 2318
rect 2283 2314 2351 2318
rect 2355 2314 2359 2318
rect 2363 2314 2439 2318
rect 2443 2314 2463 2318
rect 2467 2314 2519 2318
rect 2523 2314 2583 2318
rect 2587 2314 2599 2318
rect 2603 2314 2679 2318
rect 2683 2314 2711 2318
rect 2715 2314 2759 2318
rect 2763 2314 2847 2318
rect 2851 2314 2855 2318
rect 2859 2314 2935 2318
rect 2939 2314 3015 2318
rect 3019 2314 3183 2318
rect 3187 2314 3359 2318
rect 3363 2314 3511 2318
rect 3515 2314 3591 2318
rect 3595 2314 3631 2318
rect 1861 2313 3631 2314
rect 3637 2313 3638 2319
rect 84 2253 85 2259
rect 91 2258 1843 2259
rect 91 2254 111 2258
rect 115 2254 351 2258
rect 355 2254 375 2258
rect 379 2254 431 2258
rect 435 2254 455 2258
rect 459 2254 511 2258
rect 515 2254 535 2258
rect 539 2254 591 2258
rect 595 2254 615 2258
rect 619 2254 671 2258
rect 675 2254 695 2258
rect 699 2254 751 2258
rect 755 2254 775 2258
rect 779 2254 831 2258
rect 835 2254 855 2258
rect 859 2254 911 2258
rect 915 2254 935 2258
rect 939 2254 991 2258
rect 995 2254 1015 2258
rect 1019 2254 1071 2258
rect 1075 2254 1095 2258
rect 1099 2254 1151 2258
rect 1155 2254 1175 2258
rect 1179 2254 1231 2258
rect 1235 2254 1255 2258
rect 1259 2254 1311 2258
rect 1315 2254 1831 2258
rect 1835 2254 1843 2258
rect 91 2253 1843 2254
rect 1849 2253 1850 2259
rect 1842 2237 1843 2243
rect 1849 2242 3619 2243
rect 1849 2238 1871 2242
rect 1875 2238 2271 2242
rect 2275 2238 2311 2242
rect 2315 2238 2351 2242
rect 2355 2238 2399 2242
rect 2403 2238 2431 2242
rect 2435 2238 2495 2242
rect 2499 2238 2511 2242
rect 2515 2238 2591 2242
rect 2595 2238 2599 2242
rect 2603 2238 2671 2242
rect 2675 2238 2719 2242
rect 2723 2238 2751 2242
rect 2755 2238 2839 2242
rect 2843 2238 2855 2242
rect 2859 2238 2927 2242
rect 2931 2238 3007 2242
rect 3011 2238 3175 2242
rect 3179 2238 3351 2242
rect 3355 2238 3503 2242
rect 3507 2238 3591 2242
rect 3595 2238 3619 2242
rect 1849 2237 3619 2238
rect 3625 2237 3626 2243
rect 2734 2180 2740 2181
rect 3082 2180 3088 2181
rect 2734 2176 2735 2180
rect 2739 2176 3083 2180
rect 3087 2176 3088 2180
rect 2734 2175 2740 2176
rect 3082 2175 3088 2176
rect 96 2165 97 2171
rect 103 2170 1855 2171
rect 103 2166 111 2170
rect 115 2166 311 2170
rect 315 2166 383 2170
rect 387 2166 407 2170
rect 411 2166 463 2170
rect 467 2166 503 2170
rect 507 2166 543 2170
rect 547 2166 599 2170
rect 603 2166 623 2170
rect 627 2166 687 2170
rect 691 2166 703 2170
rect 707 2166 775 2170
rect 779 2166 783 2170
rect 787 2166 863 2170
rect 867 2166 943 2170
rect 947 2166 951 2170
rect 955 2166 1023 2170
rect 1027 2166 1039 2170
rect 1043 2166 1103 2170
rect 1107 2166 1127 2170
rect 1131 2166 1183 2170
rect 1187 2166 1223 2170
rect 1227 2166 1263 2170
rect 1267 2166 1831 2170
rect 1835 2166 1855 2170
rect 103 2165 1855 2166
rect 1861 2165 1862 2171
rect 1854 2163 1862 2165
rect 1854 2157 1855 2163
rect 1861 2162 3631 2163
rect 1861 2158 1871 2162
rect 1875 2158 1903 2162
rect 1907 2158 1983 2162
rect 1987 2158 2111 2162
rect 2115 2158 2247 2162
rect 2251 2158 2319 2162
rect 2323 2158 2391 2162
rect 2395 2158 2407 2162
rect 2411 2158 2503 2162
rect 2507 2158 2543 2162
rect 2547 2158 2607 2162
rect 2611 2158 2695 2162
rect 2699 2158 2727 2162
rect 2731 2158 2847 2162
rect 2851 2158 2863 2162
rect 2867 2158 3007 2162
rect 3011 2158 3015 2162
rect 3019 2158 3175 2162
rect 3179 2158 3183 2162
rect 3187 2158 3351 2162
rect 3355 2158 3359 2162
rect 3363 2158 3511 2162
rect 3515 2158 3591 2162
rect 3595 2158 3631 2162
rect 1861 2157 3631 2158
rect 3637 2157 3638 2163
rect 84 2077 85 2083
rect 91 2082 1843 2083
rect 91 2078 111 2082
rect 115 2078 207 2082
rect 211 2078 303 2082
rect 307 2078 327 2082
rect 331 2078 399 2082
rect 403 2078 447 2082
rect 451 2078 495 2082
rect 499 2078 575 2082
rect 579 2078 591 2082
rect 595 2078 679 2082
rect 683 2078 703 2082
rect 707 2078 767 2082
rect 771 2078 823 2082
rect 827 2078 855 2082
rect 859 2078 943 2082
rect 947 2078 1031 2082
rect 1035 2078 1063 2082
rect 1067 2078 1119 2082
rect 1123 2078 1175 2082
rect 1179 2078 1215 2082
rect 1219 2078 1279 2082
rect 1283 2078 1375 2082
rect 1379 2078 1471 2082
rect 1475 2078 1567 2082
rect 1571 2078 1663 2082
rect 1667 2078 1743 2082
rect 1747 2078 1831 2082
rect 1835 2078 1843 2082
rect 91 2077 1843 2078
rect 1849 2079 1850 2083
rect 1849 2078 3626 2079
rect 1849 2077 1871 2078
rect 1842 2074 1871 2077
rect 1875 2074 1895 2078
rect 1899 2074 1967 2078
rect 1971 2074 1975 2078
rect 1979 2074 2103 2078
rect 2107 2074 2215 2078
rect 2219 2074 2239 2078
rect 2243 2074 2383 2078
rect 2387 2074 2447 2078
rect 2451 2074 2535 2078
rect 2539 2074 2655 2078
rect 2659 2074 2687 2078
rect 2691 2074 2839 2078
rect 2843 2074 2999 2078
rect 3003 2074 3143 2078
rect 3147 2074 3167 2078
rect 3171 2074 3271 2078
rect 3275 2074 3343 2078
rect 3347 2074 3399 2078
rect 3403 2074 3503 2078
rect 3507 2074 3591 2078
rect 3595 2074 3626 2078
rect 1842 2073 3626 2074
rect 2686 2012 2692 2013
rect 3086 2012 3092 2013
rect 2686 2008 2687 2012
rect 2691 2008 3087 2012
rect 3091 2008 3092 2012
rect 2686 2007 2692 2008
rect 3086 2007 3092 2008
rect 96 1997 97 2003
rect 103 2002 1855 2003
rect 103 1998 111 2002
rect 115 1998 191 2002
rect 195 1998 215 2002
rect 219 1998 335 2002
rect 339 1998 351 2002
rect 355 1998 455 2002
rect 459 1998 519 2002
rect 523 1998 583 2002
rect 587 1998 687 2002
rect 691 1998 711 2002
rect 715 1998 831 2002
rect 835 1998 855 2002
rect 859 1998 951 2002
rect 955 1998 1015 2002
rect 1019 1998 1071 2002
rect 1075 1998 1167 2002
rect 1171 1998 1183 2002
rect 1187 1998 1287 2002
rect 1291 1998 1311 2002
rect 1315 1998 1383 2002
rect 1387 1998 1447 2002
rect 1451 1998 1479 2002
rect 1483 1998 1575 2002
rect 1579 1998 1583 2002
rect 1587 1998 1671 2002
rect 1675 1998 1719 2002
rect 1723 1998 1751 2002
rect 1755 1998 1831 2002
rect 1835 1998 1855 2002
rect 103 1997 1855 1998
rect 1861 2002 3638 2003
rect 1861 1998 1871 2002
rect 1875 1998 1959 2002
rect 1963 1998 1975 2002
rect 1979 1998 2079 2002
rect 2083 1998 2199 2002
rect 2203 1998 2223 2002
rect 2227 1998 2319 2002
rect 2323 1998 2447 2002
rect 2451 1998 2455 2002
rect 2459 1998 2583 2002
rect 2587 1998 2663 2002
rect 2667 1998 2743 2002
rect 2747 1998 2847 2002
rect 2851 1998 2919 2002
rect 2923 1998 3007 2002
rect 3011 1998 3119 2002
rect 3123 1998 3151 2002
rect 3155 1998 3279 2002
rect 3283 1998 3327 2002
rect 3331 1998 3407 2002
rect 3411 1998 3511 2002
rect 3515 1998 3591 2002
rect 3595 1998 3638 2002
rect 1861 1997 3638 1998
rect 84 1917 85 1923
rect 91 1922 1843 1923
rect 91 1918 111 1922
rect 115 1918 135 1922
rect 139 1918 183 1922
rect 187 1918 239 1922
rect 243 1918 343 1922
rect 347 1918 375 1922
rect 379 1918 511 1922
rect 515 1918 527 1922
rect 531 1918 679 1922
rect 683 1918 687 1922
rect 691 1918 847 1922
rect 851 1918 1007 1922
rect 1011 1918 1159 1922
rect 1163 1918 1303 1922
rect 1307 1918 1439 1922
rect 1443 1918 1455 1922
rect 1459 1918 1575 1922
rect 1579 1918 1607 1922
rect 1611 1918 1711 1922
rect 1715 1918 1831 1922
rect 1835 1918 1843 1922
rect 91 1917 1843 1918
rect 1849 1919 1850 1923
rect 1849 1918 3626 1919
rect 1849 1917 1871 1918
rect 1842 1914 1871 1917
rect 1875 1914 1951 1918
rect 1955 1914 2063 1918
rect 2067 1914 2071 1918
rect 2075 1914 2151 1918
rect 2155 1914 2191 1918
rect 2195 1914 2239 1918
rect 2243 1914 2311 1918
rect 2315 1914 2319 1918
rect 2323 1914 2399 1918
rect 2403 1914 2439 1918
rect 2443 1914 2487 1918
rect 2491 1914 2575 1918
rect 2579 1914 2663 1918
rect 2667 1914 2735 1918
rect 2739 1914 2759 1918
rect 2763 1914 2871 1918
rect 2875 1914 2911 1918
rect 2915 1914 2991 1918
rect 2995 1914 3111 1918
rect 3115 1914 3119 1918
rect 3123 1914 3247 1918
rect 3251 1914 3319 1918
rect 3323 1914 3383 1918
rect 3387 1914 3503 1918
rect 3507 1914 3591 1918
rect 3595 1914 3626 1918
rect 1842 1913 3626 1914
rect 96 1837 97 1843
rect 103 1842 1855 1843
rect 103 1838 111 1842
rect 115 1838 143 1842
rect 147 1838 247 1842
rect 251 1838 287 1842
rect 291 1838 383 1842
rect 387 1838 471 1842
rect 475 1838 535 1842
rect 539 1838 663 1842
rect 667 1838 695 1842
rect 699 1838 847 1842
rect 851 1838 855 1842
rect 859 1838 1015 1842
rect 1019 1838 1023 1842
rect 1027 1838 1167 1842
rect 1171 1838 1191 1842
rect 1195 1838 1311 1842
rect 1315 1838 1351 1842
rect 1355 1838 1463 1842
rect 1467 1838 1511 1842
rect 1515 1838 1615 1842
rect 1619 1838 1679 1842
rect 1683 1838 1831 1842
rect 1835 1838 1855 1842
rect 103 1837 1855 1838
rect 1861 1837 1862 1843
rect 1854 1821 1855 1827
rect 1861 1826 3631 1827
rect 1861 1822 1871 1826
rect 1875 1822 2071 1826
rect 2075 1822 2095 1826
rect 2099 1822 2159 1826
rect 2163 1822 2239 1826
rect 2243 1822 2247 1826
rect 2251 1822 2327 1826
rect 2331 1822 2399 1826
rect 2403 1822 2407 1826
rect 2411 1822 2495 1826
rect 2499 1822 2559 1826
rect 2563 1822 2583 1826
rect 2587 1822 2671 1826
rect 2675 1822 2719 1826
rect 2723 1822 2767 1826
rect 2771 1822 2879 1826
rect 2883 1822 2999 1826
rect 3003 1822 3031 1826
rect 3035 1822 3127 1826
rect 3131 1822 3175 1826
rect 3179 1822 3255 1826
rect 3259 1822 3319 1826
rect 3323 1822 3391 1826
rect 3395 1822 3471 1826
rect 3475 1822 3511 1826
rect 3515 1822 3591 1826
rect 3595 1822 3631 1826
rect 1861 1821 3631 1822
rect 3637 1821 3638 1827
rect 84 1753 85 1759
rect 91 1758 1843 1759
rect 91 1754 111 1758
rect 115 1754 135 1758
rect 139 1754 215 1758
rect 219 1754 279 1758
rect 283 1754 343 1758
rect 347 1754 463 1758
rect 467 1754 495 1758
rect 499 1754 655 1758
rect 659 1754 663 1758
rect 667 1754 839 1758
rect 843 1754 1007 1758
rect 1011 1754 1015 1758
rect 1019 1754 1167 1758
rect 1171 1754 1183 1758
rect 1187 1754 1319 1758
rect 1323 1754 1343 1758
rect 1347 1754 1463 1758
rect 1467 1754 1503 1758
rect 1507 1754 1607 1758
rect 1611 1754 1671 1758
rect 1675 1754 1743 1758
rect 1747 1754 1831 1758
rect 1835 1754 1843 1758
rect 91 1753 1843 1754
rect 1849 1753 1850 1759
rect 1842 1741 1843 1747
rect 1849 1746 3619 1747
rect 1849 1742 1871 1746
rect 1875 1742 2087 1746
rect 2091 1742 2103 1746
rect 2107 1742 2231 1746
rect 2235 1742 2239 1746
rect 2243 1742 2383 1746
rect 2387 1742 2391 1746
rect 2395 1742 2527 1746
rect 2531 1742 2551 1746
rect 2555 1742 2663 1746
rect 2667 1742 2711 1746
rect 2715 1742 2799 1746
rect 2803 1742 2871 1746
rect 2875 1742 2927 1746
rect 2931 1742 3023 1746
rect 3027 1742 3047 1746
rect 3051 1742 3159 1746
rect 3163 1742 3167 1746
rect 3171 1742 3271 1746
rect 3275 1742 3311 1746
rect 3315 1742 3391 1746
rect 3395 1742 3463 1746
rect 3467 1742 3503 1746
rect 3507 1742 3591 1746
rect 3595 1742 3619 1746
rect 1849 1741 3619 1742
rect 3625 1741 3626 1747
rect 96 1673 97 1679
rect 103 1678 1855 1679
rect 103 1674 111 1678
rect 115 1674 143 1678
rect 147 1674 223 1678
rect 227 1674 295 1678
rect 299 1674 351 1678
rect 355 1674 479 1678
rect 483 1674 503 1678
rect 507 1674 671 1678
rect 675 1674 847 1678
rect 851 1674 855 1678
rect 859 1674 1015 1678
rect 1019 1674 1031 1678
rect 1035 1674 1175 1678
rect 1179 1674 1199 1678
rect 1203 1674 1327 1678
rect 1331 1674 1359 1678
rect 1363 1674 1471 1678
rect 1475 1674 1519 1678
rect 1523 1674 1615 1678
rect 1619 1674 1679 1678
rect 1683 1674 1751 1678
rect 1755 1674 1831 1678
rect 1835 1674 1855 1678
rect 103 1673 1855 1674
rect 1861 1673 1862 1679
rect 1854 1661 1855 1667
rect 1861 1666 3631 1667
rect 1861 1662 1871 1666
rect 1875 1662 1967 1666
rect 1971 1662 2087 1666
rect 2091 1662 2111 1666
rect 2115 1662 2215 1666
rect 2219 1662 2247 1666
rect 2251 1662 2351 1666
rect 2355 1662 2391 1666
rect 2395 1662 2495 1666
rect 2499 1662 2535 1666
rect 2539 1662 2639 1666
rect 2643 1662 2671 1666
rect 2675 1662 2783 1666
rect 2787 1662 2807 1666
rect 2811 1662 2927 1666
rect 2931 1662 2935 1666
rect 2939 1662 3055 1666
rect 3059 1662 3071 1666
rect 3075 1662 3167 1666
rect 3171 1662 3223 1666
rect 3227 1662 3279 1666
rect 3283 1662 3375 1666
rect 3379 1662 3399 1666
rect 3403 1662 3511 1666
rect 3515 1662 3591 1666
rect 3595 1662 3631 1666
rect 1861 1661 3631 1662
rect 3637 1661 3638 1667
rect 84 1597 85 1603
rect 91 1602 1843 1603
rect 91 1598 111 1602
rect 115 1598 135 1602
rect 139 1598 159 1602
rect 163 1598 287 1602
rect 291 1598 423 1602
rect 427 1598 471 1602
rect 475 1598 567 1602
rect 571 1598 663 1602
rect 667 1598 711 1602
rect 715 1598 847 1602
rect 851 1598 983 1602
rect 987 1598 1023 1602
rect 1027 1598 1119 1602
rect 1123 1598 1191 1602
rect 1195 1598 1247 1602
rect 1251 1598 1351 1602
rect 1355 1598 1375 1602
rect 1379 1598 1511 1602
rect 1515 1598 1671 1602
rect 1675 1598 1831 1602
rect 1835 1598 1843 1602
rect 91 1597 1843 1598
rect 1849 1597 1850 1603
rect 1842 1577 1843 1583
rect 1849 1582 3619 1583
rect 1849 1578 1871 1582
rect 1875 1578 1895 1582
rect 1899 1578 1959 1582
rect 1963 1578 2047 1582
rect 2051 1578 2079 1582
rect 2083 1578 2207 1582
rect 2211 1578 2343 1582
rect 2347 1578 2367 1582
rect 2371 1578 2487 1582
rect 2491 1578 2527 1582
rect 2531 1578 2631 1582
rect 2635 1578 2687 1582
rect 2691 1578 2775 1582
rect 2779 1578 2839 1582
rect 2843 1578 2919 1582
rect 2923 1578 2983 1582
rect 2987 1578 3063 1582
rect 3067 1578 3119 1582
rect 3123 1578 3215 1582
rect 3219 1578 3255 1582
rect 3259 1578 3367 1582
rect 3371 1578 3391 1582
rect 3395 1578 3503 1582
rect 3507 1578 3591 1582
rect 3595 1578 3619 1582
rect 1849 1577 3619 1578
rect 3625 1577 3626 1583
rect 96 1517 97 1523
rect 103 1522 1855 1523
rect 103 1518 111 1522
rect 115 1518 167 1522
rect 171 1518 231 1522
rect 235 1518 295 1522
rect 299 1518 375 1522
rect 379 1518 431 1522
rect 435 1518 519 1522
rect 523 1518 575 1522
rect 579 1518 655 1522
rect 659 1518 719 1522
rect 723 1518 783 1522
rect 787 1518 855 1522
rect 859 1518 903 1522
rect 907 1518 991 1522
rect 995 1518 1015 1522
rect 1019 1518 1119 1522
rect 1123 1518 1127 1522
rect 1131 1518 1215 1522
rect 1219 1518 1255 1522
rect 1259 1518 1319 1522
rect 1323 1518 1383 1522
rect 1387 1518 1423 1522
rect 1427 1518 1519 1522
rect 1523 1518 1831 1522
rect 1835 1518 1855 1522
rect 103 1517 1855 1518
rect 1861 1517 1862 1523
rect 1430 1508 1436 1509
rect 1158 1504 1431 1508
rect 1435 1504 1436 1508
rect 1158 1501 1162 1504
rect 1430 1503 1436 1504
rect 1154 1500 1162 1501
rect 1154 1496 1155 1500
rect 1159 1496 1162 1500
rect 1154 1495 1160 1496
rect 1854 1493 1855 1499
rect 1861 1498 3631 1499
rect 1861 1494 1871 1498
rect 1875 1494 1903 1498
rect 1907 1494 2007 1498
rect 2011 1494 2055 1498
rect 2059 1494 2135 1498
rect 2139 1494 2215 1498
rect 2219 1494 2271 1498
rect 2275 1494 2375 1498
rect 2379 1494 2415 1498
rect 2419 1494 2535 1498
rect 2539 1494 2567 1498
rect 2571 1494 2695 1498
rect 2699 1494 2719 1498
rect 2723 1494 2847 1498
rect 2851 1494 2879 1498
rect 2883 1494 2991 1498
rect 2995 1494 3039 1498
rect 3043 1494 3127 1498
rect 3131 1494 3199 1498
rect 3203 1494 3263 1498
rect 3267 1494 3367 1498
rect 3371 1494 3399 1498
rect 3403 1494 3511 1498
rect 3515 1494 3591 1498
rect 3595 1494 3631 1498
rect 1861 1493 3631 1494
rect 3637 1493 3638 1499
rect 84 1433 85 1439
rect 91 1438 1843 1439
rect 91 1434 111 1438
rect 115 1434 223 1438
rect 227 1434 255 1438
rect 259 1434 351 1438
rect 355 1434 367 1438
rect 371 1434 447 1438
rect 451 1434 511 1438
rect 515 1434 543 1438
rect 547 1434 631 1438
rect 635 1434 647 1438
rect 651 1434 719 1438
rect 723 1434 775 1438
rect 779 1434 807 1438
rect 811 1434 895 1438
rect 899 1434 919 1438
rect 923 1434 1007 1438
rect 1011 1434 1047 1438
rect 1051 1434 1111 1438
rect 1115 1434 1207 1438
rect 1211 1434 1311 1438
rect 1315 1434 1383 1438
rect 1387 1434 1415 1438
rect 1419 1434 1575 1438
rect 1579 1434 1743 1438
rect 1747 1434 1831 1438
rect 1835 1434 1843 1438
rect 91 1433 1843 1434
rect 1849 1433 1850 1439
rect 1842 1417 1843 1423
rect 1849 1422 3619 1423
rect 1849 1418 1871 1422
rect 1875 1418 1895 1422
rect 1899 1418 1999 1422
rect 2003 1418 2023 1422
rect 2027 1418 2127 1422
rect 2131 1418 2167 1422
rect 2171 1418 2263 1422
rect 2267 1418 2303 1422
rect 2307 1418 2407 1422
rect 2411 1418 2431 1422
rect 2435 1418 2551 1422
rect 2555 1418 2559 1422
rect 2563 1418 2671 1422
rect 2675 1418 2711 1422
rect 2715 1418 2791 1422
rect 2795 1418 2871 1422
rect 2875 1418 2911 1422
rect 2915 1418 3031 1422
rect 3035 1418 3191 1422
rect 3195 1418 3359 1422
rect 3363 1418 3503 1422
rect 3507 1418 3591 1422
rect 3595 1418 3619 1422
rect 1849 1417 3619 1418
rect 3625 1417 3626 1423
rect 1242 1372 1248 1373
rect 1518 1372 1524 1373
rect 1242 1368 1243 1372
rect 1247 1368 1519 1372
rect 1523 1368 1524 1372
rect 1242 1367 1248 1368
rect 1518 1367 1524 1368
rect 96 1357 97 1363
rect 103 1362 1855 1363
rect 103 1358 111 1362
rect 115 1358 263 1362
rect 267 1358 359 1362
rect 363 1358 455 1362
rect 459 1358 471 1362
rect 475 1358 551 1362
rect 555 1358 591 1362
rect 595 1358 639 1362
rect 643 1358 727 1362
rect 731 1358 815 1362
rect 819 1358 863 1362
rect 867 1358 927 1362
rect 931 1358 1007 1362
rect 1011 1358 1055 1362
rect 1059 1358 1143 1362
rect 1147 1358 1215 1362
rect 1219 1358 1279 1362
rect 1283 1358 1391 1362
rect 1395 1358 1407 1362
rect 1411 1358 1527 1362
rect 1531 1358 1583 1362
rect 1587 1358 1647 1362
rect 1651 1358 1751 1362
rect 1755 1358 1831 1362
rect 1835 1358 1855 1362
rect 103 1357 1855 1358
rect 1861 1357 1862 1363
rect 2618 1348 2624 1349
rect 2874 1348 2880 1349
rect 2618 1344 2619 1348
rect 2623 1344 2875 1348
rect 2879 1344 2880 1348
rect 2618 1343 2624 1344
rect 2874 1343 2880 1344
rect 1854 1333 1855 1339
rect 1861 1338 3631 1339
rect 1861 1334 1871 1338
rect 1875 1334 1903 1338
rect 1907 1334 1927 1338
rect 1931 1334 2031 1338
rect 2035 1334 2047 1338
rect 2051 1334 2175 1338
rect 2179 1334 2183 1338
rect 2187 1334 2311 1338
rect 2315 1334 2319 1338
rect 2323 1334 2439 1338
rect 2443 1334 2455 1338
rect 2459 1334 2559 1338
rect 2563 1334 2591 1338
rect 2595 1334 2679 1338
rect 2683 1334 2719 1338
rect 2723 1334 2799 1338
rect 2803 1334 2839 1338
rect 2843 1334 2919 1338
rect 2923 1334 2951 1338
rect 2955 1334 3063 1338
rect 3067 1334 3183 1338
rect 3187 1334 3591 1338
rect 3595 1334 3631 1338
rect 1861 1333 3631 1334
rect 3637 1333 3638 1339
rect 1986 1324 1992 1325
rect 2326 1324 2332 1325
rect 1986 1320 1987 1324
rect 1991 1320 2327 1324
rect 2331 1320 2332 1324
rect 1986 1319 1992 1320
rect 2326 1319 2332 1320
rect 1306 1300 1312 1301
rect 1598 1300 1604 1301
rect 1306 1296 1307 1300
rect 1311 1296 1599 1300
rect 1603 1296 1604 1300
rect 1306 1295 1312 1296
rect 1598 1295 1604 1296
rect 84 1277 85 1283
rect 91 1282 1843 1283
rect 91 1278 111 1282
rect 115 1278 311 1282
rect 315 1278 351 1282
rect 355 1278 415 1282
rect 419 1278 463 1282
rect 467 1278 535 1282
rect 539 1278 583 1282
rect 587 1278 671 1282
rect 675 1278 719 1282
rect 723 1278 815 1282
rect 819 1278 855 1282
rect 859 1278 959 1282
rect 963 1278 999 1282
rect 1003 1278 1103 1282
rect 1107 1278 1135 1282
rect 1139 1278 1239 1282
rect 1243 1278 1271 1282
rect 1275 1278 1375 1282
rect 1379 1278 1399 1282
rect 1403 1278 1503 1282
rect 1507 1278 1519 1282
rect 1523 1278 1631 1282
rect 1635 1278 1639 1282
rect 1643 1278 1743 1282
rect 1747 1278 1831 1282
rect 1835 1278 1843 1282
rect 91 1277 1843 1278
rect 1849 1277 1850 1283
rect 1842 1249 1843 1255
rect 1849 1254 3619 1255
rect 1849 1250 1871 1254
rect 1875 1250 1895 1254
rect 1899 1250 1919 1254
rect 1923 1250 2039 1254
rect 2043 1250 2071 1254
rect 2075 1250 2175 1254
rect 2179 1250 2271 1254
rect 2275 1250 2311 1254
rect 2315 1250 2447 1254
rect 2451 1250 2471 1254
rect 2475 1250 2583 1254
rect 2587 1250 2663 1254
rect 2667 1250 2711 1254
rect 2715 1250 2831 1254
rect 2835 1250 2847 1254
rect 2851 1250 2943 1254
rect 2947 1250 3023 1254
rect 3027 1250 3055 1254
rect 3059 1250 3175 1254
rect 3179 1250 3191 1254
rect 3195 1250 3359 1254
rect 3363 1250 3503 1254
rect 3507 1250 3591 1254
rect 3595 1250 3619 1254
rect 1849 1249 3619 1250
rect 3625 1249 3626 1255
rect 96 1201 97 1207
rect 103 1206 1855 1207
rect 103 1202 111 1206
rect 115 1202 239 1206
rect 243 1202 319 1206
rect 323 1202 415 1206
rect 419 1202 423 1206
rect 427 1202 543 1206
rect 547 1202 591 1206
rect 595 1202 679 1206
rect 683 1202 759 1206
rect 763 1202 823 1206
rect 827 1202 927 1206
rect 931 1202 967 1206
rect 971 1202 1079 1206
rect 1083 1202 1111 1206
rect 1115 1202 1223 1206
rect 1227 1202 1247 1206
rect 1251 1202 1367 1206
rect 1371 1202 1383 1206
rect 1387 1202 1503 1206
rect 1507 1202 1511 1206
rect 1515 1202 1639 1206
rect 1643 1202 1751 1206
rect 1755 1202 1831 1206
rect 1835 1202 1855 1206
rect 103 1201 1855 1202
rect 1861 1201 1862 1207
rect 2506 1188 2512 1189
rect 2778 1188 2784 1189
rect 2506 1184 2507 1188
rect 2511 1184 2779 1188
rect 2783 1184 2784 1188
rect 2506 1183 2512 1184
rect 2778 1183 2784 1184
rect 1854 1169 1855 1175
rect 1861 1174 3631 1175
rect 1861 1170 1871 1174
rect 1875 1170 1903 1174
rect 1907 1170 1983 1174
rect 1987 1170 2079 1174
rect 2083 1170 2087 1174
rect 2091 1170 2215 1174
rect 2219 1170 2279 1174
rect 2283 1170 2367 1174
rect 2371 1170 2479 1174
rect 2483 1170 2527 1174
rect 2531 1170 2671 1174
rect 2675 1170 2687 1174
rect 2691 1170 2839 1174
rect 2843 1170 2855 1174
rect 2859 1170 2983 1174
rect 2987 1170 3031 1174
rect 3035 1170 3127 1174
rect 3131 1170 3199 1174
rect 3203 1170 3263 1174
rect 3267 1170 3367 1174
rect 3371 1170 3399 1174
rect 3403 1170 3511 1174
rect 3515 1170 3591 1174
rect 3595 1170 3631 1174
rect 1861 1169 3631 1170
rect 3637 1169 3638 1175
rect 84 1121 85 1127
rect 91 1126 1843 1127
rect 91 1122 111 1126
rect 115 1122 143 1126
rect 147 1122 231 1126
rect 235 1122 279 1126
rect 283 1122 407 1126
rect 411 1122 423 1126
rect 427 1122 567 1126
rect 571 1122 583 1126
rect 587 1122 711 1126
rect 715 1122 751 1126
rect 755 1122 847 1126
rect 851 1122 919 1126
rect 923 1122 975 1126
rect 979 1122 1071 1126
rect 1075 1122 1103 1126
rect 1107 1122 1215 1126
rect 1219 1122 1223 1126
rect 1227 1122 1343 1126
rect 1347 1122 1359 1126
rect 1363 1122 1471 1126
rect 1475 1122 1495 1126
rect 1499 1122 1631 1126
rect 1635 1122 1743 1126
rect 1747 1122 1831 1126
rect 1835 1122 1843 1126
rect 91 1121 1843 1122
rect 1849 1121 1850 1127
rect 1842 1085 1843 1091
rect 1849 1090 3619 1091
rect 1849 1086 1871 1090
rect 1875 1086 1895 1090
rect 1899 1086 1975 1090
rect 1979 1086 2079 1090
rect 2083 1086 2167 1090
rect 2171 1086 2207 1090
rect 2211 1086 2255 1090
rect 2259 1086 2359 1090
rect 2363 1086 2479 1090
rect 2483 1086 2519 1090
rect 2523 1086 2607 1090
rect 2611 1086 2679 1090
rect 2683 1086 2751 1090
rect 2755 1086 2831 1090
rect 2835 1086 2895 1090
rect 2899 1086 2975 1090
rect 2979 1086 3047 1090
rect 3051 1086 3119 1090
rect 3123 1086 3207 1090
rect 3211 1086 3255 1090
rect 3259 1086 3367 1090
rect 3371 1086 3391 1090
rect 3395 1086 3503 1090
rect 3507 1086 3591 1090
rect 3595 1086 3619 1090
rect 1849 1085 3619 1086
rect 3625 1085 3626 1091
rect 1054 1052 1060 1053
rect 1366 1052 1372 1053
rect 1054 1048 1055 1052
rect 1059 1048 1367 1052
rect 1371 1048 1372 1052
rect 1054 1047 1060 1048
rect 1366 1047 1372 1048
rect 96 1037 97 1043
rect 103 1042 1855 1043
rect 103 1038 111 1042
rect 115 1038 143 1042
rect 147 1038 151 1042
rect 155 1038 263 1042
rect 267 1038 287 1042
rect 291 1038 407 1042
rect 411 1038 431 1042
rect 435 1038 551 1042
rect 555 1038 575 1042
rect 579 1038 687 1042
rect 691 1038 719 1042
rect 723 1038 807 1042
rect 811 1038 855 1042
rect 859 1038 927 1042
rect 931 1038 983 1042
rect 987 1038 1039 1042
rect 1043 1038 1111 1042
rect 1115 1038 1143 1042
rect 1147 1038 1231 1042
rect 1235 1038 1247 1042
rect 1251 1038 1351 1042
rect 1355 1038 1359 1042
rect 1363 1038 1479 1042
rect 1483 1038 1831 1042
rect 1835 1038 1855 1042
rect 103 1037 1855 1038
rect 1861 1037 1862 1043
rect 2346 1028 2352 1029
rect 2562 1028 2568 1029
rect 2346 1024 2347 1028
rect 2351 1024 2563 1028
rect 2567 1024 2568 1028
rect 2346 1023 2352 1024
rect 2562 1023 2568 1024
rect 1854 1009 1855 1015
rect 1861 1014 3631 1015
rect 1861 1010 1871 1014
rect 1875 1010 2175 1014
rect 2179 1010 2263 1014
rect 2267 1010 2303 1014
rect 2307 1010 2367 1014
rect 2371 1010 2383 1014
rect 2387 1010 2471 1014
rect 2475 1010 2487 1014
rect 2491 1010 2567 1014
rect 2571 1010 2615 1014
rect 2619 1010 2671 1014
rect 2675 1010 2759 1014
rect 2763 1010 2783 1014
rect 2787 1010 2903 1014
rect 2907 1010 2911 1014
rect 2915 1010 3055 1014
rect 3059 1010 3207 1014
rect 3211 1010 3215 1014
rect 3219 1010 3367 1014
rect 3371 1010 3375 1014
rect 3379 1010 3511 1014
rect 3515 1010 3591 1014
rect 3595 1010 3631 1014
rect 1861 1009 3631 1010
rect 3637 1009 3638 1015
rect 84 953 85 959
rect 91 958 1843 959
rect 91 954 111 958
rect 115 954 135 958
rect 139 954 215 958
rect 219 954 255 958
rect 259 954 327 958
rect 331 954 399 958
rect 403 954 447 958
rect 451 954 543 958
rect 547 954 567 958
rect 571 954 679 958
rect 683 954 687 958
rect 691 954 799 958
rect 803 954 911 958
rect 915 954 919 958
rect 923 954 1015 958
rect 1019 954 1031 958
rect 1035 954 1119 958
rect 1123 954 1135 958
rect 1139 954 1223 958
rect 1227 954 1239 958
rect 1243 954 1327 958
rect 1331 954 1351 958
rect 1355 954 1831 958
rect 1835 954 1843 958
rect 91 953 1843 954
rect 1849 953 1850 959
rect 1842 925 1843 931
rect 1849 930 3619 931
rect 1849 926 1871 930
rect 1875 926 2279 930
rect 2283 926 2295 930
rect 2299 926 2359 930
rect 2363 926 2375 930
rect 2379 926 2439 930
rect 2443 926 2463 930
rect 2467 926 2519 930
rect 2523 926 2559 930
rect 2563 926 2607 930
rect 2611 926 2663 930
rect 2667 926 2703 930
rect 2707 926 2775 930
rect 2779 926 2807 930
rect 2811 926 2903 930
rect 2907 926 2911 930
rect 2915 926 3015 930
rect 3019 926 3047 930
rect 3051 926 3111 930
rect 3115 926 3199 930
rect 3203 926 3215 930
rect 3219 926 3319 930
rect 3323 926 3359 930
rect 3363 926 3423 930
rect 3427 926 3503 930
rect 3507 926 3591 930
rect 3595 926 3619 930
rect 1849 925 3619 926
rect 3625 925 3626 931
rect 96 869 97 875
rect 103 874 1855 875
rect 103 870 111 874
rect 115 870 143 874
rect 147 870 223 874
rect 227 870 255 874
rect 259 870 335 874
rect 339 870 399 874
rect 403 870 455 874
rect 459 870 559 874
rect 563 870 575 874
rect 579 870 695 874
rect 699 870 719 874
rect 723 870 807 874
rect 811 870 871 874
rect 875 870 919 874
rect 923 870 1015 874
rect 1019 870 1023 874
rect 1027 870 1127 874
rect 1131 870 1151 874
rect 1155 870 1231 874
rect 1235 870 1279 874
rect 1283 870 1335 874
rect 1339 870 1399 874
rect 1403 870 1519 874
rect 1523 870 1647 874
rect 1651 870 1831 874
rect 1835 870 1855 874
rect 103 869 1855 870
rect 1861 869 1862 875
rect 1854 837 1855 843
rect 1861 842 3631 843
rect 1861 838 1871 842
rect 1875 838 2167 842
rect 2171 838 2247 842
rect 2251 838 2287 842
rect 2291 838 2327 842
rect 2331 838 2367 842
rect 2371 838 2423 842
rect 2427 838 2447 842
rect 2451 838 2527 842
rect 2531 838 2535 842
rect 2539 838 2615 842
rect 2619 838 2655 842
rect 2659 838 2711 842
rect 2715 838 2783 842
rect 2787 838 2815 842
rect 2819 838 2911 842
rect 2915 838 2919 842
rect 2923 838 3023 842
rect 3027 838 3039 842
rect 3043 838 3119 842
rect 3123 838 3159 842
rect 3163 838 3223 842
rect 3227 838 3279 842
rect 3283 838 3327 842
rect 3331 838 3407 842
rect 3411 838 3431 842
rect 3435 838 3511 842
rect 3515 838 3591 842
rect 3595 838 3631 842
rect 1861 837 3631 838
rect 3637 837 3638 843
rect 84 781 85 787
rect 91 786 1843 787
rect 91 782 111 786
rect 115 782 135 786
rect 139 782 247 786
rect 251 782 263 786
rect 267 782 391 786
rect 395 782 431 786
rect 435 782 551 786
rect 555 782 607 786
rect 611 782 711 786
rect 715 782 783 786
rect 787 782 863 786
rect 867 782 951 786
rect 955 782 1007 786
rect 1011 782 1103 786
rect 1107 782 1143 786
rect 1147 782 1247 786
rect 1251 782 1271 786
rect 1275 782 1383 786
rect 1387 782 1391 786
rect 1395 782 1511 786
rect 1515 782 1639 786
rect 1643 782 1743 786
rect 1747 782 1831 786
rect 1835 782 1843 786
rect 91 781 1843 782
rect 1849 781 1850 787
rect 1842 753 1843 759
rect 1849 758 3619 759
rect 1849 754 1871 758
rect 1875 754 1895 758
rect 1899 754 1975 758
rect 1979 754 2071 758
rect 2075 754 2159 758
rect 2163 754 2183 758
rect 2187 754 2239 758
rect 2243 754 2311 758
rect 2315 754 2319 758
rect 2323 754 2415 758
rect 2419 754 2447 758
rect 2451 754 2527 758
rect 2531 754 2591 758
rect 2595 754 2647 758
rect 2651 754 2743 758
rect 2747 754 2775 758
rect 2779 754 2895 758
rect 2899 754 2903 758
rect 2907 754 3031 758
rect 3035 754 3047 758
rect 3051 754 3151 758
rect 3155 754 3199 758
rect 3203 754 3271 758
rect 3275 754 3359 758
rect 3363 754 3399 758
rect 3403 754 3503 758
rect 3507 754 3591 758
rect 3595 754 3619 758
rect 1849 753 3619 754
rect 3625 753 3626 759
rect 96 693 97 699
rect 103 698 1855 699
rect 103 694 111 698
rect 115 694 143 698
rect 147 694 271 698
rect 275 694 295 698
rect 299 694 407 698
rect 411 694 439 698
rect 443 694 527 698
rect 531 694 615 698
rect 619 694 655 698
rect 659 694 783 698
rect 787 694 791 698
rect 795 694 903 698
rect 907 694 959 698
rect 963 694 1023 698
rect 1027 694 1111 698
rect 1115 694 1135 698
rect 1139 694 1247 698
rect 1251 694 1255 698
rect 1259 694 1351 698
rect 1355 694 1391 698
rect 1395 694 1455 698
rect 1459 694 1519 698
rect 1523 694 1559 698
rect 1563 694 1647 698
rect 1651 694 1663 698
rect 1667 694 1751 698
rect 1755 694 1831 698
rect 1835 694 1855 698
rect 103 693 1855 694
rect 1861 693 1862 699
rect 1198 684 1204 685
rect 1566 684 1572 685
rect 1198 680 1199 684
rect 1203 680 1567 684
rect 1571 680 1572 684
rect 1198 679 1204 680
rect 1566 679 1572 680
rect 1854 673 1855 679
rect 1861 678 3631 679
rect 1861 674 1871 678
rect 1875 674 1903 678
rect 1907 674 1983 678
rect 1987 674 2079 678
rect 2083 674 2095 678
rect 2099 674 2191 678
rect 2195 674 2295 678
rect 2299 674 2319 678
rect 2323 674 2455 678
rect 2459 674 2479 678
rect 2483 674 2599 678
rect 2603 674 2655 678
rect 2659 674 2751 678
rect 2755 674 2831 678
rect 2835 674 2903 678
rect 2907 674 3007 678
rect 3011 674 3055 678
rect 3059 674 3183 678
rect 3187 674 3207 678
rect 3211 674 3359 678
rect 3363 674 3367 678
rect 3371 674 3511 678
rect 3515 674 3591 678
rect 3595 674 3631 678
rect 1861 673 3631 674
rect 3637 673 3638 679
rect 1706 660 1712 661
rect 2302 660 2308 661
rect 1706 656 1707 660
rect 1711 656 2303 660
rect 2307 656 2308 660
rect 1706 655 1712 656
rect 2302 655 2308 656
rect 84 613 85 619
rect 91 618 1843 619
rect 91 614 111 618
rect 115 614 287 618
rect 291 614 311 618
rect 315 614 391 618
rect 395 614 399 618
rect 403 614 471 618
rect 475 614 519 618
rect 523 614 559 618
rect 563 614 647 618
rect 651 614 735 618
rect 739 614 775 618
rect 779 614 823 618
rect 827 614 895 618
rect 899 614 911 618
rect 915 614 999 618
rect 1003 614 1015 618
rect 1019 614 1087 618
rect 1091 614 1127 618
rect 1131 614 1175 618
rect 1179 614 1239 618
rect 1243 614 1263 618
rect 1267 614 1343 618
rect 1347 614 1447 618
rect 1451 614 1551 618
rect 1555 614 1655 618
rect 1659 614 1743 618
rect 1747 614 1831 618
rect 1835 614 1843 618
rect 91 613 1843 614
rect 1849 613 1850 619
rect 1842 593 1843 599
rect 1849 598 3619 599
rect 1849 594 1871 598
rect 1875 594 1895 598
rect 1899 594 1975 598
rect 1979 594 2087 598
rect 2091 594 2215 598
rect 2219 594 2287 598
rect 2291 594 2351 598
rect 2355 594 2471 598
rect 2475 594 2495 598
rect 2499 594 2647 598
rect 2651 594 2807 598
rect 2811 594 2823 598
rect 2827 594 2975 598
rect 2979 594 2999 598
rect 3003 594 3151 598
rect 3155 594 3175 598
rect 3179 594 3335 598
rect 3339 594 3351 598
rect 3355 594 3503 598
rect 3507 594 3591 598
rect 3595 594 3619 598
rect 1849 593 3619 594
rect 3625 593 3626 599
rect 2178 540 2184 541
rect 2450 540 2456 541
rect 2178 536 2179 540
rect 2183 536 2451 540
rect 2455 536 2456 540
rect 2178 535 2184 536
rect 2450 535 2456 536
rect 96 525 97 531
rect 103 530 1855 531
rect 103 526 111 530
rect 115 526 239 530
rect 243 526 319 530
rect 323 526 343 530
rect 347 526 399 530
rect 403 526 439 530
rect 443 526 479 530
rect 483 526 535 530
rect 539 526 567 530
rect 571 526 631 530
rect 635 526 655 530
rect 659 526 719 530
rect 723 526 743 530
rect 747 526 807 530
rect 811 526 831 530
rect 835 526 895 530
rect 899 526 919 530
rect 923 526 983 530
rect 987 526 1007 530
rect 1011 526 1071 530
rect 1075 526 1095 530
rect 1099 526 1159 530
rect 1163 526 1183 530
rect 1187 526 1247 530
rect 1251 526 1271 530
rect 1275 526 1831 530
rect 1835 526 1855 530
rect 103 525 1855 526
rect 1861 525 1862 531
rect 1854 523 1862 525
rect 1854 517 1855 523
rect 1861 522 3631 523
rect 1861 518 1871 522
rect 1875 518 1903 522
rect 1907 518 1983 522
rect 1987 518 2095 522
rect 2099 518 2151 522
rect 2155 518 2223 522
rect 2227 518 2231 522
rect 2235 518 2327 522
rect 2331 518 2359 522
rect 2363 518 2431 522
rect 2435 518 2503 522
rect 2507 518 2551 522
rect 2555 518 2655 522
rect 2659 518 2687 522
rect 2691 518 2815 522
rect 2819 518 2839 522
rect 2843 518 2983 522
rect 2987 518 2999 522
rect 3003 518 3159 522
rect 3163 518 3175 522
rect 3179 518 3343 522
rect 3347 518 3351 522
rect 3355 518 3511 522
rect 3515 518 3591 522
rect 3595 518 3631 522
rect 1861 517 3631 518
rect 3637 517 3638 523
rect 882 516 888 517
rect 1254 516 1260 517
rect 882 512 883 516
rect 887 512 1255 516
rect 1259 512 1260 516
rect 882 511 888 512
rect 1254 511 1260 512
rect 84 441 85 447
rect 91 446 1843 447
rect 91 442 111 446
rect 115 442 135 446
rect 139 442 231 446
rect 235 442 247 446
rect 251 442 335 446
rect 339 442 375 446
rect 379 442 431 446
rect 435 442 495 446
rect 499 442 527 446
rect 531 442 607 446
rect 611 442 623 446
rect 627 442 711 446
rect 715 442 719 446
rect 723 442 799 446
rect 803 442 823 446
rect 827 442 887 446
rect 891 442 919 446
rect 923 442 975 446
rect 979 442 1007 446
rect 1011 442 1063 446
rect 1067 442 1103 446
rect 1107 442 1151 446
rect 1155 442 1199 446
rect 1203 442 1239 446
rect 1243 442 1295 446
rect 1299 442 1831 446
rect 1835 442 1843 446
rect 91 441 1843 442
rect 1849 443 1850 447
rect 1849 442 3626 443
rect 1849 441 1871 442
rect 1842 438 1871 441
rect 1875 438 2143 442
rect 2147 438 2223 442
rect 2227 438 2319 442
rect 2323 438 2335 442
rect 2339 438 2415 442
rect 2419 438 2423 442
rect 2427 438 2495 442
rect 2499 438 2543 442
rect 2547 438 2583 442
rect 2587 438 2679 442
rect 2683 438 2687 442
rect 2691 438 2799 442
rect 2803 438 2831 442
rect 2835 438 2927 442
rect 2931 438 2991 442
rect 2995 438 3071 442
rect 3075 438 3167 442
rect 3171 438 3215 442
rect 3219 438 3343 442
rect 3347 438 3367 442
rect 3371 438 3503 442
rect 3507 438 3591 442
rect 3595 438 3626 442
rect 1842 437 3626 438
rect 96 353 97 359
rect 103 358 1855 359
rect 103 354 111 358
rect 115 354 143 358
rect 147 354 247 358
rect 251 354 255 358
rect 259 354 375 358
rect 379 354 383 358
rect 387 354 503 358
rect 507 354 511 358
rect 515 354 615 358
rect 619 354 647 358
rect 651 354 727 358
rect 731 354 775 358
rect 779 354 831 358
rect 835 354 895 358
rect 899 354 927 358
rect 931 354 1007 358
rect 1011 354 1015 358
rect 1019 354 1111 358
rect 1115 354 1119 358
rect 1123 354 1207 358
rect 1211 354 1223 358
rect 1227 354 1303 358
rect 1307 354 1327 358
rect 1331 354 1439 358
rect 1443 354 1831 358
rect 1835 354 1855 358
rect 103 353 1855 354
rect 1861 358 3638 359
rect 1861 354 1871 358
rect 1875 354 2079 358
rect 2083 354 2167 358
rect 2171 354 2263 358
rect 2267 354 2343 358
rect 2347 354 2375 358
rect 2379 354 2423 358
rect 2427 354 2503 358
rect 2507 354 2591 358
rect 2595 354 2639 358
rect 2643 354 2695 358
rect 2699 354 2775 358
rect 2779 354 2807 358
rect 2811 354 2911 358
rect 2915 354 2935 358
rect 2939 354 3039 358
rect 3043 354 3079 358
rect 3083 354 3167 358
rect 3171 354 3223 358
rect 3227 354 3287 358
rect 3291 354 3375 358
rect 3379 354 3407 358
rect 3411 354 3511 358
rect 3515 354 3591 358
rect 3595 354 3638 358
rect 1861 353 3638 354
rect 84 269 85 275
rect 91 274 1843 275
rect 91 270 111 274
rect 115 270 135 274
rect 139 270 223 274
rect 227 270 239 274
rect 243 270 335 274
rect 339 270 367 274
rect 371 270 463 274
rect 467 270 503 274
rect 507 270 599 274
rect 603 270 639 274
rect 643 270 735 274
rect 739 270 767 274
rect 771 270 871 274
rect 875 270 887 274
rect 891 270 999 274
rect 1003 270 1007 274
rect 1011 270 1111 274
rect 1115 270 1135 274
rect 1139 270 1215 274
rect 1219 270 1255 274
rect 1259 270 1319 274
rect 1323 270 1367 274
rect 1371 270 1431 274
rect 1435 270 1479 274
rect 1483 270 1599 274
rect 1603 270 1831 274
rect 1835 270 1843 274
rect 91 269 1843 270
rect 1849 274 3626 275
rect 1849 270 1871 274
rect 1875 270 1895 274
rect 1899 270 1983 274
rect 1987 270 2071 274
rect 2075 270 2095 274
rect 2099 270 2159 274
rect 2163 270 2223 274
rect 2227 270 2255 274
rect 2259 270 2359 274
rect 2363 270 2367 274
rect 2371 270 2495 274
rect 2499 270 2503 274
rect 2507 270 2631 274
rect 2635 270 2647 274
rect 2651 270 2767 274
rect 2771 270 2791 274
rect 2795 270 2903 274
rect 2907 270 2935 274
rect 2939 270 3031 274
rect 3035 270 3079 274
rect 3083 270 3159 274
rect 3163 270 3223 274
rect 3227 270 3279 274
rect 3283 270 3375 274
rect 3379 270 3399 274
rect 3403 270 3503 274
rect 3507 270 3591 274
rect 3595 270 3626 274
rect 1849 269 3626 270
rect 1042 212 1048 213
rect 1570 212 1576 213
rect 1042 208 1043 212
rect 1047 208 1571 212
rect 1575 208 1576 212
rect 1042 207 1048 208
rect 1570 207 1576 208
rect 1930 212 1936 213
rect 2458 212 2464 213
rect 1930 208 1931 212
rect 1935 208 2459 212
rect 2463 208 2464 212
rect 1930 207 1936 208
rect 2458 207 2464 208
rect 1854 181 1855 187
rect 1861 186 3631 187
rect 1861 182 1871 186
rect 1875 182 1903 186
rect 1907 182 1983 186
rect 1987 182 1991 186
rect 1995 182 2087 186
rect 2091 182 2103 186
rect 2107 182 2207 186
rect 2211 182 2231 186
rect 2235 182 2335 186
rect 2339 182 2367 186
rect 2371 182 2463 186
rect 2467 182 2511 186
rect 2515 182 2583 186
rect 2587 182 2655 186
rect 2659 182 2703 186
rect 2707 182 2799 186
rect 2803 182 2815 186
rect 2819 182 2919 186
rect 2923 182 2943 186
rect 2947 182 3015 186
rect 3019 182 3087 186
rect 3091 182 3111 186
rect 3115 182 3207 186
rect 3211 182 3231 186
rect 3235 182 3303 186
rect 3307 182 3383 186
rect 3387 182 3399 186
rect 3403 182 3511 186
rect 3515 182 3591 186
rect 3595 182 3631 186
rect 1861 181 3631 182
rect 3637 181 3638 187
rect 2154 172 2160 173
rect 2470 172 2476 173
rect 2154 168 2155 172
rect 2159 168 2471 172
rect 2475 168 2476 172
rect 2154 167 2160 168
rect 2470 167 2476 168
rect 96 161 97 167
rect 103 166 1855 167
rect 103 162 111 166
rect 115 162 159 166
rect 163 162 231 166
rect 235 162 239 166
rect 243 162 319 166
rect 323 162 343 166
rect 347 162 399 166
rect 403 162 471 166
rect 475 162 479 166
rect 483 162 559 166
rect 563 162 607 166
rect 611 162 647 166
rect 651 162 735 166
rect 739 162 743 166
rect 747 162 823 166
rect 827 162 879 166
rect 883 162 911 166
rect 915 162 999 166
rect 1003 162 1015 166
rect 1019 162 1087 166
rect 1091 162 1143 166
rect 1147 162 1167 166
rect 1171 162 1247 166
rect 1251 162 1263 166
rect 1267 162 1335 166
rect 1339 162 1375 166
rect 1379 162 1423 166
rect 1427 162 1487 166
rect 1491 162 1511 166
rect 1515 162 1591 166
rect 1595 162 1607 166
rect 1611 162 1671 166
rect 1675 162 1751 166
rect 1755 162 1831 166
rect 1835 162 1855 166
rect 103 161 1855 162
rect 1861 161 1862 167
rect 1842 105 1843 111
rect 1849 110 3619 111
rect 1849 106 1871 110
rect 1875 106 1895 110
rect 1899 106 1975 110
rect 1979 106 2079 110
rect 2083 106 2199 110
rect 2203 106 2327 110
rect 2331 106 2455 110
rect 2459 106 2575 110
rect 2579 106 2695 110
rect 2699 106 2807 110
rect 2811 106 2911 110
rect 2915 106 3007 110
rect 3011 106 3103 110
rect 3107 106 3199 110
rect 3203 106 3295 110
rect 3299 106 3391 110
rect 3395 106 3591 110
rect 3595 106 3619 110
rect 1849 105 3619 106
rect 3625 105 3626 111
rect 84 85 85 91
rect 91 90 1843 91
rect 91 86 111 90
rect 115 86 151 90
rect 155 86 231 90
rect 235 86 311 90
rect 315 86 391 90
rect 395 86 471 90
rect 475 86 551 90
rect 555 86 639 90
rect 643 86 727 90
rect 731 86 815 90
rect 819 86 903 90
rect 907 86 991 90
rect 995 86 1079 90
rect 1083 86 1159 90
rect 1163 86 1239 90
rect 1243 86 1327 90
rect 1331 86 1415 90
rect 1419 86 1503 90
rect 1507 86 1583 90
rect 1587 86 1663 90
rect 1667 86 1743 90
rect 1747 86 1831 90
rect 1835 86 1843 90
rect 91 85 1843 86
rect 1849 85 1850 91
<< m5c >>
rect 1843 3665 1849 3671
rect 3619 3665 3625 3671
rect 97 3637 103 3643
rect 1855 3637 1861 3643
rect 1855 3589 1861 3595
rect 3631 3589 3637 3595
rect 85 3561 91 3567
rect 1843 3561 1849 3567
rect 1843 3513 1849 3519
rect 3619 3513 3625 3519
rect 97 3477 103 3483
rect 1855 3477 1861 3483
rect 1855 3437 1861 3443
rect 3631 3437 3637 3443
rect 85 3397 91 3403
rect 1843 3397 1849 3403
rect 1843 3361 1849 3367
rect 3619 3361 3625 3367
rect 97 3317 103 3323
rect 1855 3317 1861 3323
rect 1855 3285 1861 3291
rect 3631 3285 3637 3291
rect 85 3241 91 3247
rect 1843 3241 1849 3247
rect 1843 3209 1849 3215
rect 3619 3209 3625 3215
rect 1583 3196 1589 3197
rect 1583 3192 1587 3196
rect 1587 3192 1589 3196
rect 1583 3191 1589 3192
rect 911 3172 917 3173
rect 911 3168 915 3172
rect 915 3168 917 3172
rect 911 3167 917 3168
rect 97 3157 103 3163
rect 1855 3157 1861 3163
rect 1855 3133 1861 3139
rect 3631 3133 3637 3139
rect 85 3069 91 3075
rect 1843 3069 1849 3075
rect 1843 3045 1849 3051
rect 3619 3045 3625 3051
rect 97 2981 103 2987
rect 1855 2981 1861 2987
rect 1855 2957 1861 2963
rect 3631 2957 3637 2963
rect 85 2905 91 2911
rect 1843 2905 1849 2911
rect 1843 2881 1849 2887
rect 3619 2881 3625 2887
rect 97 2825 103 2831
rect 1855 2825 1861 2831
rect 1855 2793 1861 2799
rect 3631 2793 3637 2799
rect 85 2745 91 2751
rect 1843 2745 1849 2751
rect 1843 2717 1849 2723
rect 3619 2717 3625 2723
rect 97 2661 103 2667
rect 1855 2661 1861 2667
rect 1855 2633 1861 2639
rect 3631 2633 3637 2639
rect 85 2581 91 2587
rect 1843 2581 1849 2587
rect 1843 2557 1849 2563
rect 3619 2557 3625 2563
rect 97 2501 103 2507
rect 1855 2501 1861 2507
rect 1855 2473 1861 2479
rect 3631 2473 3637 2479
rect 85 2413 91 2419
rect 1843 2413 1849 2419
rect 1843 2393 1849 2399
rect 3619 2393 3625 2399
rect 97 2329 103 2335
rect 1855 2329 1861 2335
rect 1855 2313 1861 2319
rect 3631 2313 3637 2319
rect 85 2253 91 2259
rect 1843 2253 1849 2259
rect 1843 2237 1849 2243
rect 3619 2237 3625 2243
rect 97 2165 103 2171
rect 1855 2165 1861 2171
rect 1855 2157 1861 2163
rect 3631 2157 3637 2163
rect 85 2077 91 2083
rect 1843 2077 1849 2083
rect 97 1997 103 2003
rect 1855 1997 1861 2003
rect 85 1917 91 1923
rect 1843 1917 1849 1923
rect 97 1837 103 1843
rect 1855 1837 1861 1843
rect 1855 1821 1861 1827
rect 3631 1821 3637 1827
rect 85 1753 91 1759
rect 1843 1753 1849 1759
rect 1843 1741 1849 1747
rect 3619 1741 3625 1747
rect 97 1673 103 1679
rect 1855 1673 1861 1679
rect 1855 1661 1861 1667
rect 3631 1661 3637 1667
rect 85 1597 91 1603
rect 1843 1597 1849 1603
rect 1843 1577 1849 1583
rect 3619 1577 3625 1583
rect 97 1517 103 1523
rect 1855 1517 1861 1523
rect 1855 1493 1861 1499
rect 3631 1493 3637 1499
rect 85 1433 91 1439
rect 1843 1433 1849 1439
rect 1843 1417 1849 1423
rect 3619 1417 3625 1423
rect 97 1357 103 1363
rect 1855 1357 1861 1363
rect 1855 1333 1861 1339
rect 3631 1333 3637 1339
rect 85 1277 91 1283
rect 1843 1277 1849 1283
rect 1843 1249 1849 1255
rect 3619 1249 3625 1255
rect 97 1201 103 1207
rect 1855 1201 1861 1207
rect 1855 1169 1861 1175
rect 3631 1169 3637 1175
rect 85 1121 91 1127
rect 1843 1121 1849 1127
rect 1843 1085 1849 1091
rect 3619 1085 3625 1091
rect 97 1037 103 1043
rect 1855 1037 1861 1043
rect 1855 1009 1861 1015
rect 3631 1009 3637 1015
rect 85 953 91 959
rect 1843 953 1849 959
rect 1843 925 1849 931
rect 3619 925 3625 931
rect 97 869 103 875
rect 1855 869 1861 875
rect 1855 837 1861 843
rect 3631 837 3637 843
rect 85 781 91 787
rect 1843 781 1849 787
rect 1843 753 1849 759
rect 3619 753 3625 759
rect 97 693 103 699
rect 1855 693 1861 699
rect 1855 673 1861 679
rect 3631 673 3637 679
rect 85 613 91 619
rect 1843 613 1849 619
rect 1843 593 1849 599
rect 3619 593 3625 599
rect 97 525 103 531
rect 1855 525 1861 531
rect 1855 517 1861 523
rect 3631 517 3637 523
rect 85 441 91 447
rect 1843 441 1849 447
rect 97 353 103 359
rect 1855 353 1861 359
rect 85 269 91 275
rect 1843 269 1849 275
rect 1855 181 1861 187
rect 3631 181 3637 187
rect 97 161 103 167
rect 1855 161 1861 167
rect 1843 105 1849 111
rect 3619 105 3625 111
rect 85 85 91 91
rect 1843 85 1849 91
<< m5 >>
rect 84 3567 92 3672
rect 84 3561 85 3567
rect 91 3561 92 3567
rect 84 3403 92 3561
rect 84 3397 85 3403
rect 91 3397 92 3403
rect 84 3247 92 3397
rect 84 3241 85 3247
rect 91 3241 92 3247
rect 84 3075 92 3241
rect 84 3069 85 3075
rect 91 3069 92 3075
rect 84 2911 92 3069
rect 84 2905 85 2911
rect 91 2905 92 2911
rect 84 2751 92 2905
rect 84 2745 85 2751
rect 91 2745 92 2751
rect 84 2587 92 2745
rect 84 2581 85 2587
rect 91 2581 92 2587
rect 84 2419 92 2581
rect 84 2413 85 2419
rect 91 2413 92 2419
rect 84 2259 92 2413
rect 84 2253 85 2259
rect 91 2253 92 2259
rect 84 2083 92 2253
rect 84 2077 85 2083
rect 91 2077 92 2083
rect 84 1923 92 2077
rect 84 1917 85 1923
rect 91 1917 92 1923
rect 84 1759 92 1917
rect 84 1753 85 1759
rect 91 1753 92 1759
rect 84 1603 92 1753
rect 84 1597 85 1603
rect 91 1597 92 1603
rect 84 1439 92 1597
rect 84 1433 85 1439
rect 91 1433 92 1439
rect 84 1283 92 1433
rect 84 1277 85 1283
rect 91 1277 92 1283
rect 84 1127 92 1277
rect 84 1121 85 1127
rect 91 1121 92 1127
rect 84 959 92 1121
rect 84 953 85 959
rect 91 953 92 959
rect 84 787 92 953
rect 84 781 85 787
rect 91 781 92 787
rect 84 619 92 781
rect 84 613 85 619
rect 91 613 92 619
rect 84 447 92 613
rect 84 441 85 447
rect 91 441 92 447
rect 84 275 92 441
rect 84 269 85 275
rect 91 269 92 275
rect 84 91 92 269
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 3643 104 3672
rect 96 3637 97 3643
rect 103 3637 104 3643
rect 96 3483 104 3637
rect 96 3477 97 3483
rect 103 3477 104 3483
rect 96 3323 104 3477
rect 96 3317 97 3323
rect 103 3317 104 3323
rect 96 3163 104 3317
rect 1842 3671 1850 3672
rect 1842 3665 1843 3671
rect 1849 3665 1850 3671
rect 1842 3567 1850 3665
rect 1842 3561 1843 3567
rect 1849 3561 1850 3567
rect 1842 3519 1850 3561
rect 1842 3513 1843 3519
rect 1849 3513 1850 3519
rect 1842 3403 1850 3513
rect 1842 3397 1843 3403
rect 1849 3397 1850 3403
rect 1842 3367 1850 3397
rect 1842 3361 1843 3367
rect 1849 3361 1850 3367
rect 1842 3247 1850 3361
rect 1842 3241 1843 3247
rect 1849 3241 1850 3247
rect 1842 3215 1850 3241
rect 1842 3209 1843 3215
rect 1849 3209 1850 3215
rect 1582 3197 1590 3198
rect 1582 3191 1583 3197
rect 1589 3191 1590 3197
rect 1582 3190 1590 3191
rect 910 3173 918 3174
rect 910 3171 911 3173
rect 917 3171 918 3173
rect 1584 3171 1588 3190
rect 96 3157 97 3163
rect 103 3157 104 3163
rect 96 2987 104 3157
rect 96 2981 97 2987
rect 103 2981 104 2987
rect 96 2831 104 2981
rect 96 2825 97 2831
rect 103 2825 104 2831
rect 96 2667 104 2825
rect 96 2661 97 2667
rect 103 2661 104 2667
rect 96 2507 104 2661
rect 96 2501 97 2507
rect 103 2501 104 2507
rect 96 2335 104 2501
rect 96 2329 97 2335
rect 103 2329 104 2335
rect 96 2171 104 2329
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 2003 104 2165
rect 96 1997 97 2003
rect 103 1997 104 2003
rect 96 1843 104 1997
rect 96 1837 97 1843
rect 103 1837 104 1843
rect 96 1679 104 1837
rect 96 1673 97 1679
rect 103 1673 104 1679
rect 96 1523 104 1673
rect 96 1517 97 1523
rect 103 1517 104 1523
rect 96 1363 104 1517
rect 96 1357 97 1363
rect 103 1357 104 1363
rect 96 1207 104 1357
rect 96 1201 97 1207
rect 103 1201 104 1207
rect 96 1043 104 1201
rect 96 1037 97 1043
rect 103 1037 104 1043
rect 96 875 104 1037
rect 96 869 97 875
rect 103 869 104 875
rect 96 699 104 869
rect 96 693 97 699
rect 103 693 104 699
rect 96 531 104 693
rect 96 525 97 531
rect 103 525 104 531
rect 96 359 104 525
rect 96 353 97 359
rect 103 353 104 359
rect 96 167 104 353
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 1842 3075 1850 3209
rect 1842 3069 1843 3075
rect 1849 3069 1850 3075
rect 1842 3051 1850 3069
rect 1842 3045 1843 3051
rect 1849 3045 1850 3051
rect 1842 2911 1850 3045
rect 1842 2905 1843 2911
rect 1849 2905 1850 2911
rect 1842 2887 1850 2905
rect 1842 2881 1843 2887
rect 1849 2881 1850 2887
rect 1842 2751 1850 2881
rect 1842 2745 1843 2751
rect 1849 2745 1850 2751
rect 1842 2723 1850 2745
rect 1842 2717 1843 2723
rect 1849 2717 1850 2723
rect 1842 2587 1850 2717
rect 1842 2581 1843 2587
rect 1849 2581 1850 2587
rect 1842 2563 1850 2581
rect 1842 2557 1843 2563
rect 1849 2557 1850 2563
rect 1842 2419 1850 2557
rect 1842 2413 1843 2419
rect 1849 2413 1850 2419
rect 1842 2399 1850 2413
rect 1842 2393 1843 2399
rect 1849 2393 1850 2399
rect 1842 2259 1850 2393
rect 1842 2253 1843 2259
rect 1849 2253 1850 2259
rect 1842 2243 1850 2253
rect 1842 2237 1843 2243
rect 1849 2237 1850 2243
rect 1842 2083 1850 2237
rect 1842 2077 1843 2083
rect 1849 2077 1850 2083
rect 1842 1923 1850 2077
rect 1842 1917 1843 1923
rect 1849 1917 1850 1923
rect 1842 1759 1850 1917
rect 1842 1753 1843 1759
rect 1849 1753 1850 1759
rect 1842 1747 1850 1753
rect 1842 1741 1843 1747
rect 1849 1741 1850 1747
rect 1842 1603 1850 1741
rect 1842 1597 1843 1603
rect 1849 1597 1850 1603
rect 1842 1583 1850 1597
rect 1842 1577 1843 1583
rect 1849 1577 1850 1583
rect 1842 1439 1850 1577
rect 1842 1433 1843 1439
rect 1849 1433 1850 1439
rect 1842 1423 1850 1433
rect 1842 1417 1843 1423
rect 1849 1417 1850 1423
rect 1842 1283 1850 1417
rect 1842 1277 1843 1283
rect 1849 1277 1850 1283
rect 1842 1255 1850 1277
rect 1842 1249 1843 1255
rect 1849 1249 1850 1255
rect 1842 1127 1850 1249
rect 1842 1121 1843 1127
rect 1849 1121 1850 1127
rect 1842 1091 1850 1121
rect 1842 1085 1843 1091
rect 1849 1085 1850 1091
rect 1842 959 1850 1085
rect 1842 953 1843 959
rect 1849 953 1850 959
rect 1842 931 1850 953
rect 1842 925 1843 931
rect 1849 925 1850 931
rect 1842 787 1850 925
rect 1842 781 1843 787
rect 1849 781 1850 787
rect 1842 759 1850 781
rect 1842 753 1843 759
rect 1849 753 1850 759
rect 1842 619 1850 753
rect 1842 613 1843 619
rect 1849 613 1850 619
rect 1842 599 1850 613
rect 1842 593 1843 599
rect 1849 593 1850 599
rect 1842 447 1850 593
rect 1842 441 1843 447
rect 1849 441 1850 447
rect 1842 275 1850 441
rect 1842 269 1843 275
rect 1849 269 1850 275
rect 1842 111 1850 269
rect 1842 105 1843 111
rect 1849 105 1850 111
rect 1842 91 1850 105
rect 1842 85 1843 91
rect 1849 85 1850 91
rect 1842 72 1850 85
rect 1854 3643 1862 3672
rect 1854 3637 1855 3643
rect 1861 3637 1862 3643
rect 1854 3595 1862 3637
rect 1854 3589 1855 3595
rect 1861 3589 1862 3595
rect 1854 3483 1862 3589
rect 1854 3477 1855 3483
rect 1861 3477 1862 3483
rect 1854 3443 1862 3477
rect 1854 3437 1855 3443
rect 1861 3437 1862 3443
rect 1854 3323 1862 3437
rect 1854 3317 1855 3323
rect 1861 3317 1862 3323
rect 1854 3291 1862 3317
rect 1854 3285 1855 3291
rect 1861 3285 1862 3291
rect 1854 3163 1862 3285
rect 1854 3157 1855 3163
rect 1861 3157 1862 3163
rect 1854 3139 1862 3157
rect 1854 3133 1855 3139
rect 1861 3133 1862 3139
rect 1854 2987 1862 3133
rect 1854 2981 1855 2987
rect 1861 2981 1862 2987
rect 1854 2963 1862 2981
rect 1854 2957 1855 2963
rect 1861 2957 1862 2963
rect 1854 2831 1862 2957
rect 1854 2825 1855 2831
rect 1861 2825 1862 2831
rect 1854 2799 1862 2825
rect 1854 2793 1855 2799
rect 1861 2793 1862 2799
rect 1854 2667 1862 2793
rect 1854 2661 1855 2667
rect 1861 2661 1862 2667
rect 1854 2639 1862 2661
rect 1854 2633 1855 2639
rect 1861 2633 1862 2639
rect 1854 2507 1862 2633
rect 1854 2501 1855 2507
rect 1861 2501 1862 2507
rect 1854 2479 1862 2501
rect 1854 2473 1855 2479
rect 1861 2473 1862 2479
rect 1854 2335 1862 2473
rect 1854 2329 1855 2335
rect 1861 2329 1862 2335
rect 1854 2319 1862 2329
rect 1854 2313 1855 2319
rect 1861 2313 1862 2319
rect 1854 2171 1862 2313
rect 1854 2165 1855 2171
rect 1861 2165 1862 2171
rect 1854 2163 1862 2165
rect 1854 2157 1855 2163
rect 1861 2157 1862 2163
rect 1854 2003 1862 2157
rect 1854 1997 1855 2003
rect 1861 1997 1862 2003
rect 1854 1843 1862 1997
rect 1854 1837 1855 1843
rect 1861 1837 1862 1843
rect 1854 1827 1862 1837
rect 1854 1821 1855 1827
rect 1861 1821 1862 1827
rect 1854 1679 1862 1821
rect 1854 1673 1855 1679
rect 1861 1673 1862 1679
rect 1854 1667 1862 1673
rect 1854 1661 1855 1667
rect 1861 1661 1862 1667
rect 1854 1523 1862 1661
rect 1854 1517 1855 1523
rect 1861 1517 1862 1523
rect 1854 1499 1862 1517
rect 1854 1493 1855 1499
rect 1861 1493 1862 1499
rect 1854 1363 1862 1493
rect 1854 1357 1855 1363
rect 1861 1357 1862 1363
rect 1854 1339 1862 1357
rect 1854 1333 1855 1339
rect 1861 1333 1862 1339
rect 1854 1207 1862 1333
rect 1854 1201 1855 1207
rect 1861 1201 1862 1207
rect 1854 1175 1862 1201
rect 1854 1169 1855 1175
rect 1861 1169 1862 1175
rect 1854 1043 1862 1169
rect 1854 1037 1855 1043
rect 1861 1037 1862 1043
rect 1854 1015 1862 1037
rect 1854 1009 1855 1015
rect 1861 1009 1862 1015
rect 1854 875 1862 1009
rect 1854 869 1855 875
rect 1861 869 1862 875
rect 1854 843 1862 869
rect 1854 837 1855 843
rect 1861 837 1862 843
rect 1854 699 1862 837
rect 1854 693 1855 699
rect 1861 693 1862 699
rect 1854 679 1862 693
rect 1854 673 1855 679
rect 1861 673 1862 679
rect 1854 531 1862 673
rect 1854 525 1855 531
rect 1861 525 1862 531
rect 1854 523 1862 525
rect 1854 517 1855 523
rect 1861 517 1862 523
rect 1854 359 1862 517
rect 1854 353 1855 359
rect 1861 353 1862 359
rect 1854 187 1862 353
rect 1854 181 1855 187
rect 1861 181 1862 187
rect 1854 167 1862 181
rect 1854 161 1855 167
rect 1861 161 1862 167
rect 1854 72 1862 161
rect 3618 3671 3626 3672
rect 3618 3665 3619 3671
rect 3625 3665 3626 3671
rect 3618 3519 3626 3665
rect 3618 3513 3619 3519
rect 3625 3513 3626 3519
rect 3618 3367 3626 3513
rect 3618 3361 3619 3367
rect 3625 3361 3626 3367
rect 3618 3215 3626 3361
rect 3618 3209 3619 3215
rect 3625 3209 3626 3215
rect 3618 3051 3626 3209
rect 3618 3045 3619 3051
rect 3625 3045 3626 3051
rect 3618 2887 3626 3045
rect 3618 2881 3619 2887
rect 3625 2881 3626 2887
rect 3618 2723 3626 2881
rect 3618 2717 3619 2723
rect 3625 2717 3626 2723
rect 3618 2563 3626 2717
rect 3618 2557 3619 2563
rect 3625 2557 3626 2563
rect 3618 2399 3626 2557
rect 3618 2393 3619 2399
rect 3625 2393 3626 2399
rect 3618 2243 3626 2393
rect 3618 2237 3619 2243
rect 3625 2237 3626 2243
rect 3618 1747 3626 2237
rect 3618 1741 3619 1747
rect 3625 1741 3626 1747
rect 3618 1583 3626 1741
rect 3618 1577 3619 1583
rect 3625 1577 3626 1583
rect 3618 1423 3626 1577
rect 3618 1417 3619 1423
rect 3625 1417 3626 1423
rect 3618 1255 3626 1417
rect 3618 1249 3619 1255
rect 3625 1249 3626 1255
rect 3618 1091 3626 1249
rect 3618 1085 3619 1091
rect 3625 1085 3626 1091
rect 3618 931 3626 1085
rect 3618 925 3619 931
rect 3625 925 3626 931
rect 3618 759 3626 925
rect 3618 753 3619 759
rect 3625 753 3626 759
rect 3618 599 3626 753
rect 3618 593 3619 599
rect 3625 593 3626 599
rect 3618 111 3626 593
rect 3618 105 3619 111
rect 3625 105 3626 111
rect 3618 72 3626 105
rect 3630 3595 3638 3672
rect 3630 3589 3631 3595
rect 3637 3589 3638 3595
rect 3630 3443 3638 3589
rect 3630 3437 3631 3443
rect 3637 3437 3638 3443
rect 3630 3291 3638 3437
rect 3630 3285 3631 3291
rect 3637 3285 3638 3291
rect 3630 3139 3638 3285
rect 3630 3133 3631 3139
rect 3637 3133 3638 3139
rect 3630 2963 3638 3133
rect 3630 2957 3631 2963
rect 3637 2957 3638 2963
rect 3630 2799 3638 2957
rect 3630 2793 3631 2799
rect 3637 2793 3638 2799
rect 3630 2639 3638 2793
rect 3630 2633 3631 2639
rect 3637 2633 3638 2639
rect 3630 2479 3638 2633
rect 3630 2473 3631 2479
rect 3637 2473 3638 2479
rect 3630 2319 3638 2473
rect 3630 2313 3631 2319
rect 3637 2313 3638 2319
rect 3630 2163 3638 2313
rect 3630 2157 3631 2163
rect 3637 2157 3638 2163
rect 3630 1827 3638 2157
rect 3630 1821 3631 1827
rect 3637 1821 3638 1827
rect 3630 1667 3638 1821
rect 3630 1661 3631 1667
rect 3637 1661 3638 1667
rect 3630 1499 3638 1661
rect 3630 1493 3631 1499
rect 3637 1493 3638 1499
rect 3630 1339 3638 1493
rect 3630 1333 3631 1339
rect 3637 1333 3638 1339
rect 3630 1175 3638 1333
rect 3630 1169 3631 1175
rect 3637 1169 3638 1175
rect 3630 1015 3638 1169
rect 3630 1009 3631 1015
rect 3637 1009 3638 1015
rect 3630 843 3638 1009
rect 3630 837 3631 843
rect 3637 837 3638 843
rect 3630 679 3638 837
rect 3630 673 3631 679
rect 3637 673 3638 679
rect 3630 523 3638 673
rect 3630 517 3631 523
rect 3637 517 3638 523
rect 3630 187 3638 517
rect 3630 181 3631 187
rect 3637 181 3638 187
rect 3630 72 3638 181
<< m6c >>
rect 906 3167 911 3171
rect 911 3167 917 3171
rect 917 3167 922 3171
rect 906 3155 922 3167
rect 1578 3155 1594 3171
<< m6 >>
rect 903 3171 1597 3174
rect 903 3155 906 3171
rect 922 3155 1578 3171
rect 1594 3155 1597 3171
rect 903 3152 1597 3155
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__173
timestamp 1731220585
transform 1 0 3584 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220585
transform 1 0 1864 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220585
transform 1 0 3584 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220585
transform 1 0 1864 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220585
transform 1 0 3584 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220585
transform 1 0 1864 0 -1 3496
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220585
transform 1 0 3584 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220585
transform 1 0 1864 0 1 3384
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220585
transform 1 0 3584 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220585
transform 1 0 1864 0 -1 3344
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220585
transform 1 0 3584 0 1 3232
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220585
transform 1 0 1864 0 1 3232
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220585
transform 1 0 3584 0 -1 3192
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220585
transform 1 0 1864 0 -1 3192
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220585
transform 1 0 3584 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220585
transform 1 0 1864 0 1 3080
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220585
transform 1 0 3584 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220585
transform 1 0 1864 0 -1 3028
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220585
transform 1 0 3584 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220585
transform 1 0 1864 0 1 2904
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220585
transform 1 0 3584 0 -1 2864
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220585
transform 1 0 1864 0 -1 2864
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220585
transform 1 0 3584 0 1 2740
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220585
transform 1 0 1864 0 1 2740
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220585
transform 1 0 3584 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220585
transform 1 0 1864 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220585
transform 1 0 3584 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220585
transform 1 0 1864 0 1 2580
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220585
transform 1 0 3584 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220585
transform 1 0 1864 0 -1 2540
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220585
transform 1 0 3584 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220585
transform 1 0 1864 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220585
transform 1 0 3584 0 -1 2376
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220585
transform 1 0 1864 0 -1 2376
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220585
transform 1 0 3584 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220585
transform 1 0 1864 0 1 2260
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220585
transform 1 0 3584 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220585
transform 1 0 1864 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220585
transform 1 0 3584 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220585
transform 1 0 1864 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220585
transform 1 0 3584 0 -1 2056
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220585
transform 1 0 1864 0 -1 2056
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220585
transform 1 0 3584 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220585
transform 1 0 1864 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220585
transform 1 0 3584 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220585
transform 1 0 1864 0 -1 1896
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220585
transform 1 0 3584 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220585
transform 1 0 1864 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220585
transform 1 0 3584 0 -1 1724
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220585
transform 1 0 1864 0 -1 1724
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220585
transform 1 0 3584 0 1 1608
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220585
transform 1 0 1864 0 1 1608
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220585
transform 1 0 3584 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220585
transform 1 0 1864 0 -1 1560
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220585
transform 1 0 3584 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220585
transform 1 0 1864 0 1 1440
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220585
transform 1 0 3584 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220585
transform 1 0 1864 0 -1 1400
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220585
transform 1 0 3584 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220585
transform 1 0 1864 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220585
transform 1 0 3584 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220585
transform 1 0 1864 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220585
transform 1 0 3584 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220585
transform 1 0 1864 0 1 1116
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220585
transform 1 0 3584 0 -1 1068
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220585
transform 1 0 1864 0 -1 1068
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220585
transform 1 0 3584 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220585
transform 1 0 1864 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220585
transform 1 0 3584 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220585
transform 1 0 1864 0 -1 908
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220585
transform 1 0 3584 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220585
transform 1 0 1864 0 1 784
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220585
transform 1 0 3584 0 -1 736
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220585
transform 1 0 1864 0 -1 736
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220585
transform 1 0 3584 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220585
transform 1 0 1864 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220585
transform 1 0 3584 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220585
transform 1 0 1864 0 -1 576
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220585
transform 1 0 3584 0 1 464
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220585
transform 1 0 1864 0 1 464
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220585
transform 1 0 3584 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220585
transform 1 0 1864 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220585
transform 1 0 3584 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220585
transform 1 0 1864 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220585
transform 1 0 3584 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220585
transform 1 0 1864 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220585
transform 1 0 3584 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220585
transform 1 0 1864 0 1 128
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220585
transform 1 0 1824 0 1 3584
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220585
transform 1 0 104 0 1 3584
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220585
transform 1 0 1824 0 -1 3544
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220585
transform 1 0 104 0 -1 3544
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220585
transform 1 0 1824 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220585
transform 1 0 104 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220585
transform 1 0 1824 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220585
transform 1 0 104 0 -1 3380
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220585
transform 1 0 1824 0 1 3264
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220585
transform 1 0 104 0 1 3264
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220585
transform 1 0 1824 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220585
transform 1 0 104 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220585
transform 1 0 1824 0 1 3104
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220585
transform 1 0 104 0 1 3104
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220585
transform 1 0 1824 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220585
transform 1 0 104 0 -1 3052
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220585
transform 1 0 1824 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220585
transform 1 0 104 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220585
transform 1 0 1824 0 -1 2888
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220585
transform 1 0 104 0 -1 2888
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220585
transform 1 0 1824 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220585
transform 1 0 104 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220585
transform 1 0 1824 0 -1 2728
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220585
transform 1 0 104 0 -1 2728
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220585
transform 1 0 1824 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220585
transform 1 0 104 0 1 2608
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220585
transform 1 0 1824 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220585
transform 1 0 104 0 -1 2564
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220585
transform 1 0 1824 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220585
transform 1 0 104 0 1 2448
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220585
transform 1 0 1824 0 -1 2396
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220585
transform 1 0 104 0 -1 2396
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220585
transform 1 0 1824 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220585
transform 1 0 104 0 1 2276
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220585
transform 1 0 1824 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220585
transform 1 0 104 0 -1 2236
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220585
transform 1 0 1824 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220585
transform 1 0 104 0 1 2112
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220585
transform 1 0 1824 0 -1 2060
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220585
transform 1 0 104 0 -1 2060
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220585
transform 1 0 1824 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220585
transform 1 0 104 0 1 1944
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220585
transform 1 0 1824 0 -1 1900
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220585
transform 1 0 104 0 -1 1900
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220585
transform 1 0 1824 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220585
transform 1 0 104 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220585
transform 1 0 1824 0 -1 1736
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220585
transform 1 0 104 0 -1 1736
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220585
transform 1 0 1824 0 1 1620
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220585
transform 1 0 104 0 1 1620
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220585
transform 1 0 1824 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220585
transform 1 0 104 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220585
transform 1 0 1824 0 1 1464
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220585
transform 1 0 104 0 1 1464
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220585
transform 1 0 1824 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220585
transform 1 0 104 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220585
transform 1 0 1824 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220585
transform 1 0 104 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220585
transform 1 0 1824 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220585
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220585
transform 1 0 1824 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220585
transform 1 0 104 0 1 1148
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220585
transform 1 0 1824 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220585
transform 1 0 104 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220585
transform 1 0 1824 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220585
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220585
transform 1 0 1824 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220585
transform 1 0 104 0 -1 936
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220585
transform 1 0 1824 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220585
transform 1 0 104 0 1 816
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220585
transform 1 0 1824 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220585
transform 1 0 104 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220585
transform 1 0 1824 0 1 640
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220585
transform 1 0 104 0 1 640
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220585
transform 1 0 1824 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220585
transform 1 0 104 0 -1 596
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220585
transform 1 0 1824 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220585
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220585
transform 1 0 1824 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220585
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220585
transform 1 0 1824 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220585
transform 1 0 104 0 1 300
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220585
transform 1 0 1824 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220585
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220585
transform 1 0 1824 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220585
transform 1 0 104 0 1 108
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCHINV  tst_5999_6
timestamp 1731220585
transform 1 0 3496 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5998_6
timestamp 1731220585
transform 1 0 3496 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5997_6
timestamp 1731220585
transform 1 0 3392 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5996_6
timestamp 1731220585
transform 1 0 3496 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5995_6
timestamp 1731220585
transform 1 0 3496 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5994_6
timestamp 1731220585
transform 1 0 3496 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5993_6
timestamp 1731220585
transform 1 0 3496 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5992_6
timestamp 1731220585
transform 1 0 3496 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5991_6
timestamp 1731220585
transform 1 0 3496 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5990_6
timestamp 1731220585
transform 1 0 3416 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5989_6
timestamp 1731220585
transform 1 0 3496 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5988_6
timestamp 1731220585
transform 1 0 3496 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5987_6
timestamp 1731220585
transform 1 0 3496 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5986_6
timestamp 1731220585
transform 1 0 3496 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5985_6
timestamp 1731220585
transform 1 0 3496 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5984_6
timestamp 1731220585
transform 1 0 3352 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5983_6
timestamp 1731220585
transform 1 0 3184 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5982_6
timestamp 1731220585
transform 1 0 3384 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5981_6
timestamp 1731220585
transform 1 0 3248 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5980_6
timestamp 1731220585
transform 1 0 3112 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5979_6
timestamp 1731220585
transform 1 0 2968 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5978_6
timestamp 1731220585
transform 1 0 3040 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5977_6
timestamp 1731220585
transform 1 0 3200 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5976_6
timestamp 1731220585
transform 1 0 3360 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5975_6
timestamp 1731220585
transform 1 0 3352 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5974_6
timestamp 1731220585
transform 1 0 3192 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5973_6
timestamp 1731220585
transform 1 0 3040 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5972_6
timestamp 1731220585
transform 1 0 3008 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5971_6
timestamp 1731220585
transform 1 0 3104 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5970_6
timestamp 1731220585
transform 1 0 3208 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5969_6
timestamp 1731220585
transform 1 0 3312 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5968_6
timestamp 1731220585
transform 1 0 3392 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5967_6
timestamp 1731220585
transform 1 0 3264 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5966_6
timestamp 1731220585
transform 1 0 3144 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5965_6
timestamp 1731220585
transform 1 0 3024 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5964_6
timestamp 1731220585
transform 1 0 3040 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5963_6
timestamp 1731220585
transform 1 0 3192 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5962_6
timestamp 1731220585
transform 1 0 3352 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5961_6
timestamp 1731220585
transform 1 0 3344 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5960_6
timestamp 1731220585
transform 1 0 3168 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5959_6
timestamp 1731220585
transform 1 0 2992 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5958_6
timestamp 1731220585
transform 1 0 2816 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5957_6
timestamp 1731220585
transform 1 0 2968 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5956_6
timestamp 1731220585
transform 1 0 3144 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5955_6
timestamp 1731220585
transform 1 0 3328 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5954_6
timestamp 1731220585
transform 1 0 3336 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5953_6
timestamp 1731220585
transform 1 0 3160 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5952_6
timestamp 1731220585
transform 1 0 3208 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5951_6
timestamp 1731220585
transform 1 0 3360 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5950_6
timestamp 1731220585
transform 1 0 3272 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5949_6
timestamp 1731220585
transform 1 0 3152 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5948_6
timestamp 1731220585
transform 1 0 3024 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5947_6
timestamp 1731220585
transform 1 0 3072 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5946_6
timestamp 1731220585
transform 1 0 3216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5945_6
timestamp 1731220585
transform 1 0 3368 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5944_6
timestamp 1731220585
transform 1 0 3384 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5943_6
timestamp 1731220585
transform 1 0 3288 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5942_6
timestamp 1731220585
transform 1 0 3192 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5941_6
timestamp 1731220585
transform 1 0 3096 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5940_6
timestamp 1731220585
transform 1 0 3000 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5939_6
timestamp 1731220585
transform 1 0 2904 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5938_6
timestamp 1731220585
transform 1 0 2800 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5937_6
timestamp 1731220585
transform 1 0 2688 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5936_6
timestamp 1731220585
transform 1 0 2568 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5935_6
timestamp 1731220585
transform 1 0 2640 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5934_6
timestamp 1731220585
transform 1 0 2784 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5933_6
timestamp 1731220585
transform 1 0 2928 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5932_6
timestamp 1731220585
transform 1 0 2896 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5931_6
timestamp 1731220585
transform 1 0 2760 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5930_6
timestamp 1731220585
transform 1 0 2792 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5929_6
timestamp 1731220585
transform 1 0 2920 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5928_6
timestamp 1731220585
transform 1 0 3064 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5927_6
timestamp 1731220585
transform 1 0 2984 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5926_6
timestamp 1731220585
transform 1 0 2824 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5925_6
timestamp 1731220585
transform 1 0 2800 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5924_6
timestamp 1731220585
transform 1 0 2640 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5923_6
timestamp 1731220585
transform 1 0 2640 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5922_6
timestamp 1731220585
transform 1 0 2464 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5921_6
timestamp 1731220585
transform 1 0 2584 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5920_6
timestamp 1731220585
transform 1 0 2736 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5919_6
timestamp 1731220585
transform 1 0 2888 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5918_6
timestamp 1731220585
transform 1 0 2768 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5917_6
timestamp 1731220585
transform 1 0 2896 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5916_6
timestamp 1731220585
transform 1 0 2904 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5915_6
timestamp 1731220585
transform 1 0 2800 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5914_6
timestamp 1731220585
transform 1 0 2896 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5913_6
timestamp 1731220585
transform 1 0 2768 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5912_6
timestamp 1731220585
transform 1 0 2744 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5911_6
timestamp 1731220585
transform 1 0 2888 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5910_6
timestamp 1731220585
transform 1 0 2824 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5909_6
timestamp 1731220585
transform 1 0 2672 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5908_6
timestamp 1731220585
transform 1 0 2656 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5907_6
timestamp 1731220585
transform 1 0 2464 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5906_6
timestamp 1731220585
transform 1 0 2840 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5905_6
timestamp 1731220585
transform 1 0 3016 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5904_6
timestamp 1731220585
transform 1 0 3168 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5903_6
timestamp 1731220585
transform 1 0 3048 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5902_6
timestamp 1731220585
transform 1 0 2936 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5901_6
timestamp 1731220585
transform 1 0 2824 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5900_6
timestamp 1731220585
transform 1 0 2704 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5899_6
timestamp 1731220585
transform 1 0 2576 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5898_6
timestamp 1731220585
transform 1 0 2904 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5897_6
timestamp 1731220585
transform 1 0 2784 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5896_6
timestamp 1731220585
transform 1 0 2664 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5895_6
timestamp 1731220585
transform 1 0 2544 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5894_6
timestamp 1731220585
transform 1 0 2424 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5893_6
timestamp 1731220585
transform 1 0 2552 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5892_6
timestamp 1731220585
transform 1 0 2704 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5891_6
timestamp 1731220585
transform 1 0 2864 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5890_6
timestamp 1731220585
transform 1 0 3024 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5889_6
timestamp 1731220585
transform 1 0 2976 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5888_6
timestamp 1731220585
transform 1 0 2832 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5887_6
timestamp 1731220585
transform 1 0 2680 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5886_6
timestamp 1731220585
transform 1 0 2768 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5885_6
timestamp 1731220585
transform 1 0 2912 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5884_6
timestamp 1731220585
transform 1 0 3056 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5883_6
timestamp 1731220585
transform 1 0 3040 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5882_6
timestamp 1731220585
transform 1 0 2920 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5881_6
timestamp 1731220585
transform 1 0 2792 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5880_6
timestamp 1731220585
transform 1 0 2864 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5879_6
timestamp 1731220585
transform 1 0 3016 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5878_6
timestamp 1731220585
transform 1 0 3152 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5877_6
timestamp 1731220585
transform 1 0 3264 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5876_6
timestamp 1731220585
transform 1 0 3360 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5875_6
timestamp 1731220585
transform 1 0 3208 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5874_6
timestamp 1731220585
transform 1 0 3112 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5873_6
timestamp 1731220585
transform 1 0 3248 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5872_6
timestamp 1731220585
transform 1 0 3384 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5871_6
timestamp 1731220585
transform 1 0 3352 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5870_6
timestamp 1731220585
transform 1 0 3184 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5869_6
timestamp 1731220585
transform 1 0 3496 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5868_6
timestamp 1731220585
transform 1 0 3496 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5867_6
timestamp 1731220585
transform 1 0 3496 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5866_6
timestamp 1731220585
transform 1 0 3496 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5865_6
timestamp 1731220585
transform 1 0 3384 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5864_6
timestamp 1731220585
transform 1 0 3456 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5863_6
timestamp 1731220585
transform 1 0 3304 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5862_6
timestamp 1731220585
transform 1 0 3160 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5861_6
timestamp 1731220585
transform 1 0 3240 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5860_6
timestamp 1731220585
transform 1 0 3112 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5859_6
timestamp 1731220585
transform 1 0 2984 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5858_6
timestamp 1731220585
transform 1 0 2864 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5857_6
timestamp 1731220585
transform 1 0 2752 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5856_6
timestamp 1731220585
transform 1 0 2656 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5855_6
timestamp 1731220585
transform 1 0 2568 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5854_6
timestamp 1731220585
transform 1 0 2480 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5853_6
timestamp 1731220585
transform 1 0 2392 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5852_6
timestamp 1731220585
transform 1 0 2312 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5851_6
timestamp 1731220585
transform 1 0 2432 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5850_6
timestamp 1731220585
transform 1 0 2568 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5849_6
timestamp 1731220585
transform 1 0 2728 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5848_6
timestamp 1731220585
transform 1 0 2904 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5847_6
timestamp 1731220585
transform 1 0 3312 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5846_6
timestamp 1731220585
transform 1 0 3104 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5845_6
timestamp 1731220585
transform 1 0 2992 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5844_6
timestamp 1731220585
transform 1 0 2832 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5843_6
timestamp 1731220585
transform 1 0 2648 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5842_6
timestamp 1731220585
transform 1 0 3136 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5841_6
timestamp 1731220585
transform 1 0 3264 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5840_6
timestamp 1731220585
transform 1 0 3336 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5839_6
timestamp 1731220585
transform 1 0 3160 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5838_6
timestamp 1731220585
transform 1 0 2992 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5837_6
timestamp 1731220585
transform 1 0 2832 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5836_6
timestamp 1731220585
transform 1 0 2680 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5835_6
timestamp 1731220585
transform 1 0 3168 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5834_6
timestamp 1731220585
transform 1 0 3000 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5833_6
timestamp 1731220585
transform 1 0 2848 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5832_6
timestamp 1731220585
transform 1 0 2712 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5831_6
timestamp 1731220585
transform 1 0 2592 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5830_6
timestamp 1731220585
transform 1 0 2584 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5829_6
timestamp 1731220585
transform 1 0 2664 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5828_6
timestamp 1731220585
transform 1 0 2920 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5827_6
timestamp 1731220585
transform 1 0 2832 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5826_6
timestamp 1731220585
transform 1 0 2744 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5825_6
timestamp 1731220585
transform 1 0 2696 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5824_6
timestamp 1731220585
transform 1 0 2840 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5823_6
timestamp 1731220585
transform 1 0 3168 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5822_6
timestamp 1731220585
transform 1 0 3000 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5821_6
timestamp 1731220585
transform 1 0 2848 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5820_6
timestamp 1731220585
transform 1 0 2688 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5819_6
timestamp 1731220585
transform 1 0 3176 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5818_6
timestamp 1731220585
transform 1 0 3008 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5817_6
timestamp 1731220585
transform 1 0 3112 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5816_6
timestamp 1731220585
transform 1 0 2752 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5815_6
timestamp 1731220585
transform 1 0 2616 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5814_6
timestamp 1731220585
transform 1 0 2880 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5813_6
timestamp 1731220585
transform 1 0 3000 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5812_6
timestamp 1731220585
transform 1 0 3000 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5811_6
timestamp 1731220585
transform 1 0 3272 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5810_6
timestamp 1731220585
transform 1 0 3216 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5809_6
timestamp 1731220585
transform 1 0 3312 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5808_6
timestamp 1731220585
transform 1 0 3416 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5807_6
timestamp 1731220585
transform 1 0 3344 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5806_6
timestamp 1731220585
transform 1 0 3344 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5805_6
timestamp 1731220585
transform 1 0 3344 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5804_6
timestamp 1731220585
transform 1 0 3392 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5803_6
timestamp 1731220585
transform 1 0 3376 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5802_6
timestamp 1731220585
transform 1 0 3496 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5801_6
timestamp 1731220585
transform 1 0 3496 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5800_6
timestamp 1731220585
transform 1 0 3496 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5799_6
timestamp 1731220585
transform 1 0 3496 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5798_6
timestamp 1731220585
transform 1 0 3496 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5797_6
timestamp 1731220585
transform 1 0 3496 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5796_6
timestamp 1731220585
transform 1 0 3496 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5795_6
timestamp 1731220585
transform 1 0 3496 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5794_6
timestamp 1731220585
transform 1 0 3496 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5793_6
timestamp 1731220585
transform 1 0 3496 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5792_6
timestamp 1731220585
transform 1 0 3496 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5791_6
timestamp 1731220585
transform 1 0 3480 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5790_6
timestamp 1731220585
transform 1 0 3352 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5789_6
timestamp 1731220585
transform 1 0 3368 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5788_6
timestamp 1731220585
transform 1 0 3368 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5787_6
timestamp 1731220585
transform 1 0 3216 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5786_6
timestamp 1731220585
transform 1 0 3064 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5785_6
timestamp 1731220585
transform 1 0 2904 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5784_6
timestamp 1731220585
transform 1 0 2728 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5783_6
timestamp 1731220585
transform 1 0 3216 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5782_6
timestamp 1731220585
transform 1 0 3072 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5781_6
timestamp 1731220585
transform 1 0 2928 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5780_6
timestamp 1731220585
transform 1 0 2776 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5779_6
timestamp 1731220585
transform 1 0 2624 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5778_6
timestamp 1731220585
transform 1 0 3024 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5777_6
timestamp 1731220585
transform 1 0 3184 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5776_6
timestamp 1731220585
transform 1 0 3320 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5775_6
timestamp 1731220585
transform 1 0 3168 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5774_6
timestamp 1731220585
transform 1 0 3032 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5773_6
timestamp 1731220585
transform 1 0 3176 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5772_6
timestamp 1731220585
transform 1 0 3320 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5771_6
timestamp 1731220585
transform 1 0 3184 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5770_6
timestamp 1731220585
transform 1 0 3000 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5769_6
timestamp 1731220585
transform 1 0 3376 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5768_6
timestamp 1731220585
transform 1 0 3320 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5767_6
timestamp 1731220585
transform 1 0 3144 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5766_6
timestamp 1731220585
transform 1 0 3496 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5765_6
timestamp 1731220585
transform 1 0 3496 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5764_6
timestamp 1731220585
transform 1 0 3496 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5763_6
timestamp 1731220585
transform 1 0 3496 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5762_6
timestamp 1731220585
transform 1 0 3496 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5761_6
timestamp 1731220585
transform 1 0 3408 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5760_6
timestamp 1731220585
transform 1 0 3296 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5759_6
timestamp 1731220585
transform 1 0 3184 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5758_6
timestamp 1731220585
transform 1 0 3072 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5757_6
timestamp 1731220585
transform 1 0 2952 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5756_6
timestamp 1731220585
transform 1 0 2960 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5755_6
timestamp 1731220585
transform 1 0 3248 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5754_6
timestamp 1731220585
transform 1 0 3104 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5753_6
timestamp 1731220585
transform 1 0 3008 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5752_6
timestamp 1731220585
transform 1 0 2720 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5751_6
timestamp 1731220585
transform 1 0 2432 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5750_6
timestamp 1731220585
transform 1 0 2816 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5749_6
timestamp 1731220585
transform 1 0 2680 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5748_6
timestamp 1731220585
transform 1 0 2664 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5747_6
timestamp 1731220585
transform 1 0 2816 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5746_6
timestamp 1731220585
transform 1 0 2816 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5745_6
timestamp 1731220585
transform 1 0 2984 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5744_6
timestamp 1731220585
transform 1 0 3152 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5743_6
timestamp 1731220585
transform 1 0 3328 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5742_6
timestamp 1731220585
transform 1 0 3344 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5741_6
timestamp 1731220585
transform 1 0 3176 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5740_6
timestamp 1731220585
transform 1 0 3016 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5739_6
timestamp 1731220585
transform 1 0 2864 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5738_6
timestamp 1731220585
transform 1 0 2720 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5737_6
timestamp 1731220585
transform 1 0 3296 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5736_6
timestamp 1731220585
transform 1 0 3096 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5735_6
timestamp 1731220585
transform 1 0 2904 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5734_6
timestamp 1731220585
transform 1 0 2728 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5733_6
timestamp 1731220585
transform 1 0 2576 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5732_6
timestamp 1731220585
transform 1 0 2616 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5731_6
timestamp 1731220585
transform 1 0 2792 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5730_6
timestamp 1731220585
transform 1 0 2968 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5729_6
timestamp 1731220585
transform 1 0 2816 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5728_6
timestamp 1731220585
transform 1 0 2632 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5727_6
timestamp 1731220585
transform 1 0 2616 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5726_6
timestamp 1731220585
transform 1 0 2760 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5725_6
timestamp 1731220585
transform 1 0 2896 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5724_6
timestamp 1731220585
transform 1 0 3024 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5723_6
timestamp 1731220585
transform 1 0 2896 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5722_6
timestamp 1731220585
transform 1 0 2872 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5721_6
timestamp 1731220585
transform 1 0 2720 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5720_6
timestamp 1731220585
transform 1 0 2584 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5719_6
timestamp 1731220585
transform 1 0 2776 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5718_6
timestamp 1731220585
transform 1 0 2680 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5717_6
timestamp 1731220585
transform 1 0 2592 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5716_6
timestamp 1731220585
transform 1 0 2512 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5715_6
timestamp 1731220585
transform 1 0 2432 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5714_6
timestamp 1731220585
transform 1 0 2352 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5713_6
timestamp 1731220585
transform 1 0 2272 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5712_6
timestamp 1731220585
transform 1 0 2232 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5711_6
timestamp 1731220585
transform 1 0 2336 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5710_6
timestamp 1731220585
transform 1 0 2456 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5709_6
timestamp 1731220585
transform 1 0 2472 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5708_6
timestamp 1731220585
transform 1 0 2000 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5707_6
timestamp 1731220585
transform 1 0 1888 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5706_6
timestamp 1731220585
transform 1 0 2096 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5705_6
timestamp 1731220585
transform 1 0 1888 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5704_6
timestamp 1731220585
transform 1 0 1736 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5703_6
timestamp 1731220585
transform 1 0 1600 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5702_6
timestamp 1731220585
transform 1 0 1736 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5701_6
timestamp 1731220585
transform 1 0 1632 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5700_6
timestamp 1731220585
transform 1 0 1512 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5699_6
timestamp 1731220585
transform 1 0 1392 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5698_6
timestamp 1731220585
transform 1 0 1688 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5697_6
timestamp 1731220585
transform 1 0 1584 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5696_6
timestamp 1731220585
transform 1 0 1480 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5695_6
timestamp 1731220585
transform 1 0 1384 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5694_6
timestamp 1731220585
transform 1 0 1632 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5693_6
timestamp 1731220585
transform 1 0 1520 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5692_6
timestamp 1731220585
transform 1 0 1408 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5691_6
timestamp 1731220585
transform 1 0 1296 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5690_6
timestamp 1731220585
transform 1 0 1184 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5689_6
timestamp 1731220585
transform 1 0 1064 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5688_6
timestamp 1731220585
transform 1 0 928 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5687_6
timestamp 1731220585
transform 1 0 1280 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5686_6
timestamp 1731220585
transform 1 0 1168 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5685_6
timestamp 1731220585
transform 1 0 1048 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5684_6
timestamp 1731220585
transform 1 0 920 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5683_6
timestamp 1731220585
transform 1 0 984 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5682_6
timestamp 1731220585
transform 1 0 1264 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5681_6
timestamp 1731220585
transform 1 0 1128 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5680_6
timestamp 1731220585
transform 1 0 1128 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5679_6
timestamp 1731220585
transform 1 0 968 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5678_6
timestamp 1731220585
transform 1 0 1280 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5677_6
timestamp 1731220585
transform 1 0 1440 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5676_6
timestamp 1731220585
transform 1 0 1536 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5675_6
timestamp 1731220585
transform 1 0 1384 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5674_6
timestamp 1731220585
transform 1 0 1232 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5673_6
timestamp 1731220585
transform 1 0 1088 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5672_6
timestamp 1731220585
transform 1 0 936 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5671_6
timestamp 1731220585
transform 1 0 1040 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5670_6
timestamp 1731220585
transform 1 0 1200 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5669_6
timestamp 1731220585
transform 1 0 1352 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5668_6
timestamp 1731220585
transform 1 0 1504 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5667_6
timestamp 1731220585
transform 1 0 1664 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5666_6
timestamp 1731220585
transform 1 0 1656 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5665_6
timestamp 1731220585
transform 1 0 1536 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5664_6
timestamp 1731220585
transform 1 0 1416 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5663_6
timestamp 1731220585
transform 1 0 1296 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5662_6
timestamp 1731220585
transform 1 0 1176 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5661_6
timestamp 1731220585
transform 1 0 1048 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5660_6
timestamp 1731220585
transform 1 0 1456 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5659_6
timestamp 1731220585
transform 1 0 1376 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5658_6
timestamp 1731220585
transform 1 0 1296 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5657_6
timestamp 1731220585
transform 1 0 1216 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5656_6
timestamp 1731220585
transform 1 0 1136 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5655_6
timestamp 1731220585
transform 1 0 1056 0 -1 2416
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5654_6
timestamp 1731220585
transform 1 0 1304 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5653_6
timestamp 1731220585
transform 1 0 1224 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5652_6
timestamp 1731220585
transform 1 0 1144 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5651_6
timestamp 1731220585
transform 1 0 1064 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5650_6
timestamp 1731220585
transform 1 0 984 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5649_6
timestamp 1731220585
transform 1 0 1248 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5648_6
timestamp 1731220585
transform 1 0 1168 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5647_6
timestamp 1731220585
transform 1 0 1088 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5646_6
timestamp 1731220585
transform 1 0 1008 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5645_6
timestamp 1731220585
transform 1 0 928 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5644_6
timestamp 1731220585
transform 1 0 848 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5643_6
timestamp 1731220585
transform 1 0 848 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5642_6
timestamp 1731220585
transform 1 0 936 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5641_6
timestamp 1731220585
transform 1 0 1024 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5640_6
timestamp 1731220585
transform 1 0 1112 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5639_6
timestamp 1731220585
transform 1 0 1208 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5638_6
timestamp 1731220585
transform 1 0 1168 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5637_6
timestamp 1731220585
transform 1 0 1056 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5636_6
timestamp 1731220585
transform 1 0 936 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5635_6
timestamp 1731220585
transform 1 0 1000 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5634_6
timestamp 1731220585
transform 1 0 1152 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5633_6
timestamp 1731220585
transform 1 0 1152 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5632_6
timestamp 1731220585
transform 1 0 1000 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5631_6
timestamp 1731220585
transform 1 0 1008 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5630_6
timestamp 1731220585
transform 1 0 1160 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5629_6
timestamp 1731220585
transform 1 0 1000 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5628_6
timestamp 1731220585
transform 1 0 1016 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5627_6
timestamp 1731220585
transform 1 0 1112 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5626_6
timestamp 1731220585
transform 1 0 976 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5625_6
timestamp 1731220585
transform 1 0 1000 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5624_6
timestamp 1731220585
transform 1 0 888 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5623_6
timestamp 1731220585
transform 1 0 912 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5622_6
timestamp 1731220585
transform 1 0 848 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5621_6
timestamp 1731220585
transform 1 0 992 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5620_6
timestamp 1731220585
transform 1 0 1128 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5619_6
timestamp 1731220585
transform 1 0 1096 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5618_6
timestamp 1731220585
transform 1 0 952 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5617_6
timestamp 1731220585
transform 1 0 808 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5616_6
timestamp 1731220585
transform 1 0 744 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5615_6
timestamp 1731220585
transform 1 0 912 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5614_6
timestamp 1731220585
transform 1 0 840 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5613_6
timestamp 1731220585
transform 1 0 704 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5612_6
timestamp 1731220585
transform 1 0 560 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5611_6
timestamp 1731220585
transform 1 0 536 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5610_6
timestamp 1731220585
transform 1 0 672 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5609_6
timestamp 1731220585
transform 1 0 680 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5608_6
timestamp 1731220585
transform 1 0 560 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5607_6
timestamp 1731220585
transform 1 0 544 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5606_6
timestamp 1731220585
transform 1 0 704 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5605_6
timestamp 1731220585
transform 1 0 856 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5604_6
timestamp 1731220585
transform 1 0 776 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5603_6
timestamp 1731220585
transform 1 0 944 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5602_6
timestamp 1731220585
transform 1 0 888 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5601_6
timestamp 1731220585
transform 1 0 768 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5600_6
timestamp 1731220585
transform 1 0 640 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5599_6
timestamp 1731220585
transform 1 0 728 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5598_6
timestamp 1731220585
transform 1 0 640 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5597_6
timestamp 1731220585
transform 1 0 520 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5596_6
timestamp 1731220585
transform 1 0 424 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5595_6
timestamp 1731220585
transform 1 0 488 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5594_6
timestamp 1731220585
transform 1 0 600 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5593_6
timestamp 1731220585
transform 1 0 712 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5592_6
timestamp 1731220585
transform 1 0 760 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5591_6
timestamp 1731220585
transform 1 0 632 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5590_6
timestamp 1731220585
transform 1 0 592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5589_6
timestamp 1731220585
transform 1 0 728 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5588_6
timestamp 1731220585
transform 1 0 864 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5587_6
timestamp 1731220585
transform 1 0 808 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5586_6
timestamp 1731220585
transform 1 0 720 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5585_6
timestamp 1731220585
transform 1 0 632 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5584_6
timestamp 1731220585
transform 1 0 544 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5583_6
timestamp 1731220585
transform 1 0 464 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5582_6
timestamp 1731220585
transform 1 0 384 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5581_6
timestamp 1731220585
transform 1 0 304 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5580_6
timestamp 1731220585
transform 1 0 224 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5579_6
timestamp 1731220585
transform 1 0 144 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5578_6
timestamp 1731220585
transform 1 0 216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5577_6
timestamp 1731220585
transform 1 0 328 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5576_6
timestamp 1731220585
transform 1 0 456 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5575_6
timestamp 1731220585
transform 1 0 496 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5574_6
timestamp 1731220585
transform 1 0 360 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5573_6
timestamp 1731220585
transform 1 0 232 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5572_6
timestamp 1731220585
transform 1 0 128 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5571_6
timestamp 1731220585
transform 1 0 128 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5570_6
timestamp 1731220585
transform 1 0 240 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5569_6
timestamp 1731220585
transform 1 0 368 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5568_6
timestamp 1731220585
transform 1 0 328 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5567_6
timestamp 1731220585
transform 1 0 224 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5566_6
timestamp 1731220585
transform 1 0 304 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5565_6
timestamp 1731220585
transform 1 0 384 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5564_6
timestamp 1731220585
transform 1 0 464 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5563_6
timestamp 1731220585
transform 1 0 552 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5562_6
timestamp 1731220585
transform 1 0 512 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5561_6
timestamp 1731220585
transform 1 0 392 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5560_6
timestamp 1731220585
transform 1 0 280 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5559_6
timestamp 1731220585
transform 1 0 600 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5558_6
timestamp 1731220585
transform 1 0 424 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5557_6
timestamp 1731220585
transform 1 0 256 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5556_6
timestamp 1731220585
transform 1 0 128 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5555_6
timestamp 1731220585
transform 1 0 128 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5554_6
timestamp 1731220585
transform 1 0 240 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5553_6
timestamp 1731220585
transform 1 0 384 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5552_6
timestamp 1731220585
transform 1 0 440 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5551_6
timestamp 1731220585
transform 1 0 320 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5550_6
timestamp 1731220585
transform 1 0 208 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5549_6
timestamp 1731220585
transform 1 0 128 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5548_6
timestamp 1731220585
transform 1 0 128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5547_6
timestamp 1731220585
transform 1 0 392 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5546_6
timestamp 1731220585
transform 1 0 248 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5545_6
timestamp 1731220585
transform 1 0 136 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5544_6
timestamp 1731220585
transform 1 0 272 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5543_6
timestamp 1731220585
transform 1 0 416 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5542_6
timestamp 1731220585
transform 1 0 576 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5541_6
timestamp 1731220585
transform 1 0 400 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5540_6
timestamp 1731220585
transform 1 0 224 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5539_6
timestamp 1731220585
transform 1 0 304 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5538_6
timestamp 1731220585
transform 1 0 408 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5537_6
timestamp 1731220585
transform 1 0 528 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5536_6
timestamp 1731220585
transform 1 0 664 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5535_6
timestamp 1731220585
transform 1 0 712 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5534_6
timestamp 1731220585
transform 1 0 576 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5533_6
timestamp 1731220585
transform 1 0 456 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5532_6
timestamp 1731220585
transform 1 0 344 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5531_6
timestamp 1731220585
transform 1 0 248 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5530_6
timestamp 1731220585
transform 1 0 344 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5529_6
timestamp 1731220585
transform 1 0 440 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5528_6
timestamp 1731220585
transform 1 0 360 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5527_6
timestamp 1731220585
transform 1 0 216 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5526_6
timestamp 1731220585
transform 1 0 280 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5525_6
timestamp 1731220585
transform 1 0 152 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5524_6
timestamp 1731220585
transform 1 0 128 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5523_6
timestamp 1731220585
transform 1 0 280 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5522_6
timestamp 1731220585
transform 1 0 336 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5521_6
timestamp 1731220585
transform 1 0 208 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5520_6
timestamp 1731220585
transform 1 0 128 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5519_6
timestamp 1731220585
transform 1 0 128 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5518_6
timestamp 1731220585
transform 1 0 272 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5517_6
timestamp 1731220585
transform 1 0 368 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5516_6
timestamp 1731220585
transform 1 0 232 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5515_6
timestamp 1731220585
transform 1 0 128 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5514_6
timestamp 1731220585
transform 1 0 176 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5513_6
timestamp 1731220585
transform 1 0 336 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5512_6
timestamp 1731220585
transform 1 0 440 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5511_6
timestamp 1731220585
transform 1 0 320 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5510_6
timestamp 1731220585
transform 1 0 200 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5509_6
timestamp 1731220585
transform 1 0 296 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5508_6
timestamp 1731220585
transform 1 0 392 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5507_6
timestamp 1731220585
transform 1 0 488 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5506_6
timestamp 1731220585
transform 1 0 528 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5505_6
timestamp 1731220585
transform 1 0 448 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5504_6
timestamp 1731220585
transform 1 0 368 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5503_6
timestamp 1731220585
transform 1 0 344 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5502_6
timestamp 1731220585
transform 1 0 424 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5501_6
timestamp 1731220585
transform 1 0 504 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5500_6
timestamp 1731220585
transform 1 0 584 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5499_6
timestamp 1731220585
transform 1 0 664 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5498_6
timestamp 1731220585
transform 1 0 744 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5497_6
timestamp 1731220585
transform 1 0 904 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5496_6
timestamp 1731220585
transform 1 0 824 0 1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5495_6
timestamp 1731220585
transform 1 0 768 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5494_6
timestamp 1731220585
transform 1 0 688 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5493_6
timestamp 1731220585
transform 1 0 608 0 -1 2256
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5492_6
timestamp 1731220585
transform 1 0 760 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5491_6
timestamp 1731220585
transform 1 0 672 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5490_6
timestamp 1731220585
transform 1 0 584 0 1 2092
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5489_6
timestamp 1731220585
transform 1 0 568 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5488_6
timestamp 1731220585
transform 1 0 696 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5487_6
timestamp 1731220585
transform 1 0 816 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5486_6
timestamp 1731220585
transform 1 0 840 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5485_6
timestamp 1731220585
transform 1 0 672 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5484_6
timestamp 1731220585
transform 1 0 504 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5483_6
timestamp 1731220585
transform 1 0 520 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5482_6
timestamp 1731220585
transform 1 0 680 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5481_6
timestamp 1731220585
transform 1 0 840 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5480_6
timestamp 1731220585
transform 1 0 832 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5479_6
timestamp 1731220585
transform 1 0 648 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5478_6
timestamp 1731220585
transform 1 0 456 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5477_6
timestamp 1731220585
transform 1 0 488 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5476_6
timestamp 1731220585
transform 1 0 656 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5475_6
timestamp 1731220585
transform 1 0 832 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5474_6
timestamp 1731220585
transform 1 0 656 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5473_6
timestamp 1731220585
transform 1 0 464 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5472_6
timestamp 1731220585
transform 1 0 840 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5471_6
timestamp 1731220585
transform 1 0 840 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5470_6
timestamp 1731220585
transform 1 0 704 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5469_6
timestamp 1731220585
transform 1 0 560 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5468_6
timestamp 1731220585
transform 1 0 416 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5467_6
timestamp 1731220585
transform 1 0 504 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5466_6
timestamp 1731220585
transform 1 0 768 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5465_6
timestamp 1731220585
transform 1 0 640 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5464_6
timestamp 1731220585
transform 1 0 624 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5463_6
timestamp 1731220585
transform 1 0 536 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5462_6
timestamp 1731220585
transform 1 0 712 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5461_6
timestamp 1731220585
transform 1 0 800 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5460_6
timestamp 1731220585
transform 1 0 1040 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5459_6
timestamp 1731220585
transform 1 0 1200 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5458_6
timestamp 1731220585
transform 1 0 1568 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5457_6
timestamp 1731220585
transform 1 0 1376 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5456_6
timestamp 1731220585
transform 1 0 1304 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5455_6
timestamp 1731220585
transform 1 0 1200 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5454_6
timestamp 1731220585
transform 1 0 1104 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5453_6
timestamp 1731220585
transform 1 0 1408 0 1 1444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5452_6
timestamp 1731220585
transform 1 0 1504 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5451_6
timestamp 1731220585
transform 1 0 1368 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5450_6
timestamp 1731220585
transform 1 0 1240 0 -1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5449_6
timestamp 1731220585
transform 1 0 1184 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5448_6
timestamp 1731220585
transform 1 0 1344 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5447_6
timestamp 1731220585
transform 1 0 1504 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5446_6
timestamp 1731220585
transform 1 0 1664 0 1 1600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5445_6
timestamp 1731220585
transform 1 0 1736 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5444_6
timestamp 1731220585
transform 1 0 1600 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5443_6
timestamp 1731220585
transform 1 0 1456 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5442_6
timestamp 1731220585
transform 1 0 1312 0 -1 1756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5441_6
timestamp 1731220585
transform 1 0 1664 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5440_6
timestamp 1731220585
transform 1 0 1496 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5439_6
timestamp 1731220585
transform 1 0 1336 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5438_6
timestamp 1731220585
transform 1 0 1176 0 1 1764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5437_6
timestamp 1731220585
transform 1 0 1296 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5436_6
timestamp 1731220585
transform 1 0 1448 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5435_6
timestamp 1731220585
transform 1 0 1600 0 -1 1920
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5434_6
timestamp 1731220585
transform 1 0 1704 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5433_6
timestamp 1731220585
transform 1 0 1568 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5432_6
timestamp 1731220585
transform 1 0 1432 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5431_6
timestamp 1731220585
transform 1 0 1296 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5430_6
timestamp 1731220585
transform 1 0 1272 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5429_6
timestamp 1731220585
transform 1 0 1368 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5428_6
timestamp 1731220585
transform 1 0 1464 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5427_6
timestamp 1731220585
transform 1 0 1560 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5426_6
timestamp 1731220585
transform 1 0 1656 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5425_6
timestamp 1731220585
transform 1 0 1736 0 -1 2080
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5424_6
timestamp 1731220585
transform 1 0 1888 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5423_6
timestamp 1731220585
transform 1 0 1968 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5422_6
timestamp 1731220585
transform 1 0 2376 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5421_6
timestamp 1731220585
transform 1 0 2232 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5420_6
timestamp 1731220585
transform 1 0 2096 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5419_6
timestamp 1731220585
transform 1 0 1960 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5418_6
timestamp 1731220585
transform 1 0 1944 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5417_6
timestamp 1731220585
transform 1 0 2064 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5416_6
timestamp 1731220585
transform 1 0 2184 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5415_6
timestamp 1731220585
transform 1 0 2144 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5414_6
timestamp 1731220585
transform 1 0 2056 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5413_6
timestamp 1731220585
transform 1 0 2080 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5412_6
timestamp 1731220585
transform 1 0 2224 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5411_6
timestamp 1731220585
transform 1 0 2384 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5410_6
timestamp 1731220585
transform 1 0 2376 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5409_6
timestamp 1731220585
transform 1 0 2232 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5408_6
timestamp 1731220585
transform 1 0 2096 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5407_6
timestamp 1731220585
transform 1 0 2336 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5406_6
timestamp 1731220585
transform 1 0 2200 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5405_6
timestamp 1731220585
transform 1 0 2072 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5404_6
timestamp 1731220585
transform 1 0 1952 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5403_6
timestamp 1731220585
transform 1 0 1888 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5402_6
timestamp 1731220585
transform 1 0 2040 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5401_6
timestamp 1731220585
transform 1 0 2200 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5400_6
timestamp 1731220585
transform 1 0 2120 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5399_6
timestamp 1731220585
transform 1 0 1992 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5398_6
timestamp 1731220585
transform 1 0 1888 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5397_6
timestamp 1731220585
transform 1 0 1888 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5396_6
timestamp 1731220585
transform 1 0 1736 0 -1 1436
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5395_6
timestamp 1731220585
transform 1 0 1736 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5394_6
timestamp 1731220585
transform 1 0 1632 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5393_6
timestamp 1731220585
transform 1 0 1512 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5392_6
timestamp 1731220585
transform 1 0 1392 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5391_6
timestamp 1731220585
transform 1 0 1264 0 1 1284
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5390_6
timestamp 1731220585
transform 1 0 1624 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5389_6
timestamp 1731220585
transform 1 0 1496 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5388_6
timestamp 1731220585
transform 1 0 1368 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5387_6
timestamp 1731220585
transform 1 0 1232 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5386_6
timestamp 1731220585
transform 1 0 1624 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5385_6
timestamp 1731220585
transform 1 0 1488 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5384_6
timestamp 1731220585
transform 1 0 1352 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5383_6
timestamp 1731220585
transform 1 0 1208 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5382_6
timestamp 1731220585
transform 1 0 1064 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5381_6
timestamp 1731220585
transform 1 0 1464 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5380_6
timestamp 1731220585
transform 1 0 1336 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5379_6
timestamp 1731220585
transform 1 0 1216 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5378_6
timestamp 1731220585
transform 1 0 1096 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5377_6
timestamp 1731220585
transform 1 0 968 0 -1 1124
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5376_6
timestamp 1731220585
transform 1 0 1344 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5375_6
timestamp 1731220585
transform 1 0 1232 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5374_6
timestamp 1731220585
transform 1 0 1128 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5373_6
timestamp 1731220585
transform 1 0 1024 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5372_6
timestamp 1731220585
transform 1 0 912 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5371_6
timestamp 1731220585
transform 1 0 792 0 1 964
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5370_6
timestamp 1731220585
transform 1 0 792 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5369_6
timestamp 1731220585
transform 1 0 904 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5368_6
timestamp 1731220585
transform 1 0 1008 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5367_6
timestamp 1731220585
transform 1 0 1112 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5366_6
timestamp 1731220585
transform 1 0 1320 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5365_6
timestamp 1731220585
transform 1 0 1216 0 -1 956
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5364_6
timestamp 1731220585
transform 1 0 1136 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5363_6
timestamp 1731220585
transform 1 0 1000 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5362_6
timestamp 1731220585
transform 1 0 1264 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5361_6
timestamp 1731220585
transform 1 0 1384 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5360_6
timestamp 1731220585
transform 1 0 1504 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5359_6
timestamp 1731220585
transform 1 0 1632 0 1 796
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5358_6
timestamp 1731220585
transform 1 0 1736 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5357_6
timestamp 1731220585
transform 1 0 1632 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5356_6
timestamp 1731220585
transform 1 0 1504 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5355_6
timestamp 1731220585
transform 1 0 1376 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5354_6
timestamp 1731220585
transform 1 0 1240 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5353_6
timestamp 1731220585
transform 1 0 1096 0 -1 784
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5352_6
timestamp 1731220585
transform 1 0 1544 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5351_6
timestamp 1731220585
transform 1 0 1440 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5350_6
timestamp 1731220585
transform 1 0 1336 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5349_6
timestamp 1731220585
transform 1 0 1232 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5348_6
timestamp 1731220585
transform 1 0 1120 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5347_6
timestamp 1731220585
transform 1 0 1008 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5346_6
timestamp 1731220585
transform 1 0 1256 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5345_6
timestamp 1731220585
transform 1 0 1168 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5344_6
timestamp 1731220585
transform 1 0 1080 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5343_6
timestamp 1731220585
transform 1 0 992 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5342_6
timestamp 1731220585
transform 1 0 904 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5341_6
timestamp 1731220585
transform 1 0 816 0 -1 616
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5340_6
timestamp 1731220585
transform 1 0 1232 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5339_6
timestamp 1731220585
transform 1 0 1144 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5338_6
timestamp 1731220585
transform 1 0 1056 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5337_6
timestamp 1731220585
transform 1 0 968 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5336_6
timestamp 1731220585
transform 1 0 880 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5335_6
timestamp 1731220585
transform 1 0 792 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5334_6
timestamp 1731220585
transform 1 0 704 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5333_6
timestamp 1731220585
transform 1 0 616 0 1 452
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5332_6
timestamp 1731220585
transform 1 0 816 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5331_6
timestamp 1731220585
transform 1 0 912 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5330_6
timestamp 1731220585
transform 1 0 1000 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5329_6
timestamp 1731220585
transform 1 0 1096 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5328_6
timestamp 1731220585
transform 1 0 1288 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5327_6
timestamp 1731220585
transform 1 0 1192 0 -1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5326_6
timestamp 1731220585
transform 1 0 1104 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5325_6
timestamp 1731220585
transform 1 0 992 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5324_6
timestamp 1731220585
transform 1 0 880 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5323_6
timestamp 1731220585
transform 1 0 1208 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5322_6
timestamp 1731220585
transform 1 0 1424 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5321_6
timestamp 1731220585
transform 1 0 1312 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5320_6
timestamp 1731220585
transform 1 0 1248 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5319_6
timestamp 1731220585
transform 1 0 1128 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5318_6
timestamp 1731220585
transform 1 0 1000 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5317_6
timestamp 1731220585
transform 1 0 1592 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5316_6
timestamp 1731220585
transform 1 0 1472 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5315_6
timestamp 1731220585
transform 1 0 1360 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5314_6
timestamp 1731220585
transform 1 0 1072 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5313_6
timestamp 1731220585
transform 1 0 984 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5312_6
timestamp 1731220585
transform 1 0 896 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5311_6
timestamp 1731220585
transform 1 0 1152 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5310_6
timestamp 1731220585
transform 1 0 1232 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5309_6
timestamp 1731220585
transform 1 0 1320 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5308_6
timestamp 1731220585
transform 1 0 1408 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5307_6
timestamp 1731220585
transform 1 0 1496 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5306_6
timestamp 1731220585
transform 1 0 1576 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5305_6
timestamp 1731220585
transform 1 0 1656 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5304_6
timestamp 1731220585
transform 1 0 1736 0 1 88
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5303_6
timestamp 1731220585
transform 1 0 1888 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5302_6
timestamp 1731220585
transform 1 0 1968 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5301_6
timestamp 1731220585
transform 1 0 2072 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5300_6
timestamp 1731220585
transform 1 0 2448 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5299_6
timestamp 1731220585
transform 1 0 2320 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5298_6
timestamp 1731220585
transform 1 0 2192 0 1 108
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5297_6
timestamp 1731220585
transform 1 0 2088 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5296_6
timestamp 1731220585
transform 1 0 1976 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5295_6
timestamp 1731220585
transform 1 0 1888 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5294_6
timestamp 1731220585
transform 1 0 2496 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5293_6
timestamp 1731220585
transform 1 0 2352 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5292_6
timestamp 1731220585
transform 1 0 2216 0 -1 272
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5291_6
timestamp 1731220585
transform 1 0 2152 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5290_6
timestamp 1731220585
transform 1 0 2064 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5289_6
timestamp 1731220585
transform 1 0 2248 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5288_6
timestamp 1731220585
transform 1 0 2360 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5287_6
timestamp 1731220585
transform 1 0 2624 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5286_6
timestamp 1731220585
transform 1 0 2488 0 1 280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5285_6
timestamp 1731220585
transform 1 0 2408 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5284_6
timestamp 1731220585
transform 1 0 2328 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5283_6
timestamp 1731220585
transform 1 0 2488 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5282_6
timestamp 1731220585
transform 1 0 2576 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5281_6
timestamp 1731220585
transform 1 0 2680 0 -1 440
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5280_6
timestamp 1731220585
transform 1 0 2672 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5279_6
timestamp 1731220585
transform 1 0 2536 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5278_6
timestamp 1731220585
transform 1 0 2416 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5277_6
timestamp 1731220585
transform 1 0 2312 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5276_6
timestamp 1731220585
transform 1 0 2216 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5275_6
timestamp 1731220585
transform 1 0 2136 0 1 444
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5274_6
timestamp 1731220585
transform 1 0 2488 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5273_6
timestamp 1731220585
transform 1 0 2344 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5272_6
timestamp 1731220585
transform 1 0 2208 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5271_6
timestamp 1731220585
transform 1 0 2080 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5270_6
timestamp 1731220585
transform 1 0 1968 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5269_6
timestamp 1731220585
transform 1 0 1888 0 -1 596
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5268_6
timestamp 1731220585
transform 1 0 1888 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5267_6
timestamp 1731220585
transform 1 0 1736 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5266_6
timestamp 1731220585
transform 1 0 1648 0 1 620
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5265_6
timestamp 1731220585
transform 1 0 2280 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5264_6
timestamp 1731220585
transform 1 0 2080 0 1 600
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5263_6
timestamp 1731220585
transform 1 0 2064 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5262_6
timestamp 1731220585
transform 1 0 1968 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5261_6
timestamp 1731220585
transform 1 0 1888 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5260_6
timestamp 1731220585
transform 1 0 2176 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5259_6
timestamp 1731220585
transform 1 0 2440 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5258_6
timestamp 1731220585
transform 1 0 2304 0 -1 756
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5257_6
timestamp 1731220585
transform 1 0 2232 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5256_6
timestamp 1731220585
transform 1 0 2152 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5255_6
timestamp 1731220585
transform 1 0 2312 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5254_6
timestamp 1731220585
transform 1 0 2640 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5253_6
timestamp 1731220585
transform 1 0 2520 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5252_6
timestamp 1731220585
transform 1 0 2408 0 1 764
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5251_6
timestamp 1731220585
transform 1 0 2352 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5250_6
timestamp 1731220585
transform 1 0 2272 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5249_6
timestamp 1731220585
transform 1 0 2432 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5248_6
timestamp 1731220585
transform 1 0 2512 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5247_6
timestamp 1731220585
transform 1 0 2600 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5246_6
timestamp 1731220585
transform 1 0 2696 0 -1 928
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5245_6
timestamp 1731220585
transform 1 0 2656 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5244_6
timestamp 1731220585
transform 1 0 2552 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5243_6
timestamp 1731220585
transform 1 0 2456 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5242_6
timestamp 1731220585
transform 1 0 2368 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5241_6
timestamp 1731220585
transform 1 0 2288 0 1 936
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5240_6
timestamp 1731220585
transform 1 0 2600 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5239_6
timestamp 1731220585
transform 1 0 2472 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5238_6
timestamp 1731220585
transform 1 0 2352 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5237_6
timestamp 1731220585
transform 1 0 2248 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5236_6
timestamp 1731220585
transform 1 0 2160 0 -1 1088
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5235_6
timestamp 1731220585
transform 1 0 2512 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5234_6
timestamp 1731220585
transform 1 0 2352 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5233_6
timestamp 1731220585
transform 1 0 2200 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5232_6
timestamp 1731220585
transform 1 0 2072 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5231_6
timestamp 1731220585
transform 1 0 1968 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5230_6
timestamp 1731220585
transform 1 0 1888 0 1 1096
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5229_6
timestamp 1731220585
transform 1 0 1888 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5228_6
timestamp 1731220585
transform 1 0 1736 0 1 1128
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5227_6
timestamp 1731220585
transform 1 0 1736 0 -1 1280
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5226_6
timestamp 1731220585
transform 1 0 2064 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5225_6
timestamp 1731220585
transform 1 0 2264 0 -1 1252
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5224_6
timestamp 1731220585
transform 1 0 2168 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5223_6
timestamp 1731220585
transform 1 0 2032 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5222_6
timestamp 1731220585
transform 1 0 1912 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5221_6
timestamp 1731220585
transform 1 0 2304 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5220_6
timestamp 1731220585
transform 1 0 2440 0 1 1260
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5219_6
timestamp 1731220585
transform 1 0 2296 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5218_6
timestamp 1731220585
transform 1 0 2160 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5217_6
timestamp 1731220585
transform 1 0 2016 0 -1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5216_6
timestamp 1731220585
transform 1 0 2256 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5215_6
timestamp 1731220585
transform 1 0 2400 0 1 1420
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5214_6
timestamp 1731220585
transform 1 0 2360 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5213_6
timestamp 1731220585
transform 1 0 2520 0 -1 1580
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5212_6
timestamp 1731220585
transform 1 0 2480 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5211_6
timestamp 1731220585
transform 1 0 2624 0 1 1588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5210_6
timestamp 1731220585
transform 1 0 2520 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5209_6
timestamp 1731220585
transform 1 0 2656 0 -1 1744
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5208_6
timestamp 1731220585
transform 1 0 2704 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5207_6
timestamp 1731220585
transform 1 0 2544 0 1 1748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5206_6
timestamp 1731220585
transform 1 0 2232 0 -1 1916
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5205_6
timestamp 1731220585
transform 1 0 2304 0 1 1924
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5204_6
timestamp 1731220585
transform 1 0 2208 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5203_6
timestamp 1731220585
transform 1 0 2440 0 -1 2076
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5202_6
timestamp 1731220585
transform 1 0 2528 0 1 2084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5201_6
timestamp 1731220585
transform 1 0 2488 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5200_6
timestamp 1731220585
transform 1 0 2392 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5199_6
timestamp 1731220585
transform 1 0 2304 0 -1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5198_6
timestamp 1731220585
transform 1 0 2504 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5197_6
timestamp 1731220585
transform 1 0 2424 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5196_6
timestamp 1731220585
transform 1 0 2344 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5195_6
timestamp 1731220585
transform 1 0 2264 0 1 2240
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5194_6
timestamp 1731220585
transform 1 0 2568 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5193_6
timestamp 1731220585
transform 1 0 2448 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5192_6
timestamp 1731220585
transform 1 0 2336 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5191_6
timestamp 1731220585
transform 1 0 2232 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5190_6
timestamp 1731220585
transform 1 0 2136 0 -1 2396
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5189_6
timestamp 1731220585
transform 1 0 2536 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5188_6
timestamp 1731220585
transform 1 0 2392 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5187_6
timestamp 1731220585
transform 1 0 2248 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5186_6
timestamp 1731220585
transform 1 0 2112 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5185_6
timestamp 1731220585
transform 1 0 1984 0 1 2400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5184_6
timestamp 1731220585
transform 1 0 2464 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5183_6
timestamp 1731220585
transform 1 0 2312 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5182_6
timestamp 1731220585
transform 1 0 2152 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5181_6
timestamp 1731220585
transform 1 0 2000 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5180_6
timestamp 1731220585
transform 1 0 1888 0 -1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5179_6
timestamp 1731220585
transform 1 0 2736 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5178_6
timestamp 1731220585
transform 1 0 2480 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5177_6
timestamp 1731220585
transform 1 0 2248 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5176_6
timestamp 1731220585
transform 1 0 2040 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5175_6
timestamp 1731220585
transform 1 0 1888 0 1 2560
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5174_6
timestamp 1731220585
transform 1 0 2528 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5173_6
timestamp 1731220585
transform 1 0 2320 0 -1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5172_6
timestamp 1731220585
transform 1 0 2312 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5171_6
timestamp 1731220585
transform 1 0 2152 0 1 2720
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5170_6
timestamp 1731220585
transform 1 0 2128 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5169_6
timestamp 1731220585
transform 1 0 2040 0 -1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5168_6
timestamp 1731220585
transform 1 0 2112 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5167_6
timestamp 1731220585
transform 1 0 2192 0 1 2884
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5166_6
timestamp 1731220585
transform 1 0 2192 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5165_6
timestamp 1731220585
transform 1 0 2472 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5164_6
timestamp 1731220585
transform 1 0 2328 0 -1 3048
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5163_6
timestamp 1731220585
transform 1 0 2248 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5162_6
timestamp 1731220585
transform 1 0 2056 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5161_6
timestamp 1731220585
transform 1 0 2440 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5160_6
timestamp 1731220585
transform 1 0 2448 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5159_6
timestamp 1731220585
transform 1 0 2288 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5158_6
timestamp 1731220585
transform 1 0 2304 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5157_6
timestamp 1731220585
transform 1 0 2432 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5156_6
timestamp 1731220585
transform 1 0 2432 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5155_6
timestamp 1731220585
transform 1 0 2576 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5154_6
timestamp 1731220585
transform 1 0 2664 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5153_6
timestamp 1731220585
transform 1 0 2520 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5152_6
timestamp 1731220585
transform 1 0 2376 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5151_6
timestamp 1731220585
transform 1 0 2328 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5150_6
timestamp 1731220585
transform 1 0 2504 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5149_6
timestamp 1731220585
transform 1 0 2544 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5148_6
timestamp 1731220585
transform 1 0 2408 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5147_6
timestamp 1731220585
transform 1 0 2280 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5146_6
timestamp 1731220585
transform 1 0 2144 0 -1 3668
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5145_6
timestamp 1731220585
transform 1 0 2160 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5144_6
timestamp 1731220585
transform 1 0 2056 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5143_6
timestamp 1731220585
transform 1 0 1968 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5142_6
timestamp 1731220585
transform 1 0 1888 0 1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5141_6
timestamp 1731220585
transform 1 0 1960 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5140_6
timestamp 1731220585
transform 1 0 2144 0 -1 3516
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5139_6
timestamp 1731220585
transform 1 0 2112 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5138_6
timestamp 1731220585
transform 1 0 1992 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5137_6
timestamp 1731220585
transform 1 0 2240 0 1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5136_6
timestamp 1731220585
transform 1 0 2288 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5135_6
timestamp 1731220585
transform 1 0 2144 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5134_6
timestamp 1731220585
transform 1 0 2008 0 -1 3364
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5133_6
timestamp 1731220585
transform 1 0 1912 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5132_6
timestamp 1731220585
transform 1 0 2048 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5131_6
timestamp 1731220585
transform 1 0 2176 0 1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5130_6
timestamp 1731220585
transform 1 0 2136 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5129_6
timestamp 1731220585
transform 1 0 2000 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5128_6
timestamp 1731220585
transform 1 0 1888 0 -1 3212
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5127_6
timestamp 1731220585
transform 1 0 1888 0 1 3060
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5126_6
timestamp 1731220585
transform 1 0 1736 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5125_6
timestamp 1731220585
transform 1 0 1656 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5124_6
timestamp 1731220585
transform 1 0 1568 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5123_6
timestamp 1731220585
transform 1 0 1480 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5122_6
timestamp 1731220585
transform 1 0 1392 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5121_6
timestamp 1731220585
transform 1 0 1296 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5120_6
timestamp 1731220585
transform 1 0 1192 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5119_6
timestamp 1731220585
transform 1 0 1088 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5118_6
timestamp 1731220585
transform 1 0 976 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5117_6
timestamp 1731220585
transform 1 0 856 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5116_6
timestamp 1731220585
transform 1 0 1600 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5115_6
timestamp 1731220585
transform 1 0 1456 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5114_6
timestamp 1731220585
transform 1 0 1320 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5113_6
timestamp 1731220585
transform 1 0 1184 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5112_6
timestamp 1731220585
transform 1 0 1040 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5111_6
timestamp 1731220585
transform 1 0 1456 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5110_6
timestamp 1731220585
transform 1 0 1328 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5109_6
timestamp 1731220585
transform 1 0 1200 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5108_6
timestamp 1731220585
transform 1 0 1072 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5107_6
timestamp 1731220585
transform 1 0 936 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5106_6
timestamp 1731220585
transform 1 0 1344 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5105_6
timestamp 1731220585
transform 1 0 1232 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5104_6
timestamp 1731220585
transform 1 0 1120 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5103_6
timestamp 1731220585
transform 1 0 1008 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5102_6
timestamp 1731220585
transform 1 0 888 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5101_6
timestamp 1731220585
transform 1 0 1312 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_5100_6
timestamp 1731220585
transform 1 0 1216 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_599_6
timestamp 1731220585
transform 1 0 1120 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_598_6
timestamp 1731220585
transform 1 0 1024 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_597_6
timestamp 1731220585
transform 1 0 928 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_596_6
timestamp 1731220585
transform 1 0 1440 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_595_6
timestamp 1731220585
transform 1 0 1352 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_594_6
timestamp 1731220585
transform 1 0 1264 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_593_6
timestamp 1731220585
transform 1 0 1176 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_592_6
timestamp 1731220585
transform 1 0 1088 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_591_6
timestamp 1731220585
transform 1 0 1000 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_590_6
timestamp 1731220585
transform 1 0 1184 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_589_6
timestamp 1731220585
transform 1 0 1040 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_588_6
timestamp 1731220585
transform 1 0 896 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_587_6
timestamp 1731220585
transform 1 0 760 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_586_6
timestamp 1731220585
transform 1 0 912 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_585_6
timestamp 1731220585
transform 1 0 824 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_584_6
timestamp 1731220585
transform 1 0 728 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_583_6
timestamp 1731220585
transform 1 0 624 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_582_6
timestamp 1731220585
transform 1 0 520 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_581_6
timestamp 1731220585
transform 1 0 824 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_580_6
timestamp 1731220585
transform 1 0 720 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_579_6
timestamp 1731220585
transform 1 0 608 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_578_6
timestamp 1731220585
transform 1 0 488 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_577_6
timestamp 1731220585
transform 1 0 504 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_576_6
timestamp 1731220585
transform 1 0 640 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_575_6
timestamp 1731220585
transform 1 0 768 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_574_6
timestamp 1731220585
transform 1 0 800 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_573_6
timestamp 1731220585
transform 1 0 656 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_572_6
timestamp 1731220585
transform 1 0 504 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_571_6
timestamp 1731220585
transform 1 0 568 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_570_6
timestamp 1731220585
transform 1 0 728 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_569_6
timestamp 1731220585
transform 1 0 888 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_568_6
timestamp 1731220585
transform 1 0 728 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_567_6
timestamp 1731220585
transform 1 0 592 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_566_6
timestamp 1731220585
transform 1 0 448 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_565_6
timestamp 1731220585
transform 1 0 432 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_564_6
timestamp 1731220585
transform 1 0 544 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_563_6
timestamp 1731220585
transform 1 0 656 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_562_6
timestamp 1731220585
transform 1 0 784 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_561_6
timestamp 1731220585
transform 1 0 632 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_560_6
timestamp 1731220585
transform 1 0 472 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_559_6
timestamp 1731220585
transform 1 0 464 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_558_6
timestamp 1731220585
transform 1 0 624 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_557_6
timestamp 1731220585
transform 1 0 776 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_556_6
timestamp 1731220585
transform 1 0 832 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_555_6
timestamp 1731220585
transform 1 0 672 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_554_6
timestamp 1731220585
transform 1 0 520 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_553_6
timestamp 1731220585
transform 1 0 504 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_552_6
timestamp 1731220585
transform 1 0 656 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_551_6
timestamp 1731220585
transform 1 0 808 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_550_6
timestamp 1731220585
transform 1 0 776 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_549_6
timestamp 1731220585
transform 1 0 608 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_548_6
timestamp 1731220585
transform 1 0 520 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_547_6
timestamp 1731220585
transform 1 0 696 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_546_6
timestamp 1731220585
transform 1 0 872 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_545_6
timestamp 1731220585
transform 1 0 912 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_544_6
timestamp 1731220585
transform 1 0 768 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_543_6
timestamp 1731220585
transform 1 0 632 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_542_6
timestamp 1731220585
transform 1 0 496 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_541_6
timestamp 1731220585
transform 1 0 376 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_540_6
timestamp 1731220585
transform 1 0 288 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_539_6
timestamp 1731220585
transform 1 0 208 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_538_6
timestamp 1731220585
transform 1 0 128 0 1 2428
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_537_6
timestamp 1731220585
transform 1 0 128 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_536_6
timestamp 1731220585
transform 1 0 216 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_535_6
timestamp 1731220585
transform 1 0 360 0 -1 2584
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_534_6
timestamp 1731220585
transform 1 0 432 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_533_6
timestamp 1731220585
transform 1 0 264 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_532_6
timestamp 1731220585
transform 1 0 128 0 1 2588
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_531_6
timestamp 1731220585
transform 1 0 128 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_530_6
timestamp 1731220585
transform 1 0 224 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_529_6
timestamp 1731220585
transform 1 0 360 0 -1 2748
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_528_6
timestamp 1731220585
transform 1 0 368 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_527_6
timestamp 1731220585
transform 1 0 232 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_526_6
timestamp 1731220585
transform 1 0 128 0 1 2752
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_525_6
timestamp 1731220585
transform 1 0 144 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_524_6
timestamp 1731220585
transform 1 0 304 0 -1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_523_6
timestamp 1731220585
transform 1 0 304 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_522_6
timestamp 1731220585
transform 1 0 144 0 1 2908
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_521_6
timestamp 1731220585
transform 1 0 128 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_520_6
timestamp 1731220585
transform 1 0 216 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_519_6
timestamp 1731220585
transform 1 0 320 0 -1 3072
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_518_6
timestamp 1731220585
transform 1 0 304 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_517_6
timestamp 1731220585
transform 1 0 160 0 1 3084
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_516_6
timestamp 1731220585
transform 1 0 128 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_515_6
timestamp 1731220585
transform 1 0 408 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_514_6
timestamp 1731220585
transform 1 0 264 0 -1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_513_6
timestamp 1731220585
transform 1 0 192 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_512_6
timestamp 1731220585
transform 1 0 352 0 1 3244
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_511_6
timestamp 1731220585
transform 1 0 360 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_510_6
timestamp 1731220585
transform 1 0 208 0 -1 3400
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_59_6
timestamp 1731220585
transform 1 0 216 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_58_6
timestamp 1731220585
transform 1 0 352 0 1 3404
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_57_6
timestamp 1731220585
transform 1 0 296 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_56_6
timestamp 1731220585
transform 1 0 176 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_55_6
timestamp 1731220585
transform 1 0 408 0 -1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_54_6
timestamp 1731220585
transform 1 0 624 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_53_6
timestamp 1731220585
transform 1 0 488 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_52_6
timestamp 1731220585
transform 1 0 352 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_51_6
timestamp 1731220585
transform 1 0 224 0 1 3564
box 8 4 70 72
use _0_0std_0_0cells_0_0LATCHINV  tst_50_6
timestamp 1731220585
transform 1 0 128 0 1 3564
box 8 4 70 72
<< end >>
