magic
tech sky130l
timestamp 1731220370
<< m1 >>
rect 3416 3843 3420 3867
rect 2168 3735 2172 3759
rect 1104 3679 1108 3731
rect 2624 3679 2628 3703
rect 936 3651 940 3675
rect 3424 3567 3428 3591
rect 2776 3375 2780 3423
rect 720 3315 724 3339
rect 2552 3235 2556 3259
rect 744 3191 748 3223
rect 2856 3191 2860 3227
rect 3128 3191 3132 3215
rect 3424 2919 3428 3027
rect 2600 2699 2604 2723
rect 2792 2699 2796 2739
rect 3256 2423 3260 2447
rect 816 2195 820 2219
rect 776 2063 780 2111
rect 2624 2031 2628 2055
rect 3560 2031 3564 2055
rect 3512 1919 3516 1943
rect 760 1867 764 1891
rect 872 1867 876 1911
rect 1168 1867 1172 1911
rect 2744 1871 2748 1895
rect 1616 1759 1620 1783
rect 2608 1763 2612 1787
rect 1296 1603 1300 1627
rect 3128 1611 3132 1635
rect 3640 1587 3644 1635
rect 976 1447 980 1471
rect 2896 1459 2900 1555
rect 1800 1291 1804 1315
rect 3568 1291 3572 1315
rect 512 1243 516 1267
rect 1888 1243 1892 1283
rect 3232 1247 3236 1279
rect 1048 1135 1052 1159
rect 1536 1115 1540 1159
rect 3224 1139 3228 1239
rect 2448 959 2452 1003
rect 3592 979 3596 1003
rect 3224 931 3228 955
rect 3400 931 3404 955
rect 944 823 948 847
rect 2336 807 2340 847
rect 256 775 260 799
rect 1104 667 1108 691
rect 2200 667 2204 691
rect 2680 667 2684 775
rect 1392 623 1396 659
rect 472 495 476 535
rect 576 511 580 535
rect 1520 511 1524 535
rect 2184 511 2188 535
rect 2696 511 2700 535
rect 3448 511 3452 535
rect 3584 511 3588 535
rect 1032 359 1036 383
rect 152 311 156 351
rect 376 223 380 335
rect 640 195 644 219
rect 1296 195 1300 219
rect 1472 195 1476 219
rect 3416 127 3420 151
rect 3624 127 3628 151
rect 3632 127 3636 195
<< m2c >>
rect 2108 4019 2112 4023
rect 316 3999 320 4003
rect 468 3999 472 4003
rect 644 3999 648 4003
rect 828 3999 832 4003
rect 1012 3999 1016 4003
rect 1188 3997 1192 4001
rect 1348 3999 1352 4003
rect 1508 3999 1512 4003
rect 1660 3999 1664 4003
rect 1812 3999 1816 4003
rect 1940 3999 1944 4003
rect 2116 3883 2120 3887
rect 2252 3883 2256 3887
rect 2396 3883 2400 3887
rect 2540 3883 2544 3887
rect 2684 3883 2688 3887
rect 2964 3883 2968 3887
rect 3092 3883 3096 3887
rect 3212 3883 3216 3887
rect 3332 3883 3336 3887
rect 3452 3883 3456 3887
rect 3572 3883 3576 3887
rect 2828 3879 2832 3883
rect 340 3863 344 3867
rect 460 3863 464 3867
rect 588 3863 592 3867
rect 724 3863 728 3867
rect 852 3863 856 3867
rect 1108 3863 1112 3867
rect 1236 3863 1240 3867
rect 1364 3863 1368 3867
rect 1500 3863 1504 3867
rect 2292 3865 2296 3869
rect 2420 3867 2424 3871
rect 2556 3867 2560 3871
rect 2708 3867 2712 3871
rect 2868 3867 2872 3871
rect 3028 3867 3032 3871
rect 3196 3867 3200 3871
rect 3364 3867 3368 3871
rect 3416 3867 3420 3871
rect 3532 3867 3536 3871
rect 3700 3867 3704 3871
rect 980 3859 984 3863
rect 452 3845 456 3849
rect 604 3843 608 3847
rect 764 3843 768 3847
rect 924 3843 928 3847
rect 1076 3843 1080 3847
rect 1228 3843 1232 3847
rect 1380 3843 1384 3847
rect 1532 3843 1536 3847
rect 1684 3843 1688 3847
rect 3416 3839 3420 3843
rect 2168 3759 2172 3763
rect 1104 3731 1108 3735
rect 2108 3731 2112 3735
rect 2168 3731 2172 3735
rect 2236 3731 2240 3735
rect 2412 3731 2416 3735
rect 2596 3731 2600 3735
rect 2788 3731 2792 3735
rect 2988 3731 2992 3735
rect 3372 3731 3376 3735
rect 3572 3731 3576 3735
rect 3772 3731 3776 3735
rect 436 3703 440 3707
rect 604 3703 608 3707
rect 788 3703 792 3707
rect 972 3703 976 3707
rect 404 3677 408 3681
rect 3180 3727 3184 3731
rect 1164 3703 1168 3707
rect 1348 3703 1352 3707
rect 1540 3703 1544 3707
rect 1732 3703 1736 3707
rect 2108 3703 2112 3707
rect 2300 3703 2304 3707
rect 2516 3703 2520 3707
rect 2624 3703 2628 3707
rect 2732 3703 2736 3707
rect 1924 3699 1928 3703
rect 556 3675 560 3679
rect 716 3675 720 3679
rect 884 3675 888 3679
rect 936 3675 940 3679
rect 1052 3675 1056 3679
rect 1104 3675 1108 3679
rect 1212 3677 1216 3681
rect 2948 3701 2952 3705
rect 3156 3703 3160 3707
rect 3356 3701 3360 3705
rect 3556 3703 3560 3707
rect 3764 3703 3768 3707
rect 1364 3675 1368 3679
rect 1516 3675 1520 3679
rect 1668 3675 1672 3679
rect 1828 3675 1832 3679
rect 2624 3675 2628 3679
rect 936 3647 940 3651
rect 3424 3591 3428 3595
rect 2148 3563 2152 3567
rect 2308 3563 2312 3567
rect 2492 3563 2496 3567
rect 2692 3563 2696 3567
rect 2908 3563 2912 3567
rect 3364 3563 3368 3567
rect 3424 3563 3428 3567
rect 3604 3563 3608 3567
rect 3132 3559 3136 3563
rect 308 3531 312 3535
rect 452 3531 456 3535
rect 612 3531 616 3535
rect 772 3531 776 3535
rect 932 3531 936 3535
rect 1252 3531 1256 3535
rect 1412 3531 1416 3535
rect 1580 3531 1584 3535
rect 2324 3531 2328 3535
rect 2420 3531 2424 3535
rect 2516 3531 2520 3535
rect 2612 3531 2616 3535
rect 2708 3531 2712 3535
rect 2804 3531 2808 3535
rect 2908 3531 2912 3535
rect 3020 3531 3024 3535
rect 3140 3531 3144 3535
rect 3260 3531 3264 3535
rect 3388 3531 3392 3535
rect 3524 3531 3528 3535
rect 1092 3527 1096 3531
rect 196 3505 200 3509
rect 324 3507 328 3511
rect 460 3507 464 3511
rect 596 3507 600 3511
rect 732 3507 736 3511
rect 868 3507 872 3511
rect 1004 3507 1008 3511
rect 1132 3507 1136 3511
rect 1268 3507 1272 3511
rect 1404 3507 1408 3511
rect 2776 3423 2780 3427
rect 2524 3395 2528 3399
rect 2620 3395 2624 3399
rect 2716 3395 2720 3399
rect 2820 3395 2824 3399
rect 2932 3395 2936 3399
rect 3052 3395 3056 3399
rect 3308 3395 3312 3399
rect 3444 3395 3448 3399
rect 3180 3391 3184 3395
rect 2388 3369 2392 3373
rect 2516 3371 2520 3375
rect 2652 3371 2656 3375
rect 2776 3371 2780 3375
rect 2788 3371 2792 3375
rect 2924 3371 2928 3375
rect 3060 3371 3064 3375
rect 3196 3371 3200 3375
rect 3340 3371 3344 3375
rect 172 3363 176 3367
rect 284 3363 288 3367
rect 420 3363 424 3367
rect 564 3363 568 3367
rect 708 3363 712 3367
rect 852 3363 856 3367
rect 1004 3363 1008 3367
rect 1308 3363 1312 3367
rect 1156 3359 1160 3363
rect 172 3339 176 3343
rect 300 3339 304 3343
rect 468 3339 472 3343
rect 636 3339 640 3343
rect 720 3339 724 3343
rect 804 3339 808 3343
rect 964 3337 968 3341
rect 1124 3339 1128 3343
rect 1276 3339 1280 3343
rect 1428 3339 1432 3343
rect 1588 3339 1592 3343
rect 720 3311 724 3315
rect 2552 3259 2556 3263
rect 2164 3231 2168 3235
rect 2332 3231 2336 3235
rect 2492 3231 2496 3235
rect 2552 3231 2556 3235
rect 2652 3231 2656 3235
rect 2972 3231 2976 3235
rect 3132 3231 3136 3235
rect 3300 3231 3304 3235
rect 2812 3227 2816 3231
rect 2856 3227 2860 3231
rect 744 3223 748 3227
rect 180 3195 184 3199
rect 332 3195 336 3199
rect 492 3195 496 3199
rect 660 3195 664 3199
rect 2108 3213 2112 3217
rect 2244 3215 2248 3219
rect 2412 3215 2416 3219
rect 2580 3215 2584 3219
rect 2740 3215 2744 3219
rect 828 3195 832 3199
rect 1164 3195 1168 3199
rect 1340 3195 1344 3199
rect 1516 3195 1520 3199
rect 996 3191 1000 3195
rect 2900 3215 2904 3219
rect 3052 3215 3056 3219
rect 3128 3215 3132 3219
rect 3204 3215 3208 3219
rect 3364 3215 3368 3219
rect 744 3187 748 3191
rect 2856 3187 2860 3191
rect 3128 3187 3132 3191
rect 332 3181 336 3185
rect 468 3179 472 3183
rect 604 3179 608 3183
rect 740 3179 744 3183
rect 892 3179 896 3183
rect 1068 3179 1072 3183
rect 1268 3179 1272 3183
rect 1492 3179 1496 3183
rect 1724 3179 1728 3183
rect 1940 3179 1944 3183
rect 2108 3075 2112 3079
rect 2668 3075 2672 3079
rect 2940 3075 2944 3079
rect 3212 3075 3216 3079
rect 3484 3075 3488 3079
rect 2380 3071 2384 3075
rect 2524 3055 2528 3059
rect 2652 3055 2656 3059
rect 2780 3055 2784 3059
rect 2900 3055 2904 3059
rect 3020 3055 3024 3059
rect 3140 3055 3144 3059
rect 3252 3055 3256 3059
rect 3364 3055 3368 3059
rect 3468 3055 3472 3059
rect 3572 3055 3576 3059
rect 3676 3055 3680 3059
rect 3780 3055 3784 3059
rect 3876 3055 3880 3059
rect 348 3043 352 3047
rect 444 3043 448 3047
rect 540 3043 544 3047
rect 636 3043 640 3047
rect 732 3043 736 3047
rect 844 3043 848 3047
rect 1124 3043 1128 3047
rect 1284 3043 1288 3047
rect 1444 3043 1448 3047
rect 1612 3043 1616 3047
rect 1788 3043 1792 3047
rect 1940 3043 1944 3047
rect 980 3039 984 3043
rect 460 3027 464 3031
rect 556 3027 560 3031
rect 652 3027 656 3031
rect 748 3027 752 3031
rect 852 3027 856 3031
rect 972 3027 976 3031
rect 1092 3027 1096 3031
rect 1220 3027 1224 3031
rect 1348 3027 1352 3031
rect 1468 3027 1472 3031
rect 1588 3027 1592 3031
rect 1708 3025 1712 3029
rect 1836 3027 1840 3031
rect 1940 3027 1944 3031
rect 3424 3027 3428 3031
rect 2444 2915 2448 2919
rect 2612 2915 2616 2919
rect 2804 2915 2808 2919
rect 3004 2915 3008 2919
rect 3424 2915 3428 2919
rect 3436 2915 3440 2919
rect 3660 2915 3664 2919
rect 3876 2915 3880 2919
rect 3220 2911 3224 2915
rect 2588 2881 2592 2885
rect 2708 2883 2712 2887
rect 2836 2883 2840 2887
rect 2964 2883 2968 2887
rect 3092 2883 3096 2887
rect 3220 2883 3224 2887
rect 3348 2881 3352 2885
rect 3476 2883 3480 2887
rect 3612 2883 3616 2887
rect 1516 2867 1520 2871
rect 1612 2867 1616 2871
rect 1708 2867 1712 2871
rect 1804 2867 1808 2871
rect 1900 2867 1904 2871
rect 484 2845 488 2849
rect 316 2841 320 2845
rect 668 2843 672 2847
rect 852 2843 856 2847
rect 1036 2843 1040 2847
rect 1220 2841 1224 2845
rect 1396 2843 1400 2847
rect 1564 2843 1568 2847
rect 1732 2843 1736 2847
rect 1900 2843 1904 2847
rect 2604 2747 2608 2751
rect 2732 2747 2736 2751
rect 2868 2747 2872 2751
rect 3004 2747 3008 2751
rect 3140 2747 3144 2751
rect 3284 2747 3288 2751
rect 3428 2747 3432 2751
rect 3580 2747 3584 2751
rect 3876 2747 3880 2751
rect 2476 2743 2480 2747
rect 3740 2743 3744 2747
rect 2792 2739 2796 2743
rect 2372 2723 2376 2727
rect 2532 2723 2536 2727
rect 2600 2723 2604 2727
rect 2700 2723 2704 2727
rect 388 2707 392 2711
rect 508 2707 512 2711
rect 644 2707 648 2711
rect 780 2707 784 2711
rect 916 2707 920 2711
rect 1052 2707 1056 2711
rect 1188 2707 1192 2711
rect 1324 2707 1328 2711
rect 1460 2707 1464 2711
rect 1604 2707 1608 2711
rect 276 2703 280 2707
rect 2600 2695 2604 2699
rect 2868 2723 2872 2727
rect 3036 2721 3040 2725
rect 3204 2723 3208 2727
rect 3372 2723 3376 2727
rect 3548 2723 3552 2727
rect 3724 2723 3728 2727
rect 3876 2723 3880 2727
rect 2792 2695 2796 2699
rect 260 2691 264 2695
rect 404 2691 408 2695
rect 540 2691 544 2695
rect 676 2691 680 2695
rect 804 2691 808 2695
rect 924 2691 928 2695
rect 1036 2691 1040 2695
rect 1148 2689 1152 2693
rect 1268 2691 1272 2695
rect 1388 2691 1392 2695
rect 2316 2583 2320 2587
rect 2484 2583 2488 2587
rect 2660 2583 2664 2587
rect 2844 2583 2848 2587
rect 3028 2583 3032 2587
rect 3212 2583 3216 2587
rect 3388 2583 3392 2587
rect 3556 2583 3560 2587
rect 3876 2583 3880 2587
rect 2164 2579 2168 2583
rect 3724 2579 3728 2583
rect 404 2555 408 2559
rect 580 2555 584 2559
rect 748 2555 752 2559
rect 900 2555 904 2559
rect 1044 2555 1048 2559
rect 1180 2555 1184 2559
rect 1316 2555 1320 2559
rect 1460 2555 1464 2559
rect 2108 2557 2112 2561
rect 2220 2559 2224 2563
rect 2356 2559 2360 2563
rect 2508 2559 2512 2563
rect 2676 2559 2680 2563
rect 2860 2559 2864 2563
rect 3068 2559 3072 2563
rect 3300 2559 3304 2563
rect 3540 2559 3544 2563
rect 3780 2559 3784 2563
rect 212 2551 216 2555
rect 172 2535 176 2539
rect 308 2535 312 2539
rect 476 2535 480 2539
rect 644 2535 648 2539
rect 812 2535 816 2539
rect 964 2535 968 2539
rect 1116 2537 1120 2541
rect 1260 2535 1264 2539
rect 1396 2535 1400 2539
rect 1532 2535 1536 2539
rect 1676 2535 1680 2539
rect 3256 2447 3260 2451
rect 2108 2419 2112 2423
rect 2252 2419 2256 2423
rect 2420 2419 2424 2423
rect 2596 2419 2600 2423
rect 2788 2419 2792 2423
rect 2988 2419 2992 2423
rect 3204 2419 3208 2423
rect 3256 2419 3260 2423
rect 3428 2419 3432 2423
rect 3876 2419 3880 2423
rect 3660 2415 3664 2419
rect 348 2395 352 2399
rect 548 2395 552 2399
rect 748 2395 752 2399
rect 940 2395 944 2399
rect 1116 2395 1120 2399
rect 1276 2395 1280 2399
rect 1428 2395 1432 2399
rect 1564 2395 1568 2399
rect 1828 2395 1832 2399
rect 1940 2395 1944 2399
rect 172 2391 176 2395
rect 1700 2391 1704 2395
rect 2108 2387 2112 2391
rect 2284 2387 2288 2391
rect 2468 2387 2472 2391
rect 2644 2387 2648 2391
rect 2812 2387 2816 2391
rect 2972 2387 2976 2391
rect 3140 2387 3144 2391
rect 172 2379 176 2383
rect 364 2379 368 2383
rect 588 2379 592 2383
rect 804 2379 808 2383
rect 1012 2379 1016 2383
rect 1212 2381 1216 2385
rect 1404 2379 1408 2383
rect 1588 2379 1592 2383
rect 1772 2379 1776 2383
rect 1940 2379 1944 2383
rect 2108 2251 2112 2255
rect 2212 2251 2216 2255
rect 2348 2251 2352 2255
rect 2628 2251 2632 2255
rect 2788 2251 2792 2255
rect 2972 2251 2976 2255
rect 3180 2251 3184 2255
rect 3412 2251 3416 2255
rect 3652 2251 3656 2255
rect 3876 2251 3880 2255
rect 2484 2247 2488 2251
rect 172 2235 176 2239
rect 308 2235 312 2239
rect 628 2235 632 2239
rect 788 2235 792 2239
rect 1124 2235 1128 2239
rect 1300 2235 1304 2239
rect 1484 2235 1488 2239
rect 1668 2235 1672 2239
rect 1852 2235 1856 2239
rect 468 2231 472 2235
rect 956 2231 960 2235
rect 2148 2225 2152 2229
rect 2292 2227 2296 2231
rect 2444 2227 2448 2231
rect 2596 2227 2600 2231
rect 2756 2227 2760 2231
rect 2916 2229 2920 2233
rect 3084 2227 3088 2231
rect 3260 2227 3264 2231
rect 3444 2227 3448 2231
rect 3628 2227 3632 2231
rect 3820 2227 3824 2231
rect 196 2217 200 2221
rect 364 2219 368 2223
rect 532 2219 536 2223
rect 716 2219 720 2223
rect 816 2219 820 2223
rect 916 2219 920 2223
rect 1132 2219 1136 2223
rect 1364 2219 1368 2223
rect 1604 2219 1608 2223
rect 1852 2219 1856 2223
rect 816 2191 820 2195
rect 776 2111 780 2115
rect 260 2083 264 2087
rect 396 2083 400 2087
rect 532 2083 536 2087
rect 676 2079 680 2083
rect 820 2083 824 2087
rect 1132 2083 1136 2087
rect 1300 2083 1304 2087
rect 1484 2083 1488 2087
rect 1668 2083 1672 2087
rect 1860 2083 1864 2087
rect 972 2079 976 2083
rect 2324 2079 2328 2083
rect 2468 2079 2472 2083
rect 2620 2079 2624 2083
rect 2772 2079 2776 2083
rect 3084 2079 3088 2083
rect 3244 2079 3248 2083
rect 3404 2079 3408 2083
rect 3564 2079 3568 2083
rect 3732 2079 3736 2083
rect 3876 2079 3880 2083
rect 2924 2075 2928 2079
rect 412 2059 416 2063
rect 532 2059 536 2063
rect 652 2059 656 2063
rect 776 2059 780 2063
rect 788 2059 792 2063
rect 932 2059 936 2063
rect 1084 2059 1088 2063
rect 1252 2059 1256 2063
rect 1436 2059 1440 2063
rect 1620 2059 1624 2063
rect 1812 2059 1816 2063
rect 2540 2055 2544 2059
rect 2624 2055 2628 2059
rect 2708 2055 2712 2059
rect 2876 2055 2880 2059
rect 3044 2055 3048 2059
rect 3204 2057 3208 2061
rect 3348 2055 3352 2059
rect 3492 2055 3496 2059
rect 3560 2055 3564 2059
rect 3628 2055 3632 2059
rect 3764 2055 3768 2059
rect 3876 2055 3880 2059
rect 2624 2027 2628 2031
rect 3560 2027 3564 2031
rect 3512 1943 3516 1947
rect 548 1915 552 1919
rect 660 1915 664 1919
rect 908 1915 912 1919
rect 1044 1915 1048 1919
rect 1316 1915 1320 1919
rect 1452 1915 1456 1919
rect 1596 1915 1600 1919
rect 1740 1915 1744 1919
rect 2532 1915 2536 1919
rect 2628 1915 2632 1919
rect 2732 1915 2736 1919
rect 2844 1915 2848 1919
rect 3084 1915 3088 1919
rect 3212 1915 3216 1919
rect 3332 1915 3336 1919
rect 3452 1915 3456 1919
rect 3512 1915 3516 1919
rect 3580 1915 3584 1919
rect 3708 1915 3712 1919
rect 780 1911 784 1915
rect 872 1911 876 1915
rect 588 1891 592 1895
rect 700 1891 704 1895
rect 760 1891 764 1895
rect 820 1891 824 1895
rect 760 1863 764 1867
rect 1168 1911 1172 1915
rect 1180 1911 1184 1915
rect 2964 1911 2968 1915
rect 3836 1911 3840 1915
rect 948 1891 952 1895
rect 1084 1891 1088 1895
rect 872 1863 876 1867
rect 2108 1895 2112 1899
rect 1212 1891 1216 1895
rect 1348 1891 1352 1895
rect 1484 1891 1488 1895
rect 1620 1891 1624 1895
rect 1756 1891 1760 1895
rect 2284 1893 2288 1897
rect 2476 1895 2480 1899
rect 2660 1895 2664 1899
rect 2744 1895 2748 1899
rect 2828 1895 2832 1899
rect 2996 1897 3000 1901
rect 3164 1895 3168 1899
rect 3340 1895 3344 1899
rect 3524 1895 3528 1899
rect 3708 1895 3712 1899
rect 3876 1895 3880 1899
rect 2744 1867 2748 1871
rect 1168 1863 1172 1867
rect 2608 1787 2612 1791
rect 1616 1783 1620 1787
rect 2132 1759 2136 1763
rect 2268 1759 2272 1763
rect 2404 1759 2408 1763
rect 2548 1759 2552 1763
rect 2608 1759 2612 1763
rect 2892 1759 2896 1763
rect 3108 1759 3112 1763
rect 3340 1759 3344 1763
rect 3580 1759 3584 1763
rect 540 1755 544 1759
rect 652 1755 656 1759
rect 900 1755 904 1759
rect 1036 1755 1040 1759
rect 1188 1755 1192 1759
rect 1524 1755 1528 1759
rect 1616 1755 1620 1759
rect 1700 1755 1704 1759
rect 1884 1755 1888 1759
rect 2708 1755 2712 1759
rect 3828 1755 3832 1759
rect 772 1751 776 1755
rect 1356 1751 1360 1755
rect 380 1737 384 1741
rect 500 1739 504 1743
rect 628 1739 632 1743
rect 756 1739 760 1743
rect 884 1741 888 1745
rect 2220 1743 2224 1747
rect 2324 1743 2328 1747
rect 2428 1745 2432 1749
rect 1020 1739 1024 1743
rect 1164 1739 1168 1743
rect 1316 1739 1320 1743
rect 1476 1739 1480 1743
rect 1636 1739 1640 1743
rect 2532 1741 2536 1745
rect 2636 1743 2640 1747
rect 2740 1743 2744 1747
rect 2844 1743 2848 1747
rect 2948 1743 2952 1747
rect 3052 1743 3056 1747
rect 3164 1743 3168 1747
rect 3128 1635 3132 1639
rect 1296 1627 1300 1631
rect 3640 1635 3644 1639
rect 2268 1607 2272 1611
rect 2404 1607 2408 1611
rect 2556 1607 2560 1611
rect 2716 1607 2720 1611
rect 3060 1607 3064 1611
rect 3128 1607 3132 1611
rect 3228 1607 3232 1611
rect 3564 1607 3568 1611
rect 2884 1603 2888 1607
rect 3396 1603 3400 1607
rect 332 1599 336 1603
rect 492 1599 496 1603
rect 660 1599 664 1603
rect 836 1599 840 1603
rect 1020 1599 1024 1603
rect 1204 1599 1208 1603
rect 1296 1599 1300 1603
rect 1580 1599 1584 1603
rect 1772 1599 1776 1603
rect 196 1595 200 1599
rect 1388 1595 1392 1599
rect 3732 1607 3736 1611
rect 3876 1607 3880 1611
rect 172 1583 176 1587
rect 292 1583 296 1587
rect 460 1583 464 1587
rect 644 1583 648 1587
rect 836 1583 840 1587
rect 1028 1583 1032 1587
rect 1220 1583 1224 1587
rect 1404 1583 1408 1587
rect 1588 1583 1592 1587
rect 1772 1583 1776 1587
rect 1940 1581 1944 1585
rect 2108 1583 2112 1587
rect 2308 1583 2312 1587
rect 2532 1583 2536 1587
rect 2748 1583 2752 1587
rect 2948 1583 2952 1587
rect 3132 1583 3136 1587
rect 3300 1583 3304 1587
rect 3460 1583 3464 1587
rect 3604 1583 3608 1587
rect 3640 1583 3644 1587
rect 3748 1583 3752 1587
rect 3876 1583 3880 1587
rect 2896 1555 2900 1559
rect 976 1471 980 1475
rect 2896 1455 2900 1459
rect 2108 1447 2112 1451
rect 2468 1447 2472 1451
rect 2828 1447 2832 1451
rect 3500 1447 3504 1451
rect 3836 1447 3840 1451
rect 284 1443 288 1447
rect 436 1443 440 1447
rect 596 1443 600 1447
rect 756 1443 760 1447
rect 916 1443 920 1447
rect 976 1443 980 1447
rect 1076 1443 1080 1447
rect 1356 1443 1360 1447
rect 1484 1443 1488 1447
rect 1604 1443 1608 1447
rect 1724 1443 1728 1447
rect 1844 1443 1848 1447
rect 1940 1443 1944 1447
rect 3164 1443 3168 1447
rect 172 1439 176 1443
rect 1220 1439 1224 1443
rect 172 1427 176 1431
rect 300 1427 304 1431
rect 468 1425 472 1429
rect 644 1427 648 1431
rect 828 1427 832 1431
rect 1012 1427 1016 1431
rect 1196 1427 1200 1431
rect 1388 1427 1392 1431
rect 1580 1427 1584 1431
rect 1772 1427 1776 1431
rect 1940 1427 1944 1431
rect 2108 1423 2112 1427
rect 2308 1423 2312 1427
rect 2532 1423 2536 1427
rect 2748 1423 2752 1427
rect 2948 1423 2952 1427
rect 3132 1423 3136 1427
rect 3308 1423 3312 1427
rect 3476 1423 3480 1427
rect 3644 1423 3648 1427
rect 3820 1423 3824 1427
rect 1800 1315 1804 1319
rect 3568 1315 3572 1319
rect 196 1287 200 1291
rect 516 1287 520 1291
rect 892 1287 896 1291
rect 1084 1287 1088 1291
rect 1284 1287 1288 1291
rect 1484 1287 1488 1291
rect 1692 1287 1696 1291
rect 1800 1287 1804 1291
rect 2108 1287 2112 1291
rect 2244 1287 2248 1291
rect 2420 1287 2424 1291
rect 2604 1287 2608 1291
rect 2788 1287 2792 1291
rect 2972 1287 2976 1291
rect 3148 1287 3152 1291
rect 3316 1287 3320 1291
rect 3484 1287 3488 1291
rect 3568 1287 3572 1291
rect 348 1283 352 1287
rect 700 1283 704 1287
rect 1888 1283 1892 1287
rect 1900 1283 1904 1287
rect 3660 1283 3664 1287
rect 444 1267 448 1271
rect 512 1267 516 1271
rect 580 1267 584 1271
rect 732 1267 736 1271
rect 892 1267 896 1271
rect 1060 1267 1064 1271
rect 1228 1267 1232 1271
rect 1404 1267 1408 1271
rect 1580 1267 1584 1271
rect 1756 1267 1760 1271
rect 512 1239 516 1243
rect 3232 1279 3236 1283
rect 2188 1273 2192 1277
rect 2324 1271 2328 1275
rect 2468 1271 2472 1275
rect 2620 1271 2624 1275
rect 2780 1271 2784 1275
rect 2940 1271 2944 1275
rect 3108 1271 3112 1275
rect 1932 1267 1936 1271
rect 3284 1271 3288 1275
rect 3468 1271 3472 1275
rect 3652 1271 3656 1275
rect 3844 1271 3848 1275
rect 3232 1243 3236 1247
rect 1888 1239 1892 1243
rect 3224 1239 3228 1243
rect 1048 1159 1052 1163
rect 1536 1159 1540 1163
rect 628 1131 632 1135
rect 796 1131 800 1135
rect 964 1131 968 1135
rect 1048 1131 1052 1135
rect 1284 1131 1288 1135
rect 1436 1131 1440 1135
rect 460 1127 464 1131
rect 1132 1127 1136 1131
rect 412 1111 416 1115
rect 524 1113 528 1117
rect 2348 1135 2352 1139
rect 2452 1135 2456 1139
rect 2564 1135 2568 1139
rect 2676 1135 2680 1139
rect 2804 1135 2808 1139
rect 2948 1135 2952 1139
rect 3108 1135 3112 1139
rect 3224 1135 3228 1139
rect 3284 1135 3288 1139
rect 3476 1135 3480 1139
rect 3868 1135 3872 1139
rect 1724 1131 1728 1135
rect 1876 1131 1880 1135
rect 3668 1131 3672 1135
rect 1580 1127 1584 1131
rect 2444 1115 2448 1119
rect 2540 1115 2544 1119
rect 2636 1115 2640 1119
rect 2732 1115 2736 1119
rect 2844 1115 2848 1119
rect 636 1111 640 1115
rect 748 1111 752 1115
rect 868 1109 872 1113
rect 1004 1111 1008 1115
rect 1156 1111 1160 1115
rect 1316 1111 1320 1115
rect 1484 1111 1488 1115
rect 1536 1111 1540 1115
rect 1660 1111 1664 1115
rect 2980 1113 2984 1117
rect 3132 1115 3136 1119
rect 3300 1115 3304 1119
rect 3484 1115 3488 1119
rect 3676 1115 3680 1119
rect 3876 1115 3880 1119
rect 2448 1003 2452 1007
rect 340 975 344 979
rect 628 975 632 979
rect 764 975 768 979
rect 892 975 896 979
rect 1124 975 1128 979
rect 1236 975 1240 979
rect 1348 975 1352 979
rect 1468 975 1472 979
rect 484 971 488 975
rect 1012 971 1016 975
rect 292 959 296 963
rect 484 959 488 963
rect 668 959 672 963
rect 844 959 848 963
rect 1012 959 1016 963
rect 1164 959 1168 963
rect 1308 959 1312 963
rect 1452 959 1456 963
rect 1588 959 1592 963
rect 1732 959 1736 963
rect 3592 1003 3596 1007
rect 2492 975 2496 979
rect 2588 975 2592 979
rect 2684 975 2688 979
rect 2924 975 2928 979
rect 3220 975 3224 979
rect 3380 975 3384 979
rect 3540 975 3544 979
rect 3592 975 3596 979
rect 3876 975 3880 979
rect 2796 971 2800 975
rect 3068 971 3072 975
rect 3708 971 3712 975
rect 2448 955 2452 959
rect 2460 955 2464 959
rect 2556 955 2560 959
rect 2652 955 2656 959
rect 2748 955 2752 959
rect 2860 955 2864 959
rect 2988 955 2992 959
rect 3140 955 3144 959
rect 3224 955 3228 959
rect 3308 955 3312 959
rect 3400 955 3404 959
rect 3492 955 3496 959
rect 3684 955 3688 959
rect 3876 955 3880 959
rect 3224 927 3228 931
rect 3400 927 3404 931
rect 944 847 948 851
rect 2336 847 2340 851
rect 484 819 488 823
rect 676 819 680 823
rect 860 819 864 823
rect 944 819 948 823
rect 1036 819 1040 823
rect 1364 819 1368 823
rect 1516 819 1520 823
rect 1668 819 1672 823
rect 1820 819 1824 823
rect 292 815 296 819
rect 1204 815 1208 819
rect 2380 819 2384 823
rect 2476 819 2480 823
rect 2572 819 2576 823
rect 2668 819 2672 823
rect 2772 819 2776 823
rect 2900 819 2904 823
rect 3052 819 3056 823
rect 3228 819 3232 823
rect 3428 819 3432 823
rect 3644 819 3648 823
rect 3860 819 3864 823
rect 2336 803 2340 807
rect 2348 803 2352 807
rect 2532 803 2536 807
rect 2724 803 2728 807
rect 2916 805 2920 809
rect 3116 803 3120 807
rect 3324 803 3328 807
rect 3540 803 3544 807
rect 3756 803 3760 807
rect 196 799 200 803
rect 256 799 260 803
rect 348 799 352 803
rect 508 799 512 803
rect 660 799 664 803
rect 812 799 816 803
rect 972 799 976 803
rect 1132 799 1136 803
rect 1292 799 1296 803
rect 1452 799 1456 803
rect 1620 799 1624 803
rect 1788 799 1792 803
rect 1940 799 1944 803
rect 256 771 260 775
rect 2680 775 2684 779
rect 1104 691 1108 695
rect 2200 691 2204 695
rect 300 663 304 667
rect 468 663 472 667
rect 660 663 664 667
rect 860 663 864 667
rect 1052 663 1056 667
rect 1104 663 1108 667
rect 1428 663 1432 667
rect 1604 663 1608 667
rect 1780 663 1784 667
rect 1940 663 1944 667
rect 2108 663 2112 667
rect 2200 663 2204 667
rect 2292 663 2296 667
rect 2680 663 2684 667
rect 2692 663 2696 667
rect 2892 663 2896 667
rect 3084 663 3088 667
rect 3276 663 3280 667
rect 3476 663 3480 667
rect 3676 663 3680 667
rect 3876 663 3880 667
rect 172 659 176 663
rect 1244 659 1248 663
rect 1392 659 1396 663
rect 2492 659 2496 663
rect 172 647 176 651
rect 284 647 288 651
rect 420 647 424 651
rect 564 647 568 651
rect 724 647 728 651
rect 908 647 912 651
rect 1116 647 1120 651
rect 1340 647 1344 651
rect 1580 647 1584 651
rect 1820 647 1824 651
rect 2108 647 2112 651
rect 2268 647 2272 651
rect 2468 647 2472 651
rect 2668 647 2672 651
rect 2868 647 2872 651
rect 3060 649 3064 653
rect 3244 647 3248 651
rect 3412 647 3416 651
rect 3572 647 3576 651
rect 3732 647 3736 651
rect 3876 647 3880 651
rect 1392 619 1396 623
rect 472 535 476 539
rect 332 507 336 511
rect 172 503 176 507
rect 576 535 580 539
rect 1520 535 1524 539
rect 2184 535 2188 539
rect 2696 535 2700 539
rect 3448 535 3452 539
rect 3584 535 3588 539
rect 516 507 520 511
rect 576 507 580 511
rect 700 507 704 511
rect 884 507 888 511
rect 1252 507 1256 511
rect 1436 507 1440 511
rect 1520 507 1524 511
rect 1628 507 1632 511
rect 1820 507 1824 511
rect 2108 507 2112 511
rect 2184 507 2188 511
rect 2252 507 2256 511
rect 2436 507 2440 511
rect 2620 507 2624 511
rect 2696 507 2700 511
rect 2996 507 3000 511
rect 3180 507 3184 511
rect 3356 507 3360 511
rect 3448 507 3452 511
rect 3532 507 3536 511
rect 3584 507 3588 511
rect 3716 507 3720 511
rect 3876 507 3880 511
rect 1068 503 1072 507
rect 2812 503 2816 507
rect 172 491 176 495
rect 324 491 328 495
rect 472 491 476 495
rect 492 491 496 495
rect 652 491 656 495
rect 804 491 808 495
rect 940 491 944 495
rect 1068 489 1072 493
rect 1196 491 1200 495
rect 1324 491 1328 495
rect 1452 491 1456 495
rect 2108 487 2112 491
rect 2260 487 2264 491
rect 2428 487 2432 491
rect 2596 487 2600 491
rect 2764 487 2768 491
rect 2932 487 2936 491
rect 3100 487 3104 491
rect 3260 487 3264 491
rect 3420 487 3424 491
rect 3580 485 3584 489
rect 3740 487 3744 491
rect 3876 487 3880 491
rect 1032 383 1036 387
rect 324 355 328 359
rect 484 355 488 359
rect 636 355 640 359
rect 788 355 792 359
rect 940 355 944 359
rect 1032 355 1036 359
rect 1116 355 1120 359
rect 1516 355 1520 359
rect 1740 355 1744 359
rect 1940 355 1944 359
rect 152 351 156 355
rect 172 351 176 355
rect 1308 351 1312 355
rect 2500 351 2504 355
rect 2596 351 2600 355
rect 2692 351 2696 355
rect 2884 351 2888 355
rect 2980 351 2984 355
rect 3076 351 3080 355
rect 3172 351 3176 355
rect 3268 351 3272 355
rect 2788 347 2792 351
rect 196 335 200 339
rect 376 335 380 339
rect 388 335 392 339
rect 588 335 592 339
rect 796 335 800 339
rect 996 335 1000 339
rect 1196 337 1200 341
rect 152 307 156 311
rect 1380 333 1384 337
rect 1564 335 1568 339
rect 1748 335 1752 339
rect 1932 335 1936 339
rect 2436 335 2440 339
rect 2540 335 2544 339
rect 2660 335 2664 339
rect 2796 335 2800 339
rect 2948 335 2952 339
rect 3108 335 3112 339
rect 3284 335 3288 339
rect 3460 335 3464 339
rect 3644 333 3648 337
rect 3828 335 3832 339
rect 376 219 380 223
rect 640 219 644 223
rect 1296 219 1300 223
rect 1472 219 1476 223
rect 2388 199 2392 203
rect 2556 199 2560 203
rect 2724 199 2728 203
rect 2892 199 2896 203
rect 3068 199 3072 203
rect 3252 199 3256 203
rect 3444 199 3448 203
rect 3844 199 3848 203
rect 2228 195 2232 199
rect 3632 195 3636 199
rect 3644 195 3648 199
rect 420 191 424 195
rect 580 191 584 195
rect 640 191 644 195
rect 740 191 744 195
rect 900 191 904 195
rect 1068 191 1072 195
rect 1236 191 1240 195
rect 1296 191 1300 195
rect 1404 191 1408 195
rect 1472 191 1476 195
rect 1580 191 1584 195
rect 1764 191 1768 195
rect 260 187 264 191
rect 1940 187 1944 191
rect 172 153 176 157
rect 268 155 272 159
rect 364 155 368 159
rect 460 155 464 159
rect 564 153 568 157
rect 684 155 688 159
rect 812 155 816 159
rect 940 155 944 159
rect 1068 155 1072 159
rect 1188 155 1192 159
rect 1308 155 1312 159
rect 1420 155 1424 159
rect 1524 155 1528 159
rect 1628 155 1632 159
rect 1740 155 1744 159
rect 1844 155 1848 159
rect 1940 155 1944 159
rect 2108 151 2112 155
rect 2204 151 2208 155
rect 2300 151 2304 155
rect 2404 151 2408 155
rect 2524 151 2528 155
rect 2652 151 2656 155
rect 2780 151 2784 155
rect 2908 153 2912 157
rect 3028 151 3032 155
rect 3148 151 3152 155
rect 3260 151 3264 155
rect 3364 151 3368 155
rect 3416 151 3420 155
rect 3468 151 3472 155
rect 3572 151 3576 155
rect 3624 151 3628 155
rect 3416 123 3420 127
rect 3624 123 3628 127
rect 3676 151 3680 155
rect 3780 151 3784 155
rect 3876 151 3880 155
rect 3632 123 3636 127
<< m2 >>
rect 1978 4023 1984 4024
rect 1978 4019 1979 4023
rect 1983 4022 1984 4023
rect 2107 4023 2113 4024
rect 2107 4022 2108 4023
rect 1983 4020 2108 4022
rect 1983 4019 1984 4020
rect 1978 4018 1984 4019
rect 2107 4019 2108 4020
rect 2112 4019 2113 4023
rect 2107 4018 2113 4019
rect 2046 4004 2052 4005
rect 3942 4004 3948 4005
rect 226 4003 232 4004
rect 226 3999 227 4003
rect 231 4002 232 4003
rect 315 4003 321 4004
rect 315 4002 316 4003
rect 231 4000 316 4002
rect 231 3999 232 4000
rect 226 3998 232 3999
rect 315 3999 316 4000
rect 320 3999 321 4003
rect 315 3998 321 3999
rect 354 4003 360 4004
rect 354 3999 355 4003
rect 359 4002 360 4003
rect 467 4003 473 4004
rect 467 4002 468 4003
rect 359 4000 468 4002
rect 359 3999 360 4000
rect 354 3998 360 3999
rect 467 3999 468 4000
rect 472 3999 473 4003
rect 467 3998 473 3999
rect 506 4003 512 4004
rect 506 3999 507 4003
rect 511 4002 512 4003
rect 643 4003 649 4004
rect 643 4002 644 4003
rect 511 4000 644 4002
rect 511 3999 512 4000
rect 506 3998 512 3999
rect 643 3999 644 4000
rect 648 3999 649 4003
rect 643 3998 649 3999
rect 682 4003 688 4004
rect 682 3999 683 4003
rect 687 4002 688 4003
rect 827 4003 833 4004
rect 827 4002 828 4003
rect 687 4000 828 4002
rect 687 3999 688 4000
rect 682 3998 688 3999
rect 827 3999 828 4000
rect 832 3999 833 4003
rect 827 3998 833 3999
rect 866 4003 872 4004
rect 866 3999 867 4003
rect 871 4002 872 4003
rect 1011 4003 1017 4004
rect 1011 4002 1012 4003
rect 871 4000 1012 4002
rect 871 3999 872 4000
rect 866 3998 872 3999
rect 1011 3999 1012 4000
rect 1016 3999 1017 4003
rect 1226 4003 1232 4004
rect 1011 3998 1017 3999
rect 1187 4001 1193 4002
rect 1187 3997 1188 4001
rect 1192 3997 1193 4001
rect 1226 3999 1227 4003
rect 1231 4002 1232 4003
rect 1347 4003 1353 4004
rect 1347 4002 1348 4003
rect 1231 4000 1348 4002
rect 1231 3999 1232 4000
rect 1226 3998 1232 3999
rect 1347 3999 1348 4000
rect 1352 3999 1353 4003
rect 1347 3998 1353 3999
rect 1386 4003 1392 4004
rect 1386 3999 1387 4003
rect 1391 4002 1392 4003
rect 1507 4003 1513 4004
rect 1507 4002 1508 4003
rect 1391 4000 1508 4002
rect 1391 3999 1392 4000
rect 1386 3998 1392 3999
rect 1507 3999 1508 4000
rect 1512 3999 1513 4003
rect 1507 3998 1513 3999
rect 1546 4003 1552 4004
rect 1546 3999 1547 4003
rect 1551 4002 1552 4003
rect 1659 4003 1665 4004
rect 1659 4002 1660 4003
rect 1551 4000 1660 4002
rect 1551 3999 1552 4000
rect 1546 3998 1552 3999
rect 1659 3999 1660 4000
rect 1664 3999 1665 4003
rect 1659 3998 1665 3999
rect 1698 4003 1704 4004
rect 1698 3999 1699 4003
rect 1703 4002 1704 4003
rect 1811 4003 1817 4004
rect 1811 4002 1812 4003
rect 1703 4000 1812 4002
rect 1703 3999 1704 4000
rect 1698 3998 1704 3999
rect 1811 3999 1812 4000
rect 1816 3999 1817 4003
rect 1811 3998 1817 3999
rect 1850 4003 1856 4004
rect 1850 3999 1851 4003
rect 1855 4002 1856 4003
rect 1939 4003 1945 4004
rect 1939 4002 1940 4003
rect 1855 4000 1940 4002
rect 1855 3999 1856 4000
rect 1850 3998 1856 3999
rect 1939 3999 1940 4000
rect 1944 3999 1945 4003
rect 2046 4000 2047 4004
rect 2051 4000 2052 4004
rect 2046 3999 2052 4000
rect 2070 4003 2076 4004
rect 2070 3999 2071 4003
rect 2075 3999 2076 4003
rect 3942 4000 3943 4004
rect 3947 4000 3948 4004
rect 3942 3999 3948 4000
rect 1939 3998 1945 3999
rect 2070 3998 2076 3999
rect 1187 3996 1193 3997
rect 1188 3994 1190 3996
rect 1410 3995 1416 3996
rect 1410 3994 1411 3995
rect 1188 3992 1411 3994
rect 1410 3991 1411 3992
rect 1415 3991 1416 3995
rect 1410 3990 1416 3991
rect 2146 3991 2152 3992
rect 2046 3987 2052 3988
rect 110 3984 116 3985
rect 2006 3984 2012 3985
rect 110 3980 111 3984
rect 115 3980 116 3984
rect 110 3979 116 3980
rect 150 3983 156 3984
rect 150 3979 151 3983
rect 155 3979 156 3983
rect 150 3978 156 3979
rect 278 3983 284 3984
rect 278 3979 279 3983
rect 283 3979 284 3983
rect 278 3978 284 3979
rect 430 3983 436 3984
rect 430 3979 431 3983
rect 435 3979 436 3983
rect 430 3978 436 3979
rect 606 3983 612 3984
rect 606 3979 607 3983
rect 611 3979 612 3983
rect 606 3978 612 3979
rect 790 3983 796 3984
rect 790 3979 791 3983
rect 795 3979 796 3983
rect 790 3978 796 3979
rect 974 3983 980 3984
rect 974 3979 975 3983
rect 979 3979 980 3983
rect 974 3978 980 3979
rect 1150 3983 1156 3984
rect 1150 3979 1151 3983
rect 1155 3979 1156 3983
rect 1150 3978 1156 3979
rect 1310 3983 1316 3984
rect 1310 3979 1311 3983
rect 1315 3979 1316 3983
rect 1310 3978 1316 3979
rect 1470 3983 1476 3984
rect 1470 3979 1471 3983
rect 1475 3979 1476 3983
rect 1470 3978 1476 3979
rect 1622 3983 1628 3984
rect 1622 3979 1623 3983
rect 1627 3979 1628 3983
rect 1622 3978 1628 3979
rect 1774 3983 1780 3984
rect 1774 3979 1775 3983
rect 1779 3979 1780 3983
rect 1774 3978 1780 3979
rect 1902 3983 1908 3984
rect 1902 3979 1903 3983
rect 1907 3979 1908 3983
rect 2006 3980 2007 3984
rect 2011 3980 2012 3984
rect 2046 3983 2047 3987
rect 2051 3983 2052 3987
rect 2146 3987 2147 3991
rect 2151 3987 2152 3991
rect 2146 3986 2152 3987
rect 3942 3987 3948 3988
rect 2046 3982 2052 3983
rect 2070 3984 2076 3985
rect 2006 3979 2012 3980
rect 2070 3980 2071 3984
rect 2075 3980 2076 3984
rect 3942 3983 3943 3987
rect 3947 3983 3948 3987
rect 3942 3982 3948 3983
rect 2070 3979 2076 3980
rect 1902 3978 1908 3979
rect 226 3975 232 3976
rect 226 3971 227 3975
rect 231 3971 232 3975
rect 226 3970 232 3971
rect 354 3975 360 3976
rect 354 3971 355 3975
rect 359 3971 360 3975
rect 354 3970 360 3971
rect 506 3975 512 3976
rect 506 3971 507 3975
rect 511 3971 512 3975
rect 506 3970 512 3971
rect 682 3975 688 3976
rect 682 3971 683 3975
rect 687 3971 688 3975
rect 682 3970 688 3971
rect 866 3975 872 3976
rect 866 3971 867 3975
rect 871 3971 872 3975
rect 866 3970 872 3971
rect 918 3975 924 3976
rect 918 3971 919 3975
rect 923 3974 924 3975
rect 1226 3975 1232 3976
rect 923 3972 1017 3974
rect 923 3971 924 3972
rect 918 3970 924 3971
rect 1226 3971 1227 3975
rect 1231 3971 1232 3975
rect 1226 3970 1232 3971
rect 1386 3975 1392 3976
rect 1386 3971 1387 3975
rect 1391 3971 1392 3975
rect 1386 3970 1392 3971
rect 1546 3975 1552 3976
rect 1546 3971 1547 3975
rect 1551 3971 1552 3975
rect 1546 3970 1552 3971
rect 1698 3975 1704 3976
rect 1698 3971 1699 3975
rect 1703 3971 1704 3975
rect 1698 3970 1704 3971
rect 1850 3975 1856 3976
rect 1850 3971 1851 3975
rect 1855 3971 1856 3975
rect 1850 3970 1856 3971
rect 1978 3975 1984 3976
rect 1978 3971 1979 3975
rect 1983 3971 1984 3975
rect 1978 3970 1984 3971
rect 110 3967 116 3968
rect 110 3963 111 3967
rect 115 3963 116 3967
rect 2006 3967 2012 3968
rect 110 3962 116 3963
rect 150 3964 156 3965
rect 150 3960 151 3964
rect 155 3960 156 3964
rect 150 3959 156 3960
rect 278 3964 284 3965
rect 278 3960 279 3964
rect 283 3960 284 3964
rect 278 3959 284 3960
rect 430 3964 436 3965
rect 430 3960 431 3964
rect 435 3960 436 3964
rect 430 3959 436 3960
rect 606 3964 612 3965
rect 606 3960 607 3964
rect 611 3960 612 3964
rect 606 3959 612 3960
rect 790 3964 796 3965
rect 790 3960 791 3964
rect 795 3960 796 3964
rect 790 3959 796 3960
rect 974 3964 980 3965
rect 974 3960 975 3964
rect 979 3960 980 3964
rect 974 3959 980 3960
rect 1150 3964 1156 3965
rect 1150 3960 1151 3964
rect 1155 3960 1156 3964
rect 1150 3959 1156 3960
rect 1310 3964 1316 3965
rect 1310 3960 1311 3964
rect 1315 3960 1316 3964
rect 1310 3959 1316 3960
rect 1470 3964 1476 3965
rect 1470 3960 1471 3964
rect 1475 3960 1476 3964
rect 1470 3959 1476 3960
rect 1622 3964 1628 3965
rect 1622 3960 1623 3964
rect 1627 3960 1628 3964
rect 1622 3959 1628 3960
rect 1774 3964 1780 3965
rect 1774 3960 1775 3964
rect 1779 3960 1780 3964
rect 1774 3959 1780 3960
rect 1902 3964 1908 3965
rect 1902 3960 1903 3964
rect 1907 3960 1908 3964
rect 2006 3963 2007 3967
rect 2011 3963 2012 3967
rect 2006 3962 2012 3963
rect 1902 3959 1908 3960
rect 2078 3924 2084 3925
rect 2046 3921 2052 3922
rect 2046 3917 2047 3921
rect 2051 3917 2052 3921
rect 2078 3920 2079 3924
rect 2083 3920 2084 3924
rect 2078 3919 2084 3920
rect 2214 3924 2220 3925
rect 2214 3920 2215 3924
rect 2219 3920 2220 3924
rect 2214 3919 2220 3920
rect 2358 3924 2364 3925
rect 2358 3920 2359 3924
rect 2363 3920 2364 3924
rect 2358 3919 2364 3920
rect 2502 3924 2508 3925
rect 2502 3920 2503 3924
rect 2507 3920 2508 3924
rect 2502 3919 2508 3920
rect 2646 3924 2652 3925
rect 2646 3920 2647 3924
rect 2651 3920 2652 3924
rect 2646 3919 2652 3920
rect 2790 3924 2796 3925
rect 2790 3920 2791 3924
rect 2795 3920 2796 3924
rect 2790 3919 2796 3920
rect 2926 3924 2932 3925
rect 2926 3920 2927 3924
rect 2931 3920 2932 3924
rect 2926 3919 2932 3920
rect 3054 3924 3060 3925
rect 3054 3920 3055 3924
rect 3059 3920 3060 3924
rect 3054 3919 3060 3920
rect 3174 3924 3180 3925
rect 3174 3920 3175 3924
rect 3179 3920 3180 3924
rect 3174 3919 3180 3920
rect 3294 3924 3300 3925
rect 3294 3920 3295 3924
rect 3299 3920 3300 3924
rect 3294 3919 3300 3920
rect 3414 3924 3420 3925
rect 3414 3920 3415 3924
rect 3419 3920 3420 3924
rect 3414 3919 3420 3920
rect 3534 3924 3540 3925
rect 3534 3920 3535 3924
rect 3539 3920 3540 3924
rect 3534 3919 3540 3920
rect 3942 3921 3948 3922
rect 2046 3916 2052 3917
rect 3942 3917 3943 3921
rect 3947 3917 3948 3921
rect 3942 3916 3948 3917
rect 2154 3915 2160 3916
rect 2154 3911 2155 3915
rect 2159 3911 2160 3915
rect 2154 3910 2160 3911
rect 2290 3915 2296 3916
rect 2290 3911 2291 3915
rect 2295 3911 2296 3915
rect 2290 3910 2296 3911
rect 2434 3915 2440 3916
rect 2434 3911 2435 3915
rect 2439 3911 2440 3915
rect 2434 3910 2440 3911
rect 2578 3915 2584 3916
rect 2578 3911 2579 3915
rect 2583 3911 2584 3915
rect 2578 3910 2584 3911
rect 2714 3915 2720 3916
rect 2714 3911 2715 3915
rect 2719 3911 2720 3915
rect 2714 3910 2720 3911
rect 2866 3915 2872 3916
rect 2866 3911 2867 3915
rect 2871 3911 2872 3915
rect 2866 3910 2872 3911
rect 3002 3915 3008 3916
rect 3002 3911 3003 3915
rect 3007 3911 3008 3915
rect 3002 3910 3008 3911
rect 3130 3915 3136 3916
rect 3130 3911 3131 3915
rect 3135 3911 3136 3915
rect 3130 3910 3136 3911
rect 3250 3915 3256 3916
rect 3250 3911 3251 3915
rect 3255 3911 3256 3915
rect 3250 3910 3256 3911
rect 3370 3915 3376 3916
rect 3370 3911 3371 3915
rect 3375 3911 3376 3915
rect 3370 3910 3376 3911
rect 3490 3915 3496 3916
rect 3490 3911 3491 3915
rect 3495 3911 3496 3915
rect 3490 3910 3496 3911
rect 3610 3915 3616 3916
rect 3610 3911 3611 3915
rect 3615 3911 3616 3915
rect 3610 3910 3616 3911
rect 2078 3905 2084 3906
rect 302 3904 308 3905
rect 110 3901 116 3902
rect 110 3897 111 3901
rect 115 3897 116 3901
rect 302 3900 303 3904
rect 307 3900 308 3904
rect 302 3899 308 3900
rect 422 3904 428 3905
rect 422 3900 423 3904
rect 427 3900 428 3904
rect 422 3899 428 3900
rect 550 3904 556 3905
rect 550 3900 551 3904
rect 555 3900 556 3904
rect 550 3899 556 3900
rect 686 3904 692 3905
rect 686 3900 687 3904
rect 691 3900 692 3904
rect 686 3899 692 3900
rect 814 3904 820 3905
rect 814 3900 815 3904
rect 819 3900 820 3904
rect 814 3899 820 3900
rect 942 3904 948 3905
rect 942 3900 943 3904
rect 947 3900 948 3904
rect 942 3899 948 3900
rect 1070 3904 1076 3905
rect 1070 3900 1071 3904
rect 1075 3900 1076 3904
rect 1070 3899 1076 3900
rect 1198 3904 1204 3905
rect 1198 3900 1199 3904
rect 1203 3900 1204 3904
rect 1198 3899 1204 3900
rect 1326 3904 1332 3905
rect 1326 3900 1327 3904
rect 1331 3900 1332 3904
rect 1326 3899 1332 3900
rect 1462 3904 1468 3905
rect 1462 3900 1463 3904
rect 1467 3900 1468 3904
rect 2046 3904 2052 3905
rect 1462 3899 1468 3900
rect 2006 3901 2012 3902
rect 110 3896 116 3897
rect 2006 3897 2007 3901
rect 2011 3897 2012 3901
rect 2046 3900 2047 3904
rect 2051 3900 2052 3904
rect 2078 3901 2079 3905
rect 2083 3901 2084 3905
rect 2078 3900 2084 3901
rect 2214 3905 2220 3906
rect 2214 3901 2215 3905
rect 2219 3901 2220 3905
rect 2214 3900 2220 3901
rect 2358 3905 2364 3906
rect 2358 3901 2359 3905
rect 2363 3901 2364 3905
rect 2358 3900 2364 3901
rect 2502 3905 2508 3906
rect 2502 3901 2503 3905
rect 2507 3901 2508 3905
rect 2502 3900 2508 3901
rect 2646 3905 2652 3906
rect 2646 3901 2647 3905
rect 2651 3901 2652 3905
rect 2646 3900 2652 3901
rect 2790 3905 2796 3906
rect 2790 3901 2791 3905
rect 2795 3901 2796 3905
rect 2790 3900 2796 3901
rect 2926 3905 2932 3906
rect 2926 3901 2927 3905
rect 2931 3901 2932 3905
rect 2926 3900 2932 3901
rect 3054 3905 3060 3906
rect 3054 3901 3055 3905
rect 3059 3901 3060 3905
rect 3054 3900 3060 3901
rect 3174 3905 3180 3906
rect 3174 3901 3175 3905
rect 3179 3901 3180 3905
rect 3174 3900 3180 3901
rect 3294 3905 3300 3906
rect 3294 3901 3295 3905
rect 3299 3901 3300 3905
rect 3294 3900 3300 3901
rect 3414 3905 3420 3906
rect 3414 3901 3415 3905
rect 3419 3901 3420 3905
rect 3414 3900 3420 3901
rect 3534 3905 3540 3906
rect 3534 3901 3535 3905
rect 3539 3901 3540 3905
rect 3534 3900 3540 3901
rect 3942 3904 3948 3905
rect 3942 3900 3943 3904
rect 3947 3900 3948 3904
rect 2046 3899 2052 3900
rect 3942 3899 3948 3900
rect 2006 3896 2012 3897
rect 378 3895 384 3896
rect 378 3891 379 3895
rect 383 3891 384 3895
rect 378 3890 384 3891
rect 498 3895 504 3896
rect 498 3891 499 3895
rect 503 3891 504 3895
rect 498 3890 504 3891
rect 626 3895 632 3896
rect 626 3891 627 3895
rect 631 3891 632 3895
rect 626 3890 632 3891
rect 762 3895 768 3896
rect 762 3891 763 3895
rect 767 3891 768 3895
rect 762 3890 768 3891
rect 770 3895 776 3896
rect 770 3891 771 3895
rect 775 3894 776 3895
rect 1018 3895 1024 3896
rect 775 3892 857 3894
rect 775 3891 776 3892
rect 770 3890 776 3891
rect 1018 3891 1019 3895
rect 1023 3891 1024 3895
rect 1018 3890 1024 3891
rect 1146 3895 1152 3896
rect 1146 3891 1147 3895
rect 1151 3891 1152 3895
rect 1146 3890 1152 3891
rect 1274 3895 1280 3896
rect 1274 3891 1275 3895
rect 1279 3891 1280 3895
rect 1274 3890 1280 3891
rect 1402 3895 1408 3896
rect 1402 3891 1403 3895
rect 1407 3891 1408 3895
rect 1402 3890 1408 3891
rect 1410 3895 1416 3896
rect 1410 3891 1411 3895
rect 1415 3894 1416 3895
rect 1415 3892 1505 3894
rect 1415 3891 1416 3892
rect 1410 3890 1416 3891
rect 2115 3887 2121 3888
rect 302 3885 308 3886
rect 110 3884 116 3885
rect 110 3880 111 3884
rect 115 3880 116 3884
rect 302 3881 303 3885
rect 307 3881 308 3885
rect 302 3880 308 3881
rect 422 3885 428 3886
rect 422 3881 423 3885
rect 427 3881 428 3885
rect 422 3880 428 3881
rect 550 3885 556 3886
rect 550 3881 551 3885
rect 555 3881 556 3885
rect 550 3880 556 3881
rect 686 3885 692 3886
rect 686 3881 687 3885
rect 691 3881 692 3885
rect 686 3880 692 3881
rect 814 3885 820 3886
rect 814 3881 815 3885
rect 819 3881 820 3885
rect 814 3880 820 3881
rect 942 3885 948 3886
rect 942 3881 943 3885
rect 947 3881 948 3885
rect 942 3880 948 3881
rect 1070 3885 1076 3886
rect 1070 3881 1071 3885
rect 1075 3881 1076 3885
rect 1070 3880 1076 3881
rect 1198 3885 1204 3886
rect 1198 3881 1199 3885
rect 1203 3881 1204 3885
rect 1198 3880 1204 3881
rect 1326 3885 1332 3886
rect 1326 3881 1327 3885
rect 1331 3881 1332 3885
rect 1326 3880 1332 3881
rect 1462 3885 1468 3886
rect 1462 3881 1463 3885
rect 1467 3881 1468 3885
rect 1462 3880 1468 3881
rect 2006 3884 2012 3885
rect 2006 3880 2007 3884
rect 2011 3880 2012 3884
rect 2115 3883 2116 3887
rect 2120 3886 2121 3887
rect 2146 3887 2152 3888
rect 2146 3886 2147 3887
rect 2120 3884 2147 3886
rect 2120 3883 2121 3884
rect 2115 3882 2121 3883
rect 2146 3883 2147 3884
rect 2151 3883 2152 3887
rect 2146 3882 2152 3883
rect 2154 3887 2160 3888
rect 2154 3883 2155 3887
rect 2159 3886 2160 3887
rect 2251 3887 2257 3888
rect 2251 3886 2252 3887
rect 2159 3884 2252 3886
rect 2159 3883 2160 3884
rect 2154 3882 2160 3883
rect 2251 3883 2252 3884
rect 2256 3883 2257 3887
rect 2251 3882 2257 3883
rect 2290 3887 2296 3888
rect 2290 3883 2291 3887
rect 2295 3886 2296 3887
rect 2395 3887 2401 3888
rect 2395 3886 2396 3887
rect 2295 3884 2396 3886
rect 2295 3883 2296 3884
rect 2290 3882 2296 3883
rect 2395 3883 2396 3884
rect 2400 3883 2401 3887
rect 2395 3882 2401 3883
rect 2434 3887 2440 3888
rect 2434 3883 2435 3887
rect 2439 3886 2440 3887
rect 2539 3887 2545 3888
rect 2539 3886 2540 3887
rect 2439 3884 2540 3886
rect 2439 3883 2440 3884
rect 2434 3882 2440 3883
rect 2539 3883 2540 3884
rect 2544 3883 2545 3887
rect 2539 3882 2545 3883
rect 2578 3887 2584 3888
rect 2578 3883 2579 3887
rect 2583 3886 2584 3887
rect 2683 3887 2689 3888
rect 2683 3886 2684 3887
rect 2583 3884 2684 3886
rect 2583 3883 2584 3884
rect 2578 3882 2584 3883
rect 2683 3883 2684 3884
rect 2688 3883 2689 3887
rect 2866 3887 2872 3888
rect 2683 3882 2689 3883
rect 2827 3883 2833 3884
rect 110 3879 116 3880
rect 2006 3879 2012 3880
rect 2827 3879 2828 3883
rect 2832 3882 2833 3883
rect 2866 3883 2867 3887
rect 2871 3886 2872 3887
rect 2963 3887 2969 3888
rect 2963 3886 2964 3887
rect 2871 3884 2964 3886
rect 2871 3883 2872 3884
rect 2866 3882 2872 3883
rect 2963 3883 2964 3884
rect 2968 3883 2969 3887
rect 2963 3882 2969 3883
rect 3002 3887 3008 3888
rect 3002 3883 3003 3887
rect 3007 3886 3008 3887
rect 3091 3887 3097 3888
rect 3091 3886 3092 3887
rect 3007 3884 3092 3886
rect 3007 3883 3008 3884
rect 3002 3882 3008 3883
rect 3091 3883 3092 3884
rect 3096 3883 3097 3887
rect 3091 3882 3097 3883
rect 3130 3887 3136 3888
rect 3130 3883 3131 3887
rect 3135 3886 3136 3887
rect 3211 3887 3217 3888
rect 3211 3886 3212 3887
rect 3135 3884 3212 3886
rect 3135 3883 3136 3884
rect 3130 3882 3136 3883
rect 3211 3883 3212 3884
rect 3216 3883 3217 3887
rect 3211 3882 3217 3883
rect 3250 3887 3256 3888
rect 3250 3883 3251 3887
rect 3255 3886 3256 3887
rect 3331 3887 3337 3888
rect 3331 3886 3332 3887
rect 3255 3884 3332 3886
rect 3255 3883 3256 3884
rect 3250 3882 3256 3883
rect 3331 3883 3332 3884
rect 3336 3883 3337 3887
rect 3331 3882 3337 3883
rect 3370 3887 3376 3888
rect 3370 3883 3371 3887
rect 3375 3886 3376 3887
rect 3451 3887 3457 3888
rect 3451 3886 3452 3887
rect 3375 3884 3452 3886
rect 3375 3883 3376 3884
rect 3370 3882 3376 3883
rect 3451 3883 3452 3884
rect 3456 3883 3457 3887
rect 3451 3882 3457 3883
rect 3490 3887 3496 3888
rect 3490 3883 3491 3887
rect 3495 3886 3496 3887
rect 3571 3887 3577 3888
rect 3571 3886 3572 3887
rect 3495 3884 3572 3886
rect 3495 3883 3496 3884
rect 3490 3882 3496 3883
rect 3571 3883 3572 3884
rect 3576 3883 3577 3887
rect 3571 3882 3577 3883
rect 2832 3880 2841 3882
rect 2832 3879 2833 3880
rect 2827 3878 2833 3879
rect 2839 3878 2841 3880
rect 3078 3879 3084 3880
rect 3078 3878 3079 3879
rect 2839 3876 3079 3878
rect 918 3875 924 3876
rect 918 3874 919 3875
rect 372 3872 919 3874
rect 339 3867 345 3868
rect 339 3863 340 3867
rect 344 3866 345 3867
rect 372 3866 374 3872
rect 918 3871 919 3872
rect 923 3871 924 3875
rect 3078 3875 3079 3876
rect 3083 3875 3084 3879
rect 3078 3874 3084 3875
rect 918 3870 924 3871
rect 2330 3871 2336 3872
rect 2291 3869 2297 3870
rect 344 3864 374 3866
rect 378 3867 384 3868
rect 344 3863 345 3864
rect 339 3862 345 3863
rect 378 3863 379 3867
rect 383 3866 384 3867
rect 459 3867 465 3868
rect 459 3866 460 3867
rect 383 3864 460 3866
rect 383 3863 384 3864
rect 378 3862 384 3863
rect 459 3863 460 3864
rect 464 3863 465 3867
rect 459 3862 465 3863
rect 498 3867 504 3868
rect 498 3863 499 3867
rect 503 3866 504 3867
rect 587 3867 593 3868
rect 587 3866 588 3867
rect 503 3864 588 3866
rect 503 3863 504 3864
rect 498 3862 504 3863
rect 587 3863 588 3864
rect 592 3863 593 3867
rect 587 3862 593 3863
rect 626 3867 632 3868
rect 626 3863 627 3867
rect 631 3866 632 3867
rect 723 3867 729 3868
rect 723 3866 724 3867
rect 631 3864 724 3866
rect 631 3863 632 3864
rect 626 3862 632 3863
rect 723 3863 724 3864
rect 728 3863 729 3867
rect 723 3862 729 3863
rect 762 3867 768 3868
rect 762 3863 763 3867
rect 767 3866 768 3867
rect 851 3867 857 3868
rect 851 3866 852 3867
rect 767 3864 852 3866
rect 767 3863 768 3864
rect 762 3862 768 3863
rect 851 3863 852 3864
rect 856 3863 857 3867
rect 1018 3867 1024 3868
rect 851 3862 857 3863
rect 979 3863 988 3864
rect 979 3859 980 3863
rect 987 3859 988 3863
rect 1018 3863 1019 3867
rect 1023 3866 1024 3867
rect 1107 3867 1113 3868
rect 1107 3866 1108 3867
rect 1023 3864 1108 3866
rect 1023 3863 1024 3864
rect 1018 3862 1024 3863
rect 1107 3863 1108 3864
rect 1112 3863 1113 3867
rect 1107 3862 1113 3863
rect 1146 3867 1152 3868
rect 1146 3863 1147 3867
rect 1151 3866 1152 3867
rect 1235 3867 1241 3868
rect 1235 3866 1236 3867
rect 1151 3864 1236 3866
rect 1151 3863 1152 3864
rect 1146 3862 1152 3863
rect 1235 3863 1236 3864
rect 1240 3863 1241 3867
rect 1235 3862 1241 3863
rect 1274 3867 1280 3868
rect 1274 3863 1275 3867
rect 1279 3866 1280 3867
rect 1363 3867 1369 3868
rect 1363 3866 1364 3867
rect 1279 3864 1364 3866
rect 1279 3863 1280 3864
rect 1274 3862 1280 3863
rect 1363 3863 1364 3864
rect 1368 3863 1369 3867
rect 1363 3862 1369 3863
rect 1402 3867 1408 3868
rect 1402 3863 1403 3867
rect 1407 3866 1408 3867
rect 1499 3867 1505 3868
rect 1499 3866 1500 3867
rect 1407 3864 1500 3866
rect 1407 3863 1408 3864
rect 1402 3862 1408 3863
rect 1499 3863 1500 3864
rect 1504 3863 1505 3867
rect 2291 3865 2292 3869
rect 2296 3865 2297 3869
rect 2330 3867 2331 3871
rect 2335 3870 2336 3871
rect 2419 3871 2425 3872
rect 2419 3870 2420 3871
rect 2335 3868 2420 3870
rect 2335 3867 2336 3868
rect 2330 3866 2336 3867
rect 2419 3867 2420 3868
rect 2424 3867 2425 3871
rect 2419 3866 2425 3867
rect 2458 3871 2464 3872
rect 2458 3867 2459 3871
rect 2463 3870 2464 3871
rect 2555 3871 2561 3872
rect 2555 3870 2556 3871
rect 2463 3868 2556 3870
rect 2463 3867 2464 3868
rect 2458 3866 2464 3867
rect 2555 3867 2556 3868
rect 2560 3867 2561 3871
rect 2555 3866 2561 3867
rect 2707 3871 2716 3872
rect 2707 3867 2708 3871
rect 2715 3867 2716 3871
rect 2707 3866 2716 3867
rect 2746 3871 2752 3872
rect 2746 3867 2747 3871
rect 2751 3870 2752 3871
rect 2867 3871 2873 3872
rect 2867 3870 2868 3871
rect 2751 3868 2868 3870
rect 2751 3867 2752 3868
rect 2746 3866 2752 3867
rect 2867 3867 2868 3868
rect 2872 3867 2873 3871
rect 2867 3866 2873 3867
rect 3026 3871 3033 3872
rect 3026 3867 3027 3871
rect 3032 3867 3033 3871
rect 3026 3866 3033 3867
rect 3066 3871 3072 3872
rect 3066 3867 3067 3871
rect 3071 3870 3072 3871
rect 3195 3871 3201 3872
rect 3195 3870 3196 3871
rect 3071 3868 3196 3870
rect 3071 3867 3072 3868
rect 3066 3866 3072 3867
rect 3195 3867 3196 3868
rect 3200 3867 3201 3871
rect 3195 3866 3201 3867
rect 3363 3871 3369 3872
rect 3363 3867 3364 3871
rect 3368 3870 3369 3871
rect 3415 3871 3421 3872
rect 3415 3870 3416 3871
rect 3368 3868 3416 3870
rect 3368 3867 3369 3868
rect 3363 3866 3369 3867
rect 3415 3867 3416 3868
rect 3420 3867 3421 3871
rect 3415 3866 3421 3867
rect 3531 3871 3537 3872
rect 3531 3867 3532 3871
rect 3536 3870 3537 3871
rect 3602 3871 3608 3872
rect 3602 3870 3603 3871
rect 3536 3868 3603 3870
rect 3536 3867 3537 3868
rect 3531 3866 3537 3867
rect 3602 3867 3603 3868
rect 3607 3867 3608 3871
rect 3602 3866 3608 3867
rect 3610 3871 3616 3872
rect 3610 3867 3611 3871
rect 3615 3870 3616 3871
rect 3699 3871 3705 3872
rect 3699 3870 3700 3871
rect 3615 3868 3700 3870
rect 3615 3867 3616 3868
rect 3610 3866 3616 3867
rect 3699 3867 3700 3868
rect 3704 3867 3705 3871
rect 3699 3866 3705 3867
rect 2291 3864 2297 3865
rect 1499 3862 1505 3863
rect 2292 3862 2294 3864
rect 2778 3863 2784 3864
rect 2778 3862 2779 3863
rect 2292 3860 2779 3862
rect 979 3858 988 3859
rect 2778 3859 2779 3860
rect 2783 3859 2784 3863
rect 2778 3858 2784 3859
rect 770 3855 776 3856
rect 770 3854 771 3855
rect 452 3852 771 3854
rect 452 3850 454 3852
rect 770 3851 771 3852
rect 775 3851 776 3855
rect 770 3850 776 3851
rect 2046 3852 2052 3853
rect 3942 3852 3948 3853
rect 451 3849 457 3850
rect 451 3845 452 3849
rect 456 3845 457 3849
rect 2046 3848 2047 3852
rect 2051 3848 2052 3852
rect 451 3844 457 3845
rect 490 3847 496 3848
rect 490 3843 491 3847
rect 495 3846 496 3847
rect 603 3847 609 3848
rect 603 3846 604 3847
rect 495 3844 604 3846
rect 495 3843 496 3844
rect 490 3842 496 3843
rect 603 3843 604 3844
rect 608 3843 609 3847
rect 603 3842 609 3843
rect 642 3847 648 3848
rect 642 3843 643 3847
rect 647 3846 648 3847
rect 763 3847 769 3848
rect 763 3846 764 3847
rect 647 3844 764 3846
rect 647 3843 648 3844
rect 642 3842 648 3843
rect 763 3843 764 3844
rect 768 3843 769 3847
rect 763 3842 769 3843
rect 802 3847 808 3848
rect 802 3843 803 3847
rect 807 3846 808 3847
rect 923 3847 929 3848
rect 923 3846 924 3847
rect 807 3844 924 3846
rect 807 3843 808 3844
rect 802 3842 808 3843
rect 923 3843 924 3844
rect 928 3843 929 3847
rect 923 3842 929 3843
rect 1075 3847 1081 3848
rect 1075 3843 1076 3847
rect 1080 3846 1081 3847
rect 1138 3847 1144 3848
rect 1138 3846 1139 3847
rect 1080 3844 1139 3846
rect 1080 3843 1081 3844
rect 1075 3842 1081 3843
rect 1138 3843 1139 3844
rect 1143 3843 1144 3847
rect 1138 3842 1144 3843
rect 1227 3847 1233 3848
rect 1227 3843 1228 3847
rect 1232 3846 1233 3847
rect 1274 3847 1280 3848
rect 1274 3846 1275 3847
rect 1232 3844 1275 3846
rect 1232 3843 1233 3844
rect 1227 3842 1233 3843
rect 1274 3843 1275 3844
rect 1279 3843 1280 3847
rect 1274 3842 1280 3843
rect 1379 3847 1385 3848
rect 1379 3843 1380 3847
rect 1384 3846 1385 3847
rect 1426 3847 1432 3848
rect 1426 3846 1427 3847
rect 1384 3844 1427 3846
rect 1384 3843 1385 3844
rect 1379 3842 1385 3843
rect 1426 3843 1427 3844
rect 1431 3843 1432 3847
rect 1426 3842 1432 3843
rect 1531 3847 1537 3848
rect 1531 3843 1532 3847
rect 1536 3846 1537 3847
rect 1562 3847 1568 3848
rect 1562 3846 1563 3847
rect 1536 3844 1563 3846
rect 1536 3843 1537 3844
rect 1531 3842 1537 3843
rect 1562 3843 1563 3844
rect 1567 3843 1568 3847
rect 1562 3842 1568 3843
rect 1578 3847 1584 3848
rect 1578 3843 1579 3847
rect 1583 3846 1584 3847
rect 1683 3847 1689 3848
rect 2046 3847 2052 3848
rect 2254 3851 2260 3852
rect 2254 3847 2255 3851
rect 2259 3847 2260 3851
rect 1683 3846 1684 3847
rect 1583 3844 1684 3846
rect 1583 3843 1584 3844
rect 1578 3842 1584 3843
rect 1683 3843 1684 3844
rect 1688 3843 1689 3847
rect 2254 3846 2260 3847
rect 2382 3851 2388 3852
rect 2382 3847 2383 3851
rect 2387 3847 2388 3851
rect 2382 3846 2388 3847
rect 2518 3851 2524 3852
rect 2518 3847 2519 3851
rect 2523 3847 2524 3851
rect 2518 3846 2524 3847
rect 2670 3851 2676 3852
rect 2670 3847 2671 3851
rect 2675 3847 2676 3851
rect 2670 3846 2676 3847
rect 2830 3851 2836 3852
rect 2830 3847 2831 3851
rect 2835 3847 2836 3851
rect 2830 3846 2836 3847
rect 2990 3851 2996 3852
rect 2990 3847 2991 3851
rect 2995 3847 2996 3851
rect 2990 3846 2996 3847
rect 3158 3851 3164 3852
rect 3158 3847 3159 3851
rect 3163 3847 3164 3851
rect 3158 3846 3164 3847
rect 3326 3851 3332 3852
rect 3326 3847 3327 3851
rect 3331 3847 3332 3851
rect 3326 3846 3332 3847
rect 3494 3851 3500 3852
rect 3494 3847 3495 3851
rect 3499 3847 3500 3851
rect 3494 3846 3500 3847
rect 3662 3851 3668 3852
rect 3662 3847 3663 3851
rect 3667 3847 3668 3851
rect 3942 3848 3943 3852
rect 3947 3848 3948 3852
rect 3942 3847 3948 3848
rect 3662 3846 3668 3847
rect 1683 3842 1689 3843
rect 2330 3843 2336 3844
rect 2330 3839 2331 3843
rect 2335 3839 2336 3843
rect 2330 3838 2336 3839
rect 2458 3843 2464 3844
rect 2458 3839 2459 3843
rect 2463 3839 2464 3843
rect 2746 3843 2752 3844
rect 2458 3838 2464 3839
rect 2594 3839 2600 3840
rect 2046 3835 2052 3836
rect 2046 3831 2047 3835
rect 2051 3831 2052 3835
rect 2594 3835 2595 3839
rect 2599 3835 2600 3839
rect 2746 3839 2747 3843
rect 2751 3839 2752 3843
rect 2746 3838 2752 3839
rect 2778 3843 2784 3844
rect 2778 3839 2779 3843
rect 2783 3842 2784 3843
rect 3066 3843 3072 3844
rect 2783 3840 2873 3842
rect 2783 3839 2784 3840
rect 2778 3838 2784 3839
rect 3066 3839 3067 3843
rect 3071 3839 3072 3843
rect 3066 3838 3072 3839
rect 3078 3843 3084 3844
rect 3078 3839 3079 3843
rect 3083 3842 3084 3843
rect 3415 3843 3421 3844
rect 3083 3840 3201 3842
rect 3083 3839 3084 3840
rect 3078 3838 3084 3839
rect 3402 3839 3408 3840
rect 2594 3834 2600 3835
rect 3402 3835 3403 3839
rect 3407 3835 3408 3839
rect 3415 3839 3416 3843
rect 3420 3842 3421 3843
rect 3602 3843 3608 3844
rect 3420 3840 3537 3842
rect 3420 3839 3421 3840
rect 3415 3838 3421 3839
rect 3602 3839 3603 3843
rect 3607 3842 3608 3843
rect 3607 3840 3705 3842
rect 3607 3839 3608 3840
rect 3602 3838 3608 3839
rect 3402 3834 3408 3835
rect 3942 3835 3948 3836
rect 2046 3830 2052 3831
rect 2254 3832 2260 3833
rect 110 3828 116 3829
rect 2006 3828 2012 3829
rect 110 3824 111 3828
rect 115 3824 116 3828
rect 110 3823 116 3824
rect 414 3827 420 3828
rect 414 3823 415 3827
rect 419 3823 420 3827
rect 414 3822 420 3823
rect 566 3827 572 3828
rect 566 3823 567 3827
rect 571 3823 572 3827
rect 566 3822 572 3823
rect 726 3827 732 3828
rect 726 3823 727 3827
rect 731 3823 732 3827
rect 726 3822 732 3823
rect 886 3827 892 3828
rect 886 3823 887 3827
rect 891 3823 892 3827
rect 886 3822 892 3823
rect 1038 3827 1044 3828
rect 1038 3823 1039 3827
rect 1043 3823 1044 3827
rect 1038 3822 1044 3823
rect 1190 3827 1196 3828
rect 1190 3823 1191 3827
rect 1195 3823 1196 3827
rect 1190 3822 1196 3823
rect 1342 3827 1348 3828
rect 1342 3823 1343 3827
rect 1347 3823 1348 3827
rect 1342 3822 1348 3823
rect 1494 3827 1500 3828
rect 1494 3823 1495 3827
rect 1499 3823 1500 3827
rect 1646 3827 1652 3828
rect 1494 3822 1500 3823
rect 1562 3823 1568 3824
rect 490 3819 496 3820
rect 490 3815 491 3819
rect 495 3815 496 3819
rect 490 3814 496 3815
rect 642 3819 648 3820
rect 642 3815 643 3819
rect 647 3815 648 3819
rect 642 3814 648 3815
rect 802 3819 808 3820
rect 802 3815 803 3819
rect 807 3815 808 3819
rect 802 3814 808 3815
rect 858 3819 864 3820
rect 858 3815 859 3819
rect 863 3818 864 3819
rect 982 3819 988 3820
rect 863 3816 929 3818
rect 863 3815 864 3816
rect 858 3814 864 3815
rect 982 3815 983 3819
rect 987 3818 988 3819
rect 1138 3819 1144 3820
rect 987 3816 1081 3818
rect 987 3815 988 3816
rect 982 3814 988 3815
rect 1138 3815 1139 3819
rect 1143 3818 1144 3819
rect 1274 3819 1280 3820
rect 1143 3816 1233 3818
rect 1143 3815 1144 3816
rect 1138 3814 1144 3815
rect 1274 3815 1275 3819
rect 1279 3818 1280 3819
rect 1426 3819 1432 3820
rect 1279 3816 1385 3818
rect 1279 3815 1280 3816
rect 1274 3814 1280 3815
rect 1426 3815 1427 3819
rect 1431 3818 1432 3819
rect 1562 3819 1563 3823
rect 1567 3822 1568 3823
rect 1646 3823 1647 3827
rect 1651 3823 1652 3827
rect 2006 3824 2007 3828
rect 2011 3824 2012 3828
rect 2254 3828 2255 3832
rect 2259 3828 2260 3832
rect 2254 3827 2260 3828
rect 2382 3832 2388 3833
rect 2382 3828 2383 3832
rect 2387 3828 2388 3832
rect 2382 3827 2388 3828
rect 2518 3832 2524 3833
rect 2518 3828 2519 3832
rect 2523 3828 2524 3832
rect 2518 3827 2524 3828
rect 2670 3832 2676 3833
rect 2670 3828 2671 3832
rect 2675 3828 2676 3832
rect 2670 3827 2676 3828
rect 2830 3832 2836 3833
rect 2830 3828 2831 3832
rect 2835 3828 2836 3832
rect 2830 3827 2836 3828
rect 2990 3832 2996 3833
rect 2990 3828 2991 3832
rect 2995 3828 2996 3832
rect 2990 3827 2996 3828
rect 3158 3832 3164 3833
rect 3158 3828 3159 3832
rect 3163 3828 3164 3832
rect 3158 3827 3164 3828
rect 3326 3832 3332 3833
rect 3326 3828 3327 3832
rect 3331 3828 3332 3832
rect 3326 3827 3332 3828
rect 3494 3832 3500 3833
rect 3494 3828 3495 3832
rect 3499 3828 3500 3832
rect 3494 3827 3500 3828
rect 3662 3832 3668 3833
rect 3662 3828 3663 3832
rect 3667 3828 3668 3832
rect 3942 3831 3943 3835
rect 3947 3831 3948 3835
rect 3942 3830 3948 3831
rect 3662 3827 3668 3828
rect 2006 3823 2012 3824
rect 1646 3822 1652 3823
rect 1567 3820 1582 3822
rect 1567 3819 1568 3820
rect 1562 3818 1568 3819
rect 1580 3818 1582 3820
rect 1431 3816 1537 3818
rect 1580 3816 1689 3818
rect 1431 3815 1432 3816
rect 1426 3814 1432 3815
rect 110 3811 116 3812
rect 110 3807 111 3811
rect 115 3807 116 3811
rect 2006 3811 2012 3812
rect 110 3806 116 3807
rect 414 3808 420 3809
rect 414 3804 415 3808
rect 419 3804 420 3808
rect 414 3803 420 3804
rect 566 3808 572 3809
rect 566 3804 567 3808
rect 571 3804 572 3808
rect 566 3803 572 3804
rect 726 3808 732 3809
rect 726 3804 727 3808
rect 731 3804 732 3808
rect 726 3803 732 3804
rect 886 3808 892 3809
rect 886 3804 887 3808
rect 891 3804 892 3808
rect 886 3803 892 3804
rect 1038 3808 1044 3809
rect 1038 3804 1039 3808
rect 1043 3804 1044 3808
rect 1038 3803 1044 3804
rect 1190 3808 1196 3809
rect 1190 3804 1191 3808
rect 1195 3804 1196 3808
rect 1190 3803 1196 3804
rect 1342 3808 1348 3809
rect 1342 3804 1343 3808
rect 1347 3804 1348 3808
rect 1342 3803 1348 3804
rect 1494 3808 1500 3809
rect 1494 3804 1495 3808
rect 1499 3804 1500 3808
rect 1494 3803 1500 3804
rect 1646 3808 1652 3809
rect 1646 3804 1647 3808
rect 1651 3804 1652 3808
rect 2006 3807 2007 3811
rect 2011 3807 2012 3811
rect 2006 3806 2012 3807
rect 1646 3803 1652 3804
rect 2070 3772 2076 3773
rect 2046 3769 2052 3770
rect 2046 3765 2047 3769
rect 2051 3765 2052 3769
rect 2070 3768 2071 3772
rect 2075 3768 2076 3772
rect 2070 3767 2076 3768
rect 2198 3772 2204 3773
rect 2198 3768 2199 3772
rect 2203 3768 2204 3772
rect 2198 3767 2204 3768
rect 2374 3772 2380 3773
rect 2374 3768 2375 3772
rect 2379 3768 2380 3772
rect 2374 3767 2380 3768
rect 2558 3772 2564 3773
rect 2558 3768 2559 3772
rect 2563 3768 2564 3772
rect 2558 3767 2564 3768
rect 2750 3772 2756 3773
rect 2750 3768 2751 3772
rect 2755 3768 2756 3772
rect 2750 3767 2756 3768
rect 2950 3772 2956 3773
rect 2950 3768 2951 3772
rect 2955 3768 2956 3772
rect 2950 3767 2956 3768
rect 3142 3772 3148 3773
rect 3142 3768 3143 3772
rect 3147 3768 3148 3772
rect 3142 3767 3148 3768
rect 3334 3772 3340 3773
rect 3334 3768 3335 3772
rect 3339 3768 3340 3772
rect 3334 3767 3340 3768
rect 3534 3772 3540 3773
rect 3534 3768 3535 3772
rect 3539 3768 3540 3772
rect 3534 3767 3540 3768
rect 3734 3772 3740 3773
rect 3734 3768 3735 3772
rect 3739 3768 3740 3772
rect 3734 3767 3740 3768
rect 3942 3769 3948 3770
rect 2046 3764 2052 3765
rect 3942 3765 3943 3769
rect 3947 3765 3948 3769
rect 3942 3764 3948 3765
rect 2138 3763 2144 3764
rect 2138 3759 2139 3763
rect 2143 3759 2144 3763
rect 2138 3758 2144 3759
rect 2167 3763 2173 3764
rect 2167 3759 2168 3763
rect 2172 3762 2173 3763
rect 2302 3763 2308 3764
rect 2172 3760 2241 3762
rect 2172 3759 2173 3760
rect 2167 3758 2173 3759
rect 2302 3759 2303 3763
rect 2307 3762 2308 3763
rect 2634 3763 2640 3764
rect 2307 3760 2417 3762
rect 2307 3759 2308 3760
rect 2302 3758 2308 3759
rect 2634 3759 2635 3763
rect 2639 3759 2640 3763
rect 2634 3758 2640 3759
rect 2642 3763 2648 3764
rect 2642 3759 2643 3763
rect 2647 3762 2648 3763
rect 3026 3763 3032 3764
rect 2647 3760 2793 3762
rect 2647 3759 2648 3760
rect 2642 3758 2648 3759
rect 3026 3759 3027 3763
rect 3031 3759 3032 3763
rect 3026 3758 3032 3759
rect 3046 3763 3052 3764
rect 3046 3759 3047 3763
rect 3051 3762 3052 3763
rect 3410 3763 3416 3764
rect 3051 3760 3185 3762
rect 3051 3759 3052 3760
rect 3046 3758 3052 3759
rect 3410 3759 3411 3763
rect 3415 3759 3416 3763
rect 3410 3758 3416 3759
rect 3610 3763 3616 3764
rect 3610 3759 3611 3763
rect 3615 3759 3616 3763
rect 3610 3758 3616 3759
rect 3802 3763 3808 3764
rect 3802 3759 3803 3763
rect 3807 3759 3808 3763
rect 3802 3758 3808 3759
rect 438 3755 444 3756
rect 438 3751 439 3755
rect 443 3754 444 3755
rect 858 3755 864 3756
rect 858 3754 859 3755
rect 443 3752 859 3754
rect 443 3751 444 3752
rect 438 3750 444 3751
rect 858 3751 859 3752
rect 863 3751 864 3755
rect 2070 3753 2076 3754
rect 858 3750 864 3751
rect 2046 3752 2052 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2070 3749 2071 3753
rect 2075 3749 2076 3753
rect 2070 3748 2076 3749
rect 2198 3753 2204 3754
rect 2198 3749 2199 3753
rect 2203 3749 2204 3753
rect 2198 3748 2204 3749
rect 2374 3753 2380 3754
rect 2374 3749 2375 3753
rect 2379 3749 2380 3753
rect 2374 3748 2380 3749
rect 2558 3753 2564 3754
rect 2558 3749 2559 3753
rect 2563 3749 2564 3753
rect 2558 3748 2564 3749
rect 2750 3753 2756 3754
rect 2750 3749 2751 3753
rect 2755 3749 2756 3753
rect 2750 3748 2756 3749
rect 2950 3753 2956 3754
rect 2950 3749 2951 3753
rect 2955 3749 2956 3753
rect 2950 3748 2956 3749
rect 3142 3753 3148 3754
rect 3142 3749 3143 3753
rect 3147 3749 3148 3753
rect 3142 3748 3148 3749
rect 3334 3753 3340 3754
rect 3334 3749 3335 3753
rect 3339 3749 3340 3753
rect 3334 3748 3340 3749
rect 3534 3753 3540 3754
rect 3534 3749 3535 3753
rect 3539 3749 3540 3753
rect 3534 3748 3540 3749
rect 3734 3753 3740 3754
rect 3734 3749 3735 3753
rect 3739 3749 3740 3753
rect 3734 3748 3740 3749
rect 3942 3752 3948 3753
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 2046 3747 2052 3748
rect 3942 3747 3948 3748
rect 398 3744 404 3745
rect 110 3741 116 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 398 3740 399 3744
rect 403 3740 404 3744
rect 398 3739 404 3740
rect 566 3744 572 3745
rect 566 3740 567 3744
rect 571 3740 572 3744
rect 566 3739 572 3740
rect 750 3744 756 3745
rect 750 3740 751 3744
rect 755 3740 756 3744
rect 750 3739 756 3740
rect 934 3744 940 3745
rect 934 3740 935 3744
rect 939 3740 940 3744
rect 934 3739 940 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1310 3744 1316 3745
rect 1310 3740 1311 3744
rect 1315 3740 1316 3744
rect 1310 3739 1316 3740
rect 1502 3744 1508 3745
rect 1502 3740 1503 3744
rect 1507 3740 1508 3744
rect 1502 3739 1508 3740
rect 1694 3744 1700 3745
rect 1694 3740 1695 3744
rect 1699 3740 1700 3744
rect 1694 3739 1700 3740
rect 1886 3744 1892 3745
rect 1886 3740 1887 3744
rect 1891 3740 1892 3744
rect 2642 3743 2648 3744
rect 2642 3742 2643 3743
rect 1886 3739 1892 3740
rect 2006 3741 2012 3742
rect 110 3736 116 3737
rect 2006 3737 2007 3741
rect 2011 3737 2012 3741
rect 2006 3736 2012 3737
rect 2588 3740 2643 3742
rect 474 3735 480 3736
rect 474 3731 475 3735
rect 479 3731 480 3735
rect 474 3730 480 3731
rect 642 3735 648 3736
rect 642 3731 643 3735
rect 647 3731 648 3735
rect 642 3730 648 3731
rect 826 3735 832 3736
rect 826 3731 827 3735
rect 831 3731 832 3735
rect 826 3730 832 3731
rect 1010 3735 1016 3736
rect 1010 3731 1011 3735
rect 1015 3731 1016 3735
rect 1010 3730 1016 3731
rect 1103 3735 1109 3736
rect 1103 3731 1104 3735
rect 1108 3734 1109 3735
rect 1386 3735 1392 3736
rect 1108 3732 1169 3734
rect 1108 3731 1109 3732
rect 1103 3730 1109 3731
rect 1386 3731 1387 3735
rect 1391 3731 1392 3735
rect 1386 3730 1392 3731
rect 1578 3735 1584 3736
rect 1578 3731 1579 3735
rect 1583 3731 1584 3735
rect 1578 3730 1584 3731
rect 1586 3735 1592 3736
rect 1586 3731 1587 3735
rect 1591 3734 1592 3735
rect 1798 3735 1804 3736
rect 1591 3732 1737 3734
rect 1591 3731 1592 3732
rect 1586 3730 1592 3731
rect 1798 3731 1799 3735
rect 1803 3734 1804 3735
rect 2107 3735 2113 3736
rect 1803 3732 1929 3734
rect 1803 3731 1804 3732
rect 1798 3730 1804 3731
rect 2107 3731 2108 3735
rect 2112 3734 2113 3735
rect 2167 3735 2173 3736
rect 2167 3734 2168 3735
rect 2112 3732 2168 3734
rect 2112 3731 2113 3732
rect 2107 3730 2113 3731
rect 2167 3731 2168 3732
rect 2172 3731 2173 3735
rect 2167 3730 2173 3731
rect 2235 3735 2241 3736
rect 2235 3731 2236 3735
rect 2240 3734 2241 3735
rect 2302 3735 2308 3736
rect 2302 3734 2303 3735
rect 2240 3732 2303 3734
rect 2240 3731 2241 3732
rect 2235 3730 2241 3731
rect 2302 3731 2303 3732
rect 2307 3731 2308 3735
rect 2302 3730 2308 3731
rect 2411 3735 2417 3736
rect 2411 3731 2412 3735
rect 2416 3734 2417 3735
rect 2588 3734 2590 3740
rect 2642 3739 2643 3740
rect 2647 3739 2648 3743
rect 2642 3738 2648 3739
rect 2416 3732 2590 3734
rect 2594 3735 2601 3736
rect 2416 3731 2417 3732
rect 2411 3730 2417 3731
rect 2594 3731 2595 3735
rect 2600 3731 2601 3735
rect 2594 3730 2601 3731
rect 2634 3735 2640 3736
rect 2634 3731 2635 3735
rect 2639 3734 2640 3735
rect 2787 3735 2793 3736
rect 2787 3734 2788 3735
rect 2639 3732 2788 3734
rect 2639 3731 2640 3732
rect 2634 3730 2640 3731
rect 2787 3731 2788 3732
rect 2792 3731 2793 3735
rect 2787 3730 2793 3731
rect 2987 3735 2993 3736
rect 2987 3731 2988 3735
rect 2992 3734 2993 3735
rect 3046 3735 3052 3736
rect 3046 3734 3047 3735
rect 2992 3732 3047 3734
rect 2992 3731 2993 3732
rect 2987 3730 2993 3731
rect 3046 3731 3047 3732
rect 3051 3731 3052 3735
rect 3371 3735 3377 3736
rect 3046 3730 3052 3731
rect 3179 3731 3185 3732
rect 3179 3727 3180 3731
rect 3184 3730 3185 3731
rect 3194 3731 3200 3732
rect 3194 3730 3195 3731
rect 3184 3728 3195 3730
rect 3184 3727 3185 3728
rect 3179 3726 3185 3727
rect 3194 3727 3195 3728
rect 3199 3727 3200 3731
rect 3371 3731 3372 3735
rect 3376 3734 3377 3735
rect 3402 3735 3408 3736
rect 3402 3734 3403 3735
rect 3376 3732 3403 3734
rect 3376 3731 3377 3732
rect 3371 3730 3377 3731
rect 3402 3731 3403 3732
rect 3407 3731 3408 3735
rect 3402 3730 3408 3731
rect 3410 3735 3416 3736
rect 3410 3731 3411 3735
rect 3415 3734 3416 3735
rect 3571 3735 3577 3736
rect 3571 3734 3572 3735
rect 3415 3732 3572 3734
rect 3415 3731 3416 3732
rect 3410 3730 3416 3731
rect 3571 3731 3572 3732
rect 3576 3731 3577 3735
rect 3571 3730 3577 3731
rect 3610 3735 3616 3736
rect 3610 3731 3611 3735
rect 3615 3734 3616 3735
rect 3771 3735 3777 3736
rect 3771 3734 3772 3735
rect 3615 3732 3772 3734
rect 3615 3731 3616 3732
rect 3610 3730 3616 3731
rect 3771 3731 3772 3732
rect 3776 3731 3777 3735
rect 3771 3730 3777 3731
rect 3194 3726 3200 3727
rect 398 3725 404 3726
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 398 3721 399 3725
rect 403 3721 404 3725
rect 398 3720 404 3721
rect 566 3725 572 3726
rect 566 3721 567 3725
rect 571 3721 572 3725
rect 566 3720 572 3721
rect 750 3725 756 3726
rect 750 3721 751 3725
rect 755 3721 756 3725
rect 750 3720 756 3721
rect 934 3725 940 3726
rect 934 3721 935 3725
rect 939 3721 940 3725
rect 934 3720 940 3721
rect 1126 3725 1132 3726
rect 1126 3721 1127 3725
rect 1131 3721 1132 3725
rect 1126 3720 1132 3721
rect 1310 3725 1316 3726
rect 1310 3721 1311 3725
rect 1315 3721 1316 3725
rect 1310 3720 1316 3721
rect 1502 3725 1508 3726
rect 1502 3721 1503 3725
rect 1507 3721 1508 3725
rect 1502 3720 1508 3721
rect 1694 3725 1700 3726
rect 1694 3721 1695 3725
rect 1699 3721 1700 3725
rect 1694 3720 1700 3721
rect 1886 3725 1892 3726
rect 1886 3721 1887 3725
rect 1891 3721 1892 3725
rect 1886 3720 1892 3721
rect 2006 3724 2012 3725
rect 2006 3720 2007 3724
rect 2011 3720 2012 3724
rect 110 3719 116 3720
rect 2006 3719 2012 3720
rect 1586 3715 1592 3716
rect 1586 3714 1587 3715
rect 1380 3712 1587 3714
rect 435 3707 444 3708
rect 435 3703 436 3707
rect 443 3703 444 3707
rect 435 3702 444 3703
rect 474 3707 480 3708
rect 474 3703 475 3707
rect 479 3706 480 3707
rect 603 3707 609 3708
rect 603 3706 604 3707
rect 479 3704 604 3706
rect 479 3703 480 3704
rect 474 3702 480 3703
rect 603 3703 604 3704
rect 608 3703 609 3707
rect 603 3702 609 3703
rect 642 3707 648 3708
rect 642 3703 643 3707
rect 647 3706 648 3707
rect 787 3707 793 3708
rect 787 3706 788 3707
rect 647 3704 788 3706
rect 647 3703 648 3704
rect 642 3702 648 3703
rect 787 3703 788 3704
rect 792 3703 793 3707
rect 787 3702 793 3703
rect 826 3707 832 3708
rect 826 3703 827 3707
rect 831 3706 832 3707
rect 971 3707 977 3708
rect 971 3706 972 3707
rect 831 3704 972 3706
rect 831 3703 832 3704
rect 826 3702 832 3703
rect 971 3703 972 3704
rect 976 3703 977 3707
rect 971 3702 977 3703
rect 1010 3707 1016 3708
rect 1010 3703 1011 3707
rect 1015 3706 1016 3707
rect 1163 3707 1169 3708
rect 1163 3706 1164 3707
rect 1015 3704 1164 3706
rect 1015 3703 1016 3704
rect 1010 3702 1016 3703
rect 1163 3703 1164 3704
rect 1168 3703 1169 3707
rect 1163 3702 1169 3703
rect 1347 3707 1353 3708
rect 1347 3703 1348 3707
rect 1352 3706 1353 3707
rect 1380 3706 1382 3712
rect 1586 3711 1587 3712
rect 1591 3711 1592 3715
rect 1586 3710 1592 3711
rect 1352 3704 1382 3706
rect 1386 3707 1392 3708
rect 1352 3703 1353 3704
rect 1347 3702 1353 3703
rect 1386 3703 1387 3707
rect 1391 3706 1392 3707
rect 1539 3707 1545 3708
rect 1539 3706 1540 3707
rect 1391 3704 1540 3706
rect 1391 3703 1392 3704
rect 1386 3702 1392 3703
rect 1539 3703 1540 3704
rect 1544 3703 1545 3707
rect 1539 3702 1545 3703
rect 1731 3707 1737 3708
rect 1731 3703 1732 3707
rect 1736 3706 1737 3707
rect 1798 3707 1804 3708
rect 1798 3706 1799 3707
rect 1736 3704 1799 3706
rect 1736 3703 1737 3704
rect 1731 3702 1737 3703
rect 1798 3703 1799 3704
rect 1803 3703 1804 3707
rect 2107 3707 2113 3708
rect 1798 3702 1804 3703
rect 1866 3703 1872 3704
rect 1866 3699 1867 3703
rect 1871 3702 1872 3703
rect 1923 3703 1929 3704
rect 1923 3702 1924 3703
rect 1871 3700 1924 3702
rect 1871 3699 1872 3700
rect 1866 3698 1872 3699
rect 1923 3699 1924 3700
rect 1928 3699 1929 3703
rect 2107 3703 2108 3707
rect 2112 3706 2113 3707
rect 2138 3707 2144 3708
rect 2138 3706 2139 3707
rect 2112 3704 2139 3706
rect 2112 3703 2113 3704
rect 2107 3702 2113 3703
rect 2138 3703 2139 3704
rect 2143 3703 2144 3707
rect 2138 3702 2144 3703
rect 2146 3707 2152 3708
rect 2146 3703 2147 3707
rect 2151 3706 2152 3707
rect 2299 3707 2305 3708
rect 2299 3706 2300 3707
rect 2151 3704 2300 3706
rect 2151 3703 2152 3704
rect 2146 3702 2152 3703
rect 2299 3703 2300 3704
rect 2304 3703 2305 3707
rect 2299 3702 2305 3703
rect 2338 3707 2344 3708
rect 2338 3703 2339 3707
rect 2343 3706 2344 3707
rect 2515 3707 2521 3708
rect 2515 3706 2516 3707
rect 2343 3704 2516 3706
rect 2343 3703 2344 3704
rect 2338 3702 2344 3703
rect 2515 3703 2516 3704
rect 2520 3703 2521 3707
rect 2515 3702 2521 3703
rect 2623 3707 2629 3708
rect 2623 3703 2624 3707
rect 2628 3706 2629 3707
rect 2731 3707 2737 3708
rect 2731 3706 2732 3707
rect 2628 3704 2732 3706
rect 2628 3703 2629 3704
rect 2623 3702 2629 3703
rect 2731 3703 2732 3704
rect 2736 3703 2737 3707
rect 2986 3707 2992 3708
rect 2731 3702 2737 3703
rect 2947 3705 2953 3706
rect 2947 3701 2948 3705
rect 2952 3701 2953 3705
rect 2986 3703 2987 3707
rect 2991 3706 2992 3707
rect 3155 3707 3161 3708
rect 3155 3706 3156 3707
rect 2991 3704 3156 3706
rect 2991 3703 2992 3704
rect 2986 3702 2992 3703
rect 3155 3703 3156 3704
rect 3160 3703 3161 3707
rect 3394 3707 3400 3708
rect 3155 3702 3161 3703
rect 3355 3705 3361 3706
rect 2947 3700 2953 3701
rect 3355 3701 3356 3705
rect 3360 3701 3361 3705
rect 3394 3703 3395 3707
rect 3399 3706 3400 3707
rect 3555 3707 3561 3708
rect 3555 3706 3556 3707
rect 3399 3704 3556 3706
rect 3399 3703 3400 3704
rect 3394 3702 3400 3703
rect 3555 3703 3556 3704
rect 3560 3703 3561 3707
rect 3555 3702 3561 3703
rect 3763 3707 3769 3708
rect 3763 3703 3764 3707
rect 3768 3706 3769 3707
rect 3802 3707 3808 3708
rect 3802 3706 3803 3707
rect 3768 3704 3803 3706
rect 3768 3703 3769 3704
rect 3763 3702 3769 3703
rect 3802 3703 3803 3704
rect 3807 3703 3808 3707
rect 3802 3702 3808 3703
rect 3355 3700 3361 3701
rect 1923 3698 1929 3699
rect 2948 3698 2950 3700
rect 3018 3699 3024 3700
rect 3018 3698 3019 3699
rect 2948 3696 3019 3698
rect 3018 3695 3019 3696
rect 3023 3695 3024 3699
rect 3356 3698 3358 3700
rect 3618 3699 3624 3700
rect 3618 3698 3619 3699
rect 3356 3696 3619 3698
rect 3018 3694 3024 3695
rect 3618 3695 3619 3696
rect 3623 3695 3624 3699
rect 3618 3694 3624 3695
rect 2046 3688 2052 3689
rect 3942 3688 3948 3689
rect 618 3687 624 3688
rect 618 3686 619 3687
rect 404 3684 619 3686
rect 404 3682 406 3684
rect 618 3683 619 3684
rect 623 3683 624 3687
rect 1458 3687 1464 3688
rect 1458 3686 1459 3687
rect 618 3682 624 3683
rect 1212 3684 1459 3686
rect 1212 3682 1214 3684
rect 1458 3683 1459 3684
rect 1463 3683 1464 3687
rect 2046 3684 2047 3688
rect 2051 3684 2052 3688
rect 2046 3683 2052 3684
rect 2070 3687 2076 3688
rect 2070 3683 2071 3687
rect 2075 3683 2076 3687
rect 1458 3682 1464 3683
rect 2070 3682 2076 3683
rect 2262 3687 2268 3688
rect 2262 3683 2263 3687
rect 2267 3683 2268 3687
rect 2262 3682 2268 3683
rect 2478 3687 2484 3688
rect 2478 3683 2479 3687
rect 2483 3683 2484 3687
rect 2478 3682 2484 3683
rect 2694 3687 2700 3688
rect 2694 3683 2695 3687
rect 2699 3683 2700 3687
rect 2694 3682 2700 3683
rect 2910 3687 2916 3688
rect 2910 3683 2911 3687
rect 2915 3683 2916 3687
rect 2910 3682 2916 3683
rect 3118 3687 3124 3688
rect 3118 3683 3119 3687
rect 3123 3683 3124 3687
rect 3118 3682 3124 3683
rect 3318 3687 3324 3688
rect 3318 3683 3319 3687
rect 3323 3683 3324 3687
rect 3318 3682 3324 3683
rect 3518 3687 3524 3688
rect 3518 3683 3519 3687
rect 3523 3683 3524 3687
rect 3518 3682 3524 3683
rect 3726 3687 3732 3688
rect 3726 3683 3727 3687
rect 3731 3683 3732 3687
rect 3942 3684 3943 3688
rect 3947 3684 3948 3688
rect 3942 3683 3948 3684
rect 3726 3682 3732 3683
rect 403 3681 409 3682
rect 403 3677 404 3681
rect 408 3677 409 3681
rect 1211 3681 1217 3682
rect 403 3676 409 3677
rect 442 3679 448 3680
rect 442 3675 443 3679
rect 447 3678 448 3679
rect 555 3679 561 3680
rect 555 3678 556 3679
rect 447 3676 556 3678
rect 447 3675 448 3676
rect 442 3674 448 3675
rect 555 3675 556 3676
rect 560 3675 561 3679
rect 555 3674 561 3675
rect 715 3679 721 3680
rect 715 3675 716 3679
rect 720 3678 721 3679
rect 762 3679 768 3680
rect 762 3678 763 3679
rect 720 3676 763 3678
rect 720 3675 721 3676
rect 715 3674 721 3675
rect 762 3675 763 3676
rect 767 3675 768 3679
rect 762 3674 768 3675
rect 883 3679 889 3680
rect 883 3675 884 3679
rect 888 3678 889 3679
rect 935 3679 941 3680
rect 935 3678 936 3679
rect 888 3676 936 3678
rect 888 3675 889 3676
rect 883 3674 889 3675
rect 935 3675 936 3676
rect 940 3675 941 3679
rect 935 3674 941 3675
rect 1051 3679 1057 3680
rect 1051 3675 1052 3679
rect 1056 3678 1057 3679
rect 1103 3679 1109 3680
rect 1103 3678 1104 3679
rect 1056 3676 1104 3678
rect 1056 3675 1057 3676
rect 1051 3674 1057 3675
rect 1103 3675 1104 3676
rect 1108 3675 1109 3679
rect 1211 3677 1212 3681
rect 1216 3677 1217 3681
rect 1211 3676 1217 3677
rect 1250 3679 1256 3680
rect 1103 3674 1109 3675
rect 1250 3675 1251 3679
rect 1255 3678 1256 3679
rect 1363 3679 1369 3680
rect 1363 3678 1364 3679
rect 1255 3676 1364 3678
rect 1255 3675 1256 3676
rect 1250 3674 1256 3675
rect 1363 3675 1364 3676
rect 1368 3675 1369 3679
rect 1363 3674 1369 3675
rect 1402 3679 1408 3680
rect 1402 3675 1403 3679
rect 1407 3678 1408 3679
rect 1515 3679 1521 3680
rect 1515 3678 1516 3679
rect 1407 3676 1516 3678
rect 1407 3675 1408 3676
rect 1402 3674 1408 3675
rect 1515 3675 1516 3676
rect 1520 3675 1521 3679
rect 1515 3674 1521 3675
rect 1554 3679 1560 3680
rect 1554 3675 1555 3679
rect 1559 3678 1560 3679
rect 1667 3679 1673 3680
rect 1667 3678 1668 3679
rect 1559 3676 1668 3678
rect 1559 3675 1560 3676
rect 1554 3674 1560 3675
rect 1667 3675 1668 3676
rect 1672 3675 1673 3679
rect 1667 3674 1673 3675
rect 1706 3679 1712 3680
rect 1706 3675 1707 3679
rect 1711 3678 1712 3679
rect 1827 3679 1833 3680
rect 1827 3678 1828 3679
rect 1711 3676 1828 3678
rect 1711 3675 1712 3676
rect 1706 3674 1712 3675
rect 1827 3675 1828 3676
rect 1832 3675 1833 3679
rect 1827 3674 1833 3675
rect 2146 3679 2152 3680
rect 2146 3675 2147 3679
rect 2151 3675 2152 3679
rect 2146 3674 2152 3675
rect 2338 3679 2344 3680
rect 2338 3675 2339 3679
rect 2343 3675 2344 3679
rect 2623 3679 2629 3680
rect 2623 3678 2624 3679
rect 2557 3676 2624 3678
rect 2338 3674 2344 3675
rect 2623 3675 2624 3676
rect 2628 3675 2629 3679
rect 2623 3674 2629 3675
rect 2662 3679 2668 3680
rect 2662 3675 2663 3679
rect 2667 3678 2668 3679
rect 2986 3679 2992 3680
rect 2667 3676 2737 3678
rect 2667 3675 2668 3676
rect 2662 3674 2668 3675
rect 2986 3675 2987 3679
rect 2991 3675 2992 3679
rect 2986 3674 2992 3675
rect 3194 3679 3200 3680
rect 3194 3675 3195 3679
rect 3199 3675 3200 3679
rect 3194 3674 3200 3675
rect 3394 3679 3400 3680
rect 3394 3675 3395 3679
rect 3399 3675 3400 3679
rect 3618 3679 3624 3680
rect 3394 3674 3400 3675
rect 3594 3675 3600 3676
rect 2046 3671 2052 3672
rect 2046 3667 2047 3671
rect 2051 3667 2052 3671
rect 3594 3671 3595 3675
rect 3599 3671 3600 3675
rect 3618 3675 3619 3679
rect 3623 3678 3624 3679
rect 3623 3676 3769 3678
rect 3623 3675 3624 3676
rect 3618 3674 3624 3675
rect 3594 3670 3600 3671
rect 3942 3671 3948 3672
rect 2046 3666 2052 3667
rect 2070 3668 2076 3669
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 2262 3668 2268 3669
rect 2262 3664 2263 3668
rect 2267 3664 2268 3668
rect 2262 3663 2268 3664
rect 2478 3668 2484 3669
rect 2478 3664 2479 3668
rect 2483 3664 2484 3668
rect 2478 3663 2484 3664
rect 2694 3668 2700 3669
rect 2694 3664 2695 3668
rect 2699 3664 2700 3668
rect 2694 3663 2700 3664
rect 2910 3668 2916 3669
rect 2910 3664 2911 3668
rect 2915 3664 2916 3668
rect 2910 3663 2916 3664
rect 3118 3668 3124 3669
rect 3118 3664 3119 3668
rect 3123 3664 3124 3668
rect 3118 3663 3124 3664
rect 3318 3668 3324 3669
rect 3318 3664 3319 3668
rect 3323 3664 3324 3668
rect 3318 3663 3324 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3726 3668 3732 3669
rect 3726 3664 3727 3668
rect 3731 3664 3732 3668
rect 3942 3667 3943 3671
rect 3947 3667 3948 3671
rect 3942 3666 3948 3667
rect 3726 3663 3732 3664
rect 110 3660 116 3661
rect 2006 3660 2012 3661
rect 110 3656 111 3660
rect 115 3656 116 3660
rect 110 3655 116 3656
rect 366 3659 372 3660
rect 366 3655 367 3659
rect 371 3655 372 3659
rect 366 3654 372 3655
rect 518 3659 524 3660
rect 518 3655 519 3659
rect 523 3655 524 3659
rect 518 3654 524 3655
rect 678 3659 684 3660
rect 678 3655 679 3659
rect 683 3655 684 3659
rect 678 3654 684 3655
rect 846 3659 852 3660
rect 846 3655 847 3659
rect 851 3655 852 3659
rect 846 3654 852 3655
rect 1014 3659 1020 3660
rect 1014 3655 1015 3659
rect 1019 3655 1020 3659
rect 1014 3654 1020 3655
rect 1174 3659 1180 3660
rect 1174 3655 1175 3659
rect 1179 3655 1180 3659
rect 1174 3654 1180 3655
rect 1326 3659 1332 3660
rect 1326 3655 1327 3659
rect 1331 3655 1332 3659
rect 1326 3654 1332 3655
rect 1478 3659 1484 3660
rect 1478 3655 1479 3659
rect 1483 3655 1484 3659
rect 1478 3654 1484 3655
rect 1630 3659 1636 3660
rect 1630 3655 1631 3659
rect 1635 3655 1636 3659
rect 1630 3654 1636 3655
rect 1790 3659 1796 3660
rect 1790 3655 1791 3659
rect 1795 3655 1796 3659
rect 2006 3656 2007 3660
rect 2011 3656 2012 3660
rect 2006 3655 2012 3656
rect 1790 3654 1796 3655
rect 442 3651 448 3652
rect 442 3647 443 3651
rect 447 3647 448 3651
rect 618 3651 624 3652
rect 442 3646 448 3647
rect 594 3647 600 3648
rect 110 3643 116 3644
rect 110 3639 111 3643
rect 115 3639 116 3643
rect 594 3643 595 3647
rect 599 3643 600 3647
rect 618 3647 619 3651
rect 623 3650 624 3651
rect 762 3651 768 3652
rect 623 3648 721 3650
rect 623 3647 624 3648
rect 618 3646 624 3647
rect 762 3647 763 3651
rect 767 3650 768 3651
rect 935 3651 941 3652
rect 767 3648 889 3650
rect 767 3647 768 3648
rect 762 3646 768 3647
rect 935 3647 936 3651
rect 940 3650 941 3651
rect 1250 3651 1256 3652
rect 940 3648 1057 3650
rect 940 3647 941 3648
rect 935 3646 941 3647
rect 1250 3647 1251 3651
rect 1255 3647 1256 3651
rect 1250 3646 1256 3647
rect 1402 3651 1408 3652
rect 1402 3647 1403 3651
rect 1407 3647 1408 3651
rect 1402 3646 1408 3647
rect 1554 3651 1560 3652
rect 1554 3647 1555 3651
rect 1559 3647 1560 3651
rect 1554 3646 1560 3647
rect 1706 3651 1712 3652
rect 1706 3647 1707 3651
rect 1711 3647 1712 3651
rect 1706 3646 1712 3647
rect 1866 3651 1872 3652
rect 1866 3647 1867 3651
rect 1871 3647 1872 3651
rect 1866 3646 1872 3647
rect 594 3642 600 3643
rect 2006 3643 2012 3644
rect 110 3638 116 3639
rect 366 3640 372 3641
rect 366 3636 367 3640
rect 371 3636 372 3640
rect 366 3635 372 3636
rect 518 3640 524 3641
rect 518 3636 519 3640
rect 523 3636 524 3640
rect 518 3635 524 3636
rect 678 3640 684 3641
rect 678 3636 679 3640
rect 683 3636 684 3640
rect 678 3635 684 3636
rect 846 3640 852 3641
rect 846 3636 847 3640
rect 851 3636 852 3640
rect 846 3635 852 3636
rect 1014 3640 1020 3641
rect 1014 3636 1015 3640
rect 1019 3636 1020 3640
rect 1014 3635 1020 3636
rect 1174 3640 1180 3641
rect 1174 3636 1175 3640
rect 1179 3636 1180 3640
rect 1174 3635 1180 3636
rect 1326 3640 1332 3641
rect 1326 3636 1327 3640
rect 1331 3636 1332 3640
rect 1326 3635 1332 3636
rect 1478 3640 1484 3641
rect 1478 3636 1479 3640
rect 1483 3636 1484 3640
rect 1478 3635 1484 3636
rect 1630 3640 1636 3641
rect 1630 3636 1631 3640
rect 1635 3636 1636 3640
rect 1630 3635 1636 3636
rect 1790 3640 1796 3641
rect 1790 3636 1791 3640
rect 1795 3636 1796 3640
rect 2006 3639 2007 3643
rect 2011 3639 2012 3643
rect 2006 3638 2012 3639
rect 1790 3635 1796 3636
rect 2110 3604 2116 3605
rect 2046 3601 2052 3602
rect 2046 3597 2047 3601
rect 2051 3597 2052 3601
rect 2110 3600 2111 3604
rect 2115 3600 2116 3604
rect 2110 3599 2116 3600
rect 2270 3604 2276 3605
rect 2270 3600 2271 3604
rect 2275 3600 2276 3604
rect 2270 3599 2276 3600
rect 2454 3604 2460 3605
rect 2454 3600 2455 3604
rect 2459 3600 2460 3604
rect 2454 3599 2460 3600
rect 2654 3604 2660 3605
rect 2654 3600 2655 3604
rect 2659 3600 2660 3604
rect 2654 3599 2660 3600
rect 2870 3604 2876 3605
rect 2870 3600 2871 3604
rect 2875 3600 2876 3604
rect 2870 3599 2876 3600
rect 3094 3604 3100 3605
rect 3094 3600 3095 3604
rect 3099 3600 3100 3604
rect 3094 3599 3100 3600
rect 3326 3604 3332 3605
rect 3326 3600 3327 3604
rect 3331 3600 3332 3604
rect 3326 3599 3332 3600
rect 3566 3604 3572 3605
rect 3566 3600 3567 3604
rect 3571 3600 3572 3604
rect 3566 3599 3572 3600
rect 3942 3601 3948 3602
rect 2046 3596 2052 3597
rect 3942 3597 3943 3601
rect 3947 3597 3948 3601
rect 3942 3596 3948 3597
rect 2186 3595 2192 3596
rect 2186 3591 2187 3595
rect 2191 3591 2192 3595
rect 2186 3590 2192 3591
rect 2346 3595 2352 3596
rect 2346 3591 2347 3595
rect 2351 3591 2352 3595
rect 2346 3590 2352 3591
rect 2530 3595 2536 3596
rect 2530 3591 2531 3595
rect 2535 3591 2536 3595
rect 2530 3590 2536 3591
rect 2730 3595 2736 3596
rect 2730 3591 2731 3595
rect 2735 3591 2736 3595
rect 2730 3590 2736 3591
rect 2862 3595 2868 3596
rect 2862 3591 2863 3595
rect 2867 3594 2868 3595
rect 3018 3595 3024 3596
rect 2867 3592 2913 3594
rect 2867 3591 2868 3592
rect 2862 3590 2868 3591
rect 3018 3591 3019 3595
rect 3023 3594 3024 3595
rect 3394 3595 3400 3596
rect 3023 3592 3137 3594
rect 3023 3591 3024 3592
rect 3018 3590 3024 3591
rect 3394 3591 3395 3595
rect 3399 3591 3400 3595
rect 3394 3590 3400 3591
rect 3423 3595 3429 3596
rect 3423 3591 3424 3595
rect 3428 3594 3429 3595
rect 3428 3592 3609 3594
rect 3428 3591 3429 3592
rect 3423 3590 3429 3591
rect 2110 3585 2116 3586
rect 2046 3584 2052 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2110 3581 2111 3585
rect 2115 3581 2116 3585
rect 2110 3580 2116 3581
rect 2270 3585 2276 3586
rect 2270 3581 2271 3585
rect 2275 3581 2276 3585
rect 2270 3580 2276 3581
rect 2454 3585 2460 3586
rect 2454 3581 2455 3585
rect 2459 3581 2460 3585
rect 2454 3580 2460 3581
rect 2654 3585 2660 3586
rect 2654 3581 2655 3585
rect 2659 3581 2660 3585
rect 2654 3580 2660 3581
rect 2870 3585 2876 3586
rect 2870 3581 2871 3585
rect 2875 3581 2876 3585
rect 2870 3580 2876 3581
rect 3094 3585 3100 3586
rect 3094 3581 3095 3585
rect 3099 3581 3100 3585
rect 3094 3580 3100 3581
rect 3326 3585 3332 3586
rect 3326 3581 3327 3585
rect 3331 3581 3332 3585
rect 3326 3580 3332 3581
rect 3566 3585 3572 3586
rect 3566 3581 3567 3585
rect 3571 3581 3572 3585
rect 3566 3580 3572 3581
rect 3942 3584 3948 3585
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 2046 3579 2052 3580
rect 3942 3579 3948 3580
rect 2662 3575 2668 3576
rect 2662 3574 2663 3575
rect 270 3572 276 3573
rect 110 3569 116 3570
rect 110 3565 111 3569
rect 115 3565 116 3569
rect 270 3568 271 3572
rect 275 3568 276 3572
rect 270 3567 276 3568
rect 414 3572 420 3573
rect 414 3568 415 3572
rect 419 3568 420 3572
rect 414 3567 420 3568
rect 574 3572 580 3573
rect 574 3568 575 3572
rect 579 3568 580 3572
rect 574 3567 580 3568
rect 734 3572 740 3573
rect 734 3568 735 3572
rect 739 3568 740 3572
rect 734 3567 740 3568
rect 894 3572 900 3573
rect 894 3568 895 3572
rect 899 3568 900 3572
rect 894 3567 900 3568
rect 1054 3572 1060 3573
rect 1054 3568 1055 3572
rect 1059 3568 1060 3572
rect 1054 3567 1060 3568
rect 1214 3572 1220 3573
rect 1214 3568 1215 3572
rect 1219 3568 1220 3572
rect 1214 3567 1220 3568
rect 1374 3572 1380 3573
rect 1374 3568 1375 3572
rect 1379 3568 1380 3572
rect 1374 3567 1380 3568
rect 1542 3572 1548 3573
rect 1542 3568 1543 3572
rect 1547 3568 1548 3572
rect 2180 3572 2663 3574
rect 1542 3567 1548 3568
rect 2006 3569 2012 3570
rect 110 3564 116 3565
rect 2006 3565 2007 3569
rect 2011 3565 2012 3569
rect 2006 3564 2012 3565
rect 2147 3567 2153 3568
rect 346 3563 352 3564
rect 346 3559 347 3563
rect 351 3559 352 3563
rect 346 3558 352 3559
rect 482 3563 488 3564
rect 482 3559 483 3563
rect 487 3559 488 3563
rect 482 3558 488 3559
rect 650 3563 656 3564
rect 650 3559 651 3563
rect 655 3559 656 3563
rect 650 3558 656 3559
rect 810 3563 816 3564
rect 810 3559 811 3563
rect 815 3559 816 3563
rect 810 3558 816 3559
rect 818 3563 824 3564
rect 818 3559 819 3563
rect 823 3562 824 3563
rect 1130 3563 1136 3564
rect 823 3560 937 3562
rect 823 3559 824 3560
rect 818 3558 824 3559
rect 1130 3559 1131 3563
rect 1135 3559 1136 3563
rect 1130 3558 1136 3559
rect 1290 3563 1296 3564
rect 1290 3559 1291 3563
rect 1295 3559 1296 3563
rect 1290 3558 1296 3559
rect 1450 3563 1456 3564
rect 1450 3559 1451 3563
rect 1455 3559 1456 3563
rect 1450 3558 1456 3559
rect 1458 3563 1464 3564
rect 1458 3559 1459 3563
rect 1463 3562 1464 3563
rect 2147 3563 2148 3567
rect 2152 3566 2153 3567
rect 2180 3566 2182 3572
rect 2662 3571 2663 3572
rect 2667 3571 2668 3575
rect 2662 3570 2668 3571
rect 2152 3564 2182 3566
rect 2186 3567 2192 3568
rect 2152 3563 2153 3564
rect 2147 3562 2153 3563
rect 2186 3563 2187 3567
rect 2191 3566 2192 3567
rect 2307 3567 2313 3568
rect 2307 3566 2308 3567
rect 2191 3564 2308 3566
rect 2191 3563 2192 3564
rect 2186 3562 2192 3563
rect 2307 3563 2308 3564
rect 2312 3563 2313 3567
rect 2307 3562 2313 3563
rect 2346 3567 2352 3568
rect 2346 3563 2347 3567
rect 2351 3566 2352 3567
rect 2491 3567 2497 3568
rect 2491 3566 2492 3567
rect 2351 3564 2492 3566
rect 2351 3563 2352 3564
rect 2346 3562 2352 3563
rect 2491 3563 2492 3564
rect 2496 3563 2497 3567
rect 2491 3562 2497 3563
rect 2530 3567 2536 3568
rect 2530 3563 2531 3567
rect 2535 3566 2536 3567
rect 2691 3567 2697 3568
rect 2691 3566 2692 3567
rect 2535 3564 2692 3566
rect 2535 3563 2536 3564
rect 2530 3562 2536 3563
rect 2691 3563 2692 3564
rect 2696 3563 2697 3567
rect 2691 3562 2697 3563
rect 2730 3567 2736 3568
rect 2730 3563 2731 3567
rect 2735 3566 2736 3567
rect 2907 3567 2913 3568
rect 2907 3566 2908 3567
rect 2735 3564 2908 3566
rect 2735 3563 2736 3564
rect 2730 3562 2736 3563
rect 2907 3563 2908 3564
rect 2912 3563 2913 3567
rect 3363 3567 3369 3568
rect 2907 3562 2913 3563
rect 3131 3563 3137 3564
rect 1463 3560 1585 3562
rect 1463 3559 1464 3560
rect 1458 3558 1464 3559
rect 3131 3559 3132 3563
rect 3136 3562 3137 3563
rect 3190 3563 3196 3564
rect 3190 3562 3191 3563
rect 3136 3560 3191 3562
rect 3136 3559 3137 3560
rect 3131 3558 3137 3559
rect 3190 3559 3191 3560
rect 3195 3559 3196 3563
rect 3363 3563 3364 3567
rect 3368 3566 3369 3567
rect 3423 3567 3429 3568
rect 3423 3566 3424 3567
rect 3368 3564 3424 3566
rect 3368 3563 3369 3564
rect 3363 3562 3369 3563
rect 3423 3563 3424 3564
rect 3428 3563 3429 3567
rect 3423 3562 3429 3563
rect 3594 3567 3600 3568
rect 3594 3563 3595 3567
rect 3599 3566 3600 3567
rect 3603 3567 3609 3568
rect 3603 3566 3604 3567
rect 3599 3564 3604 3566
rect 3599 3563 3600 3564
rect 3594 3562 3600 3563
rect 3603 3563 3604 3564
rect 3608 3563 3609 3567
rect 3603 3562 3609 3563
rect 3190 3558 3196 3559
rect 270 3553 276 3554
rect 110 3552 116 3553
rect 110 3548 111 3552
rect 115 3548 116 3552
rect 270 3549 271 3553
rect 275 3549 276 3553
rect 270 3548 276 3549
rect 414 3553 420 3554
rect 414 3549 415 3553
rect 419 3549 420 3553
rect 414 3548 420 3549
rect 574 3553 580 3554
rect 574 3549 575 3553
rect 579 3549 580 3553
rect 574 3548 580 3549
rect 734 3553 740 3554
rect 734 3549 735 3553
rect 739 3549 740 3553
rect 734 3548 740 3549
rect 894 3553 900 3554
rect 894 3549 895 3553
rect 899 3549 900 3553
rect 894 3548 900 3549
rect 1054 3553 1060 3554
rect 1054 3549 1055 3553
rect 1059 3549 1060 3553
rect 1054 3548 1060 3549
rect 1214 3553 1220 3554
rect 1214 3549 1215 3553
rect 1219 3549 1220 3553
rect 1214 3548 1220 3549
rect 1374 3553 1380 3554
rect 1374 3549 1375 3553
rect 1379 3549 1380 3553
rect 1374 3548 1380 3549
rect 1542 3553 1548 3554
rect 1542 3549 1543 3553
rect 1547 3549 1548 3553
rect 1542 3548 1548 3549
rect 2006 3552 2012 3553
rect 2006 3548 2007 3552
rect 2011 3548 2012 3552
rect 110 3547 116 3548
rect 2006 3547 2012 3548
rect 818 3543 824 3544
rect 818 3542 819 3543
rect 319 3540 819 3542
rect 307 3535 313 3536
rect 307 3531 308 3535
rect 312 3534 313 3535
rect 319 3534 321 3540
rect 818 3539 819 3540
rect 823 3539 824 3543
rect 818 3538 824 3539
rect 1130 3539 1136 3540
rect 312 3532 321 3534
rect 346 3535 352 3536
rect 312 3531 313 3532
rect 307 3530 313 3531
rect 346 3531 347 3535
rect 351 3534 352 3535
rect 451 3535 457 3536
rect 451 3534 452 3535
rect 351 3532 452 3534
rect 351 3531 352 3532
rect 346 3530 352 3531
rect 451 3531 452 3532
rect 456 3531 457 3535
rect 451 3530 457 3531
rect 594 3535 600 3536
rect 594 3531 595 3535
rect 599 3534 600 3535
rect 611 3535 617 3536
rect 611 3534 612 3535
rect 599 3532 612 3534
rect 599 3531 600 3532
rect 594 3530 600 3531
rect 611 3531 612 3532
rect 616 3531 617 3535
rect 611 3530 617 3531
rect 650 3535 656 3536
rect 650 3531 651 3535
rect 655 3534 656 3535
rect 771 3535 777 3536
rect 771 3534 772 3535
rect 655 3532 772 3534
rect 655 3531 656 3532
rect 650 3530 656 3531
rect 771 3531 772 3532
rect 776 3531 777 3535
rect 771 3530 777 3531
rect 810 3535 816 3536
rect 810 3531 811 3535
rect 815 3534 816 3535
rect 931 3535 937 3536
rect 931 3534 932 3535
rect 815 3532 932 3534
rect 815 3531 816 3532
rect 810 3530 816 3531
rect 931 3531 932 3532
rect 936 3531 937 3535
rect 1130 3535 1131 3539
rect 1135 3535 1136 3539
rect 1130 3534 1136 3535
rect 1251 3535 1257 3536
rect 1251 3534 1252 3535
rect 1132 3532 1252 3534
rect 931 3530 937 3531
rect 1091 3531 1097 3532
rect 1091 3527 1092 3531
rect 1096 3530 1097 3531
rect 1251 3531 1252 3532
rect 1256 3531 1257 3535
rect 1251 3530 1257 3531
rect 1290 3535 1296 3536
rect 1290 3531 1291 3535
rect 1295 3534 1296 3535
rect 1411 3535 1417 3536
rect 1411 3534 1412 3535
rect 1295 3532 1412 3534
rect 1295 3531 1296 3532
rect 1290 3530 1296 3531
rect 1411 3531 1412 3532
rect 1416 3531 1417 3535
rect 1411 3530 1417 3531
rect 1450 3535 1456 3536
rect 1450 3531 1451 3535
rect 1455 3534 1456 3535
rect 1579 3535 1585 3536
rect 1579 3534 1580 3535
rect 1455 3532 1580 3534
rect 1455 3531 1456 3532
rect 1450 3530 1456 3531
rect 1579 3531 1580 3532
rect 1584 3531 1585 3535
rect 1579 3530 1585 3531
rect 2323 3535 2329 3536
rect 2323 3531 2324 3535
rect 2328 3534 2329 3535
rect 2354 3535 2360 3536
rect 2354 3534 2355 3535
rect 2328 3532 2355 3534
rect 2328 3531 2329 3532
rect 2323 3530 2329 3531
rect 2354 3531 2355 3532
rect 2359 3531 2360 3535
rect 2354 3530 2360 3531
rect 2362 3535 2368 3536
rect 2362 3531 2363 3535
rect 2367 3534 2368 3535
rect 2419 3535 2425 3536
rect 2419 3534 2420 3535
rect 2367 3532 2420 3534
rect 2367 3531 2368 3532
rect 2362 3530 2368 3531
rect 2419 3531 2420 3532
rect 2424 3531 2425 3535
rect 2419 3530 2425 3531
rect 2466 3535 2472 3536
rect 2466 3531 2467 3535
rect 2471 3534 2472 3535
rect 2515 3535 2521 3536
rect 2515 3534 2516 3535
rect 2471 3532 2516 3534
rect 2471 3531 2472 3532
rect 2466 3530 2472 3531
rect 2515 3531 2516 3532
rect 2520 3531 2521 3535
rect 2515 3530 2521 3531
rect 2554 3535 2560 3536
rect 2554 3531 2555 3535
rect 2559 3534 2560 3535
rect 2611 3535 2617 3536
rect 2611 3534 2612 3535
rect 2559 3532 2612 3534
rect 2559 3531 2560 3532
rect 2554 3530 2560 3531
rect 2611 3531 2612 3532
rect 2616 3531 2617 3535
rect 2611 3530 2617 3531
rect 2707 3535 2713 3536
rect 2707 3531 2708 3535
rect 2712 3534 2713 3535
rect 2738 3535 2744 3536
rect 2738 3534 2739 3535
rect 2712 3532 2739 3534
rect 2712 3531 2713 3532
rect 2707 3530 2713 3531
rect 2738 3531 2739 3532
rect 2743 3531 2744 3535
rect 2738 3530 2744 3531
rect 2746 3535 2752 3536
rect 2746 3531 2747 3535
rect 2751 3534 2752 3535
rect 2803 3535 2809 3536
rect 2803 3534 2804 3535
rect 2751 3532 2804 3534
rect 2751 3531 2752 3532
rect 2746 3530 2752 3531
rect 2803 3531 2804 3532
rect 2808 3531 2809 3535
rect 2803 3530 2809 3531
rect 2842 3535 2848 3536
rect 2842 3531 2843 3535
rect 2847 3534 2848 3535
rect 2907 3535 2913 3536
rect 2907 3534 2908 3535
rect 2847 3532 2908 3534
rect 2847 3531 2848 3532
rect 2842 3530 2848 3531
rect 2907 3531 2908 3532
rect 2912 3531 2913 3535
rect 2907 3530 2913 3531
rect 2946 3535 2952 3536
rect 2946 3531 2947 3535
rect 2951 3534 2952 3535
rect 3019 3535 3025 3536
rect 3019 3534 3020 3535
rect 2951 3532 3020 3534
rect 2951 3531 2952 3532
rect 2946 3530 2952 3531
rect 3019 3531 3020 3532
rect 3024 3531 3025 3535
rect 3019 3530 3025 3531
rect 3058 3535 3064 3536
rect 3058 3531 3059 3535
rect 3063 3534 3064 3535
rect 3139 3535 3145 3536
rect 3139 3534 3140 3535
rect 3063 3532 3140 3534
rect 3063 3531 3064 3532
rect 3058 3530 3064 3531
rect 3139 3531 3140 3532
rect 3144 3531 3145 3535
rect 3139 3530 3145 3531
rect 3230 3535 3236 3536
rect 3230 3531 3231 3535
rect 3235 3534 3236 3535
rect 3259 3535 3265 3536
rect 3259 3534 3260 3535
rect 3235 3532 3260 3534
rect 3235 3531 3236 3532
rect 3230 3530 3236 3531
rect 3259 3531 3260 3532
rect 3264 3531 3265 3535
rect 3259 3530 3265 3531
rect 3387 3535 3396 3536
rect 3387 3531 3388 3535
rect 3395 3531 3396 3535
rect 3387 3530 3396 3531
rect 3426 3535 3432 3536
rect 3426 3531 3427 3535
rect 3431 3534 3432 3535
rect 3523 3535 3529 3536
rect 3523 3534 3524 3535
rect 3431 3532 3524 3534
rect 3431 3531 3432 3532
rect 3426 3530 3432 3531
rect 3523 3531 3524 3532
rect 3528 3531 3529 3535
rect 3523 3530 3529 3531
rect 1096 3528 1161 3530
rect 1096 3527 1097 3528
rect 1091 3526 1097 3527
rect 1159 3526 1161 3528
rect 1338 3527 1344 3528
rect 1338 3526 1339 3527
rect 1159 3524 1339 3526
rect 1338 3523 1339 3524
rect 1343 3523 1344 3527
rect 1338 3522 1344 3523
rect 2046 3516 2052 3517
rect 3942 3516 3948 3517
rect 2046 3512 2047 3516
rect 2051 3512 2052 3516
rect 234 3511 240 3512
rect 195 3509 201 3510
rect 195 3505 196 3509
rect 200 3505 201 3509
rect 234 3507 235 3511
rect 239 3510 240 3511
rect 323 3511 329 3512
rect 323 3510 324 3511
rect 239 3508 324 3510
rect 239 3507 240 3508
rect 234 3506 240 3507
rect 323 3507 324 3508
rect 328 3507 329 3511
rect 323 3506 329 3507
rect 459 3511 465 3512
rect 459 3507 460 3511
rect 464 3510 465 3511
rect 482 3511 488 3512
rect 482 3510 483 3511
rect 464 3508 483 3510
rect 464 3507 465 3508
rect 459 3506 465 3507
rect 482 3507 483 3508
rect 487 3507 488 3511
rect 482 3506 488 3507
rect 498 3511 504 3512
rect 498 3507 499 3511
rect 503 3510 504 3511
rect 595 3511 601 3512
rect 595 3510 596 3511
rect 503 3508 596 3510
rect 503 3507 504 3508
rect 498 3506 504 3507
rect 595 3507 596 3508
rect 600 3507 601 3511
rect 595 3506 601 3507
rect 634 3511 640 3512
rect 634 3507 635 3511
rect 639 3510 640 3511
rect 731 3511 737 3512
rect 731 3510 732 3511
rect 639 3508 732 3510
rect 639 3507 640 3508
rect 634 3506 640 3507
rect 731 3507 732 3508
rect 736 3507 737 3511
rect 731 3506 737 3507
rect 867 3511 873 3512
rect 867 3507 868 3511
rect 872 3510 873 3511
rect 882 3511 888 3512
rect 882 3510 883 3511
rect 872 3508 883 3510
rect 872 3507 873 3508
rect 867 3506 873 3507
rect 882 3507 883 3508
rect 887 3507 888 3511
rect 882 3506 888 3507
rect 906 3511 912 3512
rect 906 3507 907 3511
rect 911 3510 912 3511
rect 1003 3511 1009 3512
rect 1003 3510 1004 3511
rect 911 3508 1004 3510
rect 911 3507 912 3508
rect 906 3506 912 3507
rect 1003 3507 1004 3508
rect 1008 3507 1009 3511
rect 1003 3506 1009 3507
rect 1042 3511 1048 3512
rect 1042 3507 1043 3511
rect 1047 3510 1048 3511
rect 1131 3511 1137 3512
rect 1131 3510 1132 3511
rect 1047 3508 1132 3510
rect 1047 3507 1048 3508
rect 1042 3506 1048 3507
rect 1131 3507 1132 3508
rect 1136 3507 1137 3511
rect 1131 3506 1137 3507
rect 1170 3511 1176 3512
rect 1170 3507 1171 3511
rect 1175 3510 1176 3511
rect 1267 3511 1273 3512
rect 1267 3510 1268 3511
rect 1175 3508 1268 3510
rect 1175 3507 1176 3508
rect 1170 3506 1176 3507
rect 1267 3507 1268 3508
rect 1272 3507 1273 3511
rect 1267 3506 1273 3507
rect 1306 3511 1312 3512
rect 1306 3507 1307 3511
rect 1311 3510 1312 3511
rect 1403 3511 1409 3512
rect 2046 3511 2052 3512
rect 2286 3515 2292 3516
rect 2286 3511 2287 3515
rect 2291 3511 2292 3515
rect 1403 3510 1404 3511
rect 1311 3508 1404 3510
rect 1311 3507 1312 3508
rect 1306 3506 1312 3507
rect 1403 3507 1404 3508
rect 1408 3507 1409 3511
rect 2286 3510 2292 3511
rect 2382 3515 2388 3516
rect 2382 3511 2383 3515
rect 2387 3511 2388 3515
rect 2382 3510 2388 3511
rect 2478 3515 2484 3516
rect 2478 3511 2479 3515
rect 2483 3511 2484 3515
rect 2478 3510 2484 3511
rect 2574 3515 2580 3516
rect 2574 3511 2575 3515
rect 2579 3511 2580 3515
rect 2574 3510 2580 3511
rect 2670 3515 2676 3516
rect 2670 3511 2671 3515
rect 2675 3511 2676 3515
rect 2670 3510 2676 3511
rect 2766 3515 2772 3516
rect 2766 3511 2767 3515
rect 2771 3511 2772 3515
rect 2766 3510 2772 3511
rect 2870 3515 2876 3516
rect 2870 3511 2871 3515
rect 2875 3511 2876 3515
rect 2870 3510 2876 3511
rect 2982 3515 2988 3516
rect 2982 3511 2983 3515
rect 2987 3511 2988 3515
rect 2982 3510 2988 3511
rect 3102 3515 3108 3516
rect 3102 3511 3103 3515
rect 3107 3511 3108 3515
rect 3102 3510 3108 3511
rect 3222 3515 3228 3516
rect 3222 3511 3223 3515
rect 3227 3511 3228 3515
rect 3222 3510 3228 3511
rect 3350 3515 3356 3516
rect 3350 3511 3351 3515
rect 3355 3511 3356 3515
rect 3350 3510 3356 3511
rect 3486 3515 3492 3516
rect 3486 3511 3487 3515
rect 3491 3511 3492 3515
rect 3942 3512 3943 3516
rect 3947 3512 3948 3516
rect 3942 3511 3948 3512
rect 3486 3510 3492 3511
rect 1403 3506 1409 3507
rect 2362 3507 2368 3508
rect 195 3504 201 3505
rect 196 3502 198 3504
rect 642 3503 648 3504
rect 642 3502 643 3503
rect 196 3500 643 3502
rect 642 3499 643 3500
rect 647 3499 648 3503
rect 2362 3503 2363 3507
rect 2367 3503 2368 3507
rect 2466 3507 2472 3508
rect 2466 3506 2467 3507
rect 2461 3504 2467 3506
rect 2362 3502 2368 3503
rect 2466 3503 2467 3504
rect 2471 3503 2472 3507
rect 2466 3502 2472 3503
rect 2554 3507 2560 3508
rect 2554 3503 2555 3507
rect 2559 3503 2560 3507
rect 2746 3507 2752 3508
rect 2554 3502 2560 3503
rect 2568 3504 2617 3506
rect 642 3498 648 3499
rect 2046 3499 2052 3500
rect 2046 3495 2047 3499
rect 2051 3495 2052 3499
rect 2546 3499 2552 3500
rect 2046 3494 2052 3495
rect 2286 3496 2292 3497
rect 110 3492 116 3493
rect 2006 3492 2012 3493
rect 110 3488 111 3492
rect 115 3488 116 3492
rect 110 3487 116 3488
rect 158 3491 164 3492
rect 158 3487 159 3491
rect 163 3487 164 3491
rect 158 3486 164 3487
rect 286 3491 292 3492
rect 286 3487 287 3491
rect 291 3487 292 3491
rect 286 3486 292 3487
rect 422 3491 428 3492
rect 422 3487 423 3491
rect 427 3487 428 3491
rect 422 3486 428 3487
rect 558 3491 564 3492
rect 558 3487 559 3491
rect 563 3487 564 3491
rect 558 3486 564 3487
rect 694 3491 700 3492
rect 694 3487 695 3491
rect 699 3487 700 3491
rect 694 3486 700 3487
rect 830 3491 836 3492
rect 830 3487 831 3491
rect 835 3487 836 3491
rect 830 3486 836 3487
rect 966 3491 972 3492
rect 966 3487 967 3491
rect 971 3487 972 3491
rect 966 3486 972 3487
rect 1094 3491 1100 3492
rect 1094 3487 1095 3491
rect 1099 3487 1100 3491
rect 1094 3486 1100 3487
rect 1230 3491 1236 3492
rect 1230 3487 1231 3491
rect 1235 3487 1236 3491
rect 1230 3486 1236 3487
rect 1366 3491 1372 3492
rect 1366 3487 1367 3491
rect 1371 3487 1372 3491
rect 2006 3488 2007 3492
rect 2011 3488 2012 3492
rect 2286 3492 2287 3496
rect 2291 3492 2292 3496
rect 2286 3491 2292 3492
rect 2382 3496 2388 3497
rect 2382 3492 2383 3496
rect 2387 3492 2388 3496
rect 2382 3491 2388 3492
rect 2478 3496 2484 3497
rect 2478 3492 2479 3496
rect 2483 3492 2484 3496
rect 2546 3495 2547 3499
rect 2551 3498 2552 3499
rect 2568 3498 2570 3504
rect 2746 3503 2747 3507
rect 2751 3503 2752 3507
rect 2746 3502 2752 3503
rect 2842 3507 2848 3508
rect 2842 3503 2843 3507
rect 2847 3503 2848 3507
rect 2842 3502 2848 3503
rect 2946 3507 2952 3508
rect 2946 3503 2947 3507
rect 2951 3503 2952 3507
rect 2946 3502 2952 3503
rect 3058 3507 3064 3508
rect 3058 3503 3059 3507
rect 3063 3503 3064 3507
rect 3058 3502 3064 3503
rect 3066 3507 3072 3508
rect 3066 3503 3067 3507
rect 3071 3506 3072 3507
rect 3190 3507 3196 3508
rect 3071 3504 3145 3506
rect 3071 3503 3072 3504
rect 3066 3502 3072 3503
rect 3190 3503 3191 3507
rect 3195 3506 3196 3507
rect 3426 3507 3432 3508
rect 3195 3504 3265 3506
rect 3195 3503 3196 3504
rect 3190 3502 3196 3503
rect 3426 3503 3427 3507
rect 3431 3503 3432 3507
rect 3426 3502 3432 3503
rect 3466 3507 3472 3508
rect 3466 3503 3467 3507
rect 3471 3506 3472 3507
rect 3471 3504 3529 3506
rect 3471 3503 3472 3504
rect 3466 3502 3472 3503
rect 2551 3496 2570 3498
rect 3942 3499 3948 3500
rect 2574 3496 2580 3497
rect 2551 3495 2552 3496
rect 2546 3494 2552 3495
rect 2478 3491 2484 3492
rect 2574 3492 2575 3496
rect 2579 3492 2580 3496
rect 2574 3491 2580 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2766 3496 2772 3497
rect 2766 3492 2767 3496
rect 2771 3492 2772 3496
rect 2766 3491 2772 3492
rect 2870 3496 2876 3497
rect 2870 3492 2871 3496
rect 2875 3492 2876 3496
rect 2870 3491 2876 3492
rect 2982 3496 2988 3497
rect 2982 3492 2983 3496
rect 2987 3492 2988 3496
rect 2982 3491 2988 3492
rect 3102 3496 3108 3497
rect 3102 3492 3103 3496
rect 3107 3492 3108 3496
rect 3102 3491 3108 3492
rect 3222 3496 3228 3497
rect 3222 3492 3223 3496
rect 3227 3492 3228 3496
rect 3222 3491 3228 3492
rect 3350 3496 3356 3497
rect 3350 3492 3351 3496
rect 3355 3492 3356 3496
rect 3350 3491 3356 3492
rect 3486 3496 3492 3497
rect 3486 3492 3487 3496
rect 3491 3492 3492 3496
rect 3942 3495 3943 3499
rect 3947 3495 3948 3499
rect 3942 3494 3948 3495
rect 3486 3491 3492 3492
rect 2006 3487 2012 3488
rect 1366 3486 1372 3487
rect 234 3483 240 3484
rect 234 3479 235 3483
rect 239 3479 240 3483
rect 498 3483 504 3484
rect 234 3478 240 3479
rect 362 3479 368 3480
rect 110 3475 116 3476
rect 110 3471 111 3475
rect 115 3471 116 3475
rect 362 3475 363 3479
rect 367 3475 368 3479
rect 498 3479 499 3483
rect 503 3479 504 3483
rect 498 3478 504 3479
rect 634 3483 640 3484
rect 634 3479 635 3483
rect 639 3479 640 3483
rect 634 3478 640 3479
rect 642 3483 648 3484
rect 642 3479 643 3483
rect 647 3482 648 3483
rect 906 3483 912 3484
rect 647 3480 737 3482
rect 647 3479 648 3480
rect 642 3478 648 3479
rect 906 3479 907 3483
rect 911 3479 912 3483
rect 906 3478 912 3479
rect 1042 3483 1048 3484
rect 1042 3479 1043 3483
rect 1047 3479 1048 3483
rect 1042 3478 1048 3479
rect 1170 3483 1176 3484
rect 1170 3479 1171 3483
rect 1175 3479 1176 3483
rect 1170 3478 1176 3479
rect 1306 3483 1312 3484
rect 1306 3479 1307 3483
rect 1311 3479 1312 3483
rect 1306 3478 1312 3479
rect 1338 3483 1344 3484
rect 1338 3479 1339 3483
rect 1343 3482 1344 3483
rect 1343 3480 1409 3482
rect 1343 3479 1344 3480
rect 1338 3478 1344 3479
rect 362 3474 368 3475
rect 2006 3475 2012 3476
rect 110 3470 116 3471
rect 158 3472 164 3473
rect 158 3468 159 3472
rect 163 3468 164 3472
rect 158 3467 164 3468
rect 286 3472 292 3473
rect 286 3468 287 3472
rect 291 3468 292 3472
rect 286 3467 292 3468
rect 422 3472 428 3473
rect 422 3468 423 3472
rect 427 3468 428 3472
rect 422 3467 428 3468
rect 558 3472 564 3473
rect 558 3468 559 3472
rect 563 3468 564 3472
rect 558 3467 564 3468
rect 694 3472 700 3473
rect 694 3468 695 3472
rect 699 3468 700 3472
rect 694 3467 700 3468
rect 830 3472 836 3473
rect 830 3468 831 3472
rect 835 3468 836 3472
rect 830 3467 836 3468
rect 966 3472 972 3473
rect 966 3468 967 3472
rect 971 3468 972 3472
rect 966 3467 972 3468
rect 1094 3472 1100 3473
rect 1094 3468 1095 3472
rect 1099 3468 1100 3472
rect 1094 3467 1100 3468
rect 1230 3472 1236 3473
rect 1230 3468 1231 3472
rect 1235 3468 1236 3472
rect 1230 3467 1236 3468
rect 1366 3472 1372 3473
rect 1366 3468 1367 3472
rect 1371 3468 1372 3472
rect 2006 3471 2007 3475
rect 2011 3471 2012 3475
rect 2006 3470 2012 3471
rect 1366 3467 1372 3468
rect 2486 3436 2492 3437
rect 2046 3433 2052 3434
rect 2046 3429 2047 3433
rect 2051 3429 2052 3433
rect 2486 3432 2487 3436
rect 2491 3432 2492 3436
rect 2486 3431 2492 3432
rect 2582 3436 2588 3437
rect 2582 3432 2583 3436
rect 2587 3432 2588 3436
rect 2582 3431 2588 3432
rect 2678 3436 2684 3437
rect 2678 3432 2679 3436
rect 2683 3432 2684 3436
rect 2678 3431 2684 3432
rect 2782 3436 2788 3437
rect 2782 3432 2783 3436
rect 2787 3432 2788 3436
rect 2782 3431 2788 3432
rect 2894 3436 2900 3437
rect 2894 3432 2895 3436
rect 2899 3432 2900 3436
rect 2894 3431 2900 3432
rect 3014 3436 3020 3437
rect 3014 3432 3015 3436
rect 3019 3432 3020 3436
rect 3014 3431 3020 3432
rect 3142 3436 3148 3437
rect 3142 3432 3143 3436
rect 3147 3432 3148 3436
rect 3142 3431 3148 3432
rect 3270 3436 3276 3437
rect 3270 3432 3271 3436
rect 3275 3432 3276 3436
rect 3270 3431 3276 3432
rect 3406 3436 3412 3437
rect 3406 3432 3407 3436
rect 3411 3432 3412 3436
rect 3406 3431 3412 3432
rect 3942 3433 3948 3434
rect 2046 3428 2052 3429
rect 3942 3429 3943 3433
rect 3947 3429 3948 3433
rect 3942 3428 3948 3429
rect 2562 3427 2568 3428
rect 2562 3423 2563 3427
rect 2567 3423 2568 3427
rect 2562 3422 2568 3423
rect 2658 3427 2664 3428
rect 2658 3423 2659 3427
rect 2663 3423 2664 3427
rect 2658 3422 2664 3423
rect 2746 3427 2752 3428
rect 2746 3423 2747 3427
rect 2751 3423 2752 3427
rect 2746 3422 2752 3423
rect 2775 3427 2781 3428
rect 2775 3423 2776 3427
rect 2780 3426 2781 3427
rect 2886 3427 2892 3428
rect 2780 3424 2825 3426
rect 2780 3423 2781 3424
rect 2775 3422 2781 3423
rect 2886 3423 2887 3427
rect 2891 3426 2892 3427
rect 2990 3427 2996 3428
rect 2891 3424 2937 3426
rect 2891 3423 2892 3424
rect 2886 3422 2892 3423
rect 2990 3423 2991 3427
rect 2995 3426 2996 3427
rect 3230 3427 3236 3428
rect 3230 3426 3231 3427
rect 2995 3424 3057 3426
rect 3221 3424 3231 3426
rect 2995 3423 2996 3424
rect 2990 3422 2996 3423
rect 3230 3423 3231 3424
rect 3235 3423 3236 3427
rect 3230 3422 3236 3423
rect 3338 3427 3344 3428
rect 3338 3423 3339 3427
rect 3343 3423 3344 3427
rect 3338 3422 3344 3423
rect 3378 3427 3384 3428
rect 3378 3423 3379 3427
rect 3383 3426 3384 3427
rect 3383 3424 3449 3426
rect 3383 3423 3384 3424
rect 3378 3422 3384 3423
rect 2486 3417 2492 3418
rect 2046 3416 2052 3417
rect 2046 3412 2047 3416
rect 2051 3412 2052 3416
rect 2486 3413 2487 3417
rect 2491 3413 2492 3417
rect 2486 3412 2492 3413
rect 2582 3417 2588 3418
rect 2582 3413 2583 3417
rect 2587 3413 2588 3417
rect 2582 3412 2588 3413
rect 2678 3417 2684 3418
rect 2678 3413 2679 3417
rect 2683 3413 2684 3417
rect 2678 3412 2684 3413
rect 2782 3417 2788 3418
rect 2782 3413 2783 3417
rect 2787 3413 2788 3417
rect 2782 3412 2788 3413
rect 2894 3417 2900 3418
rect 2894 3413 2895 3417
rect 2899 3413 2900 3417
rect 2894 3412 2900 3413
rect 3014 3417 3020 3418
rect 3014 3413 3015 3417
rect 3019 3413 3020 3417
rect 3014 3412 3020 3413
rect 3142 3417 3148 3418
rect 3142 3413 3143 3417
rect 3147 3413 3148 3417
rect 3142 3412 3148 3413
rect 3270 3417 3276 3418
rect 3270 3413 3271 3417
rect 3275 3413 3276 3417
rect 3270 3412 3276 3413
rect 3406 3417 3412 3418
rect 3406 3413 3407 3417
rect 3411 3413 3412 3417
rect 3406 3412 3412 3413
rect 3942 3416 3948 3417
rect 3942 3412 3943 3416
rect 3947 3412 3948 3416
rect 2046 3411 2052 3412
rect 3942 3411 3948 3412
rect 134 3404 140 3405
rect 110 3401 116 3402
rect 110 3397 111 3401
rect 115 3397 116 3401
rect 134 3400 135 3404
rect 139 3400 140 3404
rect 134 3399 140 3400
rect 246 3404 252 3405
rect 246 3400 247 3404
rect 251 3400 252 3404
rect 246 3399 252 3400
rect 382 3404 388 3405
rect 382 3400 383 3404
rect 387 3400 388 3404
rect 382 3399 388 3400
rect 526 3404 532 3405
rect 526 3400 527 3404
rect 531 3400 532 3404
rect 526 3399 532 3400
rect 670 3404 676 3405
rect 670 3400 671 3404
rect 675 3400 676 3404
rect 670 3399 676 3400
rect 814 3404 820 3405
rect 814 3400 815 3404
rect 819 3400 820 3404
rect 814 3399 820 3400
rect 966 3404 972 3405
rect 966 3400 967 3404
rect 971 3400 972 3404
rect 966 3399 972 3400
rect 1118 3404 1124 3405
rect 1118 3400 1119 3404
rect 1123 3400 1124 3404
rect 1118 3399 1124 3400
rect 1270 3404 1276 3405
rect 1270 3400 1271 3404
rect 1275 3400 1276 3404
rect 1270 3399 1276 3400
rect 2006 3401 2012 3402
rect 110 3396 116 3397
rect 2006 3397 2007 3401
rect 2011 3397 2012 3401
rect 2006 3396 2012 3397
rect 2523 3399 2529 3400
rect 202 3395 208 3396
rect 202 3391 203 3395
rect 207 3391 208 3395
rect 202 3390 208 3391
rect 218 3395 224 3396
rect 218 3391 219 3395
rect 223 3394 224 3395
rect 458 3395 464 3396
rect 223 3392 289 3394
rect 223 3391 224 3392
rect 218 3390 224 3391
rect 458 3391 459 3395
rect 463 3391 464 3395
rect 458 3390 464 3391
rect 602 3395 608 3396
rect 602 3391 603 3395
rect 607 3391 608 3395
rect 602 3390 608 3391
rect 610 3395 616 3396
rect 610 3391 611 3395
rect 615 3394 616 3395
rect 882 3395 888 3396
rect 615 3392 713 3394
rect 615 3391 616 3392
rect 610 3390 616 3391
rect 882 3391 883 3395
rect 887 3391 888 3395
rect 882 3390 888 3391
rect 902 3395 908 3396
rect 902 3391 903 3395
rect 907 3394 908 3395
rect 1194 3395 1200 3396
rect 907 3392 1009 3394
rect 907 3391 908 3392
rect 902 3390 908 3391
rect 1194 3391 1195 3395
rect 1199 3391 1200 3395
rect 1194 3390 1200 3391
rect 1234 3395 1240 3396
rect 1234 3391 1235 3395
rect 1239 3394 1240 3395
rect 2523 3395 2524 3399
rect 2528 3398 2529 3399
rect 2546 3399 2552 3400
rect 2546 3398 2547 3399
rect 2528 3396 2547 3398
rect 2528 3395 2529 3396
rect 2523 3394 2529 3395
rect 2546 3395 2547 3396
rect 2551 3395 2552 3399
rect 2546 3394 2552 3395
rect 2562 3399 2568 3400
rect 2562 3395 2563 3399
rect 2567 3398 2568 3399
rect 2619 3399 2625 3400
rect 2619 3398 2620 3399
rect 2567 3396 2620 3398
rect 2567 3395 2568 3396
rect 2562 3394 2568 3395
rect 2619 3395 2620 3396
rect 2624 3395 2625 3399
rect 2619 3394 2625 3395
rect 2658 3399 2664 3400
rect 2658 3395 2659 3399
rect 2663 3398 2664 3399
rect 2715 3399 2721 3400
rect 2715 3398 2716 3399
rect 2663 3396 2716 3398
rect 2663 3395 2664 3396
rect 2658 3394 2664 3395
rect 2715 3395 2716 3396
rect 2720 3395 2721 3399
rect 2715 3394 2721 3395
rect 2819 3399 2825 3400
rect 2819 3395 2820 3399
rect 2824 3398 2825 3399
rect 2886 3399 2892 3400
rect 2886 3398 2887 3399
rect 2824 3396 2887 3398
rect 2824 3395 2825 3396
rect 2819 3394 2825 3395
rect 2886 3395 2887 3396
rect 2891 3395 2892 3399
rect 2886 3394 2892 3395
rect 2931 3399 2937 3400
rect 2931 3395 2932 3399
rect 2936 3398 2937 3399
rect 2990 3399 2996 3400
rect 2990 3398 2991 3399
rect 2936 3396 2991 3398
rect 2936 3395 2937 3396
rect 2931 3394 2937 3395
rect 2990 3395 2991 3396
rect 2995 3395 2996 3399
rect 2990 3394 2996 3395
rect 3051 3399 3057 3400
rect 3051 3395 3052 3399
rect 3056 3398 3057 3399
rect 3066 3399 3072 3400
rect 3066 3398 3067 3399
rect 3056 3396 3067 3398
rect 3056 3395 3057 3396
rect 3051 3394 3057 3395
rect 3066 3395 3067 3396
rect 3071 3395 3072 3399
rect 3307 3399 3313 3400
rect 3066 3394 3072 3395
rect 3098 3395 3104 3396
rect 1239 3392 1313 3394
rect 1239 3391 1240 3392
rect 1234 3390 1240 3391
rect 3098 3391 3099 3395
rect 3103 3394 3104 3395
rect 3179 3395 3185 3396
rect 3179 3394 3180 3395
rect 3103 3392 3180 3394
rect 3103 3391 3104 3392
rect 3098 3390 3104 3391
rect 3179 3391 3180 3392
rect 3184 3391 3185 3395
rect 3307 3395 3308 3399
rect 3312 3398 3313 3399
rect 3378 3399 3384 3400
rect 3378 3398 3379 3399
rect 3312 3396 3379 3398
rect 3312 3395 3313 3396
rect 3307 3394 3313 3395
rect 3378 3395 3379 3396
rect 3383 3395 3384 3399
rect 3378 3394 3384 3395
rect 3443 3399 3449 3400
rect 3443 3395 3444 3399
rect 3448 3398 3449 3399
rect 3466 3399 3472 3400
rect 3466 3398 3467 3399
rect 3448 3396 3467 3398
rect 3448 3395 3449 3396
rect 3443 3394 3449 3395
rect 3466 3395 3467 3396
rect 3471 3395 3472 3399
rect 3466 3394 3472 3395
rect 3179 3390 3185 3391
rect 134 3385 140 3386
rect 110 3384 116 3385
rect 110 3380 111 3384
rect 115 3380 116 3384
rect 134 3381 135 3385
rect 139 3381 140 3385
rect 134 3380 140 3381
rect 246 3385 252 3386
rect 246 3381 247 3385
rect 251 3381 252 3385
rect 246 3380 252 3381
rect 382 3385 388 3386
rect 382 3381 383 3385
rect 387 3381 388 3385
rect 382 3380 388 3381
rect 526 3385 532 3386
rect 526 3381 527 3385
rect 531 3381 532 3385
rect 526 3380 532 3381
rect 670 3385 676 3386
rect 670 3381 671 3385
rect 675 3381 676 3385
rect 670 3380 676 3381
rect 814 3385 820 3386
rect 814 3381 815 3385
rect 819 3381 820 3385
rect 814 3380 820 3381
rect 966 3385 972 3386
rect 966 3381 967 3385
rect 971 3381 972 3385
rect 966 3380 972 3381
rect 1118 3385 1124 3386
rect 1118 3381 1119 3385
rect 1123 3381 1124 3385
rect 1118 3380 1124 3381
rect 1270 3385 1276 3386
rect 1270 3381 1271 3385
rect 1275 3381 1276 3385
rect 1270 3380 1276 3381
rect 2006 3384 2012 3385
rect 2006 3380 2007 3384
rect 2011 3380 2012 3384
rect 110 3379 116 3380
rect 2006 3379 2012 3380
rect 610 3375 616 3376
rect 610 3374 611 3375
rect 319 3372 611 3374
rect 171 3367 177 3368
rect 171 3363 172 3367
rect 176 3366 177 3367
rect 218 3367 224 3368
rect 218 3366 219 3367
rect 176 3364 219 3366
rect 176 3363 177 3364
rect 171 3362 177 3363
rect 218 3363 219 3364
rect 223 3363 224 3367
rect 218 3362 224 3363
rect 283 3367 289 3368
rect 283 3363 284 3367
rect 288 3366 289 3367
rect 319 3366 321 3372
rect 610 3371 611 3372
rect 615 3371 616 3375
rect 1234 3375 1240 3376
rect 1234 3374 1235 3375
rect 610 3370 616 3371
rect 1159 3372 1235 3374
rect 1159 3370 1161 3372
rect 1234 3371 1235 3372
rect 1239 3371 1240 3375
rect 2426 3375 2432 3376
rect 1234 3370 1240 3371
rect 2387 3373 2393 3374
rect 1080 3368 1161 3370
rect 2387 3369 2388 3373
rect 2392 3369 2393 3373
rect 2426 3371 2427 3375
rect 2431 3374 2432 3375
rect 2515 3375 2521 3376
rect 2515 3374 2516 3375
rect 2431 3372 2516 3374
rect 2431 3371 2432 3372
rect 2426 3370 2432 3371
rect 2515 3371 2516 3372
rect 2520 3371 2521 3375
rect 2515 3370 2521 3371
rect 2554 3375 2560 3376
rect 2554 3371 2555 3375
rect 2559 3374 2560 3375
rect 2651 3375 2657 3376
rect 2651 3374 2652 3375
rect 2559 3372 2652 3374
rect 2559 3371 2560 3372
rect 2554 3370 2560 3371
rect 2651 3371 2652 3372
rect 2656 3371 2657 3375
rect 2651 3370 2657 3371
rect 2775 3375 2781 3376
rect 2775 3371 2776 3375
rect 2780 3374 2781 3375
rect 2787 3375 2793 3376
rect 2787 3374 2788 3375
rect 2780 3372 2788 3374
rect 2780 3371 2781 3372
rect 2775 3370 2781 3371
rect 2787 3371 2788 3372
rect 2792 3371 2793 3375
rect 2787 3370 2793 3371
rect 2850 3375 2856 3376
rect 2850 3371 2851 3375
rect 2855 3374 2856 3375
rect 2923 3375 2929 3376
rect 2923 3374 2924 3375
rect 2855 3372 2924 3374
rect 2855 3371 2856 3372
rect 2850 3370 2856 3371
rect 2923 3371 2924 3372
rect 2928 3371 2929 3375
rect 2923 3370 2929 3371
rect 2962 3375 2968 3376
rect 2962 3371 2963 3375
rect 2967 3374 2968 3375
rect 3059 3375 3065 3376
rect 3059 3374 3060 3375
rect 2967 3372 3060 3374
rect 2967 3371 2968 3372
rect 2962 3370 2968 3371
rect 3059 3371 3060 3372
rect 3064 3371 3065 3375
rect 3059 3370 3065 3371
rect 3195 3375 3201 3376
rect 3195 3371 3196 3375
rect 3200 3374 3201 3375
rect 3242 3375 3248 3376
rect 3242 3374 3243 3375
rect 3200 3372 3243 3374
rect 3200 3371 3201 3372
rect 3195 3370 3201 3371
rect 3242 3371 3243 3372
rect 3247 3371 3248 3375
rect 3242 3370 3248 3371
rect 3338 3375 3345 3376
rect 3338 3371 3339 3375
rect 3344 3371 3345 3375
rect 3338 3370 3345 3371
rect 2387 3368 2393 3369
rect 288 3364 321 3366
rect 362 3367 368 3368
rect 288 3363 289 3364
rect 283 3362 289 3363
rect 362 3363 363 3367
rect 367 3366 368 3367
rect 419 3367 425 3368
rect 419 3366 420 3367
rect 367 3364 420 3366
rect 367 3363 368 3364
rect 362 3362 368 3363
rect 419 3363 420 3364
rect 424 3363 425 3367
rect 419 3362 425 3363
rect 458 3367 464 3368
rect 458 3363 459 3367
rect 463 3366 464 3367
rect 563 3367 569 3368
rect 563 3366 564 3367
rect 463 3364 564 3366
rect 463 3363 464 3364
rect 458 3362 464 3363
rect 563 3363 564 3364
rect 568 3363 569 3367
rect 563 3362 569 3363
rect 602 3367 608 3368
rect 602 3363 603 3367
rect 607 3366 608 3367
rect 707 3367 713 3368
rect 707 3366 708 3367
rect 607 3364 708 3366
rect 607 3363 608 3364
rect 602 3362 608 3363
rect 707 3363 708 3364
rect 712 3363 713 3367
rect 707 3362 713 3363
rect 851 3367 857 3368
rect 851 3363 852 3367
rect 856 3366 857 3367
rect 902 3367 908 3368
rect 902 3366 903 3367
rect 856 3364 903 3366
rect 856 3363 857 3364
rect 851 3362 857 3363
rect 902 3363 903 3364
rect 907 3363 908 3367
rect 902 3362 908 3363
rect 1003 3367 1009 3368
rect 1003 3363 1004 3367
rect 1008 3366 1009 3367
rect 1080 3366 1082 3368
rect 1008 3364 1082 3366
rect 1194 3367 1200 3368
rect 1008 3363 1009 3364
rect 1003 3362 1009 3363
rect 1155 3363 1164 3364
rect 1155 3359 1156 3363
rect 1163 3359 1164 3363
rect 1194 3363 1195 3367
rect 1199 3366 1200 3367
rect 1307 3367 1313 3368
rect 1307 3366 1308 3367
rect 1199 3364 1308 3366
rect 1199 3363 1200 3364
rect 1194 3362 1200 3363
rect 1307 3363 1308 3364
rect 1312 3363 1313 3367
rect 2388 3366 2390 3368
rect 2718 3367 2724 3368
rect 2718 3366 2719 3367
rect 2388 3364 2719 3366
rect 1307 3362 1313 3363
rect 2718 3363 2719 3364
rect 2723 3363 2724 3367
rect 2718 3362 2724 3363
rect 1155 3358 1164 3359
rect 2046 3356 2052 3357
rect 3942 3356 3948 3357
rect 2046 3352 2047 3356
rect 2051 3352 2052 3356
rect 2046 3351 2052 3352
rect 2350 3355 2356 3356
rect 2350 3351 2351 3355
rect 2355 3351 2356 3355
rect 2350 3350 2356 3351
rect 2478 3355 2484 3356
rect 2478 3351 2479 3355
rect 2483 3351 2484 3355
rect 2478 3350 2484 3351
rect 2614 3355 2620 3356
rect 2614 3351 2615 3355
rect 2619 3351 2620 3355
rect 2614 3350 2620 3351
rect 2750 3355 2756 3356
rect 2750 3351 2751 3355
rect 2755 3351 2756 3355
rect 2750 3350 2756 3351
rect 2886 3355 2892 3356
rect 2886 3351 2887 3355
rect 2891 3351 2892 3355
rect 2886 3350 2892 3351
rect 3022 3355 3028 3356
rect 3022 3351 3023 3355
rect 3027 3351 3028 3355
rect 3022 3350 3028 3351
rect 3158 3355 3164 3356
rect 3158 3351 3159 3355
rect 3163 3351 3164 3355
rect 3158 3350 3164 3351
rect 3302 3355 3308 3356
rect 3302 3351 3303 3355
rect 3307 3351 3308 3355
rect 3942 3352 3943 3356
rect 3947 3352 3948 3356
rect 3942 3351 3948 3352
rect 3302 3350 3308 3351
rect 2426 3347 2432 3348
rect 171 3343 177 3344
rect 171 3339 172 3343
rect 176 3342 177 3343
rect 202 3343 208 3344
rect 202 3342 203 3343
rect 176 3340 203 3342
rect 176 3339 177 3340
rect 171 3338 177 3339
rect 202 3339 203 3340
rect 207 3339 208 3343
rect 202 3338 208 3339
rect 210 3343 216 3344
rect 210 3339 211 3343
rect 215 3342 216 3343
rect 299 3343 305 3344
rect 299 3342 300 3343
rect 215 3340 300 3342
rect 215 3339 216 3340
rect 210 3338 216 3339
rect 299 3339 300 3340
rect 304 3339 305 3343
rect 299 3338 305 3339
rect 338 3343 344 3344
rect 338 3339 339 3343
rect 343 3342 344 3343
rect 467 3343 473 3344
rect 467 3342 468 3343
rect 343 3340 468 3342
rect 343 3339 344 3340
rect 338 3338 344 3339
rect 467 3339 468 3340
rect 472 3339 473 3343
rect 467 3338 473 3339
rect 506 3343 512 3344
rect 506 3339 507 3343
rect 511 3342 512 3343
rect 635 3343 641 3344
rect 635 3342 636 3343
rect 511 3340 636 3342
rect 511 3339 512 3340
rect 506 3338 512 3339
rect 635 3339 636 3340
rect 640 3339 641 3343
rect 635 3338 641 3339
rect 719 3343 725 3344
rect 719 3339 720 3343
rect 724 3342 725 3343
rect 803 3343 809 3344
rect 803 3342 804 3343
rect 724 3340 804 3342
rect 724 3339 725 3340
rect 719 3338 725 3339
rect 803 3339 804 3340
rect 808 3339 809 3343
rect 1002 3343 1008 3344
rect 803 3338 809 3339
rect 963 3341 969 3342
rect 963 3337 964 3341
rect 968 3337 969 3341
rect 1002 3339 1003 3343
rect 1007 3342 1008 3343
rect 1123 3343 1129 3344
rect 1123 3342 1124 3343
rect 1007 3340 1124 3342
rect 1007 3339 1008 3340
rect 1002 3338 1008 3339
rect 1123 3339 1124 3340
rect 1128 3339 1129 3343
rect 1123 3338 1129 3339
rect 1275 3343 1281 3344
rect 1275 3339 1276 3343
rect 1280 3342 1281 3343
rect 1322 3343 1328 3344
rect 1322 3342 1323 3343
rect 1280 3340 1323 3342
rect 1280 3339 1281 3340
rect 1275 3338 1281 3339
rect 1322 3339 1323 3340
rect 1327 3339 1328 3343
rect 1322 3338 1328 3339
rect 1427 3343 1433 3344
rect 1427 3339 1428 3343
rect 1432 3342 1433 3343
rect 1474 3343 1480 3344
rect 1474 3342 1475 3343
rect 1432 3340 1475 3342
rect 1432 3339 1433 3340
rect 1427 3338 1433 3339
rect 1474 3339 1475 3340
rect 1479 3339 1480 3343
rect 1474 3338 1480 3339
rect 1562 3343 1568 3344
rect 1562 3339 1563 3343
rect 1567 3342 1568 3343
rect 1587 3343 1593 3344
rect 1587 3342 1588 3343
rect 1567 3340 1588 3342
rect 1567 3339 1568 3340
rect 1562 3338 1568 3339
rect 1587 3339 1588 3340
rect 1592 3339 1593 3343
rect 2426 3343 2427 3347
rect 2431 3343 2432 3347
rect 2426 3342 2432 3343
rect 2554 3347 2560 3348
rect 2554 3343 2555 3347
rect 2559 3343 2560 3347
rect 2554 3342 2560 3343
rect 2718 3347 2724 3348
rect 2718 3343 2719 3347
rect 2723 3346 2724 3347
rect 2962 3347 2968 3348
rect 2723 3344 2793 3346
rect 2723 3343 2724 3344
rect 2718 3342 2724 3343
rect 2962 3343 2963 3347
rect 2967 3343 2968 3347
rect 2962 3342 2968 3343
rect 3098 3347 3104 3348
rect 3098 3343 3099 3347
rect 3103 3343 3104 3347
rect 3242 3347 3248 3348
rect 3098 3342 3104 3343
rect 3234 3343 3240 3344
rect 1587 3338 1593 3339
rect 2046 3339 2052 3340
rect 963 3336 969 3337
rect 964 3334 966 3336
rect 1218 3335 1224 3336
rect 1218 3334 1219 3335
rect 964 3332 1219 3334
rect 1218 3331 1219 3332
rect 1223 3331 1224 3335
rect 2046 3335 2047 3339
rect 2051 3335 2052 3339
rect 2682 3339 2688 3340
rect 2046 3334 2052 3335
rect 2350 3336 2356 3337
rect 2350 3332 2351 3336
rect 2355 3332 2356 3336
rect 2350 3331 2356 3332
rect 2478 3336 2484 3337
rect 2478 3332 2479 3336
rect 2483 3332 2484 3336
rect 2478 3331 2484 3332
rect 2614 3336 2620 3337
rect 2614 3332 2615 3336
rect 2619 3332 2620 3336
rect 2682 3335 2683 3339
rect 2687 3338 2688 3339
rect 2692 3338 2694 3341
rect 3234 3339 3235 3343
rect 3239 3339 3240 3343
rect 3242 3343 3243 3347
rect 3247 3346 3248 3347
rect 3247 3344 3345 3346
rect 3247 3343 3248 3344
rect 3242 3342 3248 3343
rect 3234 3338 3240 3339
rect 3942 3339 3948 3340
rect 2687 3336 2694 3338
rect 2750 3336 2756 3337
rect 2687 3335 2688 3336
rect 2682 3334 2688 3335
rect 2614 3331 2620 3332
rect 2750 3332 2751 3336
rect 2755 3332 2756 3336
rect 2750 3331 2756 3332
rect 2886 3336 2892 3337
rect 2886 3332 2887 3336
rect 2891 3332 2892 3336
rect 2886 3331 2892 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3158 3336 3164 3337
rect 3158 3332 3159 3336
rect 3163 3332 3164 3336
rect 3158 3331 3164 3332
rect 3302 3336 3308 3337
rect 3302 3332 3303 3336
rect 3307 3332 3308 3336
rect 3942 3335 3943 3339
rect 3947 3335 3948 3339
rect 3942 3334 3948 3335
rect 3302 3331 3308 3332
rect 1218 3330 1224 3331
rect 110 3324 116 3325
rect 2006 3324 2012 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 134 3323 140 3324
rect 134 3319 135 3323
rect 139 3319 140 3323
rect 134 3318 140 3319
rect 262 3323 268 3324
rect 262 3319 263 3323
rect 267 3319 268 3323
rect 262 3318 268 3319
rect 430 3323 436 3324
rect 430 3319 431 3323
rect 435 3319 436 3323
rect 430 3318 436 3319
rect 598 3323 604 3324
rect 598 3319 599 3323
rect 603 3319 604 3323
rect 598 3318 604 3319
rect 766 3323 772 3324
rect 766 3319 767 3323
rect 771 3319 772 3323
rect 766 3318 772 3319
rect 926 3323 932 3324
rect 926 3319 927 3323
rect 931 3319 932 3323
rect 926 3318 932 3319
rect 1086 3323 1092 3324
rect 1086 3319 1087 3323
rect 1091 3319 1092 3323
rect 1086 3318 1092 3319
rect 1238 3323 1244 3324
rect 1238 3319 1239 3323
rect 1243 3319 1244 3323
rect 1238 3318 1244 3319
rect 1390 3323 1396 3324
rect 1390 3319 1391 3323
rect 1395 3319 1396 3323
rect 1390 3318 1396 3319
rect 1550 3323 1556 3324
rect 1550 3319 1551 3323
rect 1555 3319 1556 3323
rect 2006 3320 2007 3324
rect 2011 3320 2012 3324
rect 2006 3319 2012 3320
rect 1550 3318 1556 3319
rect 210 3315 216 3316
rect 210 3311 211 3315
rect 215 3311 216 3315
rect 210 3310 216 3311
rect 338 3315 344 3316
rect 338 3311 339 3315
rect 343 3311 344 3315
rect 338 3310 344 3311
rect 506 3315 512 3316
rect 506 3311 507 3315
rect 511 3311 512 3315
rect 719 3315 725 3316
rect 719 3314 720 3315
rect 677 3312 720 3314
rect 506 3310 512 3311
rect 719 3311 720 3312
rect 724 3311 725 3315
rect 719 3310 725 3311
rect 738 3315 744 3316
rect 738 3311 739 3315
rect 743 3314 744 3315
rect 1002 3315 1008 3316
rect 743 3312 809 3314
rect 743 3311 744 3312
rect 738 3310 744 3311
rect 1002 3311 1003 3315
rect 1007 3311 1008 3315
rect 1002 3310 1008 3311
rect 1162 3315 1168 3316
rect 1162 3311 1163 3315
rect 1167 3311 1168 3315
rect 1162 3310 1168 3311
rect 1218 3315 1224 3316
rect 1218 3311 1219 3315
rect 1223 3314 1224 3315
rect 1322 3315 1328 3316
rect 1223 3312 1281 3314
rect 1223 3311 1224 3312
rect 1218 3310 1224 3311
rect 1322 3311 1323 3315
rect 1327 3314 1328 3315
rect 1474 3315 1480 3316
rect 1327 3312 1433 3314
rect 1327 3311 1328 3312
rect 1322 3310 1328 3311
rect 1474 3311 1475 3315
rect 1479 3314 1480 3315
rect 1479 3312 1593 3314
rect 1479 3311 1480 3312
rect 1474 3310 1480 3311
rect 110 3307 116 3308
rect 110 3303 111 3307
rect 115 3303 116 3307
rect 2006 3307 2012 3308
rect 110 3302 116 3303
rect 134 3304 140 3305
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 262 3304 268 3305
rect 262 3300 263 3304
rect 267 3300 268 3304
rect 262 3299 268 3300
rect 430 3304 436 3305
rect 430 3300 431 3304
rect 435 3300 436 3304
rect 430 3299 436 3300
rect 598 3304 604 3305
rect 598 3300 599 3304
rect 603 3300 604 3304
rect 598 3299 604 3300
rect 766 3304 772 3305
rect 766 3300 767 3304
rect 771 3300 772 3304
rect 766 3299 772 3300
rect 926 3304 932 3305
rect 926 3300 927 3304
rect 931 3300 932 3304
rect 926 3299 932 3300
rect 1086 3304 1092 3305
rect 1086 3300 1087 3304
rect 1091 3300 1092 3304
rect 1086 3299 1092 3300
rect 1238 3304 1244 3305
rect 1238 3300 1239 3304
rect 1243 3300 1244 3304
rect 1238 3299 1244 3300
rect 1390 3304 1396 3305
rect 1390 3300 1391 3304
rect 1395 3300 1396 3304
rect 1390 3299 1396 3300
rect 1550 3304 1556 3305
rect 1550 3300 1551 3304
rect 1555 3300 1556 3304
rect 2006 3303 2007 3307
rect 2011 3303 2012 3307
rect 2006 3302 2012 3303
rect 1550 3299 1556 3300
rect 2126 3272 2132 3273
rect 2046 3269 2052 3270
rect 2046 3265 2047 3269
rect 2051 3265 2052 3269
rect 2126 3268 2127 3272
rect 2131 3268 2132 3272
rect 2126 3267 2132 3268
rect 2294 3272 2300 3273
rect 2294 3268 2295 3272
rect 2299 3268 2300 3272
rect 2294 3267 2300 3268
rect 2454 3272 2460 3273
rect 2454 3268 2455 3272
rect 2459 3268 2460 3272
rect 2454 3267 2460 3268
rect 2614 3272 2620 3273
rect 2614 3268 2615 3272
rect 2619 3268 2620 3272
rect 2614 3267 2620 3268
rect 2774 3272 2780 3273
rect 2774 3268 2775 3272
rect 2779 3268 2780 3272
rect 2774 3267 2780 3268
rect 2934 3272 2940 3273
rect 2934 3268 2935 3272
rect 2939 3268 2940 3272
rect 2934 3267 2940 3268
rect 3094 3272 3100 3273
rect 3094 3268 3095 3272
rect 3099 3268 3100 3272
rect 3094 3267 3100 3268
rect 3262 3272 3268 3273
rect 3262 3268 3263 3272
rect 3267 3268 3268 3272
rect 3262 3267 3268 3268
rect 3942 3269 3948 3270
rect 2046 3264 2052 3265
rect 3942 3265 3943 3269
rect 3947 3265 3948 3269
rect 3942 3264 3948 3265
rect 2214 3263 2220 3264
rect 2214 3262 2215 3263
rect 2205 3260 2215 3262
rect 2214 3259 2215 3260
rect 2219 3259 2220 3263
rect 2214 3258 2220 3259
rect 2222 3263 2228 3264
rect 2222 3259 2223 3263
rect 2227 3262 2228 3263
rect 2398 3263 2404 3264
rect 2227 3260 2337 3262
rect 2227 3259 2228 3260
rect 2222 3258 2228 3259
rect 2398 3259 2399 3263
rect 2403 3262 2404 3263
rect 2551 3263 2557 3264
rect 2403 3260 2497 3262
rect 2403 3259 2404 3260
rect 2398 3258 2404 3259
rect 2551 3259 2552 3263
rect 2556 3262 2557 3263
rect 2850 3263 2856 3264
rect 2556 3260 2657 3262
rect 2556 3259 2557 3260
rect 2551 3258 2557 3259
rect 2850 3259 2851 3263
rect 2855 3259 2856 3263
rect 3022 3263 3028 3264
rect 3022 3262 3023 3263
rect 3013 3260 3023 3262
rect 2850 3258 2856 3259
rect 3022 3259 3023 3260
rect 3027 3259 3028 3263
rect 3022 3258 3028 3259
rect 3030 3263 3036 3264
rect 3030 3259 3031 3263
rect 3035 3262 3036 3263
rect 3178 3263 3184 3264
rect 3035 3260 3137 3262
rect 3035 3259 3036 3260
rect 3030 3258 3036 3259
rect 3178 3259 3179 3263
rect 3183 3262 3184 3263
rect 3183 3260 3305 3262
rect 3183 3259 3184 3260
rect 3178 3258 3184 3259
rect 2126 3253 2132 3254
rect 2046 3252 2052 3253
rect 2046 3248 2047 3252
rect 2051 3248 2052 3252
rect 2126 3249 2127 3253
rect 2131 3249 2132 3253
rect 2126 3248 2132 3249
rect 2294 3253 2300 3254
rect 2294 3249 2295 3253
rect 2299 3249 2300 3253
rect 2294 3248 2300 3249
rect 2454 3253 2460 3254
rect 2454 3249 2455 3253
rect 2459 3249 2460 3253
rect 2454 3248 2460 3249
rect 2614 3253 2620 3254
rect 2614 3249 2615 3253
rect 2619 3249 2620 3253
rect 2614 3248 2620 3249
rect 2774 3253 2780 3254
rect 2774 3249 2775 3253
rect 2779 3249 2780 3253
rect 2774 3248 2780 3249
rect 2934 3253 2940 3254
rect 2934 3249 2935 3253
rect 2939 3249 2940 3253
rect 2934 3248 2940 3249
rect 3094 3253 3100 3254
rect 3094 3249 3095 3253
rect 3099 3249 3100 3253
rect 3094 3248 3100 3249
rect 3262 3253 3268 3254
rect 3262 3249 3263 3253
rect 3267 3249 3268 3253
rect 3262 3248 3268 3249
rect 3942 3252 3948 3253
rect 3942 3248 3943 3252
rect 3947 3248 3948 3252
rect 2046 3247 2052 3248
rect 3942 3247 3948 3248
rect 142 3236 148 3237
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 142 3232 143 3236
rect 147 3232 148 3236
rect 142 3231 148 3232
rect 294 3236 300 3237
rect 294 3232 295 3236
rect 299 3232 300 3236
rect 294 3231 300 3232
rect 454 3236 460 3237
rect 454 3232 455 3236
rect 459 3232 460 3236
rect 454 3231 460 3232
rect 622 3236 628 3237
rect 622 3232 623 3236
rect 627 3232 628 3236
rect 622 3231 628 3232
rect 790 3236 796 3237
rect 790 3232 791 3236
rect 795 3232 796 3236
rect 790 3231 796 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 958 3231 964 3232
rect 1126 3236 1132 3237
rect 1126 3232 1127 3236
rect 1131 3232 1132 3236
rect 1126 3231 1132 3232
rect 1302 3236 1308 3237
rect 1302 3232 1303 3236
rect 1307 3232 1308 3236
rect 1302 3231 1308 3232
rect 1478 3236 1484 3237
rect 1478 3232 1479 3236
rect 1483 3232 1484 3236
rect 2163 3235 2169 3236
rect 1478 3231 1484 3232
rect 2006 3233 2012 3234
rect 110 3228 116 3229
rect 2006 3229 2007 3233
rect 2011 3229 2012 3233
rect 2163 3231 2164 3235
rect 2168 3234 2169 3235
rect 2222 3235 2228 3236
rect 2222 3234 2223 3235
rect 2168 3232 2223 3234
rect 2168 3231 2169 3232
rect 2163 3230 2169 3231
rect 2222 3231 2223 3232
rect 2227 3231 2228 3235
rect 2222 3230 2228 3231
rect 2331 3235 2337 3236
rect 2331 3231 2332 3235
rect 2336 3234 2337 3235
rect 2398 3235 2404 3236
rect 2398 3234 2399 3235
rect 2336 3232 2399 3234
rect 2336 3231 2337 3232
rect 2331 3230 2337 3231
rect 2398 3231 2399 3232
rect 2403 3231 2404 3235
rect 2398 3230 2404 3231
rect 2491 3235 2497 3236
rect 2491 3231 2492 3235
rect 2496 3234 2497 3235
rect 2551 3235 2557 3236
rect 2551 3234 2552 3235
rect 2496 3232 2552 3234
rect 2496 3231 2497 3232
rect 2491 3230 2497 3231
rect 2551 3231 2552 3232
rect 2556 3231 2557 3235
rect 2551 3230 2557 3231
rect 2651 3235 2657 3236
rect 2651 3231 2652 3235
rect 2656 3234 2657 3235
rect 2682 3235 2688 3236
rect 2682 3234 2683 3235
rect 2656 3232 2683 3234
rect 2656 3231 2657 3232
rect 2651 3230 2657 3231
rect 2682 3231 2683 3232
rect 2687 3231 2688 3235
rect 2971 3235 2977 3236
rect 2682 3230 2688 3231
rect 2811 3231 2817 3232
rect 2006 3228 2012 3229
rect 218 3227 224 3228
rect 218 3223 219 3227
rect 223 3223 224 3227
rect 218 3222 224 3223
rect 370 3227 376 3228
rect 370 3223 371 3227
rect 375 3223 376 3227
rect 370 3222 376 3223
rect 530 3227 536 3228
rect 530 3223 531 3227
rect 535 3223 536 3227
rect 530 3222 536 3223
rect 698 3227 704 3228
rect 698 3223 699 3227
rect 703 3223 704 3227
rect 698 3222 704 3223
rect 743 3227 749 3228
rect 743 3223 744 3227
rect 748 3226 749 3227
rect 1034 3227 1040 3228
rect 748 3224 833 3226
rect 748 3223 749 3224
rect 743 3222 749 3223
rect 1034 3223 1035 3227
rect 1039 3223 1040 3227
rect 1034 3222 1040 3223
rect 1202 3227 1208 3228
rect 1202 3223 1203 3227
rect 1207 3223 1208 3227
rect 1202 3222 1208 3223
rect 1378 3227 1384 3228
rect 1378 3223 1379 3227
rect 1383 3223 1384 3227
rect 1562 3227 1568 3228
rect 1562 3226 1563 3227
rect 1557 3224 1563 3226
rect 1378 3222 1384 3223
rect 1562 3223 1563 3224
rect 1567 3223 1568 3227
rect 2811 3227 2812 3231
rect 2816 3230 2817 3231
rect 2855 3231 2861 3232
rect 2855 3230 2856 3231
rect 2816 3228 2856 3230
rect 2816 3227 2817 3228
rect 2811 3226 2817 3227
rect 2855 3227 2856 3228
rect 2860 3227 2861 3231
rect 2971 3231 2972 3235
rect 2976 3234 2977 3235
rect 3030 3235 3036 3236
rect 3030 3234 3031 3235
rect 2976 3232 3031 3234
rect 2976 3231 2977 3232
rect 2971 3230 2977 3231
rect 3030 3231 3031 3232
rect 3035 3231 3036 3235
rect 3030 3230 3036 3231
rect 3131 3235 3137 3236
rect 3131 3231 3132 3235
rect 3136 3234 3137 3235
rect 3178 3235 3184 3236
rect 3178 3234 3179 3235
rect 3136 3232 3179 3234
rect 3136 3231 3137 3232
rect 3131 3230 3137 3231
rect 3178 3231 3179 3232
rect 3183 3231 3184 3235
rect 3178 3230 3184 3231
rect 3234 3235 3240 3236
rect 3234 3231 3235 3235
rect 3239 3234 3240 3235
rect 3299 3235 3305 3236
rect 3299 3234 3300 3235
rect 3239 3232 3300 3234
rect 3239 3231 3240 3232
rect 3234 3230 3240 3231
rect 3299 3231 3300 3232
rect 3304 3231 3305 3235
rect 3299 3230 3305 3231
rect 2855 3226 2861 3227
rect 1562 3222 1568 3223
rect 2214 3219 2220 3220
rect 142 3217 148 3218
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 142 3213 143 3217
rect 147 3213 148 3217
rect 142 3212 148 3213
rect 294 3217 300 3218
rect 294 3213 295 3217
rect 299 3213 300 3217
rect 294 3212 300 3213
rect 454 3217 460 3218
rect 454 3213 455 3217
rect 459 3213 460 3217
rect 454 3212 460 3213
rect 622 3217 628 3218
rect 622 3213 623 3217
rect 627 3213 628 3217
rect 622 3212 628 3213
rect 790 3217 796 3218
rect 790 3213 791 3217
rect 795 3213 796 3217
rect 790 3212 796 3213
rect 958 3217 964 3218
rect 958 3213 959 3217
rect 963 3213 964 3217
rect 958 3212 964 3213
rect 1126 3217 1132 3218
rect 1126 3213 1127 3217
rect 1131 3213 1132 3217
rect 1126 3212 1132 3213
rect 1302 3217 1308 3218
rect 1302 3213 1303 3217
rect 1307 3213 1308 3217
rect 1302 3212 1308 3213
rect 1478 3217 1484 3218
rect 2107 3217 2113 3218
rect 1478 3213 1479 3217
rect 1483 3213 1484 3217
rect 1478 3212 1484 3213
rect 2006 3216 2012 3217
rect 2006 3212 2007 3216
rect 2011 3212 2012 3216
rect 2107 3213 2108 3217
rect 2112 3213 2113 3217
rect 2214 3215 2215 3219
rect 2219 3218 2220 3219
rect 2243 3219 2249 3220
rect 2243 3218 2244 3219
rect 2219 3216 2244 3218
rect 2219 3215 2220 3216
rect 2214 3214 2220 3215
rect 2243 3215 2244 3216
rect 2248 3215 2249 3219
rect 2243 3214 2249 3215
rect 2282 3219 2288 3220
rect 2282 3215 2283 3219
rect 2287 3218 2288 3219
rect 2411 3219 2417 3220
rect 2411 3218 2412 3219
rect 2287 3216 2412 3218
rect 2287 3215 2288 3216
rect 2282 3214 2288 3215
rect 2411 3215 2412 3216
rect 2416 3215 2417 3219
rect 2411 3214 2417 3215
rect 2494 3219 2500 3220
rect 2494 3215 2495 3219
rect 2499 3218 2500 3219
rect 2579 3219 2585 3220
rect 2579 3218 2580 3219
rect 2499 3216 2580 3218
rect 2499 3215 2500 3216
rect 2494 3214 2500 3215
rect 2579 3215 2580 3216
rect 2584 3215 2585 3219
rect 2579 3214 2585 3215
rect 2714 3219 2720 3220
rect 2714 3215 2715 3219
rect 2719 3218 2720 3219
rect 2739 3219 2745 3220
rect 2739 3218 2740 3219
rect 2719 3216 2740 3218
rect 2719 3215 2720 3216
rect 2714 3214 2720 3215
rect 2739 3215 2740 3216
rect 2744 3215 2745 3219
rect 2739 3214 2745 3215
rect 2790 3219 2796 3220
rect 2790 3215 2791 3219
rect 2795 3218 2796 3219
rect 2899 3219 2905 3220
rect 2899 3218 2900 3219
rect 2795 3216 2900 3218
rect 2795 3215 2796 3216
rect 2790 3214 2796 3215
rect 2899 3215 2900 3216
rect 2904 3215 2905 3219
rect 2899 3214 2905 3215
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3218 3028 3219
rect 3051 3219 3057 3220
rect 3051 3218 3052 3219
rect 3027 3216 3052 3218
rect 3027 3215 3028 3216
rect 3022 3214 3028 3215
rect 3051 3215 3052 3216
rect 3056 3215 3057 3219
rect 3051 3214 3057 3215
rect 3127 3219 3133 3220
rect 3127 3215 3128 3219
rect 3132 3218 3133 3219
rect 3203 3219 3209 3220
rect 3203 3218 3204 3219
rect 3132 3216 3204 3218
rect 3132 3215 3133 3216
rect 3127 3214 3133 3215
rect 3203 3215 3204 3216
rect 3208 3215 3209 3219
rect 3203 3214 3209 3215
rect 3242 3219 3248 3220
rect 3242 3215 3243 3219
rect 3247 3218 3248 3219
rect 3363 3219 3369 3220
rect 3363 3218 3364 3219
rect 3247 3216 3364 3218
rect 3247 3215 3248 3216
rect 3242 3214 3248 3215
rect 3363 3215 3364 3216
rect 3368 3215 3369 3219
rect 3363 3214 3369 3215
rect 2107 3212 2113 3213
rect 110 3211 116 3212
rect 2006 3211 2012 3212
rect 2108 3210 2110 3212
rect 2502 3211 2508 3212
rect 2502 3210 2503 3211
rect 2108 3208 2503 3210
rect 2502 3207 2503 3208
rect 2507 3207 2508 3211
rect 2502 3206 2508 3207
rect 1034 3203 1040 3204
rect 179 3199 188 3200
rect 179 3195 180 3199
rect 187 3195 188 3199
rect 179 3194 188 3195
rect 218 3199 224 3200
rect 218 3195 219 3199
rect 223 3198 224 3199
rect 331 3199 337 3200
rect 331 3198 332 3199
rect 223 3196 332 3198
rect 223 3195 224 3196
rect 218 3194 224 3195
rect 331 3195 332 3196
rect 336 3195 337 3199
rect 331 3194 337 3195
rect 370 3199 376 3200
rect 370 3195 371 3199
rect 375 3198 376 3199
rect 491 3199 497 3200
rect 491 3198 492 3199
rect 375 3196 492 3198
rect 375 3195 376 3196
rect 370 3194 376 3195
rect 491 3195 492 3196
rect 496 3195 497 3199
rect 491 3194 497 3195
rect 530 3199 536 3200
rect 530 3195 531 3199
rect 535 3198 536 3199
rect 659 3199 665 3200
rect 659 3198 660 3199
rect 535 3196 660 3198
rect 535 3195 536 3196
rect 530 3194 536 3195
rect 659 3195 660 3196
rect 664 3195 665 3199
rect 659 3194 665 3195
rect 698 3199 704 3200
rect 698 3195 699 3199
rect 703 3198 704 3199
rect 827 3199 833 3200
rect 827 3198 828 3199
rect 703 3196 828 3198
rect 703 3195 704 3196
rect 698 3194 704 3195
rect 827 3195 828 3196
rect 832 3195 833 3199
rect 1034 3199 1035 3203
rect 1039 3199 1040 3203
rect 2046 3200 2052 3201
rect 3942 3200 3948 3201
rect 1034 3198 1040 3199
rect 1163 3199 1169 3200
rect 1163 3198 1164 3199
rect 1036 3196 1164 3198
rect 827 3194 833 3195
rect 995 3195 1001 3196
rect 743 3191 749 3192
rect 743 3190 744 3191
rect 332 3188 744 3190
rect 332 3186 334 3188
rect 743 3187 744 3188
rect 748 3187 749 3191
rect 995 3191 996 3195
rect 1000 3194 1001 3195
rect 1163 3195 1164 3196
rect 1168 3195 1169 3199
rect 1163 3194 1169 3195
rect 1202 3199 1208 3200
rect 1202 3195 1203 3199
rect 1207 3198 1208 3199
rect 1339 3199 1345 3200
rect 1339 3198 1340 3199
rect 1207 3196 1340 3198
rect 1207 3195 1208 3196
rect 1202 3194 1208 3195
rect 1339 3195 1340 3196
rect 1344 3195 1345 3199
rect 1339 3194 1345 3195
rect 1378 3199 1384 3200
rect 1378 3195 1379 3199
rect 1383 3198 1384 3199
rect 1515 3199 1521 3200
rect 1515 3198 1516 3199
rect 1383 3196 1516 3198
rect 1383 3195 1384 3196
rect 1378 3194 1384 3195
rect 1515 3195 1516 3196
rect 1520 3195 1521 3199
rect 2046 3196 2047 3200
rect 2051 3196 2052 3200
rect 2046 3195 2052 3196
rect 2070 3199 2076 3200
rect 2070 3195 2071 3199
rect 2075 3195 2076 3199
rect 1515 3194 1521 3195
rect 2070 3194 2076 3195
rect 2206 3199 2212 3200
rect 2206 3195 2207 3199
rect 2211 3195 2212 3199
rect 2206 3194 2212 3195
rect 2374 3199 2380 3200
rect 2374 3195 2375 3199
rect 2379 3195 2380 3199
rect 2374 3194 2380 3195
rect 2542 3199 2548 3200
rect 2542 3195 2543 3199
rect 2547 3195 2548 3199
rect 2542 3194 2548 3195
rect 2702 3199 2708 3200
rect 2702 3195 2703 3199
rect 2707 3195 2708 3199
rect 2702 3194 2708 3195
rect 2862 3199 2868 3200
rect 2862 3195 2863 3199
rect 2867 3195 2868 3199
rect 2862 3194 2868 3195
rect 3014 3199 3020 3200
rect 3014 3195 3015 3199
rect 3019 3195 3020 3199
rect 3014 3194 3020 3195
rect 3166 3199 3172 3200
rect 3166 3195 3167 3199
rect 3171 3195 3172 3199
rect 3166 3194 3172 3195
rect 3326 3199 3332 3200
rect 3326 3195 3327 3199
rect 3331 3195 3332 3199
rect 3942 3196 3943 3200
rect 3947 3196 3948 3200
rect 3942 3195 3948 3196
rect 3326 3194 3332 3195
rect 1000 3192 1161 3194
rect 1000 3191 1001 3192
rect 995 3190 1001 3191
rect 1159 3190 1161 3192
rect 1638 3191 1644 3192
rect 1638 3190 1639 3191
rect 1159 3188 1639 3190
rect 743 3186 749 3187
rect 1638 3187 1639 3188
rect 1643 3187 1644 3191
rect 2282 3191 2288 3192
rect 1638 3186 1644 3187
rect 2146 3187 2152 3188
rect 331 3185 337 3186
rect 331 3181 332 3185
rect 336 3181 337 3185
rect 331 3180 337 3181
rect 370 3183 376 3184
rect 370 3179 371 3183
rect 375 3182 376 3183
rect 467 3183 473 3184
rect 467 3182 468 3183
rect 375 3180 468 3182
rect 375 3179 376 3180
rect 370 3178 376 3179
rect 467 3179 468 3180
rect 472 3179 473 3183
rect 467 3178 473 3179
rect 506 3183 512 3184
rect 506 3179 507 3183
rect 511 3182 512 3183
rect 603 3183 609 3184
rect 603 3182 604 3183
rect 511 3180 604 3182
rect 511 3179 512 3180
rect 506 3178 512 3179
rect 603 3179 604 3180
rect 608 3179 609 3183
rect 603 3178 609 3179
rect 642 3183 648 3184
rect 642 3179 643 3183
rect 647 3182 648 3183
rect 739 3183 745 3184
rect 739 3182 740 3183
rect 647 3180 740 3182
rect 647 3179 648 3180
rect 642 3178 648 3179
rect 739 3179 740 3180
rect 744 3179 745 3183
rect 739 3178 745 3179
rect 891 3183 897 3184
rect 891 3179 892 3183
rect 896 3182 897 3183
rect 922 3183 928 3184
rect 922 3182 923 3183
rect 896 3180 923 3182
rect 896 3179 897 3180
rect 891 3178 897 3179
rect 922 3179 923 3180
rect 927 3179 928 3183
rect 922 3178 928 3179
rect 930 3183 936 3184
rect 930 3179 931 3183
rect 935 3182 936 3183
rect 1067 3183 1073 3184
rect 1067 3182 1068 3183
rect 935 3180 1068 3182
rect 935 3179 936 3180
rect 930 3178 936 3179
rect 1067 3179 1068 3180
rect 1072 3179 1073 3183
rect 1067 3178 1073 3179
rect 1106 3183 1112 3184
rect 1106 3179 1107 3183
rect 1111 3182 1112 3183
rect 1267 3183 1273 3184
rect 1267 3182 1268 3183
rect 1111 3180 1268 3182
rect 1111 3179 1112 3180
rect 1106 3178 1112 3179
rect 1267 3179 1268 3180
rect 1272 3179 1273 3183
rect 1267 3178 1273 3179
rect 1382 3183 1388 3184
rect 1382 3179 1383 3183
rect 1387 3182 1388 3183
rect 1491 3183 1497 3184
rect 1491 3182 1492 3183
rect 1387 3180 1492 3182
rect 1387 3179 1388 3180
rect 1382 3178 1388 3179
rect 1491 3179 1492 3180
rect 1496 3179 1497 3183
rect 1491 3178 1497 3179
rect 1530 3183 1536 3184
rect 1530 3179 1531 3183
rect 1535 3182 1536 3183
rect 1723 3183 1729 3184
rect 1723 3182 1724 3183
rect 1535 3180 1724 3182
rect 1535 3179 1536 3180
rect 1530 3178 1536 3179
rect 1723 3179 1724 3180
rect 1728 3179 1729 3183
rect 1723 3178 1729 3179
rect 1939 3183 1945 3184
rect 1939 3179 1940 3183
rect 1944 3182 1945 3183
rect 1962 3183 1968 3184
rect 1962 3182 1963 3183
rect 1944 3180 1963 3182
rect 1944 3179 1945 3180
rect 1939 3178 1945 3179
rect 1962 3179 1963 3180
rect 1967 3179 1968 3183
rect 1962 3178 1968 3179
rect 2046 3183 2052 3184
rect 2046 3179 2047 3183
rect 2051 3179 2052 3183
rect 2146 3183 2147 3187
rect 2151 3183 2152 3187
rect 2282 3187 2283 3191
rect 2287 3187 2288 3191
rect 2494 3191 2500 3192
rect 2494 3190 2495 3191
rect 2453 3188 2495 3190
rect 2282 3186 2288 3187
rect 2494 3187 2495 3188
rect 2499 3187 2500 3191
rect 2494 3186 2500 3187
rect 2502 3191 2508 3192
rect 2502 3187 2503 3191
rect 2507 3190 2508 3191
rect 2790 3191 2796 3192
rect 2790 3190 2791 3191
rect 2507 3188 2585 3190
rect 2781 3188 2791 3190
rect 2507 3187 2508 3188
rect 2502 3186 2508 3187
rect 2790 3187 2791 3188
rect 2795 3187 2796 3191
rect 2790 3186 2796 3187
rect 2855 3191 2861 3192
rect 2855 3187 2856 3191
rect 2860 3190 2861 3191
rect 3127 3191 3133 3192
rect 3127 3190 3128 3191
rect 2860 3188 2905 3190
rect 3093 3188 3128 3190
rect 2860 3187 2861 3188
rect 2855 3186 2861 3187
rect 3127 3187 3128 3188
rect 3132 3187 3133 3191
rect 3127 3186 3133 3187
rect 3242 3191 3248 3192
rect 3242 3187 3243 3191
rect 3247 3187 3248 3191
rect 3242 3186 3248 3187
rect 3402 3187 3408 3188
rect 2146 3182 2152 3183
rect 3402 3183 3403 3187
rect 3407 3183 3408 3187
rect 3402 3182 3408 3183
rect 3942 3183 3948 3184
rect 2046 3178 2052 3179
rect 2070 3180 2076 3181
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2206 3180 2212 3181
rect 2206 3176 2207 3180
rect 2211 3176 2212 3180
rect 2206 3175 2212 3176
rect 2374 3180 2380 3181
rect 2374 3176 2375 3180
rect 2379 3176 2380 3180
rect 2374 3175 2380 3176
rect 2542 3180 2548 3181
rect 2542 3176 2543 3180
rect 2547 3176 2548 3180
rect 2542 3175 2548 3176
rect 2702 3180 2708 3181
rect 2702 3176 2703 3180
rect 2707 3176 2708 3180
rect 2702 3175 2708 3176
rect 2862 3180 2868 3181
rect 2862 3176 2863 3180
rect 2867 3176 2868 3180
rect 2862 3175 2868 3176
rect 3014 3180 3020 3181
rect 3014 3176 3015 3180
rect 3019 3176 3020 3180
rect 3014 3175 3020 3176
rect 3166 3180 3172 3181
rect 3166 3176 3167 3180
rect 3171 3176 3172 3180
rect 3166 3175 3172 3176
rect 3326 3180 3332 3181
rect 3326 3176 3327 3180
rect 3331 3176 3332 3180
rect 3942 3179 3943 3183
rect 3947 3179 3948 3183
rect 3942 3178 3948 3179
rect 3326 3175 3332 3176
rect 110 3164 116 3165
rect 2006 3164 2012 3165
rect 110 3160 111 3164
rect 115 3160 116 3164
rect 110 3159 116 3160
rect 294 3163 300 3164
rect 294 3159 295 3163
rect 299 3159 300 3163
rect 294 3158 300 3159
rect 430 3163 436 3164
rect 430 3159 431 3163
rect 435 3159 436 3163
rect 430 3158 436 3159
rect 566 3163 572 3164
rect 566 3159 567 3163
rect 571 3159 572 3163
rect 566 3158 572 3159
rect 702 3163 708 3164
rect 702 3159 703 3163
rect 707 3159 708 3163
rect 702 3158 708 3159
rect 854 3163 860 3164
rect 854 3159 855 3163
rect 859 3159 860 3163
rect 854 3158 860 3159
rect 1030 3163 1036 3164
rect 1030 3159 1031 3163
rect 1035 3159 1036 3163
rect 1030 3158 1036 3159
rect 1230 3163 1236 3164
rect 1230 3159 1231 3163
rect 1235 3159 1236 3163
rect 1230 3158 1236 3159
rect 1454 3163 1460 3164
rect 1454 3159 1455 3163
rect 1459 3159 1460 3163
rect 1454 3158 1460 3159
rect 1686 3163 1692 3164
rect 1686 3159 1687 3163
rect 1691 3159 1692 3163
rect 1686 3158 1692 3159
rect 1902 3163 1908 3164
rect 1902 3159 1903 3163
rect 1907 3159 1908 3163
rect 2006 3160 2007 3164
rect 2011 3160 2012 3164
rect 2006 3159 2012 3160
rect 1902 3158 1908 3159
rect 370 3155 376 3156
rect 370 3151 371 3155
rect 375 3151 376 3155
rect 370 3150 376 3151
rect 506 3155 512 3156
rect 506 3151 507 3155
rect 511 3151 512 3155
rect 506 3150 512 3151
rect 642 3155 648 3156
rect 642 3151 643 3155
rect 647 3151 648 3155
rect 642 3150 648 3151
rect 650 3155 656 3156
rect 650 3151 651 3155
rect 655 3154 656 3155
rect 930 3155 936 3156
rect 655 3152 745 3154
rect 655 3151 656 3152
rect 650 3150 656 3151
rect 930 3151 931 3155
rect 935 3151 936 3155
rect 930 3150 936 3151
rect 1106 3155 1112 3156
rect 1106 3151 1107 3155
rect 1111 3151 1112 3155
rect 1382 3155 1388 3156
rect 1382 3154 1383 3155
rect 1309 3152 1383 3154
rect 1106 3150 1112 3151
rect 1382 3151 1383 3152
rect 1387 3151 1388 3155
rect 1382 3150 1388 3151
rect 1530 3155 1536 3156
rect 1530 3151 1531 3155
rect 1535 3151 1536 3155
rect 1530 3150 1536 3151
rect 1638 3155 1644 3156
rect 1638 3151 1639 3155
rect 1643 3154 1644 3155
rect 1643 3152 1729 3154
rect 1643 3151 1644 3152
rect 1638 3150 1644 3151
rect 110 3147 116 3148
rect 110 3143 111 3147
rect 115 3143 116 3147
rect 1970 3147 1976 3148
rect 110 3142 116 3143
rect 294 3144 300 3145
rect 294 3140 295 3144
rect 299 3140 300 3144
rect 294 3139 300 3140
rect 430 3144 436 3145
rect 430 3140 431 3144
rect 435 3140 436 3144
rect 430 3139 436 3140
rect 566 3144 572 3145
rect 566 3140 567 3144
rect 571 3140 572 3144
rect 566 3139 572 3140
rect 702 3144 708 3145
rect 702 3140 703 3144
rect 707 3140 708 3144
rect 702 3139 708 3140
rect 854 3144 860 3145
rect 854 3140 855 3144
rect 859 3140 860 3144
rect 854 3139 860 3140
rect 1030 3144 1036 3145
rect 1030 3140 1031 3144
rect 1035 3140 1036 3144
rect 1030 3139 1036 3140
rect 1230 3144 1236 3145
rect 1230 3140 1231 3144
rect 1235 3140 1236 3144
rect 1230 3139 1236 3140
rect 1454 3144 1460 3145
rect 1454 3140 1455 3144
rect 1459 3140 1460 3144
rect 1454 3139 1460 3140
rect 1686 3144 1692 3145
rect 1686 3140 1687 3144
rect 1691 3140 1692 3144
rect 1686 3139 1692 3140
rect 1902 3144 1908 3145
rect 1902 3140 1903 3144
rect 1907 3140 1908 3144
rect 1970 3143 1971 3147
rect 1975 3146 1976 3147
rect 1980 3146 1982 3149
rect 1975 3144 1982 3146
rect 2006 3147 2012 3148
rect 1975 3143 1976 3144
rect 1970 3142 1976 3143
rect 2006 3143 2007 3147
rect 2011 3143 2012 3147
rect 2006 3142 2012 3143
rect 1902 3139 1908 3140
rect 2070 3116 2076 3117
rect 2046 3113 2052 3114
rect 2046 3109 2047 3113
rect 2051 3109 2052 3113
rect 2070 3112 2071 3116
rect 2075 3112 2076 3116
rect 2070 3111 2076 3112
rect 2342 3116 2348 3117
rect 2342 3112 2343 3116
rect 2347 3112 2348 3116
rect 2342 3111 2348 3112
rect 2630 3116 2636 3117
rect 2630 3112 2631 3116
rect 2635 3112 2636 3116
rect 2630 3111 2636 3112
rect 2902 3116 2908 3117
rect 2902 3112 2903 3116
rect 2907 3112 2908 3116
rect 2902 3111 2908 3112
rect 3174 3116 3180 3117
rect 3174 3112 3175 3116
rect 3179 3112 3180 3116
rect 3174 3111 3180 3112
rect 3446 3116 3452 3117
rect 3446 3112 3447 3116
rect 3451 3112 3452 3116
rect 3446 3111 3452 3112
rect 3942 3113 3948 3114
rect 2046 3108 2052 3109
rect 3942 3109 3943 3113
rect 3947 3109 3948 3113
rect 3942 3108 3948 3109
rect 1962 3107 1968 3108
rect 350 3103 356 3104
rect 350 3099 351 3103
rect 355 3102 356 3103
rect 650 3103 656 3104
rect 650 3102 651 3103
rect 355 3100 651 3102
rect 355 3099 356 3100
rect 350 3098 356 3099
rect 650 3099 651 3100
rect 655 3099 656 3103
rect 1962 3103 1963 3107
rect 1967 3106 1968 3107
rect 2418 3107 2424 3108
rect 1967 3104 2113 3106
rect 1967 3103 1968 3104
rect 1962 3102 1968 3103
rect 2418 3103 2419 3107
rect 2423 3103 2424 3107
rect 2714 3107 2720 3108
rect 2714 3106 2715 3107
rect 2709 3104 2715 3106
rect 2418 3102 2424 3103
rect 2714 3103 2715 3104
rect 2719 3103 2720 3107
rect 2990 3107 2996 3108
rect 2990 3106 2991 3107
rect 2981 3104 2991 3106
rect 2714 3102 2720 3103
rect 2990 3103 2991 3104
rect 2995 3103 2996 3107
rect 2990 3102 2996 3103
rect 3006 3107 3012 3108
rect 3006 3103 3007 3107
rect 3011 3106 3012 3107
rect 3258 3107 3264 3108
rect 3011 3104 3217 3106
rect 3011 3103 3012 3104
rect 3006 3102 3012 3103
rect 3258 3103 3259 3107
rect 3263 3106 3264 3107
rect 3263 3104 3489 3106
rect 3263 3103 3264 3104
rect 3258 3102 3264 3103
rect 650 3098 656 3099
rect 2070 3097 2076 3098
rect 2046 3096 2052 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2070 3093 2071 3097
rect 2075 3093 2076 3097
rect 2070 3092 2076 3093
rect 2342 3097 2348 3098
rect 2342 3093 2343 3097
rect 2347 3093 2348 3097
rect 2342 3092 2348 3093
rect 2630 3097 2636 3098
rect 2630 3093 2631 3097
rect 2635 3093 2636 3097
rect 2630 3092 2636 3093
rect 2902 3097 2908 3098
rect 2902 3093 2903 3097
rect 2907 3093 2908 3097
rect 2902 3092 2908 3093
rect 3174 3097 3180 3098
rect 3174 3093 3175 3097
rect 3179 3093 3180 3097
rect 3174 3092 3180 3093
rect 3446 3097 3452 3098
rect 3446 3093 3447 3097
rect 3451 3093 3452 3097
rect 3446 3092 3452 3093
rect 3942 3096 3948 3097
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 922 3091 928 3092
rect 2046 3091 2052 3092
rect 3942 3091 3948 3092
rect 922 3087 923 3091
rect 927 3090 928 3091
rect 927 3088 1334 3090
rect 927 3087 928 3088
rect 922 3086 928 3087
rect 310 3084 316 3085
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 310 3080 311 3084
rect 315 3080 316 3084
rect 310 3079 316 3080
rect 406 3084 412 3085
rect 406 3080 407 3084
rect 411 3080 412 3084
rect 406 3079 412 3080
rect 502 3084 508 3085
rect 502 3080 503 3084
rect 507 3080 508 3084
rect 502 3079 508 3080
rect 598 3084 604 3085
rect 598 3080 599 3084
rect 603 3080 604 3084
rect 598 3079 604 3080
rect 694 3084 700 3085
rect 694 3080 695 3084
rect 699 3080 700 3084
rect 694 3079 700 3080
rect 806 3084 812 3085
rect 806 3080 807 3084
rect 811 3080 812 3084
rect 806 3079 812 3080
rect 942 3084 948 3085
rect 942 3080 943 3084
rect 947 3080 948 3084
rect 942 3079 948 3080
rect 1086 3084 1092 3085
rect 1086 3080 1087 3084
rect 1091 3080 1092 3084
rect 1086 3079 1092 3080
rect 1246 3084 1252 3085
rect 1246 3080 1247 3084
rect 1251 3080 1252 3084
rect 1246 3079 1252 3080
rect 110 3076 116 3077
rect 386 3075 392 3076
rect 386 3071 387 3075
rect 391 3071 392 3075
rect 386 3070 392 3071
rect 482 3075 488 3076
rect 482 3071 483 3075
rect 487 3071 488 3075
rect 482 3070 488 3071
rect 578 3075 584 3076
rect 578 3071 579 3075
rect 583 3071 584 3075
rect 578 3070 584 3071
rect 674 3075 680 3076
rect 674 3071 675 3075
rect 679 3071 680 3075
rect 674 3070 680 3071
rect 770 3075 776 3076
rect 770 3071 771 3075
rect 775 3071 776 3075
rect 770 3070 776 3071
rect 778 3075 784 3076
rect 778 3071 779 3075
rect 783 3074 784 3075
rect 1018 3075 1024 3076
rect 783 3072 849 3074
rect 783 3071 784 3072
rect 778 3070 784 3071
rect 1018 3071 1019 3075
rect 1023 3071 1024 3075
rect 1018 3070 1024 3071
rect 1162 3075 1168 3076
rect 1162 3071 1163 3075
rect 1167 3071 1168 3075
rect 1162 3070 1168 3071
rect 1322 3075 1328 3076
rect 1322 3071 1323 3075
rect 1327 3071 1328 3075
rect 1332 3074 1334 3088
rect 1406 3084 1412 3085
rect 1406 3080 1407 3084
rect 1411 3080 1412 3084
rect 1406 3079 1412 3080
rect 1574 3084 1580 3085
rect 1574 3080 1575 3084
rect 1579 3080 1580 3084
rect 1574 3079 1580 3080
rect 1750 3084 1756 3085
rect 1750 3080 1751 3084
rect 1755 3080 1756 3084
rect 1750 3079 1756 3080
rect 1902 3084 1908 3085
rect 1902 3080 1903 3084
rect 1907 3080 1908 3084
rect 1902 3079 1908 3080
rect 2006 3081 2012 3082
rect 2006 3077 2007 3081
rect 2011 3077 2012 3081
rect 2006 3076 2012 3077
rect 2107 3079 2113 3080
rect 1650 3075 1656 3076
rect 1332 3072 1449 3074
rect 1322 3070 1328 3071
rect 1650 3071 1651 3075
rect 1655 3071 1656 3075
rect 1650 3070 1656 3071
rect 1826 3075 1832 3076
rect 1826 3071 1827 3075
rect 1831 3071 1832 3075
rect 1826 3070 1832 3071
rect 1834 3075 1840 3076
rect 1834 3071 1835 3075
rect 1839 3074 1840 3075
rect 2107 3075 2108 3079
rect 2112 3078 2113 3079
rect 2146 3079 2152 3080
rect 2146 3078 2147 3079
rect 2112 3076 2147 3078
rect 2112 3075 2113 3076
rect 2107 3074 2113 3075
rect 2146 3075 2147 3076
rect 2151 3075 2152 3079
rect 2418 3079 2424 3080
rect 2146 3074 2152 3075
rect 2379 3075 2385 3076
rect 1839 3072 1945 3074
rect 1839 3071 1840 3072
rect 1834 3070 1840 3071
rect 2379 3071 2380 3075
rect 2384 3074 2385 3075
rect 2418 3075 2419 3079
rect 2423 3078 2424 3079
rect 2667 3079 2673 3080
rect 2667 3078 2668 3079
rect 2423 3076 2668 3078
rect 2423 3075 2424 3076
rect 2418 3074 2424 3075
rect 2667 3075 2668 3076
rect 2672 3075 2673 3079
rect 2667 3074 2673 3075
rect 2939 3079 2945 3080
rect 2939 3075 2940 3079
rect 2944 3078 2945 3079
rect 3006 3079 3012 3080
rect 3006 3078 3007 3079
rect 2944 3076 3007 3078
rect 2944 3075 2945 3076
rect 2939 3074 2945 3075
rect 3006 3075 3007 3076
rect 3011 3075 3012 3079
rect 3006 3074 3012 3075
rect 3211 3079 3217 3080
rect 3211 3075 3212 3079
rect 3216 3078 3217 3079
rect 3258 3079 3264 3080
rect 3258 3078 3259 3079
rect 3216 3076 3259 3078
rect 3216 3075 3217 3076
rect 3211 3074 3217 3075
rect 3258 3075 3259 3076
rect 3263 3075 3264 3079
rect 3258 3074 3264 3075
rect 3402 3079 3408 3080
rect 3402 3075 3403 3079
rect 3407 3078 3408 3079
rect 3483 3079 3489 3080
rect 3483 3078 3484 3079
rect 3407 3076 3484 3078
rect 3407 3075 3408 3076
rect 3402 3074 3408 3075
rect 3483 3075 3484 3076
rect 3488 3075 3489 3079
rect 3483 3074 3489 3075
rect 2384 3072 2414 3074
rect 2384 3071 2385 3072
rect 2379 3070 2385 3071
rect 2412 3070 2414 3072
rect 2826 3071 2832 3072
rect 2826 3070 2827 3071
rect 2412 3068 2827 3070
rect 2826 3067 2827 3068
rect 2831 3067 2832 3071
rect 2826 3066 2832 3067
rect 310 3065 316 3066
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 310 3061 311 3065
rect 315 3061 316 3065
rect 310 3060 316 3061
rect 406 3065 412 3066
rect 406 3061 407 3065
rect 411 3061 412 3065
rect 406 3060 412 3061
rect 502 3065 508 3066
rect 502 3061 503 3065
rect 507 3061 508 3065
rect 502 3060 508 3061
rect 598 3065 604 3066
rect 598 3061 599 3065
rect 603 3061 604 3065
rect 598 3060 604 3061
rect 694 3065 700 3066
rect 694 3061 695 3065
rect 699 3061 700 3065
rect 694 3060 700 3061
rect 806 3065 812 3066
rect 806 3061 807 3065
rect 811 3061 812 3065
rect 806 3060 812 3061
rect 942 3065 948 3066
rect 942 3061 943 3065
rect 947 3061 948 3065
rect 942 3060 948 3061
rect 1086 3065 1092 3066
rect 1086 3061 1087 3065
rect 1091 3061 1092 3065
rect 1086 3060 1092 3061
rect 1246 3065 1252 3066
rect 1246 3061 1247 3065
rect 1251 3061 1252 3065
rect 1246 3060 1252 3061
rect 1406 3065 1412 3066
rect 1406 3061 1407 3065
rect 1411 3061 1412 3065
rect 1406 3060 1412 3061
rect 1574 3065 1580 3066
rect 1574 3061 1575 3065
rect 1579 3061 1580 3065
rect 1574 3060 1580 3061
rect 1750 3065 1756 3066
rect 1750 3061 1751 3065
rect 1755 3061 1756 3065
rect 1750 3060 1756 3061
rect 1902 3065 1908 3066
rect 1902 3061 1903 3065
rect 1907 3061 1908 3065
rect 1902 3060 1908 3061
rect 2006 3064 2012 3065
rect 2006 3060 2007 3064
rect 2011 3060 2012 3064
rect 110 3059 116 3060
rect 2006 3059 2012 3060
rect 2494 3059 2500 3060
rect 1834 3055 1840 3056
rect 1834 3054 1835 3055
rect 1644 3052 1835 3054
rect 347 3047 356 3048
rect 347 3043 348 3047
rect 355 3043 356 3047
rect 347 3042 356 3043
rect 386 3047 392 3048
rect 386 3043 387 3047
rect 391 3046 392 3047
rect 443 3047 449 3048
rect 443 3046 444 3047
rect 391 3044 444 3046
rect 391 3043 392 3044
rect 386 3042 392 3043
rect 443 3043 444 3044
rect 448 3043 449 3047
rect 443 3042 449 3043
rect 482 3047 488 3048
rect 482 3043 483 3047
rect 487 3046 488 3047
rect 539 3047 545 3048
rect 539 3046 540 3047
rect 487 3044 540 3046
rect 487 3043 488 3044
rect 482 3042 488 3043
rect 539 3043 540 3044
rect 544 3043 545 3047
rect 539 3042 545 3043
rect 578 3047 584 3048
rect 578 3043 579 3047
rect 583 3046 584 3047
rect 635 3047 641 3048
rect 635 3046 636 3047
rect 583 3044 636 3046
rect 583 3043 584 3044
rect 578 3042 584 3043
rect 635 3043 636 3044
rect 640 3043 641 3047
rect 635 3042 641 3043
rect 674 3047 680 3048
rect 674 3043 675 3047
rect 679 3046 680 3047
rect 731 3047 737 3048
rect 731 3046 732 3047
rect 679 3044 732 3046
rect 679 3043 680 3044
rect 674 3042 680 3043
rect 731 3043 732 3044
rect 736 3043 737 3047
rect 731 3042 737 3043
rect 770 3047 776 3048
rect 770 3043 771 3047
rect 775 3046 776 3047
rect 843 3047 849 3048
rect 843 3046 844 3047
rect 775 3044 844 3046
rect 775 3043 776 3044
rect 770 3042 776 3043
rect 843 3043 844 3044
rect 848 3043 849 3047
rect 1018 3047 1024 3048
rect 843 3042 849 3043
rect 979 3043 985 3044
rect 979 3039 980 3043
rect 984 3042 985 3043
rect 1018 3043 1019 3047
rect 1023 3046 1024 3047
rect 1123 3047 1129 3048
rect 1123 3046 1124 3047
rect 1023 3044 1124 3046
rect 1023 3043 1024 3044
rect 1018 3042 1024 3043
rect 1123 3043 1124 3044
rect 1128 3043 1129 3047
rect 1123 3042 1129 3043
rect 1162 3047 1168 3048
rect 1162 3043 1163 3047
rect 1167 3046 1168 3047
rect 1283 3047 1289 3048
rect 1283 3046 1284 3047
rect 1167 3044 1284 3046
rect 1167 3043 1168 3044
rect 1162 3042 1168 3043
rect 1283 3043 1284 3044
rect 1288 3043 1289 3047
rect 1283 3042 1289 3043
rect 1322 3047 1328 3048
rect 1322 3043 1323 3047
rect 1327 3046 1328 3047
rect 1443 3047 1449 3048
rect 1443 3046 1444 3047
rect 1327 3044 1444 3046
rect 1327 3043 1328 3044
rect 1322 3042 1328 3043
rect 1443 3043 1444 3044
rect 1448 3043 1449 3047
rect 1443 3042 1449 3043
rect 1611 3047 1617 3048
rect 1611 3043 1612 3047
rect 1616 3046 1617 3047
rect 1644 3046 1646 3052
rect 1834 3051 1835 3052
rect 1839 3051 1840 3055
rect 2494 3055 2495 3059
rect 2499 3058 2500 3059
rect 2523 3059 2529 3060
rect 2523 3058 2524 3059
rect 2499 3056 2524 3058
rect 2499 3055 2500 3056
rect 2494 3054 2500 3055
rect 2523 3055 2524 3056
rect 2528 3055 2529 3059
rect 2523 3054 2529 3055
rect 2562 3059 2568 3060
rect 2562 3055 2563 3059
rect 2567 3058 2568 3059
rect 2651 3059 2657 3060
rect 2651 3058 2652 3059
rect 2567 3056 2652 3058
rect 2567 3055 2568 3056
rect 2562 3054 2568 3055
rect 2651 3055 2652 3056
rect 2656 3055 2657 3059
rect 2651 3054 2657 3055
rect 2690 3059 2696 3060
rect 2690 3055 2691 3059
rect 2695 3058 2696 3059
rect 2779 3059 2785 3060
rect 2779 3058 2780 3059
rect 2695 3056 2780 3058
rect 2695 3055 2696 3056
rect 2690 3054 2696 3055
rect 2779 3055 2780 3056
rect 2784 3055 2785 3059
rect 2779 3054 2785 3055
rect 2818 3059 2824 3060
rect 2818 3055 2819 3059
rect 2823 3058 2824 3059
rect 2899 3059 2905 3060
rect 2899 3058 2900 3059
rect 2823 3056 2900 3058
rect 2823 3055 2824 3056
rect 2818 3054 2824 3055
rect 2899 3055 2900 3056
rect 2904 3055 2905 3059
rect 2899 3054 2905 3055
rect 2990 3059 2996 3060
rect 2990 3055 2991 3059
rect 2995 3058 2996 3059
rect 3019 3059 3025 3060
rect 3019 3058 3020 3059
rect 2995 3056 3020 3058
rect 2995 3055 2996 3056
rect 2990 3054 2996 3055
rect 3019 3055 3020 3056
rect 3024 3055 3025 3059
rect 3019 3054 3025 3055
rect 3058 3059 3064 3060
rect 3058 3055 3059 3059
rect 3063 3058 3064 3059
rect 3139 3059 3145 3060
rect 3139 3058 3140 3059
rect 3063 3056 3140 3058
rect 3063 3055 3064 3056
rect 3058 3054 3064 3055
rect 3139 3055 3140 3056
rect 3144 3055 3145 3059
rect 3139 3054 3145 3055
rect 3198 3059 3204 3060
rect 3198 3055 3199 3059
rect 3203 3058 3204 3059
rect 3251 3059 3257 3060
rect 3251 3058 3252 3059
rect 3203 3056 3252 3058
rect 3203 3055 3204 3056
rect 3198 3054 3204 3055
rect 3251 3055 3252 3056
rect 3256 3055 3257 3059
rect 3251 3054 3257 3055
rect 3290 3059 3296 3060
rect 3290 3055 3291 3059
rect 3295 3058 3296 3059
rect 3363 3059 3369 3060
rect 3363 3058 3364 3059
rect 3295 3056 3364 3058
rect 3295 3055 3296 3056
rect 3290 3054 3296 3055
rect 3363 3055 3364 3056
rect 3368 3055 3369 3059
rect 3363 3054 3369 3055
rect 3402 3059 3408 3060
rect 3402 3055 3403 3059
rect 3407 3058 3408 3059
rect 3467 3059 3473 3060
rect 3467 3058 3468 3059
rect 3407 3056 3468 3058
rect 3407 3055 3408 3056
rect 3402 3054 3408 3055
rect 3467 3055 3468 3056
rect 3472 3055 3473 3059
rect 3467 3054 3473 3055
rect 3571 3059 3577 3060
rect 3571 3055 3572 3059
rect 3576 3058 3577 3059
rect 3602 3059 3608 3060
rect 3602 3058 3603 3059
rect 3576 3056 3603 3058
rect 3576 3055 3577 3056
rect 3571 3054 3577 3055
rect 3602 3055 3603 3056
rect 3607 3055 3608 3059
rect 3602 3054 3608 3055
rect 3610 3059 3616 3060
rect 3610 3055 3611 3059
rect 3615 3058 3616 3059
rect 3675 3059 3681 3060
rect 3675 3058 3676 3059
rect 3615 3056 3676 3058
rect 3615 3055 3616 3056
rect 3610 3054 3616 3055
rect 3675 3055 3676 3056
rect 3680 3055 3681 3059
rect 3675 3054 3681 3055
rect 3714 3059 3720 3060
rect 3714 3055 3715 3059
rect 3719 3058 3720 3059
rect 3779 3059 3785 3060
rect 3779 3058 3780 3059
rect 3719 3056 3780 3058
rect 3719 3055 3720 3056
rect 3714 3054 3720 3055
rect 3779 3055 3780 3056
rect 3784 3055 3785 3059
rect 3779 3054 3785 3055
rect 3818 3059 3824 3060
rect 3818 3055 3819 3059
rect 3823 3058 3824 3059
rect 3875 3059 3881 3060
rect 3875 3058 3876 3059
rect 3823 3056 3876 3058
rect 3823 3055 3824 3056
rect 3818 3054 3824 3055
rect 3875 3055 3876 3056
rect 3880 3055 3881 3059
rect 3875 3054 3881 3055
rect 1834 3050 1840 3051
rect 1616 3044 1646 3046
rect 1650 3047 1656 3048
rect 1616 3043 1617 3044
rect 1611 3042 1617 3043
rect 1650 3043 1651 3047
rect 1655 3046 1656 3047
rect 1787 3047 1793 3048
rect 1787 3046 1788 3047
rect 1655 3044 1788 3046
rect 1655 3043 1656 3044
rect 1650 3042 1656 3043
rect 1787 3043 1788 3044
rect 1792 3043 1793 3047
rect 1787 3042 1793 3043
rect 1939 3047 1945 3048
rect 1939 3043 1940 3047
rect 1944 3046 1945 3047
rect 1970 3047 1976 3048
rect 1970 3046 1971 3047
rect 1944 3044 1971 3046
rect 1944 3043 1945 3044
rect 1939 3042 1945 3043
rect 1970 3043 1971 3044
rect 1975 3043 1976 3047
rect 1970 3042 1976 3043
rect 984 3040 1014 3042
rect 2046 3040 2052 3041
rect 3942 3040 3948 3041
rect 984 3039 985 3040
rect 979 3038 985 3039
rect 1012 3038 1014 3040
rect 1278 3039 1284 3040
rect 1278 3038 1279 3039
rect 1012 3036 1279 3038
rect 1278 3035 1279 3036
rect 1283 3035 1284 3039
rect 2046 3036 2047 3040
rect 2051 3036 2052 3040
rect 2046 3035 2052 3036
rect 2486 3039 2492 3040
rect 2486 3035 2487 3039
rect 2491 3035 2492 3039
rect 1278 3034 1284 3035
rect 2486 3034 2492 3035
rect 2614 3039 2620 3040
rect 2614 3035 2615 3039
rect 2619 3035 2620 3039
rect 2614 3034 2620 3035
rect 2742 3039 2748 3040
rect 2742 3035 2743 3039
rect 2747 3035 2748 3039
rect 2742 3034 2748 3035
rect 2862 3039 2868 3040
rect 2862 3035 2863 3039
rect 2867 3035 2868 3039
rect 2862 3034 2868 3035
rect 2982 3039 2988 3040
rect 2982 3035 2983 3039
rect 2987 3035 2988 3039
rect 2982 3034 2988 3035
rect 3102 3039 3108 3040
rect 3102 3035 3103 3039
rect 3107 3035 3108 3039
rect 3102 3034 3108 3035
rect 3214 3039 3220 3040
rect 3214 3035 3215 3039
rect 3219 3035 3220 3039
rect 3214 3034 3220 3035
rect 3326 3039 3332 3040
rect 3326 3035 3327 3039
rect 3331 3035 3332 3039
rect 3326 3034 3332 3035
rect 3430 3039 3436 3040
rect 3430 3035 3431 3039
rect 3435 3035 3436 3039
rect 3430 3034 3436 3035
rect 3534 3039 3540 3040
rect 3534 3035 3535 3039
rect 3539 3035 3540 3039
rect 3534 3034 3540 3035
rect 3638 3039 3644 3040
rect 3638 3035 3639 3039
rect 3643 3035 3644 3039
rect 3638 3034 3644 3035
rect 3742 3039 3748 3040
rect 3742 3035 3743 3039
rect 3747 3035 3748 3039
rect 3742 3034 3748 3035
rect 3838 3039 3844 3040
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3942 3036 3943 3040
rect 3947 3036 3948 3040
rect 3942 3035 3948 3036
rect 3838 3034 3844 3035
rect 459 3031 468 3032
rect 459 3027 460 3031
rect 467 3027 468 3031
rect 459 3026 468 3027
rect 510 3031 516 3032
rect 510 3027 511 3031
rect 515 3030 516 3031
rect 555 3031 561 3032
rect 555 3030 556 3031
rect 515 3028 556 3030
rect 515 3027 516 3028
rect 510 3026 516 3027
rect 555 3027 556 3028
rect 560 3027 561 3031
rect 555 3026 561 3027
rect 606 3031 612 3032
rect 606 3027 607 3031
rect 611 3030 612 3031
rect 651 3031 657 3032
rect 651 3030 652 3031
rect 611 3028 652 3030
rect 611 3027 612 3028
rect 606 3026 612 3027
rect 651 3027 652 3028
rect 656 3027 657 3031
rect 651 3026 657 3027
rect 702 3031 708 3032
rect 702 3027 703 3031
rect 707 3030 708 3031
rect 747 3031 753 3032
rect 747 3030 748 3031
rect 707 3028 748 3030
rect 707 3027 708 3028
rect 702 3026 708 3027
rect 747 3027 748 3028
rect 752 3027 753 3031
rect 747 3026 753 3027
rect 786 3031 792 3032
rect 786 3027 787 3031
rect 791 3030 792 3031
rect 851 3031 857 3032
rect 851 3030 852 3031
rect 791 3028 852 3030
rect 791 3027 792 3028
rect 786 3026 792 3027
rect 851 3027 852 3028
rect 856 3027 857 3031
rect 851 3026 857 3027
rect 890 3031 896 3032
rect 890 3027 891 3031
rect 895 3030 896 3031
rect 971 3031 977 3032
rect 971 3030 972 3031
rect 895 3028 972 3030
rect 895 3027 896 3028
rect 890 3026 896 3027
rect 971 3027 972 3028
rect 976 3027 977 3031
rect 971 3026 977 3027
rect 1010 3031 1016 3032
rect 1010 3027 1011 3031
rect 1015 3030 1016 3031
rect 1091 3031 1097 3032
rect 1091 3030 1092 3031
rect 1015 3028 1092 3030
rect 1015 3027 1016 3028
rect 1010 3026 1016 3027
rect 1091 3027 1092 3028
rect 1096 3027 1097 3031
rect 1091 3026 1097 3027
rect 1130 3031 1136 3032
rect 1130 3027 1131 3031
rect 1135 3030 1136 3031
rect 1219 3031 1225 3032
rect 1219 3030 1220 3031
rect 1135 3028 1220 3030
rect 1135 3027 1136 3028
rect 1130 3026 1136 3027
rect 1219 3027 1220 3028
rect 1224 3027 1225 3031
rect 1219 3026 1225 3027
rect 1258 3031 1264 3032
rect 1258 3027 1259 3031
rect 1263 3030 1264 3031
rect 1347 3031 1353 3032
rect 1347 3030 1348 3031
rect 1263 3028 1348 3030
rect 1263 3027 1264 3028
rect 1258 3026 1264 3027
rect 1347 3027 1348 3028
rect 1352 3027 1353 3031
rect 1347 3026 1353 3027
rect 1467 3031 1473 3032
rect 1467 3027 1468 3031
rect 1472 3030 1473 3031
rect 1514 3031 1520 3032
rect 1514 3030 1515 3031
rect 1472 3028 1515 3030
rect 1472 3027 1473 3028
rect 1467 3026 1473 3027
rect 1514 3027 1515 3028
rect 1519 3027 1520 3031
rect 1514 3026 1520 3027
rect 1587 3031 1593 3032
rect 1587 3027 1588 3031
rect 1592 3030 1593 3031
rect 1634 3031 1640 3032
rect 1634 3030 1635 3031
rect 1592 3028 1635 3030
rect 1592 3027 1593 3028
rect 1587 3026 1593 3027
rect 1634 3027 1635 3028
rect 1639 3027 1640 3031
rect 1826 3031 1832 3032
rect 1634 3026 1640 3027
rect 1707 3029 1713 3030
rect 1707 3025 1708 3029
rect 1712 3025 1713 3029
rect 1826 3027 1827 3031
rect 1831 3030 1832 3031
rect 1835 3031 1841 3032
rect 1835 3030 1836 3031
rect 1831 3028 1836 3030
rect 1831 3027 1832 3028
rect 1826 3026 1832 3027
rect 1835 3027 1836 3028
rect 1840 3027 1841 3031
rect 1835 3026 1841 3027
rect 1874 3031 1880 3032
rect 1874 3027 1875 3031
rect 1879 3030 1880 3031
rect 1939 3031 1945 3032
rect 1939 3030 1940 3031
rect 1879 3028 1940 3030
rect 1879 3027 1880 3028
rect 1874 3026 1880 3027
rect 1939 3027 1940 3028
rect 1944 3027 1945 3031
rect 1939 3026 1945 3027
rect 2562 3031 2568 3032
rect 2562 3027 2563 3031
rect 2567 3027 2568 3031
rect 2562 3026 2568 3027
rect 2690 3031 2696 3032
rect 2690 3027 2691 3031
rect 2695 3027 2696 3031
rect 2690 3026 2696 3027
rect 2818 3031 2824 3032
rect 2818 3027 2819 3031
rect 2823 3027 2824 3031
rect 2818 3026 2824 3027
rect 2826 3031 2832 3032
rect 2826 3027 2827 3031
rect 2831 3030 2832 3031
rect 3058 3031 3064 3032
rect 2831 3028 2905 3030
rect 2831 3027 2832 3028
rect 2826 3026 2832 3027
rect 3058 3027 3059 3031
rect 3063 3027 3064 3031
rect 3198 3031 3204 3032
rect 3198 3030 3199 3031
rect 3181 3028 3199 3030
rect 3058 3026 3064 3027
rect 3198 3027 3199 3028
rect 3203 3027 3204 3031
rect 3198 3026 3204 3027
rect 3290 3031 3296 3032
rect 3290 3027 3291 3031
rect 3295 3027 3296 3031
rect 3290 3026 3296 3027
rect 3402 3031 3408 3032
rect 3402 3027 3403 3031
rect 3407 3027 3408 3031
rect 3402 3026 3408 3027
rect 3423 3031 3429 3032
rect 3423 3027 3424 3031
rect 3428 3030 3429 3031
rect 3610 3031 3616 3032
rect 3428 3028 3473 3030
rect 3428 3027 3429 3028
rect 3423 3026 3429 3027
rect 3610 3027 3611 3031
rect 3615 3027 3616 3031
rect 3610 3026 3616 3027
rect 3714 3031 3720 3032
rect 3714 3027 3715 3031
rect 3719 3027 3720 3031
rect 3714 3026 3720 3027
rect 3818 3031 3824 3032
rect 3818 3027 3819 3031
rect 3823 3027 3824 3031
rect 3818 3026 3824 3027
rect 1707 3024 1713 3025
rect 1708 3022 1710 3024
rect 1882 3023 1888 3024
rect 1882 3022 1883 3023
rect 1708 3020 1883 3022
rect 1882 3019 1883 3020
rect 1887 3019 1888 3023
rect 1882 3018 1888 3019
rect 2046 3023 2052 3024
rect 2046 3019 2047 3023
rect 2051 3019 2052 3023
rect 3906 3023 3912 3024
rect 2046 3018 2052 3019
rect 2486 3020 2492 3021
rect 2486 3016 2487 3020
rect 2491 3016 2492 3020
rect 2486 3015 2492 3016
rect 2614 3020 2620 3021
rect 2614 3016 2615 3020
rect 2619 3016 2620 3020
rect 2614 3015 2620 3016
rect 2742 3020 2748 3021
rect 2742 3016 2743 3020
rect 2747 3016 2748 3020
rect 2742 3015 2748 3016
rect 2862 3020 2868 3021
rect 2862 3016 2863 3020
rect 2867 3016 2868 3020
rect 2862 3015 2868 3016
rect 2982 3020 2988 3021
rect 2982 3016 2983 3020
rect 2987 3016 2988 3020
rect 2982 3015 2988 3016
rect 3102 3020 3108 3021
rect 3102 3016 3103 3020
rect 3107 3016 3108 3020
rect 3102 3015 3108 3016
rect 3214 3020 3220 3021
rect 3214 3016 3215 3020
rect 3219 3016 3220 3020
rect 3214 3015 3220 3016
rect 3326 3020 3332 3021
rect 3326 3016 3327 3020
rect 3331 3016 3332 3020
rect 3326 3015 3332 3016
rect 3430 3020 3436 3021
rect 3430 3016 3431 3020
rect 3435 3016 3436 3020
rect 3430 3015 3436 3016
rect 3534 3020 3540 3021
rect 3534 3016 3535 3020
rect 3539 3016 3540 3020
rect 3534 3015 3540 3016
rect 3638 3020 3644 3021
rect 3638 3016 3639 3020
rect 3643 3016 3644 3020
rect 3638 3015 3644 3016
rect 3742 3020 3748 3021
rect 3742 3016 3743 3020
rect 3747 3016 3748 3020
rect 3742 3015 3748 3016
rect 3838 3020 3844 3021
rect 3838 3016 3839 3020
rect 3843 3016 3844 3020
rect 3906 3019 3907 3023
rect 3911 3022 3912 3023
rect 3916 3022 3918 3025
rect 3911 3020 3918 3022
rect 3942 3023 3948 3024
rect 3911 3019 3912 3020
rect 3906 3018 3912 3019
rect 3942 3019 3943 3023
rect 3947 3019 3948 3023
rect 3942 3018 3948 3019
rect 3838 3015 3844 3016
rect 110 3012 116 3013
rect 2006 3012 2012 3013
rect 110 3008 111 3012
rect 115 3008 116 3012
rect 110 3007 116 3008
rect 422 3011 428 3012
rect 422 3007 423 3011
rect 427 3007 428 3011
rect 422 3006 428 3007
rect 518 3011 524 3012
rect 518 3007 519 3011
rect 523 3007 524 3011
rect 518 3006 524 3007
rect 614 3011 620 3012
rect 614 3007 615 3011
rect 619 3007 620 3011
rect 614 3006 620 3007
rect 710 3011 716 3012
rect 710 3007 711 3011
rect 715 3007 716 3011
rect 710 3006 716 3007
rect 814 3011 820 3012
rect 814 3007 815 3011
rect 819 3007 820 3011
rect 814 3006 820 3007
rect 934 3011 940 3012
rect 934 3007 935 3011
rect 939 3007 940 3011
rect 934 3006 940 3007
rect 1054 3011 1060 3012
rect 1054 3007 1055 3011
rect 1059 3007 1060 3011
rect 1054 3006 1060 3007
rect 1182 3011 1188 3012
rect 1182 3007 1183 3011
rect 1187 3007 1188 3011
rect 1182 3006 1188 3007
rect 1310 3011 1316 3012
rect 1310 3007 1311 3011
rect 1315 3007 1316 3011
rect 1310 3006 1316 3007
rect 1430 3011 1436 3012
rect 1430 3007 1431 3011
rect 1435 3007 1436 3011
rect 1430 3006 1436 3007
rect 1550 3011 1556 3012
rect 1550 3007 1551 3011
rect 1555 3007 1556 3011
rect 1550 3006 1556 3007
rect 1670 3011 1676 3012
rect 1670 3007 1671 3011
rect 1675 3007 1676 3011
rect 1670 3006 1676 3007
rect 1798 3011 1804 3012
rect 1798 3007 1799 3011
rect 1803 3007 1804 3011
rect 1798 3006 1804 3007
rect 1902 3011 1908 3012
rect 1902 3007 1903 3011
rect 1907 3007 1908 3011
rect 2006 3008 2007 3012
rect 2011 3008 2012 3012
rect 2006 3007 2012 3008
rect 1902 3006 1908 3007
rect 510 3003 516 3004
rect 510 3002 511 3003
rect 501 3000 511 3002
rect 510 2999 511 3000
rect 515 2999 516 3003
rect 606 3003 612 3004
rect 606 3002 607 3003
rect 597 3000 607 3002
rect 510 2998 516 2999
rect 606 2999 607 3000
rect 611 2999 612 3003
rect 702 3003 708 3004
rect 702 3002 703 3003
rect 693 3000 703 3002
rect 606 2998 612 2999
rect 702 2999 703 3000
rect 707 2999 708 3003
rect 702 2998 708 2999
rect 786 3003 792 3004
rect 786 2999 787 3003
rect 791 2999 792 3003
rect 786 2998 792 2999
rect 890 3003 896 3004
rect 890 2999 891 3003
rect 895 2999 896 3003
rect 890 2998 896 2999
rect 1010 3003 1016 3004
rect 1010 2999 1011 3003
rect 1015 2999 1016 3003
rect 1010 2998 1016 2999
rect 1130 3003 1136 3004
rect 1130 2999 1131 3003
rect 1135 2999 1136 3003
rect 1130 2998 1136 2999
rect 1258 3003 1264 3004
rect 1258 2999 1259 3003
rect 1263 2999 1264 3003
rect 1258 2998 1264 2999
rect 1278 3003 1284 3004
rect 1278 2999 1279 3003
rect 1283 3002 1284 3003
rect 1514 3003 1520 3004
rect 1283 3000 1353 3002
rect 1283 2999 1284 3000
rect 1278 2998 1284 2999
rect 1506 2999 1512 3000
rect 110 2995 116 2996
rect 110 2991 111 2995
rect 115 2991 116 2995
rect 1506 2995 1507 2999
rect 1511 2995 1512 2999
rect 1514 2999 1515 3003
rect 1519 3002 1520 3003
rect 1634 3003 1640 3004
rect 1519 3000 1593 3002
rect 1519 2999 1520 3000
rect 1514 2998 1520 2999
rect 1634 2999 1635 3003
rect 1639 3002 1640 3003
rect 1874 3003 1880 3004
rect 1639 3000 1713 3002
rect 1639 2999 1640 3000
rect 1634 2998 1640 2999
rect 1874 2999 1875 3003
rect 1879 2999 1880 3003
rect 1874 2998 1880 2999
rect 1882 3003 1888 3004
rect 1882 2999 1883 3003
rect 1887 3002 1888 3003
rect 1887 3000 1945 3002
rect 1887 2999 1888 3000
rect 1882 2998 1888 2999
rect 1506 2994 1512 2995
rect 2006 2995 2012 2996
rect 110 2990 116 2991
rect 422 2992 428 2993
rect 422 2988 423 2992
rect 427 2988 428 2992
rect 422 2987 428 2988
rect 518 2992 524 2993
rect 518 2988 519 2992
rect 523 2988 524 2992
rect 518 2987 524 2988
rect 614 2992 620 2993
rect 614 2988 615 2992
rect 619 2988 620 2992
rect 614 2987 620 2988
rect 710 2992 716 2993
rect 710 2988 711 2992
rect 715 2988 716 2992
rect 710 2987 716 2988
rect 814 2992 820 2993
rect 814 2988 815 2992
rect 819 2988 820 2992
rect 814 2987 820 2988
rect 934 2992 940 2993
rect 934 2988 935 2992
rect 939 2988 940 2992
rect 934 2987 940 2988
rect 1054 2992 1060 2993
rect 1054 2988 1055 2992
rect 1059 2988 1060 2992
rect 1054 2987 1060 2988
rect 1182 2992 1188 2993
rect 1182 2988 1183 2992
rect 1187 2988 1188 2992
rect 1182 2987 1188 2988
rect 1310 2992 1316 2993
rect 1310 2988 1311 2992
rect 1315 2988 1316 2992
rect 1310 2987 1316 2988
rect 1430 2992 1436 2993
rect 1430 2988 1431 2992
rect 1435 2988 1436 2992
rect 1430 2987 1436 2988
rect 1550 2992 1556 2993
rect 1550 2988 1551 2992
rect 1555 2988 1556 2992
rect 1550 2987 1556 2988
rect 1670 2992 1676 2993
rect 1670 2988 1671 2992
rect 1675 2988 1676 2992
rect 1670 2987 1676 2988
rect 1798 2992 1804 2993
rect 1798 2988 1799 2992
rect 1803 2988 1804 2992
rect 1798 2987 1804 2988
rect 1902 2992 1908 2993
rect 1902 2988 1903 2992
rect 1907 2988 1908 2992
rect 2006 2991 2007 2995
rect 2011 2991 2012 2995
rect 2006 2990 2012 2991
rect 1902 2987 1908 2988
rect 2406 2956 2412 2957
rect 2046 2953 2052 2954
rect 2046 2949 2047 2953
rect 2051 2949 2052 2953
rect 2406 2952 2407 2956
rect 2411 2952 2412 2956
rect 2406 2951 2412 2952
rect 2574 2956 2580 2957
rect 2574 2952 2575 2956
rect 2579 2952 2580 2956
rect 2574 2951 2580 2952
rect 2766 2956 2772 2957
rect 2766 2952 2767 2956
rect 2771 2952 2772 2956
rect 2766 2951 2772 2952
rect 2966 2956 2972 2957
rect 2966 2952 2967 2956
rect 2971 2952 2972 2956
rect 2966 2951 2972 2952
rect 3182 2956 3188 2957
rect 3182 2952 3183 2956
rect 3187 2952 3188 2956
rect 3182 2951 3188 2952
rect 3398 2956 3404 2957
rect 3398 2952 3399 2956
rect 3403 2952 3404 2956
rect 3398 2951 3404 2952
rect 3622 2956 3628 2957
rect 3622 2952 3623 2956
rect 3627 2952 3628 2956
rect 3622 2951 3628 2952
rect 3838 2956 3844 2957
rect 3838 2952 3839 2956
rect 3843 2952 3844 2956
rect 3838 2951 3844 2952
rect 3942 2953 3948 2954
rect 2046 2948 2052 2949
rect 3942 2949 3943 2953
rect 3947 2949 3948 2953
rect 3942 2948 3948 2949
rect 2494 2947 2500 2948
rect 2494 2946 2495 2947
rect 2485 2944 2495 2946
rect 2494 2943 2495 2944
rect 2499 2943 2500 2947
rect 2494 2942 2500 2943
rect 2502 2947 2508 2948
rect 2502 2943 2503 2947
rect 2507 2946 2508 2947
rect 2694 2947 2700 2948
rect 2507 2944 2617 2946
rect 2507 2943 2508 2944
rect 2502 2942 2508 2943
rect 2694 2943 2695 2947
rect 2699 2946 2700 2947
rect 2922 2947 2928 2948
rect 2699 2944 2809 2946
rect 2699 2943 2700 2944
rect 2694 2942 2700 2943
rect 2922 2943 2923 2947
rect 2927 2946 2928 2947
rect 3114 2947 3120 2948
rect 2927 2944 3009 2946
rect 2927 2943 2928 2944
rect 2922 2942 2928 2943
rect 3114 2943 3115 2947
rect 3119 2946 3120 2947
rect 3474 2947 3480 2948
rect 3119 2944 3225 2946
rect 3119 2943 3120 2944
rect 3114 2942 3120 2943
rect 3474 2943 3475 2947
rect 3479 2943 3480 2947
rect 3474 2942 3480 2943
rect 3602 2947 3608 2948
rect 3602 2943 3603 2947
rect 3607 2946 3608 2947
rect 3914 2947 3920 2948
rect 3607 2944 3665 2946
rect 3607 2943 3608 2944
rect 3602 2942 3608 2943
rect 3914 2943 3915 2947
rect 3919 2943 3920 2947
rect 3914 2942 3920 2943
rect 2406 2937 2412 2938
rect 2046 2936 2052 2937
rect 2046 2932 2047 2936
rect 2051 2932 2052 2936
rect 2406 2933 2407 2937
rect 2411 2933 2412 2937
rect 2406 2932 2412 2933
rect 2574 2937 2580 2938
rect 2574 2933 2575 2937
rect 2579 2933 2580 2937
rect 2574 2932 2580 2933
rect 2766 2937 2772 2938
rect 2766 2933 2767 2937
rect 2771 2933 2772 2937
rect 2766 2932 2772 2933
rect 2966 2937 2972 2938
rect 2966 2933 2967 2937
rect 2971 2933 2972 2937
rect 2966 2932 2972 2933
rect 3182 2937 3188 2938
rect 3182 2933 3183 2937
rect 3187 2933 3188 2937
rect 3182 2932 3188 2933
rect 3398 2937 3404 2938
rect 3398 2933 3399 2937
rect 3403 2933 3404 2937
rect 3398 2932 3404 2933
rect 3622 2937 3628 2938
rect 3622 2933 3623 2937
rect 3627 2933 3628 2937
rect 3622 2932 3628 2933
rect 3838 2937 3844 2938
rect 3838 2933 3839 2937
rect 3843 2933 3844 2937
rect 3838 2932 3844 2933
rect 3942 2936 3948 2937
rect 3942 2932 3943 2936
rect 3947 2932 3948 2936
rect 2046 2931 2052 2932
rect 3942 2931 3948 2932
rect 2443 2919 2449 2920
rect 2443 2915 2444 2919
rect 2448 2918 2449 2919
rect 2502 2919 2508 2920
rect 2502 2918 2503 2919
rect 2448 2916 2503 2918
rect 2448 2915 2449 2916
rect 2443 2914 2449 2915
rect 2502 2915 2503 2916
rect 2507 2915 2508 2919
rect 2502 2914 2508 2915
rect 2611 2919 2617 2920
rect 2611 2915 2612 2919
rect 2616 2918 2617 2919
rect 2694 2919 2700 2920
rect 2694 2918 2695 2919
rect 2616 2916 2695 2918
rect 2616 2915 2617 2916
rect 2611 2914 2617 2915
rect 2694 2915 2695 2916
rect 2699 2915 2700 2919
rect 2694 2914 2700 2915
rect 2803 2919 2809 2920
rect 2803 2915 2804 2919
rect 2808 2918 2809 2919
rect 2922 2919 2928 2920
rect 2922 2918 2923 2919
rect 2808 2916 2923 2918
rect 2808 2915 2809 2916
rect 2803 2914 2809 2915
rect 2922 2915 2923 2916
rect 2927 2915 2928 2919
rect 2922 2914 2928 2915
rect 3003 2919 3009 2920
rect 3003 2915 3004 2919
rect 3008 2918 3009 2919
rect 3114 2919 3120 2920
rect 3114 2918 3115 2919
rect 3008 2916 3115 2918
rect 3008 2915 3009 2916
rect 3003 2914 3009 2915
rect 3114 2915 3115 2916
rect 3119 2915 3120 2919
rect 3423 2919 3429 2920
rect 3114 2914 3120 2915
rect 3130 2915 3136 2916
rect 3130 2911 3131 2915
rect 3135 2914 3136 2915
rect 3219 2915 3225 2916
rect 3219 2914 3220 2915
rect 3135 2912 3220 2914
rect 3135 2911 3136 2912
rect 3130 2910 3136 2911
rect 3219 2911 3220 2912
rect 3224 2911 3225 2915
rect 3423 2915 3424 2919
rect 3428 2918 3429 2919
rect 3435 2919 3441 2920
rect 3435 2918 3436 2919
rect 3428 2916 3436 2918
rect 3428 2915 3429 2916
rect 3423 2914 3429 2915
rect 3435 2915 3436 2916
rect 3440 2915 3441 2919
rect 3435 2914 3441 2915
rect 3474 2919 3480 2920
rect 3474 2915 3475 2919
rect 3479 2918 3480 2919
rect 3659 2919 3665 2920
rect 3659 2918 3660 2919
rect 3479 2916 3660 2918
rect 3479 2915 3480 2916
rect 3474 2914 3480 2915
rect 3659 2915 3660 2916
rect 3664 2915 3665 2919
rect 3659 2914 3665 2915
rect 3875 2919 3881 2920
rect 3875 2915 3876 2919
rect 3880 2918 3881 2919
rect 3906 2919 3912 2920
rect 3906 2918 3907 2919
rect 3880 2916 3907 2918
rect 3880 2915 3881 2916
rect 3875 2914 3881 2915
rect 3906 2915 3907 2916
rect 3911 2915 3912 2919
rect 3906 2914 3912 2915
rect 3219 2910 3225 2911
rect 1478 2908 1484 2909
rect 110 2905 116 2906
rect 110 2901 111 2905
rect 115 2901 116 2905
rect 1478 2904 1479 2908
rect 1483 2904 1484 2908
rect 1478 2903 1484 2904
rect 1574 2908 1580 2909
rect 1574 2904 1575 2908
rect 1579 2904 1580 2908
rect 1574 2903 1580 2904
rect 1670 2908 1676 2909
rect 1670 2904 1671 2908
rect 1675 2904 1676 2908
rect 1670 2903 1676 2904
rect 1766 2908 1772 2909
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1862 2908 1868 2909
rect 1862 2904 1863 2908
rect 1867 2904 1868 2908
rect 1862 2903 1868 2904
rect 2006 2905 2012 2906
rect 110 2900 116 2901
rect 2006 2901 2007 2905
rect 2011 2901 2012 2905
rect 2006 2900 2012 2901
rect 1554 2899 1560 2900
rect 1554 2895 1555 2899
rect 1559 2895 1560 2899
rect 1554 2894 1560 2895
rect 1650 2899 1656 2900
rect 1650 2895 1651 2899
rect 1655 2895 1656 2899
rect 1650 2894 1656 2895
rect 1746 2899 1752 2900
rect 1746 2895 1747 2899
rect 1751 2895 1752 2899
rect 1746 2894 1752 2895
rect 1842 2899 1848 2900
rect 1842 2895 1843 2899
rect 1847 2895 1848 2899
rect 1842 2894 1848 2895
rect 1930 2899 1936 2900
rect 1930 2895 1931 2899
rect 1935 2895 1936 2899
rect 1930 2894 1936 2895
rect 1478 2889 1484 2890
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 1478 2885 1479 2889
rect 1483 2885 1484 2889
rect 1478 2884 1484 2885
rect 1574 2889 1580 2890
rect 1574 2885 1575 2889
rect 1579 2885 1580 2889
rect 1574 2884 1580 2885
rect 1670 2889 1676 2890
rect 1670 2885 1671 2889
rect 1675 2885 1676 2889
rect 1670 2884 1676 2885
rect 1766 2889 1772 2890
rect 1766 2885 1767 2889
rect 1771 2885 1772 2889
rect 1766 2884 1772 2885
rect 1862 2889 1868 2890
rect 1862 2885 1863 2889
rect 1867 2885 1868 2889
rect 1862 2884 1868 2885
rect 2006 2888 2012 2889
rect 2006 2884 2007 2888
rect 2011 2884 2012 2888
rect 2626 2887 2632 2888
rect 110 2883 116 2884
rect 2006 2883 2012 2884
rect 2587 2885 2593 2886
rect 2587 2881 2588 2885
rect 2592 2881 2593 2885
rect 2626 2883 2627 2887
rect 2631 2886 2632 2887
rect 2707 2887 2713 2888
rect 2707 2886 2708 2887
rect 2631 2884 2708 2886
rect 2631 2883 2632 2884
rect 2626 2882 2632 2883
rect 2707 2883 2708 2884
rect 2712 2883 2713 2887
rect 2707 2882 2713 2883
rect 2746 2887 2752 2888
rect 2746 2883 2747 2887
rect 2751 2886 2752 2887
rect 2835 2887 2841 2888
rect 2835 2886 2836 2887
rect 2751 2884 2836 2886
rect 2751 2883 2752 2884
rect 2746 2882 2752 2883
rect 2835 2883 2836 2884
rect 2840 2883 2841 2887
rect 2835 2882 2841 2883
rect 2874 2887 2880 2888
rect 2874 2883 2875 2887
rect 2879 2886 2880 2887
rect 2963 2887 2969 2888
rect 2963 2886 2964 2887
rect 2879 2884 2964 2886
rect 2879 2883 2880 2884
rect 2874 2882 2880 2883
rect 2963 2883 2964 2884
rect 2968 2883 2969 2887
rect 2963 2882 2969 2883
rect 3002 2887 3008 2888
rect 3002 2883 3003 2887
rect 3007 2886 3008 2887
rect 3091 2887 3097 2888
rect 3091 2886 3092 2887
rect 3007 2884 3092 2886
rect 3007 2883 3008 2884
rect 3002 2882 3008 2883
rect 3091 2883 3092 2884
rect 3096 2883 3097 2887
rect 3091 2882 3097 2883
rect 3219 2887 3225 2888
rect 3219 2883 3220 2887
rect 3224 2886 3225 2887
rect 3266 2887 3272 2888
rect 3266 2886 3267 2887
rect 3224 2884 3267 2886
rect 3224 2883 3225 2884
rect 3219 2882 3225 2883
rect 3266 2883 3267 2884
rect 3271 2883 3272 2887
rect 3466 2887 3472 2888
rect 3266 2882 3272 2883
rect 3347 2885 3353 2886
rect 2587 2880 2593 2881
rect 3347 2881 3348 2885
rect 3352 2881 3353 2885
rect 3466 2883 3467 2887
rect 3471 2886 3472 2887
rect 3475 2887 3481 2888
rect 3475 2886 3476 2887
rect 3471 2884 3476 2886
rect 3471 2883 3472 2884
rect 3466 2882 3472 2883
rect 3475 2883 3476 2884
rect 3480 2883 3481 2887
rect 3475 2882 3481 2883
rect 3514 2887 3520 2888
rect 3514 2883 3515 2887
rect 3519 2886 3520 2887
rect 3611 2887 3617 2888
rect 3611 2886 3612 2887
rect 3519 2884 3612 2886
rect 3519 2883 3520 2884
rect 3514 2882 3520 2883
rect 3611 2883 3612 2884
rect 3616 2883 3617 2887
rect 3611 2882 3617 2883
rect 3347 2880 3353 2881
rect 2588 2878 2590 2880
rect 2914 2879 2920 2880
rect 2914 2878 2915 2879
rect 2588 2876 2915 2878
rect 2914 2875 2915 2876
rect 2919 2875 2920 2879
rect 3348 2878 3350 2880
rect 3522 2879 3528 2880
rect 3522 2878 3523 2879
rect 3348 2876 3523 2878
rect 2914 2874 2920 2875
rect 3522 2875 3523 2876
rect 3527 2875 3528 2879
rect 3522 2874 3528 2875
rect 1506 2871 1512 2872
rect 1506 2867 1507 2871
rect 1511 2870 1512 2871
rect 1515 2871 1521 2872
rect 1515 2870 1516 2871
rect 1511 2868 1516 2870
rect 1511 2867 1512 2868
rect 1506 2866 1512 2867
rect 1515 2867 1516 2868
rect 1520 2867 1521 2871
rect 1515 2866 1521 2867
rect 1554 2871 1560 2872
rect 1554 2867 1555 2871
rect 1559 2870 1560 2871
rect 1611 2871 1617 2872
rect 1611 2870 1612 2871
rect 1559 2868 1612 2870
rect 1559 2867 1560 2868
rect 1554 2866 1560 2867
rect 1611 2867 1612 2868
rect 1616 2867 1617 2871
rect 1611 2866 1617 2867
rect 1650 2871 1656 2872
rect 1650 2867 1651 2871
rect 1655 2870 1656 2871
rect 1707 2871 1713 2872
rect 1707 2870 1708 2871
rect 1655 2868 1708 2870
rect 1655 2867 1656 2868
rect 1650 2866 1656 2867
rect 1707 2867 1708 2868
rect 1712 2867 1713 2871
rect 1707 2866 1713 2867
rect 1746 2871 1752 2872
rect 1746 2867 1747 2871
rect 1751 2870 1752 2871
rect 1803 2871 1809 2872
rect 1803 2870 1804 2871
rect 1751 2868 1804 2870
rect 1751 2867 1752 2868
rect 1746 2866 1752 2867
rect 1803 2867 1804 2868
rect 1808 2867 1809 2871
rect 1803 2866 1809 2867
rect 1842 2871 1848 2872
rect 1842 2867 1843 2871
rect 1847 2870 1848 2871
rect 1899 2871 1905 2872
rect 1899 2870 1900 2871
rect 1847 2868 1900 2870
rect 1847 2867 1848 2868
rect 1842 2866 1848 2867
rect 1899 2867 1900 2868
rect 1904 2867 1905 2871
rect 1899 2866 1905 2867
rect 2046 2868 2052 2869
rect 3942 2868 3948 2869
rect 2046 2864 2047 2868
rect 2051 2864 2052 2868
rect 2046 2863 2052 2864
rect 2550 2867 2556 2868
rect 2550 2863 2551 2867
rect 2555 2863 2556 2867
rect 2550 2862 2556 2863
rect 2670 2867 2676 2868
rect 2670 2863 2671 2867
rect 2675 2863 2676 2867
rect 2670 2862 2676 2863
rect 2798 2867 2804 2868
rect 2798 2863 2799 2867
rect 2803 2863 2804 2867
rect 2798 2862 2804 2863
rect 2926 2867 2932 2868
rect 2926 2863 2927 2867
rect 2931 2863 2932 2867
rect 2926 2862 2932 2863
rect 3054 2867 3060 2868
rect 3054 2863 3055 2867
rect 3059 2863 3060 2867
rect 3054 2862 3060 2863
rect 3182 2867 3188 2868
rect 3182 2863 3183 2867
rect 3187 2863 3188 2867
rect 3182 2862 3188 2863
rect 3310 2867 3316 2868
rect 3310 2863 3311 2867
rect 3315 2863 3316 2867
rect 3310 2862 3316 2863
rect 3438 2867 3444 2868
rect 3438 2863 3439 2867
rect 3443 2863 3444 2867
rect 3438 2862 3444 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3942 2864 3943 2868
rect 3947 2864 3948 2868
rect 3942 2863 3948 2864
rect 3574 2862 3580 2863
rect 2626 2859 2632 2860
rect 2626 2855 2627 2859
rect 2631 2855 2632 2859
rect 2626 2854 2632 2855
rect 2746 2859 2752 2860
rect 2746 2855 2747 2859
rect 2751 2855 2752 2859
rect 2746 2854 2752 2855
rect 2874 2859 2880 2860
rect 2874 2855 2875 2859
rect 2879 2855 2880 2859
rect 2874 2854 2880 2855
rect 3002 2859 3008 2860
rect 3002 2855 3003 2859
rect 3007 2855 3008 2859
rect 3002 2854 3008 2855
rect 3130 2859 3136 2860
rect 3130 2855 3131 2859
rect 3135 2855 3136 2859
rect 3130 2854 3136 2855
rect 3142 2859 3148 2860
rect 3142 2855 3143 2859
rect 3147 2858 3148 2859
rect 3266 2859 3272 2860
rect 3147 2856 3225 2858
rect 3147 2855 3148 2856
rect 3142 2854 3148 2855
rect 3266 2855 3267 2859
rect 3271 2858 3272 2859
rect 3514 2859 3520 2860
rect 3271 2856 3353 2858
rect 3271 2855 3272 2856
rect 3266 2854 3272 2855
rect 3514 2855 3515 2859
rect 3519 2855 3520 2859
rect 3514 2854 3520 2855
rect 3522 2859 3528 2860
rect 3522 2855 3523 2859
rect 3527 2858 3528 2859
rect 3527 2856 3617 2858
rect 3527 2855 3528 2856
rect 3522 2854 3528 2855
rect 354 2851 360 2852
rect 354 2847 355 2851
rect 359 2850 360 2851
rect 2046 2851 2052 2852
rect 359 2849 489 2850
rect 359 2848 484 2849
rect 359 2847 360 2848
rect 354 2846 360 2847
rect 315 2845 321 2846
rect 315 2841 316 2845
rect 320 2842 321 2845
rect 483 2845 484 2848
rect 488 2845 489 2849
rect 483 2844 489 2845
rect 522 2847 528 2848
rect 438 2843 444 2844
rect 438 2842 439 2843
rect 320 2841 439 2842
rect 315 2840 439 2841
rect 438 2839 439 2840
rect 443 2839 444 2843
rect 522 2843 523 2847
rect 527 2846 528 2847
rect 667 2847 673 2848
rect 667 2846 668 2847
rect 527 2844 668 2846
rect 527 2843 528 2844
rect 522 2842 528 2843
rect 667 2843 668 2844
rect 672 2843 673 2847
rect 667 2842 673 2843
rect 706 2847 712 2848
rect 706 2843 707 2847
rect 711 2846 712 2847
rect 851 2847 857 2848
rect 851 2846 852 2847
rect 711 2844 852 2846
rect 711 2843 712 2844
rect 706 2842 712 2843
rect 851 2843 852 2844
rect 856 2843 857 2847
rect 851 2842 857 2843
rect 890 2847 896 2848
rect 890 2843 891 2847
rect 895 2846 896 2847
rect 1035 2847 1041 2848
rect 1035 2846 1036 2847
rect 895 2844 1036 2846
rect 895 2843 896 2844
rect 890 2842 896 2843
rect 1035 2843 1036 2844
rect 1040 2843 1041 2847
rect 1258 2847 1264 2848
rect 1035 2842 1041 2843
rect 1219 2845 1225 2846
rect 1219 2841 1220 2845
rect 1224 2841 1225 2845
rect 1258 2843 1259 2847
rect 1263 2846 1264 2847
rect 1395 2847 1401 2848
rect 1395 2846 1396 2847
rect 1263 2844 1396 2846
rect 1263 2843 1264 2844
rect 1258 2842 1264 2843
rect 1395 2843 1396 2844
rect 1400 2843 1401 2847
rect 1395 2842 1401 2843
rect 1563 2847 1569 2848
rect 1563 2843 1564 2847
rect 1568 2846 1569 2847
rect 1610 2847 1616 2848
rect 1610 2846 1611 2847
rect 1568 2844 1611 2846
rect 1568 2843 1569 2844
rect 1563 2842 1569 2843
rect 1610 2843 1611 2844
rect 1615 2843 1616 2847
rect 1610 2842 1616 2843
rect 1731 2847 1737 2848
rect 1731 2843 1732 2847
rect 1736 2846 1737 2847
rect 1778 2847 1784 2848
rect 1778 2846 1779 2847
rect 1736 2844 1779 2846
rect 1736 2843 1737 2844
rect 1731 2842 1737 2843
rect 1778 2843 1779 2844
rect 1783 2843 1784 2847
rect 1778 2842 1784 2843
rect 1899 2847 1905 2848
rect 1899 2843 1900 2847
rect 1904 2846 1905 2847
rect 1930 2847 1936 2848
rect 1930 2846 1931 2847
rect 1904 2844 1931 2846
rect 1904 2843 1905 2844
rect 1899 2842 1905 2843
rect 1930 2843 1931 2844
rect 1935 2843 1936 2847
rect 2046 2847 2047 2851
rect 2051 2847 2052 2851
rect 3942 2851 3948 2852
rect 2046 2846 2052 2847
rect 2550 2848 2556 2849
rect 2550 2844 2551 2848
rect 2555 2844 2556 2848
rect 2550 2843 2556 2844
rect 2670 2848 2676 2849
rect 2670 2844 2671 2848
rect 2675 2844 2676 2848
rect 2670 2843 2676 2844
rect 2798 2848 2804 2849
rect 2798 2844 2799 2848
rect 2803 2844 2804 2848
rect 2798 2843 2804 2844
rect 2926 2848 2932 2849
rect 2926 2844 2927 2848
rect 2931 2844 2932 2848
rect 2926 2843 2932 2844
rect 3054 2848 3060 2849
rect 3054 2844 3055 2848
rect 3059 2844 3060 2848
rect 3054 2843 3060 2844
rect 3182 2848 3188 2849
rect 3182 2844 3183 2848
rect 3187 2844 3188 2848
rect 3182 2843 3188 2844
rect 3310 2848 3316 2849
rect 3310 2844 3311 2848
rect 3315 2844 3316 2848
rect 3310 2843 3316 2844
rect 3438 2848 3444 2849
rect 3438 2844 3439 2848
rect 3443 2844 3444 2848
rect 3438 2843 3444 2844
rect 3574 2848 3580 2849
rect 3574 2844 3575 2848
rect 3579 2844 3580 2848
rect 3942 2847 3943 2851
rect 3947 2847 3948 2851
rect 3942 2846 3948 2847
rect 3574 2843 3580 2844
rect 1930 2842 1936 2843
rect 1219 2840 1225 2841
rect 438 2838 444 2839
rect 1220 2838 1222 2840
rect 1458 2839 1464 2840
rect 1458 2838 1459 2839
rect 1220 2836 1459 2838
rect 1458 2835 1459 2836
rect 1463 2835 1464 2839
rect 1458 2834 1464 2835
rect 110 2828 116 2829
rect 2006 2828 2012 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 110 2823 116 2824
rect 278 2827 284 2828
rect 278 2823 279 2827
rect 283 2823 284 2827
rect 278 2822 284 2823
rect 446 2827 452 2828
rect 446 2823 447 2827
rect 451 2823 452 2827
rect 446 2822 452 2823
rect 630 2827 636 2828
rect 630 2823 631 2827
rect 635 2823 636 2827
rect 630 2822 636 2823
rect 814 2827 820 2828
rect 814 2823 815 2827
rect 819 2823 820 2827
rect 814 2822 820 2823
rect 998 2827 1004 2828
rect 998 2823 999 2827
rect 1003 2823 1004 2827
rect 998 2822 1004 2823
rect 1182 2827 1188 2828
rect 1182 2823 1183 2827
rect 1187 2823 1188 2827
rect 1182 2822 1188 2823
rect 1358 2827 1364 2828
rect 1358 2823 1359 2827
rect 1363 2823 1364 2827
rect 1358 2822 1364 2823
rect 1526 2827 1532 2828
rect 1526 2823 1527 2827
rect 1531 2823 1532 2827
rect 1526 2822 1532 2823
rect 1694 2827 1700 2828
rect 1694 2823 1695 2827
rect 1699 2823 1700 2827
rect 1694 2822 1700 2823
rect 1862 2827 1868 2828
rect 1862 2823 1863 2827
rect 1867 2823 1868 2827
rect 2006 2824 2007 2828
rect 2011 2824 2012 2828
rect 2006 2823 2012 2824
rect 1862 2822 1868 2823
rect 354 2819 360 2820
rect 354 2815 355 2819
rect 359 2815 360 2819
rect 354 2814 360 2815
rect 522 2819 528 2820
rect 522 2815 523 2819
rect 527 2815 528 2819
rect 522 2814 528 2815
rect 706 2819 712 2820
rect 706 2815 707 2819
rect 711 2815 712 2819
rect 706 2814 712 2815
rect 890 2819 896 2820
rect 890 2815 891 2819
rect 895 2815 896 2819
rect 890 2814 896 2815
rect 966 2819 972 2820
rect 966 2815 967 2819
rect 971 2818 972 2819
rect 1258 2819 1264 2820
rect 971 2816 1041 2818
rect 971 2815 972 2816
rect 966 2814 972 2815
rect 1258 2815 1259 2819
rect 1263 2815 1264 2819
rect 1458 2819 1464 2820
rect 1258 2814 1264 2815
rect 1434 2815 1440 2816
rect 110 2811 116 2812
rect 110 2807 111 2811
rect 115 2807 116 2811
rect 1434 2811 1435 2815
rect 1439 2811 1440 2815
rect 1458 2815 1459 2819
rect 1463 2818 1464 2819
rect 1610 2819 1616 2820
rect 1463 2816 1569 2818
rect 1463 2815 1464 2816
rect 1458 2814 1464 2815
rect 1610 2815 1611 2819
rect 1615 2818 1616 2819
rect 1778 2819 1784 2820
rect 1615 2816 1737 2818
rect 1615 2815 1616 2816
rect 1610 2814 1616 2815
rect 1778 2815 1779 2819
rect 1783 2818 1784 2819
rect 1783 2816 1905 2818
rect 1783 2815 1784 2816
rect 1778 2814 1784 2815
rect 1434 2810 1440 2811
rect 2006 2811 2012 2812
rect 110 2806 116 2807
rect 278 2808 284 2809
rect 278 2804 279 2808
rect 283 2804 284 2808
rect 278 2803 284 2804
rect 446 2808 452 2809
rect 446 2804 447 2808
rect 451 2804 452 2808
rect 446 2803 452 2804
rect 630 2808 636 2809
rect 630 2804 631 2808
rect 635 2804 636 2808
rect 630 2803 636 2804
rect 814 2808 820 2809
rect 814 2804 815 2808
rect 819 2804 820 2808
rect 814 2803 820 2804
rect 998 2808 1004 2809
rect 998 2804 999 2808
rect 1003 2804 1004 2808
rect 998 2803 1004 2804
rect 1182 2808 1188 2809
rect 1182 2804 1183 2808
rect 1187 2804 1188 2808
rect 1182 2803 1188 2804
rect 1358 2808 1364 2809
rect 1358 2804 1359 2808
rect 1363 2804 1364 2808
rect 1358 2803 1364 2804
rect 1526 2808 1532 2809
rect 1526 2804 1527 2808
rect 1531 2804 1532 2808
rect 1526 2803 1532 2804
rect 1694 2808 1700 2809
rect 1694 2804 1695 2808
rect 1699 2804 1700 2808
rect 1694 2803 1700 2804
rect 1862 2808 1868 2809
rect 1862 2804 1863 2808
rect 1867 2804 1868 2808
rect 2006 2807 2007 2811
rect 2011 2807 2012 2811
rect 2006 2806 2012 2807
rect 1862 2803 1868 2804
rect 2438 2788 2444 2789
rect 2046 2785 2052 2786
rect 2046 2781 2047 2785
rect 2051 2781 2052 2785
rect 2438 2784 2439 2788
rect 2443 2784 2444 2788
rect 2438 2783 2444 2784
rect 2566 2788 2572 2789
rect 2566 2784 2567 2788
rect 2571 2784 2572 2788
rect 2566 2783 2572 2784
rect 2694 2788 2700 2789
rect 2694 2784 2695 2788
rect 2699 2784 2700 2788
rect 2694 2783 2700 2784
rect 2830 2788 2836 2789
rect 2830 2784 2831 2788
rect 2835 2784 2836 2788
rect 2830 2783 2836 2784
rect 2966 2788 2972 2789
rect 2966 2784 2967 2788
rect 2971 2784 2972 2788
rect 2966 2783 2972 2784
rect 3102 2788 3108 2789
rect 3102 2784 3103 2788
rect 3107 2784 3108 2788
rect 3102 2783 3108 2784
rect 3246 2788 3252 2789
rect 3246 2784 3247 2788
rect 3251 2784 3252 2788
rect 3246 2783 3252 2784
rect 3390 2788 3396 2789
rect 3390 2784 3391 2788
rect 3395 2784 3396 2788
rect 3390 2783 3396 2784
rect 3542 2788 3548 2789
rect 3542 2784 3543 2788
rect 3547 2784 3548 2788
rect 3542 2783 3548 2784
rect 3702 2788 3708 2789
rect 3702 2784 3703 2788
rect 3707 2784 3708 2788
rect 3702 2783 3708 2784
rect 3838 2788 3844 2789
rect 3838 2784 3839 2788
rect 3843 2784 3844 2788
rect 3838 2783 3844 2784
rect 3942 2785 3948 2786
rect 2046 2780 2052 2781
rect 3942 2781 3943 2785
rect 3947 2781 3948 2785
rect 3942 2780 3948 2781
rect 2514 2779 2520 2780
rect 2514 2775 2515 2779
rect 2519 2775 2520 2779
rect 2514 2774 2520 2775
rect 2642 2779 2648 2780
rect 2642 2775 2643 2779
rect 2647 2775 2648 2779
rect 2642 2774 2648 2775
rect 2770 2779 2776 2780
rect 2770 2775 2771 2779
rect 2775 2775 2776 2779
rect 2770 2774 2776 2775
rect 2906 2779 2912 2780
rect 2906 2775 2907 2779
rect 2911 2775 2912 2779
rect 2906 2774 2912 2775
rect 2914 2779 2920 2780
rect 2914 2775 2915 2779
rect 2919 2778 2920 2779
rect 3178 2779 3184 2780
rect 2919 2776 3009 2778
rect 2919 2775 2920 2776
rect 2914 2774 2920 2775
rect 3178 2775 3179 2779
rect 3183 2775 3184 2779
rect 3178 2774 3184 2775
rect 3322 2779 3328 2780
rect 3322 2775 3323 2779
rect 3327 2775 3328 2779
rect 3322 2774 3328 2775
rect 3466 2779 3472 2780
rect 3466 2775 3467 2779
rect 3471 2775 3472 2779
rect 3466 2774 3472 2775
rect 3474 2779 3480 2780
rect 3474 2775 3475 2779
rect 3479 2778 3480 2779
rect 3630 2779 3636 2780
rect 3479 2776 3585 2778
rect 3479 2775 3480 2776
rect 3474 2774 3480 2775
rect 3630 2775 3631 2779
rect 3635 2778 3636 2779
rect 3906 2779 3912 2780
rect 3635 2776 3745 2778
rect 3635 2775 3636 2776
rect 3630 2774 3636 2775
rect 3906 2775 3907 2779
rect 3911 2775 3912 2779
rect 3906 2774 3912 2775
rect 2438 2769 2444 2770
rect 2046 2768 2052 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2438 2765 2439 2769
rect 2443 2765 2444 2769
rect 2438 2764 2444 2765
rect 2566 2769 2572 2770
rect 2566 2765 2567 2769
rect 2571 2765 2572 2769
rect 2566 2764 2572 2765
rect 2694 2769 2700 2770
rect 2694 2765 2695 2769
rect 2699 2765 2700 2769
rect 2694 2764 2700 2765
rect 2830 2769 2836 2770
rect 2830 2765 2831 2769
rect 2835 2765 2836 2769
rect 2830 2764 2836 2765
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2966 2764 2972 2765
rect 3102 2769 3108 2770
rect 3102 2765 3103 2769
rect 3107 2765 3108 2769
rect 3102 2764 3108 2765
rect 3246 2769 3252 2770
rect 3246 2765 3247 2769
rect 3251 2765 3252 2769
rect 3246 2764 3252 2765
rect 3390 2769 3396 2770
rect 3390 2765 3391 2769
rect 3395 2765 3396 2769
rect 3390 2764 3396 2765
rect 3542 2769 3548 2770
rect 3542 2765 3543 2769
rect 3547 2765 3548 2769
rect 3542 2764 3548 2765
rect 3702 2769 3708 2770
rect 3702 2765 3703 2769
rect 3707 2765 3708 2769
rect 3702 2764 3708 2765
rect 3838 2769 3844 2770
rect 3838 2765 3839 2769
rect 3843 2765 3844 2769
rect 3838 2764 3844 2765
rect 3942 2768 3948 2769
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 2046 2763 2052 2764
rect 3942 2763 3948 2764
rect 2514 2751 2520 2752
rect 238 2748 244 2749
rect 110 2745 116 2746
rect 110 2741 111 2745
rect 115 2741 116 2745
rect 238 2744 239 2748
rect 243 2744 244 2748
rect 238 2743 244 2744
rect 350 2748 356 2749
rect 350 2744 351 2748
rect 355 2744 356 2748
rect 350 2743 356 2744
rect 470 2748 476 2749
rect 470 2744 471 2748
rect 475 2744 476 2748
rect 470 2743 476 2744
rect 606 2748 612 2749
rect 606 2744 607 2748
rect 611 2744 612 2748
rect 606 2743 612 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 878 2748 884 2749
rect 878 2744 879 2748
rect 883 2744 884 2748
rect 878 2743 884 2744
rect 1014 2748 1020 2749
rect 1014 2744 1015 2748
rect 1019 2744 1020 2748
rect 1014 2743 1020 2744
rect 1150 2748 1156 2749
rect 1150 2744 1151 2748
rect 1155 2744 1156 2748
rect 1150 2743 1156 2744
rect 1286 2748 1292 2749
rect 1286 2744 1287 2748
rect 1291 2744 1292 2748
rect 1286 2743 1292 2744
rect 1422 2748 1428 2749
rect 1422 2744 1423 2748
rect 1427 2744 1428 2748
rect 1422 2743 1428 2744
rect 1566 2748 1572 2749
rect 1566 2744 1567 2748
rect 1571 2744 1572 2748
rect 2475 2747 2481 2748
rect 1566 2743 1572 2744
rect 2006 2745 2012 2746
rect 110 2740 116 2741
rect 2006 2741 2007 2745
rect 2011 2741 2012 2745
rect 2475 2743 2476 2747
rect 2480 2746 2481 2747
rect 2514 2747 2515 2751
rect 2519 2750 2520 2751
rect 2603 2751 2609 2752
rect 2603 2750 2604 2751
rect 2519 2748 2604 2750
rect 2519 2747 2520 2748
rect 2514 2746 2520 2747
rect 2603 2747 2604 2748
rect 2608 2747 2609 2751
rect 2603 2746 2609 2747
rect 2642 2751 2648 2752
rect 2642 2747 2643 2751
rect 2647 2750 2648 2751
rect 2731 2751 2737 2752
rect 2731 2750 2732 2751
rect 2647 2748 2732 2750
rect 2647 2747 2648 2748
rect 2642 2746 2648 2747
rect 2731 2747 2732 2748
rect 2736 2747 2737 2751
rect 2731 2746 2737 2747
rect 2770 2751 2776 2752
rect 2770 2747 2771 2751
rect 2775 2750 2776 2751
rect 2867 2751 2873 2752
rect 2867 2750 2868 2751
rect 2775 2748 2868 2750
rect 2775 2747 2776 2748
rect 2770 2746 2776 2747
rect 2867 2747 2868 2748
rect 2872 2747 2873 2751
rect 2867 2746 2873 2747
rect 2906 2751 2912 2752
rect 2906 2747 2907 2751
rect 2911 2750 2912 2751
rect 3003 2751 3009 2752
rect 3003 2750 3004 2751
rect 2911 2748 3004 2750
rect 2911 2747 2912 2748
rect 2906 2746 2912 2747
rect 3003 2747 3004 2748
rect 3008 2747 3009 2751
rect 3003 2746 3009 2747
rect 3139 2751 3148 2752
rect 3139 2747 3140 2751
rect 3147 2747 3148 2751
rect 3139 2746 3148 2747
rect 3178 2751 3184 2752
rect 3178 2747 3179 2751
rect 3183 2750 3184 2751
rect 3283 2751 3289 2752
rect 3283 2750 3284 2751
rect 3183 2748 3284 2750
rect 3183 2747 3184 2748
rect 3178 2746 3184 2747
rect 3283 2747 3284 2748
rect 3288 2747 3289 2751
rect 3283 2746 3289 2747
rect 3427 2751 3433 2752
rect 3427 2747 3428 2751
rect 3432 2750 3433 2751
rect 3474 2751 3480 2752
rect 3474 2750 3475 2751
rect 3432 2748 3475 2750
rect 3432 2747 3433 2748
rect 3427 2746 3433 2747
rect 3474 2747 3475 2748
rect 3479 2747 3480 2751
rect 3474 2746 3480 2747
rect 3579 2751 3585 2752
rect 3579 2747 3580 2751
rect 3584 2750 3585 2751
rect 3630 2751 3636 2752
rect 3630 2750 3631 2751
rect 3584 2748 3631 2750
rect 3584 2747 3585 2748
rect 3579 2746 3585 2747
rect 3630 2747 3631 2748
rect 3635 2747 3636 2751
rect 3875 2751 3881 2752
rect 3630 2746 3636 2747
rect 3739 2747 3745 2748
rect 2480 2744 2510 2746
rect 2480 2743 2481 2744
rect 2475 2742 2481 2743
rect 2508 2742 2510 2744
rect 2791 2743 2797 2744
rect 2791 2742 2792 2743
rect 2006 2740 2012 2741
rect 2508 2740 2792 2742
rect 314 2739 320 2740
rect 314 2735 315 2739
rect 319 2735 320 2739
rect 314 2734 320 2735
rect 426 2739 432 2740
rect 426 2735 427 2739
rect 431 2735 432 2739
rect 426 2734 432 2735
rect 438 2739 444 2740
rect 438 2735 439 2739
rect 443 2738 444 2739
rect 554 2739 560 2740
rect 443 2736 513 2738
rect 443 2735 444 2736
rect 438 2734 444 2735
rect 554 2735 555 2739
rect 559 2738 560 2739
rect 726 2739 732 2740
rect 559 2736 649 2738
rect 559 2735 560 2736
rect 554 2734 560 2735
rect 726 2735 727 2739
rect 731 2738 732 2739
rect 850 2739 856 2740
rect 731 2736 785 2738
rect 731 2735 732 2736
rect 726 2734 732 2735
rect 850 2735 851 2739
rect 855 2738 856 2739
rect 1090 2739 1096 2740
rect 855 2736 921 2738
rect 855 2735 856 2736
rect 850 2734 856 2735
rect 1090 2735 1091 2739
rect 1095 2735 1096 2739
rect 1238 2739 1244 2740
rect 1238 2738 1239 2739
rect 1229 2736 1239 2738
rect 1090 2734 1096 2735
rect 1238 2735 1239 2736
rect 1243 2735 1244 2739
rect 1238 2734 1244 2735
rect 1246 2739 1252 2740
rect 1246 2735 1247 2739
rect 1251 2738 1252 2739
rect 1498 2739 1504 2740
rect 1251 2736 1329 2738
rect 1251 2735 1252 2736
rect 1246 2734 1252 2735
rect 1498 2735 1499 2739
rect 1503 2735 1504 2739
rect 1498 2734 1504 2735
rect 1506 2739 1512 2740
rect 1506 2735 1507 2739
rect 1511 2738 1512 2739
rect 2791 2739 2792 2740
rect 2796 2739 2797 2743
rect 3739 2743 3740 2747
rect 3744 2746 3745 2747
rect 3762 2747 3768 2748
rect 3762 2746 3763 2747
rect 3744 2744 3763 2746
rect 3744 2743 3745 2744
rect 3739 2742 3745 2743
rect 3762 2743 3763 2744
rect 3767 2743 3768 2747
rect 3875 2747 3876 2751
rect 3880 2750 3881 2751
rect 3914 2751 3920 2752
rect 3914 2750 3915 2751
rect 3880 2748 3915 2750
rect 3880 2747 3881 2748
rect 3875 2746 3881 2747
rect 3914 2747 3915 2748
rect 3919 2747 3920 2751
rect 3914 2746 3920 2747
rect 3762 2742 3768 2743
rect 2791 2738 2797 2739
rect 1511 2736 1609 2738
rect 1511 2735 1512 2736
rect 1506 2734 1512 2735
rect 238 2729 244 2730
rect 110 2728 116 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 238 2725 239 2729
rect 243 2725 244 2729
rect 238 2724 244 2725
rect 350 2729 356 2730
rect 350 2725 351 2729
rect 355 2725 356 2729
rect 350 2724 356 2725
rect 470 2729 476 2730
rect 470 2725 471 2729
rect 475 2725 476 2729
rect 470 2724 476 2725
rect 606 2729 612 2730
rect 606 2725 607 2729
rect 611 2725 612 2729
rect 606 2724 612 2725
rect 742 2729 748 2730
rect 742 2725 743 2729
rect 747 2725 748 2729
rect 742 2724 748 2725
rect 878 2729 884 2730
rect 878 2725 879 2729
rect 883 2725 884 2729
rect 878 2724 884 2725
rect 1014 2729 1020 2730
rect 1014 2725 1015 2729
rect 1019 2725 1020 2729
rect 1014 2724 1020 2725
rect 1150 2729 1156 2730
rect 1150 2725 1151 2729
rect 1155 2725 1156 2729
rect 1150 2724 1156 2725
rect 1286 2729 1292 2730
rect 1286 2725 1287 2729
rect 1291 2725 1292 2729
rect 1286 2724 1292 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1566 2729 1572 2730
rect 1566 2725 1567 2729
rect 1571 2725 1572 2729
rect 1566 2724 1572 2725
rect 2006 2728 2012 2729
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 110 2723 116 2724
rect 2006 2723 2012 2724
rect 2371 2727 2377 2728
rect 2371 2723 2372 2727
rect 2376 2726 2377 2727
rect 2402 2727 2408 2728
rect 2402 2726 2403 2727
rect 2376 2724 2403 2726
rect 2376 2723 2377 2724
rect 2371 2722 2377 2723
rect 2402 2723 2403 2724
rect 2407 2723 2408 2727
rect 2402 2722 2408 2723
rect 2410 2727 2416 2728
rect 2410 2723 2411 2727
rect 2415 2726 2416 2727
rect 2531 2727 2537 2728
rect 2531 2726 2532 2727
rect 2415 2724 2532 2726
rect 2415 2723 2416 2724
rect 2410 2722 2416 2723
rect 2531 2723 2532 2724
rect 2536 2723 2537 2727
rect 2531 2722 2537 2723
rect 2599 2727 2605 2728
rect 2599 2723 2600 2727
rect 2604 2726 2605 2727
rect 2699 2727 2705 2728
rect 2699 2726 2700 2727
rect 2604 2724 2700 2726
rect 2604 2723 2605 2724
rect 2599 2722 2605 2723
rect 2699 2723 2700 2724
rect 2704 2723 2705 2727
rect 2699 2722 2705 2723
rect 2738 2727 2744 2728
rect 2738 2723 2739 2727
rect 2743 2726 2744 2727
rect 2867 2727 2873 2728
rect 2867 2726 2868 2727
rect 2743 2724 2868 2726
rect 2743 2723 2744 2724
rect 2738 2722 2744 2723
rect 2867 2723 2868 2724
rect 2872 2723 2873 2727
rect 3074 2727 3080 2728
rect 2867 2722 2873 2723
rect 3035 2725 3041 2726
rect 3035 2721 3036 2725
rect 3040 2721 3041 2725
rect 3074 2723 3075 2727
rect 3079 2726 3080 2727
rect 3203 2727 3209 2728
rect 3203 2726 3204 2727
rect 3079 2724 3204 2726
rect 3079 2723 3080 2724
rect 3074 2722 3080 2723
rect 3203 2723 3204 2724
rect 3208 2723 3209 2727
rect 3203 2722 3209 2723
rect 3322 2727 3328 2728
rect 3322 2723 3323 2727
rect 3327 2726 3328 2727
rect 3371 2727 3377 2728
rect 3371 2726 3372 2727
rect 3327 2724 3372 2726
rect 3327 2723 3328 2724
rect 3322 2722 3328 2723
rect 3371 2723 3372 2724
rect 3376 2723 3377 2727
rect 3371 2722 3377 2723
rect 3547 2727 3553 2728
rect 3547 2723 3548 2727
rect 3552 2726 3553 2727
rect 3578 2727 3584 2728
rect 3578 2726 3579 2727
rect 3552 2724 3579 2726
rect 3552 2723 3553 2724
rect 3547 2722 3553 2723
rect 3578 2723 3579 2724
rect 3583 2723 3584 2727
rect 3578 2722 3584 2723
rect 3586 2727 3592 2728
rect 3586 2723 3587 2727
rect 3591 2726 3592 2727
rect 3723 2727 3729 2728
rect 3723 2726 3724 2727
rect 3591 2724 3724 2726
rect 3591 2723 3592 2724
rect 3586 2722 3592 2723
rect 3723 2723 3724 2724
rect 3728 2723 3729 2727
rect 3723 2722 3729 2723
rect 3875 2727 3881 2728
rect 3875 2723 3876 2727
rect 3880 2726 3881 2727
rect 3906 2727 3912 2728
rect 3906 2726 3907 2727
rect 3880 2724 3907 2726
rect 3880 2723 3881 2724
rect 3875 2722 3881 2723
rect 3906 2723 3907 2724
rect 3911 2723 3912 2727
rect 3906 2722 3912 2723
rect 3035 2720 3041 2721
rect 1246 2719 1252 2720
rect 1246 2718 1247 2719
rect 1084 2716 1247 2718
rect 314 2711 320 2712
rect 275 2707 281 2708
rect 275 2703 276 2707
rect 280 2706 281 2707
rect 298 2707 304 2708
rect 298 2706 299 2707
rect 280 2704 299 2706
rect 280 2703 281 2704
rect 275 2702 281 2703
rect 298 2703 299 2704
rect 303 2703 304 2707
rect 314 2707 315 2711
rect 319 2710 320 2711
rect 387 2711 393 2712
rect 387 2710 388 2711
rect 319 2708 388 2710
rect 319 2707 320 2708
rect 314 2706 320 2707
rect 387 2707 388 2708
rect 392 2707 393 2711
rect 387 2706 393 2707
rect 426 2711 432 2712
rect 426 2707 427 2711
rect 431 2710 432 2711
rect 507 2711 513 2712
rect 507 2710 508 2711
rect 431 2708 508 2710
rect 431 2707 432 2708
rect 426 2706 432 2707
rect 507 2707 508 2708
rect 512 2707 513 2711
rect 507 2706 513 2707
rect 643 2711 649 2712
rect 643 2707 644 2711
rect 648 2710 649 2711
rect 726 2711 732 2712
rect 726 2710 727 2711
rect 648 2708 727 2710
rect 648 2707 649 2708
rect 643 2706 649 2707
rect 726 2707 727 2708
rect 731 2707 732 2711
rect 726 2706 732 2707
rect 779 2711 785 2712
rect 779 2707 780 2711
rect 784 2710 785 2711
rect 850 2711 856 2712
rect 850 2710 851 2711
rect 784 2708 851 2710
rect 784 2707 785 2708
rect 779 2706 785 2707
rect 850 2707 851 2708
rect 855 2707 856 2711
rect 850 2706 856 2707
rect 915 2711 921 2712
rect 915 2707 916 2711
rect 920 2710 921 2711
rect 966 2711 972 2712
rect 966 2710 967 2711
rect 920 2708 967 2710
rect 920 2707 921 2708
rect 915 2706 921 2707
rect 966 2707 967 2708
rect 971 2707 972 2711
rect 966 2706 972 2707
rect 1051 2711 1057 2712
rect 1051 2707 1052 2711
rect 1056 2710 1057 2711
rect 1084 2710 1086 2716
rect 1246 2715 1247 2716
rect 1251 2715 1252 2719
rect 1506 2719 1512 2720
rect 1506 2718 1507 2719
rect 1246 2714 1252 2715
rect 1428 2716 1507 2718
rect 1056 2708 1086 2710
rect 1090 2711 1096 2712
rect 1056 2707 1057 2708
rect 1051 2706 1057 2707
rect 1090 2707 1091 2711
rect 1095 2710 1096 2711
rect 1187 2711 1193 2712
rect 1187 2710 1188 2711
rect 1095 2708 1188 2710
rect 1095 2707 1096 2708
rect 1090 2706 1096 2707
rect 1187 2707 1188 2708
rect 1192 2707 1193 2711
rect 1187 2706 1193 2707
rect 1323 2711 1329 2712
rect 1323 2707 1324 2711
rect 1328 2710 1329 2711
rect 1428 2710 1430 2716
rect 1506 2715 1507 2716
rect 1511 2715 1512 2719
rect 3036 2718 3038 2720
rect 3258 2719 3264 2720
rect 3258 2718 3259 2719
rect 3036 2716 3259 2718
rect 1506 2714 1512 2715
rect 3258 2715 3259 2716
rect 3263 2715 3264 2719
rect 3258 2714 3264 2715
rect 1328 2708 1430 2710
rect 1434 2711 1440 2712
rect 1328 2707 1329 2708
rect 1323 2706 1329 2707
rect 1434 2707 1435 2711
rect 1439 2710 1440 2711
rect 1459 2711 1465 2712
rect 1459 2710 1460 2711
rect 1439 2708 1460 2710
rect 1439 2707 1440 2708
rect 1434 2706 1440 2707
rect 1459 2707 1460 2708
rect 1464 2707 1465 2711
rect 1459 2706 1465 2707
rect 1498 2711 1504 2712
rect 1498 2707 1499 2711
rect 1503 2710 1504 2711
rect 1603 2711 1609 2712
rect 1603 2710 1604 2711
rect 1503 2708 1604 2710
rect 1503 2707 1504 2708
rect 1498 2706 1504 2707
rect 1603 2707 1604 2708
rect 1608 2707 1609 2711
rect 1603 2706 1609 2707
rect 2046 2708 2052 2709
rect 3942 2708 3948 2709
rect 2046 2704 2047 2708
rect 2051 2704 2052 2708
rect 2046 2703 2052 2704
rect 2334 2707 2340 2708
rect 2334 2703 2335 2707
rect 2339 2703 2340 2707
rect 298 2702 304 2703
rect 2334 2702 2340 2703
rect 2494 2707 2500 2708
rect 2494 2703 2495 2707
rect 2499 2703 2500 2707
rect 2494 2702 2500 2703
rect 2662 2707 2668 2708
rect 2662 2703 2663 2707
rect 2667 2703 2668 2707
rect 2662 2702 2668 2703
rect 2830 2707 2836 2708
rect 2830 2703 2831 2707
rect 2835 2703 2836 2707
rect 2830 2702 2836 2703
rect 2998 2707 3004 2708
rect 2998 2703 2999 2707
rect 3003 2703 3004 2707
rect 2998 2702 3004 2703
rect 3166 2707 3172 2708
rect 3166 2703 3167 2707
rect 3171 2703 3172 2707
rect 3166 2702 3172 2703
rect 3334 2707 3340 2708
rect 3334 2703 3335 2707
rect 3339 2703 3340 2707
rect 3334 2702 3340 2703
rect 3510 2707 3516 2708
rect 3510 2703 3511 2707
rect 3515 2703 3516 2707
rect 3510 2702 3516 2703
rect 3686 2707 3692 2708
rect 3686 2703 3687 2707
rect 3691 2703 3692 2707
rect 3686 2702 3692 2703
rect 3838 2707 3844 2708
rect 3838 2703 3839 2707
rect 3843 2703 3844 2707
rect 3942 2704 3943 2708
rect 3947 2704 3948 2708
rect 3942 2703 3948 2704
rect 3838 2702 3844 2703
rect 2410 2699 2416 2700
rect 259 2695 265 2696
rect 259 2691 260 2695
rect 264 2694 265 2695
rect 306 2695 312 2696
rect 306 2694 307 2695
rect 264 2692 307 2694
rect 264 2691 265 2692
rect 259 2690 265 2691
rect 306 2691 307 2692
rect 311 2691 312 2695
rect 306 2690 312 2691
rect 403 2695 409 2696
rect 403 2691 404 2695
rect 408 2694 409 2695
rect 434 2695 440 2696
rect 434 2694 435 2695
rect 408 2692 435 2694
rect 408 2691 409 2692
rect 403 2690 409 2691
rect 434 2691 435 2692
rect 439 2691 440 2695
rect 434 2690 440 2691
rect 539 2695 545 2696
rect 539 2691 540 2695
rect 544 2694 545 2695
rect 554 2695 560 2696
rect 554 2694 555 2695
rect 544 2692 555 2694
rect 544 2691 545 2692
rect 539 2690 545 2691
rect 554 2691 555 2692
rect 559 2691 560 2695
rect 554 2690 560 2691
rect 578 2695 584 2696
rect 578 2691 579 2695
rect 583 2694 584 2695
rect 675 2695 681 2696
rect 675 2694 676 2695
rect 583 2692 676 2694
rect 583 2691 584 2692
rect 578 2690 584 2691
rect 675 2691 676 2692
rect 680 2691 681 2695
rect 675 2690 681 2691
rect 714 2695 720 2696
rect 714 2691 715 2695
rect 719 2694 720 2695
rect 803 2695 809 2696
rect 803 2694 804 2695
rect 719 2692 804 2694
rect 719 2691 720 2692
rect 714 2690 720 2691
rect 803 2691 804 2692
rect 808 2691 809 2695
rect 803 2690 809 2691
rect 923 2695 929 2696
rect 923 2691 924 2695
rect 928 2694 929 2695
rect 970 2695 976 2696
rect 970 2694 971 2695
rect 928 2692 971 2694
rect 928 2691 929 2692
rect 923 2690 929 2691
rect 970 2691 971 2692
rect 975 2691 976 2695
rect 970 2690 976 2691
rect 1035 2695 1041 2696
rect 1035 2691 1036 2695
rect 1040 2694 1041 2695
rect 1082 2695 1088 2696
rect 1082 2694 1083 2695
rect 1040 2692 1083 2694
rect 1040 2691 1041 2692
rect 1035 2690 1041 2691
rect 1082 2691 1083 2692
rect 1087 2691 1088 2695
rect 1238 2695 1244 2696
rect 1082 2690 1088 2691
rect 1147 2693 1153 2694
rect 1147 2689 1148 2693
rect 1152 2689 1153 2693
rect 1238 2691 1239 2695
rect 1243 2694 1244 2695
rect 1267 2695 1273 2696
rect 1267 2694 1268 2695
rect 1243 2692 1268 2694
rect 1243 2691 1244 2692
rect 1238 2690 1244 2691
rect 1267 2691 1268 2692
rect 1272 2691 1273 2695
rect 1267 2690 1273 2691
rect 1306 2695 1312 2696
rect 1306 2691 1307 2695
rect 1311 2694 1312 2695
rect 1387 2695 1393 2696
rect 1387 2694 1388 2695
rect 1311 2692 1388 2694
rect 1311 2691 1312 2692
rect 1306 2690 1312 2691
rect 1387 2691 1388 2692
rect 1392 2691 1393 2695
rect 2410 2695 2411 2699
rect 2415 2695 2416 2699
rect 2599 2699 2605 2700
rect 2599 2698 2600 2699
rect 2573 2696 2600 2698
rect 2410 2694 2416 2695
rect 2599 2695 2600 2696
rect 2604 2695 2605 2699
rect 2599 2694 2605 2695
rect 2738 2699 2744 2700
rect 2738 2695 2739 2699
rect 2743 2695 2744 2699
rect 2738 2694 2744 2695
rect 2791 2699 2797 2700
rect 2791 2695 2792 2699
rect 2796 2698 2797 2699
rect 3074 2699 3080 2700
rect 2796 2696 2873 2698
rect 2796 2695 2797 2696
rect 2791 2694 2797 2695
rect 3074 2695 3075 2699
rect 3079 2695 3080 2699
rect 3258 2699 3264 2700
rect 3074 2694 3080 2695
rect 3242 2695 3248 2696
rect 1387 2690 1393 2691
rect 2046 2691 2052 2692
rect 1147 2688 1153 2689
rect 1148 2686 1150 2688
rect 1314 2687 1320 2688
rect 1314 2686 1315 2687
rect 1148 2684 1315 2686
rect 1314 2683 1315 2684
rect 1319 2683 1320 2687
rect 2046 2687 2047 2691
rect 2051 2687 2052 2691
rect 3242 2691 3243 2695
rect 3247 2691 3248 2695
rect 3258 2695 3259 2699
rect 3263 2698 3264 2699
rect 3586 2699 3592 2700
rect 3263 2696 3377 2698
rect 3263 2695 3264 2696
rect 3258 2694 3264 2695
rect 3586 2695 3587 2699
rect 3591 2695 3592 2699
rect 3586 2694 3592 2695
rect 3762 2699 3768 2700
rect 3762 2695 3763 2699
rect 3767 2695 3768 2699
rect 3762 2694 3768 2695
rect 3242 2690 3248 2691
rect 3906 2691 3912 2692
rect 2046 2686 2052 2687
rect 2334 2688 2340 2689
rect 2334 2684 2335 2688
rect 2339 2684 2340 2688
rect 2334 2683 2340 2684
rect 2494 2688 2500 2689
rect 2494 2684 2495 2688
rect 2499 2684 2500 2688
rect 2494 2683 2500 2684
rect 2662 2688 2668 2689
rect 2662 2684 2663 2688
rect 2667 2684 2668 2688
rect 2662 2683 2668 2684
rect 2830 2688 2836 2689
rect 2830 2684 2831 2688
rect 2835 2684 2836 2688
rect 2830 2683 2836 2684
rect 2998 2688 3004 2689
rect 2998 2684 2999 2688
rect 3003 2684 3004 2688
rect 2998 2683 3004 2684
rect 3166 2688 3172 2689
rect 3166 2684 3167 2688
rect 3171 2684 3172 2688
rect 3166 2683 3172 2684
rect 3334 2688 3340 2689
rect 3334 2684 3335 2688
rect 3339 2684 3340 2688
rect 3334 2683 3340 2684
rect 3510 2688 3516 2689
rect 3510 2684 3511 2688
rect 3515 2684 3516 2688
rect 3510 2683 3516 2684
rect 3686 2688 3692 2689
rect 3686 2684 3687 2688
rect 3691 2684 3692 2688
rect 3686 2683 3692 2684
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3906 2687 3907 2691
rect 3911 2690 3912 2691
rect 3916 2690 3918 2693
rect 3911 2688 3918 2690
rect 3942 2691 3948 2692
rect 3911 2687 3912 2688
rect 3906 2686 3912 2687
rect 3942 2687 3943 2691
rect 3947 2687 3948 2691
rect 3942 2686 3948 2687
rect 3838 2683 3844 2684
rect 1314 2682 1320 2683
rect 110 2676 116 2677
rect 2006 2676 2012 2677
rect 110 2672 111 2676
rect 115 2672 116 2676
rect 110 2671 116 2672
rect 222 2675 228 2676
rect 222 2671 223 2675
rect 227 2671 228 2675
rect 222 2670 228 2671
rect 366 2675 372 2676
rect 366 2671 367 2675
rect 371 2671 372 2675
rect 366 2670 372 2671
rect 502 2675 508 2676
rect 502 2671 503 2675
rect 507 2671 508 2675
rect 502 2670 508 2671
rect 638 2675 644 2676
rect 638 2671 639 2675
rect 643 2671 644 2675
rect 638 2670 644 2671
rect 766 2675 772 2676
rect 766 2671 767 2675
rect 771 2671 772 2675
rect 766 2670 772 2671
rect 886 2675 892 2676
rect 886 2671 887 2675
rect 891 2671 892 2675
rect 886 2670 892 2671
rect 998 2675 1004 2676
rect 998 2671 999 2675
rect 1003 2671 1004 2675
rect 998 2670 1004 2671
rect 1110 2675 1116 2676
rect 1110 2671 1111 2675
rect 1115 2671 1116 2675
rect 1110 2670 1116 2671
rect 1230 2675 1236 2676
rect 1230 2671 1231 2675
rect 1235 2671 1236 2675
rect 1230 2670 1236 2671
rect 1350 2675 1356 2676
rect 1350 2671 1351 2675
rect 1355 2671 1356 2675
rect 2006 2672 2007 2676
rect 2011 2672 2012 2676
rect 2006 2671 2012 2672
rect 1350 2670 1356 2671
rect 298 2667 304 2668
rect 298 2663 299 2667
rect 303 2663 304 2667
rect 298 2662 304 2663
rect 306 2667 312 2668
rect 306 2663 307 2667
rect 311 2666 312 2667
rect 578 2667 584 2668
rect 311 2664 409 2666
rect 311 2663 312 2664
rect 306 2662 312 2663
rect 578 2663 579 2667
rect 583 2663 584 2667
rect 578 2662 584 2663
rect 714 2667 720 2668
rect 714 2663 715 2667
rect 719 2663 720 2667
rect 714 2662 720 2663
rect 750 2667 756 2668
rect 750 2663 751 2667
rect 755 2666 756 2667
rect 878 2667 884 2668
rect 755 2664 809 2666
rect 755 2663 756 2664
rect 750 2662 756 2663
rect 878 2663 879 2667
rect 883 2666 884 2667
rect 970 2667 976 2668
rect 883 2664 929 2666
rect 883 2663 884 2664
rect 878 2662 884 2663
rect 970 2663 971 2667
rect 975 2666 976 2667
rect 1082 2667 1088 2668
rect 975 2664 1041 2666
rect 975 2663 976 2664
rect 970 2662 976 2663
rect 1082 2663 1083 2667
rect 1087 2666 1088 2667
rect 1306 2667 1312 2668
rect 1087 2664 1153 2666
rect 1087 2663 1088 2664
rect 1082 2662 1088 2663
rect 1306 2663 1307 2667
rect 1311 2663 1312 2667
rect 1306 2662 1312 2663
rect 1314 2667 1320 2668
rect 1314 2663 1315 2667
rect 1319 2666 1320 2667
rect 1319 2664 1393 2666
rect 1319 2663 1320 2664
rect 1314 2662 1320 2663
rect 110 2659 116 2660
rect 110 2655 111 2659
rect 115 2655 116 2659
rect 2006 2659 2012 2660
rect 110 2654 116 2655
rect 222 2656 228 2657
rect 222 2652 223 2656
rect 227 2652 228 2656
rect 222 2651 228 2652
rect 366 2656 372 2657
rect 366 2652 367 2656
rect 371 2652 372 2656
rect 366 2651 372 2652
rect 502 2656 508 2657
rect 502 2652 503 2656
rect 507 2652 508 2656
rect 502 2651 508 2652
rect 638 2656 644 2657
rect 638 2652 639 2656
rect 643 2652 644 2656
rect 638 2651 644 2652
rect 766 2656 772 2657
rect 766 2652 767 2656
rect 771 2652 772 2656
rect 766 2651 772 2652
rect 886 2656 892 2657
rect 886 2652 887 2656
rect 891 2652 892 2656
rect 886 2651 892 2652
rect 998 2656 1004 2657
rect 998 2652 999 2656
rect 1003 2652 1004 2656
rect 998 2651 1004 2652
rect 1110 2656 1116 2657
rect 1110 2652 1111 2656
rect 1115 2652 1116 2656
rect 1110 2651 1116 2652
rect 1230 2656 1236 2657
rect 1230 2652 1231 2656
rect 1235 2652 1236 2656
rect 1230 2651 1236 2652
rect 1350 2656 1356 2657
rect 1350 2652 1351 2656
rect 1355 2652 1356 2656
rect 2006 2655 2007 2659
rect 2011 2655 2012 2659
rect 2006 2654 2012 2655
rect 1350 2651 1356 2652
rect 2402 2631 2408 2632
rect 2402 2627 2403 2631
rect 2407 2630 2408 2631
rect 2407 2628 2710 2630
rect 2407 2627 2408 2628
rect 2402 2626 2408 2627
rect 2126 2624 2132 2625
rect 2046 2621 2052 2622
rect 2046 2617 2047 2621
rect 2051 2617 2052 2621
rect 2126 2620 2127 2624
rect 2131 2620 2132 2624
rect 2126 2619 2132 2620
rect 2278 2624 2284 2625
rect 2278 2620 2279 2624
rect 2283 2620 2284 2624
rect 2278 2619 2284 2620
rect 2446 2624 2452 2625
rect 2446 2620 2447 2624
rect 2451 2620 2452 2624
rect 2446 2619 2452 2620
rect 2622 2624 2628 2625
rect 2622 2620 2623 2624
rect 2627 2620 2628 2624
rect 2622 2619 2628 2620
rect 2046 2616 2052 2617
rect 2202 2615 2208 2616
rect 2202 2611 2203 2615
rect 2207 2611 2208 2615
rect 2202 2610 2208 2611
rect 2354 2615 2360 2616
rect 2354 2611 2355 2615
rect 2359 2611 2360 2615
rect 2354 2610 2360 2611
rect 2522 2615 2528 2616
rect 2522 2611 2523 2615
rect 2527 2611 2528 2615
rect 2522 2610 2528 2611
rect 2698 2615 2704 2616
rect 2698 2611 2699 2615
rect 2703 2611 2704 2615
rect 2708 2614 2710 2628
rect 2806 2624 2812 2625
rect 2806 2620 2807 2624
rect 2811 2620 2812 2624
rect 2806 2619 2812 2620
rect 2990 2624 2996 2625
rect 2990 2620 2991 2624
rect 2995 2620 2996 2624
rect 2990 2619 2996 2620
rect 3174 2624 3180 2625
rect 3174 2620 3175 2624
rect 3179 2620 3180 2624
rect 3174 2619 3180 2620
rect 3350 2624 3356 2625
rect 3350 2620 3351 2624
rect 3355 2620 3356 2624
rect 3350 2619 3356 2620
rect 3518 2624 3524 2625
rect 3518 2620 3519 2624
rect 3523 2620 3524 2624
rect 3518 2619 3524 2620
rect 3686 2624 3692 2625
rect 3686 2620 3687 2624
rect 3691 2620 3692 2624
rect 3686 2619 3692 2620
rect 3838 2624 3844 2625
rect 3838 2620 3839 2624
rect 3843 2620 3844 2624
rect 3838 2619 3844 2620
rect 3942 2621 3948 2622
rect 3942 2617 3943 2621
rect 3947 2617 3948 2621
rect 3942 2616 3948 2617
rect 2890 2615 2896 2616
rect 2708 2612 2849 2614
rect 2698 2610 2704 2611
rect 2890 2611 2891 2615
rect 2895 2614 2896 2615
rect 3102 2615 3108 2616
rect 2895 2612 3033 2614
rect 2895 2611 2896 2612
rect 2890 2610 2896 2611
rect 3102 2611 3103 2615
rect 3107 2614 3108 2615
rect 3426 2615 3432 2616
rect 3107 2612 3217 2614
rect 3107 2611 3108 2612
rect 3102 2610 3108 2611
rect 3426 2611 3427 2615
rect 3431 2611 3432 2615
rect 3426 2610 3432 2611
rect 3586 2615 3592 2616
rect 3586 2611 3587 2615
rect 3591 2611 3592 2615
rect 3586 2610 3592 2611
rect 3618 2615 3624 2616
rect 3618 2611 3619 2615
rect 3623 2614 3624 2615
rect 3922 2615 3928 2616
rect 3922 2614 3923 2615
rect 3623 2612 3729 2614
rect 3917 2612 3923 2614
rect 3623 2611 3624 2612
rect 3618 2610 3624 2611
rect 3922 2611 3923 2612
rect 3927 2611 3928 2615
rect 3922 2610 3928 2611
rect 2126 2605 2132 2606
rect 2046 2604 2052 2605
rect 2046 2600 2047 2604
rect 2051 2600 2052 2604
rect 2126 2601 2127 2605
rect 2131 2601 2132 2605
rect 2126 2600 2132 2601
rect 2278 2605 2284 2606
rect 2278 2601 2279 2605
rect 2283 2601 2284 2605
rect 2278 2600 2284 2601
rect 2446 2605 2452 2606
rect 2446 2601 2447 2605
rect 2451 2601 2452 2605
rect 2446 2600 2452 2601
rect 2622 2605 2628 2606
rect 2622 2601 2623 2605
rect 2627 2601 2628 2605
rect 2622 2600 2628 2601
rect 2806 2605 2812 2606
rect 2806 2601 2807 2605
rect 2811 2601 2812 2605
rect 2806 2600 2812 2601
rect 2990 2605 2996 2606
rect 2990 2601 2991 2605
rect 2995 2601 2996 2605
rect 2990 2600 2996 2601
rect 3174 2605 3180 2606
rect 3174 2601 3175 2605
rect 3179 2601 3180 2605
rect 3174 2600 3180 2601
rect 3350 2605 3356 2606
rect 3350 2601 3351 2605
rect 3355 2601 3356 2605
rect 3350 2600 3356 2601
rect 3518 2605 3524 2606
rect 3518 2601 3519 2605
rect 3523 2601 3524 2605
rect 3518 2600 3524 2601
rect 3686 2605 3692 2606
rect 3686 2601 3687 2605
rect 3691 2601 3692 2605
rect 3686 2600 3692 2601
rect 3838 2605 3844 2606
rect 3838 2601 3839 2605
rect 3843 2601 3844 2605
rect 3838 2600 3844 2601
rect 3942 2604 3948 2605
rect 3942 2600 3943 2604
rect 3947 2600 3948 2604
rect 2046 2599 2052 2600
rect 3942 2599 3948 2600
rect 174 2596 180 2597
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 174 2592 175 2596
rect 179 2592 180 2596
rect 174 2591 180 2592
rect 366 2596 372 2597
rect 366 2592 367 2596
rect 371 2592 372 2596
rect 366 2591 372 2592
rect 542 2596 548 2597
rect 542 2592 543 2596
rect 547 2592 548 2596
rect 542 2591 548 2592
rect 710 2596 716 2597
rect 710 2592 711 2596
rect 715 2592 716 2596
rect 710 2591 716 2592
rect 862 2596 868 2597
rect 862 2592 863 2596
rect 867 2592 868 2596
rect 862 2591 868 2592
rect 1006 2596 1012 2597
rect 1006 2592 1007 2596
rect 1011 2592 1012 2596
rect 1006 2591 1012 2592
rect 1142 2596 1148 2597
rect 1142 2592 1143 2596
rect 1147 2592 1148 2596
rect 1142 2591 1148 2592
rect 1278 2596 1284 2597
rect 1278 2592 1279 2596
rect 1283 2592 1284 2596
rect 1278 2591 1284 2592
rect 1422 2596 1428 2597
rect 1422 2592 1423 2596
rect 1427 2592 1428 2596
rect 3618 2595 3624 2596
rect 3618 2594 3619 2595
rect 1422 2591 1428 2592
rect 2006 2593 2012 2594
rect 110 2588 116 2589
rect 2006 2589 2007 2593
rect 2011 2589 2012 2593
rect 2006 2588 2012 2589
rect 3420 2592 3619 2594
rect 250 2587 256 2588
rect 250 2583 251 2587
rect 255 2583 256 2587
rect 250 2582 256 2583
rect 434 2587 440 2588
rect 434 2583 435 2587
rect 439 2583 440 2587
rect 434 2582 440 2583
rect 618 2587 624 2588
rect 618 2583 619 2587
rect 623 2583 624 2587
rect 618 2582 624 2583
rect 630 2587 636 2588
rect 630 2583 631 2587
rect 635 2586 636 2587
rect 938 2587 944 2588
rect 635 2584 753 2586
rect 635 2583 636 2584
rect 630 2582 636 2583
rect 938 2583 939 2587
rect 943 2583 944 2587
rect 938 2582 944 2583
rect 1082 2587 1088 2588
rect 1082 2583 1083 2587
rect 1087 2583 1088 2587
rect 1082 2582 1088 2583
rect 1218 2587 1224 2588
rect 1218 2583 1219 2587
rect 1223 2583 1224 2587
rect 1218 2582 1224 2583
rect 1354 2587 1360 2588
rect 1354 2583 1355 2587
rect 1359 2583 1360 2587
rect 1354 2582 1360 2583
rect 1366 2587 1372 2588
rect 1366 2583 1367 2587
rect 1371 2586 1372 2587
rect 2202 2587 2208 2588
rect 1371 2584 1465 2586
rect 1371 2583 1372 2584
rect 1366 2582 1372 2583
rect 2163 2583 2172 2584
rect 2163 2579 2164 2583
rect 2171 2579 2172 2583
rect 2202 2583 2203 2587
rect 2207 2586 2208 2587
rect 2315 2587 2321 2588
rect 2315 2586 2316 2587
rect 2207 2584 2316 2586
rect 2207 2583 2208 2584
rect 2202 2582 2208 2583
rect 2315 2583 2316 2584
rect 2320 2583 2321 2587
rect 2315 2582 2321 2583
rect 2354 2587 2360 2588
rect 2354 2583 2355 2587
rect 2359 2586 2360 2587
rect 2483 2587 2489 2588
rect 2483 2586 2484 2587
rect 2359 2584 2484 2586
rect 2359 2583 2360 2584
rect 2354 2582 2360 2583
rect 2483 2583 2484 2584
rect 2488 2583 2489 2587
rect 2483 2582 2489 2583
rect 2522 2587 2528 2588
rect 2522 2583 2523 2587
rect 2527 2586 2528 2587
rect 2659 2587 2665 2588
rect 2659 2586 2660 2587
rect 2527 2584 2660 2586
rect 2527 2583 2528 2584
rect 2522 2582 2528 2583
rect 2659 2583 2660 2584
rect 2664 2583 2665 2587
rect 2659 2582 2665 2583
rect 2698 2587 2704 2588
rect 2698 2583 2699 2587
rect 2703 2586 2704 2587
rect 2843 2587 2849 2588
rect 2843 2586 2844 2587
rect 2703 2584 2844 2586
rect 2703 2583 2704 2584
rect 2698 2582 2704 2583
rect 2843 2583 2844 2584
rect 2848 2583 2849 2587
rect 2843 2582 2849 2583
rect 3027 2587 3033 2588
rect 3027 2583 3028 2587
rect 3032 2586 3033 2587
rect 3102 2587 3108 2588
rect 3102 2586 3103 2587
rect 3032 2584 3103 2586
rect 3032 2583 3033 2584
rect 3027 2582 3033 2583
rect 3102 2583 3103 2584
rect 3107 2583 3108 2587
rect 3102 2582 3108 2583
rect 3211 2587 3217 2588
rect 3211 2583 3212 2587
rect 3216 2586 3217 2587
rect 3242 2587 3248 2588
rect 3242 2586 3243 2587
rect 3216 2584 3243 2586
rect 3216 2583 3217 2584
rect 3211 2582 3217 2583
rect 3242 2583 3243 2584
rect 3247 2583 3248 2587
rect 3242 2582 3248 2583
rect 3387 2587 3393 2588
rect 3387 2583 3388 2587
rect 3392 2586 3393 2587
rect 3420 2586 3422 2592
rect 3618 2591 3619 2592
rect 3623 2591 3624 2595
rect 3618 2590 3624 2591
rect 3392 2584 3422 2586
rect 3426 2587 3432 2588
rect 3392 2583 3393 2584
rect 3387 2582 3393 2583
rect 3426 2583 3427 2587
rect 3431 2586 3432 2587
rect 3555 2587 3561 2588
rect 3555 2586 3556 2587
rect 3431 2584 3556 2586
rect 3431 2583 3432 2584
rect 3426 2582 3432 2583
rect 3555 2583 3556 2584
rect 3560 2583 3561 2587
rect 3875 2587 3881 2588
rect 3555 2582 3561 2583
rect 3723 2583 3732 2584
rect 2163 2578 2172 2579
rect 3723 2579 3724 2583
rect 3731 2579 3732 2583
rect 3875 2583 3876 2587
rect 3880 2586 3881 2587
rect 3906 2587 3912 2588
rect 3906 2586 3907 2587
rect 3880 2584 3907 2586
rect 3880 2583 3881 2584
rect 3875 2582 3881 2583
rect 3906 2583 3907 2584
rect 3911 2583 3912 2587
rect 3906 2582 3912 2583
rect 3723 2578 3732 2579
rect 174 2577 180 2578
rect 110 2576 116 2577
rect 110 2572 111 2576
rect 115 2572 116 2576
rect 174 2573 175 2577
rect 179 2573 180 2577
rect 174 2572 180 2573
rect 366 2577 372 2578
rect 366 2573 367 2577
rect 371 2573 372 2577
rect 366 2572 372 2573
rect 542 2577 548 2578
rect 542 2573 543 2577
rect 547 2573 548 2577
rect 542 2572 548 2573
rect 710 2577 716 2578
rect 710 2573 711 2577
rect 715 2573 716 2577
rect 710 2572 716 2573
rect 862 2577 868 2578
rect 862 2573 863 2577
rect 867 2573 868 2577
rect 862 2572 868 2573
rect 1006 2577 1012 2578
rect 1006 2573 1007 2577
rect 1011 2573 1012 2577
rect 1006 2572 1012 2573
rect 1142 2577 1148 2578
rect 1142 2573 1143 2577
rect 1147 2573 1148 2577
rect 1142 2572 1148 2573
rect 1278 2577 1284 2578
rect 1278 2573 1279 2577
rect 1283 2573 1284 2577
rect 1278 2572 1284 2573
rect 1422 2577 1428 2578
rect 1422 2573 1423 2577
rect 1427 2573 1428 2577
rect 1422 2572 1428 2573
rect 2006 2576 2012 2577
rect 2006 2572 2007 2576
rect 2011 2572 2012 2576
rect 110 2571 116 2572
rect 2006 2571 2012 2572
rect 2146 2563 2152 2564
rect 2107 2561 2113 2562
rect 250 2559 256 2560
rect 210 2555 217 2556
rect 210 2551 211 2555
rect 216 2551 217 2555
rect 250 2555 251 2559
rect 255 2558 256 2559
rect 403 2559 409 2560
rect 403 2558 404 2559
rect 255 2556 404 2558
rect 255 2555 256 2556
rect 250 2554 256 2555
rect 403 2555 404 2556
rect 408 2555 409 2559
rect 403 2554 409 2555
rect 579 2559 585 2560
rect 579 2555 580 2559
rect 584 2558 585 2559
rect 630 2559 636 2560
rect 630 2558 631 2559
rect 584 2556 631 2558
rect 584 2555 585 2556
rect 579 2554 585 2555
rect 630 2555 631 2556
rect 635 2555 636 2559
rect 630 2554 636 2555
rect 747 2559 756 2560
rect 747 2555 748 2559
rect 755 2555 756 2559
rect 747 2554 756 2555
rect 878 2559 884 2560
rect 878 2555 879 2559
rect 883 2558 884 2559
rect 899 2559 905 2560
rect 899 2558 900 2559
rect 883 2556 900 2558
rect 883 2555 884 2556
rect 878 2554 884 2555
rect 899 2555 900 2556
rect 904 2555 905 2559
rect 899 2554 905 2555
rect 938 2559 944 2560
rect 938 2555 939 2559
rect 943 2558 944 2559
rect 1043 2559 1049 2560
rect 1043 2558 1044 2559
rect 943 2556 1044 2558
rect 943 2555 944 2556
rect 938 2554 944 2555
rect 1043 2555 1044 2556
rect 1048 2555 1049 2559
rect 1043 2554 1049 2555
rect 1082 2559 1088 2560
rect 1082 2555 1083 2559
rect 1087 2558 1088 2559
rect 1179 2559 1185 2560
rect 1179 2558 1180 2559
rect 1087 2556 1180 2558
rect 1087 2555 1088 2556
rect 1082 2554 1088 2555
rect 1179 2555 1180 2556
rect 1184 2555 1185 2559
rect 1179 2554 1185 2555
rect 1218 2559 1224 2560
rect 1218 2555 1219 2559
rect 1223 2558 1224 2559
rect 1315 2559 1321 2560
rect 1315 2558 1316 2559
rect 1223 2556 1316 2558
rect 1223 2555 1224 2556
rect 1218 2554 1224 2555
rect 1315 2555 1316 2556
rect 1320 2555 1321 2559
rect 1315 2554 1321 2555
rect 1354 2559 1360 2560
rect 1354 2555 1355 2559
rect 1359 2558 1360 2559
rect 1459 2559 1465 2560
rect 1459 2558 1460 2559
rect 1359 2556 1460 2558
rect 1359 2555 1360 2556
rect 1354 2554 1360 2555
rect 1459 2555 1460 2556
rect 1464 2555 1465 2559
rect 2107 2557 2108 2561
rect 2112 2557 2113 2561
rect 2146 2559 2147 2563
rect 2151 2562 2152 2563
rect 2219 2563 2225 2564
rect 2219 2562 2220 2563
rect 2151 2560 2220 2562
rect 2151 2559 2152 2560
rect 2146 2558 2152 2559
rect 2219 2559 2220 2560
rect 2224 2559 2225 2563
rect 2219 2558 2225 2559
rect 2258 2563 2264 2564
rect 2258 2559 2259 2563
rect 2263 2562 2264 2563
rect 2355 2563 2361 2564
rect 2355 2562 2356 2563
rect 2263 2560 2356 2562
rect 2263 2559 2264 2560
rect 2258 2558 2264 2559
rect 2355 2559 2356 2560
rect 2360 2559 2361 2563
rect 2355 2558 2361 2559
rect 2394 2563 2400 2564
rect 2394 2559 2395 2563
rect 2399 2562 2400 2563
rect 2507 2563 2513 2564
rect 2507 2562 2508 2563
rect 2399 2560 2508 2562
rect 2399 2559 2400 2560
rect 2394 2558 2400 2559
rect 2507 2559 2508 2560
rect 2512 2559 2513 2563
rect 2507 2558 2513 2559
rect 2546 2563 2552 2564
rect 2546 2559 2547 2563
rect 2551 2562 2552 2563
rect 2675 2563 2681 2564
rect 2675 2562 2676 2563
rect 2551 2560 2676 2562
rect 2551 2559 2552 2560
rect 2546 2558 2552 2559
rect 2675 2559 2676 2560
rect 2680 2559 2681 2563
rect 2675 2558 2681 2559
rect 2859 2563 2865 2564
rect 2859 2559 2860 2563
rect 2864 2562 2865 2563
rect 2890 2563 2896 2564
rect 2890 2562 2891 2563
rect 2864 2560 2891 2562
rect 2864 2559 2865 2560
rect 2859 2558 2865 2559
rect 2890 2559 2891 2560
rect 2895 2559 2896 2563
rect 2890 2558 2896 2559
rect 2898 2563 2904 2564
rect 2898 2559 2899 2563
rect 2903 2562 2904 2563
rect 3067 2563 3073 2564
rect 3067 2562 3068 2563
rect 2903 2560 3068 2562
rect 2903 2559 2904 2560
rect 2898 2558 2904 2559
rect 3067 2559 3068 2560
rect 3072 2559 3073 2563
rect 3067 2558 3073 2559
rect 3106 2563 3112 2564
rect 3106 2559 3107 2563
rect 3111 2562 3112 2563
rect 3299 2563 3305 2564
rect 3299 2562 3300 2563
rect 3111 2560 3300 2562
rect 3111 2559 3112 2560
rect 3106 2558 3112 2559
rect 3299 2559 3300 2560
rect 3304 2559 3305 2563
rect 3299 2558 3305 2559
rect 3338 2563 3344 2564
rect 3338 2559 3339 2563
rect 3343 2562 3344 2563
rect 3539 2563 3545 2564
rect 3539 2562 3540 2563
rect 3343 2560 3540 2562
rect 3343 2559 3344 2560
rect 3338 2558 3344 2559
rect 3539 2559 3540 2560
rect 3544 2559 3545 2563
rect 3539 2558 3545 2559
rect 3698 2563 3704 2564
rect 3698 2559 3699 2563
rect 3703 2562 3704 2563
rect 3779 2563 3785 2564
rect 3779 2562 3780 2563
rect 3703 2560 3780 2562
rect 3703 2559 3704 2560
rect 3698 2558 3704 2559
rect 3779 2559 3780 2560
rect 3784 2559 3785 2563
rect 3779 2558 3785 2559
rect 2107 2556 2113 2557
rect 1459 2554 1465 2555
rect 2108 2554 2110 2556
rect 2298 2555 2304 2556
rect 2298 2554 2299 2555
rect 2108 2552 2299 2554
rect 210 2550 217 2551
rect 2298 2551 2299 2552
rect 2303 2551 2304 2555
rect 2298 2550 2304 2551
rect 1366 2547 1372 2548
rect 1366 2546 1367 2547
rect 1116 2544 1367 2546
rect 1116 2542 1118 2544
rect 1366 2543 1367 2544
rect 1371 2543 1372 2547
rect 1366 2542 1372 2543
rect 2046 2544 2052 2545
rect 3942 2544 3948 2545
rect 1115 2541 1121 2542
rect 171 2539 177 2540
rect 171 2535 172 2539
rect 176 2538 177 2539
rect 218 2539 224 2540
rect 218 2538 219 2539
rect 176 2536 219 2538
rect 176 2535 177 2536
rect 171 2534 177 2535
rect 218 2535 219 2536
rect 223 2535 224 2539
rect 218 2534 224 2535
rect 307 2539 313 2540
rect 307 2535 308 2539
rect 312 2538 313 2539
rect 354 2539 360 2540
rect 354 2538 355 2539
rect 312 2536 355 2538
rect 312 2535 313 2536
rect 307 2534 313 2535
rect 354 2535 355 2536
rect 359 2535 360 2539
rect 354 2534 360 2535
rect 475 2539 484 2540
rect 475 2535 476 2539
rect 483 2535 484 2539
rect 475 2534 484 2535
rect 618 2539 624 2540
rect 618 2535 619 2539
rect 623 2538 624 2539
rect 643 2539 649 2540
rect 643 2538 644 2539
rect 623 2536 644 2538
rect 623 2535 624 2536
rect 618 2534 624 2535
rect 643 2535 644 2536
rect 648 2535 649 2539
rect 643 2534 649 2535
rect 682 2539 688 2540
rect 682 2535 683 2539
rect 687 2538 688 2539
rect 811 2539 817 2540
rect 811 2538 812 2539
rect 687 2536 812 2538
rect 687 2535 688 2536
rect 682 2534 688 2535
rect 811 2535 812 2536
rect 816 2535 817 2539
rect 811 2534 817 2535
rect 850 2539 856 2540
rect 850 2535 851 2539
rect 855 2538 856 2539
rect 963 2539 969 2540
rect 963 2538 964 2539
rect 855 2536 964 2538
rect 855 2535 856 2536
rect 850 2534 856 2535
rect 963 2535 964 2536
rect 968 2535 969 2539
rect 1115 2537 1116 2541
rect 1120 2537 1121 2541
rect 2046 2540 2047 2544
rect 2051 2540 2052 2544
rect 1115 2536 1121 2537
rect 1154 2539 1160 2540
rect 963 2534 969 2535
rect 1154 2535 1155 2539
rect 1159 2538 1160 2539
rect 1259 2539 1265 2540
rect 1259 2538 1260 2539
rect 1159 2536 1260 2538
rect 1159 2535 1160 2536
rect 1154 2534 1160 2535
rect 1259 2535 1260 2536
rect 1264 2535 1265 2539
rect 1259 2534 1265 2535
rect 1298 2539 1304 2540
rect 1298 2535 1299 2539
rect 1303 2538 1304 2539
rect 1395 2539 1401 2540
rect 1395 2538 1396 2539
rect 1303 2536 1396 2538
rect 1303 2535 1304 2536
rect 1298 2534 1304 2535
rect 1395 2535 1396 2536
rect 1400 2535 1401 2539
rect 1395 2534 1401 2535
rect 1434 2539 1440 2540
rect 1434 2535 1435 2539
rect 1439 2538 1440 2539
rect 1531 2539 1537 2540
rect 1531 2538 1532 2539
rect 1439 2536 1532 2538
rect 1439 2535 1440 2536
rect 1434 2534 1440 2535
rect 1531 2535 1532 2536
rect 1536 2535 1537 2539
rect 1531 2534 1537 2535
rect 1570 2539 1576 2540
rect 1570 2535 1571 2539
rect 1575 2538 1576 2539
rect 1675 2539 1681 2540
rect 2046 2539 2052 2540
rect 2070 2543 2076 2544
rect 2070 2539 2071 2543
rect 2075 2539 2076 2543
rect 1675 2538 1676 2539
rect 1575 2536 1676 2538
rect 1575 2535 1576 2536
rect 1570 2534 1576 2535
rect 1675 2535 1676 2536
rect 1680 2535 1681 2539
rect 2070 2538 2076 2539
rect 2182 2543 2188 2544
rect 2182 2539 2183 2543
rect 2187 2539 2188 2543
rect 2182 2538 2188 2539
rect 2318 2543 2324 2544
rect 2318 2539 2319 2543
rect 2323 2539 2324 2543
rect 2318 2538 2324 2539
rect 2470 2543 2476 2544
rect 2470 2539 2471 2543
rect 2475 2539 2476 2543
rect 2470 2538 2476 2539
rect 2638 2543 2644 2544
rect 2638 2539 2639 2543
rect 2643 2539 2644 2543
rect 2638 2538 2644 2539
rect 2822 2543 2828 2544
rect 2822 2539 2823 2543
rect 2827 2539 2828 2543
rect 2822 2538 2828 2539
rect 3030 2543 3036 2544
rect 3030 2539 3031 2543
rect 3035 2539 3036 2543
rect 3030 2538 3036 2539
rect 3262 2543 3268 2544
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3502 2543 3508 2544
rect 3502 2539 3503 2543
rect 3507 2539 3508 2543
rect 3502 2538 3508 2539
rect 3742 2543 3748 2544
rect 3742 2539 3743 2543
rect 3747 2539 3748 2543
rect 3942 2540 3943 2544
rect 3947 2540 3948 2544
rect 3942 2539 3948 2540
rect 3742 2538 3748 2539
rect 1675 2534 1681 2535
rect 2146 2535 2152 2536
rect 2146 2531 2147 2535
rect 2151 2531 2152 2535
rect 2146 2530 2152 2531
rect 2258 2535 2264 2536
rect 2258 2531 2259 2535
rect 2263 2531 2264 2535
rect 2258 2530 2264 2531
rect 2394 2535 2400 2536
rect 2394 2531 2395 2535
rect 2399 2531 2400 2535
rect 2394 2530 2400 2531
rect 2546 2535 2552 2536
rect 2546 2531 2547 2535
rect 2551 2531 2552 2535
rect 2546 2530 2552 2531
rect 2598 2535 2604 2536
rect 2598 2531 2599 2535
rect 2603 2534 2604 2535
rect 2898 2535 2904 2536
rect 2603 2532 2681 2534
rect 2603 2531 2604 2532
rect 2598 2530 2604 2531
rect 2898 2531 2899 2535
rect 2903 2531 2904 2535
rect 2898 2530 2904 2531
rect 3106 2535 3112 2536
rect 3106 2531 3107 2535
rect 3111 2531 3112 2535
rect 3106 2530 3112 2531
rect 3338 2535 3344 2536
rect 3338 2531 3339 2535
rect 3343 2531 3344 2535
rect 3338 2530 3344 2531
rect 3450 2535 3456 2536
rect 3450 2531 3451 2535
rect 3455 2534 3456 2535
rect 3726 2535 3732 2536
rect 3455 2532 3545 2534
rect 3455 2531 3456 2532
rect 3450 2530 3456 2531
rect 3726 2531 3727 2535
rect 3731 2534 3732 2535
rect 3731 2532 3785 2534
rect 3731 2531 3732 2532
rect 3726 2530 3732 2531
rect 2046 2527 2052 2528
rect 2046 2523 2047 2527
rect 2051 2523 2052 2527
rect 3942 2527 3948 2528
rect 2046 2522 2052 2523
rect 2070 2524 2076 2525
rect 110 2520 116 2521
rect 2006 2520 2012 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 134 2519 140 2520
rect 134 2515 135 2519
rect 139 2515 140 2519
rect 134 2514 140 2515
rect 270 2519 276 2520
rect 270 2515 271 2519
rect 275 2515 276 2519
rect 270 2514 276 2515
rect 438 2519 444 2520
rect 438 2515 439 2519
rect 443 2515 444 2519
rect 438 2514 444 2515
rect 606 2519 612 2520
rect 606 2515 607 2519
rect 611 2515 612 2519
rect 606 2514 612 2515
rect 774 2519 780 2520
rect 774 2515 775 2519
rect 779 2515 780 2519
rect 774 2514 780 2515
rect 926 2519 932 2520
rect 926 2515 927 2519
rect 931 2515 932 2519
rect 926 2514 932 2515
rect 1078 2519 1084 2520
rect 1078 2515 1079 2519
rect 1083 2515 1084 2519
rect 1078 2514 1084 2515
rect 1222 2519 1228 2520
rect 1222 2515 1223 2519
rect 1227 2515 1228 2519
rect 1222 2514 1228 2515
rect 1358 2519 1364 2520
rect 1358 2515 1359 2519
rect 1363 2515 1364 2519
rect 1358 2514 1364 2515
rect 1494 2519 1500 2520
rect 1494 2515 1495 2519
rect 1499 2515 1500 2519
rect 1494 2514 1500 2515
rect 1638 2519 1644 2520
rect 1638 2515 1639 2519
rect 1643 2515 1644 2519
rect 2006 2516 2007 2520
rect 2011 2516 2012 2520
rect 2070 2520 2071 2524
rect 2075 2520 2076 2524
rect 2070 2519 2076 2520
rect 2182 2524 2188 2525
rect 2182 2520 2183 2524
rect 2187 2520 2188 2524
rect 2182 2519 2188 2520
rect 2318 2524 2324 2525
rect 2318 2520 2319 2524
rect 2323 2520 2324 2524
rect 2318 2519 2324 2520
rect 2470 2524 2476 2525
rect 2470 2520 2471 2524
rect 2475 2520 2476 2524
rect 2470 2519 2476 2520
rect 2638 2524 2644 2525
rect 2638 2520 2639 2524
rect 2643 2520 2644 2524
rect 2638 2519 2644 2520
rect 2822 2524 2828 2525
rect 2822 2520 2823 2524
rect 2827 2520 2828 2524
rect 2822 2519 2828 2520
rect 3030 2524 3036 2525
rect 3030 2520 3031 2524
rect 3035 2520 3036 2524
rect 3030 2519 3036 2520
rect 3262 2524 3268 2525
rect 3262 2520 3263 2524
rect 3267 2520 3268 2524
rect 3262 2519 3268 2520
rect 3502 2524 3508 2525
rect 3502 2520 3503 2524
rect 3507 2520 3508 2524
rect 3502 2519 3508 2520
rect 3742 2524 3748 2525
rect 3742 2520 3743 2524
rect 3747 2520 3748 2524
rect 3942 2523 3943 2527
rect 3947 2523 3948 2527
rect 3942 2522 3948 2523
rect 3742 2519 3748 2520
rect 2006 2515 2012 2516
rect 1638 2514 1644 2515
rect 210 2511 216 2512
rect 210 2507 211 2511
rect 215 2507 216 2511
rect 210 2506 216 2507
rect 218 2511 224 2512
rect 218 2507 219 2511
rect 223 2510 224 2511
rect 354 2511 360 2512
rect 223 2508 313 2510
rect 223 2507 224 2508
rect 218 2506 224 2507
rect 354 2507 355 2511
rect 359 2510 360 2511
rect 682 2511 688 2512
rect 359 2508 481 2510
rect 359 2507 360 2508
rect 354 2506 360 2507
rect 682 2507 683 2511
rect 687 2507 688 2511
rect 682 2506 688 2507
rect 850 2511 856 2512
rect 850 2507 851 2511
rect 855 2507 856 2511
rect 1154 2511 1160 2512
rect 850 2506 856 2507
rect 1002 2507 1008 2508
rect 110 2503 116 2504
rect 110 2499 111 2503
rect 115 2499 116 2503
rect 1002 2503 1003 2507
rect 1007 2503 1008 2507
rect 1154 2507 1155 2511
rect 1159 2507 1160 2511
rect 1154 2506 1160 2507
rect 1298 2511 1304 2512
rect 1298 2507 1299 2511
rect 1303 2507 1304 2511
rect 1298 2506 1304 2507
rect 1434 2511 1440 2512
rect 1434 2507 1435 2511
rect 1439 2507 1440 2511
rect 1434 2506 1440 2507
rect 1570 2511 1576 2512
rect 1570 2507 1571 2511
rect 1575 2507 1576 2511
rect 1570 2506 1576 2507
rect 1578 2511 1584 2512
rect 1578 2507 1579 2511
rect 1583 2510 1584 2511
rect 1583 2508 1681 2510
rect 1583 2507 1584 2508
rect 1578 2506 1584 2507
rect 1002 2502 1008 2503
rect 2006 2503 2012 2504
rect 110 2498 116 2499
rect 134 2500 140 2501
rect 134 2496 135 2500
rect 139 2496 140 2500
rect 134 2495 140 2496
rect 270 2500 276 2501
rect 270 2496 271 2500
rect 275 2496 276 2500
rect 270 2495 276 2496
rect 438 2500 444 2501
rect 438 2496 439 2500
rect 443 2496 444 2500
rect 438 2495 444 2496
rect 606 2500 612 2501
rect 606 2496 607 2500
rect 611 2496 612 2500
rect 606 2495 612 2496
rect 774 2500 780 2501
rect 774 2496 775 2500
rect 779 2496 780 2500
rect 774 2495 780 2496
rect 926 2500 932 2501
rect 926 2496 927 2500
rect 931 2496 932 2500
rect 926 2495 932 2496
rect 1078 2500 1084 2501
rect 1078 2496 1079 2500
rect 1083 2496 1084 2500
rect 1078 2495 1084 2496
rect 1222 2500 1228 2501
rect 1222 2496 1223 2500
rect 1227 2496 1228 2500
rect 1222 2495 1228 2496
rect 1358 2500 1364 2501
rect 1358 2496 1359 2500
rect 1363 2496 1364 2500
rect 1358 2495 1364 2496
rect 1494 2500 1500 2501
rect 1494 2496 1495 2500
rect 1499 2496 1500 2500
rect 1494 2495 1500 2496
rect 1638 2500 1644 2501
rect 1638 2496 1639 2500
rect 1643 2496 1644 2500
rect 2006 2499 2007 2503
rect 2011 2499 2012 2503
rect 2006 2498 2012 2499
rect 1638 2495 1644 2496
rect 2070 2460 2076 2461
rect 2046 2457 2052 2458
rect 2046 2453 2047 2457
rect 2051 2453 2052 2457
rect 2070 2456 2071 2460
rect 2075 2456 2076 2460
rect 2070 2455 2076 2456
rect 2214 2460 2220 2461
rect 2214 2456 2215 2460
rect 2219 2456 2220 2460
rect 2214 2455 2220 2456
rect 2382 2460 2388 2461
rect 2382 2456 2383 2460
rect 2387 2456 2388 2460
rect 2382 2455 2388 2456
rect 2558 2460 2564 2461
rect 2558 2456 2559 2460
rect 2563 2456 2564 2460
rect 2558 2455 2564 2456
rect 2750 2460 2756 2461
rect 2750 2456 2751 2460
rect 2755 2456 2756 2460
rect 2750 2455 2756 2456
rect 2950 2460 2956 2461
rect 2950 2456 2951 2460
rect 2955 2456 2956 2460
rect 2950 2455 2956 2456
rect 3166 2460 3172 2461
rect 3166 2456 3167 2460
rect 3171 2456 3172 2460
rect 3166 2455 3172 2456
rect 3390 2460 3396 2461
rect 3390 2456 3391 2460
rect 3395 2456 3396 2460
rect 3390 2455 3396 2456
rect 3622 2460 3628 2461
rect 3622 2456 3623 2460
rect 3627 2456 3628 2460
rect 3622 2455 3628 2456
rect 3838 2460 3844 2461
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3838 2455 3844 2456
rect 3942 2457 3948 2458
rect 2046 2452 2052 2453
rect 3942 2453 3943 2457
rect 3947 2453 3948 2457
rect 3942 2452 3948 2453
rect 2146 2451 2152 2452
rect 2146 2447 2147 2451
rect 2151 2447 2152 2451
rect 2146 2446 2152 2447
rect 2290 2451 2296 2452
rect 2290 2447 2291 2451
rect 2295 2447 2296 2451
rect 2290 2446 2296 2447
rect 2298 2451 2304 2452
rect 2298 2447 2299 2451
rect 2303 2450 2304 2451
rect 2470 2451 2476 2452
rect 2303 2448 2425 2450
rect 2303 2447 2304 2448
rect 2298 2446 2304 2447
rect 2470 2447 2471 2451
rect 2475 2450 2476 2451
rect 2642 2451 2648 2452
rect 2475 2448 2601 2450
rect 2475 2447 2476 2448
rect 2470 2446 2476 2447
rect 2642 2447 2643 2451
rect 2647 2450 2648 2451
rect 2898 2451 2904 2452
rect 2647 2448 2793 2450
rect 2647 2447 2648 2448
rect 2642 2446 2648 2447
rect 2898 2447 2899 2451
rect 2903 2450 2904 2451
rect 3034 2451 3040 2452
rect 2903 2448 2993 2450
rect 2903 2447 2904 2448
rect 2898 2446 2904 2447
rect 3034 2447 3035 2451
rect 3039 2450 3040 2451
rect 3255 2451 3261 2452
rect 3039 2448 3209 2450
rect 3039 2447 3040 2448
rect 3034 2446 3040 2447
rect 3255 2447 3256 2451
rect 3260 2450 3261 2451
rect 3698 2451 3704 2452
rect 3260 2448 3433 2450
rect 3260 2447 3261 2448
rect 3255 2446 3261 2447
rect 3698 2447 3699 2451
rect 3703 2447 3704 2451
rect 3698 2446 3704 2447
rect 3906 2451 3912 2452
rect 3906 2447 3907 2451
rect 3911 2447 3912 2451
rect 3906 2446 3912 2447
rect 2070 2441 2076 2442
rect 2046 2440 2052 2441
rect 134 2436 140 2437
rect 110 2433 116 2434
rect 110 2429 111 2433
rect 115 2429 116 2433
rect 134 2432 135 2436
rect 139 2432 140 2436
rect 134 2431 140 2432
rect 310 2436 316 2437
rect 310 2432 311 2436
rect 315 2432 316 2436
rect 310 2431 316 2432
rect 510 2436 516 2437
rect 510 2432 511 2436
rect 515 2432 516 2436
rect 510 2431 516 2432
rect 710 2436 716 2437
rect 710 2432 711 2436
rect 715 2432 716 2436
rect 710 2431 716 2432
rect 902 2436 908 2437
rect 902 2432 903 2436
rect 907 2432 908 2436
rect 902 2431 908 2432
rect 1078 2436 1084 2437
rect 1078 2432 1079 2436
rect 1083 2432 1084 2436
rect 1078 2431 1084 2432
rect 1238 2436 1244 2437
rect 1238 2432 1239 2436
rect 1243 2432 1244 2436
rect 1238 2431 1244 2432
rect 1390 2436 1396 2437
rect 1390 2432 1391 2436
rect 1395 2432 1396 2436
rect 1390 2431 1396 2432
rect 1526 2436 1532 2437
rect 1526 2432 1527 2436
rect 1531 2432 1532 2436
rect 1526 2431 1532 2432
rect 1662 2436 1668 2437
rect 1662 2432 1663 2436
rect 1667 2432 1668 2436
rect 1662 2431 1668 2432
rect 1790 2436 1796 2437
rect 1790 2432 1791 2436
rect 1795 2432 1796 2436
rect 1790 2431 1796 2432
rect 1902 2436 1908 2437
rect 1902 2432 1903 2436
rect 1907 2432 1908 2436
rect 2046 2436 2047 2440
rect 2051 2436 2052 2440
rect 2070 2437 2071 2441
rect 2075 2437 2076 2441
rect 2070 2436 2076 2437
rect 2214 2441 2220 2442
rect 2214 2437 2215 2441
rect 2219 2437 2220 2441
rect 2214 2436 2220 2437
rect 2382 2441 2388 2442
rect 2382 2437 2383 2441
rect 2387 2437 2388 2441
rect 2382 2436 2388 2437
rect 2558 2441 2564 2442
rect 2558 2437 2559 2441
rect 2563 2437 2564 2441
rect 2558 2436 2564 2437
rect 2750 2441 2756 2442
rect 2750 2437 2751 2441
rect 2755 2437 2756 2441
rect 2750 2436 2756 2437
rect 2950 2441 2956 2442
rect 2950 2437 2951 2441
rect 2955 2437 2956 2441
rect 2950 2436 2956 2437
rect 3166 2441 3172 2442
rect 3166 2437 3167 2441
rect 3171 2437 3172 2441
rect 3166 2436 3172 2437
rect 3390 2441 3396 2442
rect 3390 2437 3391 2441
rect 3395 2437 3396 2441
rect 3390 2436 3396 2437
rect 3622 2441 3628 2442
rect 3622 2437 3623 2441
rect 3627 2437 3628 2441
rect 3622 2436 3628 2437
rect 3838 2441 3844 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3942 2440 3948 2441
rect 3942 2436 3943 2440
rect 3947 2436 3948 2440
rect 2046 2435 2052 2436
rect 3942 2435 3948 2436
rect 1902 2431 1908 2432
rect 2006 2433 2012 2434
rect 110 2428 116 2429
rect 1976 2428 2001 2430
rect 2006 2429 2007 2433
rect 2011 2429 2012 2433
rect 2006 2428 2012 2429
rect 210 2427 216 2428
rect 210 2423 211 2427
rect 215 2423 216 2427
rect 210 2422 216 2423
rect 386 2427 392 2428
rect 386 2423 387 2427
rect 391 2423 392 2427
rect 386 2422 392 2423
rect 478 2427 484 2428
rect 478 2423 479 2427
rect 483 2426 484 2427
rect 618 2427 624 2428
rect 483 2424 553 2426
rect 483 2423 484 2424
rect 478 2422 484 2423
rect 618 2423 619 2427
rect 623 2426 624 2427
rect 846 2427 852 2428
rect 623 2424 753 2426
rect 623 2423 624 2424
rect 618 2422 624 2423
rect 846 2423 847 2427
rect 851 2426 852 2427
rect 1154 2427 1160 2428
rect 851 2424 945 2426
rect 851 2423 852 2424
rect 846 2422 852 2423
rect 1154 2423 1155 2427
rect 1159 2423 1160 2427
rect 1154 2422 1160 2423
rect 1314 2427 1320 2428
rect 1314 2423 1315 2427
rect 1319 2423 1320 2427
rect 1314 2422 1320 2423
rect 1466 2427 1472 2428
rect 1466 2423 1467 2427
rect 1471 2423 1472 2427
rect 1466 2422 1472 2423
rect 1474 2427 1480 2428
rect 1474 2423 1475 2427
rect 1479 2426 1480 2427
rect 1738 2427 1744 2428
rect 1479 2424 1569 2426
rect 1479 2423 1480 2424
rect 1474 2422 1480 2423
rect 1738 2423 1739 2427
rect 1743 2423 1744 2427
rect 1738 2422 1744 2423
rect 1866 2427 1872 2428
rect 1866 2423 1867 2427
rect 1871 2423 1872 2427
rect 1976 2425 1978 2428
rect 1866 2422 1872 2423
rect 1999 2422 2001 2428
rect 2107 2423 2113 2424
rect 2107 2422 2108 2423
rect 1999 2420 2108 2422
rect 2107 2419 2108 2420
rect 2112 2419 2113 2423
rect 2107 2418 2113 2419
rect 2146 2423 2152 2424
rect 2146 2419 2147 2423
rect 2151 2422 2152 2423
rect 2251 2423 2257 2424
rect 2251 2422 2252 2423
rect 2151 2420 2252 2422
rect 2151 2419 2152 2420
rect 2146 2418 2152 2419
rect 2251 2419 2252 2420
rect 2256 2419 2257 2423
rect 2251 2418 2257 2419
rect 2290 2423 2296 2424
rect 2290 2419 2291 2423
rect 2295 2422 2296 2423
rect 2419 2423 2425 2424
rect 2419 2422 2420 2423
rect 2295 2420 2420 2422
rect 2295 2419 2296 2420
rect 2290 2418 2296 2419
rect 2419 2419 2420 2420
rect 2424 2419 2425 2423
rect 2419 2418 2425 2419
rect 2595 2423 2601 2424
rect 2595 2419 2596 2423
rect 2600 2422 2601 2423
rect 2642 2423 2648 2424
rect 2642 2422 2643 2423
rect 2600 2420 2643 2422
rect 2600 2419 2601 2420
rect 2595 2418 2601 2419
rect 2642 2419 2643 2420
rect 2647 2419 2648 2423
rect 2642 2418 2648 2419
rect 2787 2423 2793 2424
rect 2787 2419 2788 2423
rect 2792 2422 2793 2423
rect 2898 2423 2904 2424
rect 2898 2422 2899 2423
rect 2792 2420 2899 2422
rect 2792 2419 2793 2420
rect 2787 2418 2793 2419
rect 2898 2419 2899 2420
rect 2903 2419 2904 2423
rect 2898 2418 2904 2419
rect 2987 2423 2993 2424
rect 2987 2419 2988 2423
rect 2992 2422 2993 2423
rect 3034 2423 3040 2424
rect 3034 2422 3035 2423
rect 2992 2420 3035 2422
rect 2992 2419 2993 2420
rect 2987 2418 2993 2419
rect 3034 2419 3035 2420
rect 3039 2419 3040 2423
rect 3034 2418 3040 2419
rect 3203 2423 3209 2424
rect 3203 2419 3204 2423
rect 3208 2422 3209 2423
rect 3255 2423 3261 2424
rect 3255 2422 3256 2423
rect 3208 2420 3256 2422
rect 3208 2419 3209 2420
rect 3203 2418 3209 2419
rect 3255 2419 3256 2420
rect 3260 2419 3261 2423
rect 3255 2418 3261 2419
rect 3427 2423 3433 2424
rect 3427 2419 3428 2423
rect 3432 2422 3433 2423
rect 3450 2423 3456 2424
rect 3450 2422 3451 2423
rect 3432 2420 3451 2422
rect 3432 2419 3433 2420
rect 3427 2418 3433 2419
rect 3450 2419 3451 2420
rect 3455 2419 3456 2423
rect 3875 2423 3881 2424
rect 3450 2418 3456 2419
rect 3659 2419 3665 2420
rect 134 2417 140 2418
rect 110 2416 116 2417
rect 110 2412 111 2416
rect 115 2412 116 2416
rect 134 2413 135 2417
rect 139 2413 140 2417
rect 134 2412 140 2413
rect 310 2417 316 2418
rect 310 2413 311 2417
rect 315 2413 316 2417
rect 310 2412 316 2413
rect 510 2417 516 2418
rect 510 2413 511 2417
rect 515 2413 516 2417
rect 510 2412 516 2413
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 902 2417 908 2418
rect 902 2413 903 2417
rect 907 2413 908 2417
rect 902 2412 908 2413
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1238 2417 1244 2418
rect 1238 2413 1239 2417
rect 1243 2413 1244 2417
rect 1238 2412 1244 2413
rect 1390 2417 1396 2418
rect 1390 2413 1391 2417
rect 1395 2413 1396 2417
rect 1390 2412 1396 2413
rect 1526 2417 1532 2418
rect 1526 2413 1527 2417
rect 1531 2413 1532 2417
rect 1526 2412 1532 2413
rect 1662 2417 1668 2418
rect 1662 2413 1663 2417
rect 1667 2413 1668 2417
rect 1662 2412 1668 2413
rect 1790 2417 1796 2418
rect 1790 2413 1791 2417
rect 1795 2413 1796 2417
rect 1790 2412 1796 2413
rect 1902 2417 1908 2418
rect 1902 2413 1903 2417
rect 1907 2413 1908 2417
rect 1902 2412 1908 2413
rect 2006 2416 2012 2417
rect 2006 2412 2007 2416
rect 2011 2412 2012 2416
rect 3659 2415 3660 2419
rect 3664 2418 3665 2419
rect 3746 2419 3752 2420
rect 3746 2418 3747 2419
rect 3664 2416 3747 2418
rect 3664 2415 3665 2416
rect 3659 2414 3665 2415
rect 3746 2415 3747 2416
rect 3751 2415 3752 2419
rect 3875 2419 3876 2423
rect 3880 2422 3881 2423
rect 3922 2423 3928 2424
rect 3922 2422 3923 2423
rect 3880 2420 3923 2422
rect 3880 2419 3881 2420
rect 3875 2418 3881 2419
rect 3922 2419 3923 2420
rect 3927 2419 3928 2423
rect 3922 2418 3928 2419
rect 3746 2414 3752 2415
rect 110 2411 116 2412
rect 2006 2411 2012 2412
rect 1578 2407 1584 2408
rect 1578 2406 1579 2407
rect 1148 2404 1579 2406
rect 210 2399 216 2400
rect 171 2395 177 2396
rect 171 2391 172 2395
rect 176 2394 177 2395
rect 210 2395 211 2399
rect 215 2398 216 2399
rect 347 2399 353 2400
rect 347 2398 348 2399
rect 215 2396 348 2398
rect 215 2395 216 2396
rect 210 2394 216 2395
rect 347 2395 348 2396
rect 352 2395 353 2399
rect 347 2394 353 2395
rect 386 2399 392 2400
rect 386 2395 387 2399
rect 391 2398 392 2399
rect 547 2399 553 2400
rect 547 2398 548 2399
rect 391 2396 548 2398
rect 391 2395 392 2396
rect 386 2394 392 2395
rect 547 2395 548 2396
rect 552 2395 553 2399
rect 547 2394 553 2395
rect 747 2399 753 2400
rect 747 2395 748 2399
rect 752 2398 753 2399
rect 846 2399 852 2400
rect 846 2398 847 2399
rect 752 2396 847 2398
rect 752 2395 753 2396
rect 747 2394 753 2395
rect 846 2395 847 2396
rect 851 2395 852 2399
rect 846 2394 852 2395
rect 939 2399 945 2400
rect 939 2395 940 2399
rect 944 2398 945 2399
rect 1002 2399 1008 2400
rect 1002 2398 1003 2399
rect 944 2396 1003 2398
rect 944 2395 945 2396
rect 939 2394 945 2395
rect 1002 2395 1003 2396
rect 1007 2395 1008 2399
rect 1002 2394 1008 2395
rect 1115 2399 1121 2400
rect 1115 2395 1116 2399
rect 1120 2398 1121 2399
rect 1148 2398 1150 2404
rect 1578 2403 1579 2404
rect 1583 2403 1584 2407
rect 1578 2402 1584 2403
rect 1120 2396 1150 2398
rect 1154 2399 1160 2400
rect 1120 2395 1121 2396
rect 1115 2394 1121 2395
rect 1154 2395 1155 2399
rect 1159 2398 1160 2399
rect 1275 2399 1281 2400
rect 1275 2398 1276 2399
rect 1159 2396 1276 2398
rect 1159 2395 1160 2396
rect 1154 2394 1160 2395
rect 1275 2395 1276 2396
rect 1280 2395 1281 2399
rect 1275 2394 1281 2395
rect 1314 2399 1320 2400
rect 1314 2395 1315 2399
rect 1319 2398 1320 2399
rect 1427 2399 1433 2400
rect 1427 2398 1428 2399
rect 1319 2396 1428 2398
rect 1319 2395 1320 2396
rect 1314 2394 1320 2395
rect 1427 2395 1428 2396
rect 1432 2395 1433 2399
rect 1427 2394 1433 2395
rect 1466 2399 1472 2400
rect 1466 2395 1467 2399
rect 1471 2398 1472 2399
rect 1563 2399 1569 2400
rect 1563 2398 1564 2399
rect 1471 2396 1564 2398
rect 1471 2395 1472 2396
rect 1466 2394 1472 2395
rect 1563 2395 1564 2396
rect 1568 2395 1569 2399
rect 1738 2399 1744 2400
rect 1563 2394 1569 2395
rect 1699 2395 1705 2396
rect 176 2391 178 2394
rect 171 2390 178 2391
rect 210 2391 216 2392
rect 210 2390 211 2391
rect 176 2388 211 2390
rect 210 2387 211 2388
rect 215 2387 216 2391
rect 1474 2391 1480 2392
rect 1474 2390 1475 2391
rect 210 2386 216 2387
rect 1212 2388 1475 2390
rect 1212 2386 1214 2388
rect 1474 2387 1475 2388
rect 1479 2387 1480 2391
rect 1699 2391 1700 2395
rect 1704 2394 1705 2395
rect 1738 2395 1739 2399
rect 1743 2398 1744 2399
rect 1827 2399 1833 2400
rect 1827 2398 1828 2399
rect 1743 2396 1828 2398
rect 1743 2395 1744 2396
rect 1738 2394 1744 2395
rect 1827 2395 1828 2396
rect 1832 2395 1833 2399
rect 1827 2394 1833 2395
rect 1866 2399 1872 2400
rect 1866 2395 1867 2399
rect 1871 2398 1872 2399
rect 1939 2399 1945 2400
rect 1939 2398 1940 2399
rect 1871 2396 1940 2398
rect 1871 2395 1872 2396
rect 1866 2394 1872 2395
rect 1939 2395 1940 2396
rect 1944 2395 1945 2399
rect 1939 2394 1945 2395
rect 1704 2392 1735 2394
rect 1704 2391 1705 2392
rect 1699 2390 1705 2391
rect 1733 2390 1735 2392
rect 1818 2391 1824 2392
rect 1818 2390 1819 2391
rect 1733 2388 1819 2390
rect 1474 2386 1480 2387
rect 1818 2387 1819 2388
rect 1823 2387 1824 2391
rect 1818 2386 1824 2387
rect 2107 2391 2113 2392
rect 2107 2387 2108 2391
rect 2112 2390 2113 2391
rect 2154 2391 2160 2392
rect 2154 2390 2155 2391
rect 2112 2388 2155 2390
rect 2112 2387 2113 2388
rect 2107 2386 2113 2387
rect 2154 2387 2155 2388
rect 2159 2387 2160 2391
rect 2154 2386 2160 2387
rect 2258 2391 2264 2392
rect 2258 2387 2259 2391
rect 2263 2390 2264 2391
rect 2283 2391 2289 2392
rect 2283 2390 2284 2391
rect 2263 2388 2284 2390
rect 2263 2387 2264 2388
rect 2258 2386 2264 2387
rect 2283 2387 2284 2388
rect 2288 2387 2289 2391
rect 2283 2386 2289 2387
rect 2467 2391 2476 2392
rect 2467 2387 2468 2391
rect 2475 2387 2476 2391
rect 2467 2386 2476 2387
rect 2506 2391 2512 2392
rect 2506 2387 2507 2391
rect 2511 2390 2512 2391
rect 2643 2391 2649 2392
rect 2643 2390 2644 2391
rect 2511 2388 2644 2390
rect 2511 2387 2512 2388
rect 2506 2386 2512 2387
rect 2643 2387 2644 2388
rect 2648 2387 2649 2391
rect 2643 2386 2649 2387
rect 2682 2391 2688 2392
rect 2682 2387 2683 2391
rect 2687 2390 2688 2391
rect 2811 2391 2817 2392
rect 2811 2390 2812 2391
rect 2687 2388 2812 2390
rect 2687 2387 2688 2388
rect 2682 2386 2688 2387
rect 2811 2387 2812 2388
rect 2816 2387 2817 2391
rect 2811 2386 2817 2387
rect 2850 2391 2856 2392
rect 2850 2387 2851 2391
rect 2855 2390 2856 2391
rect 2971 2391 2977 2392
rect 2971 2390 2972 2391
rect 2855 2388 2972 2390
rect 2855 2387 2856 2388
rect 2850 2386 2856 2387
rect 2971 2387 2972 2388
rect 2976 2387 2977 2391
rect 2971 2386 2977 2387
rect 3010 2391 3016 2392
rect 3010 2387 3011 2391
rect 3015 2390 3016 2391
rect 3139 2391 3145 2392
rect 3139 2390 3140 2391
rect 3015 2388 3140 2390
rect 3015 2387 3016 2388
rect 3010 2386 3016 2387
rect 3139 2387 3140 2388
rect 3144 2387 3145 2391
rect 3139 2386 3145 2387
rect 1211 2385 1217 2386
rect 171 2383 177 2384
rect 171 2379 172 2383
rect 176 2382 177 2383
rect 246 2383 252 2384
rect 246 2382 247 2383
rect 176 2380 247 2382
rect 176 2379 177 2380
rect 171 2378 177 2379
rect 246 2379 247 2380
rect 251 2379 252 2383
rect 246 2378 252 2379
rect 346 2383 352 2384
rect 346 2379 347 2383
rect 351 2382 352 2383
rect 363 2383 369 2384
rect 363 2382 364 2383
rect 351 2380 364 2382
rect 351 2379 352 2380
rect 346 2378 352 2379
rect 363 2379 364 2380
rect 368 2379 369 2383
rect 363 2378 369 2379
rect 587 2383 593 2384
rect 587 2379 588 2383
rect 592 2382 593 2383
rect 618 2383 624 2384
rect 618 2382 619 2383
rect 592 2380 619 2382
rect 592 2379 593 2380
rect 587 2378 593 2379
rect 618 2379 619 2380
rect 623 2379 624 2383
rect 618 2378 624 2379
rect 626 2383 632 2384
rect 626 2379 627 2383
rect 631 2382 632 2383
rect 803 2383 809 2384
rect 803 2382 804 2383
rect 631 2380 804 2382
rect 631 2379 632 2380
rect 626 2378 632 2379
rect 803 2379 804 2380
rect 808 2379 809 2383
rect 803 2378 809 2379
rect 842 2383 848 2384
rect 842 2379 843 2383
rect 847 2382 848 2383
rect 1011 2383 1017 2384
rect 1011 2382 1012 2383
rect 847 2380 1012 2382
rect 847 2379 848 2380
rect 842 2378 848 2379
rect 1011 2379 1012 2380
rect 1016 2379 1017 2383
rect 1211 2381 1212 2385
rect 1216 2381 1217 2385
rect 1211 2380 1217 2381
rect 1250 2383 1256 2384
rect 1011 2378 1017 2379
rect 1250 2379 1251 2383
rect 1255 2382 1256 2383
rect 1403 2383 1409 2384
rect 1403 2382 1404 2383
rect 1255 2380 1404 2382
rect 1255 2379 1256 2380
rect 1250 2378 1256 2379
rect 1403 2379 1404 2380
rect 1408 2379 1409 2383
rect 1403 2378 1409 2379
rect 1442 2383 1448 2384
rect 1442 2379 1443 2383
rect 1447 2382 1448 2383
rect 1587 2383 1593 2384
rect 1587 2382 1588 2383
rect 1447 2380 1588 2382
rect 1447 2379 1448 2380
rect 1442 2378 1448 2379
rect 1587 2379 1588 2380
rect 1592 2379 1593 2383
rect 1587 2378 1593 2379
rect 1626 2383 1632 2384
rect 1626 2379 1627 2383
rect 1631 2382 1632 2383
rect 1771 2383 1777 2384
rect 1771 2382 1772 2383
rect 1631 2380 1772 2382
rect 1631 2379 1632 2380
rect 1626 2378 1632 2379
rect 1771 2379 1772 2380
rect 1776 2379 1777 2383
rect 1771 2378 1777 2379
rect 1939 2383 1945 2384
rect 1939 2379 1940 2383
rect 1944 2382 1945 2383
rect 2054 2383 2060 2384
rect 2054 2382 2055 2383
rect 1944 2380 2055 2382
rect 1944 2379 1945 2380
rect 1939 2378 1945 2379
rect 2054 2379 2055 2380
rect 2059 2379 2060 2383
rect 2054 2378 2060 2379
rect 2046 2372 2052 2373
rect 3942 2372 3948 2373
rect 2046 2368 2047 2372
rect 2051 2368 2052 2372
rect 2046 2367 2052 2368
rect 2070 2371 2076 2372
rect 2070 2367 2071 2371
rect 2075 2367 2076 2371
rect 2070 2366 2076 2367
rect 2246 2371 2252 2372
rect 2246 2367 2247 2371
rect 2251 2367 2252 2371
rect 2246 2366 2252 2367
rect 2430 2371 2436 2372
rect 2430 2367 2431 2371
rect 2435 2367 2436 2371
rect 2430 2366 2436 2367
rect 2606 2371 2612 2372
rect 2606 2367 2607 2371
rect 2611 2367 2612 2371
rect 2606 2366 2612 2367
rect 2774 2371 2780 2372
rect 2774 2367 2775 2371
rect 2779 2367 2780 2371
rect 2774 2366 2780 2367
rect 2934 2371 2940 2372
rect 2934 2367 2935 2371
rect 2939 2367 2940 2371
rect 2934 2366 2940 2367
rect 3102 2371 3108 2372
rect 3102 2367 3103 2371
rect 3107 2367 3108 2371
rect 3942 2368 3943 2372
rect 3947 2368 3948 2372
rect 3942 2367 3948 2368
rect 3102 2366 3108 2367
rect 110 2364 116 2365
rect 2006 2364 2012 2365
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 110 2359 116 2360
rect 134 2363 140 2364
rect 134 2359 135 2363
rect 139 2359 140 2363
rect 134 2358 140 2359
rect 326 2363 332 2364
rect 326 2359 327 2363
rect 331 2359 332 2363
rect 326 2358 332 2359
rect 550 2363 556 2364
rect 550 2359 551 2363
rect 555 2359 556 2363
rect 550 2358 556 2359
rect 766 2363 772 2364
rect 766 2359 767 2363
rect 771 2359 772 2363
rect 766 2358 772 2359
rect 974 2363 980 2364
rect 974 2359 975 2363
rect 979 2359 980 2363
rect 974 2358 980 2359
rect 1174 2363 1180 2364
rect 1174 2359 1175 2363
rect 1179 2359 1180 2363
rect 1174 2358 1180 2359
rect 1366 2363 1372 2364
rect 1366 2359 1367 2363
rect 1371 2359 1372 2363
rect 1366 2358 1372 2359
rect 1550 2363 1556 2364
rect 1550 2359 1551 2363
rect 1555 2359 1556 2363
rect 1550 2358 1556 2359
rect 1734 2363 1740 2364
rect 1734 2359 1735 2363
rect 1739 2359 1740 2363
rect 1734 2358 1740 2359
rect 1902 2363 1908 2364
rect 1902 2359 1903 2363
rect 1907 2359 1908 2363
rect 2006 2360 2007 2364
rect 2011 2360 2012 2364
rect 2006 2359 2012 2360
rect 2054 2363 2060 2364
rect 2054 2359 2055 2363
rect 2059 2362 2060 2363
rect 2154 2363 2160 2364
rect 2059 2360 2113 2362
rect 2059 2359 2060 2360
rect 1902 2358 1908 2359
rect 2054 2358 2060 2359
rect 2154 2359 2155 2363
rect 2159 2362 2160 2363
rect 2506 2363 2512 2364
rect 2159 2360 2289 2362
rect 2159 2359 2160 2360
rect 2154 2358 2160 2359
rect 2506 2359 2507 2363
rect 2511 2359 2512 2363
rect 2506 2358 2512 2359
rect 2682 2363 2688 2364
rect 2682 2359 2683 2363
rect 2687 2359 2688 2363
rect 2682 2358 2688 2359
rect 2850 2363 2856 2364
rect 2850 2359 2851 2363
rect 2855 2359 2856 2363
rect 2850 2358 2856 2359
rect 3010 2363 3016 2364
rect 3010 2359 3011 2363
rect 3015 2359 3016 2363
rect 3010 2358 3016 2359
rect 3018 2363 3024 2364
rect 3018 2359 3019 2363
rect 3023 2362 3024 2363
rect 3023 2360 3145 2362
rect 3023 2359 3024 2360
rect 3018 2358 3024 2359
rect 210 2355 216 2356
rect 210 2351 211 2355
rect 215 2351 216 2355
rect 210 2350 216 2351
rect 246 2355 252 2356
rect 246 2351 247 2355
rect 251 2354 252 2355
rect 626 2355 632 2356
rect 251 2352 369 2354
rect 251 2351 252 2352
rect 246 2350 252 2351
rect 626 2351 627 2355
rect 631 2351 632 2355
rect 626 2350 632 2351
rect 842 2355 848 2356
rect 842 2351 843 2355
rect 847 2351 848 2355
rect 842 2350 848 2351
rect 966 2355 972 2356
rect 966 2351 967 2355
rect 971 2354 972 2355
rect 1250 2355 1256 2356
rect 971 2352 1017 2354
rect 971 2351 972 2352
rect 966 2350 972 2351
rect 1250 2351 1251 2355
rect 1255 2351 1256 2355
rect 1250 2350 1256 2351
rect 1442 2355 1448 2356
rect 1442 2351 1443 2355
rect 1447 2351 1448 2355
rect 1442 2350 1448 2351
rect 1626 2355 1632 2356
rect 1626 2351 1627 2355
rect 1631 2351 1632 2355
rect 1626 2350 1632 2351
rect 1670 2355 1676 2356
rect 1670 2351 1671 2355
rect 1675 2354 1676 2355
rect 1818 2355 1824 2356
rect 1675 2352 1777 2354
rect 1675 2351 1676 2352
rect 1670 2350 1676 2351
rect 1818 2351 1819 2355
rect 1823 2354 1824 2355
rect 2046 2355 2052 2356
rect 1823 2352 1945 2354
rect 1823 2351 1824 2352
rect 1818 2350 1824 2351
rect 2046 2351 2047 2355
rect 2051 2351 2052 2355
rect 3942 2355 3948 2356
rect 2046 2350 2052 2351
rect 2070 2352 2076 2353
rect 2070 2348 2071 2352
rect 2075 2348 2076 2352
rect 110 2347 116 2348
rect 110 2343 111 2347
rect 115 2343 116 2347
rect 2006 2347 2012 2348
rect 2070 2347 2076 2348
rect 2246 2352 2252 2353
rect 2246 2348 2247 2352
rect 2251 2348 2252 2352
rect 2246 2347 2252 2348
rect 2430 2352 2436 2353
rect 2430 2348 2431 2352
rect 2435 2348 2436 2352
rect 2430 2347 2436 2348
rect 2606 2352 2612 2353
rect 2606 2348 2607 2352
rect 2611 2348 2612 2352
rect 2606 2347 2612 2348
rect 2774 2352 2780 2353
rect 2774 2348 2775 2352
rect 2779 2348 2780 2352
rect 2774 2347 2780 2348
rect 2934 2352 2940 2353
rect 2934 2348 2935 2352
rect 2939 2348 2940 2352
rect 2934 2347 2940 2348
rect 3102 2352 3108 2353
rect 3102 2348 3103 2352
rect 3107 2348 3108 2352
rect 3942 2351 3943 2355
rect 3947 2351 3948 2355
rect 3942 2350 3948 2351
rect 3102 2347 3108 2348
rect 110 2342 116 2343
rect 134 2344 140 2345
rect 134 2340 135 2344
rect 139 2340 140 2344
rect 134 2339 140 2340
rect 326 2344 332 2345
rect 326 2340 327 2344
rect 331 2340 332 2344
rect 326 2339 332 2340
rect 550 2344 556 2345
rect 550 2340 551 2344
rect 555 2340 556 2344
rect 550 2339 556 2340
rect 766 2344 772 2345
rect 766 2340 767 2344
rect 771 2340 772 2344
rect 766 2339 772 2340
rect 974 2344 980 2345
rect 974 2340 975 2344
rect 979 2340 980 2344
rect 974 2339 980 2340
rect 1174 2344 1180 2345
rect 1174 2340 1175 2344
rect 1179 2340 1180 2344
rect 1174 2339 1180 2340
rect 1366 2344 1372 2345
rect 1366 2340 1367 2344
rect 1371 2340 1372 2344
rect 1366 2339 1372 2340
rect 1550 2344 1556 2345
rect 1550 2340 1551 2344
rect 1555 2340 1556 2344
rect 1550 2339 1556 2340
rect 1734 2344 1740 2345
rect 1734 2340 1735 2344
rect 1739 2340 1740 2344
rect 1734 2339 1740 2340
rect 1902 2344 1908 2345
rect 1902 2340 1903 2344
rect 1907 2340 1908 2344
rect 2006 2343 2007 2347
rect 2011 2343 2012 2347
rect 2006 2342 2012 2343
rect 1902 2339 1908 2340
rect 2070 2292 2076 2293
rect 2046 2289 2052 2290
rect 2046 2285 2047 2289
rect 2051 2285 2052 2289
rect 2070 2288 2071 2292
rect 2075 2288 2076 2292
rect 2070 2287 2076 2288
rect 2174 2292 2180 2293
rect 2174 2288 2175 2292
rect 2179 2288 2180 2292
rect 2174 2287 2180 2288
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2446 2292 2452 2293
rect 2446 2288 2447 2292
rect 2451 2288 2452 2292
rect 2446 2287 2452 2288
rect 2590 2292 2596 2293
rect 2590 2288 2591 2292
rect 2595 2288 2596 2292
rect 2590 2287 2596 2288
rect 2750 2292 2756 2293
rect 2750 2288 2751 2292
rect 2755 2288 2756 2292
rect 2750 2287 2756 2288
rect 2934 2292 2940 2293
rect 2934 2288 2935 2292
rect 2939 2288 2940 2292
rect 2934 2287 2940 2288
rect 3142 2292 3148 2293
rect 3142 2288 3143 2292
rect 3147 2288 3148 2292
rect 3142 2287 3148 2288
rect 3374 2292 3380 2293
rect 3374 2288 3375 2292
rect 3379 2288 3380 2292
rect 3374 2287 3380 2288
rect 3614 2292 3620 2293
rect 3614 2288 3615 2292
rect 3619 2288 3620 2292
rect 3614 2287 3620 2288
rect 3838 2292 3844 2293
rect 3838 2288 3839 2292
rect 3843 2288 3844 2292
rect 3838 2287 3844 2288
rect 3942 2289 3948 2290
rect 2046 2284 2052 2285
rect 3942 2285 3943 2289
rect 3947 2285 3948 2289
rect 3942 2284 3948 2285
rect 2146 2283 2152 2284
rect 2146 2279 2147 2283
rect 2151 2279 2152 2283
rect 2258 2283 2264 2284
rect 2258 2282 2259 2283
rect 2253 2280 2259 2282
rect 2146 2278 2152 2279
rect 2258 2279 2259 2280
rect 2263 2279 2264 2283
rect 2258 2278 2264 2279
rect 2266 2283 2272 2284
rect 2266 2279 2267 2283
rect 2271 2282 2272 2283
rect 2522 2283 2528 2284
rect 2271 2280 2353 2282
rect 2271 2279 2272 2280
rect 2266 2278 2272 2279
rect 2522 2279 2523 2283
rect 2527 2279 2528 2283
rect 2522 2278 2528 2279
rect 2530 2283 2536 2284
rect 2530 2279 2531 2283
rect 2535 2282 2536 2283
rect 2826 2283 2832 2284
rect 2535 2280 2633 2282
rect 2535 2279 2536 2280
rect 2530 2278 2536 2279
rect 2826 2279 2827 2283
rect 2831 2279 2832 2283
rect 2826 2278 2832 2279
rect 3010 2283 3016 2284
rect 3010 2279 3011 2283
rect 3015 2279 3016 2283
rect 3010 2278 3016 2279
rect 3218 2283 3224 2284
rect 3218 2279 3219 2283
rect 3223 2279 3224 2283
rect 3218 2278 3224 2279
rect 3450 2283 3456 2284
rect 3450 2279 3451 2283
rect 3455 2279 3456 2283
rect 3450 2278 3456 2279
rect 3506 2283 3512 2284
rect 3506 2279 3507 2283
rect 3511 2282 3512 2283
rect 3914 2283 3920 2284
rect 3511 2280 3657 2282
rect 3511 2279 3512 2280
rect 3506 2278 3512 2279
rect 3914 2279 3915 2283
rect 3919 2279 3920 2283
rect 3914 2278 3920 2279
rect 134 2276 140 2277
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 134 2272 135 2276
rect 139 2272 140 2276
rect 134 2271 140 2272
rect 270 2276 276 2277
rect 270 2272 271 2276
rect 275 2272 276 2276
rect 270 2271 276 2272
rect 430 2276 436 2277
rect 430 2272 431 2276
rect 435 2272 436 2276
rect 430 2271 436 2272
rect 590 2276 596 2277
rect 590 2272 591 2276
rect 595 2272 596 2276
rect 590 2271 596 2272
rect 750 2276 756 2277
rect 750 2272 751 2276
rect 755 2272 756 2276
rect 750 2271 756 2272
rect 918 2276 924 2277
rect 918 2272 919 2276
rect 923 2272 924 2276
rect 918 2271 924 2272
rect 1086 2276 1092 2277
rect 1086 2272 1087 2276
rect 1091 2272 1092 2276
rect 1086 2271 1092 2272
rect 1262 2276 1268 2277
rect 1262 2272 1263 2276
rect 1267 2272 1268 2276
rect 1262 2271 1268 2272
rect 1446 2276 1452 2277
rect 1446 2272 1447 2276
rect 1451 2272 1452 2276
rect 1446 2271 1452 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1814 2271 1820 2272
rect 2006 2273 2012 2274
rect 2070 2273 2076 2274
rect 110 2268 116 2269
rect 2006 2269 2007 2273
rect 2011 2269 2012 2273
rect 2006 2268 2012 2269
rect 2046 2272 2052 2273
rect 2046 2268 2047 2272
rect 2051 2268 2052 2272
rect 2070 2269 2071 2273
rect 2075 2269 2076 2273
rect 2070 2268 2076 2269
rect 2174 2273 2180 2274
rect 2174 2269 2175 2273
rect 2179 2269 2180 2273
rect 2174 2268 2180 2269
rect 2310 2273 2316 2274
rect 2310 2269 2311 2273
rect 2315 2269 2316 2273
rect 2310 2268 2316 2269
rect 2446 2273 2452 2274
rect 2446 2269 2447 2273
rect 2451 2269 2452 2273
rect 2446 2268 2452 2269
rect 2590 2273 2596 2274
rect 2590 2269 2591 2273
rect 2595 2269 2596 2273
rect 2590 2268 2596 2269
rect 2750 2273 2756 2274
rect 2750 2269 2751 2273
rect 2755 2269 2756 2273
rect 2750 2268 2756 2269
rect 2934 2273 2940 2274
rect 2934 2269 2935 2273
rect 2939 2269 2940 2273
rect 2934 2268 2940 2269
rect 3142 2273 3148 2274
rect 3142 2269 3143 2273
rect 3147 2269 3148 2273
rect 3142 2268 3148 2269
rect 3374 2273 3380 2274
rect 3374 2269 3375 2273
rect 3379 2269 3380 2273
rect 3374 2268 3380 2269
rect 3614 2273 3620 2274
rect 3614 2269 3615 2273
rect 3619 2269 3620 2273
rect 3614 2268 3620 2269
rect 3838 2273 3844 2274
rect 3838 2269 3839 2273
rect 3843 2269 3844 2273
rect 3838 2268 3844 2269
rect 3942 2272 3948 2273
rect 3942 2268 3943 2272
rect 3947 2268 3948 2272
rect 210 2267 216 2268
rect 210 2263 211 2267
rect 215 2263 216 2267
rect 210 2262 216 2263
rect 346 2267 352 2268
rect 346 2263 347 2267
rect 351 2263 352 2267
rect 346 2262 352 2263
rect 378 2267 384 2268
rect 378 2263 379 2267
rect 383 2266 384 2267
rect 666 2267 672 2268
rect 383 2264 473 2266
rect 383 2263 384 2264
rect 378 2262 384 2263
rect 666 2263 667 2267
rect 671 2263 672 2267
rect 666 2262 672 2263
rect 734 2267 740 2268
rect 734 2263 735 2267
rect 739 2266 740 2267
rect 994 2267 1000 2268
rect 739 2264 793 2266
rect 739 2263 740 2264
rect 734 2262 740 2263
rect 994 2263 995 2267
rect 999 2263 1000 2267
rect 994 2262 1000 2263
rect 1162 2267 1168 2268
rect 1162 2263 1163 2267
rect 1167 2263 1168 2267
rect 1162 2262 1168 2263
rect 1338 2267 1344 2268
rect 1338 2263 1339 2267
rect 1343 2263 1344 2267
rect 1338 2262 1344 2263
rect 1522 2267 1528 2268
rect 1522 2263 1523 2267
rect 1527 2263 1528 2267
rect 1522 2262 1528 2263
rect 1706 2267 1712 2268
rect 1706 2263 1707 2267
rect 1711 2263 1712 2267
rect 1706 2262 1712 2263
rect 1882 2267 1888 2268
rect 2046 2267 2052 2268
rect 3942 2267 3948 2268
rect 1882 2263 1883 2267
rect 1887 2263 1888 2267
rect 1882 2262 1888 2263
rect 2266 2263 2272 2264
rect 2266 2262 2267 2263
rect 2140 2260 2267 2262
rect 134 2257 140 2258
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 134 2253 135 2257
rect 139 2253 140 2257
rect 134 2252 140 2253
rect 270 2257 276 2258
rect 270 2253 271 2257
rect 275 2253 276 2257
rect 270 2252 276 2253
rect 430 2257 436 2258
rect 430 2253 431 2257
rect 435 2253 436 2257
rect 430 2252 436 2253
rect 590 2257 596 2258
rect 590 2253 591 2257
rect 595 2253 596 2257
rect 590 2252 596 2253
rect 750 2257 756 2258
rect 750 2253 751 2257
rect 755 2253 756 2257
rect 750 2252 756 2253
rect 918 2257 924 2258
rect 918 2253 919 2257
rect 923 2253 924 2257
rect 918 2252 924 2253
rect 1086 2257 1092 2258
rect 1086 2253 1087 2257
rect 1091 2253 1092 2257
rect 1086 2252 1092 2253
rect 1262 2257 1268 2258
rect 1262 2253 1263 2257
rect 1267 2253 1268 2257
rect 1262 2252 1268 2253
rect 1446 2257 1452 2258
rect 1446 2253 1447 2257
rect 1451 2253 1452 2257
rect 1446 2252 1452 2253
rect 1630 2257 1636 2258
rect 1630 2253 1631 2257
rect 1635 2253 1636 2257
rect 1630 2252 1636 2253
rect 1814 2257 1820 2258
rect 1814 2253 1815 2257
rect 1819 2253 1820 2257
rect 1814 2252 1820 2253
rect 2006 2256 2012 2257
rect 2006 2252 2007 2256
rect 2011 2252 2012 2256
rect 110 2251 116 2252
rect 2006 2251 2012 2252
rect 2107 2255 2113 2256
rect 2107 2251 2108 2255
rect 2112 2254 2113 2255
rect 2140 2254 2142 2260
rect 2266 2259 2267 2260
rect 2271 2259 2272 2263
rect 2530 2263 2536 2264
rect 2530 2262 2531 2263
rect 2266 2258 2272 2259
rect 2464 2260 2531 2262
rect 2112 2252 2142 2254
rect 2146 2255 2152 2256
rect 2112 2251 2113 2252
rect 2107 2250 2113 2251
rect 2146 2251 2147 2255
rect 2151 2254 2152 2255
rect 2211 2255 2217 2256
rect 2211 2254 2212 2255
rect 2151 2252 2212 2254
rect 2151 2251 2152 2252
rect 2146 2250 2152 2251
rect 2211 2251 2212 2252
rect 2216 2251 2217 2255
rect 2211 2250 2217 2251
rect 2347 2255 2353 2256
rect 2347 2251 2348 2255
rect 2352 2254 2353 2255
rect 2464 2254 2466 2260
rect 2530 2259 2531 2260
rect 2535 2259 2536 2263
rect 3018 2263 3024 2264
rect 3018 2262 3019 2263
rect 2530 2258 2536 2259
rect 2839 2260 3019 2262
rect 2839 2258 2841 2260
rect 3018 2259 3019 2260
rect 3023 2259 3024 2263
rect 3018 2258 3024 2259
rect 2796 2256 2841 2258
rect 2352 2252 2466 2254
rect 2522 2255 2528 2256
rect 2352 2251 2353 2252
rect 2347 2250 2353 2251
rect 2482 2251 2489 2252
rect 378 2247 384 2248
rect 378 2246 379 2247
rect 204 2244 379 2246
rect 171 2239 177 2240
rect 171 2235 172 2239
rect 176 2238 177 2239
rect 204 2238 206 2244
rect 378 2243 379 2244
rect 383 2243 384 2247
rect 2482 2247 2483 2251
rect 2488 2247 2489 2251
rect 2522 2251 2523 2255
rect 2527 2254 2528 2255
rect 2627 2255 2633 2256
rect 2627 2254 2628 2255
rect 2527 2252 2628 2254
rect 2527 2251 2528 2252
rect 2522 2250 2528 2251
rect 2627 2251 2628 2252
rect 2632 2251 2633 2255
rect 2627 2250 2633 2251
rect 2787 2255 2793 2256
rect 2787 2251 2788 2255
rect 2792 2254 2793 2255
rect 2796 2254 2798 2256
rect 2971 2255 2977 2256
rect 2971 2254 2972 2255
rect 2792 2252 2798 2254
rect 2839 2252 2972 2254
rect 2792 2251 2793 2252
rect 2787 2250 2793 2251
rect 2826 2251 2832 2252
rect 2482 2246 2489 2247
rect 2826 2247 2827 2251
rect 2831 2250 2832 2251
rect 2839 2250 2841 2252
rect 2971 2251 2972 2252
rect 2976 2251 2977 2255
rect 2971 2250 2977 2251
rect 3010 2255 3016 2256
rect 3010 2251 3011 2255
rect 3015 2254 3016 2255
rect 3179 2255 3185 2256
rect 3179 2254 3180 2255
rect 3015 2252 3180 2254
rect 3015 2251 3016 2252
rect 3010 2250 3016 2251
rect 3179 2251 3180 2252
rect 3184 2251 3185 2255
rect 3179 2250 3185 2251
rect 3218 2255 3224 2256
rect 3218 2251 3219 2255
rect 3223 2254 3224 2255
rect 3411 2255 3417 2256
rect 3411 2254 3412 2255
rect 3223 2252 3412 2254
rect 3223 2251 3224 2252
rect 3218 2250 3224 2251
rect 3411 2251 3412 2252
rect 3416 2251 3417 2255
rect 3411 2250 3417 2251
rect 3450 2255 3456 2256
rect 3450 2251 3451 2255
rect 3455 2254 3456 2255
rect 3651 2255 3657 2256
rect 3651 2254 3652 2255
rect 3455 2252 3652 2254
rect 3455 2251 3456 2252
rect 3450 2250 3456 2251
rect 3651 2251 3652 2252
rect 3656 2251 3657 2255
rect 3651 2250 3657 2251
rect 3875 2255 3881 2256
rect 3875 2251 3876 2255
rect 3880 2254 3881 2255
rect 3906 2255 3912 2256
rect 3906 2254 3907 2255
rect 3880 2252 3907 2254
rect 3880 2251 3881 2252
rect 3875 2250 3881 2251
rect 3906 2251 3907 2252
rect 3911 2251 3912 2255
rect 3906 2250 3912 2251
rect 2831 2248 2841 2250
rect 2831 2247 2832 2248
rect 2826 2246 2832 2247
rect 378 2242 384 2243
rect 966 2243 972 2244
rect 966 2242 967 2243
rect 880 2240 967 2242
rect 176 2236 206 2238
rect 210 2239 216 2240
rect 176 2235 177 2236
rect 171 2234 177 2235
rect 210 2235 211 2239
rect 215 2238 216 2239
rect 307 2239 313 2240
rect 307 2238 308 2239
rect 215 2236 308 2238
rect 215 2235 216 2236
rect 210 2234 216 2235
rect 307 2235 308 2236
rect 312 2235 313 2239
rect 627 2239 633 2240
rect 307 2234 313 2235
rect 402 2235 408 2236
rect 402 2231 403 2235
rect 407 2234 408 2235
rect 467 2235 473 2236
rect 467 2234 468 2235
rect 407 2232 468 2234
rect 407 2231 408 2232
rect 402 2230 408 2231
rect 467 2231 468 2232
rect 472 2231 473 2235
rect 627 2235 628 2239
rect 632 2238 633 2239
rect 734 2239 740 2240
rect 734 2238 735 2239
rect 632 2236 735 2238
rect 632 2235 633 2236
rect 627 2234 633 2235
rect 734 2235 735 2236
rect 739 2235 740 2239
rect 734 2234 740 2235
rect 787 2239 793 2240
rect 787 2235 788 2239
rect 792 2238 793 2239
rect 880 2238 882 2240
rect 966 2239 967 2240
rect 971 2239 972 2243
rect 966 2238 972 2239
rect 994 2239 1000 2240
rect 792 2236 882 2238
rect 792 2235 793 2236
rect 787 2234 793 2235
rect 955 2235 961 2236
rect 467 2230 473 2231
rect 955 2231 956 2235
rect 960 2234 961 2235
rect 986 2235 992 2236
rect 986 2234 987 2235
rect 960 2232 987 2234
rect 960 2231 961 2232
rect 955 2230 961 2231
rect 986 2231 987 2232
rect 991 2231 992 2235
rect 994 2235 995 2239
rect 999 2238 1000 2239
rect 1123 2239 1129 2240
rect 1123 2238 1124 2239
rect 999 2236 1124 2238
rect 999 2235 1000 2236
rect 994 2234 1000 2235
rect 1123 2235 1124 2236
rect 1128 2235 1129 2239
rect 1123 2234 1129 2235
rect 1162 2239 1168 2240
rect 1162 2235 1163 2239
rect 1167 2238 1168 2239
rect 1299 2239 1305 2240
rect 1299 2238 1300 2239
rect 1167 2236 1300 2238
rect 1167 2235 1168 2236
rect 1162 2234 1168 2235
rect 1299 2235 1300 2236
rect 1304 2235 1305 2239
rect 1299 2234 1305 2235
rect 1338 2239 1344 2240
rect 1338 2235 1339 2239
rect 1343 2238 1344 2239
rect 1483 2239 1489 2240
rect 1483 2238 1484 2239
rect 1343 2236 1484 2238
rect 1343 2235 1344 2236
rect 1338 2234 1344 2235
rect 1483 2235 1484 2236
rect 1488 2235 1489 2239
rect 1483 2234 1489 2235
rect 1667 2239 1676 2240
rect 1667 2235 1668 2239
rect 1675 2235 1676 2239
rect 1667 2234 1676 2235
rect 1706 2239 1712 2240
rect 1706 2235 1707 2239
rect 1711 2238 1712 2239
rect 1851 2239 1857 2240
rect 1851 2238 1852 2239
rect 1711 2236 1852 2238
rect 1711 2235 1712 2236
rect 1706 2234 1712 2235
rect 1851 2235 1852 2236
rect 1856 2235 1857 2239
rect 3506 2239 3512 2240
rect 3506 2238 3507 2239
rect 1851 2234 1857 2235
rect 2916 2236 3507 2238
rect 2916 2234 2918 2236
rect 3506 2235 3507 2236
rect 3511 2235 3512 2239
rect 3506 2234 3512 2235
rect 2915 2233 2921 2234
rect 986 2230 992 2231
rect 2186 2231 2192 2232
rect 2147 2229 2153 2230
rect 2147 2225 2148 2229
rect 2152 2225 2153 2229
rect 2186 2227 2187 2231
rect 2191 2230 2192 2231
rect 2291 2231 2297 2232
rect 2291 2230 2292 2231
rect 2191 2228 2292 2230
rect 2191 2227 2192 2228
rect 2186 2226 2192 2227
rect 2291 2227 2292 2228
rect 2296 2227 2297 2231
rect 2291 2226 2297 2227
rect 2330 2231 2336 2232
rect 2330 2227 2331 2231
rect 2335 2230 2336 2231
rect 2443 2231 2449 2232
rect 2443 2230 2444 2231
rect 2335 2228 2444 2230
rect 2335 2227 2336 2228
rect 2330 2226 2336 2227
rect 2443 2227 2444 2228
rect 2448 2227 2449 2231
rect 2443 2226 2449 2227
rect 2595 2231 2601 2232
rect 2595 2227 2596 2231
rect 2600 2230 2601 2231
rect 2642 2231 2648 2232
rect 2642 2230 2643 2231
rect 2600 2228 2643 2230
rect 2600 2227 2601 2228
rect 2595 2226 2601 2227
rect 2642 2227 2643 2228
rect 2647 2227 2648 2231
rect 2642 2226 2648 2227
rect 2658 2231 2664 2232
rect 2658 2227 2659 2231
rect 2663 2230 2664 2231
rect 2755 2231 2761 2232
rect 2755 2230 2756 2231
rect 2663 2228 2756 2230
rect 2663 2227 2664 2228
rect 2658 2226 2664 2227
rect 2755 2227 2756 2228
rect 2760 2227 2761 2231
rect 2915 2229 2916 2233
rect 2920 2229 2921 2233
rect 2915 2228 2921 2229
rect 2954 2231 2960 2232
rect 2755 2226 2761 2227
rect 2954 2227 2955 2231
rect 2959 2230 2960 2231
rect 3083 2231 3089 2232
rect 3083 2230 3084 2231
rect 2959 2228 3084 2230
rect 2959 2227 2960 2228
rect 2954 2226 2960 2227
rect 3083 2227 3084 2228
rect 3088 2227 3089 2231
rect 3083 2226 3089 2227
rect 3122 2231 3128 2232
rect 3122 2227 3123 2231
rect 3127 2230 3128 2231
rect 3259 2231 3265 2232
rect 3259 2230 3260 2231
rect 3127 2228 3260 2230
rect 3127 2227 3128 2228
rect 3122 2226 3128 2227
rect 3259 2227 3260 2228
rect 3264 2227 3265 2231
rect 3259 2226 3265 2227
rect 3298 2231 3304 2232
rect 3298 2227 3299 2231
rect 3303 2230 3304 2231
rect 3443 2231 3449 2232
rect 3443 2230 3444 2231
rect 3303 2228 3444 2230
rect 3303 2227 3304 2228
rect 3298 2226 3304 2227
rect 3443 2227 3444 2228
rect 3448 2227 3449 2231
rect 3443 2226 3449 2227
rect 3482 2231 3488 2232
rect 3482 2227 3483 2231
rect 3487 2230 3488 2231
rect 3627 2231 3633 2232
rect 3627 2230 3628 2231
rect 3487 2228 3628 2230
rect 3487 2227 3488 2228
rect 3482 2226 3488 2227
rect 3627 2227 3628 2228
rect 3632 2227 3633 2231
rect 3627 2226 3633 2227
rect 3819 2231 3825 2232
rect 3819 2227 3820 2231
rect 3824 2230 3825 2231
rect 3866 2231 3872 2232
rect 3866 2230 3867 2231
rect 3824 2228 3867 2230
rect 3824 2227 3825 2228
rect 3819 2226 3825 2227
rect 3866 2227 3867 2228
rect 3871 2227 3872 2231
rect 3866 2226 3872 2227
rect 2147 2224 2153 2225
rect 234 2223 240 2224
rect 195 2221 201 2222
rect 195 2217 196 2221
rect 200 2217 201 2221
rect 234 2219 235 2223
rect 239 2222 240 2223
rect 363 2223 369 2224
rect 363 2222 364 2223
rect 239 2220 364 2222
rect 239 2219 240 2220
rect 234 2218 240 2219
rect 363 2219 364 2220
rect 368 2219 369 2223
rect 363 2218 369 2219
rect 531 2223 537 2224
rect 531 2219 532 2223
rect 536 2222 537 2223
rect 562 2223 568 2224
rect 562 2222 563 2223
rect 536 2220 563 2222
rect 536 2219 537 2220
rect 531 2218 537 2219
rect 562 2219 563 2220
rect 567 2219 568 2223
rect 562 2218 568 2219
rect 666 2223 672 2224
rect 666 2219 667 2223
rect 671 2222 672 2223
rect 715 2223 721 2224
rect 715 2222 716 2223
rect 671 2220 716 2222
rect 671 2219 672 2220
rect 666 2218 672 2219
rect 715 2219 716 2220
rect 720 2219 721 2223
rect 715 2218 721 2219
rect 815 2223 821 2224
rect 815 2219 816 2223
rect 820 2222 821 2223
rect 915 2223 921 2224
rect 915 2222 916 2223
rect 820 2220 916 2222
rect 820 2219 821 2220
rect 815 2218 821 2219
rect 915 2219 916 2220
rect 920 2219 921 2223
rect 915 2218 921 2219
rect 1131 2223 1137 2224
rect 1131 2219 1132 2223
rect 1136 2222 1137 2223
rect 1162 2223 1168 2224
rect 1162 2222 1163 2223
rect 1136 2220 1163 2222
rect 1136 2219 1137 2220
rect 1131 2218 1137 2219
rect 1162 2219 1163 2220
rect 1167 2219 1168 2223
rect 1162 2218 1168 2219
rect 1363 2223 1369 2224
rect 1363 2219 1364 2223
rect 1368 2222 1369 2223
rect 1410 2223 1416 2224
rect 1410 2222 1411 2223
rect 1368 2220 1411 2222
rect 1368 2219 1369 2220
rect 1363 2218 1369 2219
rect 1410 2219 1411 2220
rect 1415 2219 1416 2223
rect 1410 2218 1416 2219
rect 1522 2223 1528 2224
rect 1522 2219 1523 2223
rect 1527 2222 1528 2223
rect 1603 2223 1609 2224
rect 1603 2222 1604 2223
rect 1527 2220 1604 2222
rect 1527 2219 1528 2220
rect 1522 2218 1528 2219
rect 1603 2219 1604 2220
rect 1608 2219 1609 2223
rect 1603 2218 1609 2219
rect 1851 2223 1857 2224
rect 1851 2219 1852 2223
rect 1856 2222 1857 2223
rect 1882 2223 1888 2224
rect 1882 2222 1883 2223
rect 1856 2220 1883 2222
rect 1856 2219 1857 2220
rect 1851 2218 1857 2219
rect 1882 2219 1883 2220
rect 1887 2219 1888 2223
rect 2148 2222 2150 2224
rect 2490 2223 2496 2224
rect 2490 2222 2491 2223
rect 2148 2220 2491 2222
rect 1882 2218 1888 2219
rect 2490 2219 2491 2220
rect 2495 2219 2496 2223
rect 2490 2218 2496 2219
rect 195 2216 201 2217
rect 196 2214 198 2216
rect 410 2215 416 2216
rect 410 2214 411 2215
rect 196 2212 411 2214
rect 410 2211 411 2212
rect 415 2211 416 2215
rect 410 2210 416 2211
rect 2046 2212 2052 2213
rect 3942 2212 3948 2213
rect 2046 2208 2047 2212
rect 2051 2208 2052 2212
rect 2046 2207 2052 2208
rect 2110 2211 2116 2212
rect 2110 2207 2111 2211
rect 2115 2207 2116 2211
rect 2110 2206 2116 2207
rect 2254 2211 2260 2212
rect 2254 2207 2255 2211
rect 2259 2207 2260 2211
rect 2254 2206 2260 2207
rect 2406 2211 2412 2212
rect 2406 2207 2407 2211
rect 2411 2207 2412 2211
rect 2406 2206 2412 2207
rect 2558 2211 2564 2212
rect 2558 2207 2559 2211
rect 2563 2207 2564 2211
rect 2558 2206 2564 2207
rect 2718 2211 2724 2212
rect 2718 2207 2719 2211
rect 2723 2207 2724 2211
rect 2718 2206 2724 2207
rect 2878 2211 2884 2212
rect 2878 2207 2879 2211
rect 2883 2207 2884 2211
rect 2878 2206 2884 2207
rect 3046 2211 3052 2212
rect 3046 2207 3047 2211
rect 3051 2207 3052 2211
rect 3046 2206 3052 2207
rect 3222 2211 3228 2212
rect 3222 2207 3223 2211
rect 3227 2207 3228 2211
rect 3222 2206 3228 2207
rect 3406 2211 3412 2212
rect 3406 2207 3407 2211
rect 3411 2207 3412 2211
rect 3406 2206 3412 2207
rect 3590 2211 3596 2212
rect 3590 2207 3591 2211
rect 3595 2207 3596 2211
rect 3590 2206 3596 2207
rect 3782 2211 3788 2212
rect 3782 2207 3783 2211
rect 3787 2207 3788 2211
rect 3942 2208 3943 2212
rect 3947 2208 3948 2212
rect 3942 2207 3948 2208
rect 3782 2206 3788 2207
rect 110 2204 116 2205
rect 2006 2204 2012 2205
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 110 2199 116 2200
rect 158 2203 164 2204
rect 158 2199 159 2203
rect 163 2199 164 2203
rect 158 2198 164 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 678 2203 684 2204
rect 678 2199 679 2203
rect 683 2199 684 2203
rect 678 2198 684 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 1094 2203 1100 2204
rect 1094 2199 1095 2203
rect 1099 2199 1100 2203
rect 1094 2198 1100 2199
rect 1326 2203 1332 2204
rect 1326 2199 1327 2203
rect 1331 2199 1332 2203
rect 1326 2198 1332 2199
rect 1566 2203 1572 2204
rect 1566 2199 1567 2203
rect 1571 2199 1572 2203
rect 1566 2198 1572 2199
rect 1814 2203 1820 2204
rect 1814 2199 1815 2203
rect 1819 2199 1820 2203
rect 2006 2200 2007 2204
rect 2011 2200 2012 2204
rect 2006 2199 2012 2200
rect 2186 2203 2192 2204
rect 2186 2199 2187 2203
rect 2191 2199 2192 2203
rect 1814 2198 1820 2199
rect 2186 2198 2192 2199
rect 2330 2203 2336 2204
rect 2330 2199 2331 2203
rect 2335 2199 2336 2203
rect 2330 2198 2336 2199
rect 2482 2203 2488 2204
rect 2482 2199 2483 2203
rect 2487 2199 2488 2203
rect 2482 2198 2488 2199
rect 2490 2203 2496 2204
rect 2490 2199 2491 2203
rect 2495 2202 2496 2203
rect 2642 2203 2648 2204
rect 2495 2200 2601 2202
rect 2495 2199 2496 2200
rect 2490 2198 2496 2199
rect 2642 2199 2643 2203
rect 2647 2202 2648 2203
rect 2954 2203 2960 2204
rect 2647 2200 2761 2202
rect 2647 2199 2648 2200
rect 2642 2198 2648 2199
rect 2954 2199 2955 2203
rect 2959 2199 2960 2203
rect 2954 2198 2960 2199
rect 3122 2203 3128 2204
rect 3122 2199 3123 2203
rect 3127 2199 3128 2203
rect 3122 2198 3128 2199
rect 3298 2203 3304 2204
rect 3298 2199 3299 2203
rect 3303 2199 3304 2203
rect 3298 2198 3304 2199
rect 3482 2203 3488 2204
rect 3482 2199 3483 2203
rect 3487 2199 3488 2203
rect 3482 2198 3488 2199
rect 3558 2203 3564 2204
rect 3558 2199 3559 2203
rect 3563 2202 3564 2203
rect 3746 2203 3752 2204
rect 3563 2200 3633 2202
rect 3563 2199 3564 2200
rect 3558 2198 3564 2199
rect 3746 2199 3747 2203
rect 3751 2202 3752 2203
rect 3751 2200 3825 2202
rect 3751 2199 3752 2200
rect 3746 2198 3752 2199
rect 234 2195 240 2196
rect 234 2191 235 2195
rect 239 2191 240 2195
rect 234 2190 240 2191
rect 402 2195 408 2196
rect 402 2191 403 2195
rect 407 2191 408 2195
rect 402 2190 408 2191
rect 410 2195 416 2196
rect 410 2191 411 2195
rect 415 2194 416 2195
rect 815 2195 821 2196
rect 815 2194 816 2195
rect 415 2192 537 2194
rect 757 2192 816 2194
rect 415 2191 416 2192
rect 410 2190 416 2191
rect 815 2191 816 2192
rect 820 2191 821 2195
rect 815 2190 821 2191
rect 826 2195 832 2196
rect 826 2191 827 2195
rect 831 2194 832 2195
rect 986 2195 992 2196
rect 831 2192 921 2194
rect 831 2191 832 2192
rect 826 2190 832 2191
rect 986 2191 987 2195
rect 991 2194 992 2195
rect 1302 2195 1308 2196
rect 991 2192 1137 2194
rect 991 2191 992 2192
rect 986 2190 992 2191
rect 1302 2191 1303 2195
rect 1307 2194 1308 2195
rect 1410 2195 1416 2196
rect 1307 2192 1369 2194
rect 1307 2191 1308 2192
rect 1302 2190 1308 2191
rect 1410 2191 1411 2195
rect 1415 2194 1416 2195
rect 2046 2195 2052 2196
rect 1415 2192 1609 2194
rect 1415 2191 1416 2192
rect 1410 2190 1416 2191
rect 1890 2191 1896 2192
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 1890 2187 1891 2191
rect 1895 2187 1896 2191
rect 2046 2191 2047 2195
rect 2051 2191 2052 2195
rect 3942 2195 3948 2196
rect 2046 2190 2052 2191
rect 2110 2192 2116 2193
rect 2110 2188 2111 2192
rect 2115 2188 2116 2192
rect 1890 2186 1896 2187
rect 2006 2187 2012 2188
rect 2110 2187 2116 2188
rect 2254 2192 2260 2193
rect 2254 2188 2255 2192
rect 2259 2188 2260 2192
rect 2254 2187 2260 2188
rect 2406 2192 2412 2193
rect 2406 2188 2407 2192
rect 2411 2188 2412 2192
rect 2406 2187 2412 2188
rect 2558 2192 2564 2193
rect 2558 2188 2559 2192
rect 2563 2188 2564 2192
rect 2558 2187 2564 2188
rect 2718 2192 2724 2193
rect 2718 2188 2719 2192
rect 2723 2188 2724 2192
rect 2718 2187 2724 2188
rect 2878 2192 2884 2193
rect 2878 2188 2879 2192
rect 2883 2188 2884 2192
rect 2878 2187 2884 2188
rect 3046 2192 3052 2193
rect 3046 2188 3047 2192
rect 3051 2188 3052 2192
rect 3046 2187 3052 2188
rect 3222 2192 3228 2193
rect 3222 2188 3223 2192
rect 3227 2188 3228 2192
rect 3222 2187 3228 2188
rect 3406 2192 3412 2193
rect 3406 2188 3407 2192
rect 3411 2188 3412 2192
rect 3406 2187 3412 2188
rect 3590 2192 3596 2193
rect 3590 2188 3591 2192
rect 3595 2188 3596 2192
rect 3590 2187 3596 2188
rect 3782 2192 3788 2193
rect 3782 2188 3783 2192
rect 3787 2188 3788 2192
rect 3942 2191 3943 2195
rect 3947 2191 3948 2195
rect 3942 2190 3948 2191
rect 3782 2187 3788 2188
rect 110 2182 116 2183
rect 158 2184 164 2185
rect 158 2180 159 2184
rect 163 2180 164 2184
rect 158 2179 164 2180
rect 326 2184 332 2185
rect 326 2180 327 2184
rect 331 2180 332 2184
rect 326 2179 332 2180
rect 494 2184 500 2185
rect 494 2180 495 2184
rect 499 2180 500 2184
rect 494 2179 500 2180
rect 678 2184 684 2185
rect 678 2180 679 2184
rect 683 2180 684 2184
rect 678 2179 684 2180
rect 878 2184 884 2185
rect 878 2180 879 2184
rect 883 2180 884 2184
rect 878 2179 884 2180
rect 1094 2184 1100 2185
rect 1094 2180 1095 2184
rect 1099 2180 1100 2184
rect 1094 2179 1100 2180
rect 1326 2184 1332 2185
rect 1326 2180 1327 2184
rect 1331 2180 1332 2184
rect 1326 2179 1332 2180
rect 1566 2184 1572 2185
rect 1566 2180 1567 2184
rect 1571 2180 1572 2184
rect 1566 2179 1572 2180
rect 1814 2184 1820 2185
rect 1814 2180 1815 2184
rect 1819 2180 1820 2184
rect 2006 2183 2007 2187
rect 2011 2183 2012 2187
rect 2006 2182 2012 2183
rect 1814 2179 1820 2180
rect 3086 2143 3092 2144
rect 3086 2139 3087 2143
rect 3091 2142 3092 2143
rect 3558 2143 3564 2144
rect 3558 2142 3559 2143
rect 3091 2140 3559 2142
rect 3091 2139 3092 2140
rect 3086 2138 3092 2139
rect 3558 2139 3559 2140
rect 3563 2139 3564 2143
rect 3558 2138 3564 2139
rect 222 2124 228 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 222 2120 223 2124
rect 227 2120 228 2124
rect 222 2119 228 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 494 2124 500 2125
rect 494 2120 495 2124
rect 499 2120 500 2124
rect 494 2119 500 2120
rect 638 2124 644 2125
rect 638 2120 639 2124
rect 643 2120 644 2124
rect 638 2119 644 2120
rect 782 2124 788 2125
rect 782 2120 783 2124
rect 787 2120 788 2124
rect 782 2119 788 2120
rect 934 2124 940 2125
rect 934 2120 935 2124
rect 939 2120 940 2124
rect 934 2119 940 2120
rect 1094 2124 1100 2125
rect 1094 2120 1095 2124
rect 1099 2120 1100 2124
rect 1094 2119 1100 2120
rect 1262 2124 1268 2125
rect 1262 2120 1263 2124
rect 1267 2120 1268 2124
rect 1262 2119 1268 2120
rect 1446 2124 1452 2125
rect 1446 2120 1447 2124
rect 1451 2120 1452 2124
rect 1446 2119 1452 2120
rect 1630 2124 1636 2125
rect 1630 2120 1631 2124
rect 1635 2120 1636 2124
rect 1630 2119 1636 2120
rect 1822 2124 1828 2125
rect 1822 2120 1823 2124
rect 1827 2120 1828 2124
rect 1822 2119 1828 2120
rect 2006 2121 2012 2122
rect 110 2116 116 2117
rect 2006 2117 2007 2121
rect 2011 2117 2012 2121
rect 2286 2120 2292 2121
rect 2006 2116 2012 2117
rect 2046 2117 2052 2118
rect 298 2115 304 2116
rect 298 2111 299 2115
rect 303 2111 304 2115
rect 298 2110 304 2111
rect 434 2115 440 2116
rect 434 2111 435 2115
rect 439 2111 440 2115
rect 434 2110 440 2111
rect 562 2115 568 2116
rect 562 2111 563 2115
rect 567 2111 568 2115
rect 562 2110 568 2111
rect 578 2115 584 2116
rect 578 2111 579 2115
rect 583 2114 584 2115
rect 775 2115 781 2116
rect 583 2112 681 2114
rect 583 2111 584 2112
rect 578 2110 584 2111
rect 775 2111 776 2115
rect 780 2114 781 2115
rect 1010 2115 1016 2116
rect 780 2112 825 2114
rect 780 2111 781 2112
rect 775 2110 781 2111
rect 1010 2111 1011 2115
rect 1015 2111 1016 2115
rect 1010 2110 1016 2111
rect 1162 2115 1168 2116
rect 1162 2111 1163 2115
rect 1167 2111 1168 2115
rect 1162 2110 1168 2111
rect 1338 2115 1344 2116
rect 1338 2111 1339 2115
rect 1343 2111 1344 2115
rect 1338 2110 1344 2111
rect 1522 2115 1528 2116
rect 1522 2111 1523 2115
rect 1527 2111 1528 2115
rect 1522 2110 1528 2111
rect 1622 2115 1628 2116
rect 1622 2111 1623 2115
rect 1627 2114 1628 2115
rect 1814 2115 1820 2116
rect 1627 2112 1673 2114
rect 1627 2111 1628 2112
rect 1622 2110 1628 2111
rect 1814 2111 1815 2115
rect 1819 2114 1820 2115
rect 1819 2112 1865 2114
rect 2046 2113 2047 2117
rect 2051 2113 2052 2117
rect 2286 2116 2287 2120
rect 2291 2116 2292 2120
rect 2286 2115 2292 2116
rect 2430 2120 2436 2121
rect 2430 2116 2431 2120
rect 2435 2116 2436 2120
rect 2430 2115 2436 2116
rect 2582 2120 2588 2121
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2734 2120 2740 2121
rect 2734 2116 2735 2120
rect 2739 2116 2740 2120
rect 2734 2115 2740 2116
rect 2886 2120 2892 2121
rect 2886 2116 2887 2120
rect 2891 2116 2892 2120
rect 2886 2115 2892 2116
rect 3046 2120 3052 2121
rect 3046 2116 3047 2120
rect 3051 2116 3052 2120
rect 3046 2115 3052 2116
rect 3206 2120 3212 2121
rect 3206 2116 3207 2120
rect 3211 2116 3212 2120
rect 3206 2115 3212 2116
rect 3366 2120 3372 2121
rect 3366 2116 3367 2120
rect 3371 2116 3372 2120
rect 3366 2115 3372 2116
rect 3526 2120 3532 2121
rect 3526 2116 3527 2120
rect 3531 2116 3532 2120
rect 3526 2115 3532 2116
rect 3694 2120 3700 2121
rect 3694 2116 3695 2120
rect 3699 2116 3700 2120
rect 3694 2115 3700 2116
rect 3838 2120 3844 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3838 2115 3844 2116
rect 3942 2117 3948 2118
rect 2046 2112 2052 2113
rect 3942 2113 3943 2117
rect 3947 2113 3948 2117
rect 3942 2112 3948 2113
rect 1819 2111 1820 2112
rect 1814 2110 1820 2111
rect 2362 2111 2368 2112
rect 2362 2107 2363 2111
rect 2367 2107 2368 2111
rect 2362 2106 2368 2107
rect 2506 2111 2512 2112
rect 2506 2107 2507 2111
rect 2511 2107 2512 2111
rect 2506 2106 2512 2107
rect 2658 2111 2664 2112
rect 2658 2107 2659 2111
rect 2663 2107 2664 2111
rect 2658 2106 2664 2107
rect 2666 2111 2672 2112
rect 2666 2107 2667 2111
rect 2671 2110 2672 2111
rect 2818 2111 2824 2112
rect 2671 2108 2777 2110
rect 2671 2107 2672 2108
rect 2666 2106 2672 2107
rect 2818 2107 2819 2111
rect 2823 2110 2824 2111
rect 3122 2111 3128 2112
rect 2823 2108 2929 2110
rect 2823 2107 2824 2108
rect 2818 2106 2824 2107
rect 3122 2107 3123 2111
rect 3127 2107 3128 2111
rect 3122 2106 3128 2107
rect 3282 2111 3288 2112
rect 3282 2107 3283 2111
rect 3287 2107 3288 2111
rect 3282 2106 3288 2107
rect 3442 2111 3448 2112
rect 3442 2107 3443 2111
rect 3447 2107 3448 2111
rect 3442 2106 3448 2107
rect 3602 2111 3608 2112
rect 3602 2107 3603 2111
rect 3607 2107 3608 2111
rect 3602 2106 3608 2107
rect 3618 2111 3624 2112
rect 3618 2107 3619 2111
rect 3623 2110 3624 2111
rect 3906 2111 3912 2112
rect 3623 2108 3737 2110
rect 3623 2107 3624 2108
rect 3618 2106 3624 2107
rect 3906 2107 3907 2111
rect 3911 2107 3912 2111
rect 3906 2106 3912 2107
rect 222 2105 228 2106
rect 110 2104 116 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 222 2101 223 2105
rect 227 2101 228 2105
rect 222 2100 228 2101
rect 358 2105 364 2106
rect 358 2101 359 2105
rect 363 2101 364 2105
rect 358 2100 364 2101
rect 494 2105 500 2106
rect 494 2101 495 2105
rect 499 2101 500 2105
rect 494 2100 500 2101
rect 638 2105 644 2106
rect 638 2101 639 2105
rect 643 2101 644 2105
rect 638 2100 644 2101
rect 782 2105 788 2106
rect 782 2101 783 2105
rect 787 2101 788 2105
rect 782 2100 788 2101
rect 934 2105 940 2106
rect 934 2101 935 2105
rect 939 2101 940 2105
rect 934 2100 940 2101
rect 1094 2105 1100 2106
rect 1094 2101 1095 2105
rect 1099 2101 1100 2105
rect 1094 2100 1100 2101
rect 1262 2105 1268 2106
rect 1262 2101 1263 2105
rect 1267 2101 1268 2105
rect 1262 2100 1268 2101
rect 1446 2105 1452 2106
rect 1446 2101 1447 2105
rect 1451 2101 1452 2105
rect 1446 2100 1452 2101
rect 1630 2105 1636 2106
rect 1630 2101 1631 2105
rect 1635 2101 1636 2105
rect 1630 2100 1636 2101
rect 1822 2105 1828 2106
rect 1822 2101 1823 2105
rect 1827 2101 1828 2105
rect 1822 2100 1828 2101
rect 2006 2104 2012 2105
rect 2006 2100 2007 2104
rect 2011 2100 2012 2104
rect 2286 2101 2292 2102
rect 110 2099 116 2100
rect 2006 2099 2012 2100
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2286 2097 2287 2101
rect 2291 2097 2292 2101
rect 2286 2096 2292 2097
rect 2430 2101 2436 2102
rect 2430 2097 2431 2101
rect 2435 2097 2436 2101
rect 2430 2096 2436 2097
rect 2582 2101 2588 2102
rect 2582 2097 2583 2101
rect 2587 2097 2588 2101
rect 2582 2096 2588 2097
rect 2734 2101 2740 2102
rect 2734 2097 2735 2101
rect 2739 2097 2740 2101
rect 2734 2096 2740 2097
rect 2886 2101 2892 2102
rect 2886 2097 2887 2101
rect 2891 2097 2892 2101
rect 2886 2096 2892 2097
rect 3046 2101 3052 2102
rect 3046 2097 3047 2101
rect 3051 2097 3052 2101
rect 3046 2096 3052 2097
rect 3206 2101 3212 2102
rect 3206 2097 3207 2101
rect 3211 2097 3212 2101
rect 3206 2096 3212 2097
rect 3366 2101 3372 2102
rect 3366 2097 3367 2101
rect 3371 2097 3372 2101
rect 3366 2096 3372 2097
rect 3526 2101 3532 2102
rect 3526 2097 3527 2101
rect 3531 2097 3532 2101
rect 3526 2096 3532 2097
rect 3694 2101 3700 2102
rect 3694 2097 3695 2101
rect 3699 2097 3700 2101
rect 3694 2096 3700 2097
rect 3838 2101 3844 2102
rect 3838 2097 3839 2101
rect 3843 2097 3844 2101
rect 3838 2096 3844 2097
rect 3942 2100 3948 2101
rect 3942 2096 3943 2100
rect 3947 2096 3948 2100
rect 578 2095 584 2096
rect 2046 2095 2052 2096
rect 3942 2095 3948 2096
rect 578 2094 579 2095
rect 319 2092 579 2094
rect 319 2090 321 2092
rect 578 2091 579 2092
rect 583 2091 584 2095
rect 578 2090 584 2091
rect 2666 2091 2672 2092
rect 2666 2090 2667 2091
rect 288 2088 321 2090
rect 2356 2088 2667 2090
rect 259 2087 265 2088
rect 259 2083 260 2087
rect 264 2086 265 2087
rect 288 2086 290 2088
rect 395 2087 401 2088
rect 395 2086 396 2087
rect 264 2084 290 2086
rect 319 2084 396 2086
rect 264 2083 265 2084
rect 259 2082 265 2083
rect 298 2083 304 2084
rect 298 2079 299 2083
rect 303 2082 304 2083
rect 319 2082 321 2084
rect 395 2083 396 2084
rect 400 2083 401 2087
rect 395 2082 401 2083
rect 434 2087 440 2088
rect 434 2083 435 2087
rect 439 2086 440 2087
rect 531 2087 537 2088
rect 531 2086 532 2087
rect 439 2084 532 2086
rect 439 2083 440 2084
rect 434 2082 440 2083
rect 531 2083 532 2084
rect 536 2083 537 2087
rect 819 2087 828 2088
rect 531 2082 537 2083
rect 675 2083 681 2084
rect 303 2080 321 2082
rect 303 2079 304 2080
rect 298 2078 304 2079
rect 675 2079 676 2083
rect 680 2082 681 2083
rect 690 2083 696 2084
rect 690 2082 691 2083
rect 680 2080 691 2082
rect 680 2079 681 2080
rect 675 2078 681 2079
rect 690 2079 691 2080
rect 695 2079 696 2083
rect 819 2083 820 2087
rect 827 2083 828 2087
rect 1010 2087 1016 2088
rect 819 2082 828 2083
rect 971 2083 977 2084
rect 690 2078 696 2079
rect 971 2079 972 2083
rect 976 2082 977 2083
rect 1002 2083 1008 2084
rect 1002 2082 1003 2083
rect 976 2080 1003 2082
rect 976 2079 977 2080
rect 971 2078 977 2079
rect 1002 2079 1003 2080
rect 1007 2079 1008 2083
rect 1010 2083 1011 2087
rect 1015 2086 1016 2087
rect 1131 2087 1137 2088
rect 1131 2086 1132 2087
rect 1015 2084 1132 2086
rect 1015 2083 1016 2084
rect 1010 2082 1016 2083
rect 1131 2083 1132 2084
rect 1136 2083 1137 2087
rect 1131 2082 1137 2083
rect 1299 2087 1308 2088
rect 1299 2083 1300 2087
rect 1307 2083 1308 2087
rect 1299 2082 1308 2083
rect 1338 2087 1344 2088
rect 1338 2083 1339 2087
rect 1343 2086 1344 2087
rect 1483 2087 1489 2088
rect 1483 2086 1484 2087
rect 1343 2084 1484 2086
rect 1343 2083 1344 2084
rect 1338 2082 1344 2083
rect 1483 2083 1484 2084
rect 1488 2083 1489 2087
rect 1483 2082 1489 2083
rect 1522 2087 1528 2088
rect 1522 2083 1523 2087
rect 1527 2086 1528 2087
rect 1667 2087 1673 2088
rect 1667 2086 1668 2087
rect 1527 2084 1668 2086
rect 1527 2083 1528 2084
rect 1522 2082 1528 2083
rect 1667 2083 1668 2084
rect 1672 2083 1673 2087
rect 1667 2082 1673 2083
rect 1859 2087 1865 2088
rect 1859 2083 1860 2087
rect 1864 2086 1865 2087
rect 1890 2087 1896 2088
rect 1890 2086 1891 2087
rect 1864 2084 1891 2086
rect 1864 2083 1865 2084
rect 1859 2082 1865 2083
rect 1890 2083 1891 2084
rect 1895 2083 1896 2087
rect 1890 2082 1896 2083
rect 2323 2083 2329 2084
rect 1002 2078 1008 2079
rect 2323 2079 2324 2083
rect 2328 2082 2329 2083
rect 2356 2082 2358 2088
rect 2666 2087 2667 2088
rect 2671 2087 2672 2091
rect 2666 2086 2672 2087
rect 2328 2080 2358 2082
rect 2362 2083 2368 2084
rect 2328 2079 2329 2080
rect 2323 2078 2329 2079
rect 2362 2079 2363 2083
rect 2367 2082 2368 2083
rect 2467 2083 2473 2084
rect 2467 2082 2468 2083
rect 2367 2080 2468 2082
rect 2367 2079 2368 2080
rect 2362 2078 2368 2079
rect 2467 2079 2468 2080
rect 2472 2079 2473 2083
rect 2467 2078 2473 2079
rect 2506 2083 2512 2084
rect 2506 2079 2507 2083
rect 2511 2082 2512 2083
rect 2619 2083 2625 2084
rect 2619 2082 2620 2083
rect 2511 2080 2620 2082
rect 2511 2079 2512 2080
rect 2506 2078 2512 2079
rect 2619 2079 2620 2080
rect 2624 2079 2625 2083
rect 2619 2078 2625 2079
rect 2771 2083 2777 2084
rect 2771 2079 2772 2083
rect 2776 2082 2777 2083
rect 2818 2083 2824 2084
rect 2818 2082 2819 2083
rect 2776 2080 2819 2082
rect 2776 2079 2777 2080
rect 2771 2078 2777 2079
rect 2818 2079 2819 2080
rect 2823 2079 2824 2083
rect 3083 2083 3092 2084
rect 2818 2078 2824 2079
rect 2923 2079 2932 2080
rect 2923 2075 2924 2079
rect 2931 2075 2932 2079
rect 3083 2079 3084 2083
rect 3091 2079 3092 2083
rect 3083 2078 3092 2079
rect 3122 2083 3128 2084
rect 3122 2079 3123 2083
rect 3127 2082 3128 2083
rect 3243 2083 3249 2084
rect 3243 2082 3244 2083
rect 3127 2080 3244 2082
rect 3127 2079 3128 2080
rect 3122 2078 3128 2079
rect 3243 2079 3244 2080
rect 3248 2079 3249 2083
rect 3243 2078 3249 2079
rect 3282 2083 3288 2084
rect 3282 2079 3283 2083
rect 3287 2082 3288 2083
rect 3403 2083 3409 2084
rect 3403 2082 3404 2083
rect 3287 2080 3404 2082
rect 3287 2079 3288 2080
rect 3282 2078 3288 2079
rect 3403 2079 3404 2080
rect 3408 2079 3409 2083
rect 3403 2078 3409 2079
rect 3442 2083 3448 2084
rect 3442 2079 3443 2083
rect 3447 2082 3448 2083
rect 3563 2083 3569 2084
rect 3563 2082 3564 2083
rect 3447 2080 3564 2082
rect 3447 2079 3448 2080
rect 3442 2078 3448 2079
rect 3563 2079 3564 2080
rect 3568 2079 3569 2083
rect 3563 2078 3569 2079
rect 3602 2083 3608 2084
rect 3602 2079 3603 2083
rect 3607 2082 3608 2083
rect 3731 2083 3737 2084
rect 3731 2082 3732 2083
rect 3607 2080 3732 2082
rect 3607 2079 3608 2080
rect 3602 2078 3608 2079
rect 3731 2079 3732 2080
rect 3736 2079 3737 2083
rect 3731 2078 3737 2079
rect 3875 2083 3881 2084
rect 3875 2079 3876 2083
rect 3880 2082 3881 2083
rect 3914 2083 3920 2084
rect 3914 2082 3915 2083
rect 3880 2080 3915 2082
rect 3880 2079 3881 2080
rect 3875 2078 3881 2079
rect 3914 2079 3915 2080
rect 3919 2079 3920 2083
rect 3914 2078 3920 2079
rect 2923 2074 2932 2075
rect 3618 2067 3624 2068
rect 3618 2066 3619 2067
rect 3204 2064 3619 2066
rect 411 2063 420 2064
rect 411 2059 412 2063
rect 419 2059 420 2063
rect 411 2058 420 2059
rect 450 2063 456 2064
rect 450 2059 451 2063
rect 455 2062 456 2063
rect 531 2063 537 2064
rect 531 2062 532 2063
rect 455 2060 532 2062
rect 455 2059 456 2060
rect 450 2058 456 2059
rect 531 2059 532 2060
rect 536 2059 537 2063
rect 531 2058 537 2059
rect 570 2063 576 2064
rect 570 2059 571 2063
rect 575 2062 576 2063
rect 651 2063 657 2064
rect 651 2062 652 2063
rect 575 2060 652 2062
rect 575 2059 576 2060
rect 570 2058 576 2059
rect 651 2059 652 2060
rect 656 2059 657 2063
rect 651 2058 657 2059
rect 775 2063 781 2064
rect 775 2059 776 2063
rect 780 2062 781 2063
rect 787 2063 793 2064
rect 787 2062 788 2063
rect 780 2060 788 2062
rect 780 2059 781 2060
rect 775 2058 781 2059
rect 787 2059 788 2060
rect 792 2059 793 2063
rect 787 2058 793 2059
rect 826 2063 832 2064
rect 826 2059 827 2063
rect 831 2062 832 2063
rect 931 2063 937 2064
rect 931 2062 932 2063
rect 831 2060 932 2062
rect 831 2059 832 2060
rect 826 2058 832 2059
rect 931 2059 932 2060
rect 936 2059 937 2063
rect 931 2058 937 2059
rect 1083 2063 1089 2064
rect 1083 2059 1084 2063
rect 1088 2062 1089 2063
rect 1130 2063 1136 2064
rect 1130 2062 1131 2063
rect 1088 2060 1131 2062
rect 1088 2059 1089 2060
rect 1083 2058 1089 2059
rect 1130 2059 1131 2060
rect 1135 2059 1136 2063
rect 1130 2058 1136 2059
rect 1226 2063 1232 2064
rect 1226 2059 1227 2063
rect 1231 2062 1232 2063
rect 1251 2063 1257 2064
rect 1251 2062 1252 2063
rect 1231 2060 1252 2062
rect 1231 2059 1232 2060
rect 1226 2058 1232 2059
rect 1251 2059 1252 2060
rect 1256 2059 1257 2063
rect 1251 2058 1257 2059
rect 1435 2063 1441 2064
rect 1435 2059 1436 2063
rect 1440 2062 1441 2063
rect 1482 2063 1488 2064
rect 1482 2062 1483 2063
rect 1440 2060 1483 2062
rect 1440 2059 1441 2060
rect 1435 2058 1441 2059
rect 1482 2059 1483 2060
rect 1487 2059 1488 2063
rect 1482 2058 1488 2059
rect 1619 2063 1628 2064
rect 1619 2059 1620 2063
rect 1627 2059 1628 2063
rect 1619 2058 1628 2059
rect 1811 2063 1820 2064
rect 1811 2059 1812 2063
rect 1819 2059 1820 2063
rect 3204 2062 3206 2064
rect 3618 2063 3619 2064
rect 3623 2063 3624 2067
rect 3618 2062 3624 2063
rect 3203 2061 3209 2062
rect 1811 2058 1820 2059
rect 2539 2059 2545 2060
rect 2539 2055 2540 2059
rect 2544 2058 2545 2059
rect 2562 2059 2568 2060
rect 2562 2058 2563 2059
rect 2544 2056 2563 2058
rect 2544 2055 2545 2056
rect 2539 2054 2545 2055
rect 2562 2055 2563 2056
rect 2567 2055 2568 2059
rect 2562 2054 2568 2055
rect 2623 2059 2629 2060
rect 2623 2055 2624 2059
rect 2628 2058 2629 2059
rect 2707 2059 2713 2060
rect 2707 2058 2708 2059
rect 2628 2056 2708 2058
rect 2628 2055 2629 2056
rect 2623 2054 2629 2055
rect 2707 2055 2708 2056
rect 2712 2055 2713 2059
rect 2707 2054 2713 2055
rect 2746 2059 2752 2060
rect 2746 2055 2747 2059
rect 2751 2058 2752 2059
rect 2875 2059 2881 2060
rect 2875 2058 2876 2059
rect 2751 2056 2876 2058
rect 2751 2055 2752 2056
rect 2746 2054 2752 2055
rect 2875 2055 2876 2056
rect 2880 2055 2881 2059
rect 2875 2054 2881 2055
rect 2914 2059 2920 2060
rect 2914 2055 2915 2059
rect 2919 2058 2920 2059
rect 3043 2059 3049 2060
rect 3043 2058 3044 2059
rect 2919 2056 3044 2058
rect 2919 2055 2920 2056
rect 2914 2054 2920 2055
rect 3043 2055 3044 2056
rect 3048 2055 3049 2059
rect 3203 2057 3204 2061
rect 3208 2057 3209 2061
rect 3203 2056 3209 2057
rect 3242 2059 3248 2060
rect 3043 2054 3049 2055
rect 3242 2055 3243 2059
rect 3247 2058 3248 2059
rect 3347 2059 3353 2060
rect 3347 2058 3348 2059
rect 3247 2056 3348 2058
rect 3247 2055 3248 2056
rect 3242 2054 3248 2055
rect 3347 2055 3348 2056
rect 3352 2055 3353 2059
rect 3347 2054 3353 2055
rect 3386 2059 3392 2060
rect 3386 2055 3387 2059
rect 3391 2058 3392 2059
rect 3491 2059 3497 2060
rect 3491 2058 3492 2059
rect 3391 2056 3492 2058
rect 3391 2055 3392 2056
rect 3386 2054 3392 2055
rect 3491 2055 3492 2056
rect 3496 2055 3497 2059
rect 3491 2054 3497 2055
rect 3559 2059 3565 2060
rect 3559 2055 3560 2059
rect 3564 2058 3565 2059
rect 3627 2059 3633 2060
rect 3627 2058 3628 2059
rect 3564 2056 3628 2058
rect 3564 2055 3565 2056
rect 3559 2054 3565 2055
rect 3627 2055 3628 2056
rect 3632 2055 3633 2059
rect 3627 2054 3633 2055
rect 3666 2059 3672 2060
rect 3666 2055 3667 2059
rect 3671 2058 3672 2059
rect 3763 2059 3769 2060
rect 3763 2058 3764 2059
rect 3671 2056 3764 2058
rect 3671 2055 3672 2056
rect 3666 2054 3672 2055
rect 3763 2055 3764 2056
rect 3768 2055 3769 2059
rect 3763 2054 3769 2055
rect 3875 2059 3881 2060
rect 3875 2055 3876 2059
rect 3880 2058 3881 2059
rect 3906 2059 3912 2060
rect 3906 2058 3907 2059
rect 3880 2056 3907 2058
rect 3880 2055 3881 2056
rect 3875 2054 3881 2055
rect 3906 2055 3907 2056
rect 3911 2055 3912 2059
rect 3906 2054 3912 2055
rect 110 2044 116 2045
rect 2006 2044 2012 2045
rect 110 2040 111 2044
rect 115 2040 116 2044
rect 110 2039 116 2040
rect 374 2043 380 2044
rect 374 2039 375 2043
rect 379 2039 380 2043
rect 374 2038 380 2039
rect 494 2043 500 2044
rect 494 2039 495 2043
rect 499 2039 500 2043
rect 494 2038 500 2039
rect 614 2043 620 2044
rect 614 2039 615 2043
rect 619 2039 620 2043
rect 614 2038 620 2039
rect 750 2043 756 2044
rect 750 2039 751 2043
rect 755 2039 756 2043
rect 750 2038 756 2039
rect 894 2043 900 2044
rect 894 2039 895 2043
rect 899 2039 900 2043
rect 894 2038 900 2039
rect 1046 2043 1052 2044
rect 1046 2039 1047 2043
rect 1051 2039 1052 2043
rect 1046 2038 1052 2039
rect 1214 2043 1220 2044
rect 1214 2039 1215 2043
rect 1219 2039 1220 2043
rect 1214 2038 1220 2039
rect 1398 2043 1404 2044
rect 1398 2039 1399 2043
rect 1403 2039 1404 2043
rect 1398 2038 1404 2039
rect 1582 2043 1588 2044
rect 1582 2039 1583 2043
rect 1587 2039 1588 2043
rect 1582 2038 1588 2039
rect 1774 2043 1780 2044
rect 1774 2039 1775 2043
rect 1779 2039 1780 2043
rect 2006 2040 2007 2044
rect 2011 2040 2012 2044
rect 2006 2039 2012 2040
rect 2046 2040 2052 2041
rect 3942 2040 3948 2041
rect 1774 2038 1780 2039
rect 2046 2036 2047 2040
rect 2051 2036 2052 2040
rect 450 2035 456 2036
rect 450 2031 451 2035
rect 455 2031 456 2035
rect 450 2030 456 2031
rect 570 2035 576 2036
rect 570 2031 571 2035
rect 575 2031 576 2035
rect 570 2030 576 2031
rect 690 2035 696 2036
rect 690 2031 691 2035
rect 695 2031 696 2035
rect 690 2030 696 2031
rect 826 2035 832 2036
rect 826 2031 827 2035
rect 831 2031 832 2035
rect 826 2030 832 2031
rect 886 2035 892 2036
rect 886 2031 887 2035
rect 891 2034 892 2035
rect 1002 2035 1008 2036
rect 891 2032 937 2034
rect 891 2031 892 2032
rect 886 2030 892 2031
rect 1002 2031 1003 2035
rect 1007 2034 1008 2035
rect 1130 2035 1136 2036
rect 1007 2032 1089 2034
rect 1007 2031 1008 2032
rect 1002 2030 1008 2031
rect 1130 2031 1131 2035
rect 1135 2034 1136 2035
rect 1482 2035 1488 2036
rect 1135 2032 1257 2034
rect 1135 2031 1136 2032
rect 1130 2030 1136 2031
rect 1474 2031 1480 2032
rect 110 2027 116 2028
rect 110 2023 111 2027
rect 115 2023 116 2027
rect 1474 2027 1475 2031
rect 1479 2027 1480 2031
rect 1482 2031 1483 2035
rect 1487 2034 1488 2035
rect 1754 2035 1760 2036
rect 2046 2035 2052 2036
rect 2502 2039 2508 2040
rect 2502 2035 2503 2039
rect 2507 2035 2508 2039
rect 1487 2032 1625 2034
rect 1487 2031 1488 2032
rect 1482 2030 1488 2031
rect 1754 2031 1755 2035
rect 1759 2034 1760 2035
rect 2502 2034 2508 2035
rect 2670 2039 2676 2040
rect 2670 2035 2671 2039
rect 2675 2035 2676 2039
rect 2670 2034 2676 2035
rect 2838 2039 2844 2040
rect 2838 2035 2839 2039
rect 2843 2035 2844 2039
rect 2838 2034 2844 2035
rect 3006 2039 3012 2040
rect 3006 2035 3007 2039
rect 3011 2035 3012 2039
rect 3006 2034 3012 2035
rect 3166 2039 3172 2040
rect 3166 2035 3167 2039
rect 3171 2035 3172 2039
rect 3166 2034 3172 2035
rect 3310 2039 3316 2040
rect 3310 2035 3311 2039
rect 3315 2035 3316 2039
rect 3310 2034 3316 2035
rect 3454 2039 3460 2040
rect 3454 2035 3455 2039
rect 3459 2035 3460 2039
rect 3454 2034 3460 2035
rect 3590 2039 3596 2040
rect 3590 2035 3591 2039
rect 3595 2035 3596 2039
rect 3590 2034 3596 2035
rect 3726 2039 3732 2040
rect 3726 2035 3727 2039
rect 3731 2035 3732 2039
rect 3726 2034 3732 2035
rect 3838 2039 3844 2040
rect 3838 2035 3839 2039
rect 3843 2035 3844 2039
rect 3942 2036 3943 2040
rect 3947 2036 3948 2040
rect 3942 2035 3948 2036
rect 3838 2034 3844 2035
rect 1759 2032 1817 2034
rect 1759 2031 1760 2032
rect 1754 2030 1760 2031
rect 2623 2031 2629 2032
rect 2623 2030 2624 2031
rect 2581 2028 2624 2030
rect 1474 2026 1480 2027
rect 2006 2027 2012 2028
rect 110 2022 116 2023
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 494 2024 500 2025
rect 494 2020 495 2024
rect 499 2020 500 2024
rect 494 2019 500 2020
rect 614 2024 620 2025
rect 614 2020 615 2024
rect 619 2020 620 2024
rect 614 2019 620 2020
rect 750 2024 756 2025
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 894 2024 900 2025
rect 894 2020 895 2024
rect 899 2020 900 2024
rect 894 2019 900 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1214 2024 1220 2025
rect 1214 2020 1215 2024
rect 1219 2020 1220 2024
rect 1214 2019 1220 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1582 2024 1588 2025
rect 1582 2020 1583 2024
rect 1587 2020 1588 2024
rect 1582 2019 1588 2020
rect 1774 2024 1780 2025
rect 1774 2020 1775 2024
rect 1779 2020 1780 2024
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2623 2027 2624 2028
rect 2628 2027 2629 2031
rect 2623 2026 2629 2027
rect 2746 2031 2752 2032
rect 2746 2027 2747 2031
rect 2751 2027 2752 2031
rect 2746 2026 2752 2027
rect 2914 2031 2920 2032
rect 2914 2027 2915 2031
rect 2919 2027 2920 2031
rect 2914 2026 2920 2027
rect 2926 2031 2932 2032
rect 2926 2027 2927 2031
rect 2931 2030 2932 2031
rect 3242 2031 3248 2032
rect 2931 2028 3049 2030
rect 2931 2027 2932 2028
rect 2926 2026 2932 2027
rect 3242 2027 3243 2031
rect 3247 2027 3248 2031
rect 3242 2026 3248 2027
rect 3386 2031 3392 2032
rect 3386 2027 3387 2031
rect 3391 2027 3392 2031
rect 3559 2031 3565 2032
rect 3559 2030 3560 2031
rect 3533 2028 3560 2030
rect 3386 2026 3392 2027
rect 3559 2027 3560 2028
rect 3564 2027 3565 2031
rect 3559 2026 3565 2027
rect 3666 2031 3672 2032
rect 3666 2027 3667 2031
rect 3671 2027 3672 2031
rect 3666 2026 3672 2027
rect 3710 2031 3716 2032
rect 3710 2027 3711 2031
rect 3715 2030 3716 2031
rect 3715 2028 3769 2030
rect 3715 2027 3716 2028
rect 3710 2026 3716 2027
rect 3914 2027 3920 2028
rect 2006 2022 2012 2023
rect 2046 2023 2052 2024
rect 1774 2019 1780 2020
rect 2046 2019 2047 2023
rect 2051 2019 2052 2023
rect 3914 2023 3915 2027
rect 3919 2023 3920 2027
rect 3914 2022 3920 2023
rect 3942 2023 3948 2024
rect 2046 2018 2052 2019
rect 2502 2020 2508 2021
rect 2502 2016 2503 2020
rect 2507 2016 2508 2020
rect 2502 2015 2508 2016
rect 2670 2020 2676 2021
rect 2670 2016 2671 2020
rect 2675 2016 2676 2020
rect 2670 2015 2676 2016
rect 2838 2020 2844 2021
rect 2838 2016 2839 2020
rect 2843 2016 2844 2020
rect 2838 2015 2844 2016
rect 3006 2020 3012 2021
rect 3006 2016 3007 2020
rect 3011 2016 3012 2020
rect 3006 2015 3012 2016
rect 3166 2020 3172 2021
rect 3166 2016 3167 2020
rect 3171 2016 3172 2020
rect 3166 2015 3172 2016
rect 3310 2020 3316 2021
rect 3310 2016 3311 2020
rect 3315 2016 3316 2020
rect 3310 2015 3316 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3590 2020 3596 2021
rect 3590 2016 3591 2020
rect 3595 2016 3596 2020
rect 3590 2015 3596 2016
rect 3726 2020 3732 2021
rect 3726 2016 3727 2020
rect 3731 2016 3732 2020
rect 3726 2015 3732 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3942 2019 3943 2023
rect 3947 2019 3948 2023
rect 3942 2018 3948 2019
rect 3838 2015 3844 2016
rect 510 1956 516 1957
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 510 1952 511 1956
rect 515 1952 516 1956
rect 510 1951 516 1952
rect 622 1956 628 1957
rect 622 1952 623 1956
rect 627 1952 628 1956
rect 622 1951 628 1952
rect 742 1956 748 1957
rect 742 1952 743 1956
rect 747 1952 748 1956
rect 742 1951 748 1952
rect 870 1956 876 1957
rect 870 1952 871 1956
rect 875 1952 876 1956
rect 870 1951 876 1952
rect 1006 1956 1012 1957
rect 1006 1952 1007 1956
rect 1011 1952 1012 1956
rect 1006 1951 1012 1952
rect 1142 1956 1148 1957
rect 1142 1952 1143 1956
rect 1147 1952 1148 1956
rect 1142 1951 1148 1952
rect 1278 1956 1284 1957
rect 1278 1952 1279 1956
rect 1283 1952 1284 1956
rect 1278 1951 1284 1952
rect 1414 1956 1420 1957
rect 1414 1952 1415 1956
rect 1419 1952 1420 1956
rect 1414 1951 1420 1952
rect 1558 1956 1564 1957
rect 1558 1952 1559 1956
rect 1563 1952 1564 1956
rect 1558 1951 1564 1952
rect 1702 1956 1708 1957
rect 1702 1952 1703 1956
rect 1707 1952 1708 1956
rect 2494 1956 2500 1957
rect 1702 1951 1708 1952
rect 2006 1953 2012 1954
rect 110 1948 116 1949
rect 2006 1949 2007 1953
rect 2011 1949 2012 1953
rect 2006 1948 2012 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2494 1952 2495 1956
rect 2499 1952 2500 1956
rect 2494 1951 2500 1952
rect 2590 1956 2596 1957
rect 2590 1952 2591 1956
rect 2595 1952 2596 1956
rect 2590 1951 2596 1952
rect 2694 1956 2700 1957
rect 2694 1952 2695 1956
rect 2699 1952 2700 1956
rect 2694 1951 2700 1952
rect 2806 1956 2812 1957
rect 2806 1952 2807 1956
rect 2811 1952 2812 1956
rect 2806 1951 2812 1952
rect 2926 1956 2932 1957
rect 2926 1952 2927 1956
rect 2931 1952 2932 1956
rect 2926 1951 2932 1952
rect 3046 1956 3052 1957
rect 3046 1952 3047 1956
rect 3051 1952 3052 1956
rect 3046 1951 3052 1952
rect 3174 1956 3180 1957
rect 3174 1952 3175 1956
rect 3179 1952 3180 1956
rect 3174 1951 3180 1952
rect 3294 1956 3300 1957
rect 3294 1952 3295 1956
rect 3299 1952 3300 1956
rect 3294 1951 3300 1952
rect 3414 1956 3420 1957
rect 3414 1952 3415 1956
rect 3419 1952 3420 1956
rect 3414 1951 3420 1952
rect 3542 1956 3548 1957
rect 3542 1952 3543 1956
rect 3547 1952 3548 1956
rect 3542 1951 3548 1952
rect 3670 1956 3676 1957
rect 3670 1952 3671 1956
rect 3675 1952 3676 1956
rect 3670 1951 3676 1952
rect 3798 1956 3804 1957
rect 3798 1952 3799 1956
rect 3803 1952 3804 1956
rect 3798 1951 3804 1952
rect 3942 1953 3948 1954
rect 2046 1948 2052 1949
rect 3942 1949 3943 1953
rect 3947 1949 3948 1953
rect 3942 1948 3948 1949
rect 414 1947 420 1948
rect 414 1943 415 1947
rect 419 1946 420 1947
rect 594 1947 600 1948
rect 419 1944 553 1946
rect 419 1943 420 1944
rect 414 1942 420 1943
rect 594 1943 595 1947
rect 599 1946 600 1947
rect 718 1947 724 1948
rect 599 1944 665 1946
rect 599 1943 600 1944
rect 594 1942 600 1943
rect 718 1943 719 1947
rect 723 1946 724 1947
rect 946 1947 952 1948
rect 723 1944 785 1946
rect 723 1943 724 1944
rect 718 1942 724 1943
rect 946 1943 947 1947
rect 951 1943 952 1947
rect 946 1942 952 1943
rect 1082 1947 1088 1948
rect 1082 1943 1083 1947
rect 1087 1943 1088 1947
rect 1226 1947 1232 1948
rect 1226 1946 1227 1947
rect 1221 1944 1227 1946
rect 1082 1942 1088 1943
rect 1226 1943 1227 1944
rect 1231 1943 1232 1947
rect 1226 1942 1232 1943
rect 1346 1947 1352 1948
rect 1346 1943 1347 1947
rect 1351 1943 1352 1947
rect 1346 1942 1352 1943
rect 1490 1947 1496 1948
rect 1490 1943 1491 1947
rect 1495 1943 1496 1947
rect 1490 1942 1496 1943
rect 1518 1947 1524 1948
rect 1518 1943 1519 1947
rect 1523 1946 1524 1947
rect 1770 1947 1776 1948
rect 1523 1944 1601 1946
rect 1523 1943 1524 1944
rect 1518 1942 1524 1943
rect 1770 1943 1771 1947
rect 1775 1943 1776 1947
rect 1770 1942 1776 1943
rect 2562 1947 2568 1948
rect 2562 1943 2563 1947
rect 2567 1943 2568 1947
rect 2562 1942 2568 1943
rect 2578 1947 2584 1948
rect 2578 1943 2579 1947
rect 2583 1946 2584 1947
rect 2682 1947 2688 1948
rect 2583 1944 2633 1946
rect 2583 1943 2584 1944
rect 2578 1942 2584 1943
rect 2682 1943 2683 1947
rect 2687 1946 2688 1947
rect 2778 1947 2784 1948
rect 2687 1944 2737 1946
rect 2687 1943 2688 1944
rect 2682 1942 2688 1943
rect 2778 1943 2779 1947
rect 2783 1946 2784 1947
rect 3002 1947 3008 1948
rect 2783 1944 2849 1946
rect 2783 1943 2784 1944
rect 2778 1942 2784 1943
rect 3002 1943 3003 1947
rect 3007 1943 3008 1947
rect 3002 1942 3008 1943
rect 3122 1947 3128 1948
rect 3122 1943 3123 1947
rect 3127 1943 3128 1947
rect 3122 1942 3128 1943
rect 3130 1947 3136 1948
rect 3130 1943 3131 1947
rect 3135 1946 3136 1947
rect 3258 1947 3264 1948
rect 3135 1944 3217 1946
rect 3135 1943 3136 1944
rect 3130 1942 3136 1943
rect 3258 1943 3259 1947
rect 3263 1946 3264 1947
rect 3386 1947 3392 1948
rect 3263 1944 3337 1946
rect 3263 1943 3264 1944
rect 3258 1942 3264 1943
rect 3386 1943 3387 1947
rect 3391 1946 3392 1947
rect 3511 1947 3517 1948
rect 3391 1944 3457 1946
rect 3391 1943 3392 1944
rect 3386 1942 3392 1943
rect 3511 1943 3512 1947
rect 3516 1946 3517 1947
rect 3630 1947 3636 1948
rect 3516 1944 3585 1946
rect 3516 1943 3517 1944
rect 3511 1942 3517 1943
rect 3630 1943 3631 1947
rect 3635 1946 3636 1947
rect 3866 1947 3872 1948
rect 3635 1944 3713 1946
rect 3635 1943 3636 1944
rect 3630 1942 3636 1943
rect 3866 1943 3867 1947
rect 3871 1943 3872 1947
rect 3866 1942 3872 1943
rect 510 1937 516 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 510 1933 511 1937
rect 515 1933 516 1937
rect 510 1932 516 1933
rect 622 1937 628 1938
rect 622 1933 623 1937
rect 627 1933 628 1937
rect 622 1932 628 1933
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 870 1937 876 1938
rect 870 1933 871 1937
rect 875 1933 876 1937
rect 870 1932 876 1933
rect 1006 1937 1012 1938
rect 1006 1933 1007 1937
rect 1011 1933 1012 1937
rect 1006 1932 1012 1933
rect 1142 1937 1148 1938
rect 1142 1933 1143 1937
rect 1147 1933 1148 1937
rect 1142 1932 1148 1933
rect 1278 1937 1284 1938
rect 1278 1933 1279 1937
rect 1283 1933 1284 1937
rect 1278 1932 1284 1933
rect 1414 1937 1420 1938
rect 1414 1933 1415 1937
rect 1419 1933 1420 1937
rect 1414 1932 1420 1933
rect 1558 1937 1564 1938
rect 1558 1933 1559 1937
rect 1563 1933 1564 1937
rect 1558 1932 1564 1933
rect 1702 1937 1708 1938
rect 2494 1937 2500 1938
rect 1702 1933 1703 1937
rect 1707 1933 1708 1937
rect 1702 1932 1708 1933
rect 2006 1936 2012 1937
rect 2006 1932 2007 1936
rect 2011 1932 2012 1936
rect 110 1931 116 1932
rect 2006 1931 2012 1932
rect 2046 1936 2052 1937
rect 2046 1932 2047 1936
rect 2051 1932 2052 1936
rect 2494 1933 2495 1937
rect 2499 1933 2500 1937
rect 2494 1932 2500 1933
rect 2590 1937 2596 1938
rect 2590 1933 2591 1937
rect 2595 1933 2596 1937
rect 2590 1932 2596 1933
rect 2694 1937 2700 1938
rect 2694 1933 2695 1937
rect 2699 1933 2700 1937
rect 2694 1932 2700 1933
rect 2806 1937 2812 1938
rect 2806 1933 2807 1937
rect 2811 1933 2812 1937
rect 2806 1932 2812 1933
rect 2926 1937 2932 1938
rect 2926 1933 2927 1937
rect 2931 1933 2932 1937
rect 2926 1932 2932 1933
rect 3046 1937 3052 1938
rect 3046 1933 3047 1937
rect 3051 1933 3052 1937
rect 3046 1932 3052 1933
rect 3174 1937 3180 1938
rect 3174 1933 3175 1937
rect 3179 1933 3180 1937
rect 3174 1932 3180 1933
rect 3294 1937 3300 1938
rect 3294 1933 3295 1937
rect 3299 1933 3300 1937
rect 3294 1932 3300 1933
rect 3414 1937 3420 1938
rect 3414 1933 3415 1937
rect 3419 1933 3420 1937
rect 3414 1932 3420 1933
rect 3542 1937 3548 1938
rect 3542 1933 3543 1937
rect 3547 1933 3548 1937
rect 3542 1932 3548 1933
rect 3670 1937 3676 1938
rect 3670 1933 3671 1937
rect 3675 1933 3676 1937
rect 3670 1932 3676 1933
rect 3798 1937 3804 1938
rect 3798 1933 3799 1937
rect 3803 1933 3804 1937
rect 3798 1932 3804 1933
rect 3942 1936 3948 1937
rect 3942 1932 3943 1936
rect 3947 1932 3948 1936
rect 2046 1931 2052 1932
rect 3942 1931 3948 1932
rect 1518 1927 1524 1928
rect 1518 1926 1519 1927
rect 1444 1924 1519 1926
rect 547 1919 553 1920
rect 547 1915 548 1919
rect 552 1918 553 1919
rect 594 1919 600 1920
rect 594 1918 595 1919
rect 552 1916 595 1918
rect 552 1915 553 1916
rect 547 1914 553 1915
rect 594 1915 595 1916
rect 599 1915 600 1919
rect 594 1914 600 1915
rect 659 1919 665 1920
rect 659 1915 660 1919
rect 664 1918 665 1919
rect 718 1919 724 1920
rect 718 1918 719 1919
rect 664 1916 719 1918
rect 664 1915 665 1916
rect 659 1914 665 1915
rect 718 1915 719 1916
rect 723 1915 724 1919
rect 886 1919 892 1920
rect 718 1914 724 1915
rect 779 1915 785 1916
rect 779 1911 780 1915
rect 784 1914 785 1915
rect 871 1915 877 1916
rect 871 1914 872 1915
rect 784 1912 872 1914
rect 784 1911 785 1912
rect 779 1910 785 1911
rect 871 1911 872 1912
rect 876 1911 877 1915
rect 886 1915 887 1919
rect 891 1918 892 1919
rect 907 1919 913 1920
rect 907 1918 908 1919
rect 891 1916 908 1918
rect 891 1915 892 1916
rect 886 1914 892 1915
rect 907 1915 908 1916
rect 912 1915 913 1919
rect 907 1914 913 1915
rect 946 1919 952 1920
rect 946 1915 947 1919
rect 951 1918 952 1919
rect 1043 1919 1049 1920
rect 1043 1918 1044 1919
rect 951 1916 1044 1918
rect 951 1915 952 1916
rect 946 1914 952 1915
rect 1043 1915 1044 1916
rect 1048 1915 1049 1919
rect 1315 1919 1321 1920
rect 1043 1914 1049 1915
rect 1167 1915 1173 1916
rect 871 1910 877 1911
rect 1167 1911 1168 1915
rect 1172 1914 1173 1915
rect 1179 1915 1185 1916
rect 1179 1914 1180 1915
rect 1172 1912 1180 1914
rect 1172 1911 1173 1912
rect 1167 1910 1173 1911
rect 1179 1911 1180 1912
rect 1184 1911 1185 1915
rect 1315 1915 1316 1919
rect 1320 1918 1321 1919
rect 1444 1918 1446 1924
rect 1518 1923 1519 1924
rect 1523 1923 1524 1927
rect 3130 1927 3136 1928
rect 3130 1926 3131 1927
rect 1518 1922 1524 1923
rect 2860 1924 3131 1926
rect 1320 1916 1446 1918
rect 1451 1919 1457 1920
rect 1320 1915 1321 1916
rect 1315 1914 1321 1915
rect 1451 1915 1452 1919
rect 1456 1918 1457 1919
rect 1474 1919 1480 1920
rect 1474 1918 1475 1919
rect 1456 1916 1475 1918
rect 1456 1915 1457 1916
rect 1451 1914 1457 1915
rect 1474 1915 1475 1916
rect 1479 1915 1480 1919
rect 1474 1914 1480 1915
rect 1490 1919 1496 1920
rect 1490 1915 1491 1919
rect 1495 1918 1496 1919
rect 1595 1919 1601 1920
rect 1595 1918 1596 1919
rect 1495 1916 1596 1918
rect 1495 1915 1496 1916
rect 1490 1914 1496 1915
rect 1595 1915 1596 1916
rect 1600 1915 1601 1919
rect 1595 1914 1601 1915
rect 1739 1919 1745 1920
rect 1739 1915 1740 1919
rect 1744 1918 1745 1919
rect 1754 1919 1760 1920
rect 1754 1918 1755 1919
rect 1744 1916 1755 1918
rect 1744 1915 1745 1916
rect 1739 1914 1745 1915
rect 1754 1915 1755 1916
rect 1759 1915 1760 1919
rect 1754 1914 1760 1915
rect 2531 1919 2537 1920
rect 2531 1915 2532 1919
rect 2536 1918 2537 1919
rect 2578 1919 2584 1920
rect 2578 1918 2579 1919
rect 2536 1916 2579 1918
rect 2536 1915 2537 1916
rect 2531 1914 2537 1915
rect 2578 1915 2579 1916
rect 2583 1915 2584 1919
rect 2578 1914 2584 1915
rect 2627 1919 2633 1920
rect 2627 1915 2628 1919
rect 2632 1918 2633 1919
rect 2682 1919 2688 1920
rect 2682 1918 2683 1919
rect 2632 1916 2683 1918
rect 2632 1915 2633 1916
rect 2627 1914 2633 1915
rect 2682 1915 2683 1916
rect 2687 1915 2688 1919
rect 2682 1914 2688 1915
rect 2731 1919 2737 1920
rect 2731 1915 2732 1919
rect 2736 1918 2737 1919
rect 2778 1919 2784 1920
rect 2778 1918 2779 1919
rect 2736 1916 2779 1918
rect 2736 1915 2737 1916
rect 2731 1914 2737 1915
rect 2778 1915 2779 1916
rect 2783 1915 2784 1919
rect 2778 1914 2784 1915
rect 2843 1919 2849 1920
rect 2843 1915 2844 1919
rect 2848 1918 2849 1919
rect 2860 1918 2862 1924
rect 3130 1923 3131 1924
rect 3135 1923 3136 1927
rect 3130 1922 3136 1923
rect 2848 1916 2862 1918
rect 3002 1919 3008 1920
rect 2848 1915 2849 1916
rect 2843 1914 2849 1915
rect 2866 1915 2872 1916
rect 1179 1910 1185 1911
rect 2866 1911 2867 1915
rect 2871 1914 2872 1915
rect 2963 1915 2969 1916
rect 2963 1914 2964 1915
rect 2871 1912 2964 1914
rect 2871 1911 2872 1912
rect 2866 1910 2872 1911
rect 2963 1911 2964 1912
rect 2968 1911 2969 1915
rect 3002 1915 3003 1919
rect 3007 1918 3008 1919
rect 3083 1919 3089 1920
rect 3083 1918 3084 1919
rect 3007 1916 3084 1918
rect 3007 1915 3008 1916
rect 3002 1914 3008 1915
rect 3083 1915 3084 1916
rect 3088 1915 3089 1919
rect 3083 1914 3089 1915
rect 3122 1919 3128 1920
rect 3122 1915 3123 1919
rect 3127 1918 3128 1919
rect 3211 1919 3217 1920
rect 3211 1918 3212 1919
rect 3127 1916 3212 1918
rect 3127 1915 3128 1916
rect 3122 1914 3128 1915
rect 3211 1915 3212 1916
rect 3216 1915 3217 1919
rect 3211 1914 3217 1915
rect 3331 1919 3337 1920
rect 3331 1915 3332 1919
rect 3336 1918 3337 1919
rect 3386 1919 3392 1920
rect 3386 1918 3387 1919
rect 3336 1916 3387 1918
rect 3336 1915 3337 1916
rect 3331 1914 3337 1915
rect 3386 1915 3387 1916
rect 3391 1915 3392 1919
rect 3386 1914 3392 1915
rect 3451 1919 3457 1920
rect 3451 1915 3452 1919
rect 3456 1918 3457 1919
rect 3511 1919 3517 1920
rect 3511 1918 3512 1919
rect 3456 1916 3512 1918
rect 3456 1915 3457 1916
rect 3451 1914 3457 1915
rect 3511 1915 3512 1916
rect 3516 1915 3517 1919
rect 3511 1914 3517 1915
rect 3579 1919 3585 1920
rect 3579 1915 3580 1919
rect 3584 1918 3585 1919
rect 3630 1919 3636 1920
rect 3630 1918 3631 1919
rect 3584 1916 3631 1918
rect 3584 1915 3585 1916
rect 3579 1914 3585 1915
rect 3630 1915 3631 1916
rect 3635 1915 3636 1919
rect 3630 1914 3636 1915
rect 3707 1919 3716 1920
rect 3707 1915 3708 1919
rect 3715 1915 3716 1919
rect 3707 1914 3716 1915
rect 3835 1915 3841 1916
rect 2963 1910 2969 1911
rect 3835 1911 3836 1915
rect 3840 1914 3841 1915
rect 3858 1915 3864 1916
rect 3858 1914 3859 1915
rect 3840 1912 3859 1914
rect 3840 1911 3841 1912
rect 3835 1910 3841 1911
rect 3858 1911 3859 1912
rect 3863 1911 3864 1915
rect 3858 1910 3864 1911
rect 3258 1907 3264 1908
rect 3258 1906 3259 1907
rect 2996 1904 3259 1906
rect 2996 1902 2998 1904
rect 3258 1903 3259 1904
rect 3263 1903 3264 1907
rect 3258 1902 3264 1903
rect 2995 1901 3001 1902
rect 1922 1899 1928 1900
rect 578 1895 584 1896
rect 578 1891 579 1895
rect 583 1894 584 1895
rect 587 1895 593 1896
rect 587 1894 588 1895
rect 583 1892 588 1894
rect 583 1891 584 1892
rect 578 1890 584 1891
rect 587 1891 588 1892
rect 592 1891 593 1895
rect 587 1890 593 1891
rect 646 1895 652 1896
rect 646 1891 647 1895
rect 651 1894 652 1895
rect 699 1895 705 1896
rect 699 1894 700 1895
rect 651 1892 700 1894
rect 651 1891 652 1892
rect 646 1890 652 1891
rect 699 1891 700 1892
rect 704 1891 705 1895
rect 699 1890 705 1891
rect 759 1895 765 1896
rect 759 1891 760 1895
rect 764 1894 765 1895
rect 819 1895 825 1896
rect 819 1894 820 1895
rect 764 1892 820 1894
rect 764 1891 765 1892
rect 759 1890 765 1891
rect 819 1891 820 1892
rect 824 1891 825 1895
rect 819 1890 825 1891
rect 858 1895 864 1896
rect 858 1891 859 1895
rect 863 1894 864 1895
rect 947 1895 953 1896
rect 947 1894 948 1895
rect 863 1892 948 1894
rect 863 1891 864 1892
rect 858 1890 864 1891
rect 947 1891 948 1892
rect 952 1891 953 1895
rect 947 1890 953 1891
rect 1082 1895 1089 1896
rect 1082 1891 1083 1895
rect 1088 1891 1089 1895
rect 1082 1890 1089 1891
rect 1211 1895 1220 1896
rect 1211 1891 1212 1895
rect 1219 1891 1220 1895
rect 1211 1890 1220 1891
rect 1346 1895 1353 1896
rect 1346 1891 1347 1895
rect 1352 1891 1353 1895
rect 1346 1890 1353 1891
rect 1386 1895 1392 1896
rect 1386 1891 1387 1895
rect 1391 1894 1392 1895
rect 1483 1895 1489 1896
rect 1483 1894 1484 1895
rect 1391 1892 1484 1894
rect 1391 1891 1392 1892
rect 1386 1890 1392 1891
rect 1483 1891 1484 1892
rect 1488 1891 1489 1895
rect 1483 1890 1489 1891
rect 1522 1895 1528 1896
rect 1522 1891 1523 1895
rect 1527 1894 1528 1895
rect 1619 1895 1625 1896
rect 1619 1894 1620 1895
rect 1527 1892 1620 1894
rect 1527 1891 1528 1892
rect 1522 1890 1528 1891
rect 1619 1891 1620 1892
rect 1624 1891 1625 1895
rect 1619 1890 1625 1891
rect 1755 1895 1761 1896
rect 1755 1891 1756 1895
rect 1760 1894 1761 1895
rect 1770 1895 1776 1896
rect 1770 1894 1771 1895
rect 1760 1892 1771 1894
rect 1760 1891 1761 1892
rect 1755 1890 1761 1891
rect 1770 1891 1771 1892
rect 1775 1891 1776 1895
rect 1922 1895 1923 1899
rect 1927 1898 1928 1899
rect 2107 1899 2113 1900
rect 2107 1898 2108 1899
rect 1927 1896 2108 1898
rect 1927 1895 1928 1896
rect 1922 1894 1928 1895
rect 2107 1895 2108 1896
rect 2112 1895 2113 1899
rect 2322 1899 2328 1900
rect 2107 1894 2113 1895
rect 2283 1897 2289 1898
rect 2283 1893 2284 1897
rect 2288 1893 2289 1897
rect 2322 1895 2323 1899
rect 2327 1898 2328 1899
rect 2475 1899 2481 1900
rect 2475 1898 2476 1899
rect 2327 1896 2476 1898
rect 2327 1895 2328 1896
rect 2322 1894 2328 1895
rect 2475 1895 2476 1896
rect 2480 1895 2481 1899
rect 2475 1894 2481 1895
rect 2514 1899 2520 1900
rect 2514 1895 2515 1899
rect 2519 1898 2520 1899
rect 2659 1899 2665 1900
rect 2659 1898 2660 1899
rect 2519 1896 2660 1898
rect 2519 1895 2520 1896
rect 2514 1894 2520 1895
rect 2659 1895 2660 1896
rect 2664 1895 2665 1899
rect 2659 1894 2665 1895
rect 2743 1899 2749 1900
rect 2743 1895 2744 1899
rect 2748 1898 2749 1899
rect 2827 1899 2833 1900
rect 2827 1898 2828 1899
rect 2748 1896 2828 1898
rect 2748 1895 2749 1896
rect 2743 1894 2749 1895
rect 2827 1895 2828 1896
rect 2832 1895 2833 1899
rect 2995 1897 2996 1901
rect 3000 1897 3001 1901
rect 2995 1896 3001 1897
rect 3034 1899 3040 1900
rect 2827 1894 2833 1895
rect 3034 1895 3035 1899
rect 3039 1898 3040 1899
rect 3163 1899 3169 1900
rect 3163 1898 3164 1899
rect 3039 1896 3164 1898
rect 3039 1895 3040 1896
rect 3034 1894 3040 1895
rect 3163 1895 3164 1896
rect 3168 1895 3169 1899
rect 3163 1894 3169 1895
rect 3202 1899 3208 1900
rect 3202 1895 3203 1899
rect 3207 1898 3208 1899
rect 3339 1899 3345 1900
rect 3339 1898 3340 1899
rect 3207 1896 3340 1898
rect 3207 1895 3208 1896
rect 3202 1894 3208 1895
rect 3339 1895 3340 1896
rect 3344 1895 3345 1899
rect 3339 1894 3345 1895
rect 3378 1899 3384 1900
rect 3378 1895 3379 1899
rect 3383 1898 3384 1899
rect 3523 1899 3529 1900
rect 3523 1898 3524 1899
rect 3383 1896 3524 1898
rect 3383 1895 3384 1896
rect 3378 1894 3384 1895
rect 3523 1895 3524 1896
rect 3528 1895 3529 1899
rect 3523 1894 3529 1895
rect 3562 1899 3568 1900
rect 3562 1895 3563 1899
rect 3567 1898 3568 1899
rect 3707 1899 3713 1900
rect 3707 1898 3708 1899
rect 3567 1896 3708 1898
rect 3567 1895 3568 1896
rect 3562 1894 3568 1895
rect 3707 1895 3708 1896
rect 3712 1895 3713 1899
rect 3707 1894 3713 1895
rect 3875 1899 3881 1900
rect 3875 1895 3876 1899
rect 3880 1898 3881 1899
rect 3914 1899 3920 1900
rect 3914 1898 3915 1899
rect 3880 1896 3915 1898
rect 3880 1895 3881 1896
rect 3875 1894 3881 1895
rect 3914 1895 3915 1896
rect 3919 1895 3920 1899
rect 3914 1894 3920 1895
rect 2283 1892 2289 1893
rect 1770 1890 1776 1891
rect 2284 1890 2286 1892
rect 2478 1891 2484 1892
rect 2478 1890 2479 1891
rect 2284 1888 2479 1890
rect 2478 1887 2479 1888
rect 2483 1887 2484 1891
rect 2478 1886 2484 1887
rect 2046 1880 2052 1881
rect 3942 1880 3948 1881
rect 110 1876 116 1877
rect 2006 1876 2012 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 550 1875 556 1876
rect 550 1871 551 1875
rect 555 1871 556 1875
rect 550 1870 556 1871
rect 662 1875 668 1876
rect 662 1871 663 1875
rect 667 1871 668 1875
rect 662 1870 668 1871
rect 782 1875 788 1876
rect 782 1871 783 1875
rect 787 1871 788 1875
rect 782 1870 788 1871
rect 910 1875 916 1876
rect 910 1871 911 1875
rect 915 1871 916 1875
rect 910 1870 916 1871
rect 1046 1875 1052 1876
rect 1046 1871 1047 1875
rect 1051 1871 1052 1875
rect 1046 1870 1052 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1174 1870 1180 1871
rect 1310 1875 1316 1876
rect 1310 1871 1311 1875
rect 1315 1871 1316 1875
rect 1310 1870 1316 1871
rect 1446 1875 1452 1876
rect 1446 1871 1447 1875
rect 1451 1871 1452 1875
rect 1446 1870 1452 1871
rect 1582 1875 1588 1876
rect 1582 1871 1583 1875
rect 1587 1871 1588 1875
rect 1582 1870 1588 1871
rect 1718 1875 1724 1876
rect 1718 1871 1719 1875
rect 1723 1871 1724 1875
rect 2006 1872 2007 1876
rect 2011 1872 2012 1876
rect 2046 1876 2047 1880
rect 2051 1876 2052 1880
rect 2046 1875 2052 1876
rect 2070 1879 2076 1880
rect 2070 1875 2071 1879
rect 2075 1875 2076 1879
rect 2070 1874 2076 1875
rect 2246 1879 2252 1880
rect 2246 1875 2247 1879
rect 2251 1875 2252 1879
rect 2246 1874 2252 1875
rect 2438 1879 2444 1880
rect 2438 1875 2439 1879
rect 2443 1875 2444 1879
rect 2438 1874 2444 1875
rect 2622 1879 2628 1880
rect 2622 1875 2623 1879
rect 2627 1875 2628 1879
rect 2622 1874 2628 1875
rect 2790 1879 2796 1880
rect 2790 1875 2791 1879
rect 2795 1875 2796 1879
rect 2790 1874 2796 1875
rect 2958 1879 2964 1880
rect 2958 1875 2959 1879
rect 2963 1875 2964 1879
rect 2958 1874 2964 1875
rect 3126 1879 3132 1880
rect 3126 1875 3127 1879
rect 3131 1875 3132 1879
rect 3126 1874 3132 1875
rect 3302 1879 3308 1880
rect 3302 1875 3303 1879
rect 3307 1875 3308 1879
rect 3302 1874 3308 1875
rect 3486 1879 3492 1880
rect 3486 1875 3487 1879
rect 3491 1875 3492 1879
rect 3486 1874 3492 1875
rect 3670 1879 3676 1880
rect 3670 1875 3671 1879
rect 3675 1875 3676 1879
rect 3670 1874 3676 1875
rect 3838 1879 3844 1880
rect 3838 1875 3839 1879
rect 3843 1875 3844 1879
rect 3942 1876 3943 1880
rect 3947 1876 3948 1880
rect 3942 1875 3948 1876
rect 3838 1874 3844 1875
rect 2006 1871 2012 1872
rect 2322 1871 2328 1872
rect 1718 1870 1724 1871
rect 646 1867 652 1868
rect 646 1866 647 1867
rect 629 1864 647 1866
rect 646 1863 647 1864
rect 651 1863 652 1867
rect 759 1867 765 1868
rect 759 1866 760 1867
rect 741 1864 760 1866
rect 646 1862 652 1863
rect 759 1863 760 1864
rect 764 1863 765 1867
rect 759 1862 765 1863
rect 858 1867 864 1868
rect 858 1863 859 1867
rect 863 1863 864 1867
rect 858 1862 864 1863
rect 871 1867 877 1868
rect 871 1863 872 1867
rect 876 1866 877 1867
rect 1038 1867 1044 1868
rect 876 1864 953 1866
rect 876 1863 877 1864
rect 871 1862 877 1863
rect 1038 1863 1039 1867
rect 1043 1866 1044 1867
rect 1167 1867 1173 1868
rect 1043 1864 1089 1866
rect 1043 1863 1044 1864
rect 1038 1862 1044 1863
rect 1167 1863 1168 1867
rect 1172 1866 1173 1867
rect 1386 1867 1392 1868
rect 1172 1864 1217 1866
rect 1172 1863 1173 1864
rect 1167 1862 1173 1863
rect 1386 1863 1387 1867
rect 1391 1863 1392 1867
rect 1386 1862 1392 1863
rect 1522 1867 1528 1868
rect 1522 1863 1523 1867
rect 1527 1863 1528 1867
rect 1522 1862 1528 1863
rect 1702 1867 1708 1868
rect 1702 1863 1703 1867
rect 1707 1866 1708 1867
rect 2146 1867 2152 1868
rect 1707 1864 1761 1866
rect 1707 1863 1708 1864
rect 1702 1862 1708 1863
rect 2046 1863 2052 1864
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 1660 1858 1662 1861
rect 1710 1859 1716 1860
rect 1710 1858 1711 1859
rect 110 1854 116 1855
rect 550 1856 556 1857
rect 550 1852 551 1856
rect 555 1852 556 1856
rect 550 1851 556 1852
rect 662 1856 668 1857
rect 662 1852 663 1856
rect 667 1852 668 1856
rect 662 1851 668 1852
rect 782 1856 788 1857
rect 782 1852 783 1856
rect 787 1852 788 1856
rect 782 1851 788 1852
rect 910 1856 916 1857
rect 910 1852 911 1856
rect 915 1852 916 1856
rect 910 1851 916 1852
rect 1046 1856 1052 1857
rect 1046 1852 1047 1856
rect 1051 1852 1052 1856
rect 1046 1851 1052 1852
rect 1174 1856 1180 1857
rect 1174 1852 1175 1856
rect 1179 1852 1180 1856
rect 1174 1851 1180 1852
rect 1310 1856 1316 1857
rect 1310 1852 1311 1856
rect 1315 1852 1316 1856
rect 1310 1851 1316 1852
rect 1446 1856 1452 1857
rect 1446 1852 1447 1856
rect 1451 1852 1452 1856
rect 1446 1851 1452 1852
rect 1582 1856 1588 1857
rect 1660 1856 1711 1858
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1710 1855 1711 1856
rect 1715 1855 1716 1859
rect 2006 1859 2012 1860
rect 1710 1854 1716 1855
rect 1718 1856 1724 1857
rect 1582 1851 1588 1852
rect 1718 1852 1719 1856
rect 1723 1852 1724 1856
rect 2006 1855 2007 1859
rect 2011 1855 2012 1859
rect 2046 1859 2047 1863
rect 2051 1859 2052 1863
rect 2146 1863 2147 1867
rect 2151 1863 2152 1867
rect 2322 1867 2323 1871
rect 2327 1867 2328 1871
rect 2322 1866 2328 1867
rect 2514 1871 2520 1872
rect 2514 1867 2515 1871
rect 2519 1867 2520 1871
rect 2743 1871 2749 1872
rect 2743 1870 2744 1871
rect 2701 1868 2744 1870
rect 2514 1866 2520 1867
rect 2743 1867 2744 1868
rect 2748 1867 2749 1871
rect 2743 1866 2749 1867
rect 2866 1871 2872 1872
rect 2866 1867 2867 1871
rect 2871 1867 2872 1871
rect 2866 1866 2872 1867
rect 3034 1871 3040 1872
rect 3034 1867 3035 1871
rect 3039 1867 3040 1871
rect 3034 1866 3040 1867
rect 3202 1871 3208 1872
rect 3202 1867 3203 1871
rect 3207 1867 3208 1871
rect 3202 1866 3208 1867
rect 3378 1871 3384 1872
rect 3378 1867 3379 1871
rect 3383 1867 3384 1871
rect 3378 1866 3384 1867
rect 3562 1871 3568 1872
rect 3562 1867 3563 1871
rect 3567 1867 3568 1871
rect 3562 1866 3568 1867
rect 3606 1871 3612 1872
rect 3606 1867 3607 1871
rect 3611 1870 3612 1871
rect 3611 1868 3713 1870
rect 3611 1867 3612 1868
rect 3606 1866 3612 1867
rect 3914 1867 3920 1868
rect 2146 1862 2152 1863
rect 3914 1863 3915 1867
rect 3919 1863 3920 1867
rect 3914 1862 3920 1863
rect 3942 1863 3948 1864
rect 2046 1858 2052 1859
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2070 1855 2076 1856
rect 2246 1860 2252 1861
rect 2246 1856 2247 1860
rect 2251 1856 2252 1860
rect 2246 1855 2252 1856
rect 2438 1860 2444 1861
rect 2438 1856 2439 1860
rect 2443 1856 2444 1860
rect 2438 1855 2444 1856
rect 2622 1860 2628 1861
rect 2622 1856 2623 1860
rect 2627 1856 2628 1860
rect 2622 1855 2628 1856
rect 2790 1860 2796 1861
rect 2790 1856 2791 1860
rect 2795 1856 2796 1860
rect 2790 1855 2796 1856
rect 2958 1860 2964 1861
rect 2958 1856 2959 1860
rect 2963 1856 2964 1860
rect 2958 1855 2964 1856
rect 3126 1860 3132 1861
rect 3126 1856 3127 1860
rect 3131 1856 3132 1860
rect 3126 1855 3132 1856
rect 3302 1860 3308 1861
rect 3302 1856 3303 1860
rect 3307 1856 3308 1860
rect 3302 1855 3308 1856
rect 3486 1860 3492 1861
rect 3486 1856 3487 1860
rect 3491 1856 3492 1860
rect 3486 1855 3492 1856
rect 3670 1860 3676 1861
rect 3670 1856 3671 1860
rect 3675 1856 3676 1860
rect 3670 1855 3676 1856
rect 3838 1860 3844 1861
rect 3838 1856 3839 1860
rect 3843 1856 3844 1860
rect 3942 1859 3943 1863
rect 3947 1859 3948 1863
rect 3942 1858 3948 1859
rect 3838 1855 3844 1856
rect 2006 1854 2012 1855
rect 1718 1851 1724 1852
rect 2094 1800 2100 1801
rect 2046 1797 2052 1798
rect 502 1796 508 1797
rect 110 1793 116 1794
rect 110 1789 111 1793
rect 115 1789 116 1793
rect 502 1792 503 1796
rect 507 1792 508 1796
rect 502 1791 508 1792
rect 614 1796 620 1797
rect 614 1792 615 1796
rect 619 1792 620 1796
rect 614 1791 620 1792
rect 734 1796 740 1797
rect 734 1792 735 1796
rect 739 1792 740 1796
rect 734 1791 740 1792
rect 862 1796 868 1797
rect 862 1792 863 1796
rect 867 1792 868 1796
rect 862 1791 868 1792
rect 998 1796 1004 1797
rect 998 1792 999 1796
rect 1003 1792 1004 1796
rect 998 1791 1004 1792
rect 1150 1796 1156 1797
rect 1150 1792 1151 1796
rect 1155 1792 1156 1796
rect 1150 1791 1156 1792
rect 1318 1796 1324 1797
rect 1318 1792 1319 1796
rect 1323 1792 1324 1796
rect 1318 1791 1324 1792
rect 1486 1796 1492 1797
rect 1486 1792 1487 1796
rect 1491 1792 1492 1796
rect 1486 1791 1492 1792
rect 1662 1796 1668 1797
rect 1662 1792 1663 1796
rect 1667 1792 1668 1796
rect 1662 1791 1668 1792
rect 1846 1796 1852 1797
rect 1846 1792 1847 1796
rect 1851 1792 1852 1796
rect 1846 1791 1852 1792
rect 2006 1793 2012 1794
rect 110 1788 116 1789
rect 2006 1789 2007 1793
rect 2011 1789 2012 1793
rect 2046 1793 2047 1797
rect 2051 1793 2052 1797
rect 2094 1796 2095 1800
rect 2099 1796 2100 1800
rect 2094 1795 2100 1796
rect 2230 1800 2236 1801
rect 2230 1796 2231 1800
rect 2235 1796 2236 1800
rect 2230 1795 2236 1796
rect 2366 1800 2372 1801
rect 2366 1796 2367 1800
rect 2371 1796 2372 1800
rect 2366 1795 2372 1796
rect 2510 1800 2516 1801
rect 2510 1796 2511 1800
rect 2515 1796 2516 1800
rect 2510 1795 2516 1796
rect 2670 1800 2676 1801
rect 2670 1796 2671 1800
rect 2675 1796 2676 1800
rect 2670 1795 2676 1796
rect 2854 1800 2860 1801
rect 2854 1796 2855 1800
rect 2859 1796 2860 1800
rect 2854 1795 2860 1796
rect 3070 1800 3076 1801
rect 3070 1796 3071 1800
rect 3075 1796 3076 1800
rect 3070 1795 3076 1796
rect 3302 1800 3308 1801
rect 3302 1796 3303 1800
rect 3307 1796 3308 1800
rect 3302 1795 3308 1796
rect 3542 1800 3548 1801
rect 3542 1796 3543 1800
rect 3547 1796 3548 1800
rect 3542 1795 3548 1796
rect 3790 1800 3796 1801
rect 3790 1796 3791 1800
rect 3795 1796 3796 1800
rect 3790 1795 3796 1796
rect 3942 1797 3948 1798
rect 2046 1792 2052 1793
rect 3942 1793 3943 1797
rect 3947 1793 3948 1797
rect 3942 1792 3948 1793
rect 2006 1788 2012 1789
rect 2170 1791 2176 1792
rect 578 1787 584 1788
rect 578 1783 579 1787
rect 583 1783 584 1787
rect 578 1782 584 1783
rect 590 1787 596 1788
rect 590 1783 591 1787
rect 595 1786 596 1787
rect 710 1787 716 1788
rect 595 1784 657 1786
rect 595 1783 596 1784
rect 590 1782 596 1783
rect 710 1783 711 1787
rect 715 1786 716 1787
rect 930 1787 936 1788
rect 715 1784 777 1786
rect 715 1783 716 1784
rect 710 1782 716 1783
rect 930 1783 931 1787
rect 935 1783 936 1787
rect 930 1782 936 1783
rect 970 1787 976 1788
rect 970 1783 971 1787
rect 975 1786 976 1787
rect 1218 1787 1224 1788
rect 975 1784 1041 1786
rect 975 1783 976 1784
rect 970 1782 976 1783
rect 1218 1783 1219 1787
rect 1223 1783 1224 1787
rect 1218 1782 1224 1783
rect 1262 1787 1268 1788
rect 1262 1783 1263 1787
rect 1267 1786 1268 1787
rect 1562 1787 1568 1788
rect 1267 1784 1361 1786
rect 1267 1783 1268 1784
rect 1262 1782 1268 1783
rect 1562 1783 1563 1787
rect 1567 1783 1568 1787
rect 1562 1782 1568 1783
rect 1615 1787 1621 1788
rect 1615 1783 1616 1787
rect 1620 1786 1621 1787
rect 1922 1787 1928 1788
rect 1620 1784 1705 1786
rect 1620 1783 1621 1784
rect 1615 1782 1621 1783
rect 1922 1783 1923 1787
rect 1927 1783 1928 1787
rect 2170 1787 2171 1791
rect 2175 1787 2176 1791
rect 2170 1786 2176 1787
rect 2306 1791 2312 1792
rect 2306 1787 2307 1791
rect 2311 1787 2312 1791
rect 2306 1786 2312 1787
rect 2434 1791 2440 1792
rect 2434 1787 2435 1791
rect 2439 1787 2440 1791
rect 2434 1786 2440 1787
rect 2478 1791 2484 1792
rect 2478 1787 2479 1791
rect 2483 1790 2484 1791
rect 2607 1791 2613 1792
rect 2483 1788 2553 1790
rect 2483 1787 2484 1788
rect 2478 1786 2484 1787
rect 2607 1787 2608 1791
rect 2612 1790 2613 1791
rect 2770 1791 2776 1792
rect 2612 1788 2713 1790
rect 2612 1787 2613 1788
rect 2607 1786 2613 1787
rect 2770 1787 2771 1791
rect 2775 1790 2776 1791
rect 2938 1791 2944 1792
rect 2775 1788 2897 1790
rect 2775 1787 2776 1788
rect 2770 1786 2776 1787
rect 2938 1787 2939 1791
rect 2943 1790 2944 1791
rect 3166 1791 3172 1792
rect 2943 1788 3113 1790
rect 2943 1787 2944 1788
rect 2938 1786 2944 1787
rect 3166 1787 3167 1791
rect 3171 1790 3172 1791
rect 3422 1791 3428 1792
rect 3171 1788 3345 1790
rect 3171 1787 3172 1788
rect 3166 1786 3172 1787
rect 3422 1787 3423 1791
rect 3427 1790 3428 1791
rect 3858 1791 3864 1792
rect 3427 1788 3585 1790
rect 3427 1787 3428 1788
rect 3422 1786 3428 1787
rect 3858 1787 3859 1791
rect 3863 1787 3864 1791
rect 3858 1786 3864 1787
rect 1922 1782 1928 1783
rect 2094 1781 2100 1782
rect 2046 1780 2052 1781
rect 502 1777 508 1778
rect 110 1776 116 1777
rect 110 1772 111 1776
rect 115 1772 116 1776
rect 502 1773 503 1777
rect 507 1773 508 1777
rect 502 1772 508 1773
rect 614 1777 620 1778
rect 614 1773 615 1777
rect 619 1773 620 1777
rect 614 1772 620 1773
rect 734 1777 740 1778
rect 734 1773 735 1777
rect 739 1773 740 1777
rect 734 1772 740 1773
rect 862 1777 868 1778
rect 862 1773 863 1777
rect 867 1773 868 1777
rect 862 1772 868 1773
rect 998 1777 1004 1778
rect 998 1773 999 1777
rect 1003 1773 1004 1777
rect 998 1772 1004 1773
rect 1150 1777 1156 1778
rect 1150 1773 1151 1777
rect 1155 1773 1156 1777
rect 1150 1772 1156 1773
rect 1318 1777 1324 1778
rect 1318 1773 1319 1777
rect 1323 1773 1324 1777
rect 1318 1772 1324 1773
rect 1486 1777 1492 1778
rect 1486 1773 1487 1777
rect 1491 1773 1492 1777
rect 1486 1772 1492 1773
rect 1662 1777 1668 1778
rect 1662 1773 1663 1777
rect 1667 1773 1668 1777
rect 1662 1772 1668 1773
rect 1846 1777 1852 1778
rect 1846 1773 1847 1777
rect 1851 1773 1852 1777
rect 1846 1772 1852 1773
rect 2006 1776 2012 1777
rect 2006 1772 2007 1776
rect 2011 1772 2012 1776
rect 2046 1776 2047 1780
rect 2051 1776 2052 1780
rect 2094 1777 2095 1781
rect 2099 1777 2100 1781
rect 2094 1776 2100 1777
rect 2230 1781 2236 1782
rect 2230 1777 2231 1781
rect 2235 1777 2236 1781
rect 2230 1776 2236 1777
rect 2366 1781 2372 1782
rect 2366 1777 2367 1781
rect 2371 1777 2372 1781
rect 2366 1776 2372 1777
rect 2510 1781 2516 1782
rect 2510 1777 2511 1781
rect 2515 1777 2516 1781
rect 2510 1776 2516 1777
rect 2670 1781 2676 1782
rect 2670 1777 2671 1781
rect 2675 1777 2676 1781
rect 2670 1776 2676 1777
rect 2854 1781 2860 1782
rect 2854 1777 2855 1781
rect 2859 1777 2860 1781
rect 2854 1776 2860 1777
rect 3070 1781 3076 1782
rect 3070 1777 3071 1781
rect 3075 1777 3076 1781
rect 3070 1776 3076 1777
rect 3302 1781 3308 1782
rect 3302 1777 3303 1781
rect 3307 1777 3308 1781
rect 3302 1776 3308 1777
rect 3542 1781 3548 1782
rect 3542 1777 3543 1781
rect 3547 1777 3548 1781
rect 3542 1776 3548 1777
rect 3790 1781 3796 1782
rect 3790 1777 3791 1781
rect 3795 1777 3796 1781
rect 3790 1776 3796 1777
rect 3942 1780 3948 1781
rect 3942 1776 3943 1780
rect 3947 1776 3948 1780
rect 2046 1775 2052 1776
rect 3942 1775 3948 1776
rect 110 1771 116 1772
rect 2006 1771 2012 1772
rect 2131 1763 2137 1764
rect 539 1759 545 1760
rect 539 1755 540 1759
rect 544 1758 545 1759
rect 590 1759 596 1760
rect 590 1758 591 1759
rect 544 1756 591 1758
rect 544 1755 545 1756
rect 539 1754 545 1755
rect 590 1755 591 1756
rect 595 1755 596 1759
rect 590 1754 596 1755
rect 651 1759 657 1760
rect 651 1755 652 1759
rect 656 1758 657 1759
rect 710 1759 716 1760
rect 710 1758 711 1759
rect 656 1756 711 1758
rect 656 1755 657 1756
rect 651 1754 657 1755
rect 710 1755 711 1756
rect 715 1755 716 1759
rect 899 1759 905 1760
rect 710 1754 716 1755
rect 771 1755 777 1756
rect 771 1751 772 1755
rect 776 1754 777 1755
rect 794 1755 800 1756
rect 794 1754 795 1755
rect 776 1752 795 1754
rect 776 1751 777 1752
rect 771 1750 777 1751
rect 794 1751 795 1752
rect 799 1751 800 1755
rect 899 1755 900 1759
rect 904 1758 905 1759
rect 970 1759 976 1760
rect 970 1758 971 1759
rect 904 1756 971 1758
rect 904 1755 905 1756
rect 899 1754 905 1755
rect 970 1755 971 1756
rect 975 1755 976 1759
rect 970 1754 976 1755
rect 1035 1759 1044 1760
rect 1035 1755 1036 1759
rect 1043 1755 1044 1759
rect 1035 1754 1044 1755
rect 1187 1759 1193 1760
rect 1187 1755 1188 1759
rect 1192 1758 1193 1759
rect 1262 1759 1268 1760
rect 1262 1758 1263 1759
rect 1192 1756 1263 1758
rect 1192 1755 1193 1756
rect 1187 1754 1193 1755
rect 1262 1755 1263 1756
rect 1267 1755 1268 1759
rect 1523 1759 1529 1760
rect 1262 1754 1268 1755
rect 1355 1755 1364 1756
rect 794 1750 800 1751
rect 930 1751 936 1752
rect 930 1750 931 1751
rect 908 1748 931 1750
rect 908 1746 910 1748
rect 930 1747 931 1748
rect 935 1747 936 1751
rect 1355 1751 1356 1755
rect 1363 1751 1364 1755
rect 1523 1755 1524 1759
rect 1528 1758 1529 1759
rect 1615 1759 1621 1760
rect 1615 1758 1616 1759
rect 1528 1756 1616 1758
rect 1528 1755 1529 1756
rect 1523 1754 1529 1755
rect 1615 1755 1616 1756
rect 1620 1755 1621 1759
rect 1615 1754 1621 1755
rect 1699 1759 1708 1760
rect 1699 1755 1700 1759
rect 1707 1755 1708 1759
rect 1699 1754 1708 1755
rect 1710 1759 1716 1760
rect 1710 1755 1711 1759
rect 1715 1758 1716 1759
rect 1883 1759 1889 1760
rect 1883 1758 1884 1759
rect 1715 1756 1884 1758
rect 1715 1755 1716 1756
rect 1710 1754 1716 1755
rect 1883 1755 1884 1756
rect 1888 1755 1889 1759
rect 2131 1759 2132 1763
rect 2136 1762 2137 1763
rect 2146 1763 2152 1764
rect 2146 1762 2147 1763
rect 2136 1760 2147 1762
rect 2136 1759 2137 1760
rect 2131 1758 2137 1759
rect 2146 1759 2147 1760
rect 2151 1759 2152 1763
rect 2146 1758 2152 1759
rect 2170 1763 2176 1764
rect 2170 1759 2171 1763
rect 2175 1762 2176 1763
rect 2267 1763 2273 1764
rect 2267 1762 2268 1763
rect 2175 1760 2268 1762
rect 2175 1759 2176 1760
rect 2170 1758 2176 1759
rect 2267 1759 2268 1760
rect 2272 1759 2273 1763
rect 2267 1758 2273 1759
rect 2306 1763 2312 1764
rect 2306 1759 2307 1763
rect 2311 1762 2312 1763
rect 2403 1763 2409 1764
rect 2403 1762 2404 1763
rect 2311 1760 2404 1762
rect 2311 1759 2312 1760
rect 2306 1758 2312 1759
rect 2403 1759 2404 1760
rect 2408 1759 2409 1763
rect 2403 1758 2409 1759
rect 2547 1763 2553 1764
rect 2547 1759 2548 1763
rect 2552 1762 2553 1763
rect 2607 1763 2613 1764
rect 2607 1762 2608 1763
rect 2552 1760 2608 1762
rect 2552 1759 2553 1760
rect 2547 1758 2553 1759
rect 2607 1759 2608 1760
rect 2612 1759 2613 1763
rect 2891 1763 2897 1764
rect 2607 1758 2613 1759
rect 2682 1759 2688 1760
rect 1883 1754 1889 1755
rect 2682 1755 2683 1759
rect 2687 1758 2688 1759
rect 2707 1759 2713 1760
rect 2707 1758 2708 1759
rect 2687 1756 2708 1758
rect 2687 1755 2688 1756
rect 2682 1754 2688 1755
rect 2707 1755 2708 1756
rect 2712 1755 2713 1759
rect 2891 1759 2892 1763
rect 2896 1762 2897 1763
rect 2938 1763 2944 1764
rect 2938 1762 2939 1763
rect 2896 1760 2939 1762
rect 2896 1759 2897 1760
rect 2891 1758 2897 1759
rect 2938 1759 2939 1760
rect 2943 1759 2944 1763
rect 2938 1758 2944 1759
rect 3107 1763 3113 1764
rect 3107 1759 3108 1763
rect 3112 1762 3113 1763
rect 3166 1763 3172 1764
rect 3166 1762 3167 1763
rect 3112 1760 3167 1762
rect 3112 1759 3113 1760
rect 3107 1758 3113 1759
rect 3166 1759 3167 1760
rect 3171 1759 3172 1763
rect 3166 1758 3172 1759
rect 3339 1763 3345 1764
rect 3339 1759 3340 1763
rect 3344 1762 3345 1763
rect 3422 1763 3428 1764
rect 3422 1762 3423 1763
rect 3344 1760 3423 1762
rect 3344 1759 3345 1760
rect 3339 1758 3345 1759
rect 3422 1759 3423 1760
rect 3427 1759 3428 1763
rect 3422 1758 3428 1759
rect 3579 1763 3585 1764
rect 3579 1759 3580 1763
rect 3584 1762 3585 1763
rect 3606 1763 3612 1764
rect 3606 1762 3607 1763
rect 3584 1760 3607 1762
rect 3584 1759 3585 1760
rect 3579 1758 3585 1759
rect 3606 1759 3607 1760
rect 3611 1759 3612 1763
rect 3606 1758 3612 1759
rect 3798 1759 3804 1760
rect 2707 1754 2713 1755
rect 3798 1755 3799 1759
rect 3803 1758 3804 1759
rect 3827 1759 3833 1760
rect 3827 1758 3828 1759
rect 3803 1756 3828 1758
rect 3803 1755 3804 1756
rect 3798 1754 3804 1755
rect 3827 1755 3828 1756
rect 3832 1755 3833 1759
rect 3827 1754 3833 1755
rect 1355 1750 1364 1751
rect 2426 1751 2432 1752
rect 930 1746 936 1747
rect 2219 1747 2225 1748
rect 883 1745 910 1746
rect 418 1743 424 1744
rect 379 1741 385 1742
rect 379 1737 380 1741
rect 384 1737 385 1741
rect 418 1739 419 1743
rect 423 1742 424 1743
rect 499 1743 505 1744
rect 499 1742 500 1743
rect 423 1740 500 1742
rect 423 1739 424 1740
rect 418 1738 424 1739
rect 499 1739 500 1740
rect 504 1739 505 1743
rect 499 1738 505 1739
rect 538 1743 544 1744
rect 538 1739 539 1743
rect 543 1742 544 1743
rect 627 1743 633 1744
rect 627 1742 628 1743
rect 543 1740 628 1742
rect 543 1739 544 1740
rect 538 1738 544 1739
rect 627 1739 628 1740
rect 632 1739 633 1743
rect 627 1738 633 1739
rect 666 1743 672 1744
rect 666 1739 667 1743
rect 671 1742 672 1743
rect 755 1743 761 1744
rect 755 1742 756 1743
rect 671 1740 756 1742
rect 671 1739 672 1740
rect 666 1738 672 1739
rect 755 1739 756 1740
rect 760 1739 761 1743
rect 883 1741 884 1745
rect 888 1744 910 1745
rect 888 1741 889 1744
rect 883 1740 889 1741
rect 922 1743 928 1744
rect 755 1738 761 1739
rect 922 1739 923 1743
rect 927 1742 928 1743
rect 1019 1743 1025 1744
rect 1019 1742 1020 1743
rect 927 1740 1020 1742
rect 927 1739 928 1740
rect 922 1738 928 1739
rect 1019 1739 1020 1740
rect 1024 1739 1025 1743
rect 1019 1738 1025 1739
rect 1158 1743 1169 1744
rect 1158 1739 1159 1743
rect 1163 1739 1164 1743
rect 1168 1739 1169 1743
rect 1158 1738 1169 1739
rect 1202 1743 1208 1744
rect 1202 1739 1203 1743
rect 1207 1742 1208 1743
rect 1315 1743 1321 1744
rect 1315 1742 1316 1743
rect 1207 1740 1316 1742
rect 1207 1739 1208 1740
rect 1202 1738 1208 1739
rect 1315 1739 1316 1740
rect 1320 1739 1321 1743
rect 1315 1738 1321 1739
rect 1354 1743 1360 1744
rect 1354 1739 1355 1743
rect 1359 1742 1360 1743
rect 1475 1743 1481 1744
rect 1475 1742 1476 1743
rect 1359 1740 1476 1742
rect 1359 1739 1360 1740
rect 1354 1738 1360 1739
rect 1475 1739 1476 1740
rect 1480 1739 1481 1743
rect 1475 1738 1481 1739
rect 1562 1743 1568 1744
rect 1562 1739 1563 1743
rect 1567 1742 1568 1743
rect 1635 1743 1641 1744
rect 1635 1742 1636 1743
rect 1567 1740 1636 1742
rect 1567 1739 1568 1740
rect 1562 1738 1568 1739
rect 1635 1739 1636 1740
rect 1640 1739 1641 1743
rect 2219 1743 2220 1747
rect 2224 1746 2225 1747
rect 2266 1747 2272 1748
rect 2266 1746 2267 1747
rect 2224 1744 2267 1746
rect 2224 1743 2225 1744
rect 2219 1742 2225 1743
rect 2266 1743 2267 1744
rect 2271 1743 2272 1747
rect 2266 1742 2272 1743
rect 2323 1747 2329 1748
rect 2323 1743 2324 1747
rect 2328 1746 2329 1747
rect 2374 1747 2380 1748
rect 2374 1746 2375 1747
rect 2328 1744 2375 1746
rect 2328 1743 2329 1744
rect 2323 1742 2329 1743
rect 2374 1743 2375 1744
rect 2379 1743 2380 1747
rect 2426 1747 2427 1751
rect 2431 1750 2432 1751
rect 2431 1749 2433 1750
rect 2426 1746 2428 1747
rect 2427 1745 2428 1746
rect 2432 1745 2433 1749
rect 2570 1747 2576 1748
rect 2427 1744 2433 1745
rect 2531 1745 2537 1746
rect 2374 1742 2380 1743
rect 2531 1741 2532 1745
rect 2536 1741 2537 1745
rect 2570 1743 2571 1747
rect 2575 1746 2576 1747
rect 2635 1747 2641 1748
rect 2635 1746 2636 1747
rect 2575 1744 2636 1746
rect 2575 1743 2576 1744
rect 2570 1742 2576 1743
rect 2635 1743 2636 1744
rect 2640 1743 2641 1747
rect 2635 1742 2641 1743
rect 2739 1747 2745 1748
rect 2739 1743 2740 1747
rect 2744 1746 2745 1747
rect 2770 1747 2776 1748
rect 2770 1746 2771 1747
rect 2744 1744 2771 1746
rect 2744 1743 2745 1744
rect 2739 1742 2745 1743
rect 2770 1743 2771 1744
rect 2775 1743 2776 1747
rect 2770 1742 2776 1743
rect 2778 1747 2784 1748
rect 2778 1743 2779 1747
rect 2783 1746 2784 1747
rect 2843 1747 2849 1748
rect 2843 1746 2844 1747
rect 2783 1744 2844 1746
rect 2783 1743 2784 1744
rect 2778 1742 2784 1743
rect 2843 1743 2844 1744
rect 2848 1743 2849 1747
rect 2843 1742 2849 1743
rect 2882 1747 2888 1748
rect 2882 1743 2883 1747
rect 2887 1746 2888 1747
rect 2947 1747 2953 1748
rect 2947 1746 2948 1747
rect 2887 1744 2948 1746
rect 2887 1743 2888 1744
rect 2882 1742 2888 1743
rect 2947 1743 2948 1744
rect 2952 1743 2953 1747
rect 2947 1742 2953 1743
rect 2986 1747 2992 1748
rect 2986 1743 2987 1747
rect 2991 1746 2992 1747
rect 3051 1747 3057 1748
rect 3051 1746 3052 1747
rect 2991 1744 3052 1746
rect 2991 1743 2992 1744
rect 2986 1742 2992 1743
rect 3051 1743 3052 1744
rect 3056 1743 3057 1747
rect 3051 1742 3057 1743
rect 3090 1747 3096 1748
rect 3090 1743 3091 1747
rect 3095 1746 3096 1747
rect 3163 1747 3169 1748
rect 3163 1746 3164 1747
rect 3095 1744 3164 1746
rect 3095 1743 3096 1744
rect 3090 1742 3096 1743
rect 3163 1743 3164 1744
rect 3168 1743 3169 1747
rect 3163 1742 3169 1743
rect 2531 1740 2537 1741
rect 1635 1738 1641 1739
rect 2532 1738 2534 1740
rect 2626 1739 2632 1740
rect 2626 1738 2627 1739
rect 379 1736 385 1737
rect 2532 1736 2627 1738
rect 380 1734 382 1736
rect 738 1735 744 1736
rect 738 1734 739 1735
rect 380 1732 739 1734
rect 738 1731 739 1732
rect 743 1731 744 1735
rect 2626 1735 2627 1736
rect 2631 1735 2632 1739
rect 2626 1734 2632 1735
rect 738 1730 744 1731
rect 2046 1728 2052 1729
rect 3942 1728 3948 1729
rect 110 1724 116 1725
rect 2006 1724 2012 1725
rect 110 1720 111 1724
rect 115 1720 116 1724
rect 110 1719 116 1720
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1719 348 1723
rect 342 1718 348 1719
rect 462 1723 468 1724
rect 462 1719 463 1723
rect 467 1719 468 1723
rect 462 1718 468 1719
rect 590 1723 596 1724
rect 590 1719 591 1723
rect 595 1719 596 1723
rect 590 1718 596 1719
rect 718 1723 724 1724
rect 718 1719 719 1723
rect 723 1719 724 1723
rect 718 1718 724 1719
rect 846 1723 852 1724
rect 846 1719 847 1723
rect 851 1719 852 1723
rect 846 1718 852 1719
rect 982 1723 988 1724
rect 982 1719 983 1723
rect 987 1719 988 1723
rect 982 1718 988 1719
rect 1126 1723 1132 1724
rect 1126 1719 1127 1723
rect 1131 1719 1132 1723
rect 1126 1718 1132 1719
rect 1278 1723 1284 1724
rect 1278 1719 1279 1723
rect 1283 1719 1284 1723
rect 1278 1718 1284 1719
rect 1438 1723 1444 1724
rect 1438 1719 1439 1723
rect 1443 1719 1444 1723
rect 1438 1718 1444 1719
rect 1598 1723 1604 1724
rect 1598 1719 1599 1723
rect 1603 1719 1604 1723
rect 2006 1720 2007 1724
rect 2011 1720 2012 1724
rect 2046 1724 2047 1728
rect 2051 1724 2052 1728
rect 2046 1723 2052 1724
rect 2182 1727 2188 1728
rect 2182 1723 2183 1727
rect 2187 1723 2188 1727
rect 2182 1722 2188 1723
rect 2286 1727 2292 1728
rect 2286 1723 2287 1727
rect 2291 1723 2292 1727
rect 2286 1722 2292 1723
rect 2390 1727 2396 1728
rect 2390 1723 2391 1727
rect 2395 1723 2396 1727
rect 2390 1722 2396 1723
rect 2494 1727 2500 1728
rect 2494 1723 2495 1727
rect 2499 1723 2500 1727
rect 2494 1722 2500 1723
rect 2598 1727 2604 1728
rect 2598 1723 2599 1727
rect 2603 1723 2604 1727
rect 2598 1722 2604 1723
rect 2702 1727 2708 1728
rect 2702 1723 2703 1727
rect 2707 1723 2708 1727
rect 2702 1722 2708 1723
rect 2806 1727 2812 1728
rect 2806 1723 2807 1727
rect 2811 1723 2812 1727
rect 2806 1722 2812 1723
rect 2910 1727 2916 1728
rect 2910 1723 2911 1727
rect 2915 1723 2916 1727
rect 2910 1722 2916 1723
rect 3014 1727 3020 1728
rect 3014 1723 3015 1727
rect 3019 1723 3020 1727
rect 3014 1722 3020 1723
rect 3126 1727 3132 1728
rect 3126 1723 3127 1727
rect 3131 1723 3132 1727
rect 3942 1724 3943 1728
rect 3947 1724 3948 1728
rect 3942 1723 3948 1724
rect 3126 1722 3132 1723
rect 2006 1719 2012 1720
rect 2266 1719 2272 1720
rect 1598 1718 1604 1719
rect 418 1715 424 1716
rect 418 1711 419 1715
rect 423 1711 424 1715
rect 418 1710 424 1711
rect 538 1715 544 1716
rect 538 1711 539 1715
rect 543 1711 544 1715
rect 538 1710 544 1711
rect 666 1715 672 1716
rect 666 1711 667 1715
rect 671 1711 672 1715
rect 666 1710 672 1711
rect 794 1715 800 1716
rect 794 1711 795 1715
rect 799 1711 800 1715
rect 794 1710 800 1711
rect 922 1715 928 1716
rect 922 1711 923 1715
rect 927 1711 928 1715
rect 1202 1715 1208 1716
rect 922 1710 928 1711
rect 1058 1711 1064 1712
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 1058 1707 1059 1711
rect 1063 1707 1064 1711
rect 1202 1711 1203 1715
rect 1207 1711 1208 1715
rect 1202 1710 1208 1711
rect 1354 1715 1360 1716
rect 1354 1711 1355 1715
rect 1359 1711 1360 1715
rect 1354 1710 1360 1711
rect 1362 1715 1368 1716
rect 1362 1711 1363 1715
rect 1367 1714 1368 1715
rect 1582 1715 1588 1716
rect 1367 1712 1481 1714
rect 1367 1711 1368 1712
rect 1362 1710 1368 1711
rect 1582 1711 1583 1715
rect 1587 1714 1588 1715
rect 2258 1715 2264 1716
rect 1587 1712 1641 1714
rect 1587 1711 1588 1712
rect 1582 1710 1588 1711
rect 2046 1711 2052 1712
rect 1058 1706 1064 1707
rect 2006 1707 2012 1708
rect 110 1702 116 1703
rect 342 1704 348 1705
rect 342 1700 343 1704
rect 347 1700 348 1704
rect 342 1699 348 1700
rect 462 1704 468 1705
rect 462 1700 463 1704
rect 467 1700 468 1704
rect 462 1699 468 1700
rect 590 1704 596 1705
rect 590 1700 591 1704
rect 595 1700 596 1704
rect 590 1699 596 1700
rect 718 1704 724 1705
rect 718 1700 719 1704
rect 723 1700 724 1704
rect 718 1699 724 1700
rect 846 1704 852 1705
rect 846 1700 847 1704
rect 851 1700 852 1704
rect 846 1699 852 1700
rect 982 1704 988 1705
rect 982 1700 983 1704
rect 987 1700 988 1704
rect 982 1699 988 1700
rect 1126 1704 1132 1705
rect 1126 1700 1127 1704
rect 1131 1700 1132 1704
rect 1126 1699 1132 1700
rect 1278 1704 1284 1705
rect 1278 1700 1279 1704
rect 1283 1700 1284 1704
rect 1278 1699 1284 1700
rect 1438 1704 1444 1705
rect 1438 1700 1439 1704
rect 1443 1700 1444 1704
rect 1438 1699 1444 1700
rect 1598 1704 1604 1705
rect 1598 1700 1599 1704
rect 1603 1700 1604 1704
rect 2006 1703 2007 1707
rect 2011 1703 2012 1707
rect 2046 1707 2047 1711
rect 2051 1707 2052 1711
rect 2258 1711 2259 1715
rect 2263 1711 2264 1715
rect 2266 1715 2267 1719
rect 2271 1718 2272 1719
rect 2374 1719 2380 1720
rect 2271 1716 2329 1718
rect 2271 1715 2272 1716
rect 2266 1714 2272 1715
rect 2374 1715 2375 1719
rect 2379 1718 2380 1719
rect 2570 1719 2576 1720
rect 2379 1716 2433 1718
rect 2379 1715 2380 1716
rect 2374 1714 2380 1715
rect 2570 1715 2571 1719
rect 2575 1715 2576 1719
rect 2682 1719 2688 1720
rect 2682 1718 2683 1719
rect 2677 1716 2683 1718
rect 2570 1714 2576 1715
rect 2682 1715 2683 1716
rect 2687 1715 2688 1719
rect 2682 1714 2688 1715
rect 2778 1719 2784 1720
rect 2778 1715 2779 1719
rect 2783 1715 2784 1719
rect 2778 1714 2784 1715
rect 2882 1719 2888 1720
rect 2882 1715 2883 1719
rect 2887 1715 2888 1719
rect 2882 1714 2888 1715
rect 2986 1719 2992 1720
rect 2986 1715 2987 1719
rect 2991 1715 2992 1719
rect 2986 1714 2992 1715
rect 3090 1719 3096 1720
rect 3090 1715 3091 1719
rect 3095 1715 3096 1719
rect 3090 1714 3096 1715
rect 3202 1715 3208 1716
rect 2258 1710 2264 1711
rect 3202 1711 3203 1715
rect 3207 1711 3208 1715
rect 3202 1710 3208 1711
rect 3942 1711 3948 1712
rect 2046 1706 2052 1707
rect 2182 1708 2188 1709
rect 2182 1704 2183 1708
rect 2187 1704 2188 1708
rect 2182 1703 2188 1704
rect 2286 1708 2292 1709
rect 2286 1704 2287 1708
rect 2291 1704 2292 1708
rect 2286 1703 2292 1704
rect 2390 1708 2396 1709
rect 2390 1704 2391 1708
rect 2395 1704 2396 1708
rect 2390 1703 2396 1704
rect 2494 1708 2500 1709
rect 2494 1704 2495 1708
rect 2499 1704 2500 1708
rect 2494 1703 2500 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2702 1708 2708 1709
rect 2702 1704 2703 1708
rect 2707 1704 2708 1708
rect 2702 1703 2708 1704
rect 2806 1708 2812 1709
rect 2806 1704 2807 1708
rect 2811 1704 2812 1708
rect 2806 1703 2812 1704
rect 2910 1708 2916 1709
rect 2910 1704 2911 1708
rect 2915 1704 2916 1708
rect 2910 1703 2916 1704
rect 3014 1708 3020 1709
rect 3014 1704 3015 1708
rect 3019 1704 3020 1708
rect 3014 1703 3020 1704
rect 3126 1708 3132 1709
rect 3126 1704 3127 1708
rect 3131 1704 3132 1708
rect 3942 1707 3943 1711
rect 3947 1707 3948 1711
rect 3942 1706 3948 1707
rect 3126 1703 3132 1704
rect 2006 1702 2012 1703
rect 1598 1699 1604 1700
rect 2230 1648 2236 1649
rect 2046 1645 2052 1646
rect 2046 1641 2047 1645
rect 2051 1641 2052 1645
rect 2230 1644 2231 1648
rect 2235 1644 2236 1648
rect 2230 1643 2236 1644
rect 2366 1648 2372 1649
rect 2366 1644 2367 1648
rect 2371 1644 2372 1648
rect 2366 1643 2372 1644
rect 2518 1648 2524 1649
rect 2518 1644 2519 1648
rect 2523 1644 2524 1648
rect 2518 1643 2524 1644
rect 2678 1648 2684 1649
rect 2678 1644 2679 1648
rect 2683 1644 2684 1648
rect 2678 1643 2684 1644
rect 2846 1648 2852 1649
rect 2846 1644 2847 1648
rect 2851 1644 2852 1648
rect 2846 1643 2852 1644
rect 3022 1648 3028 1649
rect 3022 1644 3023 1648
rect 3027 1644 3028 1648
rect 3022 1643 3028 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3526 1648 3532 1649
rect 3526 1644 3527 1648
rect 3531 1644 3532 1648
rect 3526 1643 3532 1644
rect 3694 1648 3700 1649
rect 3694 1644 3695 1648
rect 3699 1644 3700 1648
rect 3694 1643 3700 1644
rect 3838 1648 3844 1649
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 3942 1645 3948 1646
rect 158 1640 164 1641
rect 110 1637 116 1638
rect 110 1633 111 1637
rect 115 1633 116 1637
rect 158 1636 159 1640
rect 163 1636 164 1640
rect 158 1635 164 1636
rect 294 1640 300 1641
rect 294 1636 295 1640
rect 299 1636 300 1640
rect 294 1635 300 1636
rect 454 1640 460 1641
rect 454 1636 455 1640
rect 459 1636 460 1640
rect 454 1635 460 1636
rect 622 1640 628 1641
rect 622 1636 623 1640
rect 627 1636 628 1640
rect 622 1635 628 1636
rect 798 1640 804 1641
rect 798 1636 799 1640
rect 803 1636 804 1640
rect 798 1635 804 1636
rect 982 1640 988 1641
rect 982 1636 983 1640
rect 987 1636 988 1640
rect 982 1635 988 1636
rect 1166 1640 1172 1641
rect 1166 1636 1167 1640
rect 1171 1636 1172 1640
rect 1166 1635 1172 1636
rect 1350 1640 1356 1641
rect 1350 1636 1351 1640
rect 1355 1636 1356 1640
rect 1350 1635 1356 1636
rect 1542 1640 1548 1641
rect 1542 1636 1543 1640
rect 1547 1636 1548 1640
rect 1542 1635 1548 1636
rect 1734 1640 1740 1641
rect 2046 1640 2052 1641
rect 3942 1641 3943 1645
rect 3947 1641 3948 1645
rect 3942 1640 3948 1641
rect 1734 1636 1735 1640
rect 1739 1636 1740 1640
rect 2306 1639 2312 1640
rect 1734 1635 1740 1636
rect 2006 1637 2012 1638
rect 110 1632 116 1633
rect 2006 1633 2007 1637
rect 2011 1633 2012 1637
rect 2306 1635 2307 1639
rect 2311 1635 2312 1639
rect 2306 1634 2312 1635
rect 2442 1639 2448 1640
rect 2442 1635 2443 1639
rect 2447 1635 2448 1639
rect 2442 1634 2448 1635
rect 2594 1639 2600 1640
rect 2594 1635 2595 1639
rect 2599 1635 2600 1639
rect 2594 1634 2600 1635
rect 2626 1639 2632 1640
rect 2626 1635 2627 1639
rect 2631 1638 2632 1639
rect 2762 1639 2768 1640
rect 2631 1636 2721 1638
rect 2631 1635 2632 1636
rect 2626 1634 2632 1635
rect 2762 1635 2763 1639
rect 2767 1638 2768 1639
rect 3106 1639 3112 1640
rect 3106 1638 3107 1639
rect 2767 1636 2889 1638
rect 3101 1636 3107 1638
rect 2767 1635 2768 1636
rect 2762 1634 2768 1635
rect 3106 1635 3107 1636
rect 3111 1635 3112 1639
rect 3106 1634 3112 1635
rect 3127 1639 3133 1640
rect 3127 1635 3128 1639
rect 3132 1638 3133 1639
rect 3434 1639 3440 1640
rect 3132 1636 3233 1638
rect 3132 1635 3133 1636
rect 3127 1634 3133 1635
rect 3434 1635 3435 1639
rect 3439 1635 3440 1639
rect 3434 1634 3440 1635
rect 3602 1639 3608 1640
rect 3602 1635 3603 1639
rect 3607 1635 3608 1639
rect 3602 1634 3608 1635
rect 3639 1639 3645 1640
rect 3639 1635 3640 1639
rect 3644 1638 3645 1639
rect 3906 1639 3912 1640
rect 3644 1636 3737 1638
rect 3644 1635 3645 1636
rect 3639 1634 3645 1635
rect 3906 1635 3907 1639
rect 3911 1635 3912 1639
rect 3906 1634 3912 1635
rect 2006 1632 2012 1633
rect 234 1631 240 1632
rect 234 1627 235 1631
rect 239 1627 240 1631
rect 234 1626 240 1627
rect 370 1631 376 1632
rect 370 1627 371 1631
rect 375 1627 376 1631
rect 370 1626 376 1627
rect 530 1631 536 1632
rect 530 1627 531 1631
rect 535 1627 536 1631
rect 530 1626 536 1627
rect 698 1631 704 1632
rect 698 1627 699 1631
rect 703 1627 704 1631
rect 698 1626 704 1627
rect 738 1631 744 1632
rect 738 1627 739 1631
rect 743 1630 744 1631
rect 1050 1631 1056 1632
rect 743 1628 841 1630
rect 743 1627 744 1628
rect 738 1626 744 1627
rect 1050 1627 1051 1631
rect 1055 1627 1056 1631
rect 1050 1626 1056 1627
rect 1158 1631 1164 1632
rect 1158 1627 1159 1631
rect 1163 1630 1164 1631
rect 1295 1631 1301 1632
rect 1163 1628 1209 1630
rect 1163 1627 1164 1628
rect 1158 1626 1164 1627
rect 1295 1627 1296 1631
rect 1300 1630 1301 1631
rect 1618 1631 1624 1632
rect 1300 1628 1393 1630
rect 1300 1627 1301 1628
rect 1295 1626 1301 1627
rect 1618 1627 1619 1631
rect 1623 1627 1624 1631
rect 1618 1626 1624 1627
rect 1802 1631 1808 1632
rect 1802 1627 1803 1631
rect 1807 1627 1808 1631
rect 2230 1629 2236 1630
rect 1802 1626 1808 1627
rect 2046 1628 2052 1629
rect 2046 1624 2047 1628
rect 2051 1624 2052 1628
rect 2230 1625 2231 1629
rect 2235 1625 2236 1629
rect 2230 1624 2236 1625
rect 2366 1629 2372 1630
rect 2366 1625 2367 1629
rect 2371 1625 2372 1629
rect 2366 1624 2372 1625
rect 2518 1629 2524 1630
rect 2518 1625 2519 1629
rect 2523 1625 2524 1629
rect 2518 1624 2524 1625
rect 2678 1629 2684 1630
rect 2678 1625 2679 1629
rect 2683 1625 2684 1629
rect 2678 1624 2684 1625
rect 2846 1629 2852 1630
rect 2846 1625 2847 1629
rect 2851 1625 2852 1629
rect 2846 1624 2852 1625
rect 3022 1629 3028 1630
rect 3022 1625 3023 1629
rect 3027 1625 3028 1629
rect 3022 1624 3028 1625
rect 3190 1629 3196 1630
rect 3190 1625 3191 1629
rect 3195 1625 3196 1629
rect 3190 1624 3196 1625
rect 3358 1629 3364 1630
rect 3358 1625 3359 1629
rect 3363 1625 3364 1629
rect 3358 1624 3364 1625
rect 3526 1629 3532 1630
rect 3526 1625 3527 1629
rect 3531 1625 3532 1629
rect 3526 1624 3532 1625
rect 3694 1629 3700 1630
rect 3694 1625 3695 1629
rect 3699 1625 3700 1629
rect 3694 1624 3700 1625
rect 3838 1629 3844 1630
rect 3838 1625 3839 1629
rect 3843 1625 3844 1629
rect 3838 1624 3844 1625
rect 3942 1628 3948 1629
rect 3942 1624 3943 1628
rect 3947 1624 3948 1628
rect 2046 1623 2052 1624
rect 3942 1623 3948 1624
rect 158 1621 164 1622
rect 110 1620 116 1621
rect 110 1616 111 1620
rect 115 1616 116 1620
rect 158 1617 159 1621
rect 163 1617 164 1621
rect 158 1616 164 1617
rect 294 1621 300 1622
rect 294 1617 295 1621
rect 299 1617 300 1621
rect 294 1616 300 1617
rect 454 1621 460 1622
rect 454 1617 455 1621
rect 459 1617 460 1621
rect 454 1616 460 1617
rect 622 1621 628 1622
rect 622 1617 623 1621
rect 627 1617 628 1621
rect 622 1616 628 1617
rect 798 1621 804 1622
rect 798 1617 799 1621
rect 803 1617 804 1621
rect 798 1616 804 1617
rect 982 1621 988 1622
rect 982 1617 983 1621
rect 987 1617 988 1621
rect 982 1616 988 1617
rect 1166 1621 1172 1622
rect 1166 1617 1167 1621
rect 1171 1617 1172 1621
rect 1166 1616 1172 1617
rect 1350 1621 1356 1622
rect 1350 1617 1351 1621
rect 1355 1617 1356 1621
rect 1350 1616 1356 1617
rect 1542 1621 1548 1622
rect 1542 1617 1543 1621
rect 1547 1617 1548 1621
rect 1542 1616 1548 1617
rect 1734 1621 1740 1622
rect 1734 1617 1735 1621
rect 1739 1617 1740 1621
rect 1734 1616 1740 1617
rect 2006 1620 2012 1621
rect 2006 1616 2007 1620
rect 2011 1616 2012 1620
rect 110 1615 116 1616
rect 2006 1615 2012 1616
rect 2258 1611 2264 1612
rect 234 1607 240 1608
rect 234 1603 235 1607
rect 239 1606 240 1607
rect 2258 1607 2259 1611
rect 2263 1610 2264 1611
rect 2267 1611 2273 1612
rect 2267 1610 2268 1611
rect 2263 1608 2268 1610
rect 2263 1607 2264 1608
rect 2258 1606 2264 1607
rect 2267 1607 2268 1608
rect 2272 1607 2273 1611
rect 2267 1606 2273 1607
rect 2306 1611 2312 1612
rect 2306 1607 2307 1611
rect 2311 1610 2312 1611
rect 2403 1611 2409 1612
rect 2403 1610 2404 1611
rect 2311 1608 2404 1610
rect 2311 1607 2312 1608
rect 2306 1606 2312 1607
rect 2403 1607 2404 1608
rect 2408 1607 2409 1611
rect 2403 1606 2409 1607
rect 2442 1611 2448 1612
rect 2442 1607 2443 1611
rect 2447 1610 2448 1611
rect 2555 1611 2561 1612
rect 2555 1610 2556 1611
rect 2447 1608 2556 1610
rect 2447 1607 2448 1608
rect 2442 1606 2448 1607
rect 2555 1607 2556 1608
rect 2560 1607 2561 1611
rect 2555 1606 2561 1607
rect 2715 1611 2721 1612
rect 2715 1607 2716 1611
rect 2720 1610 2721 1611
rect 2762 1611 2768 1612
rect 2762 1610 2763 1611
rect 2720 1608 2763 1610
rect 2720 1607 2721 1608
rect 2715 1606 2721 1607
rect 2762 1607 2763 1608
rect 2767 1607 2768 1611
rect 3059 1611 3065 1612
rect 2762 1606 2768 1607
rect 2786 1607 2792 1608
rect 239 1604 321 1606
rect 239 1603 240 1604
rect 234 1602 240 1603
rect 319 1602 321 1604
rect 331 1603 337 1604
rect 331 1602 332 1603
rect 319 1600 332 1602
rect 195 1599 201 1600
rect 195 1595 196 1599
rect 200 1598 201 1599
rect 331 1599 332 1600
rect 336 1599 337 1603
rect 331 1598 337 1599
rect 370 1603 376 1604
rect 370 1599 371 1603
rect 375 1602 376 1603
rect 491 1603 497 1604
rect 491 1602 492 1603
rect 375 1600 492 1602
rect 375 1599 376 1600
rect 370 1598 376 1599
rect 491 1599 492 1600
rect 496 1599 497 1603
rect 491 1598 497 1599
rect 530 1603 536 1604
rect 530 1599 531 1603
rect 535 1602 536 1603
rect 659 1603 665 1604
rect 659 1602 660 1603
rect 535 1600 660 1602
rect 535 1599 536 1600
rect 530 1598 536 1599
rect 659 1599 660 1600
rect 664 1599 665 1603
rect 659 1598 665 1599
rect 698 1603 704 1604
rect 698 1599 699 1603
rect 703 1602 704 1603
rect 835 1603 841 1604
rect 835 1602 836 1603
rect 703 1600 836 1602
rect 703 1599 704 1600
rect 698 1598 704 1599
rect 835 1599 836 1600
rect 840 1599 841 1603
rect 835 1598 841 1599
rect 1019 1603 1025 1604
rect 1019 1599 1020 1603
rect 1024 1602 1025 1603
rect 1058 1603 1064 1604
rect 1058 1602 1059 1603
rect 1024 1600 1059 1602
rect 1024 1599 1025 1600
rect 1019 1598 1025 1599
rect 1058 1599 1059 1600
rect 1063 1599 1064 1603
rect 1058 1598 1064 1599
rect 1203 1603 1209 1604
rect 1203 1599 1204 1603
rect 1208 1602 1209 1603
rect 1295 1603 1301 1604
rect 1295 1602 1296 1603
rect 1208 1600 1296 1602
rect 1208 1599 1209 1600
rect 1203 1598 1209 1599
rect 1295 1599 1296 1600
rect 1300 1599 1301 1603
rect 1579 1603 1588 1604
rect 1295 1598 1301 1599
rect 1387 1599 1393 1600
rect 200 1596 321 1598
rect 200 1595 201 1596
rect 195 1594 201 1595
rect 319 1594 321 1596
rect 738 1595 744 1596
rect 738 1594 739 1595
rect 319 1592 739 1594
rect 738 1591 739 1592
rect 743 1591 744 1595
rect 1387 1595 1388 1599
rect 1392 1598 1393 1599
rect 1442 1599 1448 1600
rect 1442 1598 1443 1599
rect 1392 1596 1443 1598
rect 1392 1595 1393 1596
rect 1387 1594 1393 1595
rect 1442 1595 1443 1596
rect 1447 1595 1448 1599
rect 1579 1599 1580 1603
rect 1587 1599 1588 1603
rect 1579 1598 1588 1599
rect 1618 1603 1624 1604
rect 1618 1599 1619 1603
rect 1623 1602 1624 1603
rect 1771 1603 1777 1604
rect 1771 1602 1772 1603
rect 1623 1600 1772 1602
rect 1623 1599 1624 1600
rect 1618 1598 1624 1599
rect 1771 1599 1772 1600
rect 1776 1599 1777 1603
rect 2786 1603 2787 1607
rect 2791 1606 2792 1607
rect 2883 1607 2889 1608
rect 2883 1606 2884 1607
rect 2791 1604 2884 1606
rect 2791 1603 2792 1604
rect 2786 1602 2792 1603
rect 2883 1603 2884 1604
rect 2888 1603 2889 1607
rect 3059 1607 3060 1611
rect 3064 1610 3065 1611
rect 3127 1611 3133 1612
rect 3127 1610 3128 1611
rect 3064 1608 3128 1610
rect 3064 1607 3065 1608
rect 3059 1606 3065 1607
rect 3127 1607 3128 1608
rect 3132 1607 3133 1611
rect 3127 1606 3133 1607
rect 3202 1611 3208 1612
rect 3202 1607 3203 1611
rect 3207 1610 3208 1611
rect 3227 1611 3233 1612
rect 3227 1610 3228 1611
rect 3207 1608 3228 1610
rect 3207 1607 3208 1608
rect 3202 1606 3208 1607
rect 3227 1607 3228 1608
rect 3232 1607 3233 1611
rect 3434 1611 3440 1612
rect 3227 1606 3233 1607
rect 3395 1607 3404 1608
rect 2883 1602 2889 1603
rect 3395 1603 3396 1607
rect 3403 1603 3404 1607
rect 3434 1607 3435 1611
rect 3439 1610 3440 1611
rect 3563 1611 3569 1612
rect 3563 1610 3564 1611
rect 3439 1608 3564 1610
rect 3439 1607 3440 1608
rect 3434 1606 3440 1607
rect 3563 1607 3564 1608
rect 3568 1607 3569 1611
rect 3563 1606 3569 1607
rect 3602 1611 3608 1612
rect 3602 1607 3603 1611
rect 3607 1610 3608 1611
rect 3731 1611 3737 1612
rect 3731 1610 3732 1611
rect 3607 1608 3732 1610
rect 3607 1607 3608 1608
rect 3602 1606 3608 1607
rect 3731 1607 3732 1608
rect 3736 1607 3737 1611
rect 3731 1606 3737 1607
rect 3875 1611 3881 1612
rect 3875 1607 3876 1611
rect 3880 1610 3881 1611
rect 3914 1611 3920 1612
rect 3914 1610 3915 1611
rect 3880 1608 3915 1610
rect 3880 1607 3881 1608
rect 3875 1606 3881 1607
rect 3914 1607 3915 1608
rect 3919 1607 3920 1611
rect 3914 1606 3920 1607
rect 3395 1602 3404 1603
rect 1771 1598 1777 1599
rect 1442 1594 1448 1595
rect 738 1590 744 1591
rect 171 1587 177 1588
rect 171 1583 172 1587
rect 176 1586 177 1587
rect 202 1587 208 1588
rect 202 1586 203 1587
rect 176 1584 203 1586
rect 176 1583 177 1584
rect 171 1582 177 1583
rect 202 1583 203 1584
rect 207 1583 208 1587
rect 202 1582 208 1583
rect 210 1587 216 1588
rect 210 1583 211 1587
rect 215 1586 216 1587
rect 291 1587 297 1588
rect 291 1586 292 1587
rect 215 1584 292 1586
rect 215 1583 216 1584
rect 210 1582 216 1583
rect 291 1583 292 1584
rect 296 1583 297 1587
rect 291 1582 297 1583
rect 330 1587 336 1588
rect 330 1583 331 1587
rect 335 1586 336 1587
rect 459 1587 465 1588
rect 459 1586 460 1587
rect 335 1584 460 1586
rect 335 1583 336 1584
rect 330 1582 336 1583
rect 459 1583 460 1584
rect 464 1583 465 1587
rect 459 1582 465 1583
rect 498 1587 504 1588
rect 498 1583 499 1587
rect 503 1586 504 1587
rect 643 1587 649 1588
rect 643 1586 644 1587
rect 503 1584 644 1586
rect 503 1583 504 1584
rect 498 1582 504 1583
rect 643 1583 644 1584
rect 648 1583 649 1587
rect 643 1582 649 1583
rect 682 1587 688 1588
rect 682 1583 683 1587
rect 687 1586 688 1587
rect 835 1587 841 1588
rect 835 1586 836 1587
rect 687 1584 836 1586
rect 687 1583 688 1584
rect 682 1582 688 1583
rect 835 1583 836 1584
rect 840 1583 841 1587
rect 835 1582 841 1583
rect 1027 1587 1033 1588
rect 1027 1583 1028 1587
rect 1032 1586 1033 1587
rect 1050 1587 1056 1588
rect 1050 1586 1051 1587
rect 1032 1584 1051 1586
rect 1032 1583 1033 1584
rect 1027 1582 1033 1583
rect 1050 1583 1051 1584
rect 1055 1583 1056 1587
rect 1050 1582 1056 1583
rect 1219 1587 1225 1588
rect 1219 1583 1220 1587
rect 1224 1586 1225 1587
rect 1250 1587 1256 1588
rect 1250 1586 1251 1587
rect 1224 1584 1251 1586
rect 1224 1583 1225 1584
rect 1219 1582 1225 1583
rect 1250 1583 1251 1584
rect 1255 1583 1256 1587
rect 1250 1582 1256 1583
rect 1258 1587 1264 1588
rect 1258 1583 1259 1587
rect 1263 1586 1264 1587
rect 1403 1587 1409 1588
rect 1403 1586 1404 1587
rect 1263 1584 1404 1586
rect 1263 1583 1264 1584
rect 1258 1582 1264 1583
rect 1403 1583 1404 1584
rect 1408 1583 1409 1587
rect 1403 1582 1409 1583
rect 1587 1587 1593 1588
rect 1587 1583 1588 1587
rect 1592 1586 1593 1587
rect 1634 1587 1640 1588
rect 1634 1586 1635 1587
rect 1592 1584 1635 1586
rect 1592 1583 1593 1584
rect 1587 1582 1593 1583
rect 1634 1583 1635 1584
rect 1639 1583 1640 1587
rect 1634 1582 1640 1583
rect 1771 1587 1777 1588
rect 1771 1583 1772 1587
rect 1776 1586 1777 1587
rect 1802 1587 1808 1588
rect 1802 1586 1803 1587
rect 1776 1584 1803 1586
rect 1776 1583 1777 1584
rect 1771 1582 1777 1583
rect 1802 1583 1803 1584
rect 1807 1583 1808 1587
rect 1978 1587 1984 1588
rect 1802 1582 1808 1583
rect 1939 1585 1945 1586
rect 1939 1581 1940 1585
rect 1944 1581 1945 1585
rect 1978 1583 1979 1587
rect 1983 1586 1984 1587
rect 2107 1587 2113 1588
rect 2107 1586 2108 1587
rect 1983 1584 2108 1586
rect 1983 1583 1984 1584
rect 1978 1582 1984 1583
rect 2107 1583 2108 1584
rect 2112 1583 2113 1587
rect 2107 1582 2113 1583
rect 2146 1587 2152 1588
rect 2146 1583 2147 1587
rect 2151 1586 2152 1587
rect 2307 1587 2313 1588
rect 2307 1586 2308 1587
rect 2151 1584 2308 1586
rect 2151 1583 2152 1584
rect 2146 1582 2152 1583
rect 2307 1583 2308 1584
rect 2312 1583 2313 1587
rect 2307 1582 2313 1583
rect 2346 1587 2352 1588
rect 2346 1583 2347 1587
rect 2351 1586 2352 1587
rect 2531 1587 2537 1588
rect 2531 1586 2532 1587
rect 2351 1584 2532 1586
rect 2351 1583 2352 1584
rect 2346 1582 2352 1583
rect 2531 1583 2532 1584
rect 2536 1583 2537 1587
rect 2531 1582 2537 1583
rect 2594 1587 2600 1588
rect 2594 1583 2595 1587
rect 2599 1586 2600 1587
rect 2747 1587 2753 1588
rect 2747 1586 2748 1587
rect 2599 1584 2748 1586
rect 2599 1583 2600 1584
rect 2594 1582 2600 1583
rect 2747 1583 2748 1584
rect 2752 1583 2753 1587
rect 2747 1582 2753 1583
rect 2947 1587 2953 1588
rect 2947 1583 2948 1587
rect 2952 1586 2953 1587
rect 2994 1587 3000 1588
rect 2994 1586 2995 1587
rect 2952 1584 2995 1586
rect 2952 1583 2953 1584
rect 2947 1582 2953 1583
rect 2994 1583 2995 1584
rect 2999 1583 3000 1587
rect 2994 1582 3000 1583
rect 3106 1587 3112 1588
rect 3106 1583 3107 1587
rect 3111 1586 3112 1587
rect 3131 1587 3137 1588
rect 3131 1586 3132 1587
rect 3111 1584 3132 1586
rect 3111 1583 3112 1584
rect 3106 1582 3112 1583
rect 3131 1583 3132 1584
rect 3136 1583 3137 1587
rect 3131 1582 3137 1583
rect 3202 1587 3208 1588
rect 3202 1583 3203 1587
rect 3207 1586 3208 1587
rect 3299 1587 3305 1588
rect 3299 1586 3300 1587
rect 3207 1584 3300 1586
rect 3207 1583 3208 1584
rect 3202 1582 3208 1583
rect 3299 1583 3300 1584
rect 3304 1583 3305 1587
rect 3299 1582 3305 1583
rect 3338 1587 3344 1588
rect 3338 1583 3339 1587
rect 3343 1586 3344 1587
rect 3459 1587 3465 1588
rect 3459 1586 3460 1587
rect 3343 1584 3460 1586
rect 3343 1583 3344 1584
rect 3338 1582 3344 1583
rect 3459 1583 3460 1584
rect 3464 1583 3465 1587
rect 3459 1582 3465 1583
rect 3603 1587 3609 1588
rect 3603 1583 3604 1587
rect 3608 1586 3609 1587
rect 3639 1587 3645 1588
rect 3639 1586 3640 1587
rect 3608 1584 3640 1586
rect 3608 1583 3609 1584
rect 3603 1582 3609 1583
rect 3639 1583 3640 1584
rect 3644 1583 3645 1587
rect 3639 1582 3645 1583
rect 3747 1587 3753 1588
rect 3747 1583 3748 1587
rect 3752 1586 3753 1587
rect 3806 1587 3812 1588
rect 3806 1586 3807 1587
rect 3752 1584 3807 1586
rect 3752 1583 3753 1584
rect 3747 1582 3753 1583
rect 3806 1583 3807 1584
rect 3811 1583 3812 1587
rect 3806 1582 3812 1583
rect 3875 1587 3881 1588
rect 3875 1583 3876 1587
rect 3880 1586 3881 1587
rect 3906 1587 3912 1588
rect 3906 1586 3907 1587
rect 3880 1584 3907 1586
rect 3880 1583 3881 1584
rect 3875 1582 3881 1583
rect 3906 1583 3907 1584
rect 3911 1583 3912 1587
rect 3906 1582 3912 1583
rect 1939 1580 1945 1581
rect 1762 1579 1768 1580
rect 1762 1575 1763 1579
rect 1767 1578 1768 1579
rect 1940 1578 1942 1580
rect 1767 1576 1942 1578
rect 1767 1575 1768 1576
rect 1762 1574 1768 1575
rect 110 1568 116 1569
rect 2006 1568 2012 1569
rect 110 1564 111 1568
rect 115 1564 116 1568
rect 110 1563 116 1564
rect 134 1567 140 1568
rect 134 1563 135 1567
rect 139 1563 140 1567
rect 134 1562 140 1563
rect 254 1567 260 1568
rect 254 1563 255 1567
rect 259 1563 260 1567
rect 254 1562 260 1563
rect 422 1567 428 1568
rect 422 1563 423 1567
rect 427 1563 428 1567
rect 422 1562 428 1563
rect 606 1567 612 1568
rect 606 1563 607 1567
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 798 1567 804 1568
rect 798 1563 799 1567
rect 803 1563 804 1567
rect 798 1562 804 1563
rect 990 1567 996 1568
rect 990 1563 991 1567
rect 995 1563 996 1567
rect 990 1562 996 1563
rect 1182 1567 1188 1568
rect 1182 1563 1183 1567
rect 1187 1563 1188 1567
rect 1182 1562 1188 1563
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 1550 1567 1556 1568
rect 1550 1563 1551 1567
rect 1555 1563 1556 1567
rect 1550 1562 1556 1563
rect 1734 1567 1740 1568
rect 1734 1563 1735 1567
rect 1739 1563 1740 1567
rect 1734 1562 1740 1563
rect 1902 1567 1908 1568
rect 1902 1563 1903 1567
rect 1907 1563 1908 1567
rect 2006 1564 2007 1568
rect 2011 1564 2012 1568
rect 2006 1563 2012 1564
rect 2046 1568 2052 1569
rect 3942 1568 3948 1569
rect 2046 1564 2047 1568
rect 2051 1564 2052 1568
rect 2046 1563 2052 1564
rect 2070 1567 2076 1568
rect 2070 1563 2071 1567
rect 2075 1563 2076 1567
rect 1902 1562 1908 1563
rect 2070 1562 2076 1563
rect 2270 1567 2276 1568
rect 2270 1563 2271 1567
rect 2275 1563 2276 1567
rect 2270 1562 2276 1563
rect 2494 1567 2500 1568
rect 2494 1563 2495 1567
rect 2499 1563 2500 1567
rect 2494 1562 2500 1563
rect 2710 1567 2716 1568
rect 2710 1563 2711 1567
rect 2715 1563 2716 1567
rect 2710 1562 2716 1563
rect 2910 1567 2916 1568
rect 2910 1563 2911 1567
rect 2915 1563 2916 1567
rect 2910 1562 2916 1563
rect 3094 1567 3100 1568
rect 3094 1563 3095 1567
rect 3099 1563 3100 1567
rect 3094 1562 3100 1563
rect 3262 1567 3268 1568
rect 3262 1563 3263 1567
rect 3267 1563 3268 1567
rect 3262 1562 3268 1563
rect 3422 1567 3428 1568
rect 3422 1563 3423 1567
rect 3427 1563 3428 1567
rect 3422 1562 3428 1563
rect 3566 1567 3572 1568
rect 3566 1563 3567 1567
rect 3571 1563 3572 1567
rect 3566 1562 3572 1563
rect 3710 1567 3716 1568
rect 3710 1563 3711 1567
rect 3715 1563 3716 1567
rect 3710 1562 3716 1563
rect 3838 1567 3844 1568
rect 3838 1563 3839 1567
rect 3843 1563 3844 1567
rect 3942 1564 3943 1568
rect 3947 1564 3948 1568
rect 3942 1563 3948 1564
rect 3838 1562 3844 1563
rect 210 1559 216 1560
rect 210 1555 211 1559
rect 215 1555 216 1559
rect 210 1554 216 1555
rect 330 1559 336 1560
rect 330 1555 331 1559
rect 335 1555 336 1559
rect 330 1554 336 1555
rect 498 1559 504 1560
rect 498 1555 499 1559
rect 503 1555 504 1559
rect 498 1554 504 1555
rect 682 1559 688 1560
rect 682 1555 683 1559
rect 687 1555 688 1559
rect 682 1554 688 1555
rect 738 1559 744 1560
rect 738 1555 739 1559
rect 743 1558 744 1559
rect 1258 1559 1264 1560
rect 743 1556 841 1558
rect 743 1555 744 1556
rect 738 1554 744 1555
rect 1066 1555 1072 1556
rect 110 1551 116 1552
rect 110 1547 111 1551
rect 115 1547 116 1551
rect 1066 1551 1067 1555
rect 1071 1551 1072 1555
rect 1258 1555 1259 1559
rect 1263 1555 1264 1559
rect 1258 1554 1264 1555
rect 1442 1559 1448 1560
rect 1442 1555 1443 1559
rect 1447 1555 1448 1559
rect 1442 1554 1448 1555
rect 1454 1559 1460 1560
rect 1454 1555 1455 1559
rect 1459 1558 1460 1559
rect 1634 1559 1640 1560
rect 1459 1556 1593 1558
rect 1459 1555 1460 1556
rect 1454 1554 1460 1555
rect 1634 1555 1635 1559
rect 1639 1558 1640 1559
rect 1978 1559 1984 1560
rect 1639 1556 1777 1558
rect 1639 1555 1640 1556
rect 1634 1554 1640 1555
rect 1978 1555 1979 1559
rect 1983 1555 1984 1559
rect 1978 1554 1984 1555
rect 2146 1559 2152 1560
rect 2146 1555 2147 1559
rect 2151 1555 2152 1559
rect 2146 1554 2152 1555
rect 2346 1559 2352 1560
rect 2346 1555 2347 1559
rect 2351 1555 2352 1559
rect 2346 1554 2352 1555
rect 2418 1559 2424 1560
rect 2418 1555 2419 1559
rect 2423 1558 2424 1559
rect 2786 1559 2792 1560
rect 2423 1556 2537 1558
rect 2423 1555 2424 1556
rect 2418 1554 2424 1555
rect 2786 1555 2787 1559
rect 2791 1555 2792 1559
rect 2786 1554 2792 1555
rect 2895 1559 2901 1560
rect 2895 1555 2896 1559
rect 2900 1558 2901 1559
rect 2994 1559 3000 1560
rect 2900 1556 2953 1558
rect 2900 1555 2901 1556
rect 2895 1554 2901 1555
rect 2994 1555 2995 1559
rect 2999 1558 3000 1559
rect 3338 1559 3344 1560
rect 2999 1556 3137 1558
rect 2999 1555 3000 1556
rect 2994 1554 3000 1555
rect 3338 1555 3339 1559
rect 3343 1555 3344 1559
rect 3338 1554 3344 1555
rect 3398 1559 3404 1560
rect 3398 1555 3399 1559
rect 3403 1558 3404 1559
rect 3506 1559 3512 1560
rect 3403 1556 3465 1558
rect 3403 1555 3404 1556
rect 3398 1554 3404 1555
rect 3506 1555 3507 1559
rect 3511 1558 3512 1559
rect 3798 1559 3804 1560
rect 3798 1558 3799 1559
rect 3511 1556 3609 1558
rect 3789 1556 3799 1558
rect 3511 1555 3512 1556
rect 3506 1554 3512 1555
rect 3798 1555 3799 1556
rect 3803 1555 3804 1559
rect 3798 1554 3804 1555
rect 3806 1559 3812 1560
rect 3806 1555 3807 1559
rect 3811 1558 3812 1559
rect 3811 1556 3881 1558
rect 3811 1555 3812 1556
rect 3806 1554 3812 1555
rect 1066 1550 1072 1551
rect 2006 1551 2012 1552
rect 110 1546 116 1547
rect 134 1548 140 1549
rect 134 1544 135 1548
rect 139 1544 140 1548
rect 134 1543 140 1544
rect 254 1548 260 1549
rect 254 1544 255 1548
rect 259 1544 260 1548
rect 254 1543 260 1544
rect 422 1548 428 1549
rect 422 1544 423 1548
rect 427 1544 428 1548
rect 422 1543 428 1544
rect 606 1548 612 1549
rect 606 1544 607 1548
rect 611 1544 612 1548
rect 606 1543 612 1544
rect 798 1548 804 1549
rect 798 1544 799 1548
rect 803 1544 804 1548
rect 798 1543 804 1544
rect 990 1548 996 1549
rect 990 1544 991 1548
rect 995 1544 996 1548
rect 990 1543 996 1544
rect 1182 1548 1188 1549
rect 1182 1544 1183 1548
rect 1187 1544 1188 1548
rect 1182 1543 1188 1544
rect 1366 1548 1372 1549
rect 1366 1544 1367 1548
rect 1371 1544 1372 1548
rect 1366 1543 1372 1544
rect 1550 1548 1556 1549
rect 1550 1544 1551 1548
rect 1555 1544 1556 1548
rect 1550 1543 1556 1544
rect 1734 1548 1740 1549
rect 1734 1544 1735 1548
rect 1739 1544 1740 1548
rect 1734 1543 1740 1544
rect 1902 1548 1908 1549
rect 1902 1544 1903 1548
rect 1907 1544 1908 1548
rect 2006 1547 2007 1551
rect 2011 1547 2012 1551
rect 2006 1546 2012 1547
rect 2046 1551 2052 1552
rect 2046 1547 2047 1551
rect 2051 1547 2052 1551
rect 3942 1551 3948 1552
rect 2046 1546 2052 1547
rect 2070 1548 2076 1549
rect 1902 1543 1908 1544
rect 2070 1544 2071 1548
rect 2075 1544 2076 1548
rect 2070 1543 2076 1544
rect 2270 1548 2276 1549
rect 2270 1544 2271 1548
rect 2275 1544 2276 1548
rect 2270 1543 2276 1544
rect 2494 1548 2500 1549
rect 2494 1544 2495 1548
rect 2499 1544 2500 1548
rect 2494 1543 2500 1544
rect 2710 1548 2716 1549
rect 2710 1544 2711 1548
rect 2715 1544 2716 1548
rect 2710 1543 2716 1544
rect 2910 1548 2916 1549
rect 2910 1544 2911 1548
rect 2915 1544 2916 1548
rect 2910 1543 2916 1544
rect 3094 1548 3100 1549
rect 3094 1544 3095 1548
rect 3099 1544 3100 1548
rect 3094 1543 3100 1544
rect 3262 1548 3268 1549
rect 3262 1544 3263 1548
rect 3267 1544 3268 1548
rect 3262 1543 3268 1544
rect 3422 1548 3428 1549
rect 3422 1544 3423 1548
rect 3427 1544 3428 1548
rect 3422 1543 3428 1544
rect 3566 1548 3572 1549
rect 3566 1544 3567 1548
rect 3571 1544 3572 1548
rect 3566 1543 3572 1544
rect 3710 1548 3716 1549
rect 3710 1544 3711 1548
rect 3715 1544 3716 1548
rect 3710 1543 3716 1544
rect 3838 1548 3844 1549
rect 3838 1544 3839 1548
rect 3843 1544 3844 1548
rect 3942 1547 3943 1551
rect 3947 1547 3948 1551
rect 3942 1546 3948 1547
rect 3838 1543 3844 1544
rect 202 1491 208 1492
rect 202 1487 203 1491
rect 207 1490 208 1491
rect 207 1488 646 1490
rect 207 1487 208 1488
rect 202 1486 208 1487
rect 134 1484 140 1485
rect 110 1481 116 1482
rect 110 1477 111 1481
rect 115 1477 116 1481
rect 134 1480 135 1484
rect 139 1480 140 1484
rect 134 1479 140 1480
rect 246 1484 252 1485
rect 246 1480 247 1484
rect 251 1480 252 1484
rect 246 1479 252 1480
rect 398 1484 404 1485
rect 398 1480 399 1484
rect 403 1480 404 1484
rect 398 1479 404 1480
rect 558 1484 564 1485
rect 558 1480 559 1484
rect 563 1480 564 1484
rect 558 1479 564 1480
rect 110 1476 116 1477
rect 210 1475 216 1476
rect 210 1471 211 1475
rect 215 1471 216 1475
rect 210 1470 216 1471
rect 322 1475 328 1476
rect 322 1471 323 1475
rect 327 1471 328 1475
rect 322 1470 328 1471
rect 474 1475 480 1476
rect 474 1471 475 1475
rect 479 1471 480 1475
rect 474 1470 480 1471
rect 634 1475 640 1476
rect 634 1471 635 1475
rect 639 1471 640 1475
rect 644 1474 646 1488
rect 2070 1488 2076 1489
rect 2046 1485 2052 1486
rect 718 1484 724 1485
rect 718 1480 719 1484
rect 723 1480 724 1484
rect 718 1479 724 1480
rect 878 1484 884 1485
rect 878 1480 879 1484
rect 883 1480 884 1484
rect 878 1479 884 1480
rect 1038 1484 1044 1485
rect 1038 1480 1039 1484
rect 1043 1480 1044 1484
rect 1038 1479 1044 1480
rect 1182 1484 1188 1485
rect 1182 1480 1183 1484
rect 1187 1480 1188 1484
rect 1182 1479 1188 1480
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1446 1484 1452 1485
rect 1446 1480 1447 1484
rect 1451 1480 1452 1484
rect 1446 1479 1452 1480
rect 1566 1484 1572 1485
rect 1566 1480 1567 1484
rect 1571 1480 1572 1484
rect 1566 1479 1572 1480
rect 1686 1484 1692 1485
rect 1686 1480 1687 1484
rect 1691 1480 1692 1484
rect 1686 1479 1692 1480
rect 1806 1484 1812 1485
rect 1806 1480 1807 1484
rect 1811 1480 1812 1484
rect 1806 1479 1812 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 2006 1481 2012 1482
rect 2006 1477 2007 1481
rect 2011 1477 2012 1481
rect 2046 1481 2047 1485
rect 2051 1481 2052 1485
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 2430 1488 2436 1489
rect 2430 1484 2431 1488
rect 2435 1484 2436 1488
rect 2430 1483 2436 1484
rect 2790 1488 2796 1489
rect 2790 1484 2791 1488
rect 2795 1484 2796 1488
rect 2790 1483 2796 1484
rect 3126 1488 3132 1489
rect 3126 1484 3127 1488
rect 3131 1484 3132 1488
rect 3126 1483 3132 1484
rect 3462 1488 3468 1489
rect 3462 1484 3463 1488
rect 3467 1484 3468 1488
rect 3462 1483 3468 1484
rect 3798 1488 3804 1489
rect 3798 1484 3799 1488
rect 3803 1484 3804 1488
rect 3798 1483 3804 1484
rect 3942 1485 3948 1486
rect 2046 1480 2052 1481
rect 3942 1481 3943 1485
rect 3947 1481 3948 1485
rect 3942 1480 3948 1481
rect 2006 1476 2012 1477
rect 2054 1479 2060 1480
rect 954 1475 960 1476
rect 644 1472 761 1474
rect 634 1470 640 1471
rect 954 1471 955 1475
rect 959 1471 960 1475
rect 954 1470 960 1471
rect 975 1475 981 1476
rect 975 1471 976 1475
rect 980 1474 981 1475
rect 1250 1475 1256 1476
rect 980 1472 1081 1474
rect 980 1471 981 1472
rect 975 1470 981 1471
rect 1250 1471 1251 1475
rect 1255 1471 1256 1475
rect 1250 1470 1256 1471
rect 1394 1475 1400 1476
rect 1394 1471 1395 1475
rect 1399 1471 1400 1475
rect 1394 1470 1400 1471
rect 1522 1475 1528 1476
rect 1522 1471 1523 1475
rect 1527 1471 1528 1475
rect 1522 1470 1528 1471
rect 1642 1475 1648 1476
rect 1642 1471 1643 1475
rect 1647 1471 1648 1475
rect 1642 1470 1648 1471
rect 1762 1475 1768 1476
rect 1762 1471 1763 1475
rect 1767 1471 1768 1475
rect 1762 1470 1768 1471
rect 1882 1475 1888 1476
rect 1882 1471 1883 1475
rect 1887 1471 1888 1475
rect 1882 1470 1888 1471
rect 1894 1475 1900 1476
rect 1894 1471 1895 1475
rect 1899 1474 1900 1475
rect 2054 1475 2055 1479
rect 2059 1478 2060 1479
rect 2718 1479 2724 1480
rect 2718 1478 2719 1479
rect 2059 1476 2113 1478
rect 2509 1476 2719 1478
rect 2059 1475 2060 1476
rect 2054 1474 2060 1475
rect 2718 1475 2719 1476
rect 2723 1475 2724 1479
rect 2718 1474 2724 1475
rect 2866 1479 2872 1480
rect 2866 1475 2867 1479
rect 2871 1475 2872 1479
rect 2866 1474 2872 1475
rect 3202 1479 3208 1480
rect 3202 1475 3203 1479
rect 3207 1475 3208 1479
rect 3202 1474 3208 1475
rect 3538 1479 3544 1480
rect 3538 1475 3539 1479
rect 3543 1475 3544 1479
rect 3538 1474 3544 1475
rect 3866 1479 3872 1480
rect 3866 1475 3867 1479
rect 3871 1475 3872 1479
rect 3866 1474 3872 1475
rect 1899 1472 1945 1474
rect 1899 1471 1900 1472
rect 1894 1470 1900 1471
rect 2070 1469 2076 1470
rect 2046 1468 2052 1469
rect 134 1465 140 1466
rect 110 1464 116 1465
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 134 1461 135 1465
rect 139 1461 140 1465
rect 134 1460 140 1461
rect 246 1465 252 1466
rect 246 1461 247 1465
rect 251 1461 252 1465
rect 246 1460 252 1461
rect 398 1465 404 1466
rect 398 1461 399 1465
rect 403 1461 404 1465
rect 398 1460 404 1461
rect 558 1465 564 1466
rect 558 1461 559 1465
rect 563 1461 564 1465
rect 558 1460 564 1461
rect 718 1465 724 1466
rect 718 1461 719 1465
rect 723 1461 724 1465
rect 718 1460 724 1461
rect 878 1465 884 1466
rect 878 1461 879 1465
rect 883 1461 884 1465
rect 878 1460 884 1461
rect 1038 1465 1044 1466
rect 1038 1461 1039 1465
rect 1043 1461 1044 1465
rect 1038 1460 1044 1461
rect 1182 1465 1188 1466
rect 1182 1461 1183 1465
rect 1187 1461 1188 1465
rect 1182 1460 1188 1461
rect 1318 1465 1324 1466
rect 1318 1461 1319 1465
rect 1323 1461 1324 1465
rect 1318 1460 1324 1461
rect 1446 1465 1452 1466
rect 1446 1461 1447 1465
rect 1451 1461 1452 1465
rect 1446 1460 1452 1461
rect 1566 1465 1572 1466
rect 1566 1461 1567 1465
rect 1571 1461 1572 1465
rect 1566 1460 1572 1461
rect 1686 1465 1692 1466
rect 1686 1461 1687 1465
rect 1691 1461 1692 1465
rect 1686 1460 1692 1461
rect 1806 1465 1812 1466
rect 1806 1461 1807 1465
rect 1811 1461 1812 1465
rect 1806 1460 1812 1461
rect 1902 1465 1908 1466
rect 1902 1461 1903 1465
rect 1907 1461 1908 1465
rect 1902 1460 1908 1461
rect 2006 1464 2012 1465
rect 2006 1460 2007 1464
rect 2011 1460 2012 1464
rect 2046 1464 2047 1468
rect 2051 1464 2052 1468
rect 2070 1465 2071 1469
rect 2075 1465 2076 1469
rect 2070 1464 2076 1465
rect 2430 1469 2436 1470
rect 2430 1465 2431 1469
rect 2435 1465 2436 1469
rect 2430 1464 2436 1465
rect 2790 1469 2796 1470
rect 2790 1465 2791 1469
rect 2795 1465 2796 1469
rect 2790 1464 2796 1465
rect 3126 1469 3132 1470
rect 3126 1465 3127 1469
rect 3131 1465 3132 1469
rect 3126 1464 3132 1465
rect 3462 1469 3468 1470
rect 3462 1465 3463 1469
rect 3467 1465 3468 1469
rect 3462 1464 3468 1465
rect 3798 1469 3804 1470
rect 3798 1465 3799 1469
rect 3803 1465 3804 1469
rect 3798 1464 3804 1465
rect 3942 1468 3948 1469
rect 3942 1464 3943 1468
rect 3947 1464 3948 1468
rect 2046 1463 2052 1464
rect 3942 1463 3948 1464
rect 110 1459 116 1460
rect 2006 1459 2012 1460
rect 2895 1459 2901 1460
rect 2895 1458 2896 1459
rect 2656 1456 2896 1458
rect 1454 1455 1460 1456
rect 1454 1454 1455 1455
rect 1388 1452 1455 1454
rect 210 1447 216 1448
rect 171 1443 177 1444
rect 171 1439 172 1443
rect 176 1442 177 1443
rect 210 1443 211 1447
rect 215 1446 216 1447
rect 283 1447 289 1448
rect 283 1446 284 1447
rect 215 1444 284 1446
rect 215 1443 216 1444
rect 210 1442 216 1443
rect 283 1443 284 1444
rect 288 1443 289 1447
rect 283 1442 289 1443
rect 322 1447 328 1448
rect 322 1443 323 1447
rect 327 1446 328 1447
rect 435 1447 441 1448
rect 435 1446 436 1447
rect 327 1444 436 1446
rect 327 1443 328 1444
rect 322 1442 328 1443
rect 435 1443 436 1444
rect 440 1443 441 1447
rect 435 1442 441 1443
rect 474 1447 480 1448
rect 474 1443 475 1447
rect 479 1446 480 1447
rect 595 1447 601 1448
rect 595 1446 596 1447
rect 479 1444 596 1446
rect 479 1443 480 1444
rect 474 1442 480 1443
rect 595 1443 596 1444
rect 600 1443 601 1447
rect 595 1442 601 1443
rect 634 1447 640 1448
rect 634 1443 635 1447
rect 639 1446 640 1447
rect 755 1447 761 1448
rect 755 1446 756 1447
rect 639 1444 756 1446
rect 639 1443 640 1444
rect 634 1442 640 1443
rect 755 1443 756 1444
rect 760 1443 761 1447
rect 755 1442 761 1443
rect 915 1447 921 1448
rect 915 1443 916 1447
rect 920 1446 921 1447
rect 975 1447 981 1448
rect 975 1446 976 1447
rect 920 1444 976 1446
rect 920 1443 921 1444
rect 915 1442 921 1443
rect 975 1443 976 1444
rect 980 1443 981 1447
rect 975 1442 981 1443
rect 1066 1447 1072 1448
rect 1066 1443 1067 1447
rect 1071 1446 1072 1447
rect 1075 1447 1081 1448
rect 1075 1446 1076 1447
rect 1071 1444 1076 1446
rect 1071 1443 1072 1444
rect 1066 1442 1072 1443
rect 1075 1443 1076 1444
rect 1080 1443 1081 1447
rect 1355 1447 1361 1448
rect 1075 1442 1081 1443
rect 1219 1443 1225 1444
rect 176 1439 178 1442
rect 171 1438 178 1439
rect 210 1439 216 1440
rect 210 1438 211 1439
rect 176 1436 211 1438
rect 210 1435 211 1436
rect 215 1435 216 1439
rect 1219 1439 1220 1443
rect 1224 1442 1225 1443
rect 1242 1443 1248 1444
rect 1242 1442 1243 1443
rect 1224 1440 1243 1442
rect 1224 1439 1225 1440
rect 1219 1438 1225 1439
rect 1242 1439 1243 1440
rect 1247 1439 1248 1443
rect 1355 1443 1356 1447
rect 1360 1446 1361 1447
rect 1388 1446 1390 1452
rect 1454 1451 1455 1452
rect 1459 1451 1460 1455
rect 1454 1450 1460 1451
rect 2107 1451 2113 1452
rect 1360 1444 1390 1446
rect 1394 1447 1400 1448
rect 1360 1443 1361 1444
rect 1355 1442 1361 1443
rect 1394 1443 1395 1447
rect 1399 1446 1400 1447
rect 1483 1447 1489 1448
rect 1483 1446 1484 1447
rect 1399 1444 1484 1446
rect 1399 1443 1400 1444
rect 1394 1442 1400 1443
rect 1483 1443 1484 1444
rect 1488 1443 1489 1447
rect 1483 1442 1489 1443
rect 1522 1447 1528 1448
rect 1522 1443 1523 1447
rect 1527 1446 1528 1447
rect 1603 1447 1609 1448
rect 1603 1446 1604 1447
rect 1527 1444 1604 1446
rect 1527 1443 1528 1444
rect 1522 1442 1528 1443
rect 1603 1443 1604 1444
rect 1608 1443 1609 1447
rect 1603 1442 1609 1443
rect 1642 1447 1648 1448
rect 1642 1443 1643 1447
rect 1647 1446 1648 1447
rect 1723 1447 1729 1448
rect 1723 1446 1724 1447
rect 1647 1444 1724 1446
rect 1647 1443 1648 1444
rect 1642 1442 1648 1443
rect 1723 1443 1724 1444
rect 1728 1443 1729 1447
rect 1723 1442 1729 1443
rect 1843 1447 1849 1448
rect 1843 1443 1844 1447
rect 1848 1446 1849 1447
rect 1894 1447 1900 1448
rect 1894 1446 1895 1447
rect 1848 1444 1895 1446
rect 1848 1443 1849 1444
rect 1843 1442 1849 1443
rect 1894 1443 1895 1444
rect 1899 1443 1900 1447
rect 1894 1442 1900 1443
rect 1939 1447 1945 1448
rect 1939 1443 1940 1447
rect 1944 1446 1945 1447
rect 2054 1447 2060 1448
rect 2054 1446 2055 1447
rect 1944 1444 2055 1446
rect 1944 1443 1945 1444
rect 1939 1442 1945 1443
rect 2054 1443 2055 1444
rect 2059 1443 2060 1447
rect 2107 1447 2108 1451
rect 2112 1450 2113 1451
rect 2418 1451 2424 1452
rect 2418 1450 2419 1451
rect 2112 1448 2419 1450
rect 2112 1447 2113 1448
rect 2107 1446 2113 1447
rect 2418 1447 2419 1448
rect 2423 1447 2424 1451
rect 2418 1446 2424 1447
rect 2467 1451 2473 1452
rect 2467 1447 2468 1451
rect 2472 1450 2473 1451
rect 2656 1450 2658 1456
rect 2895 1455 2896 1456
rect 2900 1455 2901 1459
rect 2895 1454 2901 1455
rect 2472 1448 2658 1450
rect 2718 1451 2724 1452
rect 2472 1447 2473 1448
rect 2467 1446 2473 1447
rect 2718 1447 2719 1451
rect 2723 1450 2724 1451
rect 2827 1451 2833 1452
rect 2827 1450 2828 1451
rect 2723 1448 2828 1450
rect 2723 1447 2724 1448
rect 2718 1446 2724 1447
rect 2827 1447 2828 1448
rect 2832 1447 2833 1451
rect 3499 1451 3508 1452
rect 2827 1446 2833 1447
rect 3163 1447 3172 1448
rect 2054 1442 2060 1443
rect 3163 1443 3164 1447
rect 3171 1443 3172 1447
rect 3499 1447 3500 1451
rect 3507 1447 3508 1451
rect 3499 1446 3508 1447
rect 3538 1451 3544 1452
rect 3538 1447 3539 1451
rect 3543 1450 3544 1451
rect 3835 1451 3841 1452
rect 3835 1450 3836 1451
rect 3543 1448 3836 1450
rect 3543 1447 3544 1448
rect 3538 1446 3544 1447
rect 3835 1447 3836 1448
rect 3840 1447 3841 1451
rect 3835 1446 3841 1447
rect 3163 1442 3172 1443
rect 1242 1438 1248 1439
rect 210 1434 216 1435
rect 171 1431 177 1432
rect 171 1427 172 1431
rect 176 1430 177 1431
rect 218 1431 224 1432
rect 218 1430 219 1431
rect 176 1428 219 1430
rect 176 1427 177 1428
rect 171 1426 177 1427
rect 218 1427 219 1428
rect 223 1427 224 1431
rect 218 1426 224 1427
rect 299 1431 305 1432
rect 299 1427 300 1431
rect 304 1430 305 1431
rect 366 1431 372 1432
rect 366 1430 367 1431
rect 304 1428 367 1430
rect 304 1427 305 1428
rect 299 1426 305 1427
rect 366 1427 367 1428
rect 371 1427 372 1431
rect 578 1431 584 1432
rect 366 1426 372 1427
rect 467 1429 473 1430
rect 467 1425 468 1429
rect 472 1425 473 1429
rect 578 1427 579 1431
rect 583 1430 584 1431
rect 643 1431 649 1432
rect 643 1430 644 1431
rect 583 1428 644 1430
rect 583 1427 584 1428
rect 578 1426 584 1427
rect 643 1427 644 1428
rect 648 1427 649 1431
rect 643 1426 649 1427
rect 682 1431 688 1432
rect 682 1427 683 1431
rect 687 1430 688 1431
rect 827 1431 833 1432
rect 827 1430 828 1431
rect 687 1428 828 1430
rect 687 1427 688 1428
rect 682 1426 688 1427
rect 827 1427 828 1428
rect 832 1427 833 1431
rect 827 1426 833 1427
rect 954 1431 960 1432
rect 954 1427 955 1431
rect 959 1430 960 1431
rect 1011 1431 1017 1432
rect 1011 1430 1012 1431
rect 959 1428 1012 1430
rect 959 1427 960 1428
rect 954 1426 960 1427
rect 1011 1427 1012 1428
rect 1016 1427 1017 1431
rect 1011 1426 1017 1427
rect 1050 1431 1056 1432
rect 1050 1427 1051 1431
rect 1055 1430 1056 1431
rect 1195 1431 1201 1432
rect 1195 1430 1196 1431
rect 1055 1428 1196 1430
rect 1055 1427 1056 1428
rect 1050 1426 1056 1427
rect 1195 1427 1196 1428
rect 1200 1427 1201 1431
rect 1195 1426 1201 1427
rect 1387 1431 1393 1432
rect 1387 1427 1388 1431
rect 1392 1430 1393 1431
rect 1434 1431 1440 1432
rect 1434 1430 1435 1431
rect 1392 1428 1435 1430
rect 1392 1427 1393 1428
rect 1387 1426 1393 1427
rect 1434 1427 1435 1428
rect 1439 1427 1440 1431
rect 1434 1426 1440 1427
rect 1579 1431 1585 1432
rect 1579 1427 1580 1431
rect 1584 1430 1585 1431
rect 1626 1431 1632 1432
rect 1626 1430 1627 1431
rect 1584 1428 1627 1430
rect 1584 1427 1585 1428
rect 1579 1426 1585 1427
rect 1626 1427 1627 1428
rect 1631 1427 1632 1431
rect 1626 1426 1632 1427
rect 1742 1431 1748 1432
rect 1742 1427 1743 1431
rect 1747 1430 1748 1431
rect 1771 1431 1777 1432
rect 1771 1430 1772 1431
rect 1747 1428 1772 1430
rect 1747 1427 1748 1428
rect 1742 1426 1748 1427
rect 1771 1427 1772 1428
rect 1776 1427 1777 1431
rect 1771 1426 1777 1427
rect 1882 1431 1888 1432
rect 1882 1427 1883 1431
rect 1887 1430 1888 1431
rect 1939 1431 1945 1432
rect 1939 1430 1940 1431
rect 1887 1428 1940 1430
rect 1887 1427 1888 1428
rect 1882 1426 1888 1427
rect 1939 1427 1940 1428
rect 1944 1427 1945 1431
rect 1939 1426 1945 1427
rect 1978 1427 1984 1428
rect 467 1424 473 1425
rect 468 1422 470 1424
rect 690 1423 696 1424
rect 690 1422 691 1423
rect 468 1420 691 1422
rect 690 1419 691 1420
rect 695 1419 696 1423
rect 1978 1423 1979 1427
rect 1983 1426 1984 1427
rect 2107 1427 2113 1428
rect 2107 1426 2108 1427
rect 1983 1424 2108 1426
rect 1983 1423 1984 1424
rect 1978 1422 1984 1423
rect 2107 1423 2108 1424
rect 2112 1423 2113 1427
rect 2107 1422 2113 1423
rect 2146 1427 2152 1428
rect 2146 1423 2147 1427
rect 2151 1426 2152 1427
rect 2307 1427 2313 1428
rect 2307 1426 2308 1427
rect 2151 1424 2308 1426
rect 2151 1423 2152 1424
rect 2146 1422 2152 1423
rect 2307 1423 2308 1424
rect 2312 1423 2313 1427
rect 2307 1422 2313 1423
rect 2346 1427 2352 1428
rect 2346 1423 2347 1427
rect 2351 1426 2352 1427
rect 2531 1427 2537 1428
rect 2531 1426 2532 1427
rect 2351 1424 2532 1426
rect 2351 1423 2352 1424
rect 2346 1422 2352 1423
rect 2531 1423 2532 1424
rect 2536 1423 2537 1427
rect 2531 1422 2537 1423
rect 2570 1427 2576 1428
rect 2570 1423 2571 1427
rect 2575 1426 2576 1427
rect 2747 1427 2753 1428
rect 2747 1426 2748 1427
rect 2575 1424 2748 1426
rect 2575 1423 2576 1424
rect 2570 1422 2576 1423
rect 2747 1423 2748 1424
rect 2752 1423 2753 1427
rect 2747 1422 2753 1423
rect 2866 1427 2872 1428
rect 2866 1423 2867 1427
rect 2871 1426 2872 1427
rect 2947 1427 2953 1428
rect 2947 1426 2948 1427
rect 2871 1424 2948 1426
rect 2871 1423 2872 1424
rect 2866 1422 2872 1423
rect 2947 1423 2948 1424
rect 2952 1423 2953 1427
rect 2947 1422 2953 1423
rect 2986 1427 2992 1428
rect 2986 1423 2987 1427
rect 2991 1426 2992 1427
rect 3131 1427 3137 1428
rect 3131 1426 3132 1427
rect 2991 1424 3132 1426
rect 2991 1423 2992 1424
rect 2986 1422 2992 1423
rect 3131 1423 3132 1424
rect 3136 1423 3137 1427
rect 3131 1422 3137 1423
rect 3307 1427 3313 1428
rect 3307 1423 3308 1427
rect 3312 1426 3313 1427
rect 3354 1427 3360 1428
rect 3354 1426 3355 1427
rect 3312 1424 3355 1426
rect 3312 1423 3313 1424
rect 3307 1422 3313 1423
rect 3354 1423 3355 1424
rect 3359 1423 3360 1427
rect 3354 1422 3360 1423
rect 3475 1427 3481 1428
rect 3475 1423 3476 1427
rect 3480 1426 3481 1427
rect 3506 1427 3512 1428
rect 3506 1426 3507 1427
rect 3480 1424 3507 1426
rect 3480 1423 3481 1424
rect 3475 1422 3481 1423
rect 3506 1423 3507 1424
rect 3511 1423 3512 1427
rect 3506 1422 3512 1423
rect 3522 1427 3528 1428
rect 3522 1423 3523 1427
rect 3527 1426 3528 1427
rect 3643 1427 3649 1428
rect 3643 1426 3644 1427
rect 3527 1424 3644 1426
rect 3527 1423 3528 1424
rect 3522 1422 3528 1423
rect 3643 1423 3644 1424
rect 3648 1423 3649 1427
rect 3643 1422 3649 1423
rect 3819 1427 3825 1428
rect 3819 1423 3820 1427
rect 3824 1426 3825 1427
rect 3866 1427 3872 1428
rect 3866 1426 3867 1427
rect 3824 1424 3867 1426
rect 3824 1423 3825 1424
rect 3819 1422 3825 1423
rect 3866 1423 3867 1424
rect 3871 1423 3872 1427
rect 3866 1422 3872 1423
rect 690 1418 696 1419
rect 110 1412 116 1413
rect 2006 1412 2012 1413
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 110 1407 116 1408
rect 134 1411 140 1412
rect 134 1407 135 1411
rect 139 1407 140 1411
rect 134 1406 140 1407
rect 262 1411 268 1412
rect 262 1407 263 1411
rect 267 1407 268 1411
rect 262 1406 268 1407
rect 430 1411 436 1412
rect 430 1407 431 1411
rect 435 1407 436 1411
rect 430 1406 436 1407
rect 606 1411 612 1412
rect 606 1407 607 1411
rect 611 1407 612 1411
rect 606 1406 612 1407
rect 790 1411 796 1412
rect 790 1407 791 1411
rect 795 1407 796 1411
rect 790 1406 796 1407
rect 974 1411 980 1412
rect 974 1407 975 1411
rect 979 1407 980 1411
rect 974 1406 980 1407
rect 1158 1411 1164 1412
rect 1158 1407 1159 1411
rect 1163 1407 1164 1411
rect 1158 1406 1164 1407
rect 1350 1411 1356 1412
rect 1350 1407 1351 1411
rect 1355 1407 1356 1411
rect 1350 1406 1356 1407
rect 1542 1411 1548 1412
rect 1542 1407 1543 1411
rect 1547 1407 1548 1411
rect 1542 1406 1548 1407
rect 1734 1411 1740 1412
rect 1734 1407 1735 1411
rect 1739 1407 1740 1411
rect 1734 1406 1740 1407
rect 1902 1411 1908 1412
rect 1902 1407 1903 1411
rect 1907 1407 1908 1411
rect 2006 1408 2007 1412
rect 2011 1408 2012 1412
rect 2006 1407 2012 1408
rect 2046 1408 2052 1409
rect 3942 1408 3948 1409
rect 1902 1406 1908 1407
rect 2046 1404 2047 1408
rect 2051 1404 2052 1408
rect 210 1403 216 1404
rect 210 1399 211 1403
rect 215 1399 216 1403
rect 210 1398 216 1399
rect 218 1403 224 1404
rect 218 1399 219 1403
rect 223 1402 224 1403
rect 366 1403 372 1404
rect 223 1400 305 1402
rect 223 1399 224 1400
rect 218 1398 224 1399
rect 366 1399 367 1403
rect 371 1402 372 1403
rect 682 1403 688 1404
rect 371 1400 473 1402
rect 371 1399 372 1400
rect 366 1398 372 1399
rect 682 1399 683 1403
rect 687 1399 688 1403
rect 682 1398 688 1399
rect 690 1403 696 1404
rect 690 1399 691 1403
rect 695 1402 696 1403
rect 1050 1403 1056 1404
rect 695 1400 833 1402
rect 695 1399 696 1400
rect 690 1398 696 1399
rect 1050 1399 1051 1403
rect 1055 1399 1056 1403
rect 1050 1398 1056 1399
rect 1082 1403 1088 1404
rect 1082 1399 1083 1403
rect 1087 1402 1088 1403
rect 1242 1403 1248 1404
rect 1087 1400 1201 1402
rect 1087 1399 1088 1400
rect 1082 1398 1088 1399
rect 1242 1399 1243 1403
rect 1247 1402 1248 1403
rect 1434 1403 1440 1404
rect 1247 1400 1393 1402
rect 1247 1399 1248 1400
rect 1242 1398 1248 1399
rect 1434 1399 1435 1403
rect 1439 1402 1440 1403
rect 1626 1403 1632 1404
rect 1439 1400 1585 1402
rect 1439 1399 1440 1400
rect 1434 1398 1440 1399
rect 1626 1399 1627 1403
rect 1631 1402 1632 1403
rect 1978 1403 1984 1404
rect 2046 1403 2052 1404
rect 2070 1407 2076 1408
rect 2070 1403 2071 1407
rect 2075 1403 2076 1407
rect 1631 1400 1777 1402
rect 1631 1399 1632 1400
rect 1626 1398 1632 1399
rect 1978 1399 1979 1403
rect 1983 1399 1984 1403
rect 2070 1402 2076 1403
rect 2270 1407 2276 1408
rect 2270 1403 2271 1407
rect 2275 1403 2276 1407
rect 2270 1402 2276 1403
rect 2494 1407 2500 1408
rect 2494 1403 2495 1407
rect 2499 1403 2500 1407
rect 2494 1402 2500 1403
rect 2710 1407 2716 1408
rect 2710 1403 2711 1407
rect 2715 1403 2716 1407
rect 2710 1402 2716 1403
rect 2910 1407 2916 1408
rect 2910 1403 2911 1407
rect 2915 1403 2916 1407
rect 2910 1402 2916 1403
rect 3094 1407 3100 1408
rect 3094 1403 3095 1407
rect 3099 1403 3100 1407
rect 3094 1402 3100 1403
rect 3270 1407 3276 1408
rect 3270 1403 3271 1407
rect 3275 1403 3276 1407
rect 3270 1402 3276 1403
rect 3438 1407 3444 1408
rect 3438 1403 3439 1407
rect 3443 1403 3444 1407
rect 3606 1407 3612 1408
rect 3438 1402 3444 1403
rect 3506 1403 3512 1404
rect 1978 1398 1984 1399
rect 2146 1399 2152 1400
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 2006 1395 2012 1396
rect 110 1390 116 1391
rect 134 1392 140 1393
rect 134 1388 135 1392
rect 139 1388 140 1392
rect 134 1387 140 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 430 1392 436 1393
rect 430 1388 431 1392
rect 435 1388 436 1392
rect 430 1387 436 1388
rect 606 1392 612 1393
rect 606 1388 607 1392
rect 611 1388 612 1392
rect 606 1387 612 1388
rect 790 1392 796 1393
rect 790 1388 791 1392
rect 795 1388 796 1392
rect 790 1387 796 1388
rect 974 1392 980 1393
rect 974 1388 975 1392
rect 979 1388 980 1392
rect 974 1387 980 1388
rect 1158 1392 1164 1393
rect 1158 1388 1159 1392
rect 1163 1388 1164 1392
rect 1158 1387 1164 1388
rect 1350 1392 1356 1393
rect 1350 1388 1351 1392
rect 1355 1388 1356 1392
rect 1350 1387 1356 1388
rect 1542 1392 1548 1393
rect 1542 1388 1543 1392
rect 1547 1388 1548 1392
rect 1542 1387 1548 1388
rect 1734 1392 1740 1393
rect 1734 1388 1735 1392
rect 1739 1388 1740 1392
rect 1734 1387 1740 1388
rect 1902 1392 1908 1393
rect 1902 1388 1903 1392
rect 1907 1388 1908 1392
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2146 1395 2147 1399
rect 2151 1395 2152 1399
rect 2146 1394 2152 1395
rect 2346 1399 2352 1400
rect 2346 1395 2347 1399
rect 2351 1395 2352 1399
rect 2346 1394 2352 1395
rect 2570 1399 2576 1400
rect 2570 1395 2571 1399
rect 2575 1395 2576 1399
rect 2570 1394 2576 1395
rect 2658 1399 2664 1400
rect 2658 1395 2659 1399
rect 2663 1398 2664 1399
rect 2986 1399 2992 1400
rect 2663 1396 2753 1398
rect 2663 1395 2664 1396
rect 2658 1394 2664 1395
rect 2986 1395 2987 1399
rect 2991 1395 2992 1399
rect 2986 1394 2992 1395
rect 3170 1399 3176 1400
rect 3170 1395 3171 1399
rect 3175 1395 3176 1399
rect 3170 1394 3176 1395
rect 3198 1399 3204 1400
rect 3198 1395 3199 1399
rect 3203 1398 3204 1399
rect 3354 1399 3360 1400
rect 3203 1396 3313 1398
rect 3203 1395 3204 1396
rect 3198 1394 3204 1395
rect 3354 1395 3355 1399
rect 3359 1398 3360 1399
rect 3506 1399 3507 1403
rect 3511 1402 3512 1403
rect 3606 1403 3607 1407
rect 3611 1403 3612 1407
rect 3606 1402 3612 1403
rect 3782 1407 3788 1408
rect 3782 1403 3783 1407
rect 3787 1403 3788 1407
rect 3942 1404 3943 1408
rect 3947 1404 3948 1408
rect 3942 1403 3948 1404
rect 3782 1402 3788 1403
rect 3511 1400 3526 1402
rect 3511 1399 3512 1400
rect 3506 1398 3512 1399
rect 3524 1398 3526 1400
rect 3359 1396 3481 1398
rect 3524 1396 3649 1398
rect 3359 1395 3360 1396
rect 3354 1394 3360 1395
rect 3858 1395 3864 1396
rect 2006 1390 2012 1391
rect 2046 1391 2052 1392
rect 1902 1387 1908 1388
rect 2046 1387 2047 1391
rect 2051 1387 2052 1391
rect 3858 1391 3859 1395
rect 3863 1391 3864 1395
rect 3858 1390 3864 1391
rect 3942 1391 3948 1392
rect 2046 1386 2052 1387
rect 2070 1388 2076 1389
rect 2070 1384 2071 1388
rect 2075 1384 2076 1388
rect 2070 1383 2076 1384
rect 2270 1388 2276 1389
rect 2270 1384 2271 1388
rect 2275 1384 2276 1388
rect 2270 1383 2276 1384
rect 2494 1388 2500 1389
rect 2494 1384 2495 1388
rect 2499 1384 2500 1388
rect 2494 1383 2500 1384
rect 2710 1388 2716 1389
rect 2710 1384 2711 1388
rect 2715 1384 2716 1388
rect 2710 1383 2716 1384
rect 2910 1388 2916 1389
rect 2910 1384 2911 1388
rect 2915 1384 2916 1388
rect 2910 1383 2916 1384
rect 3094 1388 3100 1389
rect 3094 1384 3095 1388
rect 3099 1384 3100 1388
rect 3094 1383 3100 1384
rect 3270 1388 3276 1389
rect 3270 1384 3271 1388
rect 3275 1384 3276 1388
rect 3270 1383 3276 1384
rect 3438 1388 3444 1389
rect 3438 1384 3439 1388
rect 3443 1384 3444 1388
rect 3438 1383 3444 1384
rect 3606 1388 3612 1389
rect 3606 1384 3607 1388
rect 3611 1384 3612 1388
rect 3606 1383 3612 1384
rect 3782 1388 3788 1389
rect 3782 1384 3783 1388
rect 3787 1384 3788 1388
rect 3942 1387 3943 1391
rect 3947 1387 3948 1391
rect 3942 1386 3948 1387
rect 3782 1383 3788 1384
rect 158 1328 164 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 158 1324 159 1328
rect 163 1324 164 1328
rect 158 1323 164 1324
rect 310 1328 316 1329
rect 310 1324 311 1328
rect 315 1324 316 1328
rect 310 1323 316 1324
rect 478 1328 484 1329
rect 478 1324 479 1328
rect 483 1324 484 1328
rect 478 1323 484 1324
rect 662 1328 668 1329
rect 662 1324 663 1328
rect 667 1324 668 1328
rect 662 1323 668 1324
rect 854 1328 860 1329
rect 854 1324 855 1328
rect 859 1324 860 1328
rect 854 1323 860 1324
rect 1046 1328 1052 1329
rect 1046 1324 1047 1328
rect 1051 1324 1052 1328
rect 1046 1323 1052 1324
rect 1246 1328 1252 1329
rect 1246 1324 1247 1328
rect 1251 1324 1252 1328
rect 1246 1323 1252 1324
rect 1446 1328 1452 1329
rect 1446 1324 1447 1328
rect 1451 1324 1452 1328
rect 1446 1323 1452 1324
rect 1654 1328 1660 1329
rect 1654 1324 1655 1328
rect 1659 1324 1660 1328
rect 1654 1323 1660 1324
rect 1862 1328 1868 1329
rect 1862 1324 1863 1328
rect 1867 1324 1868 1328
rect 2070 1328 2076 1329
rect 1862 1323 1868 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2046 1325 2052 1326
rect 2046 1321 2047 1325
rect 2051 1321 2052 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2206 1328 2212 1329
rect 2206 1324 2207 1328
rect 2211 1324 2212 1328
rect 2206 1323 2212 1324
rect 2382 1328 2388 1329
rect 2382 1324 2383 1328
rect 2387 1324 2388 1328
rect 2382 1323 2388 1324
rect 2566 1328 2572 1329
rect 2566 1324 2567 1328
rect 2571 1324 2572 1328
rect 2566 1323 2572 1324
rect 2750 1328 2756 1329
rect 2750 1324 2751 1328
rect 2755 1324 2756 1328
rect 2750 1323 2756 1324
rect 2934 1328 2940 1329
rect 2934 1324 2935 1328
rect 2939 1324 2940 1328
rect 2934 1323 2940 1324
rect 3110 1328 3116 1329
rect 3110 1324 3111 1328
rect 3115 1324 3116 1328
rect 3110 1323 3116 1324
rect 3278 1328 3284 1329
rect 3278 1324 3279 1328
rect 3283 1324 3284 1328
rect 3278 1323 3284 1324
rect 3446 1328 3452 1329
rect 3446 1324 3447 1328
rect 3451 1324 3452 1328
rect 3446 1323 3452 1324
rect 3622 1328 3628 1329
rect 3622 1324 3623 1328
rect 3627 1324 3628 1328
rect 3622 1323 3628 1324
rect 3942 1325 3948 1326
rect 2046 1320 2052 1321
rect 3942 1321 3943 1325
rect 3947 1321 3948 1325
rect 3942 1320 3948 1321
rect 262 1319 268 1320
rect 262 1318 263 1319
rect 237 1316 263 1318
rect 262 1315 263 1316
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 386 1319 392 1320
rect 386 1315 387 1319
rect 391 1315 392 1319
rect 578 1319 584 1320
rect 578 1318 579 1319
rect 557 1316 579 1318
rect 386 1314 392 1315
rect 578 1315 579 1316
rect 583 1315 584 1319
rect 578 1314 584 1315
rect 738 1319 744 1320
rect 738 1315 739 1319
rect 743 1315 744 1319
rect 738 1314 744 1315
rect 746 1319 752 1320
rect 746 1315 747 1319
rect 751 1318 752 1319
rect 1122 1319 1128 1320
rect 751 1316 897 1318
rect 751 1315 752 1316
rect 746 1314 752 1315
rect 1122 1315 1123 1319
rect 1127 1315 1128 1319
rect 1122 1314 1128 1315
rect 1322 1319 1328 1320
rect 1322 1315 1323 1319
rect 1327 1315 1328 1319
rect 1322 1314 1328 1315
rect 1522 1319 1528 1320
rect 1522 1315 1523 1319
rect 1527 1315 1528 1319
rect 1742 1319 1748 1320
rect 1742 1318 1743 1319
rect 1733 1316 1743 1318
rect 1522 1314 1528 1315
rect 1742 1315 1743 1316
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 1799 1319 1805 1320
rect 1799 1315 1800 1319
rect 1804 1318 1805 1319
rect 2146 1319 2152 1320
rect 1804 1316 1905 1318
rect 1804 1315 1805 1316
rect 1799 1314 1805 1315
rect 2146 1315 2147 1319
rect 2151 1315 2152 1319
rect 2146 1314 2152 1315
rect 2282 1319 2288 1320
rect 2282 1315 2283 1319
rect 2287 1315 2288 1319
rect 2282 1314 2288 1315
rect 2458 1319 2464 1320
rect 2458 1315 2459 1319
rect 2463 1315 2464 1319
rect 2458 1314 2464 1315
rect 2642 1319 2648 1320
rect 2642 1315 2643 1319
rect 2647 1315 2648 1319
rect 2642 1314 2648 1315
rect 2718 1319 2724 1320
rect 2718 1315 2719 1319
rect 2723 1318 2724 1319
rect 3010 1319 3016 1320
rect 2723 1316 2793 1318
rect 2723 1315 2724 1316
rect 2718 1314 2724 1315
rect 3010 1315 3011 1319
rect 3015 1315 3016 1319
rect 3010 1314 3016 1315
rect 3186 1319 3192 1320
rect 3186 1315 3187 1319
rect 3191 1315 3192 1319
rect 3186 1314 3192 1315
rect 3354 1319 3360 1320
rect 3354 1315 3355 1319
rect 3359 1315 3360 1319
rect 3354 1314 3360 1315
rect 3522 1319 3528 1320
rect 3522 1315 3523 1319
rect 3527 1315 3528 1319
rect 3522 1314 3528 1315
rect 3567 1319 3573 1320
rect 3567 1315 3568 1319
rect 3572 1318 3573 1319
rect 3572 1316 3665 1318
rect 3572 1315 3573 1316
rect 3567 1314 3573 1315
rect 158 1309 164 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 158 1305 159 1309
rect 163 1305 164 1309
rect 158 1304 164 1305
rect 310 1309 316 1310
rect 310 1305 311 1309
rect 315 1305 316 1309
rect 310 1304 316 1305
rect 478 1309 484 1310
rect 478 1305 479 1309
rect 483 1305 484 1309
rect 478 1304 484 1305
rect 662 1309 668 1310
rect 662 1305 663 1309
rect 667 1305 668 1309
rect 662 1304 668 1305
rect 854 1309 860 1310
rect 854 1305 855 1309
rect 859 1305 860 1309
rect 854 1304 860 1305
rect 1046 1309 1052 1310
rect 1046 1305 1047 1309
rect 1051 1305 1052 1309
rect 1046 1304 1052 1305
rect 1246 1309 1252 1310
rect 1246 1305 1247 1309
rect 1251 1305 1252 1309
rect 1246 1304 1252 1305
rect 1446 1309 1452 1310
rect 1446 1305 1447 1309
rect 1451 1305 1452 1309
rect 1446 1304 1452 1305
rect 1654 1309 1660 1310
rect 1654 1305 1655 1309
rect 1659 1305 1660 1309
rect 1654 1304 1660 1305
rect 1862 1309 1868 1310
rect 2070 1309 2076 1310
rect 1862 1305 1863 1309
rect 1867 1305 1868 1309
rect 1862 1304 1868 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 110 1303 116 1304
rect 2006 1303 2012 1304
rect 2046 1308 2052 1309
rect 2046 1304 2047 1308
rect 2051 1304 2052 1308
rect 2070 1305 2071 1309
rect 2075 1305 2076 1309
rect 2070 1304 2076 1305
rect 2206 1309 2212 1310
rect 2206 1305 2207 1309
rect 2211 1305 2212 1309
rect 2206 1304 2212 1305
rect 2382 1309 2388 1310
rect 2382 1305 2383 1309
rect 2387 1305 2388 1309
rect 2382 1304 2388 1305
rect 2566 1309 2572 1310
rect 2566 1305 2567 1309
rect 2571 1305 2572 1309
rect 2566 1304 2572 1305
rect 2750 1309 2756 1310
rect 2750 1305 2751 1309
rect 2755 1305 2756 1309
rect 2750 1304 2756 1305
rect 2934 1309 2940 1310
rect 2934 1305 2935 1309
rect 2939 1305 2940 1309
rect 2934 1304 2940 1305
rect 3110 1309 3116 1310
rect 3110 1305 3111 1309
rect 3115 1305 3116 1309
rect 3110 1304 3116 1305
rect 3278 1309 3284 1310
rect 3278 1305 3279 1309
rect 3283 1305 3284 1309
rect 3278 1304 3284 1305
rect 3446 1309 3452 1310
rect 3446 1305 3447 1309
rect 3451 1305 3452 1309
rect 3446 1304 3452 1305
rect 3622 1309 3628 1310
rect 3622 1305 3623 1309
rect 3627 1305 3628 1309
rect 3622 1304 3628 1305
rect 3942 1308 3948 1309
rect 3942 1304 3943 1308
rect 3947 1304 3948 1308
rect 2046 1303 2052 1304
rect 3942 1303 3948 1304
rect 746 1299 752 1300
rect 746 1298 747 1299
rect 319 1296 747 1298
rect 319 1294 321 1296
rect 746 1295 747 1296
rect 751 1295 752 1299
rect 2658 1299 2664 1300
rect 2658 1298 2659 1299
rect 746 1294 752 1295
rect 2140 1296 2659 1298
rect 256 1292 321 1294
rect 195 1291 201 1292
rect 195 1287 196 1291
rect 200 1290 201 1291
rect 256 1290 258 1292
rect 200 1288 258 1290
rect 386 1291 392 1292
rect 200 1287 201 1288
rect 195 1286 201 1287
rect 262 1287 268 1288
rect 262 1283 263 1287
rect 267 1286 268 1287
rect 347 1287 353 1288
rect 347 1286 348 1287
rect 267 1284 348 1286
rect 267 1283 268 1284
rect 262 1282 268 1283
rect 347 1283 348 1284
rect 352 1283 353 1287
rect 386 1287 387 1291
rect 391 1290 392 1291
rect 515 1291 521 1292
rect 515 1290 516 1291
rect 391 1288 516 1290
rect 391 1287 392 1288
rect 386 1286 392 1287
rect 515 1287 516 1288
rect 520 1287 521 1291
rect 738 1291 744 1292
rect 515 1286 521 1287
rect 618 1287 624 1288
rect 347 1282 353 1283
rect 618 1283 619 1287
rect 623 1286 624 1287
rect 699 1287 705 1288
rect 699 1286 700 1287
rect 623 1284 700 1286
rect 623 1283 624 1284
rect 618 1282 624 1283
rect 699 1283 700 1284
rect 704 1283 705 1287
rect 738 1287 739 1291
rect 743 1290 744 1291
rect 891 1291 897 1292
rect 891 1290 892 1291
rect 743 1288 892 1290
rect 743 1287 744 1288
rect 738 1286 744 1287
rect 891 1287 892 1288
rect 896 1287 897 1291
rect 891 1286 897 1287
rect 1082 1291 1089 1292
rect 1082 1287 1083 1291
rect 1088 1287 1089 1291
rect 1082 1286 1089 1287
rect 1122 1291 1128 1292
rect 1122 1287 1123 1291
rect 1127 1290 1128 1291
rect 1283 1291 1289 1292
rect 1283 1290 1284 1291
rect 1127 1288 1284 1290
rect 1127 1287 1128 1288
rect 1122 1286 1128 1287
rect 1283 1287 1284 1288
rect 1288 1287 1289 1291
rect 1283 1286 1289 1287
rect 1322 1291 1328 1292
rect 1322 1287 1323 1291
rect 1327 1290 1328 1291
rect 1483 1291 1489 1292
rect 1483 1290 1484 1291
rect 1327 1288 1484 1290
rect 1327 1287 1328 1288
rect 1322 1286 1328 1287
rect 1483 1287 1484 1288
rect 1488 1287 1489 1291
rect 1483 1286 1489 1287
rect 1691 1291 1697 1292
rect 1691 1287 1692 1291
rect 1696 1290 1697 1291
rect 1799 1291 1805 1292
rect 1799 1290 1800 1291
rect 1696 1288 1800 1290
rect 1696 1287 1697 1288
rect 1691 1286 1697 1287
rect 1799 1287 1800 1288
rect 1804 1287 1805 1291
rect 2107 1291 2113 1292
rect 1799 1286 1805 1287
rect 1887 1287 1893 1288
rect 699 1282 705 1283
rect 1887 1283 1888 1287
rect 1892 1286 1893 1287
rect 1899 1287 1905 1288
rect 1899 1286 1900 1287
rect 1892 1284 1900 1286
rect 1892 1283 1893 1284
rect 1887 1282 1893 1283
rect 1899 1283 1900 1284
rect 1904 1283 1905 1287
rect 2107 1287 2108 1291
rect 2112 1290 2113 1291
rect 2140 1290 2142 1296
rect 2658 1295 2659 1296
rect 2663 1295 2664 1299
rect 3198 1299 3204 1300
rect 3198 1298 3199 1299
rect 2658 1294 2664 1295
rect 3004 1296 3199 1298
rect 2112 1288 2142 1290
rect 2146 1291 2152 1292
rect 2112 1287 2113 1288
rect 2107 1286 2113 1287
rect 2146 1287 2147 1291
rect 2151 1290 2152 1291
rect 2243 1291 2249 1292
rect 2243 1290 2244 1291
rect 2151 1288 2244 1290
rect 2151 1287 2152 1288
rect 2146 1286 2152 1287
rect 2243 1287 2244 1288
rect 2248 1287 2249 1291
rect 2243 1286 2249 1287
rect 2282 1291 2288 1292
rect 2282 1287 2283 1291
rect 2287 1290 2288 1291
rect 2419 1291 2425 1292
rect 2419 1290 2420 1291
rect 2287 1288 2420 1290
rect 2287 1287 2288 1288
rect 2282 1286 2288 1287
rect 2419 1287 2420 1288
rect 2424 1287 2425 1291
rect 2419 1286 2425 1287
rect 2458 1291 2464 1292
rect 2458 1287 2459 1291
rect 2463 1290 2464 1291
rect 2603 1291 2609 1292
rect 2603 1290 2604 1291
rect 2463 1288 2604 1290
rect 2463 1287 2464 1288
rect 2458 1286 2464 1287
rect 2603 1287 2604 1288
rect 2608 1287 2609 1291
rect 2603 1286 2609 1287
rect 2642 1291 2648 1292
rect 2642 1287 2643 1291
rect 2647 1290 2648 1291
rect 2787 1291 2793 1292
rect 2787 1290 2788 1291
rect 2647 1288 2788 1290
rect 2647 1287 2648 1288
rect 2642 1286 2648 1287
rect 2787 1287 2788 1288
rect 2792 1287 2793 1291
rect 2787 1286 2793 1287
rect 2971 1291 2977 1292
rect 2971 1287 2972 1291
rect 2976 1290 2977 1291
rect 3004 1290 3006 1296
rect 3198 1295 3199 1296
rect 3203 1295 3204 1299
rect 3198 1294 3204 1295
rect 2976 1288 3006 1290
rect 3010 1291 3016 1292
rect 2976 1287 2977 1288
rect 2971 1286 2977 1287
rect 3010 1287 3011 1291
rect 3015 1290 3016 1291
rect 3147 1291 3153 1292
rect 3147 1290 3148 1291
rect 3015 1288 3148 1290
rect 3015 1287 3016 1288
rect 3010 1286 3016 1287
rect 3147 1287 3148 1288
rect 3152 1287 3153 1291
rect 3147 1286 3153 1287
rect 3186 1291 3192 1292
rect 3186 1287 3187 1291
rect 3191 1290 3192 1291
rect 3315 1291 3321 1292
rect 3315 1290 3316 1291
rect 3191 1288 3316 1290
rect 3191 1287 3192 1288
rect 3186 1286 3192 1287
rect 3315 1287 3316 1288
rect 3320 1287 3321 1291
rect 3315 1286 3321 1287
rect 3483 1291 3489 1292
rect 3483 1287 3484 1291
rect 3488 1290 3489 1291
rect 3567 1291 3573 1292
rect 3567 1290 3568 1291
rect 3488 1288 3568 1290
rect 3488 1287 3489 1288
rect 3483 1286 3489 1287
rect 3567 1287 3568 1288
rect 3572 1287 3573 1291
rect 3567 1286 3573 1287
rect 3659 1287 3665 1288
rect 1899 1282 1905 1283
rect 2718 1283 2724 1284
rect 2718 1282 2719 1283
rect 2188 1280 2719 1282
rect 2188 1278 2190 1280
rect 2718 1279 2719 1280
rect 2723 1279 2724 1283
rect 2718 1278 2724 1279
rect 2982 1283 2988 1284
rect 2982 1279 2983 1283
rect 2987 1282 2988 1283
rect 3231 1283 3237 1284
rect 3231 1282 3232 1283
rect 2987 1280 3232 1282
rect 2987 1279 2988 1280
rect 2982 1278 2988 1279
rect 3231 1279 3232 1280
rect 3236 1279 3237 1283
rect 3659 1283 3660 1287
rect 3664 1286 3665 1287
rect 3690 1287 3696 1288
rect 3690 1286 3691 1287
rect 3664 1284 3691 1286
rect 3664 1283 3665 1284
rect 3659 1282 3665 1283
rect 3690 1283 3691 1284
rect 3695 1283 3696 1287
rect 3690 1282 3696 1283
rect 3231 1278 3237 1279
rect 2187 1277 2193 1278
rect 2187 1273 2188 1277
rect 2192 1273 2193 1277
rect 2187 1272 2193 1273
rect 2226 1275 2232 1276
rect 443 1271 452 1272
rect 443 1267 444 1271
rect 451 1267 452 1271
rect 443 1266 452 1267
rect 511 1271 517 1272
rect 511 1267 512 1271
rect 516 1270 517 1271
rect 579 1271 585 1272
rect 579 1270 580 1271
rect 516 1268 580 1270
rect 516 1267 517 1268
rect 511 1266 517 1267
rect 579 1267 580 1268
rect 584 1267 585 1271
rect 579 1266 585 1267
rect 674 1271 680 1272
rect 674 1267 675 1271
rect 679 1270 680 1271
rect 731 1271 737 1272
rect 731 1270 732 1271
rect 679 1268 732 1270
rect 679 1267 680 1268
rect 674 1266 680 1267
rect 731 1267 732 1268
rect 736 1267 737 1271
rect 731 1266 737 1267
rect 770 1271 776 1272
rect 770 1267 771 1271
rect 775 1270 776 1271
rect 891 1271 897 1272
rect 891 1270 892 1271
rect 775 1268 892 1270
rect 775 1267 776 1268
rect 770 1266 776 1267
rect 891 1267 892 1268
rect 896 1267 897 1271
rect 891 1266 897 1267
rect 930 1271 936 1272
rect 930 1267 931 1271
rect 935 1270 936 1271
rect 1059 1271 1065 1272
rect 1059 1270 1060 1271
rect 935 1268 1060 1270
rect 935 1267 936 1268
rect 930 1266 936 1267
rect 1059 1267 1060 1268
rect 1064 1267 1065 1271
rect 1059 1266 1065 1267
rect 1227 1271 1233 1272
rect 1227 1267 1228 1271
rect 1232 1270 1233 1271
rect 1274 1271 1280 1272
rect 1274 1270 1275 1271
rect 1232 1268 1275 1270
rect 1232 1267 1233 1268
rect 1227 1266 1233 1267
rect 1274 1267 1275 1268
rect 1279 1267 1280 1271
rect 1274 1266 1280 1267
rect 1403 1271 1409 1272
rect 1403 1267 1404 1271
rect 1408 1270 1409 1271
rect 1454 1271 1460 1272
rect 1454 1270 1455 1271
rect 1408 1268 1455 1270
rect 1408 1267 1409 1268
rect 1403 1266 1409 1267
rect 1454 1267 1455 1268
rect 1459 1267 1460 1271
rect 1454 1266 1460 1267
rect 1522 1271 1528 1272
rect 1522 1267 1523 1271
rect 1527 1270 1528 1271
rect 1579 1271 1585 1272
rect 1579 1270 1580 1271
rect 1527 1268 1580 1270
rect 1527 1267 1528 1268
rect 1522 1266 1528 1267
rect 1579 1267 1580 1268
rect 1584 1267 1585 1271
rect 1579 1266 1585 1267
rect 1755 1271 1761 1272
rect 1755 1267 1756 1271
rect 1760 1270 1761 1271
rect 1770 1271 1776 1272
rect 1770 1270 1771 1271
rect 1760 1268 1771 1270
rect 1760 1267 1761 1268
rect 1755 1266 1761 1267
rect 1770 1267 1771 1268
rect 1775 1267 1776 1271
rect 1770 1266 1776 1267
rect 1794 1271 1800 1272
rect 1794 1267 1795 1271
rect 1799 1270 1800 1271
rect 1931 1271 1937 1272
rect 1931 1270 1932 1271
rect 1799 1268 1932 1270
rect 1799 1267 1800 1268
rect 1794 1266 1800 1267
rect 1931 1267 1932 1268
rect 1936 1267 1937 1271
rect 2226 1271 2227 1275
rect 2231 1274 2232 1275
rect 2323 1275 2329 1276
rect 2323 1274 2324 1275
rect 2231 1272 2324 1274
rect 2231 1271 2232 1272
rect 2226 1270 2232 1271
rect 2323 1271 2324 1272
rect 2328 1271 2329 1275
rect 2323 1270 2329 1271
rect 2362 1275 2368 1276
rect 2362 1271 2363 1275
rect 2367 1274 2368 1275
rect 2467 1275 2473 1276
rect 2467 1274 2468 1275
rect 2367 1272 2468 1274
rect 2367 1271 2368 1272
rect 2362 1270 2368 1271
rect 2467 1271 2468 1272
rect 2472 1271 2473 1275
rect 2467 1270 2473 1271
rect 2506 1275 2512 1276
rect 2506 1271 2507 1275
rect 2511 1274 2512 1275
rect 2619 1275 2625 1276
rect 2619 1274 2620 1275
rect 2511 1272 2620 1274
rect 2511 1271 2512 1272
rect 2506 1270 2512 1271
rect 2619 1271 2620 1272
rect 2624 1271 2625 1275
rect 2619 1270 2625 1271
rect 2658 1275 2664 1276
rect 2658 1271 2659 1275
rect 2663 1274 2664 1275
rect 2779 1275 2785 1276
rect 2779 1274 2780 1275
rect 2663 1272 2780 1274
rect 2663 1271 2664 1272
rect 2658 1270 2664 1271
rect 2779 1271 2780 1272
rect 2784 1271 2785 1275
rect 2779 1270 2785 1271
rect 2939 1275 2945 1276
rect 2939 1271 2940 1275
rect 2944 1274 2945 1275
rect 2970 1275 2976 1276
rect 2970 1274 2971 1275
rect 2944 1272 2971 1274
rect 2944 1271 2945 1272
rect 2939 1270 2945 1271
rect 2970 1271 2971 1272
rect 2975 1271 2976 1275
rect 2970 1270 2976 1271
rect 2978 1275 2984 1276
rect 2978 1271 2979 1275
rect 2983 1274 2984 1275
rect 3107 1275 3113 1276
rect 3107 1274 3108 1275
rect 2983 1272 3108 1274
rect 2983 1271 2984 1272
rect 2978 1270 2984 1271
rect 3107 1271 3108 1272
rect 3112 1271 3113 1275
rect 3107 1270 3113 1271
rect 3283 1275 3289 1276
rect 3283 1271 3284 1275
rect 3288 1274 3289 1275
rect 3330 1275 3336 1276
rect 3330 1274 3331 1275
rect 3288 1272 3331 1274
rect 3288 1271 3289 1272
rect 3283 1270 3289 1271
rect 3330 1271 3331 1272
rect 3335 1271 3336 1275
rect 3330 1270 3336 1271
rect 3354 1275 3360 1276
rect 3354 1271 3355 1275
rect 3359 1274 3360 1275
rect 3467 1275 3473 1276
rect 3467 1274 3468 1275
rect 3359 1272 3468 1274
rect 3359 1271 3360 1272
rect 3354 1270 3360 1271
rect 3467 1271 3468 1272
rect 3472 1271 3473 1275
rect 3467 1270 3473 1271
rect 3651 1275 3657 1276
rect 3651 1271 3652 1275
rect 3656 1274 3657 1275
rect 3698 1275 3704 1276
rect 3698 1274 3699 1275
rect 3656 1272 3699 1274
rect 3656 1271 3657 1272
rect 3651 1270 3657 1271
rect 3698 1271 3699 1272
rect 3703 1271 3704 1275
rect 3698 1270 3704 1271
rect 3843 1275 3849 1276
rect 3843 1271 3844 1275
rect 3848 1274 3849 1275
rect 3858 1275 3864 1276
rect 3858 1274 3859 1275
rect 3848 1272 3859 1274
rect 3848 1271 3849 1272
rect 3843 1270 3849 1271
rect 3858 1271 3859 1272
rect 3863 1271 3864 1275
rect 3858 1270 3864 1271
rect 1931 1266 1937 1267
rect 2046 1256 2052 1257
rect 3942 1256 3948 1257
rect 110 1252 116 1253
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 406 1251 412 1252
rect 406 1247 407 1251
rect 411 1247 412 1251
rect 406 1246 412 1247
rect 542 1251 548 1252
rect 542 1247 543 1251
rect 547 1247 548 1251
rect 542 1246 548 1247
rect 694 1251 700 1252
rect 694 1247 695 1251
rect 699 1247 700 1251
rect 694 1246 700 1247
rect 854 1251 860 1252
rect 854 1247 855 1251
rect 859 1247 860 1251
rect 854 1246 860 1247
rect 1022 1251 1028 1252
rect 1022 1247 1023 1251
rect 1027 1247 1028 1251
rect 1022 1246 1028 1247
rect 1190 1251 1196 1252
rect 1190 1247 1191 1251
rect 1195 1247 1196 1251
rect 1190 1246 1196 1247
rect 1366 1251 1372 1252
rect 1366 1247 1367 1251
rect 1371 1247 1372 1251
rect 1366 1246 1372 1247
rect 1542 1251 1548 1252
rect 1542 1247 1543 1251
rect 1547 1247 1548 1251
rect 1542 1246 1548 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 1718 1246 1724 1247
rect 1894 1251 1900 1252
rect 1894 1247 1895 1251
rect 1899 1247 1900 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2046 1252 2047 1256
rect 2051 1252 2052 1256
rect 2046 1251 2052 1252
rect 2150 1255 2156 1256
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2286 1255 2292 1256
rect 2286 1251 2287 1255
rect 2291 1251 2292 1255
rect 2286 1250 2292 1251
rect 2430 1255 2436 1256
rect 2430 1251 2431 1255
rect 2435 1251 2436 1255
rect 2430 1250 2436 1251
rect 2582 1255 2588 1256
rect 2582 1251 2583 1255
rect 2587 1251 2588 1255
rect 2582 1250 2588 1251
rect 2742 1255 2748 1256
rect 2742 1251 2743 1255
rect 2747 1251 2748 1255
rect 2742 1250 2748 1251
rect 2902 1255 2908 1256
rect 2902 1251 2903 1255
rect 2907 1251 2908 1255
rect 2902 1250 2908 1251
rect 3070 1255 3076 1256
rect 3070 1251 3071 1255
rect 3075 1251 3076 1255
rect 3070 1250 3076 1251
rect 3246 1255 3252 1256
rect 3246 1251 3247 1255
rect 3251 1251 3252 1255
rect 3246 1250 3252 1251
rect 3430 1255 3436 1256
rect 3430 1251 3431 1255
rect 3435 1251 3436 1255
rect 3430 1250 3436 1251
rect 3614 1255 3620 1256
rect 3614 1251 3615 1255
rect 3619 1251 3620 1255
rect 3614 1250 3620 1251
rect 3806 1255 3812 1256
rect 3806 1251 3807 1255
rect 3811 1251 3812 1255
rect 3942 1252 3943 1256
rect 3947 1252 3948 1256
rect 3942 1251 3948 1252
rect 3806 1250 3812 1251
rect 2006 1247 2012 1248
rect 2226 1247 2232 1248
rect 1894 1246 1900 1247
rect 511 1243 517 1244
rect 511 1242 512 1243
rect 485 1240 512 1242
rect 511 1239 512 1240
rect 516 1239 517 1243
rect 511 1238 517 1239
rect 618 1243 624 1244
rect 618 1239 619 1243
rect 623 1239 624 1243
rect 618 1238 624 1239
rect 770 1243 776 1244
rect 770 1239 771 1243
rect 775 1239 776 1243
rect 770 1238 776 1239
rect 930 1243 936 1244
rect 930 1239 931 1243
rect 935 1239 936 1243
rect 930 1238 936 1239
rect 978 1243 984 1244
rect 978 1239 979 1243
rect 983 1242 984 1243
rect 1274 1243 1280 1244
rect 983 1240 1065 1242
rect 983 1239 984 1240
rect 978 1238 984 1239
rect 1266 1239 1272 1240
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1266 1235 1267 1239
rect 1271 1235 1272 1239
rect 1274 1239 1275 1243
rect 1279 1242 1280 1243
rect 1454 1243 1460 1244
rect 1279 1240 1409 1242
rect 1279 1239 1280 1240
rect 1274 1238 1280 1239
rect 1454 1239 1455 1243
rect 1459 1242 1460 1243
rect 1794 1243 1800 1244
rect 1459 1240 1585 1242
rect 1459 1239 1460 1240
rect 1454 1238 1460 1239
rect 1794 1239 1795 1243
rect 1799 1239 1800 1243
rect 1794 1238 1800 1239
rect 1887 1243 1893 1244
rect 1887 1239 1888 1243
rect 1892 1242 1893 1243
rect 2226 1243 2227 1247
rect 2231 1243 2232 1247
rect 2226 1242 2232 1243
rect 2362 1247 2368 1248
rect 2362 1243 2363 1247
rect 2367 1243 2368 1247
rect 2362 1242 2368 1243
rect 2506 1247 2512 1248
rect 2506 1243 2507 1247
rect 2511 1243 2512 1247
rect 2506 1242 2512 1243
rect 2658 1247 2664 1248
rect 2658 1243 2659 1247
rect 2663 1243 2664 1247
rect 2658 1242 2664 1243
rect 2666 1247 2672 1248
rect 2666 1243 2667 1247
rect 2671 1246 2672 1247
rect 2978 1247 2984 1248
rect 2671 1244 2785 1246
rect 2671 1243 2672 1244
rect 2666 1242 2672 1243
rect 2978 1243 2979 1247
rect 2983 1243 2984 1247
rect 3231 1247 3237 1248
rect 2978 1242 2984 1243
rect 3223 1243 3229 1244
rect 3223 1242 3224 1243
rect 1892 1240 1937 1242
rect 3149 1240 3224 1242
rect 1892 1239 1893 1240
rect 1887 1238 1893 1239
rect 2046 1239 2052 1240
rect 1266 1234 1272 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 406 1232 412 1233
rect 406 1228 407 1232
rect 411 1228 412 1232
rect 406 1227 412 1228
rect 542 1232 548 1233
rect 542 1228 543 1232
rect 547 1228 548 1232
rect 542 1227 548 1228
rect 694 1232 700 1233
rect 694 1228 695 1232
rect 699 1228 700 1232
rect 694 1227 700 1228
rect 854 1232 860 1233
rect 854 1228 855 1232
rect 859 1228 860 1232
rect 854 1227 860 1228
rect 1022 1232 1028 1233
rect 1022 1228 1023 1232
rect 1027 1228 1028 1232
rect 1022 1227 1028 1228
rect 1190 1232 1196 1233
rect 1190 1228 1191 1232
rect 1195 1228 1196 1232
rect 1190 1227 1196 1228
rect 1366 1232 1372 1233
rect 1366 1228 1367 1232
rect 1371 1228 1372 1232
rect 1366 1227 1372 1228
rect 1542 1232 1548 1233
rect 1542 1228 1543 1232
rect 1547 1228 1548 1232
rect 1542 1227 1548 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 1718 1227 1724 1228
rect 1894 1232 1900 1233
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2046 1235 2047 1239
rect 2051 1235 2052 1239
rect 3223 1239 3224 1240
rect 3228 1239 3229 1243
rect 3231 1243 3232 1247
rect 3236 1246 3237 1247
rect 3330 1247 3336 1248
rect 3236 1244 3289 1246
rect 3236 1243 3237 1244
rect 3231 1242 3237 1243
rect 3330 1243 3331 1247
rect 3335 1246 3336 1247
rect 3690 1247 3696 1248
rect 3335 1244 3473 1246
rect 3335 1243 3336 1244
rect 3330 1242 3336 1243
rect 3690 1243 3691 1247
rect 3695 1243 3696 1247
rect 3690 1242 3696 1243
rect 3882 1243 3888 1244
rect 3223 1238 3229 1239
rect 3882 1239 3883 1243
rect 3887 1239 3888 1243
rect 3882 1238 3888 1239
rect 3942 1239 3948 1240
rect 2046 1234 2052 1235
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2286 1236 2292 1237
rect 2286 1232 2287 1236
rect 2291 1232 2292 1236
rect 2286 1231 2292 1232
rect 2430 1236 2436 1237
rect 2430 1232 2431 1236
rect 2435 1232 2436 1236
rect 2430 1231 2436 1232
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 2582 1231 2588 1232
rect 2742 1236 2748 1237
rect 2742 1232 2743 1236
rect 2747 1232 2748 1236
rect 2742 1231 2748 1232
rect 2902 1236 2908 1237
rect 2902 1232 2903 1236
rect 2907 1232 2908 1236
rect 2902 1231 2908 1232
rect 3070 1236 3076 1237
rect 3070 1232 3071 1236
rect 3075 1232 3076 1236
rect 3070 1231 3076 1232
rect 3246 1236 3252 1237
rect 3246 1232 3247 1236
rect 3251 1232 3252 1236
rect 3246 1231 3252 1232
rect 3430 1236 3436 1237
rect 3430 1232 3431 1236
rect 3435 1232 3436 1236
rect 3430 1231 3436 1232
rect 3614 1236 3620 1237
rect 3614 1232 3615 1236
rect 3619 1232 3620 1236
rect 3614 1231 3620 1232
rect 3806 1236 3812 1237
rect 3806 1232 3807 1236
rect 3811 1232 3812 1236
rect 3942 1235 3943 1239
rect 3947 1235 3948 1239
rect 3942 1234 3948 1235
rect 3806 1231 3812 1232
rect 2006 1230 2012 1231
rect 1894 1227 1900 1228
rect 2350 1215 2356 1216
rect 2350 1211 2351 1215
rect 2355 1214 2356 1215
rect 2666 1215 2672 1216
rect 2666 1214 2667 1215
rect 2355 1212 2667 1214
rect 2355 1211 2356 1212
rect 2350 1210 2356 1211
rect 2666 1211 2667 1212
rect 2671 1211 2672 1215
rect 2666 1210 2672 1211
rect 2310 1176 2316 1177
rect 2046 1173 2052 1174
rect 422 1172 428 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 422 1168 423 1172
rect 427 1168 428 1172
rect 422 1167 428 1168
rect 590 1172 596 1173
rect 590 1168 591 1172
rect 595 1168 596 1172
rect 590 1167 596 1168
rect 758 1172 764 1173
rect 758 1168 759 1172
rect 763 1168 764 1172
rect 758 1167 764 1168
rect 926 1172 932 1173
rect 926 1168 927 1172
rect 931 1168 932 1172
rect 926 1167 932 1168
rect 1094 1172 1100 1173
rect 1094 1168 1095 1172
rect 1099 1168 1100 1172
rect 1094 1167 1100 1168
rect 1246 1172 1252 1173
rect 1246 1168 1247 1172
rect 1251 1168 1252 1172
rect 1246 1167 1252 1168
rect 1398 1172 1404 1173
rect 1398 1168 1399 1172
rect 1403 1168 1404 1172
rect 1398 1167 1404 1168
rect 1542 1172 1548 1173
rect 1542 1168 1543 1172
rect 1547 1168 1548 1172
rect 1542 1167 1548 1168
rect 1686 1172 1692 1173
rect 1686 1168 1687 1172
rect 1691 1168 1692 1172
rect 1686 1167 1692 1168
rect 1838 1172 1844 1173
rect 1838 1168 1839 1172
rect 1843 1168 1844 1172
rect 1838 1167 1844 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2046 1169 2047 1173
rect 2051 1169 2052 1173
rect 2310 1172 2311 1176
rect 2315 1172 2316 1176
rect 2310 1171 2316 1172
rect 2414 1176 2420 1177
rect 2414 1172 2415 1176
rect 2419 1172 2420 1176
rect 2414 1171 2420 1172
rect 2526 1176 2532 1177
rect 2526 1172 2527 1176
rect 2531 1172 2532 1176
rect 2526 1171 2532 1172
rect 2638 1176 2644 1177
rect 2638 1172 2639 1176
rect 2643 1172 2644 1176
rect 2638 1171 2644 1172
rect 2766 1176 2772 1177
rect 2766 1172 2767 1176
rect 2771 1172 2772 1176
rect 2766 1171 2772 1172
rect 2910 1176 2916 1177
rect 2910 1172 2911 1176
rect 2915 1172 2916 1176
rect 2910 1171 2916 1172
rect 3070 1176 3076 1177
rect 3070 1172 3071 1176
rect 3075 1172 3076 1176
rect 3070 1171 3076 1172
rect 3246 1176 3252 1177
rect 3246 1172 3247 1176
rect 3251 1172 3252 1176
rect 3246 1171 3252 1172
rect 3438 1176 3444 1177
rect 3438 1172 3439 1176
rect 3443 1172 3444 1176
rect 3438 1171 3444 1172
rect 3630 1176 3636 1177
rect 3630 1172 3631 1176
rect 3635 1172 3636 1176
rect 3630 1171 3636 1172
rect 3830 1176 3836 1177
rect 3830 1172 3831 1176
rect 3835 1172 3836 1176
rect 3830 1171 3836 1172
rect 3942 1173 3948 1174
rect 2046 1168 2052 1169
rect 3942 1169 3943 1173
rect 3947 1169 3948 1173
rect 3942 1168 3948 1169
rect 2006 1164 2012 1165
rect 2386 1167 2392 1168
rect 498 1163 504 1164
rect 498 1159 499 1163
rect 503 1159 504 1163
rect 674 1163 680 1164
rect 674 1162 675 1163
rect 669 1160 675 1162
rect 498 1158 504 1159
rect 674 1159 675 1160
rect 679 1159 680 1163
rect 674 1158 680 1159
rect 718 1163 724 1164
rect 718 1159 719 1163
rect 723 1162 724 1163
rect 878 1163 884 1164
rect 723 1160 801 1162
rect 723 1159 724 1160
rect 718 1158 724 1159
rect 878 1159 879 1163
rect 883 1162 884 1163
rect 1047 1163 1053 1164
rect 883 1160 969 1162
rect 883 1159 884 1160
rect 878 1158 884 1159
rect 1047 1159 1048 1163
rect 1052 1162 1053 1163
rect 1322 1163 1328 1164
rect 1052 1160 1137 1162
rect 1052 1159 1053 1160
rect 1047 1158 1053 1159
rect 1322 1159 1323 1163
rect 1327 1159 1328 1163
rect 1535 1163 1541 1164
rect 1535 1162 1536 1163
rect 1477 1160 1536 1162
rect 1322 1158 1328 1159
rect 1535 1159 1536 1160
rect 1540 1159 1541 1163
rect 1535 1158 1541 1159
rect 1618 1163 1624 1164
rect 1618 1159 1619 1163
rect 1623 1159 1624 1163
rect 1618 1158 1624 1159
rect 1762 1163 1768 1164
rect 1762 1159 1763 1163
rect 1767 1159 1768 1163
rect 1762 1158 1768 1159
rect 1770 1163 1776 1164
rect 1770 1159 1771 1163
rect 1775 1162 1776 1163
rect 2386 1163 2387 1167
rect 2391 1163 2392 1167
rect 2386 1162 2392 1163
rect 2490 1167 2496 1168
rect 2490 1163 2491 1167
rect 2495 1163 2496 1167
rect 2490 1162 2496 1163
rect 2602 1167 2608 1168
rect 2602 1163 2603 1167
rect 2607 1163 2608 1167
rect 2602 1162 2608 1163
rect 2714 1167 2720 1168
rect 2714 1163 2715 1167
rect 2719 1163 2720 1167
rect 2714 1162 2720 1163
rect 2722 1167 2728 1168
rect 2722 1163 2723 1167
rect 2727 1166 2728 1167
rect 2986 1167 2992 1168
rect 2727 1164 2809 1166
rect 2727 1163 2728 1164
rect 2722 1162 2728 1163
rect 2986 1163 2987 1167
rect 2991 1163 2992 1167
rect 2986 1162 2992 1163
rect 3138 1167 3144 1168
rect 3138 1163 3139 1167
rect 3143 1163 3144 1167
rect 3138 1162 3144 1163
rect 3322 1167 3328 1168
rect 3322 1163 3323 1167
rect 3327 1163 3328 1167
rect 3322 1162 3328 1163
rect 3378 1167 3384 1168
rect 3378 1163 3379 1167
rect 3383 1166 3384 1167
rect 3698 1167 3704 1168
rect 3383 1164 3481 1166
rect 3383 1163 3384 1164
rect 3378 1162 3384 1163
rect 3698 1163 3699 1167
rect 3703 1163 3704 1167
rect 3698 1162 3704 1163
rect 3898 1167 3904 1168
rect 3898 1163 3899 1167
rect 3903 1163 3904 1167
rect 3898 1162 3904 1163
rect 1775 1160 1881 1162
rect 1775 1159 1776 1160
rect 1770 1158 1776 1159
rect 2310 1157 2316 1158
rect 2046 1156 2052 1157
rect 422 1153 428 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 422 1149 423 1153
rect 427 1149 428 1153
rect 422 1148 428 1149
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 758 1153 764 1154
rect 758 1149 759 1153
rect 763 1149 764 1153
rect 758 1148 764 1149
rect 926 1153 932 1154
rect 926 1149 927 1153
rect 931 1149 932 1153
rect 926 1148 932 1149
rect 1094 1153 1100 1154
rect 1094 1149 1095 1153
rect 1099 1149 1100 1153
rect 1094 1148 1100 1149
rect 1246 1153 1252 1154
rect 1246 1149 1247 1153
rect 1251 1149 1252 1153
rect 1246 1148 1252 1149
rect 1398 1153 1404 1154
rect 1398 1149 1399 1153
rect 1403 1149 1404 1153
rect 1398 1148 1404 1149
rect 1542 1153 1548 1154
rect 1542 1149 1543 1153
rect 1547 1149 1548 1153
rect 1542 1148 1548 1149
rect 1686 1153 1692 1154
rect 1686 1149 1687 1153
rect 1691 1149 1692 1153
rect 1686 1148 1692 1149
rect 1838 1153 1844 1154
rect 1838 1149 1839 1153
rect 1843 1149 1844 1153
rect 1838 1148 1844 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2046 1152 2047 1156
rect 2051 1152 2052 1156
rect 2310 1153 2311 1157
rect 2315 1153 2316 1157
rect 2310 1152 2316 1153
rect 2414 1157 2420 1158
rect 2414 1153 2415 1157
rect 2419 1153 2420 1157
rect 2414 1152 2420 1153
rect 2526 1157 2532 1158
rect 2526 1153 2527 1157
rect 2531 1153 2532 1157
rect 2526 1152 2532 1153
rect 2638 1157 2644 1158
rect 2638 1153 2639 1157
rect 2643 1153 2644 1157
rect 2638 1152 2644 1153
rect 2766 1157 2772 1158
rect 2766 1153 2767 1157
rect 2771 1153 2772 1157
rect 2766 1152 2772 1153
rect 2910 1157 2916 1158
rect 2910 1153 2911 1157
rect 2915 1153 2916 1157
rect 2910 1152 2916 1153
rect 3070 1157 3076 1158
rect 3070 1153 3071 1157
rect 3075 1153 3076 1157
rect 3070 1152 3076 1153
rect 3246 1157 3252 1158
rect 3246 1153 3247 1157
rect 3251 1153 3252 1157
rect 3246 1152 3252 1153
rect 3438 1157 3444 1158
rect 3438 1153 3439 1157
rect 3443 1153 3444 1157
rect 3438 1152 3444 1153
rect 3630 1157 3636 1158
rect 3630 1153 3631 1157
rect 3635 1153 3636 1157
rect 3630 1152 3636 1153
rect 3830 1157 3836 1158
rect 3830 1153 3831 1157
rect 3835 1153 3836 1157
rect 3830 1152 3836 1153
rect 3942 1156 3948 1157
rect 3942 1152 3943 1156
rect 3947 1152 3948 1156
rect 2046 1151 2052 1152
rect 3942 1151 3948 1152
rect 110 1147 116 1148
rect 2006 1147 2012 1148
rect 3378 1147 3384 1148
rect 3378 1146 3379 1147
rect 2980 1144 3379 1146
rect 2347 1139 2356 1140
rect 498 1135 504 1136
rect 450 1131 456 1132
rect 450 1127 451 1131
rect 455 1130 456 1131
rect 459 1131 465 1132
rect 459 1130 460 1131
rect 455 1128 460 1130
rect 455 1127 456 1128
rect 450 1126 456 1127
rect 459 1127 460 1128
rect 464 1127 465 1131
rect 498 1131 499 1135
rect 503 1134 504 1135
rect 627 1135 633 1136
rect 627 1134 628 1135
rect 503 1132 628 1134
rect 503 1131 504 1132
rect 498 1130 504 1131
rect 627 1131 628 1132
rect 632 1131 633 1135
rect 627 1130 633 1131
rect 795 1135 801 1136
rect 795 1131 796 1135
rect 800 1134 801 1135
rect 878 1135 884 1136
rect 878 1134 879 1135
rect 800 1132 879 1134
rect 800 1131 801 1132
rect 795 1130 801 1131
rect 878 1131 879 1132
rect 883 1131 884 1135
rect 878 1130 884 1131
rect 963 1135 969 1136
rect 963 1131 964 1135
rect 968 1134 969 1135
rect 1047 1135 1053 1136
rect 1047 1134 1048 1135
rect 968 1132 1048 1134
rect 968 1131 969 1132
rect 963 1130 969 1131
rect 1047 1131 1048 1132
rect 1052 1131 1053 1135
rect 1266 1135 1272 1136
rect 1047 1130 1053 1131
rect 1131 1131 1137 1132
rect 459 1126 465 1127
rect 1131 1127 1132 1131
rect 1136 1130 1137 1131
rect 1194 1131 1200 1132
rect 1194 1130 1195 1131
rect 1136 1128 1195 1130
rect 1136 1127 1137 1128
rect 1131 1126 1137 1127
rect 1194 1127 1195 1128
rect 1199 1127 1200 1131
rect 1266 1131 1267 1135
rect 1271 1134 1272 1135
rect 1283 1135 1289 1136
rect 1283 1134 1284 1135
rect 1271 1132 1284 1134
rect 1271 1131 1272 1132
rect 1266 1130 1272 1131
rect 1283 1131 1284 1132
rect 1288 1131 1289 1135
rect 1283 1130 1289 1131
rect 1322 1135 1328 1136
rect 1322 1131 1323 1135
rect 1327 1134 1328 1135
rect 1435 1135 1441 1136
rect 1435 1134 1436 1135
rect 1327 1132 1436 1134
rect 1327 1131 1328 1132
rect 1322 1130 1328 1131
rect 1435 1131 1436 1132
rect 1440 1131 1441 1135
rect 1618 1135 1624 1136
rect 1435 1130 1441 1131
rect 1579 1131 1588 1132
rect 1194 1126 1200 1127
rect 1579 1127 1580 1131
rect 1587 1127 1588 1131
rect 1618 1131 1619 1135
rect 1623 1134 1624 1135
rect 1723 1135 1729 1136
rect 1723 1134 1724 1135
rect 1623 1132 1724 1134
rect 1623 1131 1624 1132
rect 1618 1130 1624 1131
rect 1723 1131 1724 1132
rect 1728 1131 1729 1135
rect 1723 1130 1729 1131
rect 1762 1135 1768 1136
rect 1762 1131 1763 1135
rect 1767 1134 1768 1135
rect 1875 1135 1881 1136
rect 1875 1134 1876 1135
rect 1767 1132 1876 1134
rect 1767 1131 1768 1132
rect 1762 1130 1768 1131
rect 1875 1131 1876 1132
rect 1880 1131 1881 1135
rect 2347 1135 2348 1139
rect 2355 1135 2356 1139
rect 2347 1134 2356 1135
rect 2386 1139 2392 1140
rect 2386 1135 2387 1139
rect 2391 1138 2392 1139
rect 2451 1139 2457 1140
rect 2451 1138 2452 1139
rect 2391 1136 2452 1138
rect 2391 1135 2392 1136
rect 2386 1134 2392 1135
rect 2451 1135 2452 1136
rect 2456 1135 2457 1139
rect 2451 1134 2457 1135
rect 2490 1139 2496 1140
rect 2490 1135 2491 1139
rect 2495 1138 2496 1139
rect 2563 1139 2569 1140
rect 2563 1138 2564 1139
rect 2495 1136 2564 1138
rect 2495 1135 2496 1136
rect 2490 1134 2496 1135
rect 2563 1135 2564 1136
rect 2568 1135 2569 1139
rect 2563 1134 2569 1135
rect 2602 1139 2608 1140
rect 2602 1135 2603 1139
rect 2607 1138 2608 1139
rect 2675 1139 2681 1140
rect 2675 1138 2676 1139
rect 2607 1136 2676 1138
rect 2607 1135 2608 1136
rect 2602 1134 2608 1135
rect 2675 1135 2676 1136
rect 2680 1135 2681 1139
rect 2675 1134 2681 1135
rect 2714 1139 2720 1140
rect 2714 1135 2715 1139
rect 2719 1138 2720 1139
rect 2803 1139 2809 1140
rect 2803 1138 2804 1139
rect 2719 1136 2804 1138
rect 2719 1135 2720 1136
rect 2714 1134 2720 1135
rect 2803 1135 2804 1136
rect 2808 1135 2809 1139
rect 2803 1134 2809 1135
rect 2947 1139 2953 1140
rect 2947 1135 2948 1139
rect 2952 1138 2953 1139
rect 2980 1138 2982 1144
rect 3378 1143 3379 1144
rect 3383 1143 3384 1147
rect 3378 1142 3384 1143
rect 2952 1136 2982 1138
rect 2986 1139 2992 1140
rect 2952 1135 2953 1136
rect 2947 1134 2953 1135
rect 2986 1135 2987 1139
rect 2991 1138 2992 1139
rect 3107 1139 3113 1140
rect 3107 1138 3108 1139
rect 2991 1136 3108 1138
rect 2991 1135 2992 1136
rect 2986 1134 2992 1135
rect 3107 1135 3108 1136
rect 3112 1135 3113 1139
rect 3107 1134 3113 1135
rect 3223 1139 3229 1140
rect 3223 1135 3224 1139
rect 3228 1138 3229 1139
rect 3283 1139 3289 1140
rect 3283 1138 3284 1139
rect 3228 1136 3284 1138
rect 3228 1135 3229 1136
rect 3223 1134 3229 1135
rect 3283 1135 3284 1136
rect 3288 1135 3289 1139
rect 3283 1134 3289 1135
rect 3322 1139 3328 1140
rect 3322 1135 3323 1139
rect 3327 1138 3328 1139
rect 3475 1139 3481 1140
rect 3475 1138 3476 1139
rect 3327 1136 3476 1138
rect 3327 1135 3328 1136
rect 3322 1134 3328 1135
rect 3475 1135 3476 1136
rect 3480 1135 3481 1139
rect 3867 1139 3873 1140
rect 3475 1134 3481 1135
rect 3667 1135 3673 1136
rect 1875 1130 1881 1131
rect 3667 1131 3668 1135
rect 3672 1134 3673 1135
rect 3714 1135 3720 1136
rect 3714 1134 3715 1135
rect 3672 1132 3715 1134
rect 3672 1131 3673 1132
rect 3667 1130 3673 1131
rect 3714 1131 3715 1132
rect 3719 1131 3720 1135
rect 3867 1135 3868 1139
rect 3872 1138 3873 1139
rect 3882 1139 3888 1140
rect 3882 1138 3883 1139
rect 3872 1136 3883 1138
rect 3872 1135 3873 1136
rect 3867 1134 3873 1135
rect 3882 1135 3883 1136
rect 3887 1135 3888 1139
rect 3882 1134 3888 1135
rect 3714 1130 3720 1131
rect 1579 1126 1588 1127
rect 718 1123 724 1124
rect 718 1122 719 1123
rect 524 1120 719 1122
rect 524 1118 526 1120
rect 718 1119 719 1120
rect 723 1119 724 1123
rect 718 1118 724 1119
rect 2443 1119 2449 1120
rect 523 1117 529 1118
rect 386 1115 392 1116
rect 386 1111 387 1115
rect 391 1114 392 1115
rect 411 1115 417 1116
rect 411 1114 412 1115
rect 391 1112 412 1114
rect 391 1111 392 1112
rect 386 1110 392 1111
rect 411 1111 412 1112
rect 416 1111 417 1115
rect 523 1113 524 1117
rect 528 1113 529 1117
rect 523 1112 529 1113
rect 562 1115 568 1116
rect 411 1110 417 1111
rect 562 1111 563 1115
rect 567 1114 568 1115
rect 635 1115 641 1116
rect 635 1114 636 1115
rect 567 1112 636 1114
rect 567 1111 568 1112
rect 562 1110 568 1111
rect 635 1111 636 1112
rect 640 1111 641 1115
rect 635 1110 641 1111
rect 674 1115 680 1116
rect 674 1111 675 1115
rect 679 1114 680 1115
rect 747 1115 753 1116
rect 747 1114 748 1115
rect 679 1112 748 1114
rect 679 1111 680 1112
rect 674 1110 680 1111
rect 747 1111 748 1112
rect 752 1111 753 1115
rect 906 1115 912 1116
rect 747 1110 753 1111
rect 867 1113 873 1114
rect 867 1109 868 1113
rect 872 1109 873 1113
rect 906 1111 907 1115
rect 911 1114 912 1115
rect 1003 1115 1009 1116
rect 1003 1114 1004 1115
rect 911 1112 1004 1114
rect 911 1111 912 1112
rect 906 1110 912 1111
rect 1003 1111 1004 1112
rect 1008 1111 1009 1115
rect 1003 1110 1009 1111
rect 1042 1115 1048 1116
rect 1042 1111 1043 1115
rect 1047 1114 1048 1115
rect 1155 1115 1161 1116
rect 1155 1114 1156 1115
rect 1047 1112 1156 1114
rect 1047 1111 1048 1112
rect 1042 1110 1048 1111
rect 1155 1111 1156 1112
rect 1160 1111 1161 1115
rect 1155 1110 1161 1111
rect 1315 1115 1321 1116
rect 1315 1111 1316 1115
rect 1320 1114 1321 1115
rect 1362 1115 1368 1116
rect 1362 1114 1363 1115
rect 1320 1112 1363 1114
rect 1320 1111 1321 1112
rect 1315 1110 1321 1111
rect 1362 1111 1363 1112
rect 1367 1111 1368 1115
rect 1362 1110 1368 1111
rect 1483 1115 1489 1116
rect 1483 1111 1484 1115
rect 1488 1114 1489 1115
rect 1498 1115 1504 1116
rect 1498 1114 1499 1115
rect 1488 1112 1499 1114
rect 1488 1111 1489 1112
rect 1483 1110 1489 1111
rect 1498 1111 1499 1112
rect 1503 1111 1504 1115
rect 1498 1110 1504 1111
rect 1535 1115 1541 1116
rect 1535 1111 1536 1115
rect 1540 1114 1541 1115
rect 1659 1115 1665 1116
rect 1659 1114 1660 1115
rect 1540 1112 1660 1114
rect 1540 1111 1541 1112
rect 1535 1110 1541 1111
rect 1659 1111 1660 1112
rect 1664 1111 1665 1115
rect 2443 1115 2444 1119
rect 2448 1118 2449 1119
rect 2474 1119 2480 1120
rect 2474 1118 2475 1119
rect 2448 1116 2475 1118
rect 2448 1115 2449 1116
rect 2443 1114 2449 1115
rect 2474 1115 2475 1116
rect 2479 1115 2480 1119
rect 2474 1114 2480 1115
rect 2482 1119 2488 1120
rect 2482 1115 2483 1119
rect 2487 1118 2488 1119
rect 2539 1119 2545 1120
rect 2539 1118 2540 1119
rect 2487 1116 2540 1118
rect 2487 1115 2488 1116
rect 2482 1114 2488 1115
rect 2539 1115 2540 1116
rect 2544 1115 2545 1119
rect 2539 1114 2545 1115
rect 2578 1119 2584 1120
rect 2578 1115 2579 1119
rect 2583 1118 2584 1119
rect 2635 1119 2641 1120
rect 2635 1118 2636 1119
rect 2583 1116 2636 1118
rect 2583 1115 2584 1116
rect 2578 1114 2584 1115
rect 2635 1115 2636 1116
rect 2640 1115 2641 1119
rect 2635 1114 2641 1115
rect 2674 1119 2680 1120
rect 2674 1115 2675 1119
rect 2679 1118 2680 1119
rect 2731 1119 2737 1120
rect 2731 1118 2732 1119
rect 2679 1116 2732 1118
rect 2679 1115 2680 1116
rect 2674 1114 2680 1115
rect 2731 1115 2732 1116
rect 2736 1115 2737 1119
rect 2731 1114 2737 1115
rect 2843 1119 2849 1120
rect 2843 1115 2844 1119
rect 2848 1118 2849 1119
rect 2902 1119 2908 1120
rect 2902 1118 2903 1119
rect 2848 1116 2903 1118
rect 2848 1115 2849 1116
rect 2843 1114 2849 1115
rect 2902 1115 2903 1116
rect 2907 1115 2908 1119
rect 3131 1119 3140 1120
rect 2902 1114 2908 1115
rect 2979 1117 2985 1118
rect 2979 1113 2980 1117
rect 2984 1113 2985 1117
rect 3131 1115 3132 1119
rect 3139 1115 3140 1119
rect 3131 1114 3140 1115
rect 3170 1119 3176 1120
rect 3170 1115 3171 1119
rect 3175 1118 3176 1119
rect 3299 1119 3305 1120
rect 3299 1118 3300 1119
rect 3175 1116 3300 1118
rect 3175 1115 3176 1116
rect 3170 1114 3176 1115
rect 3299 1115 3300 1116
rect 3304 1115 3305 1119
rect 3299 1114 3305 1115
rect 3338 1119 3344 1120
rect 3338 1115 3339 1119
rect 3343 1118 3344 1119
rect 3483 1119 3489 1120
rect 3483 1118 3484 1119
rect 3343 1116 3484 1118
rect 3343 1115 3344 1116
rect 3338 1114 3344 1115
rect 3483 1115 3484 1116
rect 3488 1115 3489 1119
rect 3483 1114 3489 1115
rect 3578 1119 3584 1120
rect 3578 1115 3579 1119
rect 3583 1118 3584 1119
rect 3675 1119 3681 1120
rect 3675 1118 3676 1119
rect 3583 1116 3676 1118
rect 3583 1115 3584 1116
rect 3578 1114 3584 1115
rect 3675 1115 3676 1116
rect 3680 1115 3681 1119
rect 3675 1114 3681 1115
rect 3875 1119 3881 1120
rect 3875 1115 3876 1119
rect 3880 1118 3881 1119
rect 3898 1119 3904 1120
rect 3898 1118 3899 1119
rect 3880 1116 3899 1118
rect 3880 1115 3881 1116
rect 3875 1114 3881 1115
rect 3898 1115 3899 1116
rect 3903 1115 3904 1119
rect 3898 1114 3904 1115
rect 2979 1112 2985 1113
rect 1659 1110 1665 1111
rect 2981 1110 2983 1112
rect 3142 1111 3148 1112
rect 3142 1110 3143 1111
rect 867 1108 873 1109
rect 2981 1108 3143 1110
rect 868 1106 870 1108
rect 1238 1107 1244 1108
rect 1238 1106 1239 1107
rect 868 1104 1239 1106
rect 1238 1103 1239 1104
rect 1243 1103 1244 1107
rect 3142 1107 3143 1108
rect 3147 1107 3148 1111
rect 3142 1106 3148 1107
rect 1238 1102 1244 1103
rect 2046 1100 2052 1101
rect 3942 1100 3948 1101
rect 110 1096 116 1097
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 486 1095 492 1096
rect 486 1091 487 1095
rect 491 1091 492 1095
rect 486 1090 492 1091
rect 598 1095 604 1096
rect 598 1091 599 1095
rect 603 1091 604 1095
rect 598 1090 604 1091
rect 710 1095 716 1096
rect 710 1091 711 1095
rect 715 1091 716 1095
rect 710 1090 716 1091
rect 830 1095 836 1096
rect 830 1091 831 1095
rect 835 1091 836 1095
rect 830 1090 836 1091
rect 966 1095 972 1096
rect 966 1091 967 1095
rect 971 1091 972 1095
rect 966 1090 972 1091
rect 1118 1095 1124 1096
rect 1118 1091 1119 1095
rect 1123 1091 1124 1095
rect 1118 1090 1124 1091
rect 1278 1095 1284 1096
rect 1278 1091 1279 1095
rect 1283 1091 1284 1095
rect 1278 1090 1284 1091
rect 1446 1095 1452 1096
rect 1446 1091 1447 1095
rect 1451 1091 1452 1095
rect 1446 1090 1452 1091
rect 1622 1095 1628 1096
rect 1622 1091 1623 1095
rect 1627 1091 1628 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2046 1096 2047 1100
rect 2051 1096 2052 1100
rect 2046 1095 2052 1096
rect 2406 1099 2412 1100
rect 2406 1095 2407 1099
rect 2411 1095 2412 1099
rect 2406 1094 2412 1095
rect 2502 1099 2508 1100
rect 2502 1095 2503 1099
rect 2507 1095 2508 1099
rect 2502 1094 2508 1095
rect 2598 1099 2604 1100
rect 2598 1095 2599 1099
rect 2603 1095 2604 1099
rect 2598 1094 2604 1095
rect 2694 1099 2700 1100
rect 2694 1095 2695 1099
rect 2699 1095 2700 1099
rect 2694 1094 2700 1095
rect 2806 1099 2812 1100
rect 2806 1095 2807 1099
rect 2811 1095 2812 1099
rect 2806 1094 2812 1095
rect 2942 1099 2948 1100
rect 2942 1095 2943 1099
rect 2947 1095 2948 1099
rect 2942 1094 2948 1095
rect 3094 1099 3100 1100
rect 3094 1095 3095 1099
rect 3099 1095 3100 1099
rect 3094 1094 3100 1095
rect 3262 1099 3268 1100
rect 3262 1095 3263 1099
rect 3267 1095 3268 1099
rect 3262 1094 3268 1095
rect 3446 1099 3452 1100
rect 3446 1095 3447 1099
rect 3451 1095 3452 1099
rect 3446 1094 3452 1095
rect 3638 1099 3644 1100
rect 3638 1095 3639 1099
rect 3643 1095 3644 1099
rect 3638 1094 3644 1095
rect 3838 1099 3844 1100
rect 3838 1095 3839 1099
rect 3843 1095 3844 1099
rect 3942 1096 3943 1100
rect 3947 1096 3948 1100
rect 3942 1095 3948 1096
rect 3838 1094 3844 1095
rect 2006 1091 2012 1092
rect 2482 1091 2488 1092
rect 1622 1090 1628 1091
rect 450 1087 456 1088
rect 450 1083 451 1087
rect 455 1083 456 1087
rect 450 1082 456 1083
rect 562 1087 568 1088
rect 562 1083 563 1087
rect 567 1083 568 1087
rect 562 1082 568 1083
rect 674 1087 680 1088
rect 674 1083 675 1087
rect 679 1083 680 1087
rect 906 1087 912 1088
rect 674 1082 680 1083
rect 786 1083 792 1084
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 786 1079 787 1083
rect 791 1079 792 1083
rect 906 1083 907 1087
rect 911 1083 912 1087
rect 906 1082 912 1083
rect 1042 1087 1048 1088
rect 1042 1083 1043 1087
rect 1047 1083 1048 1087
rect 1042 1082 1048 1083
rect 1194 1087 1200 1088
rect 1194 1083 1195 1087
rect 1199 1083 1200 1087
rect 1194 1082 1200 1083
rect 1238 1087 1244 1088
rect 1238 1083 1239 1087
rect 1243 1086 1244 1087
rect 1362 1087 1368 1088
rect 1243 1084 1321 1086
rect 1243 1083 1244 1084
rect 1238 1082 1244 1083
rect 1362 1083 1363 1087
rect 1367 1086 1368 1087
rect 1582 1087 1588 1088
rect 1367 1084 1489 1086
rect 1367 1083 1368 1084
rect 1362 1082 1368 1083
rect 1582 1083 1583 1087
rect 1587 1086 1588 1087
rect 2482 1087 2483 1091
rect 2487 1087 2488 1091
rect 2482 1086 2488 1087
rect 2578 1091 2584 1092
rect 2578 1087 2579 1091
rect 2583 1087 2584 1091
rect 2578 1086 2584 1087
rect 2674 1091 2680 1092
rect 2674 1087 2675 1091
rect 2679 1087 2680 1091
rect 2674 1086 2680 1087
rect 2682 1091 2688 1092
rect 2682 1087 2683 1091
rect 2687 1090 2688 1091
rect 2902 1091 2908 1092
rect 2687 1088 2737 1090
rect 2687 1087 2688 1088
rect 2682 1086 2688 1087
rect 2894 1087 2900 1088
rect 2894 1086 2895 1087
rect 1587 1084 1665 1086
rect 2885 1084 2895 1086
rect 1587 1083 1588 1084
rect 1582 1082 1588 1083
rect 2046 1083 2052 1084
rect 786 1078 792 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 486 1076 492 1077
rect 486 1072 487 1076
rect 491 1072 492 1076
rect 486 1071 492 1072
rect 598 1076 604 1077
rect 598 1072 599 1076
rect 603 1072 604 1076
rect 598 1071 604 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 830 1076 836 1077
rect 830 1072 831 1076
rect 835 1072 836 1076
rect 830 1071 836 1072
rect 966 1076 972 1077
rect 966 1072 967 1076
rect 971 1072 972 1076
rect 966 1071 972 1072
rect 1118 1076 1124 1077
rect 1118 1072 1119 1076
rect 1123 1072 1124 1076
rect 1118 1071 1124 1072
rect 1278 1076 1284 1077
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 1446 1076 1452 1077
rect 1446 1072 1447 1076
rect 1451 1072 1452 1076
rect 1446 1071 1452 1072
rect 1622 1076 1628 1077
rect 1622 1072 1623 1076
rect 1627 1072 1628 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2046 1079 2047 1083
rect 2051 1079 2052 1083
rect 2894 1083 2895 1084
rect 2899 1083 2900 1087
rect 2902 1087 2903 1091
rect 2907 1090 2908 1091
rect 3170 1091 3176 1092
rect 2907 1088 2985 1090
rect 2907 1087 2908 1088
rect 2902 1086 2908 1087
rect 3170 1087 3171 1091
rect 3175 1087 3176 1091
rect 3170 1086 3176 1087
rect 3338 1091 3344 1092
rect 3338 1087 3339 1091
rect 3343 1087 3344 1091
rect 3338 1086 3344 1087
rect 3382 1091 3388 1092
rect 3382 1087 3383 1091
rect 3387 1090 3388 1091
rect 3714 1091 3720 1092
rect 3387 1088 3489 1090
rect 3387 1087 3388 1088
rect 3382 1086 3388 1087
rect 3714 1087 3715 1091
rect 3719 1087 3720 1091
rect 3714 1086 3720 1087
rect 3914 1087 3920 1088
rect 2894 1082 2900 1083
rect 3914 1083 3915 1087
rect 3919 1083 3920 1087
rect 3914 1082 3920 1083
rect 3942 1083 3948 1084
rect 2046 1078 2052 1079
rect 2406 1080 2412 1081
rect 2406 1076 2407 1080
rect 2411 1076 2412 1080
rect 2406 1075 2412 1076
rect 2502 1080 2508 1081
rect 2502 1076 2503 1080
rect 2507 1076 2508 1080
rect 2502 1075 2508 1076
rect 2598 1080 2604 1081
rect 2598 1076 2599 1080
rect 2603 1076 2604 1080
rect 2598 1075 2604 1076
rect 2694 1080 2700 1081
rect 2694 1076 2695 1080
rect 2699 1076 2700 1080
rect 2694 1075 2700 1076
rect 2806 1080 2812 1081
rect 2806 1076 2807 1080
rect 2811 1076 2812 1080
rect 2806 1075 2812 1076
rect 2942 1080 2948 1081
rect 2942 1076 2943 1080
rect 2947 1076 2948 1080
rect 2942 1075 2948 1076
rect 3094 1080 3100 1081
rect 3094 1076 3095 1080
rect 3099 1076 3100 1080
rect 3094 1075 3100 1076
rect 3262 1080 3268 1081
rect 3262 1076 3263 1080
rect 3267 1076 3268 1080
rect 3262 1075 3268 1076
rect 3446 1080 3452 1081
rect 3446 1076 3447 1080
rect 3451 1076 3452 1080
rect 3446 1075 3452 1076
rect 3638 1080 3644 1081
rect 3638 1076 3639 1080
rect 3643 1076 3644 1080
rect 3638 1075 3644 1076
rect 3838 1080 3844 1081
rect 3838 1076 3839 1080
rect 3843 1076 3844 1080
rect 3942 1079 3943 1083
rect 3947 1079 3948 1083
rect 3942 1078 3948 1079
rect 3838 1075 3844 1076
rect 2006 1074 2012 1075
rect 1622 1071 1628 1072
rect 302 1016 308 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 302 1012 303 1016
rect 307 1012 308 1016
rect 302 1011 308 1012
rect 446 1016 452 1017
rect 446 1012 447 1016
rect 451 1012 452 1016
rect 446 1011 452 1012
rect 590 1016 596 1017
rect 590 1012 591 1016
rect 595 1012 596 1016
rect 590 1011 596 1012
rect 726 1016 732 1017
rect 726 1012 727 1016
rect 731 1012 732 1016
rect 726 1011 732 1012
rect 854 1016 860 1017
rect 854 1012 855 1016
rect 859 1012 860 1016
rect 854 1011 860 1012
rect 974 1016 980 1017
rect 974 1012 975 1016
rect 979 1012 980 1016
rect 974 1011 980 1012
rect 1086 1016 1092 1017
rect 1086 1012 1087 1016
rect 1091 1012 1092 1016
rect 1086 1011 1092 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1310 1016 1316 1017
rect 1310 1012 1311 1016
rect 1315 1012 1316 1016
rect 1310 1011 1316 1012
rect 1430 1016 1436 1017
rect 1430 1012 1431 1016
rect 1435 1012 1436 1016
rect 2454 1016 2460 1017
rect 1430 1011 1436 1012
rect 2006 1013 2012 1014
rect 110 1008 116 1009
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1013 2052 1014
rect 2046 1009 2047 1013
rect 2051 1009 2052 1013
rect 2454 1012 2455 1016
rect 2459 1012 2460 1016
rect 2454 1011 2460 1012
rect 2550 1016 2556 1017
rect 2550 1012 2551 1016
rect 2555 1012 2556 1016
rect 2550 1011 2556 1012
rect 2646 1016 2652 1017
rect 2646 1012 2647 1016
rect 2651 1012 2652 1016
rect 2646 1011 2652 1012
rect 2758 1016 2764 1017
rect 2758 1012 2759 1016
rect 2763 1012 2764 1016
rect 2758 1011 2764 1012
rect 2886 1016 2892 1017
rect 2886 1012 2887 1016
rect 2891 1012 2892 1016
rect 2886 1011 2892 1012
rect 3030 1016 3036 1017
rect 3030 1012 3031 1016
rect 3035 1012 3036 1016
rect 3030 1011 3036 1012
rect 3182 1016 3188 1017
rect 3182 1012 3183 1016
rect 3187 1012 3188 1016
rect 3182 1011 3188 1012
rect 3342 1016 3348 1017
rect 3342 1012 3343 1016
rect 3347 1012 3348 1016
rect 3342 1011 3348 1012
rect 3502 1016 3508 1017
rect 3502 1012 3503 1016
rect 3507 1012 3508 1016
rect 3502 1011 3508 1012
rect 3670 1016 3676 1017
rect 3670 1012 3671 1016
rect 3675 1012 3676 1016
rect 3670 1011 3676 1012
rect 3838 1016 3844 1017
rect 3838 1012 3839 1016
rect 3843 1012 3844 1016
rect 3838 1011 3844 1012
rect 3942 1013 3948 1014
rect 2046 1008 2052 1009
rect 3942 1009 3943 1013
rect 3947 1009 3948 1013
rect 3942 1008 3948 1009
rect 386 1007 392 1008
rect 386 1006 387 1007
rect 381 1004 387 1006
rect 386 1003 387 1004
rect 391 1003 392 1007
rect 386 1002 392 1003
rect 394 1007 400 1008
rect 394 1003 395 1007
rect 399 1006 400 1007
rect 666 1007 672 1008
rect 399 1004 489 1006
rect 399 1003 400 1004
rect 394 1002 400 1003
rect 666 1003 667 1007
rect 671 1003 672 1007
rect 666 1002 672 1003
rect 802 1007 808 1008
rect 802 1003 803 1007
rect 807 1003 808 1007
rect 802 1002 808 1003
rect 810 1007 816 1008
rect 810 1003 811 1007
rect 815 1006 816 1007
rect 1050 1007 1056 1008
rect 815 1004 897 1006
rect 815 1003 816 1004
rect 810 1002 816 1003
rect 1050 1003 1051 1007
rect 1055 1003 1056 1007
rect 1050 1002 1056 1003
rect 1162 1007 1168 1008
rect 1162 1003 1163 1007
rect 1167 1003 1168 1007
rect 1162 1002 1168 1003
rect 1274 1007 1280 1008
rect 1274 1003 1275 1007
rect 1279 1003 1280 1007
rect 1274 1002 1280 1003
rect 1386 1007 1392 1008
rect 1386 1003 1387 1007
rect 1391 1003 1392 1007
rect 1386 1002 1392 1003
rect 1498 1007 1504 1008
rect 1498 1003 1499 1007
rect 1503 1003 1504 1007
rect 1498 1002 1504 1003
rect 2447 1007 2453 1008
rect 2447 1003 2448 1007
rect 2452 1006 2453 1007
rect 2542 1007 2548 1008
rect 2452 1004 2497 1006
rect 2452 1003 2453 1004
rect 2447 1002 2453 1003
rect 2542 1003 2543 1007
rect 2547 1006 2548 1007
rect 2722 1007 2728 1008
rect 2547 1004 2593 1006
rect 2547 1003 2548 1004
rect 2542 1002 2548 1003
rect 2722 1003 2723 1007
rect 2727 1003 2728 1007
rect 2722 1002 2728 1003
rect 2834 1007 2840 1008
rect 2834 1003 2835 1007
rect 2839 1003 2840 1007
rect 2834 1002 2840 1003
rect 2858 1007 2864 1008
rect 2858 1003 2859 1007
rect 2863 1006 2864 1007
rect 2990 1007 2996 1008
rect 2863 1004 2929 1006
rect 2863 1003 2864 1004
rect 2858 1002 2864 1003
rect 2990 1003 2991 1007
rect 2995 1006 2996 1007
rect 3142 1007 3148 1008
rect 2995 1004 3073 1006
rect 2995 1003 2996 1004
rect 2990 1002 2996 1003
rect 3142 1003 3143 1007
rect 3147 1006 3148 1007
rect 3294 1007 3300 1008
rect 3147 1004 3225 1006
rect 3147 1003 3148 1004
rect 3142 1002 3148 1003
rect 3294 1003 3295 1007
rect 3299 1006 3300 1007
rect 3578 1007 3584 1008
rect 3299 1004 3385 1006
rect 3299 1003 3300 1004
rect 3294 1002 3300 1003
rect 3578 1003 3579 1007
rect 3583 1003 3584 1007
rect 3578 1002 3584 1003
rect 3591 1007 3597 1008
rect 3591 1003 3592 1007
rect 3596 1006 3597 1007
rect 3906 1007 3912 1008
rect 3596 1004 3713 1006
rect 3596 1003 3597 1004
rect 3591 1002 3597 1003
rect 3906 1003 3907 1007
rect 3911 1003 3912 1007
rect 3906 1002 3912 1003
rect 302 997 308 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 302 993 303 997
rect 307 993 308 997
rect 302 992 308 993
rect 446 997 452 998
rect 446 993 447 997
rect 451 993 452 997
rect 446 992 452 993
rect 590 997 596 998
rect 590 993 591 997
rect 595 993 596 997
rect 590 992 596 993
rect 726 997 732 998
rect 726 993 727 997
rect 731 993 732 997
rect 726 992 732 993
rect 854 997 860 998
rect 854 993 855 997
rect 859 993 860 997
rect 854 992 860 993
rect 974 997 980 998
rect 974 993 975 997
rect 979 993 980 997
rect 974 992 980 993
rect 1086 997 1092 998
rect 1086 993 1087 997
rect 1091 993 1092 997
rect 1086 992 1092 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1310 997 1316 998
rect 1310 993 1311 997
rect 1315 993 1316 997
rect 1310 992 1316 993
rect 1430 997 1436 998
rect 2454 997 2460 998
rect 1430 993 1431 997
rect 1435 993 1436 997
rect 1430 992 1436 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 2006 991 2012 992
rect 2046 996 2052 997
rect 2046 992 2047 996
rect 2051 992 2052 996
rect 2454 993 2455 997
rect 2459 993 2460 997
rect 2454 992 2460 993
rect 2550 997 2556 998
rect 2550 993 2551 997
rect 2555 993 2556 997
rect 2550 992 2556 993
rect 2646 997 2652 998
rect 2646 993 2647 997
rect 2651 993 2652 997
rect 2646 992 2652 993
rect 2758 997 2764 998
rect 2758 993 2759 997
rect 2763 993 2764 997
rect 2758 992 2764 993
rect 2886 997 2892 998
rect 2886 993 2887 997
rect 2891 993 2892 997
rect 2886 992 2892 993
rect 3030 997 3036 998
rect 3030 993 3031 997
rect 3035 993 3036 997
rect 3030 992 3036 993
rect 3182 997 3188 998
rect 3182 993 3183 997
rect 3187 993 3188 997
rect 3182 992 3188 993
rect 3342 997 3348 998
rect 3342 993 3343 997
rect 3347 993 3348 997
rect 3342 992 3348 993
rect 3502 997 3508 998
rect 3502 993 3503 997
rect 3507 993 3508 997
rect 3502 992 3508 993
rect 3670 997 3676 998
rect 3670 993 3671 997
rect 3675 993 3676 997
rect 3670 992 3676 993
rect 3838 997 3844 998
rect 3838 993 3839 997
rect 3843 993 3844 997
rect 3838 992 3844 993
rect 3942 996 3948 997
rect 3942 992 3943 996
rect 3947 992 3948 996
rect 2046 991 2052 992
rect 3942 991 3948 992
rect 810 987 816 988
rect 810 986 811 987
rect 756 984 811 986
rect 339 979 345 980
rect 339 975 340 979
rect 344 978 345 979
rect 394 979 400 980
rect 394 978 395 979
rect 344 976 395 978
rect 344 975 345 976
rect 339 974 345 975
rect 394 975 395 976
rect 399 975 400 979
rect 627 979 633 980
rect 394 974 400 975
rect 483 975 489 976
rect 483 971 484 975
rect 488 974 489 975
rect 522 975 528 976
rect 522 974 523 975
rect 488 972 523 974
rect 488 971 489 972
rect 483 970 489 971
rect 522 971 523 972
rect 527 971 528 975
rect 627 975 628 979
rect 632 978 633 979
rect 756 978 758 984
rect 810 983 811 984
rect 815 983 816 987
rect 2682 987 2688 988
rect 2682 986 2683 987
rect 810 982 816 983
rect 2664 984 2683 986
rect 632 976 758 978
rect 763 979 769 980
rect 632 975 633 976
rect 627 974 633 975
rect 763 975 764 979
rect 768 978 769 979
rect 786 979 792 980
rect 786 978 787 979
rect 768 976 787 978
rect 768 975 769 976
rect 763 974 769 975
rect 786 975 787 976
rect 791 975 792 979
rect 786 974 792 975
rect 802 979 808 980
rect 802 975 803 979
rect 807 978 808 979
rect 891 979 897 980
rect 891 978 892 979
rect 807 976 892 978
rect 807 975 808 976
rect 802 974 808 975
rect 891 975 892 976
rect 896 975 897 979
rect 1050 979 1056 980
rect 891 974 897 975
rect 1011 975 1017 976
rect 522 970 528 971
rect 1011 971 1012 975
rect 1016 974 1017 975
rect 1042 975 1048 976
rect 1042 974 1043 975
rect 1016 972 1043 974
rect 1016 971 1017 972
rect 1011 970 1017 971
rect 1042 971 1043 972
rect 1047 971 1048 975
rect 1050 975 1051 979
rect 1055 978 1056 979
rect 1123 979 1129 980
rect 1123 978 1124 979
rect 1055 976 1124 978
rect 1055 975 1056 976
rect 1050 974 1056 975
rect 1123 975 1124 976
rect 1128 975 1129 979
rect 1123 974 1129 975
rect 1162 979 1168 980
rect 1162 975 1163 979
rect 1167 978 1168 979
rect 1235 979 1241 980
rect 1235 978 1236 979
rect 1167 976 1236 978
rect 1167 975 1168 976
rect 1162 974 1168 975
rect 1235 975 1236 976
rect 1240 975 1241 979
rect 1235 974 1241 975
rect 1274 979 1280 980
rect 1274 975 1275 979
rect 1279 978 1280 979
rect 1347 979 1353 980
rect 1347 978 1348 979
rect 1279 976 1348 978
rect 1279 975 1280 976
rect 1274 974 1280 975
rect 1347 975 1348 976
rect 1352 975 1353 979
rect 1347 974 1353 975
rect 1386 979 1392 980
rect 1386 975 1387 979
rect 1391 978 1392 979
rect 1467 979 1473 980
rect 1467 978 1468 979
rect 1391 976 1468 978
rect 1391 975 1392 976
rect 1386 974 1392 975
rect 1467 975 1468 976
rect 1472 975 1473 979
rect 1467 974 1473 975
rect 2491 979 2497 980
rect 2491 975 2492 979
rect 2496 978 2497 979
rect 2542 979 2548 980
rect 2542 978 2543 979
rect 2496 976 2543 978
rect 2496 975 2497 976
rect 2491 974 2497 975
rect 2542 975 2543 976
rect 2547 975 2548 979
rect 2542 974 2548 975
rect 2587 979 2593 980
rect 2587 975 2588 979
rect 2592 978 2593 979
rect 2664 978 2666 984
rect 2682 983 2683 984
rect 2687 983 2688 987
rect 2682 982 2688 983
rect 2858 983 2864 984
rect 2858 982 2859 983
rect 2732 980 2859 982
rect 2592 976 2666 978
rect 2683 979 2689 980
rect 2592 975 2593 976
rect 2587 974 2593 975
rect 2683 975 2684 979
rect 2688 978 2689 979
rect 2732 978 2734 980
rect 2858 979 2859 980
rect 2863 979 2864 983
rect 2858 978 2864 979
rect 2894 979 2900 980
rect 2688 976 2734 978
rect 2688 975 2689 976
rect 2683 974 2689 975
rect 2786 975 2792 976
rect 1042 970 1048 971
rect 2786 971 2787 975
rect 2791 974 2792 975
rect 2795 975 2801 976
rect 2795 974 2796 975
rect 2791 972 2796 974
rect 2791 971 2792 972
rect 2786 970 2792 971
rect 2795 971 2796 972
rect 2800 971 2801 975
rect 2894 975 2895 979
rect 2899 978 2900 979
rect 2923 979 2929 980
rect 2923 978 2924 979
rect 2899 976 2924 978
rect 2899 975 2900 976
rect 2894 974 2900 975
rect 2923 975 2924 976
rect 2928 975 2929 979
rect 3219 979 3225 980
rect 2923 974 2929 975
rect 2942 975 2948 976
rect 2795 970 2801 971
rect 2942 971 2943 975
rect 2947 974 2948 975
rect 3067 975 3073 976
rect 3067 974 3068 975
rect 2947 972 3068 974
rect 2947 971 2948 972
rect 2942 970 2948 971
rect 3067 971 3068 972
rect 3072 971 3073 975
rect 3219 975 3220 979
rect 3224 978 3225 979
rect 3294 979 3300 980
rect 3294 978 3295 979
rect 3224 976 3295 978
rect 3224 975 3225 976
rect 3219 974 3225 975
rect 3294 975 3295 976
rect 3299 975 3300 979
rect 3294 974 3300 975
rect 3379 979 3388 980
rect 3379 975 3380 979
rect 3387 975 3388 979
rect 3379 974 3388 975
rect 3539 979 3545 980
rect 3539 975 3540 979
rect 3544 978 3545 979
rect 3591 979 3597 980
rect 3591 978 3592 979
rect 3544 976 3592 978
rect 3544 975 3545 976
rect 3539 974 3545 975
rect 3591 975 3592 976
rect 3596 975 3597 979
rect 3875 979 3881 980
rect 3591 974 3597 975
rect 3707 975 3713 976
rect 3067 970 3073 971
rect 3707 971 3708 975
rect 3712 974 3713 975
rect 3722 975 3728 976
rect 3722 974 3723 975
rect 3712 972 3723 974
rect 3712 971 3713 972
rect 3707 970 3713 971
rect 3722 971 3723 972
rect 3727 971 3728 975
rect 3875 975 3876 979
rect 3880 978 3881 979
rect 3914 979 3920 980
rect 3914 978 3915 979
rect 3880 976 3915 978
rect 3880 975 3881 976
rect 3875 974 3881 975
rect 3914 975 3915 976
rect 3919 975 3920 979
rect 3914 974 3920 975
rect 3722 970 3728 971
rect 291 963 297 964
rect 291 959 292 963
rect 296 962 297 963
rect 322 963 328 964
rect 322 962 323 963
rect 296 960 323 962
rect 296 959 297 960
rect 291 958 297 959
rect 322 959 323 960
rect 327 959 328 963
rect 322 958 328 959
rect 330 963 336 964
rect 330 959 331 963
rect 335 962 336 963
rect 483 963 489 964
rect 483 962 484 963
rect 335 960 484 962
rect 335 959 336 960
rect 330 958 336 959
rect 483 959 484 960
rect 488 959 489 963
rect 483 958 489 959
rect 666 963 673 964
rect 666 959 667 963
rect 672 959 673 963
rect 666 958 673 959
rect 706 963 712 964
rect 706 959 707 963
rect 711 962 712 963
rect 843 963 849 964
rect 843 962 844 963
rect 711 960 844 962
rect 711 959 712 960
rect 706 958 712 959
rect 843 959 844 960
rect 848 959 849 963
rect 843 958 849 959
rect 882 963 888 964
rect 882 959 883 963
rect 887 962 888 963
rect 1011 963 1017 964
rect 1011 962 1012 963
rect 887 960 1012 962
rect 887 959 888 960
rect 882 958 888 959
rect 1011 959 1012 960
rect 1016 959 1017 963
rect 1011 958 1017 959
rect 1163 963 1169 964
rect 1163 959 1164 963
rect 1168 962 1169 963
rect 1210 963 1216 964
rect 1210 962 1211 963
rect 1168 960 1211 962
rect 1168 959 1169 960
rect 1163 958 1169 959
rect 1210 959 1211 960
rect 1215 959 1216 963
rect 1210 958 1216 959
rect 1307 963 1313 964
rect 1307 959 1308 963
rect 1312 962 1313 963
rect 1354 963 1360 964
rect 1354 962 1355 963
rect 1312 960 1355 962
rect 1312 959 1313 960
rect 1307 958 1313 959
rect 1354 959 1355 960
rect 1359 959 1360 963
rect 1354 958 1360 959
rect 1451 963 1457 964
rect 1451 959 1452 963
rect 1456 962 1457 963
rect 1498 963 1504 964
rect 1498 962 1499 963
rect 1456 960 1499 962
rect 1456 959 1457 960
rect 1451 958 1457 959
rect 1498 959 1499 960
rect 1503 959 1504 963
rect 1498 958 1504 959
rect 1587 963 1593 964
rect 1587 959 1588 963
rect 1592 962 1593 963
rect 1634 963 1640 964
rect 1634 962 1635 963
rect 1592 960 1635 962
rect 1592 959 1593 960
rect 1587 958 1593 959
rect 1634 959 1635 960
rect 1639 959 1640 963
rect 1634 958 1640 959
rect 1731 963 1740 964
rect 1731 959 1732 963
rect 1739 959 1740 963
rect 1731 958 1740 959
rect 2447 959 2453 960
rect 2447 955 2448 959
rect 2452 958 2453 959
rect 2459 959 2465 960
rect 2459 958 2460 959
rect 2452 956 2460 958
rect 2452 955 2453 956
rect 2447 954 2453 955
rect 2459 955 2460 956
rect 2464 955 2465 959
rect 2459 954 2465 955
rect 2498 959 2504 960
rect 2498 955 2499 959
rect 2503 958 2504 959
rect 2555 959 2561 960
rect 2555 958 2556 959
rect 2503 956 2556 958
rect 2503 955 2504 956
rect 2498 954 2504 955
rect 2555 955 2556 956
rect 2560 955 2561 959
rect 2555 954 2561 955
rect 2594 959 2600 960
rect 2594 955 2595 959
rect 2599 958 2600 959
rect 2651 959 2657 960
rect 2651 958 2652 959
rect 2599 956 2652 958
rect 2599 955 2600 956
rect 2594 954 2600 955
rect 2651 955 2652 956
rect 2656 955 2657 959
rect 2651 954 2657 955
rect 2722 959 2728 960
rect 2722 955 2723 959
rect 2727 958 2728 959
rect 2747 959 2753 960
rect 2747 958 2748 959
rect 2727 956 2748 958
rect 2727 955 2728 956
rect 2722 954 2728 955
rect 2747 955 2748 956
rect 2752 955 2753 959
rect 2747 954 2753 955
rect 2834 959 2840 960
rect 2834 955 2835 959
rect 2839 958 2840 959
rect 2859 959 2865 960
rect 2859 958 2860 959
rect 2839 956 2860 958
rect 2839 955 2840 956
rect 2834 954 2840 955
rect 2859 955 2860 956
rect 2864 955 2865 959
rect 2859 954 2865 955
rect 2987 959 2996 960
rect 2987 955 2988 959
rect 2995 955 2996 959
rect 2987 954 2996 955
rect 3046 959 3052 960
rect 3046 955 3047 959
rect 3051 958 3052 959
rect 3139 959 3145 960
rect 3139 958 3140 959
rect 3051 956 3140 958
rect 3051 955 3052 956
rect 3046 954 3052 955
rect 3139 955 3140 956
rect 3144 955 3145 959
rect 3139 954 3145 955
rect 3223 959 3229 960
rect 3223 955 3224 959
rect 3228 958 3229 959
rect 3307 959 3313 960
rect 3307 958 3308 959
rect 3228 956 3308 958
rect 3228 955 3229 956
rect 3223 954 3229 955
rect 3307 955 3308 956
rect 3312 955 3313 959
rect 3307 954 3313 955
rect 3399 959 3405 960
rect 3399 955 3400 959
rect 3404 958 3405 959
rect 3491 959 3497 960
rect 3491 958 3492 959
rect 3404 956 3492 958
rect 3404 955 3405 956
rect 3399 954 3405 955
rect 3491 955 3492 956
rect 3496 955 3497 959
rect 3491 954 3497 955
rect 3683 959 3692 960
rect 3683 955 3684 959
rect 3691 955 3692 959
rect 3683 954 3692 955
rect 3875 959 3881 960
rect 3875 955 3876 959
rect 3880 958 3881 959
rect 3906 959 3912 960
rect 3906 958 3907 959
rect 3880 956 3907 958
rect 3880 955 3881 956
rect 3875 954 3881 955
rect 3906 955 3907 956
rect 3911 955 3912 959
rect 3906 954 3912 955
rect 110 944 116 945
rect 2006 944 2012 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 254 943 260 944
rect 254 939 255 943
rect 259 939 260 943
rect 254 938 260 939
rect 446 943 452 944
rect 446 939 447 943
rect 451 939 452 943
rect 446 938 452 939
rect 630 943 636 944
rect 630 939 631 943
rect 635 939 636 943
rect 630 938 636 939
rect 806 943 812 944
rect 806 939 807 943
rect 811 939 812 943
rect 806 938 812 939
rect 974 943 980 944
rect 974 939 975 943
rect 979 939 980 943
rect 1126 943 1132 944
rect 974 938 980 939
rect 1042 939 1048 940
rect 330 935 336 936
rect 330 931 331 935
rect 335 931 336 935
rect 330 930 336 931
rect 522 935 528 936
rect 522 931 523 935
rect 527 931 528 935
rect 522 930 528 931
rect 706 935 712 936
rect 706 931 707 935
rect 711 931 712 935
rect 706 930 712 931
rect 882 935 888 936
rect 882 931 883 935
rect 887 931 888 935
rect 1042 935 1043 939
rect 1047 938 1048 939
rect 1126 939 1127 943
rect 1131 939 1132 943
rect 1126 938 1132 939
rect 1270 943 1276 944
rect 1270 939 1271 943
rect 1275 939 1276 943
rect 1270 938 1276 939
rect 1414 943 1420 944
rect 1414 939 1415 943
rect 1419 939 1420 943
rect 1414 938 1420 939
rect 1550 943 1556 944
rect 1550 939 1551 943
rect 1555 939 1556 943
rect 1550 938 1556 939
rect 1694 943 1700 944
rect 1694 939 1695 943
rect 1699 939 1700 943
rect 2006 940 2007 944
rect 2011 940 2012 944
rect 2006 939 2012 940
rect 2046 940 2052 941
rect 3942 940 3948 941
rect 1694 938 1700 939
rect 1047 936 1102 938
rect 2046 936 2047 940
rect 2051 936 2052 940
rect 1047 935 1048 936
rect 1042 934 1048 935
rect 1100 934 1102 936
rect 1210 935 1216 936
rect 1100 932 1169 934
rect 882 930 888 931
rect 1050 931 1056 932
rect 110 927 116 928
rect 110 923 111 927
rect 115 923 116 927
rect 1050 927 1051 931
rect 1055 927 1056 931
rect 1210 931 1211 935
rect 1215 934 1216 935
rect 1354 935 1360 936
rect 1215 932 1313 934
rect 1215 931 1216 932
rect 1210 930 1216 931
rect 1354 931 1355 935
rect 1359 934 1360 935
rect 1498 935 1504 936
rect 1359 932 1457 934
rect 1359 931 1360 932
rect 1354 930 1360 931
rect 1498 931 1499 935
rect 1503 934 1504 935
rect 1634 935 1640 936
rect 2046 935 2052 936
rect 2422 939 2428 940
rect 2422 935 2423 939
rect 2427 935 2428 939
rect 1503 932 1593 934
rect 1503 931 1504 932
rect 1498 930 1504 931
rect 1634 931 1635 935
rect 1639 934 1640 935
rect 2422 934 2428 935
rect 2518 939 2524 940
rect 2518 935 2519 939
rect 2523 935 2524 939
rect 2518 934 2524 935
rect 2614 939 2620 940
rect 2614 935 2615 939
rect 2619 935 2620 939
rect 2614 934 2620 935
rect 2710 939 2716 940
rect 2710 935 2711 939
rect 2715 935 2716 939
rect 2710 934 2716 935
rect 2822 939 2828 940
rect 2822 935 2823 939
rect 2827 935 2828 939
rect 2822 934 2828 935
rect 2950 939 2956 940
rect 2950 935 2951 939
rect 2955 935 2956 939
rect 2950 934 2956 935
rect 3102 939 3108 940
rect 3102 935 3103 939
rect 3107 935 3108 939
rect 3102 934 3108 935
rect 3270 939 3276 940
rect 3270 935 3271 939
rect 3275 935 3276 939
rect 3270 934 3276 935
rect 3454 939 3460 940
rect 3454 935 3455 939
rect 3459 935 3460 939
rect 3454 934 3460 935
rect 3646 939 3652 940
rect 3646 935 3647 939
rect 3651 935 3652 939
rect 3646 934 3652 935
rect 3838 939 3844 940
rect 3838 935 3839 939
rect 3843 935 3844 939
rect 3942 936 3943 940
rect 3947 936 3948 940
rect 3942 935 3948 936
rect 3838 934 3844 935
rect 1639 932 1737 934
rect 1639 931 1640 932
rect 1634 930 1640 931
rect 2498 931 2504 932
rect 1050 926 1056 927
rect 2006 927 2012 928
rect 110 922 116 923
rect 254 924 260 925
rect 254 920 255 924
rect 259 920 260 924
rect 254 919 260 920
rect 446 924 452 925
rect 446 920 447 924
rect 451 920 452 924
rect 446 919 452 920
rect 630 924 636 925
rect 630 920 631 924
rect 635 920 636 924
rect 630 919 636 920
rect 806 924 812 925
rect 806 920 807 924
rect 811 920 812 924
rect 806 919 812 920
rect 974 924 980 925
rect 974 920 975 924
rect 979 920 980 924
rect 974 919 980 920
rect 1126 924 1132 925
rect 1126 920 1127 924
rect 1131 920 1132 924
rect 1126 919 1132 920
rect 1270 924 1276 925
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1414 924 1420 925
rect 1414 920 1415 924
rect 1419 920 1420 924
rect 1414 919 1420 920
rect 1550 924 1556 925
rect 1550 920 1551 924
rect 1555 920 1556 924
rect 1550 919 1556 920
rect 1694 924 1700 925
rect 1694 920 1695 924
rect 1699 920 1700 924
rect 2006 923 2007 927
rect 2011 923 2012 927
rect 2498 927 2499 931
rect 2503 927 2504 931
rect 2498 926 2504 927
rect 2594 931 2600 932
rect 2594 927 2595 931
rect 2599 927 2600 931
rect 2786 931 2792 932
rect 2594 926 2600 927
rect 2690 927 2696 928
rect 2006 922 2012 923
rect 2046 923 2052 924
rect 1694 919 1700 920
rect 2046 919 2047 923
rect 2051 919 2052 923
rect 2690 923 2691 927
rect 2695 923 2696 927
rect 2786 927 2787 931
rect 2791 927 2792 931
rect 2942 931 2948 932
rect 2942 930 2943 931
rect 2901 928 2943 930
rect 2786 926 2792 927
rect 2942 927 2943 928
rect 2947 927 2948 931
rect 3046 931 3052 932
rect 3046 930 3047 931
rect 3029 928 3047 930
rect 2942 926 2948 927
rect 3046 927 3047 928
rect 3051 927 3052 931
rect 3223 931 3229 932
rect 3223 930 3224 931
rect 3181 928 3224 930
rect 3046 926 3052 927
rect 3223 927 3224 928
rect 3228 927 3229 931
rect 3399 931 3405 932
rect 3399 930 3400 931
rect 3349 928 3400 930
rect 3223 926 3229 927
rect 3399 927 3400 928
rect 3404 927 3405 931
rect 3399 926 3405 927
rect 3410 931 3416 932
rect 3410 927 3411 931
rect 3415 930 3416 931
rect 3722 931 3728 932
rect 3415 928 3497 930
rect 3415 927 3416 928
rect 3410 926 3416 927
rect 3722 927 3723 931
rect 3727 927 3728 931
rect 3722 926 3728 927
rect 3914 927 3920 928
rect 2690 922 2696 923
rect 3914 923 3915 927
rect 3919 923 3920 927
rect 3914 922 3920 923
rect 3942 923 3948 924
rect 2046 918 2052 919
rect 2422 920 2428 921
rect 2422 916 2423 920
rect 2427 916 2428 920
rect 2422 915 2428 916
rect 2518 920 2524 921
rect 2518 916 2519 920
rect 2523 916 2524 920
rect 2518 915 2524 916
rect 2614 920 2620 921
rect 2614 916 2615 920
rect 2619 916 2620 920
rect 2614 915 2620 916
rect 2710 920 2716 921
rect 2710 916 2711 920
rect 2715 916 2716 920
rect 2710 915 2716 916
rect 2822 920 2828 921
rect 2822 916 2823 920
rect 2827 916 2828 920
rect 2822 915 2828 916
rect 2950 920 2956 921
rect 2950 916 2951 920
rect 2955 916 2956 920
rect 2950 915 2956 916
rect 3102 920 3108 921
rect 3102 916 3103 920
rect 3107 916 3108 920
rect 3102 915 3108 916
rect 3270 920 3276 921
rect 3270 916 3271 920
rect 3275 916 3276 920
rect 3270 915 3276 916
rect 3454 920 3460 921
rect 3454 916 3455 920
rect 3459 916 3460 920
rect 3454 915 3460 916
rect 3646 920 3652 921
rect 3646 916 3647 920
rect 3651 916 3652 920
rect 3646 915 3652 916
rect 3838 920 3844 921
rect 3838 916 3839 920
rect 3843 916 3844 920
rect 3942 919 3943 923
rect 3947 919 3948 923
rect 3942 918 3948 919
rect 3838 915 3844 916
rect 254 860 260 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 254 856 255 860
rect 259 856 260 860
rect 254 855 260 856
rect 446 860 452 861
rect 446 856 447 860
rect 451 856 452 860
rect 446 855 452 856
rect 638 860 644 861
rect 638 856 639 860
rect 643 856 644 860
rect 638 855 644 856
rect 822 860 828 861
rect 822 856 823 860
rect 827 856 828 860
rect 822 855 828 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1166 860 1172 861
rect 1166 856 1167 860
rect 1171 856 1172 860
rect 1166 855 1172 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1478 860 1484 861
rect 1478 856 1479 860
rect 1483 856 1484 860
rect 1478 855 1484 856
rect 1630 860 1636 861
rect 1630 856 1631 860
rect 1635 856 1636 860
rect 1630 855 1636 856
rect 1782 860 1788 861
rect 1782 856 1783 860
rect 1787 856 1788 860
rect 2342 860 2348 861
rect 1782 855 1788 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2006 852 2012 853
rect 2046 857 2052 858
rect 2046 853 2047 857
rect 2051 853 2052 857
rect 2342 856 2343 860
rect 2347 856 2348 860
rect 2342 855 2348 856
rect 2438 860 2444 861
rect 2438 856 2439 860
rect 2443 856 2444 860
rect 2438 855 2444 856
rect 2534 860 2540 861
rect 2534 856 2535 860
rect 2539 856 2540 860
rect 2534 855 2540 856
rect 2630 860 2636 861
rect 2630 856 2631 860
rect 2635 856 2636 860
rect 2630 855 2636 856
rect 2734 860 2740 861
rect 2734 856 2735 860
rect 2739 856 2740 860
rect 2734 855 2740 856
rect 2862 860 2868 861
rect 2862 856 2863 860
rect 2867 856 2868 860
rect 2862 855 2868 856
rect 3014 860 3020 861
rect 3014 856 3015 860
rect 3019 856 3020 860
rect 3014 855 3020 856
rect 3190 860 3196 861
rect 3190 856 3191 860
rect 3195 856 3196 860
rect 3190 855 3196 856
rect 3390 860 3396 861
rect 3390 856 3391 860
rect 3395 856 3396 860
rect 3390 855 3396 856
rect 3606 860 3612 861
rect 3606 856 3607 860
rect 3611 856 3612 860
rect 3606 855 3612 856
rect 3822 860 3828 861
rect 3822 856 3823 860
rect 3827 856 3828 860
rect 3822 855 3828 856
rect 3942 857 3948 858
rect 2046 852 2052 853
rect 3942 853 3943 857
rect 3947 853 3948 857
rect 3942 852 3948 853
rect 322 851 328 852
rect 322 847 323 851
rect 327 847 328 851
rect 322 846 328 847
rect 514 851 520 852
rect 514 847 515 851
rect 519 847 520 851
rect 514 846 520 847
rect 566 851 572 852
rect 566 847 567 851
rect 571 850 572 851
rect 770 851 776 852
rect 571 848 681 850
rect 571 847 572 848
rect 566 846 572 847
rect 770 847 771 851
rect 775 850 776 851
rect 943 851 949 852
rect 775 848 865 850
rect 775 847 776 848
rect 770 846 776 847
rect 943 847 944 851
rect 948 850 949 851
rect 1242 851 1248 852
rect 948 848 1041 850
rect 948 847 949 848
rect 943 846 949 847
rect 1242 847 1243 851
rect 1247 847 1248 851
rect 1242 846 1248 847
rect 1402 851 1408 852
rect 1402 847 1403 851
rect 1407 847 1408 851
rect 1402 846 1408 847
rect 1554 851 1560 852
rect 1554 847 1555 851
rect 1559 847 1560 851
rect 1554 846 1560 847
rect 1706 851 1712 852
rect 1706 847 1707 851
rect 1711 847 1712 851
rect 1706 846 1712 847
rect 1734 851 1740 852
rect 1734 847 1735 851
rect 1739 850 1740 851
rect 2335 851 2341 852
rect 1739 848 1825 850
rect 1739 847 1740 848
rect 1734 846 1740 847
rect 2335 847 2336 851
rect 2340 850 2341 851
rect 2430 851 2436 852
rect 2340 848 2385 850
rect 2340 847 2341 848
rect 2335 846 2341 847
rect 2430 847 2431 851
rect 2435 850 2436 851
rect 2526 851 2532 852
rect 2435 848 2481 850
rect 2435 847 2436 848
rect 2430 846 2436 847
rect 2526 847 2527 851
rect 2531 850 2532 851
rect 2706 851 2712 852
rect 2531 848 2577 850
rect 2531 847 2532 848
rect 2526 846 2532 847
rect 2706 847 2707 851
rect 2711 847 2712 851
rect 2706 846 2712 847
rect 2714 851 2720 852
rect 2714 847 2715 851
rect 2719 850 2720 851
rect 2938 851 2944 852
rect 2719 848 2777 850
rect 2719 847 2720 848
rect 2714 846 2720 847
rect 2938 847 2939 851
rect 2943 847 2944 851
rect 2938 846 2944 847
rect 3090 851 3096 852
rect 3090 847 3091 851
rect 3095 847 3096 851
rect 3090 846 3096 847
rect 3266 851 3272 852
rect 3266 847 3267 851
rect 3271 847 3272 851
rect 3266 846 3272 847
rect 3466 851 3472 852
rect 3466 847 3467 851
rect 3471 847 3472 851
rect 3466 846 3472 847
rect 3474 851 3480 852
rect 3474 847 3475 851
rect 3479 850 3480 851
rect 3890 851 3896 852
rect 3479 848 3649 850
rect 3479 847 3480 848
rect 3474 846 3480 847
rect 3890 847 3891 851
rect 3895 847 3896 851
rect 3890 846 3896 847
rect 254 841 260 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 254 837 255 841
rect 259 837 260 841
rect 254 836 260 837
rect 446 841 452 842
rect 446 837 447 841
rect 451 837 452 841
rect 446 836 452 837
rect 638 841 644 842
rect 638 837 639 841
rect 643 837 644 841
rect 638 836 644 837
rect 822 841 828 842
rect 822 837 823 841
rect 827 837 828 841
rect 822 836 828 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1166 841 1172 842
rect 1166 837 1167 841
rect 1171 837 1172 841
rect 1166 836 1172 837
rect 1326 841 1332 842
rect 1326 837 1327 841
rect 1331 837 1332 841
rect 1326 836 1332 837
rect 1478 841 1484 842
rect 1478 837 1479 841
rect 1483 837 1484 841
rect 1478 836 1484 837
rect 1630 841 1636 842
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1782 841 1788 842
rect 2342 841 2348 842
rect 1782 837 1783 841
rect 1787 837 1788 841
rect 1782 836 1788 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 110 835 116 836
rect 2006 835 2012 836
rect 2046 840 2052 841
rect 2046 836 2047 840
rect 2051 836 2052 840
rect 2342 837 2343 841
rect 2347 837 2348 841
rect 2342 836 2348 837
rect 2438 841 2444 842
rect 2438 837 2439 841
rect 2443 837 2444 841
rect 2438 836 2444 837
rect 2534 841 2540 842
rect 2534 837 2535 841
rect 2539 837 2540 841
rect 2534 836 2540 837
rect 2630 841 2636 842
rect 2630 837 2631 841
rect 2635 837 2636 841
rect 2630 836 2636 837
rect 2734 841 2740 842
rect 2734 837 2735 841
rect 2739 837 2740 841
rect 2734 836 2740 837
rect 2862 841 2868 842
rect 2862 837 2863 841
rect 2867 837 2868 841
rect 2862 836 2868 837
rect 3014 841 3020 842
rect 3014 837 3015 841
rect 3019 837 3020 841
rect 3014 836 3020 837
rect 3190 841 3196 842
rect 3190 837 3191 841
rect 3195 837 3196 841
rect 3190 836 3196 837
rect 3390 841 3396 842
rect 3390 837 3391 841
rect 3395 837 3396 841
rect 3390 836 3396 837
rect 3606 841 3612 842
rect 3606 837 3607 841
rect 3611 837 3612 841
rect 3606 836 3612 837
rect 3822 841 3828 842
rect 3822 837 3823 841
rect 3827 837 3828 841
rect 3822 836 3828 837
rect 3942 840 3948 841
rect 3942 836 3943 840
rect 3947 836 3948 840
rect 2046 835 2052 836
rect 3942 835 3948 836
rect 2714 831 2720 832
rect 2714 830 2715 831
rect 2660 828 2715 830
rect 483 823 489 824
rect 234 819 240 820
rect 234 815 235 819
rect 239 818 240 819
rect 291 819 297 820
rect 291 818 292 819
rect 239 816 292 818
rect 239 815 240 816
rect 234 814 240 815
rect 291 815 292 816
rect 296 815 297 819
rect 483 819 484 823
rect 488 822 489 823
rect 566 823 572 824
rect 566 822 567 823
rect 488 820 567 822
rect 488 819 489 820
rect 483 818 489 819
rect 566 819 567 820
rect 571 819 572 823
rect 566 818 572 819
rect 675 823 681 824
rect 675 819 676 823
rect 680 822 681 823
rect 770 823 776 824
rect 770 822 771 823
rect 680 820 771 822
rect 680 819 681 820
rect 675 818 681 819
rect 770 819 771 820
rect 775 819 776 823
rect 770 818 776 819
rect 859 823 865 824
rect 859 819 860 823
rect 864 822 865 823
rect 943 823 949 824
rect 943 822 944 823
rect 864 820 944 822
rect 864 819 865 820
rect 859 818 865 819
rect 943 819 944 820
rect 948 819 949 823
rect 943 818 949 819
rect 1035 823 1041 824
rect 1035 819 1036 823
rect 1040 822 1041 823
rect 1050 823 1056 824
rect 1050 822 1051 823
rect 1040 820 1051 822
rect 1040 819 1041 820
rect 1035 818 1041 819
rect 1050 819 1051 820
rect 1055 819 1056 823
rect 1242 823 1248 824
rect 1050 818 1056 819
rect 1203 819 1209 820
rect 291 814 297 815
rect 1203 815 1204 819
rect 1208 818 1209 819
rect 1242 819 1243 823
rect 1247 822 1248 823
rect 1363 823 1369 824
rect 1363 822 1364 823
rect 1247 820 1364 822
rect 1247 819 1248 820
rect 1242 818 1248 819
rect 1363 819 1364 820
rect 1368 819 1369 823
rect 1363 818 1369 819
rect 1402 823 1408 824
rect 1402 819 1403 823
rect 1407 822 1408 823
rect 1515 823 1521 824
rect 1515 822 1516 823
rect 1407 820 1516 822
rect 1407 819 1408 820
rect 1402 818 1408 819
rect 1515 819 1516 820
rect 1520 819 1521 823
rect 1515 818 1521 819
rect 1554 823 1560 824
rect 1554 819 1555 823
rect 1559 822 1560 823
rect 1667 823 1673 824
rect 1667 822 1668 823
rect 1559 820 1668 822
rect 1559 819 1560 820
rect 1554 818 1560 819
rect 1667 819 1668 820
rect 1672 819 1673 823
rect 1667 818 1673 819
rect 1706 823 1712 824
rect 1706 819 1707 823
rect 1711 822 1712 823
rect 1819 823 1825 824
rect 1819 822 1820 823
rect 1711 820 1820 822
rect 1711 819 1712 820
rect 1706 818 1712 819
rect 1819 819 1820 820
rect 1824 819 1825 823
rect 1819 818 1825 819
rect 2379 823 2385 824
rect 2379 819 2380 823
rect 2384 822 2385 823
rect 2430 823 2436 824
rect 2430 822 2431 823
rect 2384 820 2431 822
rect 2384 819 2385 820
rect 2379 818 2385 819
rect 2430 819 2431 820
rect 2435 819 2436 823
rect 2430 818 2436 819
rect 2475 823 2481 824
rect 2475 819 2476 823
rect 2480 822 2481 823
rect 2526 823 2532 824
rect 2526 822 2527 823
rect 2480 820 2527 822
rect 2480 819 2481 820
rect 2475 818 2481 819
rect 2526 819 2527 820
rect 2531 819 2532 823
rect 2526 818 2532 819
rect 2571 823 2577 824
rect 2571 819 2572 823
rect 2576 822 2577 823
rect 2660 822 2662 828
rect 2714 827 2715 828
rect 2719 827 2720 831
rect 3410 831 3416 832
rect 3410 830 3411 831
rect 2714 826 2720 827
rect 2932 828 3411 830
rect 2576 820 2662 822
rect 2667 823 2673 824
rect 2576 819 2577 820
rect 2571 818 2577 819
rect 2667 819 2668 823
rect 2672 822 2673 823
rect 2690 823 2696 824
rect 2690 822 2691 823
rect 2672 820 2691 822
rect 2672 819 2673 820
rect 2667 818 2673 819
rect 2690 819 2691 820
rect 2695 819 2696 823
rect 2690 818 2696 819
rect 2706 823 2712 824
rect 2706 819 2707 823
rect 2711 822 2712 823
rect 2771 823 2777 824
rect 2771 822 2772 823
rect 2711 820 2772 822
rect 2711 819 2712 820
rect 2706 818 2712 819
rect 2771 819 2772 820
rect 2776 819 2777 823
rect 2771 818 2777 819
rect 2899 823 2905 824
rect 2899 819 2900 823
rect 2904 822 2905 823
rect 2932 822 2934 828
rect 3410 827 3411 828
rect 3415 827 3416 831
rect 3410 826 3416 827
rect 2904 820 2934 822
rect 2938 823 2944 824
rect 2904 819 2905 820
rect 2899 818 2905 819
rect 2938 819 2939 823
rect 2943 822 2944 823
rect 3051 823 3057 824
rect 3051 822 3052 823
rect 2943 820 3052 822
rect 2943 819 2944 820
rect 2938 818 2944 819
rect 3051 819 3052 820
rect 3056 819 3057 823
rect 3051 818 3057 819
rect 3090 823 3096 824
rect 3090 819 3091 823
rect 3095 822 3096 823
rect 3227 823 3233 824
rect 3227 822 3228 823
rect 3095 820 3228 822
rect 3095 819 3096 820
rect 3090 818 3096 819
rect 3227 819 3228 820
rect 3232 819 3233 823
rect 3227 818 3233 819
rect 3266 823 3272 824
rect 3266 819 3267 823
rect 3271 822 3272 823
rect 3427 823 3433 824
rect 3427 822 3428 823
rect 3271 820 3428 822
rect 3271 819 3272 820
rect 3266 818 3272 819
rect 3427 819 3428 820
rect 3432 819 3433 823
rect 3427 818 3433 819
rect 3466 823 3472 824
rect 3466 819 3467 823
rect 3471 822 3472 823
rect 3643 823 3649 824
rect 3643 822 3644 823
rect 3471 820 3644 822
rect 3471 819 3472 820
rect 3466 818 3472 819
rect 3643 819 3644 820
rect 3648 819 3649 823
rect 3643 818 3649 819
rect 3859 823 3865 824
rect 3859 819 3860 823
rect 3864 822 3865 823
rect 3914 823 3920 824
rect 3914 822 3915 823
rect 3864 820 3915 822
rect 3864 819 3865 820
rect 3859 818 3865 819
rect 3914 819 3915 820
rect 3919 819 3920 823
rect 3914 818 3920 819
rect 1208 816 1238 818
rect 1208 815 1209 816
rect 1203 814 1209 815
rect 1236 814 1238 816
rect 1518 815 1524 816
rect 1518 814 1519 815
rect 1236 812 1519 814
rect 1518 811 1519 812
rect 1523 811 1524 815
rect 3474 815 3480 816
rect 3474 814 3475 815
rect 1518 810 1524 811
rect 2916 812 3475 814
rect 2916 810 2918 812
rect 3474 811 3475 812
rect 3479 811 3480 815
rect 3474 810 3480 811
rect 2915 809 2921 810
rect 2335 807 2341 808
rect 195 803 201 804
rect 195 799 196 803
rect 200 802 201 803
rect 255 803 261 804
rect 255 802 256 803
rect 200 800 256 802
rect 200 799 201 800
rect 195 798 201 799
rect 255 799 256 800
rect 260 799 261 803
rect 255 798 261 799
rect 338 803 344 804
rect 338 799 339 803
rect 343 802 344 803
rect 347 803 353 804
rect 347 802 348 803
rect 343 800 348 802
rect 343 799 344 800
rect 338 798 344 799
rect 347 799 348 800
rect 352 799 353 803
rect 347 798 353 799
rect 507 803 516 804
rect 507 799 508 803
rect 515 799 516 803
rect 507 798 516 799
rect 546 803 552 804
rect 546 799 547 803
rect 551 802 552 803
rect 659 803 665 804
rect 659 802 660 803
rect 551 800 660 802
rect 551 799 552 800
rect 546 798 552 799
rect 659 799 660 800
rect 664 799 665 803
rect 659 798 665 799
rect 698 803 704 804
rect 698 799 699 803
rect 703 802 704 803
rect 811 803 817 804
rect 811 802 812 803
rect 703 800 812 802
rect 703 799 704 800
rect 698 798 704 799
rect 811 799 812 800
rect 816 799 817 803
rect 811 798 817 799
rect 971 803 980 804
rect 971 799 972 803
rect 979 799 980 803
rect 971 798 980 799
rect 1010 803 1016 804
rect 1010 799 1011 803
rect 1015 802 1016 803
rect 1131 803 1137 804
rect 1131 802 1132 803
rect 1015 800 1132 802
rect 1015 799 1016 800
rect 1010 798 1016 799
rect 1131 799 1132 800
rect 1136 799 1137 803
rect 1131 798 1137 799
rect 1230 803 1236 804
rect 1230 799 1231 803
rect 1235 802 1236 803
rect 1291 803 1297 804
rect 1291 802 1292 803
rect 1235 800 1292 802
rect 1235 799 1236 800
rect 1230 798 1236 799
rect 1291 799 1292 800
rect 1296 799 1297 803
rect 1291 798 1297 799
rect 1374 803 1380 804
rect 1374 799 1375 803
rect 1379 802 1380 803
rect 1451 803 1457 804
rect 1451 802 1452 803
rect 1379 800 1452 802
rect 1379 799 1380 800
rect 1374 798 1380 799
rect 1451 799 1452 800
rect 1456 799 1457 803
rect 1451 798 1457 799
rect 1490 803 1496 804
rect 1490 799 1491 803
rect 1495 802 1496 803
rect 1619 803 1625 804
rect 1619 802 1620 803
rect 1495 800 1620 802
rect 1495 799 1496 800
rect 1490 798 1496 799
rect 1619 799 1620 800
rect 1624 799 1625 803
rect 1619 798 1625 799
rect 1787 803 1793 804
rect 1787 799 1788 803
rect 1792 802 1793 803
rect 1834 803 1840 804
rect 1834 802 1835 803
rect 1792 800 1835 802
rect 1792 799 1793 800
rect 1787 798 1793 799
rect 1834 799 1835 800
rect 1839 799 1840 803
rect 1834 798 1840 799
rect 1939 803 1945 804
rect 1939 799 1940 803
rect 1944 802 1945 803
rect 1986 803 1992 804
rect 1986 802 1987 803
rect 1944 800 1987 802
rect 1944 799 1945 800
rect 1939 798 1945 799
rect 1986 799 1987 800
rect 1991 799 1992 803
rect 2335 803 2336 807
rect 2340 806 2341 807
rect 2347 807 2353 808
rect 2347 806 2348 807
rect 2340 804 2348 806
rect 2340 803 2341 804
rect 2335 802 2341 803
rect 2347 803 2348 804
rect 2352 803 2353 807
rect 2347 802 2353 803
rect 2386 807 2392 808
rect 2386 803 2387 807
rect 2391 806 2392 807
rect 2531 807 2537 808
rect 2531 806 2532 807
rect 2391 804 2532 806
rect 2391 803 2392 804
rect 2386 802 2392 803
rect 2531 803 2532 804
rect 2536 803 2537 807
rect 2531 802 2537 803
rect 2570 807 2576 808
rect 2570 803 2571 807
rect 2575 806 2576 807
rect 2723 807 2729 808
rect 2723 806 2724 807
rect 2575 804 2724 806
rect 2575 803 2576 804
rect 2570 802 2576 803
rect 2723 803 2724 804
rect 2728 803 2729 807
rect 2915 805 2916 809
rect 2920 805 2921 809
rect 2915 804 2921 805
rect 2954 807 2960 808
rect 2723 802 2729 803
rect 2954 803 2955 807
rect 2959 806 2960 807
rect 3115 807 3121 808
rect 3115 806 3116 807
rect 2959 804 3116 806
rect 2959 803 2960 804
rect 2954 802 2960 803
rect 3115 803 3116 804
rect 3120 803 3121 807
rect 3115 802 3121 803
rect 3154 807 3160 808
rect 3154 803 3155 807
rect 3159 806 3160 807
rect 3323 807 3329 808
rect 3323 806 3324 807
rect 3159 804 3324 806
rect 3159 803 3160 804
rect 3154 802 3160 803
rect 3323 803 3324 804
rect 3328 803 3329 807
rect 3323 802 3329 803
rect 3362 807 3368 808
rect 3362 803 3363 807
rect 3367 806 3368 807
rect 3539 807 3545 808
rect 3539 806 3540 807
rect 3367 804 3540 806
rect 3367 803 3368 804
rect 3362 802 3368 803
rect 3539 803 3540 804
rect 3544 803 3545 807
rect 3539 802 3545 803
rect 3755 807 3761 808
rect 3755 803 3756 807
rect 3760 806 3761 807
rect 3770 807 3776 808
rect 3770 806 3771 807
rect 3760 804 3771 806
rect 3760 803 3761 804
rect 3755 802 3761 803
rect 3770 803 3771 804
rect 3775 803 3776 807
rect 3770 802 3776 803
rect 1986 798 1992 799
rect 2046 788 2052 789
rect 3942 788 3948 789
rect 110 784 116 785
rect 2006 784 2012 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 158 783 164 784
rect 158 779 159 783
rect 163 779 164 783
rect 158 778 164 779
rect 310 783 316 784
rect 310 779 311 783
rect 315 779 316 783
rect 310 778 316 779
rect 470 783 476 784
rect 470 779 471 783
rect 475 779 476 783
rect 470 778 476 779
rect 622 783 628 784
rect 622 779 623 783
rect 627 779 628 783
rect 622 778 628 779
rect 774 783 780 784
rect 774 779 775 783
rect 779 779 780 783
rect 774 778 780 779
rect 934 783 940 784
rect 934 779 935 783
rect 939 779 940 783
rect 934 778 940 779
rect 1094 783 1100 784
rect 1094 779 1095 783
rect 1099 779 1100 783
rect 1094 778 1100 779
rect 1254 783 1260 784
rect 1254 779 1255 783
rect 1259 779 1260 783
rect 1254 778 1260 779
rect 1414 783 1420 784
rect 1414 779 1415 783
rect 1419 779 1420 783
rect 1414 778 1420 779
rect 1582 783 1588 784
rect 1582 779 1583 783
rect 1587 779 1588 783
rect 1582 778 1588 779
rect 1750 783 1756 784
rect 1750 779 1751 783
rect 1755 779 1756 783
rect 1750 778 1756 779
rect 1902 783 1908 784
rect 1902 779 1903 783
rect 1907 779 1908 783
rect 2006 780 2007 784
rect 2011 780 2012 784
rect 2046 784 2047 788
rect 2051 784 2052 788
rect 2046 783 2052 784
rect 2310 787 2316 788
rect 2310 783 2311 787
rect 2315 783 2316 787
rect 2310 782 2316 783
rect 2494 787 2500 788
rect 2494 783 2495 787
rect 2499 783 2500 787
rect 2494 782 2500 783
rect 2686 787 2692 788
rect 2686 783 2687 787
rect 2691 783 2692 787
rect 2686 782 2692 783
rect 2878 787 2884 788
rect 2878 783 2879 787
rect 2883 783 2884 787
rect 2878 782 2884 783
rect 3078 787 3084 788
rect 3078 783 3079 787
rect 3083 783 3084 787
rect 3078 782 3084 783
rect 3286 787 3292 788
rect 3286 783 3287 787
rect 3291 783 3292 787
rect 3286 782 3292 783
rect 3502 787 3508 788
rect 3502 783 3503 787
rect 3507 783 3508 787
rect 3502 782 3508 783
rect 3718 787 3724 788
rect 3718 783 3719 787
rect 3723 783 3724 787
rect 3942 784 3943 788
rect 3947 784 3948 788
rect 3942 783 3948 784
rect 3718 782 3724 783
rect 2006 779 2012 780
rect 2386 779 2392 780
rect 1902 778 1908 779
rect 234 775 240 776
rect 234 771 235 775
rect 239 771 240 775
rect 234 770 240 771
rect 255 775 261 776
rect 255 771 256 775
rect 260 774 261 775
rect 546 775 552 776
rect 260 772 353 774
rect 260 771 261 772
rect 255 770 261 771
rect 546 771 547 775
rect 551 771 552 775
rect 546 770 552 771
rect 698 775 704 776
rect 698 771 699 775
rect 703 771 704 775
rect 1010 775 1016 776
rect 698 770 704 771
rect 850 771 856 772
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 850 767 851 771
rect 855 767 856 771
rect 1010 771 1011 775
rect 1015 771 1016 775
rect 1230 775 1236 776
rect 1230 774 1231 775
rect 1173 772 1231 774
rect 1010 770 1016 771
rect 1230 771 1231 772
rect 1235 771 1236 775
rect 1374 775 1380 776
rect 1374 774 1375 775
rect 1333 772 1375 774
rect 1230 770 1236 771
rect 1374 771 1375 772
rect 1379 771 1380 775
rect 1374 770 1380 771
rect 1490 775 1496 776
rect 1490 771 1491 775
rect 1495 771 1496 775
rect 1490 770 1496 771
rect 1518 775 1524 776
rect 1518 771 1519 775
rect 1523 774 1524 775
rect 1834 775 1840 776
rect 1523 772 1625 774
rect 1523 771 1524 772
rect 1518 770 1524 771
rect 1826 771 1832 772
rect 850 766 856 767
rect 1826 767 1827 771
rect 1831 767 1832 771
rect 1834 771 1835 775
rect 1839 774 1840 775
rect 2386 775 2387 779
rect 2391 775 2392 779
rect 2386 774 2392 775
rect 2570 779 2576 780
rect 2570 775 2571 779
rect 2575 775 2576 779
rect 2570 774 2576 775
rect 2679 779 2685 780
rect 2679 775 2680 779
rect 2684 778 2685 779
rect 2954 779 2960 780
rect 2684 776 2729 778
rect 2684 775 2685 776
rect 2679 774 2685 775
rect 2954 775 2955 779
rect 2959 775 2960 779
rect 2954 774 2960 775
rect 3154 779 3160 780
rect 3154 775 3155 779
rect 3159 775 3160 779
rect 3154 774 3160 775
rect 3362 779 3368 780
rect 3362 775 3363 779
rect 3367 775 3368 779
rect 3362 774 3368 775
rect 3446 779 3452 780
rect 3446 775 3447 779
rect 3451 778 3452 779
rect 3686 779 3692 780
rect 3451 776 3545 778
rect 3451 775 3452 776
rect 3446 774 3452 775
rect 3686 775 3687 779
rect 3691 778 3692 779
rect 3691 776 3761 778
rect 3691 775 3692 776
rect 3686 774 3692 775
rect 1839 772 1945 774
rect 1839 771 1840 772
rect 1834 770 1840 771
rect 2046 771 2052 772
rect 1826 766 1832 767
rect 2006 767 2012 768
rect 110 762 116 763
rect 158 764 164 765
rect 158 760 159 764
rect 163 760 164 764
rect 158 759 164 760
rect 310 764 316 765
rect 310 760 311 764
rect 315 760 316 764
rect 310 759 316 760
rect 470 764 476 765
rect 470 760 471 764
rect 475 760 476 764
rect 470 759 476 760
rect 622 764 628 765
rect 622 760 623 764
rect 627 760 628 764
rect 622 759 628 760
rect 774 764 780 765
rect 774 760 775 764
rect 779 760 780 764
rect 774 759 780 760
rect 934 764 940 765
rect 934 760 935 764
rect 939 760 940 764
rect 934 759 940 760
rect 1094 764 1100 765
rect 1094 760 1095 764
rect 1099 760 1100 764
rect 1094 759 1100 760
rect 1254 764 1260 765
rect 1254 760 1255 764
rect 1259 760 1260 764
rect 1254 759 1260 760
rect 1414 764 1420 765
rect 1414 760 1415 764
rect 1419 760 1420 764
rect 1414 759 1420 760
rect 1582 764 1588 765
rect 1582 760 1583 764
rect 1587 760 1588 764
rect 1582 759 1588 760
rect 1750 764 1756 765
rect 1750 760 1751 764
rect 1755 760 1756 764
rect 1750 759 1756 760
rect 1902 764 1908 765
rect 1902 760 1903 764
rect 1907 760 1908 764
rect 2006 763 2007 767
rect 2011 763 2012 767
rect 2046 767 2047 771
rect 2051 767 2052 771
rect 3942 771 3948 772
rect 2046 766 2052 767
rect 2310 768 2316 769
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2494 768 2500 769
rect 2494 764 2495 768
rect 2499 764 2500 768
rect 2494 763 2500 764
rect 2686 768 2692 769
rect 2686 764 2687 768
rect 2691 764 2692 768
rect 2686 763 2692 764
rect 2878 768 2884 769
rect 2878 764 2879 768
rect 2883 764 2884 768
rect 2878 763 2884 764
rect 3078 768 3084 769
rect 3078 764 3079 768
rect 3083 764 3084 768
rect 3078 763 3084 764
rect 3286 768 3292 769
rect 3286 764 3287 768
rect 3291 764 3292 768
rect 3286 763 3292 764
rect 3502 768 3508 769
rect 3502 764 3503 768
rect 3507 764 3508 768
rect 3502 763 3508 764
rect 3718 768 3724 769
rect 3718 764 3719 768
rect 3723 764 3724 768
rect 3942 767 3943 771
rect 3947 767 3948 771
rect 3942 766 3948 767
rect 3718 763 3724 764
rect 2006 762 2012 763
rect 1902 759 1908 760
rect 134 704 140 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 134 700 135 704
rect 139 700 140 704
rect 134 699 140 700
rect 262 704 268 705
rect 262 700 263 704
rect 267 700 268 704
rect 262 699 268 700
rect 430 704 436 705
rect 430 700 431 704
rect 435 700 436 704
rect 430 699 436 700
rect 622 704 628 705
rect 622 700 623 704
rect 627 700 628 704
rect 622 699 628 700
rect 822 704 828 705
rect 822 700 823 704
rect 827 700 828 704
rect 822 699 828 700
rect 1014 704 1020 705
rect 1014 700 1015 704
rect 1019 700 1020 704
rect 1014 699 1020 700
rect 1206 704 1212 705
rect 1206 700 1207 704
rect 1211 700 1212 704
rect 1206 699 1212 700
rect 1390 704 1396 705
rect 1390 700 1391 704
rect 1395 700 1396 704
rect 1390 699 1396 700
rect 1566 704 1572 705
rect 1566 700 1567 704
rect 1571 700 1572 704
rect 1566 699 1572 700
rect 1742 704 1748 705
rect 1742 700 1743 704
rect 1747 700 1748 704
rect 1742 699 1748 700
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2070 704 2076 705
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2046 701 2052 702
rect 2046 697 2047 701
rect 2051 697 2052 701
rect 2070 700 2071 704
rect 2075 700 2076 704
rect 2070 699 2076 700
rect 2254 704 2260 705
rect 2254 700 2255 704
rect 2259 700 2260 704
rect 2254 699 2260 700
rect 2454 704 2460 705
rect 2454 700 2455 704
rect 2459 700 2460 704
rect 2454 699 2460 700
rect 2654 704 2660 705
rect 2654 700 2655 704
rect 2659 700 2660 704
rect 2654 699 2660 700
rect 2854 704 2860 705
rect 2854 700 2855 704
rect 2859 700 2860 704
rect 2854 699 2860 700
rect 3046 704 3052 705
rect 3046 700 3047 704
rect 3051 700 3052 704
rect 3046 699 3052 700
rect 3238 704 3244 705
rect 3238 700 3239 704
rect 3243 700 3244 704
rect 3238 699 3244 700
rect 3438 704 3444 705
rect 3438 700 3439 704
rect 3443 700 3444 704
rect 3438 699 3444 700
rect 3638 704 3644 705
rect 3638 700 3639 704
rect 3643 700 3644 704
rect 3638 699 3644 700
rect 3838 704 3844 705
rect 3838 700 3839 704
rect 3843 700 3844 704
rect 3838 699 3844 700
rect 3942 701 3948 702
rect 2046 696 2052 697
rect 3942 697 3943 701
rect 3947 697 3948 701
rect 3942 696 3948 697
rect 210 695 216 696
rect 210 691 211 695
rect 215 691 216 695
rect 210 690 216 691
rect 338 695 344 696
rect 338 691 339 695
rect 343 691 344 695
rect 338 690 344 691
rect 422 695 428 696
rect 422 691 423 695
rect 427 694 428 695
rect 542 695 548 696
rect 427 692 473 694
rect 427 691 428 692
rect 422 690 428 691
rect 542 691 543 695
rect 547 694 548 695
rect 706 695 712 696
rect 547 692 665 694
rect 547 691 548 692
rect 542 690 548 691
rect 706 691 707 695
rect 711 694 712 695
rect 974 695 980 696
rect 711 692 865 694
rect 711 691 712 692
rect 706 690 712 691
rect 974 691 975 695
rect 979 694 980 695
rect 1103 695 1109 696
rect 979 692 1057 694
rect 979 691 980 692
rect 974 690 980 691
rect 1103 691 1104 695
rect 1108 694 1109 695
rect 1466 695 1472 696
rect 1108 692 1249 694
rect 1108 691 1109 692
rect 1103 690 1109 691
rect 1466 691 1467 695
rect 1471 691 1472 695
rect 1466 690 1472 691
rect 1642 695 1648 696
rect 1642 691 1643 695
rect 1647 691 1648 695
rect 1642 690 1648 691
rect 1650 695 1656 696
rect 1650 691 1651 695
rect 1655 694 1656 695
rect 1986 695 1992 696
rect 1655 692 1785 694
rect 1828 692 1945 694
rect 1655 691 1656 692
rect 1650 690 1656 691
rect 1810 687 1816 688
rect 134 685 140 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 134 681 135 685
rect 139 681 140 685
rect 134 680 140 681
rect 262 685 268 686
rect 262 681 263 685
rect 267 681 268 685
rect 262 680 268 681
rect 430 685 436 686
rect 430 681 431 685
rect 435 681 436 685
rect 430 680 436 681
rect 622 685 628 686
rect 622 681 623 685
rect 627 681 628 685
rect 622 680 628 681
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 1014 685 1020 686
rect 1014 681 1015 685
rect 1019 681 1020 685
rect 1014 680 1020 681
rect 1206 685 1212 686
rect 1206 681 1207 685
rect 1211 681 1212 685
rect 1206 680 1212 681
rect 1390 685 1396 686
rect 1390 681 1391 685
rect 1395 681 1396 685
rect 1390 680 1396 681
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 1742 685 1748 686
rect 1742 681 1743 685
rect 1747 681 1748 685
rect 1810 683 1811 687
rect 1815 686 1816 687
rect 1828 686 1830 692
rect 1986 691 1987 695
rect 1991 694 1992 695
rect 2199 695 2205 696
rect 1991 692 2113 694
rect 1991 691 1992 692
rect 1986 690 1992 691
rect 2199 691 2200 695
rect 2204 694 2205 695
rect 2338 695 2344 696
rect 2204 692 2297 694
rect 2204 691 2205 692
rect 2199 690 2205 691
rect 2338 691 2339 695
rect 2343 694 2344 695
rect 2730 695 2736 696
rect 2343 692 2497 694
rect 2343 691 2344 692
rect 2338 690 2344 691
rect 2730 691 2731 695
rect 2735 691 2736 695
rect 2730 690 2736 691
rect 2930 695 2936 696
rect 2930 691 2931 695
rect 2935 691 2936 695
rect 2930 690 2936 691
rect 3122 695 3128 696
rect 3122 691 3123 695
rect 3127 691 3128 695
rect 3122 690 3128 691
rect 3314 695 3320 696
rect 3314 691 3315 695
rect 3319 691 3320 695
rect 3314 690 3320 691
rect 3514 695 3520 696
rect 3514 691 3515 695
rect 3519 691 3520 695
rect 3514 690 3520 691
rect 3558 695 3564 696
rect 3558 691 3559 695
rect 3563 694 3564 695
rect 3906 695 3912 696
rect 3563 692 3681 694
rect 3563 691 3564 692
rect 3558 690 3564 691
rect 3906 691 3907 695
rect 3911 691 3912 695
rect 3906 690 3912 691
rect 1815 684 1830 686
rect 1902 685 1908 686
rect 2070 685 2076 686
rect 1815 683 1816 684
rect 1810 682 1816 683
rect 1742 680 1748 681
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 2006 679 2012 680
rect 2046 684 2052 685
rect 2046 680 2047 684
rect 2051 680 2052 684
rect 2070 681 2071 685
rect 2075 681 2076 685
rect 2070 680 2076 681
rect 2254 685 2260 686
rect 2254 681 2255 685
rect 2259 681 2260 685
rect 2254 680 2260 681
rect 2454 685 2460 686
rect 2454 681 2455 685
rect 2459 681 2460 685
rect 2454 680 2460 681
rect 2654 685 2660 686
rect 2654 681 2655 685
rect 2659 681 2660 685
rect 2654 680 2660 681
rect 2854 685 2860 686
rect 2854 681 2855 685
rect 2859 681 2860 685
rect 2854 680 2860 681
rect 3046 685 3052 686
rect 3046 681 3047 685
rect 3051 681 3052 685
rect 3046 680 3052 681
rect 3238 685 3244 686
rect 3238 681 3239 685
rect 3243 681 3244 685
rect 3238 680 3244 681
rect 3438 685 3444 686
rect 3438 681 3439 685
rect 3443 681 3444 685
rect 3438 680 3444 681
rect 3638 685 3644 686
rect 3638 681 3639 685
rect 3643 681 3644 685
rect 3638 680 3644 681
rect 3838 685 3844 686
rect 3838 681 3839 685
rect 3843 681 3844 685
rect 3838 680 3844 681
rect 3942 684 3948 685
rect 3942 680 3943 684
rect 3947 680 3948 684
rect 2046 679 2052 680
rect 3942 679 3948 680
rect 1650 675 1656 676
rect 1650 674 1651 675
rect 1460 672 1651 674
rect 210 667 216 668
rect 171 663 177 664
rect 171 659 172 663
rect 176 662 177 663
rect 210 663 211 667
rect 215 666 216 667
rect 299 667 305 668
rect 299 666 300 667
rect 215 664 300 666
rect 215 663 216 664
rect 210 662 216 663
rect 299 663 300 664
rect 304 663 305 667
rect 299 662 305 663
rect 467 667 473 668
rect 467 663 468 667
rect 472 666 473 667
rect 542 667 548 668
rect 542 666 543 667
rect 472 664 543 666
rect 472 663 473 664
rect 467 662 473 663
rect 542 663 543 664
rect 547 663 548 667
rect 542 662 548 663
rect 659 667 665 668
rect 659 663 660 667
rect 664 666 665 667
rect 706 667 712 668
rect 706 666 707 667
rect 664 664 707 666
rect 664 663 665 664
rect 659 662 665 663
rect 706 663 707 664
rect 711 663 712 667
rect 706 662 712 663
rect 850 667 856 668
rect 850 663 851 667
rect 855 666 856 667
rect 859 667 865 668
rect 859 666 860 667
rect 855 664 860 666
rect 855 663 856 664
rect 850 662 856 663
rect 859 663 860 664
rect 864 663 865 667
rect 859 662 865 663
rect 1051 667 1057 668
rect 1051 663 1052 667
rect 1056 666 1057 667
rect 1103 667 1109 668
rect 1103 666 1104 667
rect 1056 664 1104 666
rect 1056 663 1057 664
rect 1051 662 1057 663
rect 1103 663 1104 664
rect 1108 663 1109 667
rect 1427 667 1433 668
rect 1103 662 1109 663
rect 1243 663 1249 664
rect 176 659 178 662
rect 171 658 178 659
rect 210 659 216 660
rect 210 658 211 659
rect 176 656 211 658
rect 210 655 211 656
rect 215 655 216 659
rect 1243 659 1244 663
rect 1248 662 1249 663
rect 1391 663 1397 664
rect 1391 662 1392 663
rect 1248 660 1392 662
rect 1248 659 1249 660
rect 1243 658 1249 659
rect 1391 659 1392 660
rect 1396 659 1397 663
rect 1427 663 1428 667
rect 1432 666 1433 667
rect 1460 666 1462 672
rect 1650 671 1651 672
rect 1655 671 1656 675
rect 3446 675 3452 676
rect 3446 674 3447 675
rect 1650 670 1656 671
rect 2924 672 3447 674
rect 1432 664 1462 666
rect 1466 667 1472 668
rect 1432 663 1433 664
rect 1427 662 1433 663
rect 1466 663 1467 667
rect 1471 666 1472 667
rect 1603 667 1609 668
rect 1603 666 1604 667
rect 1471 664 1604 666
rect 1471 663 1472 664
rect 1466 662 1472 663
rect 1603 663 1604 664
rect 1608 663 1609 667
rect 1603 662 1609 663
rect 1779 667 1785 668
rect 1779 663 1780 667
rect 1784 666 1785 667
rect 1810 667 1816 668
rect 1810 666 1811 667
rect 1784 664 1811 666
rect 1784 663 1785 664
rect 1779 662 1785 663
rect 1810 663 1811 664
rect 1815 663 1816 667
rect 1810 662 1816 663
rect 1826 667 1832 668
rect 1826 663 1827 667
rect 1831 666 1832 667
rect 1939 667 1945 668
rect 1939 666 1940 667
rect 1831 664 1940 666
rect 1831 663 1832 664
rect 1826 662 1832 663
rect 1939 663 1940 664
rect 1944 663 1945 667
rect 1939 662 1945 663
rect 2107 667 2113 668
rect 2107 663 2108 667
rect 2112 666 2113 667
rect 2199 667 2205 668
rect 2199 666 2200 667
rect 2112 664 2200 666
rect 2112 663 2113 664
rect 2107 662 2113 663
rect 2199 663 2200 664
rect 2204 663 2205 667
rect 2199 662 2205 663
rect 2291 667 2297 668
rect 2291 663 2292 667
rect 2296 666 2297 667
rect 2338 667 2344 668
rect 2338 666 2339 667
rect 2296 664 2339 666
rect 2296 663 2297 664
rect 2291 662 2297 663
rect 2338 663 2339 664
rect 2343 663 2344 667
rect 2679 667 2685 668
rect 2338 662 2344 663
rect 2491 663 2497 664
rect 1391 658 1397 659
rect 2491 659 2492 663
rect 2496 662 2497 663
rect 2506 663 2512 664
rect 2506 662 2507 663
rect 2496 660 2507 662
rect 2496 659 2497 660
rect 2491 658 2497 659
rect 2506 659 2507 660
rect 2511 659 2512 663
rect 2679 663 2680 667
rect 2684 666 2685 667
rect 2691 667 2697 668
rect 2691 666 2692 667
rect 2684 664 2692 666
rect 2684 663 2685 664
rect 2679 662 2685 663
rect 2691 663 2692 664
rect 2696 663 2697 667
rect 2691 662 2697 663
rect 2891 667 2897 668
rect 2891 663 2892 667
rect 2896 666 2897 667
rect 2924 666 2926 672
rect 3446 671 3447 672
rect 3451 671 3452 675
rect 3446 670 3452 671
rect 2896 664 2926 666
rect 2930 667 2936 668
rect 2896 663 2897 664
rect 2891 662 2897 663
rect 2930 663 2931 667
rect 2935 666 2936 667
rect 3083 667 3089 668
rect 3083 666 3084 667
rect 2935 664 3084 666
rect 2935 663 2936 664
rect 2930 662 2936 663
rect 3083 663 3084 664
rect 3088 663 3089 667
rect 3083 662 3089 663
rect 3122 667 3128 668
rect 3122 663 3123 667
rect 3127 666 3128 667
rect 3275 667 3281 668
rect 3275 666 3276 667
rect 3127 664 3276 666
rect 3127 663 3128 664
rect 3122 662 3128 663
rect 3275 663 3276 664
rect 3280 663 3281 667
rect 3275 662 3281 663
rect 3314 667 3320 668
rect 3314 663 3315 667
rect 3319 666 3320 667
rect 3475 667 3481 668
rect 3475 666 3476 667
rect 3319 664 3476 666
rect 3319 663 3320 664
rect 3314 662 3320 663
rect 3475 663 3476 664
rect 3480 663 3481 667
rect 3475 662 3481 663
rect 3514 667 3520 668
rect 3514 663 3515 667
rect 3519 666 3520 667
rect 3675 667 3681 668
rect 3675 666 3676 667
rect 3519 664 3676 666
rect 3519 663 3520 664
rect 3514 662 3520 663
rect 3675 663 3676 664
rect 3680 663 3681 667
rect 3675 662 3681 663
rect 3875 667 3881 668
rect 3875 663 3876 667
rect 3880 666 3881 667
rect 3890 667 3896 668
rect 3890 666 3891 667
rect 3880 664 3891 666
rect 3880 663 3881 664
rect 3875 662 3881 663
rect 3890 663 3891 664
rect 3895 663 3896 667
rect 3890 662 3896 663
rect 2506 658 2512 659
rect 3558 659 3564 660
rect 3558 658 3559 659
rect 210 654 216 655
rect 3060 656 3559 658
rect 3060 654 3062 656
rect 3558 655 3559 656
rect 3563 655 3564 659
rect 3558 654 3564 655
rect 3059 653 3065 654
rect 171 651 177 652
rect 171 647 172 651
rect 176 650 177 651
rect 218 651 224 652
rect 218 650 219 651
rect 176 648 219 650
rect 176 647 177 648
rect 171 646 177 647
rect 218 647 219 648
rect 223 647 224 651
rect 218 646 224 647
rect 283 651 292 652
rect 283 647 284 651
rect 291 647 292 651
rect 283 646 292 647
rect 419 651 428 652
rect 419 647 420 651
rect 427 647 428 651
rect 419 646 428 647
rect 458 651 464 652
rect 458 647 459 651
rect 463 650 464 651
rect 563 651 569 652
rect 563 650 564 651
rect 463 648 564 650
rect 463 647 464 648
rect 458 646 464 647
rect 563 647 564 648
rect 568 647 569 651
rect 563 646 569 647
rect 602 651 608 652
rect 602 647 603 651
rect 607 650 608 651
rect 723 651 729 652
rect 723 650 724 651
rect 607 648 724 650
rect 607 647 608 648
rect 602 646 608 647
rect 723 647 724 648
rect 728 647 729 651
rect 723 646 729 647
rect 907 651 916 652
rect 907 647 908 651
rect 915 647 916 651
rect 907 646 916 647
rect 946 651 952 652
rect 946 647 947 651
rect 951 650 952 651
rect 1115 651 1121 652
rect 1115 650 1116 651
rect 951 648 1116 650
rect 951 647 952 648
rect 946 646 952 647
rect 1115 647 1116 648
rect 1120 647 1121 651
rect 1115 646 1121 647
rect 1154 651 1160 652
rect 1154 647 1155 651
rect 1159 650 1160 651
rect 1339 651 1345 652
rect 1339 650 1340 651
rect 1159 648 1340 650
rect 1159 647 1160 648
rect 1154 646 1160 647
rect 1339 647 1340 648
rect 1344 647 1345 651
rect 1339 646 1345 647
rect 1378 651 1384 652
rect 1378 647 1379 651
rect 1383 650 1384 651
rect 1579 651 1585 652
rect 1579 650 1580 651
rect 1383 648 1580 650
rect 1383 647 1384 648
rect 1378 646 1384 647
rect 1579 647 1580 648
rect 1584 647 1585 651
rect 1579 646 1585 647
rect 1642 651 1648 652
rect 1642 647 1643 651
rect 1647 650 1648 651
rect 1819 651 1825 652
rect 1819 650 1820 651
rect 1647 648 1820 650
rect 1647 647 1648 648
rect 1642 646 1648 647
rect 1819 647 1820 648
rect 1824 647 1825 651
rect 1819 646 1825 647
rect 2107 651 2116 652
rect 2107 647 2108 651
rect 2115 647 2116 651
rect 2107 646 2116 647
rect 2146 651 2152 652
rect 2146 647 2147 651
rect 2151 650 2152 651
rect 2267 651 2273 652
rect 2267 650 2268 651
rect 2151 648 2268 650
rect 2151 647 2152 648
rect 2146 646 2152 647
rect 2267 647 2268 648
rect 2272 647 2273 651
rect 2267 646 2273 647
rect 2306 651 2312 652
rect 2306 647 2307 651
rect 2311 650 2312 651
rect 2467 651 2473 652
rect 2467 650 2468 651
rect 2311 648 2468 650
rect 2311 647 2312 648
rect 2306 646 2312 647
rect 2467 647 2468 648
rect 2472 647 2473 651
rect 2467 646 2473 647
rect 2667 651 2673 652
rect 2667 647 2668 651
rect 2672 650 2673 651
rect 2722 651 2728 652
rect 2722 650 2723 651
rect 2672 648 2723 650
rect 2672 647 2673 648
rect 2667 646 2673 647
rect 2722 647 2723 648
rect 2727 647 2728 651
rect 2722 646 2728 647
rect 2730 651 2736 652
rect 2730 647 2731 651
rect 2735 650 2736 651
rect 2867 651 2873 652
rect 2867 650 2868 651
rect 2735 648 2868 650
rect 2735 647 2736 648
rect 2730 646 2736 647
rect 2867 647 2868 648
rect 2872 647 2873 651
rect 3059 649 3060 653
rect 3064 649 3065 653
rect 3059 648 3065 649
rect 3098 651 3104 652
rect 2867 646 2873 647
rect 3098 647 3099 651
rect 3103 650 3104 651
rect 3243 651 3249 652
rect 3243 650 3244 651
rect 3103 648 3244 650
rect 3103 647 3104 648
rect 3098 646 3104 647
rect 3243 647 3244 648
rect 3248 647 3249 651
rect 3243 646 3249 647
rect 3282 651 3288 652
rect 3282 647 3283 651
rect 3287 650 3288 651
rect 3411 651 3417 652
rect 3411 650 3412 651
rect 3287 648 3412 650
rect 3287 647 3288 648
rect 3282 646 3288 647
rect 3411 647 3412 648
rect 3416 647 3417 651
rect 3411 646 3417 647
rect 3450 651 3456 652
rect 3450 647 3451 651
rect 3455 650 3456 651
rect 3571 651 3577 652
rect 3571 650 3572 651
rect 3455 648 3572 650
rect 3455 647 3456 648
rect 3450 646 3456 647
rect 3571 647 3572 648
rect 3576 647 3577 651
rect 3571 646 3577 647
rect 3731 651 3737 652
rect 3731 647 3732 651
rect 3736 650 3737 651
rect 3778 651 3784 652
rect 3778 650 3779 651
rect 3736 648 3779 650
rect 3736 647 3737 648
rect 3731 646 3737 647
rect 3778 647 3779 648
rect 3783 647 3784 651
rect 3778 646 3784 647
rect 3875 651 3881 652
rect 3875 647 3876 651
rect 3880 650 3881 651
rect 3906 651 3912 652
rect 3906 650 3907 651
rect 3880 648 3907 650
rect 3880 647 3881 648
rect 3875 646 3881 647
rect 3906 647 3907 648
rect 3911 647 3912 651
rect 3906 646 3912 647
rect 110 632 116 633
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 134 631 140 632
rect 134 627 135 631
rect 139 627 140 631
rect 134 626 140 627
rect 246 631 252 632
rect 246 627 247 631
rect 251 627 252 631
rect 246 626 252 627
rect 382 631 388 632
rect 382 627 383 631
rect 387 627 388 631
rect 382 626 388 627
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 870 631 876 632
rect 870 627 871 631
rect 875 627 876 631
rect 870 626 876 627
rect 1078 631 1084 632
rect 1078 627 1079 631
rect 1083 627 1084 631
rect 1078 626 1084 627
rect 1302 631 1308 632
rect 1302 627 1303 631
rect 1307 627 1308 631
rect 1302 626 1308 627
rect 1542 631 1548 632
rect 1542 627 1543 631
rect 1547 627 1548 631
rect 1542 626 1548 627
rect 1782 631 1788 632
rect 1782 627 1783 631
rect 1787 627 1788 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 632 2052 633
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2070 631 2076 632
rect 2070 627 2071 631
rect 2075 627 2076 631
rect 1782 626 1788 627
rect 2070 626 2076 627
rect 2230 631 2236 632
rect 2230 627 2231 631
rect 2235 627 2236 631
rect 2230 626 2236 627
rect 2430 631 2436 632
rect 2430 627 2431 631
rect 2435 627 2436 631
rect 2430 626 2436 627
rect 2630 631 2636 632
rect 2630 627 2631 631
rect 2635 627 2636 631
rect 2630 626 2636 627
rect 2830 631 2836 632
rect 2830 627 2831 631
rect 2835 627 2836 631
rect 2830 626 2836 627
rect 3022 631 3028 632
rect 3022 627 3023 631
rect 3027 627 3028 631
rect 3022 626 3028 627
rect 3206 631 3212 632
rect 3206 627 3207 631
rect 3211 627 3212 631
rect 3206 626 3212 627
rect 3374 631 3380 632
rect 3374 627 3375 631
rect 3379 627 3380 631
rect 3374 626 3380 627
rect 3534 631 3540 632
rect 3534 627 3535 631
rect 3539 627 3540 631
rect 3534 626 3540 627
rect 3694 631 3700 632
rect 3694 627 3695 631
rect 3699 627 3700 631
rect 3694 626 3700 627
rect 3838 631 3844 632
rect 3838 627 3839 631
rect 3843 627 3844 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3838 626 3844 627
rect 210 623 216 624
rect 210 619 211 623
rect 215 619 216 623
rect 210 618 216 619
rect 218 623 224 624
rect 218 619 219 623
rect 223 622 224 623
rect 458 623 464 624
rect 223 620 289 622
rect 223 619 224 620
rect 218 618 224 619
rect 458 619 459 623
rect 463 619 464 623
rect 458 618 464 619
rect 602 623 608 624
rect 602 619 603 623
rect 607 619 608 623
rect 946 623 952 624
rect 602 618 608 619
rect 762 619 768 620
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 762 615 763 619
rect 767 615 768 619
rect 946 619 947 623
rect 951 619 952 623
rect 946 618 952 619
rect 1154 623 1160 624
rect 1154 619 1155 623
rect 1159 619 1160 623
rect 1154 618 1160 619
rect 1378 623 1384 624
rect 1378 619 1379 623
rect 1383 619 1384 623
rect 1378 618 1384 619
rect 1391 623 1397 624
rect 1391 619 1392 623
rect 1396 622 1397 623
rect 2146 623 2152 624
rect 1396 620 1585 622
rect 1396 619 1397 620
rect 1391 618 1397 619
rect 2146 619 2147 623
rect 2151 619 2152 623
rect 2146 618 2152 619
rect 2306 623 2312 624
rect 2306 619 2307 623
rect 2311 619 2312 623
rect 2306 618 2312 619
rect 2506 623 2512 624
rect 2506 619 2507 623
rect 2511 619 2512 623
rect 2506 618 2512 619
rect 2598 623 2604 624
rect 2598 619 2599 623
rect 2603 622 2604 623
rect 2722 623 2728 624
rect 2603 620 2673 622
rect 2603 619 2604 620
rect 2598 618 2604 619
rect 2722 619 2723 623
rect 2727 622 2728 623
rect 3098 623 3104 624
rect 2727 620 2873 622
rect 2727 619 2728 620
rect 2722 618 2728 619
rect 3098 619 3099 623
rect 3103 619 3104 623
rect 3098 618 3104 619
rect 3282 623 3288 624
rect 3282 619 3283 623
rect 3287 619 3288 623
rect 3282 618 3288 619
rect 3450 623 3456 624
rect 3450 619 3451 623
rect 3455 619 3456 623
rect 3770 623 3776 624
rect 3450 618 3456 619
rect 3610 619 3616 620
rect 762 614 768 615
rect 1850 615 1856 616
rect 110 610 116 611
rect 134 612 140 613
rect 134 608 135 612
rect 139 608 140 612
rect 134 607 140 608
rect 246 612 252 613
rect 246 608 247 612
rect 251 608 252 612
rect 246 607 252 608
rect 382 612 388 613
rect 382 608 383 612
rect 387 608 388 612
rect 382 607 388 608
rect 526 612 532 613
rect 526 608 527 612
rect 531 608 532 612
rect 526 607 532 608
rect 686 612 692 613
rect 686 608 687 612
rect 691 608 692 612
rect 686 607 692 608
rect 870 612 876 613
rect 870 608 871 612
rect 875 608 876 612
rect 870 607 876 608
rect 1078 612 1084 613
rect 1078 608 1079 612
rect 1083 608 1084 612
rect 1078 607 1084 608
rect 1302 612 1308 613
rect 1302 608 1303 612
rect 1307 608 1308 612
rect 1302 607 1308 608
rect 1542 612 1548 613
rect 1542 608 1543 612
rect 1547 608 1548 612
rect 1542 607 1548 608
rect 1782 612 1788 613
rect 1782 608 1783 612
rect 1787 608 1788 612
rect 1850 611 1851 615
rect 1855 614 1856 615
rect 1860 614 1862 617
rect 1855 612 1862 614
rect 2006 615 2012 616
rect 1855 611 1856 612
rect 1850 610 1856 611
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 615 2052 616
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 3610 615 3611 619
rect 3615 615 3616 619
rect 3770 619 3771 623
rect 3775 619 3776 623
rect 3770 618 3776 619
rect 3914 619 3920 620
rect 3610 614 3616 615
rect 3914 615 3915 619
rect 3919 615 3920 619
rect 3914 614 3920 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2070 612 2076 613
rect 1782 607 1788 608
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 2230 612 2236 613
rect 2230 608 2231 612
rect 2235 608 2236 612
rect 2230 607 2236 608
rect 2430 612 2436 613
rect 2430 608 2431 612
rect 2435 608 2436 612
rect 2430 607 2436 608
rect 2630 612 2636 613
rect 2630 608 2631 612
rect 2635 608 2636 612
rect 2630 607 2636 608
rect 2830 612 2836 613
rect 2830 608 2831 612
rect 2835 608 2836 612
rect 2830 607 2836 608
rect 3022 612 3028 613
rect 3022 608 3023 612
rect 3027 608 3028 612
rect 3022 607 3028 608
rect 3206 612 3212 613
rect 3206 608 3207 612
rect 3211 608 3212 612
rect 3206 607 3212 608
rect 3374 612 3380 613
rect 3374 608 3375 612
rect 3379 608 3380 612
rect 3374 607 3380 608
rect 3534 612 3540 613
rect 3534 608 3535 612
rect 3539 608 3540 612
rect 3534 607 3540 608
rect 3694 612 3700 613
rect 3694 608 3695 612
rect 3699 608 3700 612
rect 3694 607 3700 608
rect 3838 612 3844 613
rect 3838 608 3839 612
rect 3843 608 3844 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3838 607 3844 608
rect 2110 555 2116 556
rect 2110 551 2111 555
rect 2115 554 2116 555
rect 2115 552 2302 554
rect 2115 551 2116 552
rect 2110 550 2116 551
rect 134 548 140 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 134 544 135 548
rect 139 544 140 548
rect 134 543 140 544
rect 294 548 300 549
rect 294 544 295 548
rect 299 544 300 548
rect 294 543 300 544
rect 478 548 484 549
rect 478 544 479 548
rect 483 544 484 548
rect 478 543 484 544
rect 662 548 668 549
rect 662 544 663 548
rect 667 544 668 548
rect 662 543 668 544
rect 846 548 852 549
rect 846 544 847 548
rect 851 544 852 548
rect 846 543 852 544
rect 1030 548 1036 549
rect 1030 544 1031 548
rect 1035 544 1036 548
rect 1030 543 1036 544
rect 1214 548 1220 549
rect 1214 544 1215 548
rect 1219 544 1220 548
rect 1214 543 1220 544
rect 1398 548 1404 549
rect 1398 544 1399 548
rect 1403 544 1404 548
rect 1398 543 1404 544
rect 1590 548 1596 549
rect 1590 544 1591 548
rect 1595 544 1596 548
rect 1590 543 1596 544
rect 1782 548 1788 549
rect 1782 544 1783 548
rect 1787 544 1788 548
rect 2070 548 2076 549
rect 1782 543 1788 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2214 548 2220 549
rect 2214 544 2215 548
rect 2219 544 2220 548
rect 2214 543 2220 544
rect 2046 540 2052 541
rect 230 539 236 540
rect 230 538 231 539
rect 213 536 231 538
rect 230 535 231 536
rect 235 535 236 539
rect 230 534 236 535
rect 286 539 292 540
rect 286 535 287 539
rect 291 538 292 539
rect 471 539 477 540
rect 291 536 337 538
rect 291 535 292 536
rect 286 534 292 535
rect 471 535 472 539
rect 476 538 477 539
rect 575 539 581 540
rect 476 536 521 538
rect 476 535 477 536
rect 471 534 477 535
rect 575 535 576 539
rect 580 538 581 539
rect 914 539 920 540
rect 580 536 705 538
rect 580 535 581 536
rect 575 534 581 535
rect 914 535 915 539
rect 919 535 920 539
rect 914 534 920 535
rect 1106 539 1112 540
rect 1106 535 1107 539
rect 1111 535 1112 539
rect 1106 534 1112 535
rect 1114 539 1120 540
rect 1114 535 1115 539
rect 1119 538 1120 539
rect 1466 539 1472 540
rect 1119 536 1257 538
rect 1119 535 1120 536
rect 1114 534 1120 535
rect 1466 535 1467 539
rect 1471 535 1472 539
rect 1466 534 1472 535
rect 1519 539 1525 540
rect 1519 535 1520 539
rect 1524 538 1525 539
rect 1726 539 1732 540
rect 1524 536 1633 538
rect 1524 535 1525 536
rect 1519 534 1525 535
rect 1726 535 1727 539
rect 1731 538 1732 539
rect 2138 539 2144 540
rect 1731 536 1825 538
rect 1731 535 1732 536
rect 1726 534 1732 535
rect 2138 535 2139 539
rect 2143 535 2144 539
rect 2138 534 2144 535
rect 2183 539 2189 540
rect 2183 535 2184 539
rect 2188 538 2189 539
rect 2300 538 2302 552
rect 2398 548 2404 549
rect 2398 544 2399 548
rect 2403 544 2404 548
rect 2398 543 2404 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2774 548 2780 549
rect 2774 544 2775 548
rect 2779 544 2780 548
rect 2774 543 2780 544
rect 2958 548 2964 549
rect 2958 544 2959 548
rect 2963 544 2964 548
rect 2958 543 2964 544
rect 3142 548 3148 549
rect 3142 544 3143 548
rect 3147 544 3148 548
rect 3142 543 3148 544
rect 3318 548 3324 549
rect 3318 544 3319 548
rect 3323 544 3324 548
rect 3318 543 3324 544
rect 3494 548 3500 549
rect 3494 544 3495 548
rect 3499 544 3500 548
rect 3494 543 3500 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3678 543 3684 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 2530 539 2536 540
rect 2188 536 2257 538
rect 2300 536 2441 538
rect 2188 535 2189 536
rect 2183 534 2189 535
rect 2530 535 2531 539
rect 2535 538 2536 539
rect 2695 539 2701 540
rect 2535 536 2625 538
rect 2535 535 2536 536
rect 2530 534 2536 535
rect 2695 535 2696 539
rect 2700 538 2701 539
rect 3034 539 3040 540
rect 2700 536 2817 538
rect 2700 535 2701 536
rect 2695 534 2701 535
rect 3034 535 3035 539
rect 3039 535 3040 539
rect 3230 539 3236 540
rect 3230 538 3231 539
rect 3221 536 3231 538
rect 3034 534 3040 535
rect 3230 535 3231 536
rect 3235 535 3236 539
rect 3230 534 3236 535
rect 3238 539 3244 540
rect 3238 535 3239 539
rect 3243 538 3244 539
rect 3447 539 3453 540
rect 3243 536 3361 538
rect 3243 535 3244 536
rect 3238 534 3244 535
rect 3447 535 3448 539
rect 3452 538 3453 539
rect 3583 539 3589 540
rect 3452 536 3537 538
rect 3452 535 3453 536
rect 3447 534 3453 535
rect 3583 535 3584 539
rect 3588 538 3589 539
rect 3906 539 3912 540
rect 3588 536 3721 538
rect 3588 535 3589 536
rect 3583 534 3589 535
rect 3906 535 3907 539
rect 3911 535 3912 539
rect 3906 534 3912 535
rect 134 529 140 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 134 525 135 529
rect 139 525 140 529
rect 134 524 140 525
rect 294 529 300 530
rect 294 525 295 529
rect 299 525 300 529
rect 294 524 300 525
rect 478 529 484 530
rect 478 525 479 529
rect 483 525 484 529
rect 478 524 484 525
rect 662 529 668 530
rect 662 525 663 529
rect 667 525 668 529
rect 662 524 668 525
rect 846 529 852 530
rect 846 525 847 529
rect 851 525 852 529
rect 846 524 852 525
rect 1030 529 1036 530
rect 1030 525 1031 529
rect 1035 525 1036 529
rect 1030 524 1036 525
rect 1214 529 1220 530
rect 1214 525 1215 529
rect 1219 525 1220 529
rect 1214 524 1220 525
rect 1398 529 1404 530
rect 1398 525 1399 529
rect 1403 525 1404 529
rect 1398 524 1404 525
rect 1590 529 1596 530
rect 1590 525 1591 529
rect 1595 525 1596 529
rect 1590 524 1596 525
rect 1782 529 1788 530
rect 2070 529 2076 530
rect 1782 525 1783 529
rect 1787 525 1788 529
rect 1782 524 1788 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2214 529 2220 530
rect 2214 525 2215 529
rect 2219 525 2220 529
rect 2214 524 2220 525
rect 2398 529 2404 530
rect 2398 525 2399 529
rect 2403 525 2404 529
rect 2398 524 2404 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2774 529 2780 530
rect 2774 525 2775 529
rect 2779 525 2780 529
rect 2774 524 2780 525
rect 2958 529 2964 530
rect 2958 525 2959 529
rect 2963 525 2964 529
rect 2958 524 2964 525
rect 3142 529 3148 530
rect 3142 525 3143 529
rect 3147 525 3148 529
rect 3142 524 3148 525
rect 3318 529 3324 530
rect 3318 525 3319 529
rect 3323 525 3324 529
rect 3318 524 3324 525
rect 3494 529 3500 530
rect 3494 525 3495 529
rect 3499 525 3500 529
rect 3494 524 3500 525
rect 3678 529 3684 530
rect 3678 525 3679 529
rect 3683 525 3684 529
rect 3678 524 3684 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 1114 519 1120 520
rect 1114 518 1115 519
rect 972 516 1115 518
rect 230 511 236 512
rect 171 507 177 508
rect 171 503 172 507
rect 176 506 177 507
rect 210 507 216 508
rect 210 506 211 507
rect 176 504 211 506
rect 176 503 177 504
rect 171 502 177 503
rect 210 503 211 504
rect 215 503 216 507
rect 230 507 231 511
rect 235 510 236 511
rect 331 511 337 512
rect 331 510 332 511
rect 235 508 332 510
rect 235 507 236 508
rect 230 506 236 507
rect 331 507 332 508
rect 336 507 337 511
rect 331 506 337 507
rect 515 511 521 512
rect 515 507 516 511
rect 520 510 521 511
rect 575 511 581 512
rect 575 510 576 511
rect 520 508 576 510
rect 520 507 521 508
rect 515 506 521 507
rect 575 507 576 508
rect 580 507 581 511
rect 575 506 581 507
rect 699 511 705 512
rect 699 507 700 511
rect 704 510 705 511
rect 762 511 768 512
rect 762 510 763 511
rect 704 508 763 510
rect 704 507 705 508
rect 699 506 705 507
rect 762 507 763 508
rect 767 507 768 511
rect 762 506 768 507
rect 883 511 889 512
rect 883 507 884 511
rect 888 510 889 511
rect 972 510 974 516
rect 1114 515 1115 516
rect 1119 515 1120 519
rect 2598 519 2604 520
rect 2598 518 2599 519
rect 1114 514 1120 515
rect 2428 516 2599 518
rect 888 508 974 510
rect 1106 511 1112 512
rect 888 507 889 508
rect 883 506 889 507
rect 978 507 984 508
rect 210 502 216 503
rect 978 503 979 507
rect 983 506 984 507
rect 1067 507 1073 508
rect 1067 506 1068 507
rect 983 504 1068 506
rect 983 503 984 504
rect 978 502 984 503
rect 1067 503 1068 504
rect 1072 503 1073 507
rect 1106 507 1107 511
rect 1111 510 1112 511
rect 1251 511 1257 512
rect 1251 510 1252 511
rect 1111 508 1252 510
rect 1111 507 1112 508
rect 1106 506 1112 507
rect 1251 507 1252 508
rect 1256 507 1257 511
rect 1251 506 1257 507
rect 1435 511 1441 512
rect 1435 507 1436 511
rect 1440 510 1441 511
rect 1519 511 1525 512
rect 1519 510 1520 511
rect 1440 508 1520 510
rect 1440 507 1441 508
rect 1435 506 1441 507
rect 1519 507 1520 508
rect 1524 507 1525 511
rect 1519 506 1525 507
rect 1627 511 1633 512
rect 1627 507 1628 511
rect 1632 510 1633 511
rect 1726 511 1732 512
rect 1726 510 1727 511
rect 1632 508 1727 510
rect 1632 507 1633 508
rect 1627 506 1633 507
rect 1726 507 1727 508
rect 1731 507 1732 511
rect 1726 506 1732 507
rect 1819 511 1825 512
rect 1819 507 1820 511
rect 1824 510 1825 511
rect 1850 511 1856 512
rect 1850 510 1851 511
rect 1824 508 1851 510
rect 1824 507 1825 508
rect 1819 506 1825 507
rect 1850 507 1851 508
rect 1855 507 1856 511
rect 1850 506 1856 507
rect 2107 511 2113 512
rect 2107 507 2108 511
rect 2112 510 2113 511
rect 2183 511 2189 512
rect 2183 510 2184 511
rect 2112 508 2184 510
rect 2112 507 2113 508
rect 2107 506 2113 507
rect 2183 507 2184 508
rect 2188 507 2189 511
rect 2183 506 2189 507
rect 2251 511 2257 512
rect 2251 507 2252 511
rect 2256 510 2257 511
rect 2428 510 2430 516
rect 2598 515 2599 516
rect 2603 515 2604 519
rect 3238 519 3244 520
rect 3238 518 3239 519
rect 2598 514 2604 515
rect 3028 516 3239 518
rect 2256 508 2430 510
rect 2435 511 2441 512
rect 2256 507 2257 508
rect 2251 506 2257 507
rect 2435 507 2436 511
rect 2440 510 2441 511
rect 2530 511 2536 512
rect 2530 510 2531 511
rect 2440 508 2531 510
rect 2440 507 2441 508
rect 2435 506 2441 507
rect 2530 507 2531 508
rect 2535 507 2536 511
rect 2530 506 2536 507
rect 2619 511 2625 512
rect 2619 507 2620 511
rect 2624 510 2625 511
rect 2695 511 2701 512
rect 2695 510 2696 511
rect 2624 508 2696 510
rect 2624 507 2625 508
rect 2619 506 2625 507
rect 2695 507 2696 508
rect 2700 507 2701 511
rect 2995 511 3001 512
rect 2695 506 2701 507
rect 2802 507 2808 508
rect 1067 502 1073 503
rect 2802 503 2803 507
rect 2807 506 2808 507
rect 2811 507 2817 508
rect 2811 506 2812 507
rect 2807 504 2812 506
rect 2807 503 2808 504
rect 2802 502 2808 503
rect 2811 503 2812 504
rect 2816 503 2817 507
rect 2995 507 2996 511
rect 3000 510 3001 511
rect 3028 510 3030 516
rect 3238 515 3239 516
rect 3243 515 3244 519
rect 3238 514 3244 515
rect 3000 508 3030 510
rect 3034 511 3040 512
rect 3000 507 3001 508
rect 2995 506 3001 507
rect 3034 507 3035 511
rect 3039 510 3040 511
rect 3179 511 3185 512
rect 3179 510 3180 511
rect 3039 508 3180 510
rect 3039 507 3040 508
rect 3034 506 3040 507
rect 3179 507 3180 508
rect 3184 507 3185 511
rect 3179 506 3185 507
rect 3355 511 3361 512
rect 3355 507 3356 511
rect 3360 510 3361 511
rect 3447 511 3453 512
rect 3447 510 3448 511
rect 3360 508 3448 510
rect 3360 507 3361 508
rect 3355 506 3361 507
rect 3447 507 3448 508
rect 3452 507 3453 511
rect 3447 506 3453 507
rect 3531 511 3537 512
rect 3531 507 3532 511
rect 3536 510 3537 511
rect 3583 511 3589 512
rect 3583 510 3584 511
rect 3536 508 3584 510
rect 3536 507 3537 508
rect 3531 506 3537 507
rect 3583 507 3584 508
rect 3588 507 3589 511
rect 3583 506 3589 507
rect 3610 511 3616 512
rect 3610 507 3611 511
rect 3615 510 3616 511
rect 3715 511 3721 512
rect 3715 510 3716 511
rect 3615 508 3716 510
rect 3615 507 3616 508
rect 3610 506 3616 507
rect 3715 507 3716 508
rect 3720 507 3721 511
rect 3715 506 3721 507
rect 3875 511 3881 512
rect 3875 507 3876 511
rect 3880 510 3881 511
rect 3914 511 3920 512
rect 3914 510 3915 511
rect 3880 508 3915 510
rect 3880 507 3881 508
rect 3875 506 3881 507
rect 3914 507 3915 508
rect 3919 507 3920 511
rect 3914 506 3920 507
rect 2811 502 2817 503
rect 171 495 177 496
rect 171 491 172 495
rect 176 494 177 495
rect 246 495 252 496
rect 246 494 247 495
rect 176 492 247 494
rect 176 491 177 492
rect 171 490 177 491
rect 246 491 247 492
rect 251 491 252 495
rect 246 490 252 491
rect 323 495 329 496
rect 323 491 324 495
rect 328 494 329 495
rect 354 495 360 496
rect 354 494 355 495
rect 328 492 355 494
rect 328 491 329 492
rect 323 490 329 491
rect 354 491 355 492
rect 359 491 360 495
rect 354 490 360 491
rect 471 495 477 496
rect 471 491 472 495
rect 476 494 477 495
rect 491 495 497 496
rect 491 494 492 495
rect 476 492 492 494
rect 476 491 477 492
rect 471 490 477 491
rect 491 491 492 492
rect 496 491 497 495
rect 491 490 497 491
rect 530 495 536 496
rect 530 491 531 495
rect 535 494 536 495
rect 651 495 657 496
rect 651 494 652 495
rect 535 492 652 494
rect 535 491 536 492
rect 530 490 536 491
rect 651 491 652 492
rect 656 491 657 495
rect 651 490 657 491
rect 690 495 696 496
rect 690 491 691 495
rect 695 494 696 495
rect 803 495 809 496
rect 803 494 804 495
rect 695 492 804 494
rect 695 491 696 492
rect 690 490 696 491
rect 803 491 804 492
rect 808 491 809 495
rect 803 490 809 491
rect 939 495 945 496
rect 939 491 940 495
rect 944 494 945 495
rect 970 495 976 496
rect 970 494 971 495
rect 944 492 971 494
rect 944 491 945 492
rect 939 490 945 491
rect 970 491 971 492
rect 975 491 976 495
rect 1106 495 1112 496
rect 970 490 976 491
rect 1067 493 1073 494
rect 1067 489 1068 493
rect 1072 489 1073 493
rect 1106 491 1107 495
rect 1111 494 1112 495
rect 1195 495 1201 496
rect 1195 494 1196 495
rect 1111 492 1196 494
rect 1111 491 1112 492
rect 1106 490 1112 491
rect 1195 491 1196 492
rect 1200 491 1201 495
rect 1195 490 1201 491
rect 1234 495 1240 496
rect 1234 491 1235 495
rect 1239 494 1240 495
rect 1323 495 1329 496
rect 1323 494 1324 495
rect 1239 492 1324 494
rect 1239 491 1240 492
rect 1234 490 1240 491
rect 1323 491 1324 492
rect 1328 491 1329 495
rect 1323 490 1329 491
rect 1451 495 1457 496
rect 1451 491 1452 495
rect 1456 494 1457 495
rect 1466 495 1472 496
rect 1466 494 1467 495
rect 1456 492 1467 494
rect 1456 491 1457 492
rect 1451 490 1457 491
rect 1466 491 1467 492
rect 1471 491 1472 495
rect 1466 490 1472 491
rect 2107 491 2113 492
rect 1067 488 1073 489
rect 1068 486 1070 488
rect 1406 487 1412 488
rect 1406 486 1407 487
rect 1068 484 1407 486
rect 1406 483 1407 484
rect 1411 483 1412 487
rect 2107 487 2108 491
rect 2112 490 2113 491
rect 2138 491 2144 492
rect 2138 490 2139 491
rect 2112 488 2139 490
rect 2112 487 2113 488
rect 2107 486 2113 487
rect 2138 487 2139 488
rect 2143 487 2144 491
rect 2138 486 2144 487
rect 2259 491 2268 492
rect 2259 487 2260 491
rect 2267 487 2268 491
rect 2259 486 2268 487
rect 2298 491 2304 492
rect 2298 487 2299 491
rect 2303 490 2304 491
rect 2427 491 2433 492
rect 2427 490 2428 491
rect 2303 488 2428 490
rect 2303 487 2304 488
rect 2298 486 2304 487
rect 2427 487 2428 488
rect 2432 487 2433 491
rect 2427 486 2433 487
rect 2466 491 2472 492
rect 2466 487 2467 491
rect 2471 490 2472 491
rect 2595 491 2601 492
rect 2595 490 2596 491
rect 2471 488 2596 490
rect 2471 487 2472 488
rect 2466 486 2472 487
rect 2595 487 2596 488
rect 2600 487 2601 491
rect 2595 486 2601 487
rect 2634 491 2640 492
rect 2634 487 2635 491
rect 2639 490 2640 491
rect 2763 491 2769 492
rect 2763 490 2764 491
rect 2639 488 2764 490
rect 2639 487 2640 488
rect 2634 486 2640 487
rect 2763 487 2764 488
rect 2768 487 2769 491
rect 2763 486 2769 487
rect 2931 491 2937 492
rect 2931 487 2932 491
rect 2936 490 2937 491
rect 2978 491 2984 492
rect 2978 490 2979 491
rect 2936 488 2979 490
rect 2936 487 2937 488
rect 2931 486 2937 487
rect 2978 487 2979 488
rect 2983 487 2984 491
rect 2978 486 2984 487
rect 3099 491 3105 492
rect 3099 487 3100 491
rect 3104 490 3105 491
rect 3118 491 3124 492
rect 3118 490 3119 491
rect 3104 488 3119 490
rect 3104 487 3105 488
rect 3099 486 3105 487
rect 3118 487 3119 488
rect 3123 487 3124 491
rect 3118 486 3124 487
rect 3230 491 3236 492
rect 3230 487 3231 491
rect 3235 490 3236 491
rect 3259 491 3265 492
rect 3259 490 3260 491
rect 3235 488 3260 490
rect 3235 487 3236 488
rect 3230 486 3236 487
rect 3259 487 3260 488
rect 3264 487 3265 491
rect 3259 486 3265 487
rect 3298 491 3304 492
rect 3298 487 3299 491
rect 3303 490 3304 491
rect 3419 491 3425 492
rect 3419 490 3420 491
rect 3303 488 3420 490
rect 3303 487 3304 488
rect 3298 486 3304 487
rect 3419 487 3420 488
rect 3424 487 3425 491
rect 3618 491 3624 492
rect 3419 486 3425 487
rect 3579 489 3585 490
rect 3579 485 3580 489
rect 3584 485 3585 489
rect 3618 487 3619 491
rect 3623 490 3624 491
rect 3739 491 3745 492
rect 3739 490 3740 491
rect 3623 488 3740 490
rect 3623 487 3624 488
rect 3618 486 3624 487
rect 3739 487 3740 488
rect 3744 487 3745 491
rect 3739 486 3745 487
rect 3875 491 3881 492
rect 3875 487 3876 491
rect 3880 490 3881 491
rect 3906 491 3912 492
rect 3906 490 3907 491
rect 3880 488 3907 490
rect 3880 487 3881 488
rect 3875 486 3881 487
rect 3906 487 3907 488
rect 3911 487 3912 491
rect 3906 486 3912 487
rect 3579 484 3585 485
rect 1406 482 1412 483
rect 3580 482 3582 484
rect 3798 483 3804 484
rect 3798 482 3799 483
rect 3580 480 3799 482
rect 3798 479 3799 480
rect 3803 479 3804 483
rect 3798 478 3804 479
rect 110 476 116 477
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 454 475 460 476
rect 454 471 455 475
rect 459 471 460 475
rect 454 470 460 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 766 475 772 476
rect 766 471 767 475
rect 771 471 772 475
rect 766 470 772 471
rect 902 475 908 476
rect 902 471 903 475
rect 907 471 908 475
rect 902 470 908 471
rect 1030 475 1036 476
rect 1030 471 1031 475
rect 1035 471 1036 475
rect 1030 470 1036 471
rect 1158 475 1164 476
rect 1158 471 1159 475
rect 1163 471 1164 475
rect 1158 470 1164 471
rect 1286 475 1292 476
rect 1286 471 1287 475
rect 1291 471 1292 475
rect 1286 470 1292 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 472 2052 473
rect 3942 472 3948 473
rect 1414 470 1420 471
rect 2046 468 2047 472
rect 2051 468 2052 472
rect 210 467 216 468
rect 210 463 211 467
rect 215 463 216 467
rect 210 462 216 463
rect 246 467 252 468
rect 246 463 247 467
rect 251 466 252 467
rect 530 467 536 468
rect 251 464 329 466
rect 251 463 252 464
rect 246 462 252 463
rect 530 463 531 467
rect 535 463 536 467
rect 530 462 536 463
rect 690 467 696 468
rect 690 463 691 467
rect 695 463 696 467
rect 978 467 984 468
rect 690 462 696 463
rect 842 463 848 464
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 842 459 843 463
rect 847 459 848 463
rect 978 463 979 467
rect 983 463 984 467
rect 978 462 984 463
rect 1106 467 1112 468
rect 1106 463 1107 467
rect 1111 463 1112 467
rect 1106 462 1112 463
rect 1234 467 1240 468
rect 1234 463 1235 467
rect 1239 463 1240 467
rect 1406 467 1412 468
rect 2046 467 2052 468
rect 2070 471 2076 472
rect 2070 467 2071 471
rect 2075 467 2076 471
rect 1234 462 1240 463
rect 1398 463 1404 464
rect 1398 462 1399 463
rect 1365 460 1399 462
rect 842 458 848 459
rect 1398 459 1399 460
rect 1403 459 1404 463
rect 1406 463 1407 467
rect 1411 466 1412 467
rect 2070 466 2076 467
rect 2222 471 2228 472
rect 2222 467 2223 471
rect 2227 467 2228 471
rect 2222 466 2228 467
rect 2390 471 2396 472
rect 2390 467 2391 471
rect 2395 467 2396 471
rect 2390 466 2396 467
rect 2558 471 2564 472
rect 2558 467 2559 471
rect 2563 467 2564 471
rect 2558 466 2564 467
rect 2726 471 2732 472
rect 2726 467 2727 471
rect 2731 467 2732 471
rect 2726 466 2732 467
rect 2894 471 2900 472
rect 2894 467 2895 471
rect 2899 467 2900 471
rect 2894 466 2900 467
rect 3062 471 3068 472
rect 3062 467 3063 471
rect 3067 467 3068 471
rect 3062 466 3068 467
rect 3222 471 3228 472
rect 3222 467 3223 471
rect 3227 467 3228 471
rect 3222 466 3228 467
rect 3382 471 3388 472
rect 3382 467 3383 471
rect 3387 467 3388 471
rect 3382 466 3388 467
rect 3542 471 3548 472
rect 3542 467 3543 471
rect 3547 467 3548 471
rect 3542 466 3548 467
rect 3702 471 3708 472
rect 3702 467 3703 471
rect 3707 467 3708 471
rect 3702 466 3708 467
rect 3838 471 3844 472
rect 3838 467 3839 471
rect 3843 467 3844 471
rect 3942 468 3943 472
rect 3947 468 3948 472
rect 3942 467 3948 468
rect 3838 466 3844 467
rect 1411 464 1457 466
rect 1411 463 1412 464
rect 1406 462 1412 463
rect 2034 463 2040 464
rect 1398 458 1404 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 454 456 460 457
rect 454 452 455 456
rect 459 452 460 456
rect 454 451 460 452
rect 614 456 620 457
rect 614 452 615 456
rect 619 452 620 456
rect 614 451 620 452
rect 766 456 772 457
rect 766 452 767 456
rect 771 452 772 456
rect 766 451 772 452
rect 902 456 908 457
rect 902 452 903 456
rect 907 452 908 456
rect 902 451 908 452
rect 1030 456 1036 457
rect 1030 452 1031 456
rect 1035 452 1036 456
rect 1030 451 1036 452
rect 1158 456 1164 457
rect 1158 452 1159 456
rect 1163 452 1164 456
rect 1158 451 1164 452
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1286 451 1292 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2034 459 2035 463
rect 2039 462 2040 463
rect 2298 463 2304 464
rect 2039 460 2113 462
rect 2039 459 2040 460
rect 2034 458 2040 459
rect 2298 459 2299 463
rect 2303 459 2304 463
rect 2298 458 2304 459
rect 2466 463 2472 464
rect 2466 459 2467 463
rect 2471 459 2472 463
rect 2466 458 2472 459
rect 2634 463 2640 464
rect 2634 459 2635 463
rect 2639 459 2640 463
rect 2634 458 2640 459
rect 2802 463 2808 464
rect 2802 459 2803 463
rect 2807 459 2808 463
rect 2802 458 2808 459
rect 2886 463 2892 464
rect 2886 459 2887 463
rect 2891 462 2892 463
rect 2978 463 2984 464
rect 2891 460 2937 462
rect 2891 459 2892 460
rect 2886 458 2892 459
rect 2978 459 2979 463
rect 2983 462 2984 463
rect 3298 463 3304 464
rect 2983 460 3105 462
rect 2983 459 2984 460
rect 2978 458 2984 459
rect 3298 459 3299 463
rect 3303 459 3304 463
rect 3298 458 3304 459
rect 3318 463 3324 464
rect 3318 459 3319 463
rect 3323 462 3324 463
rect 3618 463 3624 464
rect 3323 460 3425 462
rect 3323 459 3324 460
rect 3318 458 3324 459
rect 3618 459 3619 463
rect 3623 459 3624 463
rect 3618 458 3624 459
rect 3778 463 3784 464
rect 3778 459 3779 463
rect 3783 459 3784 463
rect 3778 458 3784 459
rect 3798 463 3804 464
rect 3798 459 3799 463
rect 3803 462 3804 463
rect 3803 460 3881 462
rect 3803 459 3804 460
rect 3798 458 3804 459
rect 2006 454 2012 455
rect 2046 455 2052 456
rect 1414 451 1420 452
rect 2046 451 2047 455
rect 2051 451 2052 455
rect 3942 455 3948 456
rect 2046 450 2052 451
rect 2070 452 2076 453
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 2222 452 2228 453
rect 2222 448 2223 452
rect 2227 448 2228 452
rect 2222 447 2228 448
rect 2390 452 2396 453
rect 2390 448 2391 452
rect 2395 448 2396 452
rect 2390 447 2396 448
rect 2558 452 2564 453
rect 2558 448 2559 452
rect 2563 448 2564 452
rect 2558 447 2564 448
rect 2726 452 2732 453
rect 2726 448 2727 452
rect 2731 448 2732 452
rect 2726 447 2732 448
rect 2894 452 2900 453
rect 2894 448 2895 452
rect 2899 448 2900 452
rect 2894 447 2900 448
rect 3062 452 3068 453
rect 3062 448 3063 452
rect 3067 448 3068 452
rect 3062 447 3068 448
rect 3222 452 3228 453
rect 3222 448 3223 452
rect 3227 448 3228 452
rect 3222 447 3228 448
rect 3382 452 3388 453
rect 3382 448 3383 452
rect 3387 448 3388 452
rect 3382 447 3388 448
rect 3542 452 3548 453
rect 3542 448 3543 452
rect 3547 448 3548 452
rect 3542 447 3548 448
rect 3702 452 3708 453
rect 3702 448 3703 452
rect 3707 448 3708 452
rect 3702 447 3708 448
rect 3838 452 3844 453
rect 3838 448 3839 452
rect 3843 448 3844 452
rect 3942 451 3943 455
rect 3947 451 3948 455
rect 3942 450 3948 451
rect 3838 447 3844 448
rect 134 396 140 397
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 134 392 135 396
rect 139 392 140 396
rect 134 391 140 392
rect 286 396 292 397
rect 286 392 287 396
rect 291 392 292 396
rect 286 391 292 392
rect 446 396 452 397
rect 446 392 447 396
rect 451 392 452 396
rect 446 391 452 392
rect 598 396 604 397
rect 598 392 599 396
rect 603 392 604 396
rect 598 391 604 392
rect 750 396 756 397
rect 750 392 751 396
rect 755 392 756 396
rect 750 391 756 392
rect 902 396 908 397
rect 902 392 903 396
rect 907 392 908 396
rect 902 391 908 392
rect 1078 396 1084 397
rect 1078 392 1079 396
rect 1083 392 1084 396
rect 1078 391 1084 392
rect 1270 396 1276 397
rect 1270 392 1271 396
rect 1275 392 1276 396
rect 1270 391 1276 392
rect 1478 396 1484 397
rect 1478 392 1479 396
rect 1483 392 1484 396
rect 1478 391 1484 392
rect 1702 396 1708 397
rect 1702 392 1703 396
rect 1707 392 1708 396
rect 1702 391 1708 392
rect 1902 396 1908 397
rect 1902 392 1903 396
rect 1907 392 1908 396
rect 1902 391 1908 392
rect 2006 393 2012 394
rect 110 388 116 389
rect 2006 389 2007 393
rect 2011 389 2012 393
rect 2462 392 2468 393
rect 2006 388 2012 389
rect 2046 389 2052 390
rect 210 387 216 388
rect 210 383 211 387
rect 215 383 216 387
rect 210 382 216 383
rect 354 387 360 388
rect 354 383 355 387
rect 359 383 360 387
rect 354 382 360 383
rect 522 387 528 388
rect 522 383 523 387
rect 527 383 528 387
rect 522 382 528 383
rect 530 387 536 388
rect 530 383 531 387
rect 535 386 536 387
rect 682 387 688 388
rect 535 384 641 386
rect 535 383 536 384
rect 530 382 536 383
rect 682 383 683 387
rect 687 386 688 387
rect 970 387 976 388
rect 687 384 793 386
rect 687 383 688 384
rect 682 382 688 383
rect 970 383 971 387
rect 975 383 976 387
rect 970 382 976 383
rect 1031 387 1037 388
rect 1031 383 1032 387
rect 1036 386 1037 387
rect 1210 387 1216 388
rect 1036 384 1121 386
rect 1036 383 1037 384
rect 1031 382 1037 383
rect 1210 383 1211 387
rect 1215 386 1216 387
rect 1554 387 1560 388
rect 1215 384 1313 386
rect 1215 383 1216 384
rect 1210 382 1216 383
rect 1554 383 1555 387
rect 1559 383 1560 387
rect 1554 382 1560 383
rect 1638 387 1644 388
rect 1638 383 1639 387
rect 1643 386 1644 387
rect 1970 387 1976 388
rect 1643 384 1745 386
rect 1643 383 1644 384
rect 1638 382 1644 383
rect 1970 383 1971 387
rect 1975 383 1976 387
rect 2046 385 2047 389
rect 2051 385 2052 389
rect 2462 388 2463 392
rect 2467 388 2468 392
rect 2462 387 2468 388
rect 2558 392 2564 393
rect 2558 388 2559 392
rect 2563 388 2564 392
rect 2558 387 2564 388
rect 2654 392 2660 393
rect 2654 388 2655 392
rect 2659 388 2660 392
rect 2654 387 2660 388
rect 2750 392 2756 393
rect 2750 388 2751 392
rect 2755 388 2756 392
rect 2750 387 2756 388
rect 2846 392 2852 393
rect 2846 388 2847 392
rect 2851 388 2852 392
rect 2846 387 2852 388
rect 2942 392 2948 393
rect 2942 388 2943 392
rect 2947 388 2948 392
rect 2942 387 2948 388
rect 3038 392 3044 393
rect 3038 388 3039 392
rect 3043 388 3044 392
rect 3038 387 3044 388
rect 3134 392 3140 393
rect 3134 388 3135 392
rect 3139 388 3140 392
rect 3134 387 3140 388
rect 3230 392 3236 393
rect 3230 388 3231 392
rect 3235 388 3236 392
rect 3230 387 3236 388
rect 3942 389 3948 390
rect 2046 384 2052 385
rect 3942 385 3943 389
rect 3947 385 3948 389
rect 3942 384 3948 385
rect 1970 382 1976 383
rect 2262 383 2268 384
rect 2262 379 2263 383
rect 2267 382 2268 383
rect 2550 383 2556 384
rect 2267 380 2505 382
rect 2267 379 2268 380
rect 2262 378 2268 379
rect 2550 379 2551 383
rect 2555 382 2556 383
rect 2646 383 2652 384
rect 2555 380 2601 382
rect 2555 379 2556 380
rect 2550 378 2556 379
rect 2646 379 2647 383
rect 2651 382 2652 383
rect 2742 383 2748 384
rect 2651 380 2697 382
rect 2651 379 2652 380
rect 2646 378 2652 379
rect 2742 379 2743 383
rect 2747 382 2748 383
rect 2922 383 2928 384
rect 2747 380 2793 382
rect 2747 379 2748 380
rect 2742 378 2748 379
rect 2922 379 2923 383
rect 2927 379 2928 383
rect 2922 378 2928 379
rect 3018 383 3024 384
rect 3018 379 3019 383
rect 3023 379 3024 383
rect 3018 378 3024 379
rect 3114 383 3120 384
rect 3114 379 3115 383
rect 3119 379 3120 383
rect 3114 378 3120 379
rect 3210 383 3216 384
rect 3210 379 3211 383
rect 3215 379 3216 383
rect 3210 378 3216 379
rect 3298 383 3304 384
rect 3298 379 3299 383
rect 3303 379 3304 383
rect 3298 378 3304 379
rect 134 377 140 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 134 373 135 377
rect 139 373 140 377
rect 134 372 140 373
rect 286 377 292 378
rect 286 373 287 377
rect 291 373 292 377
rect 286 372 292 373
rect 446 377 452 378
rect 446 373 447 377
rect 451 373 452 377
rect 446 372 452 373
rect 598 377 604 378
rect 598 373 599 377
rect 603 373 604 377
rect 598 372 604 373
rect 750 377 756 378
rect 750 373 751 377
rect 755 373 756 377
rect 750 372 756 373
rect 902 377 908 378
rect 902 373 903 377
rect 907 373 908 377
rect 902 372 908 373
rect 1078 377 1084 378
rect 1078 373 1079 377
rect 1083 373 1084 377
rect 1078 372 1084 373
rect 1270 377 1276 378
rect 1270 373 1271 377
rect 1275 373 1276 377
rect 1270 372 1276 373
rect 1478 377 1484 378
rect 1478 373 1479 377
rect 1483 373 1484 377
rect 1478 372 1484 373
rect 1702 377 1708 378
rect 1702 373 1703 377
rect 1707 373 1708 377
rect 1702 372 1708 373
rect 1902 377 1908 378
rect 1902 373 1903 377
rect 1907 373 1908 377
rect 1902 372 1908 373
rect 2006 376 2012 377
rect 2006 372 2007 376
rect 2011 372 2012 376
rect 2462 373 2468 374
rect 110 371 116 372
rect 2006 371 2012 372
rect 2046 372 2052 373
rect 2046 368 2047 372
rect 2051 368 2052 372
rect 2462 369 2463 373
rect 2467 369 2468 373
rect 2462 368 2468 369
rect 2558 373 2564 374
rect 2558 369 2559 373
rect 2563 369 2564 373
rect 2558 368 2564 369
rect 2654 373 2660 374
rect 2654 369 2655 373
rect 2659 369 2660 373
rect 2654 368 2660 369
rect 2750 373 2756 374
rect 2750 369 2751 373
rect 2755 369 2756 373
rect 2750 368 2756 369
rect 2846 373 2852 374
rect 2846 369 2847 373
rect 2851 369 2852 373
rect 2846 368 2852 369
rect 2942 373 2948 374
rect 2942 369 2943 373
rect 2947 369 2948 373
rect 2942 368 2948 369
rect 3038 373 3044 374
rect 3038 369 3039 373
rect 3043 369 3044 373
rect 3038 368 3044 369
rect 3134 373 3140 374
rect 3134 369 3135 373
rect 3139 369 3140 373
rect 3134 368 3140 369
rect 3230 373 3236 374
rect 3230 369 3231 373
rect 3235 369 3236 373
rect 3230 368 3236 369
rect 3942 372 3948 373
rect 3942 368 3943 372
rect 3947 368 3948 372
rect 2046 367 2052 368
rect 3942 367 3948 368
rect 210 359 216 360
rect 151 355 157 356
rect 151 351 152 355
rect 156 354 157 355
rect 171 355 177 356
rect 171 354 172 355
rect 156 352 172 354
rect 156 351 157 352
rect 151 350 157 351
rect 171 351 172 352
rect 176 351 177 355
rect 210 355 211 359
rect 215 358 216 359
rect 323 359 329 360
rect 323 358 324 359
rect 215 356 324 358
rect 215 355 216 356
rect 210 354 216 355
rect 323 355 324 356
rect 328 355 329 359
rect 323 354 329 355
rect 483 359 489 360
rect 483 355 484 359
rect 488 358 489 359
rect 530 359 536 360
rect 530 358 531 359
rect 488 356 531 358
rect 488 355 489 356
rect 483 354 489 355
rect 530 355 531 356
rect 535 355 536 359
rect 530 354 536 355
rect 635 359 641 360
rect 635 355 636 359
rect 640 358 641 359
rect 682 359 688 360
rect 682 358 683 359
rect 640 356 683 358
rect 640 355 641 356
rect 635 354 641 355
rect 682 355 683 356
rect 687 355 688 359
rect 682 354 688 355
rect 787 359 793 360
rect 787 355 788 359
rect 792 358 793 359
rect 842 359 848 360
rect 842 358 843 359
rect 792 356 843 358
rect 792 355 793 356
rect 787 354 793 355
rect 842 355 843 356
rect 847 355 848 359
rect 842 354 848 355
rect 939 359 945 360
rect 939 355 940 359
rect 944 358 945 359
rect 1031 359 1037 360
rect 1031 358 1032 359
rect 944 356 1032 358
rect 944 355 945 356
rect 939 354 945 355
rect 1031 355 1032 356
rect 1036 355 1037 359
rect 1031 354 1037 355
rect 1115 359 1121 360
rect 1115 355 1116 359
rect 1120 358 1121 359
rect 1210 359 1216 360
rect 1210 358 1211 359
rect 1120 356 1211 358
rect 1120 355 1121 356
rect 1115 354 1121 355
rect 1210 355 1211 356
rect 1215 355 1216 359
rect 1398 359 1404 360
rect 1210 354 1216 355
rect 1234 355 1240 356
rect 171 350 177 351
rect 1234 351 1235 355
rect 1239 354 1240 355
rect 1307 355 1313 356
rect 1307 354 1308 355
rect 1239 352 1308 354
rect 1239 351 1240 352
rect 1234 350 1240 351
rect 1307 351 1308 352
rect 1312 351 1313 355
rect 1398 355 1399 359
rect 1403 358 1404 359
rect 1515 359 1521 360
rect 1515 358 1516 359
rect 1403 356 1516 358
rect 1403 355 1404 356
rect 1398 354 1404 355
rect 1515 355 1516 356
rect 1520 355 1521 359
rect 1515 354 1521 355
rect 1554 359 1560 360
rect 1554 355 1555 359
rect 1559 358 1560 359
rect 1739 359 1745 360
rect 1739 358 1740 359
rect 1559 356 1740 358
rect 1559 355 1560 356
rect 1554 354 1560 355
rect 1739 355 1740 356
rect 1744 355 1745 359
rect 1739 354 1745 355
rect 1939 359 1945 360
rect 1939 355 1940 359
rect 1944 358 1945 359
rect 2034 359 2040 360
rect 2034 358 2035 359
rect 1944 356 2035 358
rect 1944 355 1945 356
rect 1939 354 1945 355
rect 2034 355 2035 356
rect 2039 355 2040 359
rect 2034 354 2040 355
rect 2499 355 2505 356
rect 1307 350 1313 351
rect 2499 351 2500 355
rect 2504 354 2505 355
rect 2550 355 2556 356
rect 2550 354 2551 355
rect 2504 352 2551 354
rect 2504 351 2505 352
rect 2499 350 2505 351
rect 2550 351 2551 352
rect 2555 351 2556 355
rect 2550 350 2556 351
rect 2595 355 2601 356
rect 2595 351 2596 355
rect 2600 354 2601 355
rect 2646 355 2652 356
rect 2646 354 2647 355
rect 2600 352 2647 354
rect 2600 351 2601 352
rect 2595 350 2601 351
rect 2646 351 2647 352
rect 2651 351 2652 355
rect 2646 350 2652 351
rect 2691 355 2697 356
rect 2691 351 2692 355
rect 2696 354 2697 355
rect 2742 355 2748 356
rect 2742 354 2743 355
rect 2696 352 2743 354
rect 2696 351 2697 352
rect 2691 350 2697 351
rect 2742 351 2743 352
rect 2747 351 2748 355
rect 2883 355 2892 356
rect 2742 350 2748 351
rect 2787 351 2793 352
rect 1638 347 1644 348
rect 1638 346 1639 347
rect 1196 344 1639 346
rect 1196 342 1198 344
rect 1638 343 1639 344
rect 1643 343 1644 347
rect 2787 347 2788 351
rect 2792 350 2793 351
rect 2858 351 2864 352
rect 2858 350 2859 351
rect 2792 348 2859 350
rect 2792 347 2793 348
rect 2787 346 2793 347
rect 2858 347 2859 348
rect 2863 347 2864 351
rect 2883 351 2884 355
rect 2891 351 2892 355
rect 2883 350 2892 351
rect 2922 355 2928 356
rect 2922 351 2923 355
rect 2927 354 2928 355
rect 2979 355 2985 356
rect 2979 354 2980 355
rect 2927 352 2980 354
rect 2927 351 2928 352
rect 2922 350 2928 351
rect 2979 351 2980 352
rect 2984 351 2985 355
rect 2979 350 2985 351
rect 3018 355 3024 356
rect 3018 351 3019 355
rect 3023 354 3024 355
rect 3075 355 3081 356
rect 3075 354 3076 355
rect 3023 352 3076 354
rect 3023 351 3024 352
rect 3018 350 3024 351
rect 3075 351 3076 352
rect 3080 351 3081 355
rect 3075 350 3081 351
rect 3114 355 3120 356
rect 3114 351 3115 355
rect 3119 354 3120 355
rect 3171 355 3177 356
rect 3171 354 3172 355
rect 3119 352 3172 354
rect 3119 351 3120 352
rect 3114 350 3120 351
rect 3171 351 3172 352
rect 3176 351 3177 355
rect 3171 350 3177 351
rect 3210 355 3216 356
rect 3210 351 3211 355
rect 3215 354 3216 355
rect 3267 355 3273 356
rect 3267 354 3268 355
rect 3215 352 3268 354
rect 3215 351 3216 352
rect 3210 350 3216 351
rect 3267 351 3268 352
rect 3272 351 3273 355
rect 3267 350 3273 351
rect 2858 346 2864 347
rect 1638 342 1644 343
rect 1195 341 1201 342
rect 195 339 201 340
rect 195 335 196 339
rect 200 338 201 339
rect 242 339 248 340
rect 242 338 243 339
rect 200 336 243 338
rect 200 335 201 336
rect 195 334 201 335
rect 242 335 243 336
rect 247 335 248 339
rect 242 334 248 335
rect 375 339 381 340
rect 375 335 376 339
rect 380 338 381 339
rect 387 339 393 340
rect 387 338 388 339
rect 380 336 388 338
rect 380 335 381 336
rect 375 334 381 335
rect 387 335 388 336
rect 392 335 393 339
rect 387 334 393 335
rect 522 339 528 340
rect 522 335 523 339
rect 527 338 528 339
rect 587 339 593 340
rect 587 338 588 339
rect 527 336 588 338
rect 527 335 528 336
rect 522 334 528 335
rect 587 335 588 336
rect 592 335 593 339
rect 587 334 593 335
rect 626 339 632 340
rect 626 335 627 339
rect 631 338 632 339
rect 795 339 801 340
rect 795 338 796 339
rect 631 336 796 338
rect 631 335 632 336
rect 626 334 632 335
rect 795 335 796 336
rect 800 335 801 339
rect 795 334 801 335
rect 834 339 840 340
rect 834 335 835 339
rect 839 338 840 339
rect 995 339 1001 340
rect 995 338 996 339
rect 839 336 996 338
rect 839 335 840 336
rect 834 334 840 335
rect 995 335 996 336
rect 1000 335 1001 339
rect 1195 337 1196 341
rect 1200 337 1201 341
rect 1418 339 1424 340
rect 1195 336 1201 337
rect 1379 337 1385 338
rect 995 334 1001 335
rect 1379 333 1380 337
rect 1384 333 1385 337
rect 1418 335 1419 339
rect 1423 338 1424 339
rect 1563 339 1569 340
rect 1563 338 1564 339
rect 1423 336 1564 338
rect 1423 335 1424 336
rect 1418 334 1424 335
rect 1563 335 1564 336
rect 1568 335 1569 339
rect 1563 334 1569 335
rect 1602 339 1608 340
rect 1602 335 1603 339
rect 1607 338 1608 339
rect 1747 339 1753 340
rect 1747 338 1748 339
rect 1607 336 1748 338
rect 1607 335 1608 336
rect 1602 334 1608 335
rect 1747 335 1748 336
rect 1752 335 1753 339
rect 1747 334 1753 335
rect 1931 339 1937 340
rect 1931 335 1932 339
rect 1936 338 1937 339
rect 1970 339 1976 340
rect 1970 338 1971 339
rect 1936 336 1971 338
rect 1936 335 1937 336
rect 1931 334 1937 335
rect 1970 335 1971 336
rect 1975 335 1976 339
rect 1970 334 1976 335
rect 2435 339 2444 340
rect 2435 335 2436 339
rect 2443 335 2444 339
rect 2435 334 2444 335
rect 2474 339 2480 340
rect 2474 335 2475 339
rect 2479 338 2480 339
rect 2539 339 2545 340
rect 2539 338 2540 339
rect 2479 336 2540 338
rect 2479 335 2480 336
rect 2474 334 2480 335
rect 2539 335 2540 336
rect 2544 335 2545 339
rect 2539 334 2545 335
rect 2578 339 2584 340
rect 2578 335 2579 339
rect 2583 338 2584 339
rect 2659 339 2665 340
rect 2659 338 2660 339
rect 2583 336 2660 338
rect 2583 335 2584 336
rect 2578 334 2584 335
rect 2659 335 2660 336
rect 2664 335 2665 339
rect 2659 334 2665 335
rect 2698 339 2704 340
rect 2698 335 2699 339
rect 2703 338 2704 339
rect 2795 339 2801 340
rect 2795 338 2796 339
rect 2703 336 2796 338
rect 2703 335 2704 336
rect 2698 334 2704 335
rect 2795 335 2796 336
rect 2800 335 2801 339
rect 2795 334 2801 335
rect 2834 339 2840 340
rect 2834 335 2835 339
rect 2839 338 2840 339
rect 2947 339 2953 340
rect 2947 338 2948 339
rect 2839 336 2948 338
rect 2839 335 2840 336
rect 2834 334 2840 335
rect 2947 335 2948 336
rect 2952 335 2953 339
rect 2947 334 2953 335
rect 3107 339 3113 340
rect 3107 335 3108 339
rect 3112 338 3113 339
rect 3154 339 3160 340
rect 3154 338 3155 339
rect 3112 336 3155 338
rect 3112 335 3113 336
rect 3107 334 3113 335
rect 3154 335 3155 336
rect 3159 335 3160 339
rect 3154 334 3160 335
rect 3283 339 3289 340
rect 3283 335 3284 339
rect 3288 338 3289 339
rect 3298 339 3304 340
rect 3298 338 3299 339
rect 3288 336 3299 338
rect 3288 335 3289 336
rect 3283 334 3289 335
rect 3298 335 3299 336
rect 3303 335 3304 339
rect 3298 334 3304 335
rect 3459 339 3465 340
rect 3459 335 3460 339
rect 3464 338 3465 339
rect 3558 339 3564 340
rect 3558 338 3559 339
rect 3464 336 3559 338
rect 3464 335 3465 336
rect 3459 334 3465 335
rect 3558 335 3559 336
rect 3563 335 3564 339
rect 3682 339 3688 340
rect 3558 334 3564 335
rect 3643 337 3649 338
rect 1379 332 1385 333
rect 3643 333 3644 337
rect 3648 333 3649 337
rect 3682 335 3683 339
rect 3687 338 3688 339
rect 3827 339 3833 340
rect 3827 338 3828 339
rect 3687 336 3828 338
rect 3687 335 3688 336
rect 3682 334 3688 335
rect 3827 335 3828 336
rect 3832 335 3833 339
rect 3827 334 3833 335
rect 3643 332 3649 333
rect 1380 330 1382 332
rect 1818 331 1824 332
rect 1818 330 1819 331
rect 1380 328 1819 330
rect 1818 327 1819 328
rect 1823 327 1824 331
rect 1818 326 1824 327
rect 3498 331 3504 332
rect 3498 327 3499 331
rect 3503 330 3504 331
rect 3644 330 3646 332
rect 3503 328 3646 330
rect 3503 327 3504 328
rect 3498 326 3504 327
rect 110 320 116 321
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 158 319 164 320
rect 158 315 159 319
rect 163 315 164 319
rect 158 314 164 315
rect 350 319 356 320
rect 350 315 351 319
rect 355 315 356 319
rect 350 314 356 315
rect 550 319 556 320
rect 550 315 551 319
rect 555 315 556 319
rect 550 314 556 315
rect 758 319 764 320
rect 758 315 759 319
rect 763 315 764 319
rect 758 314 764 315
rect 958 319 964 320
rect 958 315 959 319
rect 963 315 964 319
rect 958 314 964 315
rect 1158 319 1164 320
rect 1158 315 1159 319
rect 1163 315 1164 319
rect 1158 314 1164 315
rect 1342 319 1348 320
rect 1342 315 1343 319
rect 1347 315 1348 319
rect 1342 314 1348 315
rect 1526 319 1532 320
rect 1526 315 1527 319
rect 1531 315 1532 319
rect 1526 314 1532 315
rect 1710 319 1716 320
rect 1710 315 1711 319
rect 1715 315 1716 319
rect 1710 314 1716 315
rect 1894 319 1900 320
rect 1894 315 1895 319
rect 1899 315 1900 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2398 319 2404 320
rect 2398 315 2399 319
rect 2403 315 2404 319
rect 1894 314 1900 315
rect 2398 314 2404 315
rect 2502 319 2508 320
rect 2502 315 2503 319
rect 2507 315 2508 319
rect 2502 314 2508 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2758 319 2764 320
rect 2758 315 2759 319
rect 2763 315 2764 319
rect 2758 314 2764 315
rect 2910 319 2916 320
rect 2910 315 2911 319
rect 2915 315 2916 319
rect 2910 314 2916 315
rect 3070 319 3076 320
rect 3070 315 3071 319
rect 3075 315 3076 319
rect 3070 314 3076 315
rect 3246 319 3252 320
rect 3246 315 3247 319
rect 3251 315 3252 319
rect 3246 314 3252 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3606 319 3612 320
rect 3606 315 3607 319
rect 3611 315 3612 319
rect 3606 314 3612 315
rect 3790 319 3796 320
rect 3790 315 3791 319
rect 3795 315 3796 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3790 314 3796 315
rect 151 311 157 312
rect 151 307 152 311
rect 156 310 157 311
rect 242 311 248 312
rect 156 308 201 310
rect 156 307 157 308
rect 151 306 157 307
rect 242 307 243 311
rect 247 310 248 311
rect 626 311 632 312
rect 247 308 393 310
rect 247 307 248 308
rect 242 306 248 307
rect 626 307 627 311
rect 631 307 632 311
rect 626 306 632 307
rect 834 311 840 312
rect 834 307 835 311
rect 839 307 840 311
rect 834 306 840 307
rect 902 311 908 312
rect 902 307 903 311
rect 907 310 908 311
rect 1234 311 1240 312
rect 907 308 1001 310
rect 907 307 908 308
rect 902 306 908 307
rect 1234 307 1235 311
rect 1239 307 1240 311
rect 1234 306 1240 307
rect 1418 311 1424 312
rect 1418 307 1419 311
rect 1423 307 1424 311
rect 1418 306 1424 307
rect 1602 311 1608 312
rect 1602 307 1603 311
rect 1607 307 1608 311
rect 1818 311 1824 312
rect 1602 306 1608 307
rect 1786 307 1792 308
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 1786 303 1787 307
rect 1791 303 1792 307
rect 1818 307 1819 311
rect 1823 310 1824 311
rect 2474 311 2480 312
rect 1823 308 1937 310
rect 1823 307 1824 308
rect 1818 306 1824 307
rect 2474 307 2475 311
rect 2479 307 2480 311
rect 2474 306 2480 307
rect 2578 311 2584 312
rect 2578 307 2579 311
rect 2583 307 2584 311
rect 2578 306 2584 307
rect 2698 311 2704 312
rect 2698 307 2699 311
rect 2703 307 2704 311
rect 2698 306 2704 307
rect 2834 311 2840 312
rect 2834 307 2835 311
rect 2839 307 2840 311
rect 2834 306 2840 307
rect 2858 311 2864 312
rect 2858 307 2859 311
rect 2863 310 2864 311
rect 3002 311 3008 312
rect 2863 308 2953 310
rect 2863 307 2864 308
rect 2858 306 2864 307
rect 3002 307 3003 311
rect 3007 310 3008 311
rect 3154 311 3160 312
rect 3007 308 3113 310
rect 3007 307 3008 308
rect 3002 306 3008 307
rect 3154 307 3155 311
rect 3159 310 3160 311
rect 3498 311 3504 312
rect 3159 308 3289 310
rect 3159 307 3160 308
rect 3154 306 3160 307
rect 3498 307 3499 311
rect 3503 307 3504 311
rect 3498 306 3504 307
rect 3682 311 3688 312
rect 3682 307 3683 311
rect 3687 307 3688 311
rect 3682 306 3688 307
rect 3866 307 3872 308
rect 1786 302 1792 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 158 300 164 301
rect 158 296 159 300
rect 163 296 164 300
rect 158 295 164 296
rect 350 300 356 301
rect 350 296 351 300
rect 355 296 356 300
rect 350 295 356 296
rect 550 300 556 301
rect 550 296 551 300
rect 555 296 556 300
rect 550 295 556 296
rect 758 300 764 301
rect 758 296 759 300
rect 763 296 764 300
rect 758 295 764 296
rect 958 300 964 301
rect 958 296 959 300
rect 963 296 964 300
rect 958 295 964 296
rect 1158 300 1164 301
rect 1158 296 1159 300
rect 1163 296 1164 300
rect 1158 295 1164 296
rect 1342 300 1348 301
rect 1342 296 1343 300
rect 1347 296 1348 300
rect 1342 295 1348 296
rect 1526 300 1532 301
rect 1526 296 1527 300
rect 1531 296 1532 300
rect 1526 295 1532 296
rect 1710 300 1716 301
rect 1710 296 1711 300
rect 1715 296 1716 300
rect 1710 295 1716 296
rect 1894 300 1900 301
rect 1894 296 1895 300
rect 1899 296 1900 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3866 303 3867 307
rect 3871 303 3872 307
rect 3866 302 3872 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2398 300 2404 301
rect 1894 295 1900 296
rect 2398 296 2399 300
rect 2403 296 2404 300
rect 2398 295 2404 296
rect 2502 300 2508 301
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2758 300 2764 301
rect 2758 296 2759 300
rect 2763 296 2764 300
rect 2758 295 2764 296
rect 2910 300 2916 301
rect 2910 296 2911 300
rect 2915 296 2916 300
rect 2910 295 2916 296
rect 3070 300 3076 301
rect 3070 296 3071 300
rect 3075 296 3076 300
rect 3070 295 3076 296
rect 3246 300 3252 301
rect 3246 296 3247 300
rect 3251 296 3252 300
rect 3246 295 3252 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3606 300 3612 301
rect 3606 296 3607 300
rect 3611 296 3612 300
rect 3606 295 3612 296
rect 3790 300 3796 301
rect 3790 296 3791 300
rect 3795 296 3796 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3790 295 3796 296
rect 2438 247 2444 248
rect 2438 243 2439 247
rect 2443 246 2444 247
rect 2443 244 2606 246
rect 2443 243 2444 244
rect 2438 242 2444 243
rect 2190 240 2196 241
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2190 236 2191 240
rect 2195 236 2196 240
rect 2190 235 2196 236
rect 2350 240 2356 241
rect 2350 236 2351 240
rect 2355 236 2356 240
rect 2350 235 2356 236
rect 2518 240 2524 241
rect 2518 236 2519 240
rect 2523 236 2524 240
rect 2518 235 2524 236
rect 222 232 228 233
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 222 228 223 232
rect 227 228 228 232
rect 222 227 228 228
rect 382 232 388 233
rect 382 228 383 232
rect 387 228 388 232
rect 382 227 388 228
rect 542 232 548 233
rect 542 228 543 232
rect 547 228 548 232
rect 542 227 548 228
rect 702 232 708 233
rect 702 228 703 232
rect 707 228 708 232
rect 702 227 708 228
rect 862 232 868 233
rect 862 228 863 232
rect 867 228 868 232
rect 862 227 868 228
rect 1030 232 1036 233
rect 1030 228 1031 232
rect 1035 228 1036 232
rect 1030 227 1036 228
rect 1198 232 1204 233
rect 1198 228 1199 232
rect 1203 228 1204 232
rect 1198 227 1204 228
rect 1366 232 1372 233
rect 1366 228 1367 232
rect 1371 228 1372 232
rect 1366 227 1372 228
rect 1542 232 1548 233
rect 1542 228 1543 232
rect 1547 228 1548 232
rect 1542 227 1548 228
rect 1726 232 1732 233
rect 1726 228 1727 232
rect 1731 228 1732 232
rect 1726 227 1732 228
rect 1902 232 1908 233
rect 2046 232 2052 233
rect 1902 228 1903 232
rect 1907 228 1908 232
rect 2266 231 2272 232
rect 1902 227 1908 228
rect 2006 229 2012 230
rect 110 224 116 225
rect 2006 225 2007 229
rect 2011 225 2012 229
rect 2266 227 2267 231
rect 2271 227 2272 231
rect 2266 226 2272 227
rect 2426 231 2432 232
rect 2426 227 2427 231
rect 2431 227 2432 231
rect 2426 226 2432 227
rect 2594 231 2600 232
rect 2594 227 2595 231
rect 2599 227 2600 231
rect 2604 230 2606 244
rect 2686 240 2692 241
rect 2686 236 2687 240
rect 2691 236 2692 240
rect 2686 235 2692 236
rect 2854 240 2860 241
rect 2854 236 2855 240
rect 2859 236 2860 240
rect 2854 235 2860 236
rect 3030 240 3036 241
rect 3030 236 3031 240
rect 3035 236 3036 240
rect 3030 235 3036 236
rect 3214 240 3220 241
rect 3214 236 3215 240
rect 3219 236 3220 240
rect 3214 235 3220 236
rect 3406 240 3412 241
rect 3406 236 3407 240
rect 3411 236 3412 240
rect 3406 235 3412 236
rect 3606 240 3612 241
rect 3606 236 3607 240
rect 3611 236 3612 240
rect 3606 235 3612 236
rect 3806 240 3812 241
rect 3806 236 3807 240
rect 3811 236 3812 240
rect 3806 235 3812 236
rect 3942 237 3948 238
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 2930 231 2936 232
rect 2604 228 2729 230
rect 2594 226 2600 227
rect 2930 227 2931 231
rect 2935 227 2936 231
rect 2930 226 2936 227
rect 3106 231 3112 232
rect 3106 227 3107 231
rect 3111 227 3112 231
rect 3106 226 3112 227
rect 3290 231 3296 232
rect 3290 227 3291 231
rect 3295 227 3296 231
rect 3290 226 3296 227
rect 3378 231 3384 232
rect 3378 227 3379 231
rect 3383 230 3384 231
rect 3558 231 3564 232
rect 3383 228 3449 230
rect 3383 227 3384 228
rect 3378 226 3384 227
rect 3558 227 3559 231
rect 3563 230 3564 231
rect 3782 231 3788 232
rect 3563 228 3649 230
rect 3563 227 3564 228
rect 3558 226 3564 227
rect 3782 227 3783 231
rect 3787 230 3788 231
rect 3787 228 3849 230
rect 3787 227 3788 228
rect 3782 226 3788 227
rect 2006 224 2012 225
rect 298 223 304 224
rect 298 219 299 223
rect 303 219 304 223
rect 298 218 304 219
rect 375 223 381 224
rect 375 219 376 223
rect 380 222 381 223
rect 618 223 624 224
rect 380 220 425 222
rect 380 219 381 220
rect 375 218 381 219
rect 618 219 619 223
rect 623 219 624 223
rect 618 218 624 219
rect 639 223 645 224
rect 639 219 640 223
rect 644 222 645 223
rect 798 223 804 224
rect 644 220 745 222
rect 644 219 645 220
rect 639 218 645 219
rect 798 219 799 223
rect 803 222 804 223
rect 1098 223 1104 224
rect 803 220 905 222
rect 803 219 804 220
rect 798 218 804 219
rect 1098 219 1099 223
rect 1103 219 1104 223
rect 1098 218 1104 219
rect 1114 223 1120 224
rect 1114 219 1115 223
rect 1119 222 1120 223
rect 1295 223 1301 224
rect 1119 220 1241 222
rect 1119 219 1120 220
rect 1114 218 1120 219
rect 1295 219 1296 223
rect 1300 222 1301 223
rect 1471 223 1477 224
rect 1300 220 1409 222
rect 1300 219 1301 220
rect 1295 218 1301 219
rect 1471 219 1472 223
rect 1476 222 1477 223
rect 1626 223 1632 224
rect 1476 220 1585 222
rect 1476 219 1477 220
rect 1471 218 1477 219
rect 1626 219 1627 223
rect 1631 222 1632 223
rect 1970 223 1976 224
rect 1631 220 1769 222
rect 1631 219 1632 220
rect 1626 218 1632 219
rect 1970 219 1971 223
rect 1975 219 1976 223
rect 2190 221 2196 222
rect 1970 218 1976 219
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2190 217 2191 221
rect 2195 217 2196 221
rect 2190 216 2196 217
rect 2350 221 2356 222
rect 2350 217 2351 221
rect 2355 217 2356 221
rect 2350 216 2356 217
rect 2518 221 2524 222
rect 2518 217 2519 221
rect 2523 217 2524 221
rect 2518 216 2524 217
rect 2686 221 2692 222
rect 2686 217 2687 221
rect 2691 217 2692 221
rect 2686 216 2692 217
rect 2854 221 2860 222
rect 2854 217 2855 221
rect 2859 217 2860 221
rect 2854 216 2860 217
rect 3030 221 3036 222
rect 3030 217 3031 221
rect 3035 217 3036 221
rect 3030 216 3036 217
rect 3214 221 3220 222
rect 3214 217 3215 221
rect 3219 217 3220 221
rect 3214 216 3220 217
rect 3406 221 3412 222
rect 3406 217 3407 221
rect 3411 217 3412 221
rect 3406 216 3412 217
rect 3606 221 3612 222
rect 3606 217 3607 221
rect 3611 217 3612 221
rect 3606 216 3612 217
rect 3806 221 3812 222
rect 3806 217 3807 221
rect 3811 217 3812 221
rect 3806 216 3812 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 222 213 228 214
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 222 209 223 213
rect 227 209 228 213
rect 222 208 228 209
rect 382 213 388 214
rect 382 209 383 213
rect 387 209 388 213
rect 382 208 388 209
rect 542 213 548 214
rect 542 209 543 213
rect 547 209 548 213
rect 542 208 548 209
rect 702 213 708 214
rect 702 209 703 213
rect 707 209 708 213
rect 702 208 708 209
rect 862 213 868 214
rect 862 209 863 213
rect 867 209 868 213
rect 862 208 868 209
rect 1030 213 1036 214
rect 1030 209 1031 213
rect 1035 209 1036 213
rect 1030 208 1036 209
rect 1198 213 1204 214
rect 1198 209 1199 213
rect 1203 209 1204 213
rect 1198 208 1204 209
rect 1366 213 1372 214
rect 1366 209 1367 213
rect 1371 209 1372 213
rect 1366 208 1372 209
rect 1542 213 1548 214
rect 1542 209 1543 213
rect 1547 209 1548 213
rect 1542 208 1548 209
rect 1726 213 1732 214
rect 1726 209 1727 213
rect 1731 209 1732 213
rect 1726 208 1732 209
rect 1902 213 1908 214
rect 1902 209 1903 213
rect 1907 209 1908 213
rect 1902 208 1908 209
rect 2006 212 2012 213
rect 2006 208 2007 212
rect 2011 208 2012 212
rect 3002 211 3008 212
rect 3002 210 3003 211
rect 110 207 116 208
rect 2006 207 2012 208
rect 2924 208 3003 210
rect 2266 203 2272 204
rect 2227 199 2233 200
rect 298 195 304 196
rect 259 191 265 192
rect 259 187 260 191
rect 264 190 265 191
rect 298 191 299 195
rect 303 194 304 195
rect 419 195 425 196
rect 419 194 420 195
rect 303 192 420 194
rect 303 191 304 192
rect 298 190 304 191
rect 419 191 420 192
rect 424 191 425 195
rect 419 190 425 191
rect 579 195 585 196
rect 579 191 580 195
rect 584 194 585 195
rect 639 195 645 196
rect 639 194 640 195
rect 584 192 640 194
rect 584 191 585 192
rect 579 190 585 191
rect 639 191 640 192
rect 644 191 645 195
rect 639 190 645 191
rect 739 195 745 196
rect 739 191 740 195
rect 744 194 745 195
rect 798 195 804 196
rect 798 194 799 195
rect 744 192 799 194
rect 744 191 745 192
rect 739 190 745 191
rect 798 191 799 192
rect 803 191 804 195
rect 798 190 804 191
rect 899 195 908 196
rect 899 191 900 195
rect 907 191 908 195
rect 899 190 908 191
rect 1067 195 1073 196
rect 1067 191 1068 195
rect 1072 194 1073 195
rect 1114 195 1120 196
rect 1114 194 1115 195
rect 1072 192 1115 194
rect 1072 191 1073 192
rect 1067 190 1073 191
rect 1114 191 1115 192
rect 1119 191 1120 195
rect 1114 190 1120 191
rect 1235 195 1241 196
rect 1235 191 1236 195
rect 1240 194 1241 195
rect 1295 195 1301 196
rect 1295 194 1296 195
rect 1240 192 1296 194
rect 1240 191 1241 192
rect 1235 190 1241 191
rect 1295 191 1296 192
rect 1300 191 1301 195
rect 1295 190 1301 191
rect 1403 195 1409 196
rect 1403 191 1404 195
rect 1408 194 1409 195
rect 1471 195 1477 196
rect 1471 194 1472 195
rect 1408 192 1472 194
rect 1408 191 1409 192
rect 1403 190 1409 191
rect 1471 191 1472 192
rect 1476 191 1477 195
rect 1471 190 1477 191
rect 1579 195 1585 196
rect 1579 191 1580 195
rect 1584 194 1585 195
rect 1626 195 1632 196
rect 1626 194 1627 195
rect 1584 192 1627 194
rect 1584 191 1585 192
rect 1579 190 1585 191
rect 1626 191 1627 192
rect 1631 191 1632 195
rect 1626 190 1632 191
rect 1763 195 1769 196
rect 1763 191 1764 195
rect 1768 194 1769 195
rect 1786 195 1792 196
rect 1786 194 1787 195
rect 1768 192 1787 194
rect 1768 191 1769 192
rect 1763 190 1769 191
rect 1786 191 1787 192
rect 1791 191 1792 195
rect 2227 195 2228 199
rect 2232 198 2233 199
rect 2266 199 2267 203
rect 2271 202 2272 203
rect 2387 203 2393 204
rect 2387 202 2388 203
rect 2271 200 2388 202
rect 2271 199 2272 200
rect 2266 198 2272 199
rect 2387 199 2388 200
rect 2392 199 2393 203
rect 2387 198 2393 199
rect 2426 203 2432 204
rect 2426 199 2427 203
rect 2431 202 2432 203
rect 2555 203 2561 204
rect 2555 202 2556 203
rect 2431 200 2556 202
rect 2431 199 2432 200
rect 2426 198 2432 199
rect 2555 199 2556 200
rect 2560 199 2561 203
rect 2555 198 2561 199
rect 2594 203 2600 204
rect 2594 199 2595 203
rect 2599 202 2600 203
rect 2723 203 2729 204
rect 2723 202 2724 203
rect 2599 200 2724 202
rect 2599 199 2600 200
rect 2594 198 2600 199
rect 2723 199 2724 200
rect 2728 199 2729 203
rect 2723 198 2729 199
rect 2891 203 2897 204
rect 2891 199 2892 203
rect 2896 202 2897 203
rect 2924 202 2926 208
rect 3002 207 3003 208
rect 3007 207 3008 211
rect 3002 206 3008 207
rect 2896 200 2926 202
rect 2930 203 2936 204
rect 2896 199 2897 200
rect 2891 198 2897 199
rect 2930 199 2931 203
rect 2935 202 2936 203
rect 3067 203 3073 204
rect 3067 202 3068 203
rect 2935 200 3068 202
rect 2935 199 2936 200
rect 2930 198 2936 199
rect 3067 199 3068 200
rect 3072 199 3073 203
rect 3067 198 3073 199
rect 3106 203 3112 204
rect 3106 199 3107 203
rect 3111 202 3112 203
rect 3251 203 3257 204
rect 3251 202 3252 203
rect 3111 200 3252 202
rect 3111 199 3112 200
rect 3106 198 3112 199
rect 3251 199 3252 200
rect 3256 199 3257 203
rect 3251 198 3257 199
rect 3290 203 3296 204
rect 3290 199 3291 203
rect 3295 202 3296 203
rect 3443 203 3449 204
rect 3443 202 3444 203
rect 3295 200 3444 202
rect 3295 199 3296 200
rect 3290 198 3296 199
rect 3443 199 3444 200
rect 3448 199 3449 203
rect 3843 203 3849 204
rect 3443 198 3449 199
rect 3631 199 3637 200
rect 2232 196 2262 198
rect 2232 195 2233 196
rect 2227 194 2233 195
rect 1786 190 1792 191
rect 1882 191 1888 192
rect 264 188 270 190
rect 264 187 265 188
rect 259 186 265 187
rect 268 186 270 188
rect 306 187 312 188
rect 306 186 307 187
rect 268 184 307 186
rect 306 183 307 184
rect 311 183 312 187
rect 1882 187 1883 191
rect 1887 190 1888 191
rect 1939 191 1945 192
rect 1939 190 1940 191
rect 1887 188 1940 190
rect 1887 187 1888 188
rect 1882 186 1888 187
rect 1939 187 1940 188
rect 1944 187 1945 191
rect 2260 190 2262 196
rect 3631 195 3632 199
rect 3636 198 3637 199
rect 3643 199 3649 200
rect 3643 198 3644 199
rect 3636 196 3644 198
rect 3636 195 3637 196
rect 3631 194 3637 195
rect 3643 195 3644 196
rect 3648 195 3649 199
rect 3843 199 3844 203
rect 3848 202 3849 203
rect 3866 203 3872 204
rect 3866 202 3867 203
rect 3848 200 3867 202
rect 3848 199 3849 200
rect 3843 198 3849 199
rect 3866 199 3867 200
rect 3871 199 3872 203
rect 3866 198 3872 199
rect 3643 194 3649 195
rect 2726 191 2732 192
rect 2726 190 2727 191
rect 2260 188 2727 190
rect 1939 186 1945 187
rect 2726 187 2727 188
rect 2731 187 2732 191
rect 2726 186 2732 187
rect 306 182 312 183
rect 3378 163 3384 164
rect 3378 162 3379 163
rect 2908 160 3379 162
rect 210 159 216 160
rect 171 157 177 158
rect 171 153 172 157
rect 176 153 177 157
rect 210 155 211 159
rect 215 158 216 159
rect 267 159 273 160
rect 267 158 268 159
rect 215 156 268 158
rect 215 155 216 156
rect 210 154 216 155
rect 267 155 268 156
rect 272 155 273 159
rect 267 154 273 155
rect 363 159 369 160
rect 363 155 364 159
rect 368 158 369 159
rect 410 159 416 160
rect 410 158 411 159
rect 368 156 411 158
rect 368 155 369 156
rect 363 154 369 155
rect 410 155 411 156
rect 415 155 416 159
rect 410 154 416 155
rect 459 159 465 160
rect 459 155 460 159
rect 464 158 465 159
rect 506 159 512 160
rect 506 158 507 159
rect 464 156 507 158
rect 464 155 465 156
rect 459 154 465 155
rect 506 155 507 156
rect 511 155 512 159
rect 618 159 624 160
rect 506 154 512 155
rect 563 157 569 158
rect 171 152 177 153
rect 563 153 564 157
rect 568 153 569 157
rect 618 155 619 159
rect 623 158 624 159
rect 683 159 689 160
rect 683 158 684 159
rect 623 156 684 158
rect 623 155 624 156
rect 618 154 624 155
rect 683 155 684 156
rect 688 155 689 159
rect 683 154 689 155
rect 722 159 728 160
rect 722 155 723 159
rect 727 158 728 159
rect 811 159 817 160
rect 811 158 812 159
rect 727 156 812 158
rect 727 155 728 156
rect 722 154 728 155
rect 811 155 812 156
rect 816 155 817 159
rect 811 154 817 155
rect 850 159 856 160
rect 850 155 851 159
rect 855 158 856 159
rect 939 159 945 160
rect 939 158 940 159
rect 855 156 940 158
rect 855 155 856 156
rect 850 154 856 155
rect 939 155 940 156
rect 944 155 945 159
rect 939 154 945 155
rect 1067 159 1073 160
rect 1067 155 1068 159
rect 1072 158 1073 159
rect 1098 159 1104 160
rect 1098 158 1099 159
rect 1072 156 1099 158
rect 1072 155 1073 156
rect 1067 154 1073 155
rect 1098 155 1099 156
rect 1103 155 1104 159
rect 1098 154 1104 155
rect 1106 159 1112 160
rect 1106 155 1107 159
rect 1111 158 1112 159
rect 1187 159 1193 160
rect 1187 158 1188 159
rect 1111 156 1188 158
rect 1111 155 1112 156
rect 1106 154 1112 155
rect 1187 155 1188 156
rect 1192 155 1193 159
rect 1187 154 1193 155
rect 1226 159 1232 160
rect 1226 155 1227 159
rect 1231 158 1232 159
rect 1307 159 1313 160
rect 1307 158 1308 159
rect 1231 156 1308 158
rect 1231 155 1232 156
rect 1226 154 1232 155
rect 1307 155 1308 156
rect 1312 155 1313 159
rect 1307 154 1313 155
rect 1346 159 1352 160
rect 1346 155 1347 159
rect 1351 158 1352 159
rect 1419 159 1425 160
rect 1419 158 1420 159
rect 1351 156 1420 158
rect 1351 155 1352 156
rect 1346 154 1352 155
rect 1419 155 1420 156
rect 1424 155 1425 159
rect 1419 154 1425 155
rect 1458 159 1464 160
rect 1458 155 1459 159
rect 1463 158 1464 159
rect 1523 159 1529 160
rect 1523 158 1524 159
rect 1463 156 1524 158
rect 1463 155 1464 156
rect 1458 154 1464 155
rect 1523 155 1524 156
rect 1528 155 1529 159
rect 1523 154 1529 155
rect 1562 159 1568 160
rect 1562 155 1563 159
rect 1567 158 1568 159
rect 1627 159 1633 160
rect 1627 158 1628 159
rect 1567 156 1628 158
rect 1567 155 1568 156
rect 1562 154 1568 155
rect 1627 155 1628 156
rect 1632 155 1633 159
rect 1627 154 1633 155
rect 1666 159 1672 160
rect 1666 155 1667 159
rect 1671 158 1672 159
rect 1739 159 1745 160
rect 1739 158 1740 159
rect 1671 156 1740 158
rect 1671 155 1672 156
rect 1666 154 1672 155
rect 1739 155 1740 156
rect 1744 155 1745 159
rect 1739 154 1745 155
rect 1778 159 1784 160
rect 1778 155 1779 159
rect 1783 158 1784 159
rect 1843 159 1849 160
rect 1843 158 1844 159
rect 1783 156 1844 158
rect 1783 155 1784 156
rect 1778 154 1784 155
rect 1843 155 1844 156
rect 1848 155 1849 159
rect 1843 154 1849 155
rect 1939 159 1945 160
rect 1939 155 1940 159
rect 1944 158 1945 159
rect 1970 159 1976 160
rect 1970 158 1971 159
rect 1944 156 1971 158
rect 1944 155 1945 156
rect 1939 154 1945 155
rect 1970 155 1971 156
rect 1975 155 1976 159
rect 2908 158 2910 160
rect 3378 159 3379 160
rect 3383 159 3384 163
rect 3378 158 3384 159
rect 2907 157 2913 158
rect 1970 154 1976 155
rect 1978 155 1984 156
rect 563 152 569 153
rect 172 150 174 152
rect 314 151 320 152
rect 314 150 315 151
rect 172 148 315 150
rect 314 147 315 148
rect 319 147 320 151
rect 564 150 566 152
rect 858 151 864 152
rect 858 150 859 151
rect 564 148 859 150
rect 314 146 320 147
rect 858 147 859 148
rect 863 147 864 151
rect 1978 151 1979 155
rect 1983 154 1984 155
rect 2107 155 2113 156
rect 2107 154 2108 155
rect 1983 152 2108 154
rect 1983 151 1984 152
rect 1978 150 1984 151
rect 2107 151 2108 152
rect 2112 151 2113 155
rect 2107 150 2113 151
rect 2146 155 2152 156
rect 2146 151 2147 155
rect 2151 154 2152 155
rect 2203 155 2209 156
rect 2203 154 2204 155
rect 2151 152 2204 154
rect 2151 151 2152 152
rect 2146 150 2152 151
rect 2203 151 2204 152
rect 2208 151 2209 155
rect 2203 150 2209 151
rect 2242 155 2248 156
rect 2242 151 2243 155
rect 2247 154 2248 155
rect 2299 155 2305 156
rect 2299 154 2300 155
rect 2247 152 2300 154
rect 2247 151 2248 152
rect 2242 150 2248 151
rect 2299 151 2300 152
rect 2304 151 2305 155
rect 2299 150 2305 151
rect 2338 155 2344 156
rect 2338 151 2339 155
rect 2343 154 2344 155
rect 2403 155 2409 156
rect 2403 154 2404 155
rect 2343 152 2404 154
rect 2343 151 2344 152
rect 2338 150 2344 151
rect 2403 151 2404 152
rect 2408 151 2409 155
rect 2403 150 2409 151
rect 2442 155 2448 156
rect 2442 151 2443 155
rect 2447 154 2448 155
rect 2523 155 2529 156
rect 2523 154 2524 155
rect 2447 152 2524 154
rect 2447 151 2448 152
rect 2442 150 2448 151
rect 2523 151 2524 152
rect 2528 151 2529 155
rect 2523 150 2529 151
rect 2562 155 2568 156
rect 2562 151 2563 155
rect 2567 154 2568 155
rect 2651 155 2657 156
rect 2651 154 2652 155
rect 2567 152 2652 154
rect 2567 151 2568 152
rect 2562 150 2568 151
rect 2651 151 2652 152
rect 2656 151 2657 155
rect 2651 150 2657 151
rect 2718 155 2724 156
rect 2718 151 2719 155
rect 2723 154 2724 155
rect 2779 155 2785 156
rect 2779 154 2780 155
rect 2723 152 2780 154
rect 2723 151 2724 152
rect 2718 150 2724 151
rect 2779 151 2780 152
rect 2784 151 2785 155
rect 2907 153 2908 157
rect 2912 153 2913 157
rect 2907 152 2913 153
rect 2946 155 2952 156
rect 2779 150 2785 151
rect 2946 151 2947 155
rect 2951 154 2952 155
rect 3027 155 3033 156
rect 3027 154 3028 155
rect 2951 152 3028 154
rect 2951 151 2952 152
rect 2946 150 2952 151
rect 3027 151 3028 152
rect 3032 151 3033 155
rect 3027 150 3033 151
rect 3066 155 3072 156
rect 3066 151 3067 155
rect 3071 154 3072 155
rect 3147 155 3153 156
rect 3147 154 3148 155
rect 3071 152 3148 154
rect 3071 151 3072 152
rect 3066 150 3072 151
rect 3147 151 3148 152
rect 3152 151 3153 155
rect 3147 150 3153 151
rect 3186 155 3192 156
rect 3186 151 3187 155
rect 3191 154 3192 155
rect 3259 155 3265 156
rect 3259 154 3260 155
rect 3191 152 3260 154
rect 3191 151 3192 152
rect 3186 150 3192 151
rect 3259 151 3260 152
rect 3264 151 3265 155
rect 3259 150 3265 151
rect 3298 155 3304 156
rect 3298 151 3299 155
rect 3303 154 3304 155
rect 3363 155 3369 156
rect 3363 154 3364 155
rect 3303 152 3364 154
rect 3303 151 3304 152
rect 3298 150 3304 151
rect 3363 151 3364 152
rect 3368 151 3369 155
rect 3363 150 3369 151
rect 3415 155 3421 156
rect 3415 151 3416 155
rect 3420 154 3421 155
rect 3467 155 3473 156
rect 3467 154 3468 155
rect 3420 152 3468 154
rect 3420 151 3421 152
rect 3415 150 3421 151
rect 3467 151 3468 152
rect 3472 151 3473 155
rect 3467 150 3473 151
rect 3506 155 3512 156
rect 3506 151 3507 155
rect 3511 154 3512 155
rect 3571 155 3577 156
rect 3571 154 3572 155
rect 3511 152 3572 154
rect 3511 151 3512 152
rect 3506 150 3512 151
rect 3571 151 3572 152
rect 3576 151 3577 155
rect 3571 150 3577 151
rect 3623 155 3629 156
rect 3623 151 3624 155
rect 3628 154 3629 155
rect 3675 155 3681 156
rect 3675 154 3676 155
rect 3628 152 3676 154
rect 3628 151 3629 152
rect 3623 150 3629 151
rect 3675 151 3676 152
rect 3680 151 3681 155
rect 3675 150 3681 151
rect 3779 155 3788 156
rect 3779 151 3780 155
rect 3787 151 3788 155
rect 3779 150 3788 151
rect 3818 155 3824 156
rect 3818 151 3819 155
rect 3823 154 3824 155
rect 3875 155 3881 156
rect 3875 154 3876 155
rect 3823 152 3876 154
rect 3823 151 3824 152
rect 3818 150 3824 151
rect 3875 151 3876 152
rect 3880 151 3881 155
rect 3875 150 3881 151
rect 858 146 864 147
rect 110 140 116 141
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2006 135 2012 136
rect 2046 136 2052 137
rect 3942 136 3948 137
rect 1902 134 1908 135
rect 2046 132 2047 136
rect 2051 132 2052 136
rect 210 131 216 132
rect 210 127 211 131
rect 215 127 216 131
rect 210 126 216 127
rect 306 131 312 132
rect 306 127 307 131
rect 311 127 312 131
rect 306 126 312 127
rect 314 131 320 132
rect 314 127 315 131
rect 319 130 320 131
rect 410 131 416 132
rect 319 128 369 130
rect 319 127 320 128
rect 314 126 320 127
rect 410 127 411 131
rect 415 130 416 131
rect 506 131 512 132
rect 415 128 465 130
rect 415 127 416 128
rect 410 126 416 127
rect 506 127 507 131
rect 511 130 512 131
rect 722 131 728 132
rect 511 128 569 130
rect 511 127 512 128
rect 506 126 512 127
rect 722 127 723 131
rect 727 127 728 131
rect 722 126 728 127
rect 850 131 856 132
rect 850 127 851 131
rect 855 127 856 131
rect 850 126 856 127
rect 858 131 864 132
rect 858 127 859 131
rect 863 130 864 131
rect 1106 131 1112 132
rect 863 128 945 130
rect 863 127 864 128
rect 858 126 864 127
rect 1106 127 1107 131
rect 1111 127 1112 131
rect 1106 126 1112 127
rect 1226 131 1232 132
rect 1226 127 1227 131
rect 1231 127 1232 131
rect 1226 126 1232 127
rect 1346 131 1352 132
rect 1346 127 1347 131
rect 1351 127 1352 131
rect 1346 126 1352 127
rect 1458 131 1464 132
rect 1458 127 1459 131
rect 1463 127 1464 131
rect 1458 126 1464 127
rect 1562 131 1568 132
rect 1562 127 1563 131
rect 1567 127 1568 131
rect 1562 126 1568 127
rect 1666 131 1672 132
rect 1666 127 1667 131
rect 1671 127 1672 131
rect 1666 126 1672 127
rect 1778 131 1784 132
rect 1778 127 1779 131
rect 1783 127 1784 131
rect 1778 126 1784 127
rect 1882 131 1888 132
rect 1882 127 1883 131
rect 1887 127 1888 131
rect 1882 126 1888 127
rect 1978 131 1984 132
rect 2046 131 2052 132
rect 2070 135 2076 136
rect 2070 131 2071 135
rect 2075 131 2076 135
rect 1978 127 1979 131
rect 1983 127 1984 131
rect 2070 130 2076 131
rect 2166 135 2172 136
rect 2166 131 2167 135
rect 2171 131 2172 135
rect 2166 130 2172 131
rect 2262 135 2268 136
rect 2262 131 2263 135
rect 2267 131 2268 135
rect 2262 130 2268 131
rect 2366 135 2372 136
rect 2366 131 2367 135
rect 2371 131 2372 135
rect 2366 130 2372 131
rect 2486 135 2492 136
rect 2486 131 2487 135
rect 2491 131 2492 135
rect 2486 130 2492 131
rect 2614 135 2620 136
rect 2614 131 2615 135
rect 2619 131 2620 135
rect 2614 130 2620 131
rect 2742 135 2748 136
rect 2742 131 2743 135
rect 2747 131 2748 135
rect 2742 130 2748 131
rect 2870 135 2876 136
rect 2870 131 2871 135
rect 2875 131 2876 135
rect 2870 130 2876 131
rect 2990 135 2996 136
rect 2990 131 2991 135
rect 2995 131 2996 135
rect 2990 130 2996 131
rect 3110 135 3116 136
rect 3110 131 3111 135
rect 3115 131 3116 135
rect 3110 130 3116 131
rect 3222 135 3228 136
rect 3222 131 3223 135
rect 3227 131 3228 135
rect 3222 130 3228 131
rect 3326 135 3332 136
rect 3326 131 3327 135
rect 3331 131 3332 135
rect 3326 130 3332 131
rect 3430 135 3436 136
rect 3430 131 3431 135
rect 3435 131 3436 135
rect 3430 130 3436 131
rect 3534 135 3540 136
rect 3534 131 3535 135
rect 3539 131 3540 135
rect 3534 130 3540 131
rect 3638 135 3644 136
rect 3638 131 3639 135
rect 3643 131 3644 135
rect 3638 130 3644 131
rect 3742 135 3748 136
rect 3742 131 3743 135
rect 3747 131 3748 135
rect 3742 130 3748 131
rect 3838 135 3844 136
rect 3838 131 3839 135
rect 3843 131 3844 135
rect 3942 132 3943 136
rect 3947 132 3948 136
rect 3942 131 3948 132
rect 3838 130 3844 131
rect 1978 126 1984 127
rect 2146 127 2152 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2146 123 2147 127
rect 2151 123 2152 127
rect 2146 122 2152 123
rect 2242 127 2248 128
rect 2242 123 2243 127
rect 2247 123 2248 127
rect 2242 122 2248 123
rect 2338 127 2344 128
rect 2338 123 2339 127
rect 2343 123 2344 127
rect 2338 122 2344 123
rect 2442 127 2448 128
rect 2442 123 2443 127
rect 2447 123 2448 127
rect 2442 122 2448 123
rect 2562 127 2568 128
rect 2562 123 2563 127
rect 2567 123 2568 127
rect 2718 127 2724 128
rect 2718 126 2719 127
rect 2693 124 2719 126
rect 2562 122 2568 123
rect 2718 123 2719 124
rect 2723 123 2724 127
rect 2718 122 2724 123
rect 2726 127 2732 128
rect 2726 123 2727 127
rect 2731 126 2732 127
rect 2946 127 2952 128
rect 2731 124 2785 126
rect 2731 123 2732 124
rect 2726 122 2732 123
rect 2946 123 2947 127
rect 2951 123 2952 127
rect 2946 122 2952 123
rect 3066 127 3072 128
rect 3066 123 3067 127
rect 3071 123 3072 127
rect 3066 122 3072 123
rect 3186 127 3192 128
rect 3186 123 3187 127
rect 3191 123 3192 127
rect 3186 122 3192 123
rect 3298 127 3304 128
rect 3298 123 3299 127
rect 3303 123 3304 127
rect 3415 127 3421 128
rect 3415 126 3416 127
rect 3405 124 3416 126
rect 3298 122 3304 123
rect 3415 123 3416 124
rect 3420 123 3421 127
rect 3415 122 3421 123
rect 3506 127 3512 128
rect 3506 123 3507 127
rect 3511 123 3512 127
rect 3623 127 3629 128
rect 3623 126 3624 127
rect 3613 124 3624 126
rect 3506 122 3512 123
rect 3623 123 3624 124
rect 3628 123 3629 127
rect 3623 122 3629 123
rect 3631 127 3637 128
rect 3631 123 3632 127
rect 3636 126 3637 127
rect 3818 127 3824 128
rect 3636 124 3681 126
rect 3636 123 3637 124
rect 3631 122 3637 123
rect 3818 123 3819 127
rect 3823 123 3824 127
rect 3818 122 3824 123
rect 2006 118 2012 119
rect 2046 119 2052 120
rect 1902 115 1908 116
rect 2046 115 2047 119
rect 2051 115 2052 119
rect 3942 119 3948 120
rect 2046 114 2052 115
rect 2070 116 2076 117
rect 2070 112 2071 116
rect 2075 112 2076 116
rect 2070 111 2076 112
rect 2166 116 2172 117
rect 2166 112 2167 116
rect 2171 112 2172 116
rect 2166 111 2172 112
rect 2262 116 2268 117
rect 2262 112 2263 116
rect 2267 112 2268 116
rect 2262 111 2268 112
rect 2366 116 2372 117
rect 2366 112 2367 116
rect 2371 112 2372 116
rect 2366 111 2372 112
rect 2486 116 2492 117
rect 2486 112 2487 116
rect 2491 112 2492 116
rect 2486 111 2492 112
rect 2614 116 2620 117
rect 2614 112 2615 116
rect 2619 112 2620 116
rect 2614 111 2620 112
rect 2742 116 2748 117
rect 2742 112 2743 116
rect 2747 112 2748 116
rect 2742 111 2748 112
rect 2870 116 2876 117
rect 2870 112 2871 116
rect 2875 112 2876 116
rect 2870 111 2876 112
rect 2990 116 2996 117
rect 2990 112 2991 116
rect 2995 112 2996 116
rect 2990 111 2996 112
rect 3110 116 3116 117
rect 3110 112 3111 116
rect 3115 112 3116 116
rect 3110 111 3116 112
rect 3222 116 3228 117
rect 3222 112 3223 116
rect 3227 112 3228 116
rect 3222 111 3228 112
rect 3326 116 3332 117
rect 3326 112 3327 116
rect 3331 112 3332 116
rect 3326 111 3332 112
rect 3430 116 3436 117
rect 3430 112 3431 116
rect 3435 112 3436 116
rect 3430 111 3436 112
rect 3534 116 3540 117
rect 3534 112 3535 116
rect 3539 112 3540 116
rect 3534 111 3540 112
rect 3638 116 3644 117
rect 3638 112 3639 116
rect 3643 112 3644 116
rect 3638 111 3644 112
rect 3742 116 3748 117
rect 3742 112 3743 116
rect 3747 112 3748 116
rect 3742 111 3748 112
rect 3838 116 3844 117
rect 3838 112 3839 116
rect 3843 112 3844 116
rect 3942 115 3943 119
rect 3947 115 3948 119
rect 3942 114 3948 115
rect 3838 111 3844 112
<< m3c >>
rect 1979 4019 1983 4023
rect 227 3999 231 4003
rect 355 3999 359 4003
rect 507 3999 511 4003
rect 683 3999 687 4003
rect 867 3999 871 4003
rect 1227 3999 1231 4003
rect 1387 3999 1391 4003
rect 1547 3999 1551 4003
rect 1699 3999 1703 4003
rect 1851 3999 1855 4003
rect 2047 4000 2051 4004
rect 2071 3999 2075 4003
rect 3943 4000 3947 4004
rect 1411 3991 1415 3995
rect 111 3980 115 3984
rect 151 3979 155 3983
rect 279 3979 283 3983
rect 431 3979 435 3983
rect 607 3979 611 3983
rect 791 3979 795 3983
rect 975 3979 979 3983
rect 1151 3979 1155 3983
rect 1311 3979 1315 3983
rect 1471 3979 1475 3983
rect 1623 3979 1627 3983
rect 1775 3979 1779 3983
rect 1903 3979 1907 3983
rect 2007 3980 2011 3984
rect 2047 3983 2051 3987
rect 2147 3987 2151 3991
rect 2071 3980 2075 3984
rect 3943 3983 3947 3987
rect 227 3971 231 3975
rect 355 3971 359 3975
rect 507 3971 511 3975
rect 683 3971 687 3975
rect 867 3971 871 3975
rect 919 3971 923 3975
rect 1227 3971 1231 3975
rect 1387 3971 1391 3975
rect 1547 3971 1551 3975
rect 1699 3971 1703 3975
rect 1851 3971 1855 3975
rect 1979 3971 1983 3975
rect 111 3963 115 3967
rect 151 3960 155 3964
rect 279 3960 283 3964
rect 431 3960 435 3964
rect 607 3960 611 3964
rect 791 3960 795 3964
rect 975 3960 979 3964
rect 1151 3960 1155 3964
rect 1311 3960 1315 3964
rect 1471 3960 1475 3964
rect 1623 3960 1627 3964
rect 1775 3960 1779 3964
rect 1903 3960 1907 3964
rect 2007 3963 2011 3967
rect 2047 3917 2051 3921
rect 2079 3920 2083 3924
rect 2215 3920 2219 3924
rect 2359 3920 2363 3924
rect 2503 3920 2507 3924
rect 2647 3920 2651 3924
rect 2791 3920 2795 3924
rect 2927 3920 2931 3924
rect 3055 3920 3059 3924
rect 3175 3920 3179 3924
rect 3295 3920 3299 3924
rect 3415 3920 3419 3924
rect 3535 3920 3539 3924
rect 3943 3917 3947 3921
rect 2155 3911 2159 3915
rect 2291 3911 2295 3915
rect 2435 3911 2439 3915
rect 2579 3911 2583 3915
rect 2715 3911 2719 3915
rect 2867 3911 2871 3915
rect 3003 3911 3007 3915
rect 3131 3911 3135 3915
rect 3251 3911 3255 3915
rect 3371 3911 3375 3915
rect 3491 3911 3495 3915
rect 3611 3911 3615 3915
rect 111 3897 115 3901
rect 303 3900 307 3904
rect 423 3900 427 3904
rect 551 3900 555 3904
rect 687 3900 691 3904
rect 815 3900 819 3904
rect 943 3900 947 3904
rect 1071 3900 1075 3904
rect 1199 3900 1203 3904
rect 1327 3900 1331 3904
rect 1463 3900 1467 3904
rect 2007 3897 2011 3901
rect 2047 3900 2051 3904
rect 2079 3901 2083 3905
rect 2215 3901 2219 3905
rect 2359 3901 2363 3905
rect 2503 3901 2507 3905
rect 2647 3901 2651 3905
rect 2791 3901 2795 3905
rect 2927 3901 2931 3905
rect 3055 3901 3059 3905
rect 3175 3901 3179 3905
rect 3295 3901 3299 3905
rect 3415 3901 3419 3905
rect 3535 3901 3539 3905
rect 3943 3900 3947 3904
rect 379 3891 383 3895
rect 499 3891 503 3895
rect 627 3891 631 3895
rect 763 3891 767 3895
rect 771 3891 775 3895
rect 1019 3891 1023 3895
rect 1147 3891 1151 3895
rect 1275 3891 1279 3895
rect 1403 3891 1407 3895
rect 1411 3891 1415 3895
rect 111 3880 115 3884
rect 303 3881 307 3885
rect 423 3881 427 3885
rect 551 3881 555 3885
rect 687 3881 691 3885
rect 815 3881 819 3885
rect 943 3881 947 3885
rect 1071 3881 1075 3885
rect 1199 3881 1203 3885
rect 1327 3881 1331 3885
rect 1463 3881 1467 3885
rect 2007 3880 2011 3884
rect 2147 3883 2151 3887
rect 2155 3883 2159 3887
rect 2291 3883 2295 3887
rect 2435 3883 2439 3887
rect 2579 3883 2583 3887
rect 2867 3883 2871 3887
rect 3003 3883 3007 3887
rect 3131 3883 3135 3887
rect 3251 3883 3255 3887
rect 3371 3883 3375 3887
rect 3491 3883 3495 3887
rect 919 3871 923 3875
rect 3079 3875 3083 3879
rect 379 3863 383 3867
rect 499 3863 503 3867
rect 627 3863 631 3867
rect 763 3863 767 3867
rect 983 3859 984 3863
rect 984 3859 987 3863
rect 1019 3863 1023 3867
rect 1147 3863 1151 3867
rect 1275 3863 1279 3867
rect 1403 3863 1407 3867
rect 2331 3867 2335 3871
rect 2459 3867 2463 3871
rect 2711 3867 2712 3871
rect 2712 3867 2715 3871
rect 2747 3867 2751 3871
rect 3027 3867 3028 3871
rect 3028 3867 3031 3871
rect 3067 3867 3071 3871
rect 3603 3867 3607 3871
rect 3611 3867 3615 3871
rect 2779 3859 2783 3863
rect 771 3851 775 3855
rect 2047 3848 2051 3852
rect 491 3843 495 3847
rect 643 3843 647 3847
rect 803 3843 807 3847
rect 1139 3843 1143 3847
rect 1275 3843 1279 3847
rect 1427 3843 1431 3847
rect 1563 3843 1567 3847
rect 1579 3843 1583 3847
rect 2255 3847 2259 3851
rect 2383 3847 2387 3851
rect 2519 3847 2523 3851
rect 2671 3847 2675 3851
rect 2831 3847 2835 3851
rect 2991 3847 2995 3851
rect 3159 3847 3163 3851
rect 3327 3847 3331 3851
rect 3495 3847 3499 3851
rect 3663 3847 3667 3851
rect 3943 3848 3947 3852
rect 2331 3839 2335 3843
rect 2459 3839 2463 3843
rect 2047 3831 2051 3835
rect 2595 3835 2599 3839
rect 2747 3839 2751 3843
rect 2779 3839 2783 3843
rect 3067 3839 3071 3843
rect 3079 3839 3083 3843
rect 3403 3835 3407 3839
rect 3603 3839 3607 3843
rect 111 3824 115 3828
rect 415 3823 419 3827
rect 567 3823 571 3827
rect 727 3823 731 3827
rect 887 3823 891 3827
rect 1039 3823 1043 3827
rect 1191 3823 1195 3827
rect 1343 3823 1347 3827
rect 1495 3823 1499 3827
rect 491 3815 495 3819
rect 643 3815 647 3819
rect 803 3815 807 3819
rect 859 3815 863 3819
rect 983 3815 987 3819
rect 1139 3815 1143 3819
rect 1275 3815 1279 3819
rect 1427 3815 1431 3819
rect 1563 3819 1567 3823
rect 1647 3823 1651 3827
rect 2007 3824 2011 3828
rect 2255 3828 2259 3832
rect 2383 3828 2387 3832
rect 2519 3828 2523 3832
rect 2671 3828 2675 3832
rect 2831 3828 2835 3832
rect 2991 3828 2995 3832
rect 3159 3828 3163 3832
rect 3327 3828 3331 3832
rect 3495 3828 3499 3832
rect 3663 3828 3667 3832
rect 3943 3831 3947 3835
rect 111 3807 115 3811
rect 415 3804 419 3808
rect 567 3804 571 3808
rect 727 3804 731 3808
rect 887 3804 891 3808
rect 1039 3804 1043 3808
rect 1191 3804 1195 3808
rect 1343 3804 1347 3808
rect 1495 3804 1499 3808
rect 1647 3804 1651 3808
rect 2007 3807 2011 3811
rect 2047 3765 2051 3769
rect 2071 3768 2075 3772
rect 2199 3768 2203 3772
rect 2375 3768 2379 3772
rect 2559 3768 2563 3772
rect 2751 3768 2755 3772
rect 2951 3768 2955 3772
rect 3143 3768 3147 3772
rect 3335 3768 3339 3772
rect 3535 3768 3539 3772
rect 3735 3768 3739 3772
rect 3943 3765 3947 3769
rect 2139 3759 2143 3763
rect 2303 3759 2307 3763
rect 2635 3759 2639 3763
rect 2643 3759 2647 3763
rect 3027 3759 3031 3763
rect 3047 3759 3051 3763
rect 3411 3759 3415 3763
rect 3611 3759 3615 3763
rect 3803 3759 3807 3763
rect 439 3751 443 3755
rect 859 3751 863 3755
rect 2047 3748 2051 3752
rect 2071 3749 2075 3753
rect 2199 3749 2203 3753
rect 2375 3749 2379 3753
rect 2559 3749 2563 3753
rect 2751 3749 2755 3753
rect 2951 3749 2955 3753
rect 3143 3749 3147 3753
rect 3335 3749 3339 3753
rect 3535 3749 3539 3753
rect 3735 3749 3739 3753
rect 3943 3748 3947 3752
rect 111 3737 115 3741
rect 399 3740 403 3744
rect 567 3740 571 3744
rect 751 3740 755 3744
rect 935 3740 939 3744
rect 1127 3740 1131 3744
rect 1311 3740 1315 3744
rect 1503 3740 1507 3744
rect 1695 3740 1699 3744
rect 1887 3740 1891 3744
rect 2007 3737 2011 3741
rect 475 3731 479 3735
rect 643 3731 647 3735
rect 827 3731 831 3735
rect 1011 3731 1015 3735
rect 1387 3731 1391 3735
rect 1579 3731 1583 3735
rect 1587 3731 1591 3735
rect 1799 3731 1803 3735
rect 2303 3731 2307 3735
rect 2643 3739 2647 3743
rect 2595 3731 2596 3735
rect 2596 3731 2599 3735
rect 2635 3731 2639 3735
rect 3047 3731 3051 3735
rect 3195 3727 3199 3731
rect 3403 3731 3407 3735
rect 3411 3731 3415 3735
rect 3611 3731 3615 3735
rect 111 3720 115 3724
rect 399 3721 403 3725
rect 567 3721 571 3725
rect 751 3721 755 3725
rect 935 3721 939 3725
rect 1127 3721 1131 3725
rect 1311 3721 1315 3725
rect 1503 3721 1507 3725
rect 1695 3721 1699 3725
rect 1887 3721 1891 3725
rect 2007 3720 2011 3724
rect 439 3703 440 3707
rect 440 3703 443 3707
rect 475 3703 479 3707
rect 643 3703 647 3707
rect 827 3703 831 3707
rect 1011 3703 1015 3707
rect 1587 3711 1591 3715
rect 1387 3703 1391 3707
rect 1799 3703 1803 3707
rect 1867 3699 1871 3703
rect 2139 3703 2143 3707
rect 2147 3703 2151 3707
rect 2339 3703 2343 3707
rect 2987 3703 2991 3707
rect 3395 3703 3399 3707
rect 3803 3703 3807 3707
rect 3019 3695 3023 3699
rect 3619 3695 3623 3699
rect 619 3683 623 3687
rect 1459 3683 1463 3687
rect 2047 3684 2051 3688
rect 2071 3683 2075 3687
rect 2263 3683 2267 3687
rect 2479 3683 2483 3687
rect 2695 3683 2699 3687
rect 2911 3683 2915 3687
rect 3119 3683 3123 3687
rect 3319 3683 3323 3687
rect 3519 3683 3523 3687
rect 3727 3683 3731 3687
rect 3943 3684 3947 3688
rect 443 3675 447 3679
rect 763 3675 767 3679
rect 1251 3675 1255 3679
rect 1403 3675 1407 3679
rect 1555 3675 1559 3679
rect 1707 3675 1711 3679
rect 2147 3675 2151 3679
rect 2339 3675 2343 3679
rect 2663 3675 2667 3679
rect 2987 3675 2991 3679
rect 3195 3675 3199 3679
rect 3395 3675 3399 3679
rect 2047 3667 2051 3671
rect 3595 3671 3599 3675
rect 3619 3675 3623 3679
rect 2071 3664 2075 3668
rect 2263 3664 2267 3668
rect 2479 3664 2483 3668
rect 2695 3664 2699 3668
rect 2911 3664 2915 3668
rect 3119 3664 3123 3668
rect 3319 3664 3323 3668
rect 3519 3664 3523 3668
rect 3727 3664 3731 3668
rect 3943 3667 3947 3671
rect 111 3656 115 3660
rect 367 3655 371 3659
rect 519 3655 523 3659
rect 679 3655 683 3659
rect 847 3655 851 3659
rect 1015 3655 1019 3659
rect 1175 3655 1179 3659
rect 1327 3655 1331 3659
rect 1479 3655 1483 3659
rect 1631 3655 1635 3659
rect 1791 3655 1795 3659
rect 2007 3656 2011 3660
rect 443 3647 447 3651
rect 111 3639 115 3643
rect 595 3643 599 3647
rect 619 3647 623 3651
rect 763 3647 767 3651
rect 1251 3647 1255 3651
rect 1403 3647 1407 3651
rect 1555 3647 1559 3651
rect 1707 3647 1711 3651
rect 1867 3647 1871 3651
rect 367 3636 371 3640
rect 519 3636 523 3640
rect 679 3636 683 3640
rect 847 3636 851 3640
rect 1015 3636 1019 3640
rect 1175 3636 1179 3640
rect 1327 3636 1331 3640
rect 1479 3636 1483 3640
rect 1631 3636 1635 3640
rect 1791 3636 1795 3640
rect 2007 3639 2011 3643
rect 2047 3597 2051 3601
rect 2111 3600 2115 3604
rect 2271 3600 2275 3604
rect 2455 3600 2459 3604
rect 2655 3600 2659 3604
rect 2871 3600 2875 3604
rect 3095 3600 3099 3604
rect 3327 3600 3331 3604
rect 3567 3600 3571 3604
rect 3943 3597 3947 3601
rect 2187 3591 2191 3595
rect 2347 3591 2351 3595
rect 2531 3591 2535 3595
rect 2731 3591 2735 3595
rect 2863 3591 2867 3595
rect 3019 3591 3023 3595
rect 3395 3591 3399 3595
rect 2047 3580 2051 3584
rect 2111 3581 2115 3585
rect 2271 3581 2275 3585
rect 2455 3581 2459 3585
rect 2655 3581 2659 3585
rect 2871 3581 2875 3585
rect 3095 3581 3099 3585
rect 3327 3581 3331 3585
rect 3567 3581 3571 3585
rect 3943 3580 3947 3584
rect 111 3565 115 3569
rect 271 3568 275 3572
rect 415 3568 419 3572
rect 575 3568 579 3572
rect 735 3568 739 3572
rect 895 3568 899 3572
rect 1055 3568 1059 3572
rect 1215 3568 1219 3572
rect 1375 3568 1379 3572
rect 1543 3568 1547 3572
rect 2007 3565 2011 3569
rect 347 3559 351 3563
rect 483 3559 487 3563
rect 651 3559 655 3563
rect 811 3559 815 3563
rect 819 3559 823 3563
rect 1131 3559 1135 3563
rect 1291 3559 1295 3563
rect 1451 3559 1455 3563
rect 1459 3559 1463 3563
rect 2663 3571 2667 3575
rect 2187 3563 2191 3567
rect 2347 3563 2351 3567
rect 2531 3563 2535 3567
rect 2731 3563 2735 3567
rect 3191 3559 3195 3563
rect 3595 3563 3599 3567
rect 111 3548 115 3552
rect 271 3549 275 3553
rect 415 3549 419 3553
rect 575 3549 579 3553
rect 735 3549 739 3553
rect 895 3549 899 3553
rect 1055 3549 1059 3553
rect 1215 3549 1219 3553
rect 1375 3549 1379 3553
rect 1543 3549 1547 3553
rect 2007 3548 2011 3552
rect 819 3539 823 3543
rect 347 3531 351 3535
rect 595 3531 599 3535
rect 651 3531 655 3535
rect 811 3531 815 3535
rect 1131 3535 1135 3539
rect 1291 3531 1295 3535
rect 1451 3531 1455 3535
rect 2355 3531 2359 3535
rect 2363 3531 2367 3535
rect 2467 3531 2471 3535
rect 2555 3531 2559 3535
rect 2739 3531 2743 3535
rect 2747 3531 2751 3535
rect 2843 3531 2847 3535
rect 2947 3531 2951 3535
rect 3059 3531 3063 3535
rect 3231 3531 3235 3535
rect 3391 3531 3392 3535
rect 3392 3531 3395 3535
rect 3427 3531 3431 3535
rect 1339 3523 1343 3527
rect 2047 3512 2051 3516
rect 235 3507 239 3511
rect 483 3507 487 3511
rect 499 3507 503 3511
rect 635 3507 639 3511
rect 883 3507 887 3511
rect 907 3507 911 3511
rect 1043 3507 1047 3511
rect 1171 3507 1175 3511
rect 1307 3507 1311 3511
rect 2287 3511 2291 3515
rect 2383 3511 2387 3515
rect 2479 3511 2483 3515
rect 2575 3511 2579 3515
rect 2671 3511 2675 3515
rect 2767 3511 2771 3515
rect 2871 3511 2875 3515
rect 2983 3511 2987 3515
rect 3103 3511 3107 3515
rect 3223 3511 3227 3515
rect 3351 3511 3355 3515
rect 3487 3511 3491 3515
rect 3943 3512 3947 3516
rect 643 3499 647 3503
rect 2363 3503 2367 3507
rect 2467 3503 2471 3507
rect 2555 3503 2559 3507
rect 2047 3495 2051 3499
rect 111 3488 115 3492
rect 159 3487 163 3491
rect 287 3487 291 3491
rect 423 3487 427 3491
rect 559 3487 563 3491
rect 695 3487 699 3491
rect 831 3487 835 3491
rect 967 3487 971 3491
rect 1095 3487 1099 3491
rect 1231 3487 1235 3491
rect 1367 3487 1371 3491
rect 2007 3488 2011 3492
rect 2287 3492 2291 3496
rect 2383 3492 2387 3496
rect 2479 3492 2483 3496
rect 2547 3495 2551 3499
rect 2747 3503 2751 3507
rect 2843 3503 2847 3507
rect 2947 3503 2951 3507
rect 3059 3503 3063 3507
rect 3067 3503 3071 3507
rect 3191 3503 3195 3507
rect 3427 3503 3431 3507
rect 3467 3503 3471 3507
rect 2575 3492 2579 3496
rect 2671 3492 2675 3496
rect 2767 3492 2771 3496
rect 2871 3492 2875 3496
rect 2983 3492 2987 3496
rect 3103 3492 3107 3496
rect 3223 3492 3227 3496
rect 3351 3492 3355 3496
rect 3487 3492 3491 3496
rect 3943 3495 3947 3499
rect 235 3479 239 3483
rect 111 3471 115 3475
rect 363 3475 367 3479
rect 499 3479 503 3483
rect 635 3479 639 3483
rect 643 3479 647 3483
rect 907 3479 911 3483
rect 1043 3479 1047 3483
rect 1171 3479 1175 3483
rect 1307 3479 1311 3483
rect 1339 3479 1343 3483
rect 159 3468 163 3472
rect 287 3468 291 3472
rect 423 3468 427 3472
rect 559 3468 563 3472
rect 695 3468 699 3472
rect 831 3468 835 3472
rect 967 3468 971 3472
rect 1095 3468 1099 3472
rect 1231 3468 1235 3472
rect 1367 3468 1371 3472
rect 2007 3471 2011 3475
rect 2047 3429 2051 3433
rect 2487 3432 2491 3436
rect 2583 3432 2587 3436
rect 2679 3432 2683 3436
rect 2783 3432 2787 3436
rect 2895 3432 2899 3436
rect 3015 3432 3019 3436
rect 3143 3432 3147 3436
rect 3271 3432 3275 3436
rect 3407 3432 3411 3436
rect 3943 3429 3947 3433
rect 2563 3423 2567 3427
rect 2659 3423 2663 3427
rect 2747 3423 2751 3427
rect 2887 3423 2891 3427
rect 2991 3423 2995 3427
rect 3231 3423 3235 3427
rect 3339 3423 3343 3427
rect 3379 3423 3383 3427
rect 2047 3412 2051 3416
rect 2487 3413 2491 3417
rect 2583 3413 2587 3417
rect 2679 3413 2683 3417
rect 2783 3413 2787 3417
rect 2895 3413 2899 3417
rect 3015 3413 3019 3417
rect 3143 3413 3147 3417
rect 3271 3413 3275 3417
rect 3407 3413 3411 3417
rect 3943 3412 3947 3416
rect 111 3397 115 3401
rect 135 3400 139 3404
rect 247 3400 251 3404
rect 383 3400 387 3404
rect 527 3400 531 3404
rect 671 3400 675 3404
rect 815 3400 819 3404
rect 967 3400 971 3404
rect 1119 3400 1123 3404
rect 1271 3400 1275 3404
rect 2007 3397 2011 3401
rect 203 3391 207 3395
rect 219 3391 223 3395
rect 459 3391 463 3395
rect 603 3391 607 3395
rect 611 3391 615 3395
rect 883 3391 887 3395
rect 903 3391 907 3395
rect 1195 3391 1199 3395
rect 1235 3391 1239 3395
rect 2547 3395 2551 3399
rect 2563 3395 2567 3399
rect 2659 3395 2663 3399
rect 2887 3395 2891 3399
rect 2991 3395 2995 3399
rect 3067 3395 3071 3399
rect 3099 3391 3103 3395
rect 3379 3395 3383 3399
rect 3467 3395 3471 3399
rect 111 3380 115 3384
rect 135 3381 139 3385
rect 247 3381 251 3385
rect 383 3381 387 3385
rect 527 3381 531 3385
rect 671 3381 675 3385
rect 815 3381 819 3385
rect 967 3381 971 3385
rect 1119 3381 1123 3385
rect 1271 3381 1275 3385
rect 2007 3380 2011 3384
rect 219 3363 223 3367
rect 611 3371 615 3375
rect 1235 3371 1239 3375
rect 2427 3371 2431 3375
rect 2555 3371 2559 3375
rect 2851 3371 2855 3375
rect 2963 3371 2967 3375
rect 3243 3371 3247 3375
rect 3339 3371 3340 3375
rect 3340 3371 3343 3375
rect 363 3363 367 3367
rect 459 3363 463 3367
rect 603 3363 607 3367
rect 903 3363 907 3367
rect 1159 3359 1160 3363
rect 1160 3359 1163 3363
rect 1195 3363 1199 3367
rect 2719 3363 2723 3367
rect 2047 3352 2051 3356
rect 2351 3351 2355 3355
rect 2479 3351 2483 3355
rect 2615 3351 2619 3355
rect 2751 3351 2755 3355
rect 2887 3351 2891 3355
rect 3023 3351 3027 3355
rect 3159 3351 3163 3355
rect 3303 3351 3307 3355
rect 3943 3352 3947 3356
rect 203 3339 207 3343
rect 211 3339 215 3343
rect 339 3339 343 3343
rect 507 3339 511 3343
rect 1003 3339 1007 3343
rect 1323 3339 1327 3343
rect 1475 3339 1479 3343
rect 1563 3339 1567 3343
rect 2427 3343 2431 3347
rect 2555 3343 2559 3347
rect 2719 3343 2723 3347
rect 2963 3343 2967 3347
rect 3099 3343 3103 3347
rect 1219 3331 1223 3335
rect 2047 3335 2051 3339
rect 2351 3332 2355 3336
rect 2479 3332 2483 3336
rect 2615 3332 2619 3336
rect 2683 3335 2687 3339
rect 3235 3339 3239 3343
rect 3243 3343 3247 3347
rect 2751 3332 2755 3336
rect 2887 3332 2891 3336
rect 3023 3332 3027 3336
rect 3159 3332 3163 3336
rect 3303 3332 3307 3336
rect 3943 3335 3947 3339
rect 111 3320 115 3324
rect 135 3319 139 3323
rect 263 3319 267 3323
rect 431 3319 435 3323
rect 599 3319 603 3323
rect 767 3319 771 3323
rect 927 3319 931 3323
rect 1087 3319 1091 3323
rect 1239 3319 1243 3323
rect 1391 3319 1395 3323
rect 1551 3319 1555 3323
rect 2007 3320 2011 3324
rect 211 3311 215 3315
rect 339 3311 343 3315
rect 507 3311 511 3315
rect 739 3311 743 3315
rect 1003 3311 1007 3315
rect 1163 3311 1167 3315
rect 1219 3311 1223 3315
rect 1323 3311 1327 3315
rect 1475 3311 1479 3315
rect 111 3303 115 3307
rect 135 3300 139 3304
rect 263 3300 267 3304
rect 431 3300 435 3304
rect 599 3300 603 3304
rect 767 3300 771 3304
rect 927 3300 931 3304
rect 1087 3300 1091 3304
rect 1239 3300 1243 3304
rect 1391 3300 1395 3304
rect 1551 3300 1555 3304
rect 2007 3303 2011 3307
rect 2047 3265 2051 3269
rect 2127 3268 2131 3272
rect 2295 3268 2299 3272
rect 2455 3268 2459 3272
rect 2615 3268 2619 3272
rect 2775 3268 2779 3272
rect 2935 3268 2939 3272
rect 3095 3268 3099 3272
rect 3263 3268 3267 3272
rect 3943 3265 3947 3269
rect 2215 3259 2219 3263
rect 2223 3259 2227 3263
rect 2399 3259 2403 3263
rect 2851 3259 2855 3263
rect 3023 3259 3027 3263
rect 3031 3259 3035 3263
rect 3179 3259 3183 3263
rect 2047 3248 2051 3252
rect 2127 3249 2131 3253
rect 2295 3249 2299 3253
rect 2455 3249 2459 3253
rect 2615 3249 2619 3253
rect 2775 3249 2779 3253
rect 2935 3249 2939 3253
rect 3095 3249 3099 3253
rect 3263 3249 3267 3253
rect 3943 3248 3947 3252
rect 111 3229 115 3233
rect 143 3232 147 3236
rect 295 3232 299 3236
rect 455 3232 459 3236
rect 623 3232 627 3236
rect 791 3232 795 3236
rect 959 3232 963 3236
rect 1127 3232 1131 3236
rect 1303 3232 1307 3236
rect 1479 3232 1483 3236
rect 2007 3229 2011 3233
rect 2223 3231 2227 3235
rect 2399 3231 2403 3235
rect 2683 3231 2687 3235
rect 219 3223 223 3227
rect 371 3223 375 3227
rect 531 3223 535 3227
rect 699 3223 703 3227
rect 1035 3223 1039 3227
rect 1203 3223 1207 3227
rect 1379 3223 1383 3227
rect 1563 3223 1567 3227
rect 3031 3231 3035 3235
rect 3179 3231 3183 3235
rect 3235 3231 3239 3235
rect 111 3212 115 3216
rect 143 3213 147 3217
rect 295 3213 299 3217
rect 455 3213 459 3217
rect 623 3213 627 3217
rect 791 3213 795 3217
rect 959 3213 963 3217
rect 1127 3213 1131 3217
rect 1303 3213 1307 3217
rect 1479 3213 1483 3217
rect 2007 3212 2011 3216
rect 2215 3215 2219 3219
rect 2283 3215 2287 3219
rect 2495 3215 2499 3219
rect 2715 3215 2719 3219
rect 2791 3215 2795 3219
rect 3023 3215 3027 3219
rect 3243 3215 3247 3219
rect 2503 3207 2507 3211
rect 183 3195 184 3199
rect 184 3195 187 3199
rect 219 3195 223 3199
rect 371 3195 375 3199
rect 531 3195 535 3199
rect 699 3195 703 3199
rect 1035 3199 1039 3203
rect 1203 3195 1207 3199
rect 1379 3195 1383 3199
rect 2047 3196 2051 3200
rect 2071 3195 2075 3199
rect 2207 3195 2211 3199
rect 2375 3195 2379 3199
rect 2543 3195 2547 3199
rect 2703 3195 2707 3199
rect 2863 3195 2867 3199
rect 3015 3195 3019 3199
rect 3167 3195 3171 3199
rect 3327 3195 3331 3199
rect 3943 3196 3947 3200
rect 1639 3187 1643 3191
rect 371 3179 375 3183
rect 507 3179 511 3183
rect 643 3179 647 3183
rect 923 3179 927 3183
rect 931 3179 935 3183
rect 1107 3179 1111 3183
rect 1383 3179 1387 3183
rect 1531 3179 1535 3183
rect 1963 3179 1967 3183
rect 2047 3179 2051 3183
rect 2147 3183 2151 3187
rect 2283 3187 2287 3191
rect 2495 3187 2499 3191
rect 2503 3187 2507 3191
rect 2791 3187 2795 3191
rect 3243 3187 3247 3191
rect 3403 3183 3407 3187
rect 2071 3176 2075 3180
rect 2207 3176 2211 3180
rect 2375 3176 2379 3180
rect 2543 3176 2547 3180
rect 2703 3176 2707 3180
rect 2863 3176 2867 3180
rect 3015 3176 3019 3180
rect 3167 3176 3171 3180
rect 3327 3176 3331 3180
rect 3943 3179 3947 3183
rect 111 3160 115 3164
rect 295 3159 299 3163
rect 431 3159 435 3163
rect 567 3159 571 3163
rect 703 3159 707 3163
rect 855 3159 859 3163
rect 1031 3159 1035 3163
rect 1231 3159 1235 3163
rect 1455 3159 1459 3163
rect 1687 3159 1691 3163
rect 1903 3159 1907 3163
rect 2007 3160 2011 3164
rect 371 3151 375 3155
rect 507 3151 511 3155
rect 643 3151 647 3155
rect 651 3151 655 3155
rect 931 3151 935 3155
rect 1107 3151 1111 3155
rect 1383 3151 1387 3155
rect 1531 3151 1535 3155
rect 1639 3151 1643 3155
rect 111 3143 115 3147
rect 295 3140 299 3144
rect 431 3140 435 3144
rect 567 3140 571 3144
rect 703 3140 707 3144
rect 855 3140 859 3144
rect 1031 3140 1035 3144
rect 1231 3140 1235 3144
rect 1455 3140 1459 3144
rect 1687 3140 1691 3144
rect 1903 3140 1907 3144
rect 1971 3143 1975 3147
rect 2007 3143 2011 3147
rect 2047 3109 2051 3113
rect 2071 3112 2075 3116
rect 2343 3112 2347 3116
rect 2631 3112 2635 3116
rect 2903 3112 2907 3116
rect 3175 3112 3179 3116
rect 3447 3112 3451 3116
rect 3943 3109 3947 3113
rect 351 3099 355 3103
rect 651 3099 655 3103
rect 1963 3103 1967 3107
rect 2419 3103 2423 3107
rect 2715 3103 2719 3107
rect 2991 3103 2995 3107
rect 3007 3103 3011 3107
rect 3259 3103 3263 3107
rect 2047 3092 2051 3096
rect 2071 3093 2075 3097
rect 2343 3093 2347 3097
rect 2631 3093 2635 3097
rect 2903 3093 2907 3097
rect 3175 3093 3179 3097
rect 3447 3093 3451 3097
rect 3943 3092 3947 3096
rect 923 3087 927 3091
rect 111 3077 115 3081
rect 311 3080 315 3084
rect 407 3080 411 3084
rect 503 3080 507 3084
rect 599 3080 603 3084
rect 695 3080 699 3084
rect 807 3080 811 3084
rect 943 3080 947 3084
rect 1087 3080 1091 3084
rect 1247 3080 1251 3084
rect 387 3071 391 3075
rect 483 3071 487 3075
rect 579 3071 583 3075
rect 675 3071 679 3075
rect 771 3071 775 3075
rect 779 3071 783 3075
rect 1019 3071 1023 3075
rect 1163 3071 1167 3075
rect 1323 3071 1327 3075
rect 1407 3080 1411 3084
rect 1575 3080 1579 3084
rect 1751 3080 1755 3084
rect 1903 3080 1907 3084
rect 2007 3077 2011 3081
rect 1651 3071 1655 3075
rect 1827 3071 1831 3075
rect 1835 3071 1839 3075
rect 2147 3075 2151 3079
rect 2419 3075 2423 3079
rect 3007 3075 3011 3079
rect 3259 3075 3263 3079
rect 3403 3075 3407 3079
rect 2827 3067 2831 3071
rect 111 3060 115 3064
rect 311 3061 315 3065
rect 407 3061 411 3065
rect 503 3061 507 3065
rect 599 3061 603 3065
rect 695 3061 699 3065
rect 807 3061 811 3065
rect 943 3061 947 3065
rect 1087 3061 1091 3065
rect 1247 3061 1251 3065
rect 1407 3061 1411 3065
rect 1575 3061 1579 3065
rect 1751 3061 1755 3065
rect 1903 3061 1907 3065
rect 2007 3060 2011 3064
rect 351 3043 352 3047
rect 352 3043 355 3047
rect 387 3043 391 3047
rect 483 3043 487 3047
rect 579 3043 583 3047
rect 675 3043 679 3047
rect 771 3043 775 3047
rect 1019 3043 1023 3047
rect 1163 3043 1167 3047
rect 1323 3043 1327 3047
rect 1835 3051 1839 3055
rect 2495 3055 2499 3059
rect 2563 3055 2567 3059
rect 2691 3055 2695 3059
rect 2819 3055 2823 3059
rect 2991 3055 2995 3059
rect 3059 3055 3063 3059
rect 3199 3055 3203 3059
rect 3291 3055 3295 3059
rect 3403 3055 3407 3059
rect 3603 3055 3607 3059
rect 3611 3055 3615 3059
rect 3715 3055 3719 3059
rect 3819 3055 3823 3059
rect 1651 3043 1655 3047
rect 1971 3043 1975 3047
rect 1279 3035 1283 3039
rect 2047 3036 2051 3040
rect 2487 3035 2491 3039
rect 2615 3035 2619 3039
rect 2743 3035 2747 3039
rect 2863 3035 2867 3039
rect 2983 3035 2987 3039
rect 3103 3035 3107 3039
rect 3215 3035 3219 3039
rect 3327 3035 3331 3039
rect 3431 3035 3435 3039
rect 3535 3035 3539 3039
rect 3639 3035 3643 3039
rect 3743 3035 3747 3039
rect 3839 3035 3843 3039
rect 3943 3036 3947 3040
rect 463 3027 464 3031
rect 464 3027 467 3031
rect 511 3027 515 3031
rect 607 3027 611 3031
rect 703 3027 707 3031
rect 787 3027 791 3031
rect 891 3027 895 3031
rect 1011 3027 1015 3031
rect 1131 3027 1135 3031
rect 1259 3027 1263 3031
rect 1515 3027 1519 3031
rect 1635 3027 1639 3031
rect 1827 3027 1831 3031
rect 1875 3027 1879 3031
rect 2563 3027 2567 3031
rect 2691 3027 2695 3031
rect 2819 3027 2823 3031
rect 2827 3027 2831 3031
rect 3059 3027 3063 3031
rect 3199 3027 3203 3031
rect 3291 3027 3295 3031
rect 3403 3027 3407 3031
rect 3611 3027 3615 3031
rect 3715 3027 3719 3031
rect 3819 3027 3823 3031
rect 1883 3019 1887 3023
rect 2047 3019 2051 3023
rect 2487 3016 2491 3020
rect 2615 3016 2619 3020
rect 2743 3016 2747 3020
rect 2863 3016 2867 3020
rect 2983 3016 2987 3020
rect 3103 3016 3107 3020
rect 3215 3016 3219 3020
rect 3327 3016 3331 3020
rect 3431 3016 3435 3020
rect 3535 3016 3539 3020
rect 3639 3016 3643 3020
rect 3743 3016 3747 3020
rect 3839 3016 3843 3020
rect 3907 3019 3911 3023
rect 3943 3019 3947 3023
rect 111 3008 115 3012
rect 423 3007 427 3011
rect 519 3007 523 3011
rect 615 3007 619 3011
rect 711 3007 715 3011
rect 815 3007 819 3011
rect 935 3007 939 3011
rect 1055 3007 1059 3011
rect 1183 3007 1187 3011
rect 1311 3007 1315 3011
rect 1431 3007 1435 3011
rect 1551 3007 1555 3011
rect 1671 3007 1675 3011
rect 1799 3007 1803 3011
rect 1903 3007 1907 3011
rect 2007 3008 2011 3012
rect 511 2999 515 3003
rect 607 2999 611 3003
rect 703 2999 707 3003
rect 787 2999 791 3003
rect 891 2999 895 3003
rect 1011 2999 1015 3003
rect 1131 2999 1135 3003
rect 1259 2999 1263 3003
rect 1279 2999 1283 3003
rect 111 2991 115 2995
rect 1507 2995 1511 2999
rect 1515 2999 1519 3003
rect 1635 2999 1639 3003
rect 1875 2999 1879 3003
rect 1883 2999 1887 3003
rect 423 2988 427 2992
rect 519 2988 523 2992
rect 615 2988 619 2992
rect 711 2988 715 2992
rect 815 2988 819 2992
rect 935 2988 939 2992
rect 1055 2988 1059 2992
rect 1183 2988 1187 2992
rect 1311 2988 1315 2992
rect 1431 2988 1435 2992
rect 1551 2988 1555 2992
rect 1671 2988 1675 2992
rect 1799 2988 1803 2992
rect 1903 2988 1907 2992
rect 2007 2991 2011 2995
rect 2047 2949 2051 2953
rect 2407 2952 2411 2956
rect 2575 2952 2579 2956
rect 2767 2952 2771 2956
rect 2967 2952 2971 2956
rect 3183 2952 3187 2956
rect 3399 2952 3403 2956
rect 3623 2952 3627 2956
rect 3839 2952 3843 2956
rect 3943 2949 3947 2953
rect 2495 2943 2499 2947
rect 2503 2943 2507 2947
rect 2695 2943 2699 2947
rect 2923 2943 2927 2947
rect 3115 2943 3119 2947
rect 3475 2943 3479 2947
rect 3603 2943 3607 2947
rect 3915 2943 3919 2947
rect 2047 2932 2051 2936
rect 2407 2933 2411 2937
rect 2575 2933 2579 2937
rect 2767 2933 2771 2937
rect 2967 2933 2971 2937
rect 3183 2933 3187 2937
rect 3399 2933 3403 2937
rect 3623 2933 3627 2937
rect 3839 2933 3843 2937
rect 3943 2932 3947 2936
rect 2503 2915 2507 2919
rect 2695 2915 2699 2919
rect 2923 2915 2927 2919
rect 3115 2915 3119 2919
rect 3131 2911 3135 2915
rect 3475 2915 3479 2919
rect 3907 2915 3911 2919
rect 111 2901 115 2905
rect 1479 2904 1483 2908
rect 1575 2904 1579 2908
rect 1671 2904 1675 2908
rect 1767 2904 1771 2908
rect 1863 2904 1867 2908
rect 2007 2901 2011 2905
rect 1555 2895 1559 2899
rect 1651 2895 1655 2899
rect 1747 2895 1751 2899
rect 1843 2895 1847 2899
rect 1931 2895 1935 2899
rect 111 2884 115 2888
rect 1479 2885 1483 2889
rect 1575 2885 1579 2889
rect 1671 2885 1675 2889
rect 1767 2885 1771 2889
rect 1863 2885 1867 2889
rect 2007 2884 2011 2888
rect 2627 2883 2631 2887
rect 2747 2883 2751 2887
rect 2875 2883 2879 2887
rect 3003 2883 3007 2887
rect 3267 2883 3271 2887
rect 3467 2883 3471 2887
rect 3515 2883 3519 2887
rect 2915 2875 2919 2879
rect 3523 2875 3527 2879
rect 1507 2867 1511 2871
rect 1555 2867 1559 2871
rect 1651 2867 1655 2871
rect 1747 2867 1751 2871
rect 1843 2867 1847 2871
rect 2047 2864 2051 2868
rect 2551 2863 2555 2867
rect 2671 2863 2675 2867
rect 2799 2863 2803 2867
rect 2927 2863 2931 2867
rect 3055 2863 3059 2867
rect 3183 2863 3187 2867
rect 3311 2863 3315 2867
rect 3439 2863 3443 2867
rect 3575 2863 3579 2867
rect 3943 2864 3947 2868
rect 2627 2855 2631 2859
rect 2747 2855 2751 2859
rect 2875 2855 2879 2859
rect 3003 2855 3007 2859
rect 3131 2855 3135 2859
rect 3143 2855 3147 2859
rect 3267 2855 3271 2859
rect 3515 2855 3519 2859
rect 3523 2855 3527 2859
rect 355 2847 359 2851
rect 439 2839 443 2843
rect 523 2843 527 2847
rect 707 2843 711 2847
rect 891 2843 895 2847
rect 1259 2843 1263 2847
rect 1611 2843 1615 2847
rect 1779 2843 1783 2847
rect 1931 2843 1935 2847
rect 2047 2847 2051 2851
rect 2551 2844 2555 2848
rect 2671 2844 2675 2848
rect 2799 2844 2803 2848
rect 2927 2844 2931 2848
rect 3055 2844 3059 2848
rect 3183 2844 3187 2848
rect 3311 2844 3315 2848
rect 3439 2844 3443 2848
rect 3575 2844 3579 2848
rect 3943 2847 3947 2851
rect 1459 2835 1463 2839
rect 111 2824 115 2828
rect 279 2823 283 2827
rect 447 2823 451 2827
rect 631 2823 635 2827
rect 815 2823 819 2827
rect 999 2823 1003 2827
rect 1183 2823 1187 2827
rect 1359 2823 1363 2827
rect 1527 2823 1531 2827
rect 1695 2823 1699 2827
rect 1863 2823 1867 2827
rect 2007 2824 2011 2828
rect 355 2815 359 2819
rect 523 2815 527 2819
rect 707 2815 711 2819
rect 891 2815 895 2819
rect 967 2815 971 2819
rect 1259 2815 1263 2819
rect 111 2807 115 2811
rect 1435 2811 1439 2815
rect 1459 2815 1463 2819
rect 1611 2815 1615 2819
rect 1779 2815 1783 2819
rect 279 2804 283 2808
rect 447 2804 451 2808
rect 631 2804 635 2808
rect 815 2804 819 2808
rect 999 2804 1003 2808
rect 1183 2804 1187 2808
rect 1359 2804 1363 2808
rect 1527 2804 1531 2808
rect 1695 2804 1699 2808
rect 1863 2804 1867 2808
rect 2007 2807 2011 2811
rect 2047 2781 2051 2785
rect 2439 2784 2443 2788
rect 2567 2784 2571 2788
rect 2695 2784 2699 2788
rect 2831 2784 2835 2788
rect 2967 2784 2971 2788
rect 3103 2784 3107 2788
rect 3247 2784 3251 2788
rect 3391 2784 3395 2788
rect 3543 2784 3547 2788
rect 3703 2784 3707 2788
rect 3839 2784 3843 2788
rect 3943 2781 3947 2785
rect 2515 2775 2519 2779
rect 2643 2775 2647 2779
rect 2771 2775 2775 2779
rect 2907 2775 2911 2779
rect 2915 2775 2919 2779
rect 3179 2775 3183 2779
rect 3323 2775 3327 2779
rect 3467 2775 3471 2779
rect 3475 2775 3479 2779
rect 3631 2775 3635 2779
rect 3907 2775 3911 2779
rect 2047 2764 2051 2768
rect 2439 2765 2443 2769
rect 2567 2765 2571 2769
rect 2695 2765 2699 2769
rect 2831 2765 2835 2769
rect 2967 2765 2971 2769
rect 3103 2765 3107 2769
rect 3247 2765 3251 2769
rect 3391 2765 3395 2769
rect 3543 2765 3547 2769
rect 3703 2765 3707 2769
rect 3839 2765 3843 2769
rect 3943 2764 3947 2768
rect 111 2741 115 2745
rect 239 2744 243 2748
rect 351 2744 355 2748
rect 471 2744 475 2748
rect 607 2744 611 2748
rect 743 2744 747 2748
rect 879 2744 883 2748
rect 1015 2744 1019 2748
rect 1151 2744 1155 2748
rect 1287 2744 1291 2748
rect 1423 2744 1427 2748
rect 1567 2744 1571 2748
rect 2007 2741 2011 2745
rect 2515 2747 2519 2751
rect 2643 2747 2647 2751
rect 2771 2747 2775 2751
rect 2907 2747 2911 2751
rect 3143 2747 3144 2751
rect 3144 2747 3147 2751
rect 3179 2747 3183 2751
rect 3475 2747 3479 2751
rect 3631 2747 3635 2751
rect 315 2735 319 2739
rect 427 2735 431 2739
rect 439 2735 443 2739
rect 555 2735 559 2739
rect 727 2735 731 2739
rect 851 2735 855 2739
rect 1091 2735 1095 2739
rect 1239 2735 1243 2739
rect 1247 2735 1251 2739
rect 1499 2735 1503 2739
rect 1507 2735 1511 2739
rect 3763 2743 3767 2747
rect 3915 2747 3919 2751
rect 111 2724 115 2728
rect 239 2725 243 2729
rect 351 2725 355 2729
rect 471 2725 475 2729
rect 607 2725 611 2729
rect 743 2725 747 2729
rect 879 2725 883 2729
rect 1015 2725 1019 2729
rect 1151 2725 1155 2729
rect 1287 2725 1291 2729
rect 1423 2725 1427 2729
rect 1567 2725 1571 2729
rect 2007 2724 2011 2728
rect 2403 2723 2407 2727
rect 2411 2723 2415 2727
rect 2739 2723 2743 2727
rect 3075 2723 3079 2727
rect 3323 2723 3327 2727
rect 3579 2723 3583 2727
rect 3587 2723 3591 2727
rect 3907 2723 3911 2727
rect 299 2703 303 2707
rect 315 2707 319 2711
rect 427 2707 431 2711
rect 727 2707 731 2711
rect 851 2707 855 2711
rect 967 2707 971 2711
rect 1247 2715 1251 2719
rect 1091 2707 1095 2711
rect 1507 2715 1511 2719
rect 3259 2715 3263 2719
rect 1435 2707 1439 2711
rect 1499 2707 1503 2711
rect 2047 2704 2051 2708
rect 2335 2703 2339 2707
rect 2495 2703 2499 2707
rect 2663 2703 2667 2707
rect 2831 2703 2835 2707
rect 2999 2703 3003 2707
rect 3167 2703 3171 2707
rect 3335 2703 3339 2707
rect 3511 2703 3515 2707
rect 3687 2703 3691 2707
rect 3839 2703 3843 2707
rect 3943 2704 3947 2708
rect 307 2691 311 2695
rect 435 2691 439 2695
rect 555 2691 559 2695
rect 579 2691 583 2695
rect 715 2691 719 2695
rect 971 2691 975 2695
rect 1083 2691 1087 2695
rect 1239 2691 1243 2695
rect 1307 2691 1311 2695
rect 2411 2695 2415 2699
rect 2739 2695 2743 2699
rect 3075 2695 3079 2699
rect 1315 2683 1319 2687
rect 2047 2687 2051 2691
rect 3243 2691 3247 2695
rect 3259 2695 3263 2699
rect 3587 2695 3591 2699
rect 3763 2695 3767 2699
rect 2335 2684 2339 2688
rect 2495 2684 2499 2688
rect 2663 2684 2667 2688
rect 2831 2684 2835 2688
rect 2999 2684 3003 2688
rect 3167 2684 3171 2688
rect 3335 2684 3339 2688
rect 3511 2684 3515 2688
rect 3687 2684 3691 2688
rect 3839 2684 3843 2688
rect 3907 2687 3911 2691
rect 3943 2687 3947 2691
rect 111 2672 115 2676
rect 223 2671 227 2675
rect 367 2671 371 2675
rect 503 2671 507 2675
rect 639 2671 643 2675
rect 767 2671 771 2675
rect 887 2671 891 2675
rect 999 2671 1003 2675
rect 1111 2671 1115 2675
rect 1231 2671 1235 2675
rect 1351 2671 1355 2675
rect 2007 2672 2011 2676
rect 299 2663 303 2667
rect 307 2663 311 2667
rect 579 2663 583 2667
rect 715 2663 719 2667
rect 751 2663 755 2667
rect 879 2663 883 2667
rect 971 2663 975 2667
rect 1083 2663 1087 2667
rect 1307 2663 1311 2667
rect 1315 2663 1319 2667
rect 111 2655 115 2659
rect 223 2652 227 2656
rect 367 2652 371 2656
rect 503 2652 507 2656
rect 639 2652 643 2656
rect 767 2652 771 2656
rect 887 2652 891 2656
rect 999 2652 1003 2656
rect 1111 2652 1115 2656
rect 1231 2652 1235 2656
rect 1351 2652 1355 2656
rect 2007 2655 2011 2659
rect 2403 2627 2407 2631
rect 2047 2617 2051 2621
rect 2127 2620 2131 2624
rect 2279 2620 2283 2624
rect 2447 2620 2451 2624
rect 2623 2620 2627 2624
rect 2203 2611 2207 2615
rect 2355 2611 2359 2615
rect 2523 2611 2527 2615
rect 2699 2611 2703 2615
rect 2807 2620 2811 2624
rect 2991 2620 2995 2624
rect 3175 2620 3179 2624
rect 3351 2620 3355 2624
rect 3519 2620 3523 2624
rect 3687 2620 3691 2624
rect 3839 2620 3843 2624
rect 3943 2617 3947 2621
rect 2891 2611 2895 2615
rect 3103 2611 3107 2615
rect 3427 2611 3431 2615
rect 3587 2611 3591 2615
rect 3619 2611 3623 2615
rect 3923 2611 3927 2615
rect 2047 2600 2051 2604
rect 2127 2601 2131 2605
rect 2279 2601 2283 2605
rect 2447 2601 2451 2605
rect 2623 2601 2627 2605
rect 2807 2601 2811 2605
rect 2991 2601 2995 2605
rect 3175 2601 3179 2605
rect 3351 2601 3355 2605
rect 3519 2601 3523 2605
rect 3687 2601 3691 2605
rect 3839 2601 3843 2605
rect 3943 2600 3947 2604
rect 111 2589 115 2593
rect 175 2592 179 2596
rect 367 2592 371 2596
rect 543 2592 547 2596
rect 711 2592 715 2596
rect 863 2592 867 2596
rect 1007 2592 1011 2596
rect 1143 2592 1147 2596
rect 1279 2592 1283 2596
rect 1423 2592 1427 2596
rect 2007 2589 2011 2593
rect 251 2583 255 2587
rect 435 2583 439 2587
rect 619 2583 623 2587
rect 631 2583 635 2587
rect 939 2583 943 2587
rect 1083 2583 1087 2587
rect 1219 2583 1223 2587
rect 1355 2583 1359 2587
rect 1367 2583 1371 2587
rect 2167 2579 2168 2583
rect 2168 2579 2171 2583
rect 2203 2583 2207 2587
rect 2355 2583 2359 2587
rect 2523 2583 2527 2587
rect 2699 2583 2703 2587
rect 3103 2583 3107 2587
rect 3243 2583 3247 2587
rect 3619 2591 3623 2595
rect 3427 2583 3431 2587
rect 3727 2579 3728 2583
rect 3728 2579 3731 2583
rect 3907 2583 3911 2587
rect 111 2572 115 2576
rect 175 2573 179 2577
rect 367 2573 371 2577
rect 543 2573 547 2577
rect 711 2573 715 2577
rect 863 2573 867 2577
rect 1007 2573 1011 2577
rect 1143 2573 1147 2577
rect 1279 2573 1283 2577
rect 1423 2573 1427 2577
rect 2007 2572 2011 2576
rect 211 2551 212 2555
rect 212 2551 215 2555
rect 251 2555 255 2559
rect 631 2555 635 2559
rect 751 2555 752 2559
rect 752 2555 755 2559
rect 879 2555 883 2559
rect 939 2555 943 2559
rect 1083 2555 1087 2559
rect 1219 2555 1223 2559
rect 1355 2555 1359 2559
rect 2147 2559 2151 2563
rect 2259 2559 2263 2563
rect 2395 2559 2399 2563
rect 2547 2559 2551 2563
rect 2891 2559 2895 2563
rect 2899 2559 2903 2563
rect 3107 2559 3111 2563
rect 3339 2559 3343 2563
rect 3699 2559 3703 2563
rect 2299 2551 2303 2555
rect 1367 2543 1371 2547
rect 219 2535 223 2539
rect 355 2535 359 2539
rect 479 2535 480 2539
rect 480 2535 483 2539
rect 619 2535 623 2539
rect 683 2535 687 2539
rect 851 2535 855 2539
rect 2047 2540 2051 2544
rect 1155 2535 1159 2539
rect 1299 2535 1303 2539
rect 1435 2535 1439 2539
rect 1571 2535 1575 2539
rect 2071 2539 2075 2543
rect 2183 2539 2187 2543
rect 2319 2539 2323 2543
rect 2471 2539 2475 2543
rect 2639 2539 2643 2543
rect 2823 2539 2827 2543
rect 3031 2539 3035 2543
rect 3263 2539 3267 2543
rect 3503 2539 3507 2543
rect 3743 2539 3747 2543
rect 3943 2540 3947 2544
rect 2147 2531 2151 2535
rect 2259 2531 2263 2535
rect 2395 2531 2399 2535
rect 2547 2531 2551 2535
rect 2599 2531 2603 2535
rect 2899 2531 2903 2535
rect 3107 2531 3111 2535
rect 3339 2531 3343 2535
rect 3451 2531 3455 2535
rect 3727 2531 3731 2535
rect 2047 2523 2051 2527
rect 111 2516 115 2520
rect 135 2515 139 2519
rect 271 2515 275 2519
rect 439 2515 443 2519
rect 607 2515 611 2519
rect 775 2515 779 2519
rect 927 2515 931 2519
rect 1079 2515 1083 2519
rect 1223 2515 1227 2519
rect 1359 2515 1363 2519
rect 1495 2515 1499 2519
rect 1639 2515 1643 2519
rect 2007 2516 2011 2520
rect 2071 2520 2075 2524
rect 2183 2520 2187 2524
rect 2319 2520 2323 2524
rect 2471 2520 2475 2524
rect 2639 2520 2643 2524
rect 2823 2520 2827 2524
rect 3031 2520 3035 2524
rect 3263 2520 3267 2524
rect 3503 2520 3507 2524
rect 3743 2520 3747 2524
rect 3943 2523 3947 2527
rect 211 2507 215 2511
rect 219 2507 223 2511
rect 355 2507 359 2511
rect 683 2507 687 2511
rect 851 2507 855 2511
rect 111 2499 115 2503
rect 1003 2503 1007 2507
rect 1155 2507 1159 2511
rect 1299 2507 1303 2511
rect 1435 2507 1439 2511
rect 1571 2507 1575 2511
rect 1579 2507 1583 2511
rect 135 2496 139 2500
rect 271 2496 275 2500
rect 439 2496 443 2500
rect 607 2496 611 2500
rect 775 2496 779 2500
rect 927 2496 931 2500
rect 1079 2496 1083 2500
rect 1223 2496 1227 2500
rect 1359 2496 1363 2500
rect 1495 2496 1499 2500
rect 1639 2496 1643 2500
rect 2007 2499 2011 2503
rect 2047 2453 2051 2457
rect 2071 2456 2075 2460
rect 2215 2456 2219 2460
rect 2383 2456 2387 2460
rect 2559 2456 2563 2460
rect 2751 2456 2755 2460
rect 2951 2456 2955 2460
rect 3167 2456 3171 2460
rect 3391 2456 3395 2460
rect 3623 2456 3627 2460
rect 3839 2456 3843 2460
rect 3943 2453 3947 2457
rect 2147 2447 2151 2451
rect 2291 2447 2295 2451
rect 2299 2447 2303 2451
rect 2471 2447 2475 2451
rect 2643 2447 2647 2451
rect 2899 2447 2903 2451
rect 3035 2447 3039 2451
rect 3699 2447 3703 2451
rect 3907 2447 3911 2451
rect 111 2429 115 2433
rect 135 2432 139 2436
rect 311 2432 315 2436
rect 511 2432 515 2436
rect 711 2432 715 2436
rect 903 2432 907 2436
rect 1079 2432 1083 2436
rect 1239 2432 1243 2436
rect 1391 2432 1395 2436
rect 1527 2432 1531 2436
rect 1663 2432 1667 2436
rect 1791 2432 1795 2436
rect 1903 2432 1907 2436
rect 2047 2436 2051 2440
rect 2071 2437 2075 2441
rect 2215 2437 2219 2441
rect 2383 2437 2387 2441
rect 2559 2437 2563 2441
rect 2751 2437 2755 2441
rect 2951 2437 2955 2441
rect 3167 2437 3171 2441
rect 3391 2437 3395 2441
rect 3623 2437 3627 2441
rect 3839 2437 3843 2441
rect 3943 2436 3947 2440
rect 2007 2429 2011 2433
rect 211 2423 215 2427
rect 387 2423 391 2427
rect 479 2423 483 2427
rect 619 2423 623 2427
rect 847 2423 851 2427
rect 1155 2423 1159 2427
rect 1315 2423 1319 2427
rect 1467 2423 1471 2427
rect 1475 2423 1479 2427
rect 1739 2423 1743 2427
rect 1867 2423 1871 2427
rect 2147 2419 2151 2423
rect 2291 2419 2295 2423
rect 2643 2419 2647 2423
rect 2899 2419 2903 2423
rect 3035 2419 3039 2423
rect 3451 2419 3455 2423
rect 111 2412 115 2416
rect 135 2413 139 2417
rect 311 2413 315 2417
rect 511 2413 515 2417
rect 711 2413 715 2417
rect 903 2413 907 2417
rect 1079 2413 1083 2417
rect 1239 2413 1243 2417
rect 1391 2413 1395 2417
rect 1527 2413 1531 2417
rect 1663 2413 1667 2417
rect 1791 2413 1795 2417
rect 1903 2413 1907 2417
rect 2007 2412 2011 2416
rect 3747 2415 3751 2419
rect 3923 2419 3927 2423
rect 211 2395 215 2399
rect 387 2395 391 2399
rect 847 2395 851 2399
rect 1003 2395 1007 2399
rect 1579 2403 1583 2407
rect 1155 2395 1159 2399
rect 1315 2395 1319 2399
rect 1467 2395 1471 2399
rect 211 2387 215 2391
rect 1475 2387 1479 2391
rect 1739 2395 1743 2399
rect 1867 2395 1871 2399
rect 1819 2387 1823 2391
rect 2155 2387 2159 2391
rect 2259 2387 2263 2391
rect 2471 2387 2472 2391
rect 2472 2387 2475 2391
rect 2507 2387 2511 2391
rect 2683 2387 2687 2391
rect 2851 2387 2855 2391
rect 3011 2387 3015 2391
rect 247 2379 251 2383
rect 347 2379 351 2383
rect 619 2379 623 2383
rect 627 2379 631 2383
rect 843 2379 847 2383
rect 1251 2379 1255 2383
rect 1443 2379 1447 2383
rect 1627 2379 1631 2383
rect 2055 2379 2059 2383
rect 2047 2368 2051 2372
rect 2071 2367 2075 2371
rect 2247 2367 2251 2371
rect 2431 2367 2435 2371
rect 2607 2367 2611 2371
rect 2775 2367 2779 2371
rect 2935 2367 2939 2371
rect 3103 2367 3107 2371
rect 3943 2368 3947 2372
rect 111 2360 115 2364
rect 135 2359 139 2363
rect 327 2359 331 2363
rect 551 2359 555 2363
rect 767 2359 771 2363
rect 975 2359 979 2363
rect 1175 2359 1179 2363
rect 1367 2359 1371 2363
rect 1551 2359 1555 2363
rect 1735 2359 1739 2363
rect 1903 2359 1907 2363
rect 2007 2360 2011 2364
rect 2055 2359 2059 2363
rect 2155 2359 2159 2363
rect 2507 2359 2511 2363
rect 2683 2359 2687 2363
rect 2851 2359 2855 2363
rect 3011 2359 3015 2363
rect 3019 2359 3023 2363
rect 211 2351 215 2355
rect 247 2351 251 2355
rect 627 2351 631 2355
rect 843 2351 847 2355
rect 967 2351 971 2355
rect 1251 2351 1255 2355
rect 1443 2351 1447 2355
rect 1627 2351 1631 2355
rect 1671 2351 1675 2355
rect 1819 2351 1823 2355
rect 2047 2351 2051 2355
rect 2071 2348 2075 2352
rect 111 2343 115 2347
rect 2247 2348 2251 2352
rect 2431 2348 2435 2352
rect 2607 2348 2611 2352
rect 2775 2348 2779 2352
rect 2935 2348 2939 2352
rect 3103 2348 3107 2352
rect 3943 2351 3947 2355
rect 135 2340 139 2344
rect 327 2340 331 2344
rect 551 2340 555 2344
rect 767 2340 771 2344
rect 975 2340 979 2344
rect 1175 2340 1179 2344
rect 1367 2340 1371 2344
rect 1551 2340 1555 2344
rect 1735 2340 1739 2344
rect 1903 2340 1907 2344
rect 2007 2343 2011 2347
rect 2047 2285 2051 2289
rect 2071 2288 2075 2292
rect 2175 2288 2179 2292
rect 2311 2288 2315 2292
rect 2447 2288 2451 2292
rect 2591 2288 2595 2292
rect 2751 2288 2755 2292
rect 2935 2288 2939 2292
rect 3143 2288 3147 2292
rect 3375 2288 3379 2292
rect 3615 2288 3619 2292
rect 3839 2288 3843 2292
rect 3943 2285 3947 2289
rect 2147 2279 2151 2283
rect 2259 2279 2263 2283
rect 2267 2279 2271 2283
rect 2523 2279 2527 2283
rect 2531 2279 2535 2283
rect 2827 2279 2831 2283
rect 3011 2279 3015 2283
rect 3219 2279 3223 2283
rect 3451 2279 3455 2283
rect 3507 2279 3511 2283
rect 3915 2279 3919 2283
rect 111 2269 115 2273
rect 135 2272 139 2276
rect 271 2272 275 2276
rect 431 2272 435 2276
rect 591 2272 595 2276
rect 751 2272 755 2276
rect 919 2272 923 2276
rect 1087 2272 1091 2276
rect 1263 2272 1267 2276
rect 1447 2272 1451 2276
rect 1631 2272 1635 2276
rect 1815 2272 1819 2276
rect 2007 2269 2011 2273
rect 2047 2268 2051 2272
rect 2071 2269 2075 2273
rect 2175 2269 2179 2273
rect 2311 2269 2315 2273
rect 2447 2269 2451 2273
rect 2591 2269 2595 2273
rect 2751 2269 2755 2273
rect 2935 2269 2939 2273
rect 3143 2269 3147 2273
rect 3375 2269 3379 2273
rect 3615 2269 3619 2273
rect 3839 2269 3843 2273
rect 3943 2268 3947 2272
rect 211 2263 215 2267
rect 347 2263 351 2267
rect 379 2263 383 2267
rect 667 2263 671 2267
rect 735 2263 739 2267
rect 995 2263 999 2267
rect 1163 2263 1167 2267
rect 1339 2263 1343 2267
rect 1523 2263 1527 2267
rect 1707 2263 1711 2267
rect 1883 2263 1887 2267
rect 111 2252 115 2256
rect 135 2253 139 2257
rect 271 2253 275 2257
rect 431 2253 435 2257
rect 591 2253 595 2257
rect 751 2253 755 2257
rect 919 2253 923 2257
rect 1087 2253 1091 2257
rect 1263 2253 1267 2257
rect 1447 2253 1451 2257
rect 1631 2253 1635 2257
rect 1815 2253 1819 2257
rect 2007 2252 2011 2256
rect 2267 2259 2271 2263
rect 2147 2251 2151 2255
rect 2531 2259 2535 2263
rect 3019 2259 3023 2263
rect 379 2243 383 2247
rect 2483 2247 2484 2251
rect 2484 2247 2487 2251
rect 2523 2251 2527 2255
rect 2827 2247 2831 2251
rect 3011 2251 3015 2255
rect 3219 2251 3223 2255
rect 3451 2251 3455 2255
rect 3907 2251 3911 2255
rect 211 2235 215 2239
rect 403 2231 407 2235
rect 735 2235 739 2239
rect 967 2239 971 2243
rect 987 2231 991 2235
rect 995 2235 999 2239
rect 1163 2235 1167 2239
rect 1339 2235 1343 2239
rect 1671 2235 1672 2239
rect 1672 2235 1675 2239
rect 1707 2235 1711 2239
rect 3507 2235 3511 2239
rect 2187 2227 2191 2231
rect 2331 2227 2335 2231
rect 2643 2227 2647 2231
rect 2659 2227 2663 2231
rect 2955 2227 2959 2231
rect 3123 2227 3127 2231
rect 3299 2227 3303 2231
rect 3483 2227 3487 2231
rect 3867 2227 3871 2231
rect 235 2219 239 2223
rect 563 2219 567 2223
rect 667 2219 671 2223
rect 1163 2219 1167 2223
rect 1411 2219 1415 2223
rect 1523 2219 1527 2223
rect 1883 2219 1887 2223
rect 2491 2219 2495 2223
rect 411 2211 415 2215
rect 2047 2208 2051 2212
rect 2111 2207 2115 2211
rect 2255 2207 2259 2211
rect 2407 2207 2411 2211
rect 2559 2207 2563 2211
rect 2719 2207 2723 2211
rect 2879 2207 2883 2211
rect 3047 2207 3051 2211
rect 3223 2207 3227 2211
rect 3407 2207 3411 2211
rect 3591 2207 3595 2211
rect 3783 2207 3787 2211
rect 3943 2208 3947 2212
rect 111 2200 115 2204
rect 159 2199 163 2203
rect 327 2199 331 2203
rect 495 2199 499 2203
rect 679 2199 683 2203
rect 879 2199 883 2203
rect 1095 2199 1099 2203
rect 1327 2199 1331 2203
rect 1567 2199 1571 2203
rect 1815 2199 1819 2203
rect 2007 2200 2011 2204
rect 2187 2199 2191 2203
rect 2331 2199 2335 2203
rect 2483 2199 2487 2203
rect 2491 2199 2495 2203
rect 2643 2199 2647 2203
rect 2955 2199 2959 2203
rect 3123 2199 3127 2203
rect 3299 2199 3303 2203
rect 3483 2199 3487 2203
rect 3559 2199 3563 2203
rect 3747 2199 3751 2203
rect 235 2191 239 2195
rect 403 2191 407 2195
rect 411 2191 415 2195
rect 827 2191 831 2195
rect 987 2191 991 2195
rect 1303 2191 1307 2195
rect 1411 2191 1415 2195
rect 111 2183 115 2187
rect 1891 2187 1895 2191
rect 2047 2191 2051 2195
rect 2111 2188 2115 2192
rect 2255 2188 2259 2192
rect 2407 2188 2411 2192
rect 2559 2188 2563 2192
rect 2719 2188 2723 2192
rect 2879 2188 2883 2192
rect 3047 2188 3051 2192
rect 3223 2188 3227 2192
rect 3407 2188 3411 2192
rect 3591 2188 3595 2192
rect 3783 2188 3787 2192
rect 3943 2191 3947 2195
rect 159 2180 163 2184
rect 327 2180 331 2184
rect 495 2180 499 2184
rect 679 2180 683 2184
rect 879 2180 883 2184
rect 1095 2180 1099 2184
rect 1327 2180 1331 2184
rect 1567 2180 1571 2184
rect 1815 2180 1819 2184
rect 2007 2183 2011 2187
rect 3087 2139 3091 2143
rect 3559 2139 3563 2143
rect 111 2117 115 2121
rect 223 2120 227 2124
rect 359 2120 363 2124
rect 495 2120 499 2124
rect 639 2120 643 2124
rect 783 2120 787 2124
rect 935 2120 939 2124
rect 1095 2120 1099 2124
rect 1263 2120 1267 2124
rect 1447 2120 1451 2124
rect 1631 2120 1635 2124
rect 1823 2120 1827 2124
rect 2007 2117 2011 2121
rect 299 2111 303 2115
rect 435 2111 439 2115
rect 563 2111 567 2115
rect 579 2111 583 2115
rect 1011 2111 1015 2115
rect 1163 2111 1167 2115
rect 1339 2111 1343 2115
rect 1523 2111 1527 2115
rect 1623 2111 1627 2115
rect 1815 2111 1819 2115
rect 2047 2113 2051 2117
rect 2287 2116 2291 2120
rect 2431 2116 2435 2120
rect 2583 2116 2587 2120
rect 2735 2116 2739 2120
rect 2887 2116 2891 2120
rect 3047 2116 3051 2120
rect 3207 2116 3211 2120
rect 3367 2116 3371 2120
rect 3527 2116 3531 2120
rect 3695 2116 3699 2120
rect 3839 2116 3843 2120
rect 3943 2113 3947 2117
rect 2363 2107 2367 2111
rect 2507 2107 2511 2111
rect 2659 2107 2663 2111
rect 2667 2107 2671 2111
rect 2819 2107 2823 2111
rect 3123 2107 3127 2111
rect 3283 2107 3287 2111
rect 3443 2107 3447 2111
rect 3603 2107 3607 2111
rect 3619 2107 3623 2111
rect 3907 2107 3911 2111
rect 111 2100 115 2104
rect 223 2101 227 2105
rect 359 2101 363 2105
rect 495 2101 499 2105
rect 639 2101 643 2105
rect 783 2101 787 2105
rect 935 2101 939 2105
rect 1095 2101 1099 2105
rect 1263 2101 1267 2105
rect 1447 2101 1451 2105
rect 1631 2101 1635 2105
rect 1823 2101 1827 2105
rect 2007 2100 2011 2104
rect 2047 2096 2051 2100
rect 2287 2097 2291 2101
rect 2431 2097 2435 2101
rect 2583 2097 2587 2101
rect 2735 2097 2739 2101
rect 2887 2097 2891 2101
rect 3047 2097 3051 2101
rect 3207 2097 3211 2101
rect 3367 2097 3371 2101
rect 3527 2097 3531 2101
rect 3695 2097 3699 2101
rect 3839 2097 3843 2101
rect 3943 2096 3947 2100
rect 579 2091 583 2095
rect 299 2079 303 2083
rect 435 2083 439 2087
rect 691 2079 695 2083
rect 823 2083 824 2087
rect 824 2083 827 2087
rect 1003 2079 1007 2083
rect 1011 2083 1015 2087
rect 1303 2083 1304 2087
rect 1304 2083 1307 2087
rect 1339 2083 1343 2087
rect 1523 2083 1527 2087
rect 1891 2083 1895 2087
rect 2667 2087 2671 2091
rect 2363 2079 2367 2083
rect 2507 2079 2511 2083
rect 2819 2079 2823 2083
rect 2927 2075 2928 2079
rect 2928 2075 2931 2079
rect 3087 2079 3088 2083
rect 3088 2079 3091 2083
rect 3123 2079 3127 2083
rect 3283 2079 3287 2083
rect 3443 2079 3447 2083
rect 3603 2079 3607 2083
rect 3915 2079 3919 2083
rect 415 2059 416 2063
rect 416 2059 419 2063
rect 451 2059 455 2063
rect 571 2059 575 2063
rect 827 2059 831 2063
rect 1131 2059 1135 2063
rect 1227 2059 1231 2063
rect 1483 2059 1487 2063
rect 1623 2059 1624 2063
rect 1624 2059 1627 2063
rect 1815 2059 1816 2063
rect 1816 2059 1819 2063
rect 3619 2063 3623 2067
rect 2563 2055 2567 2059
rect 2747 2055 2751 2059
rect 2915 2055 2919 2059
rect 3243 2055 3247 2059
rect 3387 2055 3391 2059
rect 3667 2055 3671 2059
rect 3907 2055 3911 2059
rect 111 2040 115 2044
rect 375 2039 379 2043
rect 495 2039 499 2043
rect 615 2039 619 2043
rect 751 2039 755 2043
rect 895 2039 899 2043
rect 1047 2039 1051 2043
rect 1215 2039 1219 2043
rect 1399 2039 1403 2043
rect 1583 2039 1587 2043
rect 1775 2039 1779 2043
rect 2007 2040 2011 2044
rect 2047 2036 2051 2040
rect 451 2031 455 2035
rect 571 2031 575 2035
rect 691 2031 695 2035
rect 827 2031 831 2035
rect 887 2031 891 2035
rect 1003 2031 1007 2035
rect 1131 2031 1135 2035
rect 111 2023 115 2027
rect 1475 2027 1479 2031
rect 1483 2031 1487 2035
rect 2503 2035 2507 2039
rect 1755 2031 1759 2035
rect 2671 2035 2675 2039
rect 2839 2035 2843 2039
rect 3007 2035 3011 2039
rect 3167 2035 3171 2039
rect 3311 2035 3315 2039
rect 3455 2035 3459 2039
rect 3591 2035 3595 2039
rect 3727 2035 3731 2039
rect 3839 2035 3843 2039
rect 3943 2036 3947 2040
rect 375 2020 379 2024
rect 495 2020 499 2024
rect 615 2020 619 2024
rect 751 2020 755 2024
rect 895 2020 899 2024
rect 1047 2020 1051 2024
rect 1215 2020 1219 2024
rect 1399 2020 1403 2024
rect 1583 2020 1587 2024
rect 1775 2020 1779 2024
rect 2007 2023 2011 2027
rect 2747 2027 2751 2031
rect 2915 2027 2919 2031
rect 2927 2027 2931 2031
rect 3243 2027 3247 2031
rect 3387 2027 3391 2031
rect 3667 2027 3671 2031
rect 3711 2027 3715 2031
rect 2047 2019 2051 2023
rect 3915 2023 3919 2027
rect 2503 2016 2507 2020
rect 2671 2016 2675 2020
rect 2839 2016 2843 2020
rect 3007 2016 3011 2020
rect 3167 2016 3171 2020
rect 3311 2016 3315 2020
rect 3455 2016 3459 2020
rect 3591 2016 3595 2020
rect 3727 2016 3731 2020
rect 3839 2016 3843 2020
rect 3943 2019 3947 2023
rect 111 1949 115 1953
rect 511 1952 515 1956
rect 623 1952 627 1956
rect 743 1952 747 1956
rect 871 1952 875 1956
rect 1007 1952 1011 1956
rect 1143 1952 1147 1956
rect 1279 1952 1283 1956
rect 1415 1952 1419 1956
rect 1559 1952 1563 1956
rect 1703 1952 1707 1956
rect 2007 1949 2011 1953
rect 2047 1949 2051 1953
rect 2495 1952 2499 1956
rect 2591 1952 2595 1956
rect 2695 1952 2699 1956
rect 2807 1952 2811 1956
rect 2927 1952 2931 1956
rect 3047 1952 3051 1956
rect 3175 1952 3179 1956
rect 3295 1952 3299 1956
rect 3415 1952 3419 1956
rect 3543 1952 3547 1956
rect 3671 1952 3675 1956
rect 3799 1952 3803 1956
rect 3943 1949 3947 1953
rect 415 1943 419 1947
rect 595 1943 599 1947
rect 719 1943 723 1947
rect 947 1943 951 1947
rect 1083 1943 1087 1947
rect 1227 1943 1231 1947
rect 1347 1943 1351 1947
rect 1491 1943 1495 1947
rect 1519 1943 1523 1947
rect 1771 1943 1775 1947
rect 2563 1943 2567 1947
rect 2579 1943 2583 1947
rect 2683 1943 2687 1947
rect 2779 1943 2783 1947
rect 3003 1943 3007 1947
rect 3123 1943 3127 1947
rect 3131 1943 3135 1947
rect 3259 1943 3263 1947
rect 3387 1943 3391 1947
rect 3631 1943 3635 1947
rect 3867 1943 3871 1947
rect 111 1932 115 1936
rect 511 1933 515 1937
rect 623 1933 627 1937
rect 743 1933 747 1937
rect 871 1933 875 1937
rect 1007 1933 1011 1937
rect 1143 1933 1147 1937
rect 1279 1933 1283 1937
rect 1415 1933 1419 1937
rect 1559 1933 1563 1937
rect 1703 1933 1707 1937
rect 2007 1932 2011 1936
rect 2047 1932 2051 1936
rect 2495 1933 2499 1937
rect 2591 1933 2595 1937
rect 2695 1933 2699 1937
rect 2807 1933 2811 1937
rect 2927 1933 2931 1937
rect 3047 1933 3051 1937
rect 3175 1933 3179 1937
rect 3295 1933 3299 1937
rect 3415 1933 3419 1937
rect 3543 1933 3547 1937
rect 3671 1933 3675 1937
rect 3799 1933 3803 1937
rect 3943 1932 3947 1936
rect 595 1915 599 1919
rect 719 1915 723 1919
rect 887 1915 891 1919
rect 947 1915 951 1919
rect 1519 1923 1523 1927
rect 1475 1915 1479 1919
rect 1491 1915 1495 1919
rect 1755 1915 1759 1919
rect 2579 1915 2583 1919
rect 2683 1915 2687 1919
rect 2779 1915 2783 1919
rect 3131 1923 3135 1927
rect 2867 1911 2871 1915
rect 3003 1915 3007 1919
rect 3123 1915 3127 1919
rect 3387 1915 3391 1919
rect 3631 1915 3635 1919
rect 3711 1915 3712 1919
rect 3712 1915 3715 1919
rect 3859 1911 3863 1915
rect 3259 1903 3263 1907
rect 579 1891 583 1895
rect 647 1891 651 1895
rect 859 1891 863 1895
rect 1083 1891 1084 1895
rect 1084 1891 1087 1895
rect 1215 1891 1216 1895
rect 1216 1891 1219 1895
rect 1347 1891 1348 1895
rect 1348 1891 1351 1895
rect 1387 1891 1391 1895
rect 1523 1891 1527 1895
rect 1771 1891 1775 1895
rect 1923 1895 1927 1899
rect 2323 1895 2327 1899
rect 2515 1895 2519 1899
rect 3035 1895 3039 1899
rect 3203 1895 3207 1899
rect 3379 1895 3383 1899
rect 3563 1895 3567 1899
rect 3915 1895 3919 1899
rect 2479 1887 2483 1891
rect 111 1872 115 1876
rect 551 1871 555 1875
rect 663 1871 667 1875
rect 783 1871 787 1875
rect 911 1871 915 1875
rect 1047 1871 1051 1875
rect 1175 1871 1179 1875
rect 1311 1871 1315 1875
rect 1447 1871 1451 1875
rect 1583 1871 1587 1875
rect 1719 1871 1723 1875
rect 2007 1872 2011 1876
rect 2047 1876 2051 1880
rect 2071 1875 2075 1879
rect 2247 1875 2251 1879
rect 2439 1875 2443 1879
rect 2623 1875 2627 1879
rect 2791 1875 2795 1879
rect 2959 1875 2963 1879
rect 3127 1875 3131 1879
rect 3303 1875 3307 1879
rect 3487 1875 3491 1879
rect 3671 1875 3675 1879
rect 3839 1875 3843 1879
rect 3943 1876 3947 1880
rect 647 1863 651 1867
rect 859 1863 863 1867
rect 1039 1863 1043 1867
rect 1387 1863 1391 1867
rect 1523 1863 1527 1867
rect 1703 1863 1707 1867
rect 111 1855 115 1859
rect 551 1852 555 1856
rect 663 1852 667 1856
rect 783 1852 787 1856
rect 911 1852 915 1856
rect 1047 1852 1051 1856
rect 1175 1852 1179 1856
rect 1311 1852 1315 1856
rect 1447 1852 1451 1856
rect 1583 1852 1587 1856
rect 1711 1855 1715 1859
rect 1719 1852 1723 1856
rect 2007 1855 2011 1859
rect 2047 1859 2051 1863
rect 2147 1863 2151 1867
rect 2323 1867 2327 1871
rect 2515 1867 2519 1871
rect 2867 1867 2871 1871
rect 3035 1867 3039 1871
rect 3203 1867 3207 1871
rect 3379 1867 3383 1871
rect 3563 1867 3567 1871
rect 3607 1867 3611 1871
rect 3915 1863 3919 1867
rect 2071 1856 2075 1860
rect 2247 1856 2251 1860
rect 2439 1856 2443 1860
rect 2623 1856 2627 1860
rect 2791 1856 2795 1860
rect 2959 1856 2963 1860
rect 3127 1856 3131 1860
rect 3303 1856 3307 1860
rect 3487 1856 3491 1860
rect 3671 1856 3675 1860
rect 3839 1856 3843 1860
rect 3943 1859 3947 1863
rect 111 1789 115 1793
rect 503 1792 507 1796
rect 615 1792 619 1796
rect 735 1792 739 1796
rect 863 1792 867 1796
rect 999 1792 1003 1796
rect 1151 1792 1155 1796
rect 1319 1792 1323 1796
rect 1487 1792 1491 1796
rect 1663 1792 1667 1796
rect 1847 1792 1851 1796
rect 2007 1789 2011 1793
rect 2047 1793 2051 1797
rect 2095 1796 2099 1800
rect 2231 1796 2235 1800
rect 2367 1796 2371 1800
rect 2511 1796 2515 1800
rect 2671 1796 2675 1800
rect 2855 1796 2859 1800
rect 3071 1796 3075 1800
rect 3303 1796 3307 1800
rect 3543 1796 3547 1800
rect 3791 1796 3795 1800
rect 3943 1793 3947 1797
rect 579 1783 583 1787
rect 591 1783 595 1787
rect 711 1783 715 1787
rect 931 1783 935 1787
rect 971 1783 975 1787
rect 1219 1783 1223 1787
rect 1263 1783 1267 1787
rect 1563 1783 1567 1787
rect 1923 1783 1927 1787
rect 2171 1787 2175 1791
rect 2307 1787 2311 1791
rect 2435 1787 2439 1791
rect 2479 1787 2483 1791
rect 2771 1787 2775 1791
rect 2939 1787 2943 1791
rect 3167 1787 3171 1791
rect 3423 1787 3427 1791
rect 3859 1787 3863 1791
rect 111 1772 115 1776
rect 503 1773 507 1777
rect 615 1773 619 1777
rect 735 1773 739 1777
rect 863 1773 867 1777
rect 999 1773 1003 1777
rect 1151 1773 1155 1777
rect 1319 1773 1323 1777
rect 1487 1773 1491 1777
rect 1663 1773 1667 1777
rect 1847 1773 1851 1777
rect 2007 1772 2011 1776
rect 2047 1776 2051 1780
rect 2095 1777 2099 1781
rect 2231 1777 2235 1781
rect 2367 1777 2371 1781
rect 2511 1777 2515 1781
rect 2671 1777 2675 1781
rect 2855 1777 2859 1781
rect 3071 1777 3075 1781
rect 3303 1777 3307 1781
rect 3543 1777 3547 1781
rect 3791 1777 3795 1781
rect 3943 1776 3947 1780
rect 591 1755 595 1759
rect 711 1755 715 1759
rect 795 1751 799 1755
rect 971 1755 975 1759
rect 1039 1755 1040 1759
rect 1040 1755 1043 1759
rect 1263 1755 1267 1759
rect 931 1747 935 1751
rect 1359 1751 1360 1755
rect 1360 1751 1363 1755
rect 1703 1755 1704 1759
rect 1704 1755 1707 1759
rect 1711 1755 1715 1759
rect 2147 1759 2151 1763
rect 2171 1759 2175 1763
rect 2307 1759 2311 1763
rect 2683 1755 2687 1759
rect 2939 1759 2943 1763
rect 3167 1759 3171 1763
rect 3423 1759 3427 1763
rect 3607 1759 3611 1763
rect 3799 1755 3803 1759
rect 419 1739 423 1743
rect 539 1739 543 1743
rect 667 1739 671 1743
rect 923 1739 927 1743
rect 1159 1739 1163 1743
rect 1203 1739 1207 1743
rect 1355 1739 1359 1743
rect 1563 1739 1567 1743
rect 2267 1743 2271 1747
rect 2375 1743 2379 1747
rect 2427 1749 2431 1751
rect 2427 1747 2428 1749
rect 2428 1747 2431 1749
rect 2571 1743 2575 1747
rect 2771 1743 2775 1747
rect 2779 1743 2783 1747
rect 2883 1743 2887 1747
rect 2987 1743 2991 1747
rect 3091 1743 3095 1747
rect 739 1731 743 1735
rect 2627 1735 2631 1739
rect 111 1720 115 1724
rect 343 1719 347 1723
rect 463 1719 467 1723
rect 591 1719 595 1723
rect 719 1719 723 1723
rect 847 1719 851 1723
rect 983 1719 987 1723
rect 1127 1719 1131 1723
rect 1279 1719 1283 1723
rect 1439 1719 1443 1723
rect 1599 1719 1603 1723
rect 2007 1720 2011 1724
rect 2047 1724 2051 1728
rect 2183 1723 2187 1727
rect 2287 1723 2291 1727
rect 2391 1723 2395 1727
rect 2495 1723 2499 1727
rect 2599 1723 2603 1727
rect 2703 1723 2707 1727
rect 2807 1723 2811 1727
rect 2911 1723 2915 1727
rect 3015 1723 3019 1727
rect 3127 1723 3131 1727
rect 3943 1724 3947 1728
rect 419 1711 423 1715
rect 539 1711 543 1715
rect 667 1711 671 1715
rect 795 1711 799 1715
rect 923 1711 927 1715
rect 111 1703 115 1707
rect 1059 1707 1063 1711
rect 1203 1711 1207 1715
rect 1355 1711 1359 1715
rect 1363 1711 1367 1715
rect 1583 1711 1587 1715
rect 343 1700 347 1704
rect 463 1700 467 1704
rect 591 1700 595 1704
rect 719 1700 723 1704
rect 847 1700 851 1704
rect 983 1700 987 1704
rect 1127 1700 1131 1704
rect 1279 1700 1283 1704
rect 1439 1700 1443 1704
rect 1599 1700 1603 1704
rect 2007 1703 2011 1707
rect 2047 1707 2051 1711
rect 2259 1711 2263 1715
rect 2267 1715 2271 1719
rect 2375 1715 2379 1719
rect 2571 1715 2575 1719
rect 2683 1715 2687 1719
rect 2779 1715 2783 1719
rect 2883 1715 2887 1719
rect 2987 1715 2991 1719
rect 3091 1715 3095 1719
rect 3203 1711 3207 1715
rect 2183 1704 2187 1708
rect 2287 1704 2291 1708
rect 2391 1704 2395 1708
rect 2495 1704 2499 1708
rect 2599 1704 2603 1708
rect 2703 1704 2707 1708
rect 2807 1704 2811 1708
rect 2911 1704 2915 1708
rect 3015 1704 3019 1708
rect 3127 1704 3131 1708
rect 3943 1707 3947 1711
rect 2047 1641 2051 1645
rect 2231 1644 2235 1648
rect 2367 1644 2371 1648
rect 2519 1644 2523 1648
rect 2679 1644 2683 1648
rect 2847 1644 2851 1648
rect 3023 1644 3027 1648
rect 3191 1644 3195 1648
rect 3359 1644 3363 1648
rect 3527 1644 3531 1648
rect 3695 1644 3699 1648
rect 3839 1644 3843 1648
rect 111 1633 115 1637
rect 159 1636 163 1640
rect 295 1636 299 1640
rect 455 1636 459 1640
rect 623 1636 627 1640
rect 799 1636 803 1640
rect 983 1636 987 1640
rect 1167 1636 1171 1640
rect 1351 1636 1355 1640
rect 1543 1636 1547 1640
rect 3943 1641 3947 1645
rect 1735 1636 1739 1640
rect 2007 1633 2011 1637
rect 2307 1635 2311 1639
rect 2443 1635 2447 1639
rect 2595 1635 2599 1639
rect 2627 1635 2631 1639
rect 2763 1635 2767 1639
rect 3107 1635 3111 1639
rect 3435 1635 3439 1639
rect 3603 1635 3607 1639
rect 3907 1635 3911 1639
rect 235 1627 239 1631
rect 371 1627 375 1631
rect 531 1627 535 1631
rect 699 1627 703 1631
rect 739 1627 743 1631
rect 1051 1627 1055 1631
rect 1159 1627 1163 1631
rect 1619 1627 1623 1631
rect 1803 1627 1807 1631
rect 2047 1624 2051 1628
rect 2231 1625 2235 1629
rect 2367 1625 2371 1629
rect 2519 1625 2523 1629
rect 2679 1625 2683 1629
rect 2847 1625 2851 1629
rect 3023 1625 3027 1629
rect 3191 1625 3195 1629
rect 3359 1625 3363 1629
rect 3527 1625 3531 1629
rect 3695 1625 3699 1629
rect 3839 1625 3843 1629
rect 3943 1624 3947 1628
rect 111 1616 115 1620
rect 159 1617 163 1621
rect 295 1617 299 1621
rect 455 1617 459 1621
rect 623 1617 627 1621
rect 799 1617 803 1621
rect 983 1617 987 1621
rect 1167 1617 1171 1621
rect 1351 1617 1355 1621
rect 1543 1617 1547 1621
rect 1735 1617 1739 1621
rect 2007 1616 2011 1620
rect 235 1603 239 1607
rect 2259 1607 2263 1611
rect 2307 1607 2311 1611
rect 2443 1607 2447 1611
rect 2763 1607 2767 1611
rect 371 1599 375 1603
rect 531 1599 535 1603
rect 699 1599 703 1603
rect 1059 1599 1063 1603
rect 739 1591 743 1595
rect 1443 1595 1447 1599
rect 1583 1599 1584 1603
rect 1584 1599 1587 1603
rect 1619 1599 1623 1603
rect 2787 1603 2791 1607
rect 3203 1607 3207 1611
rect 3399 1603 3400 1607
rect 3400 1603 3403 1607
rect 3435 1607 3439 1611
rect 3603 1607 3607 1611
rect 3915 1607 3919 1611
rect 203 1583 207 1587
rect 211 1583 215 1587
rect 331 1583 335 1587
rect 499 1583 503 1587
rect 683 1583 687 1587
rect 1051 1583 1055 1587
rect 1251 1583 1255 1587
rect 1259 1583 1263 1587
rect 1635 1583 1639 1587
rect 1803 1583 1807 1587
rect 1979 1583 1983 1587
rect 2147 1583 2151 1587
rect 2347 1583 2351 1587
rect 2595 1583 2599 1587
rect 2995 1583 2999 1587
rect 3107 1583 3111 1587
rect 3203 1583 3207 1587
rect 3339 1583 3343 1587
rect 3807 1583 3811 1587
rect 3907 1583 3911 1587
rect 1763 1575 1767 1579
rect 111 1564 115 1568
rect 135 1563 139 1567
rect 255 1563 259 1567
rect 423 1563 427 1567
rect 607 1563 611 1567
rect 799 1563 803 1567
rect 991 1563 995 1567
rect 1183 1563 1187 1567
rect 1367 1563 1371 1567
rect 1551 1563 1555 1567
rect 1735 1563 1739 1567
rect 1903 1563 1907 1567
rect 2007 1564 2011 1568
rect 2047 1564 2051 1568
rect 2071 1563 2075 1567
rect 2271 1563 2275 1567
rect 2495 1563 2499 1567
rect 2711 1563 2715 1567
rect 2911 1563 2915 1567
rect 3095 1563 3099 1567
rect 3263 1563 3267 1567
rect 3423 1563 3427 1567
rect 3567 1563 3571 1567
rect 3711 1563 3715 1567
rect 3839 1563 3843 1567
rect 3943 1564 3947 1568
rect 211 1555 215 1559
rect 331 1555 335 1559
rect 499 1555 503 1559
rect 683 1555 687 1559
rect 739 1555 743 1559
rect 111 1547 115 1551
rect 1067 1551 1071 1555
rect 1259 1555 1263 1559
rect 1443 1555 1447 1559
rect 1455 1555 1459 1559
rect 1635 1555 1639 1559
rect 1979 1555 1983 1559
rect 2147 1555 2151 1559
rect 2347 1555 2351 1559
rect 2419 1555 2423 1559
rect 2787 1555 2791 1559
rect 2995 1555 2999 1559
rect 3339 1555 3343 1559
rect 3399 1555 3403 1559
rect 3507 1555 3511 1559
rect 3799 1555 3803 1559
rect 3807 1555 3811 1559
rect 135 1544 139 1548
rect 255 1544 259 1548
rect 423 1544 427 1548
rect 607 1544 611 1548
rect 799 1544 803 1548
rect 991 1544 995 1548
rect 1183 1544 1187 1548
rect 1367 1544 1371 1548
rect 1551 1544 1555 1548
rect 1735 1544 1739 1548
rect 1903 1544 1907 1548
rect 2007 1547 2011 1551
rect 2047 1547 2051 1551
rect 2071 1544 2075 1548
rect 2271 1544 2275 1548
rect 2495 1544 2499 1548
rect 2711 1544 2715 1548
rect 2911 1544 2915 1548
rect 3095 1544 3099 1548
rect 3263 1544 3267 1548
rect 3423 1544 3427 1548
rect 3567 1544 3571 1548
rect 3711 1544 3715 1548
rect 3839 1544 3843 1548
rect 3943 1547 3947 1551
rect 203 1487 207 1491
rect 111 1477 115 1481
rect 135 1480 139 1484
rect 247 1480 251 1484
rect 399 1480 403 1484
rect 559 1480 563 1484
rect 211 1471 215 1475
rect 323 1471 327 1475
rect 475 1471 479 1475
rect 635 1471 639 1475
rect 719 1480 723 1484
rect 879 1480 883 1484
rect 1039 1480 1043 1484
rect 1183 1480 1187 1484
rect 1319 1480 1323 1484
rect 1447 1480 1451 1484
rect 1567 1480 1571 1484
rect 1687 1480 1691 1484
rect 1807 1480 1811 1484
rect 1903 1480 1907 1484
rect 2007 1477 2011 1481
rect 2047 1481 2051 1485
rect 2071 1484 2075 1488
rect 2431 1484 2435 1488
rect 2791 1484 2795 1488
rect 3127 1484 3131 1488
rect 3463 1484 3467 1488
rect 3799 1484 3803 1488
rect 3943 1481 3947 1485
rect 955 1471 959 1475
rect 1251 1471 1255 1475
rect 1395 1471 1399 1475
rect 1523 1471 1527 1475
rect 1643 1471 1647 1475
rect 1763 1471 1767 1475
rect 1883 1471 1887 1475
rect 1895 1471 1899 1475
rect 2055 1475 2059 1479
rect 2719 1475 2723 1479
rect 2867 1475 2871 1479
rect 3203 1475 3207 1479
rect 3539 1475 3543 1479
rect 3867 1475 3871 1479
rect 111 1460 115 1464
rect 135 1461 139 1465
rect 247 1461 251 1465
rect 399 1461 403 1465
rect 559 1461 563 1465
rect 719 1461 723 1465
rect 879 1461 883 1465
rect 1039 1461 1043 1465
rect 1183 1461 1187 1465
rect 1319 1461 1323 1465
rect 1447 1461 1451 1465
rect 1567 1461 1571 1465
rect 1687 1461 1691 1465
rect 1807 1461 1811 1465
rect 1903 1461 1907 1465
rect 2007 1460 2011 1464
rect 2047 1464 2051 1468
rect 2071 1465 2075 1469
rect 2431 1465 2435 1469
rect 2791 1465 2795 1469
rect 3127 1465 3131 1469
rect 3463 1465 3467 1469
rect 3799 1465 3803 1469
rect 3943 1464 3947 1468
rect 211 1443 215 1447
rect 323 1443 327 1447
rect 475 1443 479 1447
rect 635 1443 639 1447
rect 1067 1443 1071 1447
rect 211 1435 215 1439
rect 1243 1439 1247 1443
rect 1455 1451 1459 1455
rect 1395 1443 1399 1447
rect 1523 1443 1527 1447
rect 1643 1443 1647 1447
rect 1895 1443 1899 1447
rect 2055 1443 2059 1447
rect 2419 1447 2423 1451
rect 2719 1447 2723 1451
rect 3167 1443 3168 1447
rect 3168 1443 3171 1447
rect 3503 1447 3504 1451
rect 3504 1447 3507 1451
rect 3539 1447 3543 1451
rect 219 1427 223 1431
rect 367 1427 371 1431
rect 579 1427 583 1431
rect 683 1427 687 1431
rect 955 1427 959 1431
rect 1051 1427 1055 1431
rect 1435 1427 1439 1431
rect 1627 1427 1631 1431
rect 1743 1427 1747 1431
rect 1883 1427 1887 1431
rect 691 1419 695 1423
rect 1979 1423 1983 1427
rect 2147 1423 2151 1427
rect 2347 1423 2351 1427
rect 2571 1423 2575 1427
rect 2867 1423 2871 1427
rect 2987 1423 2991 1427
rect 3355 1423 3359 1427
rect 3507 1423 3511 1427
rect 3523 1423 3527 1427
rect 3867 1423 3871 1427
rect 111 1408 115 1412
rect 135 1407 139 1411
rect 263 1407 267 1411
rect 431 1407 435 1411
rect 607 1407 611 1411
rect 791 1407 795 1411
rect 975 1407 979 1411
rect 1159 1407 1163 1411
rect 1351 1407 1355 1411
rect 1543 1407 1547 1411
rect 1735 1407 1739 1411
rect 1903 1407 1907 1411
rect 2007 1408 2011 1412
rect 2047 1404 2051 1408
rect 211 1399 215 1403
rect 219 1399 223 1403
rect 367 1399 371 1403
rect 683 1399 687 1403
rect 691 1399 695 1403
rect 1051 1399 1055 1403
rect 1083 1399 1087 1403
rect 1243 1399 1247 1403
rect 1435 1399 1439 1403
rect 1627 1399 1631 1403
rect 2071 1403 2075 1407
rect 1979 1399 1983 1403
rect 2271 1403 2275 1407
rect 2495 1403 2499 1407
rect 2711 1403 2715 1407
rect 2911 1403 2915 1407
rect 3095 1403 3099 1407
rect 3271 1403 3275 1407
rect 3439 1403 3443 1407
rect 111 1391 115 1395
rect 135 1388 139 1392
rect 263 1388 267 1392
rect 431 1388 435 1392
rect 607 1388 611 1392
rect 791 1388 795 1392
rect 975 1388 979 1392
rect 1159 1388 1163 1392
rect 1351 1388 1355 1392
rect 1543 1388 1547 1392
rect 1735 1388 1739 1392
rect 1903 1388 1907 1392
rect 2007 1391 2011 1395
rect 2147 1395 2151 1399
rect 2347 1395 2351 1399
rect 2571 1395 2575 1399
rect 2659 1395 2663 1399
rect 2987 1395 2991 1399
rect 3171 1395 3175 1399
rect 3199 1395 3203 1399
rect 3355 1395 3359 1399
rect 3507 1399 3511 1403
rect 3607 1403 3611 1407
rect 3783 1403 3787 1407
rect 3943 1404 3947 1408
rect 2047 1387 2051 1391
rect 3859 1391 3863 1395
rect 2071 1384 2075 1388
rect 2271 1384 2275 1388
rect 2495 1384 2499 1388
rect 2711 1384 2715 1388
rect 2911 1384 2915 1388
rect 3095 1384 3099 1388
rect 3271 1384 3275 1388
rect 3439 1384 3443 1388
rect 3607 1384 3611 1388
rect 3783 1384 3787 1388
rect 3943 1387 3947 1391
rect 111 1321 115 1325
rect 159 1324 163 1328
rect 311 1324 315 1328
rect 479 1324 483 1328
rect 663 1324 667 1328
rect 855 1324 859 1328
rect 1047 1324 1051 1328
rect 1247 1324 1251 1328
rect 1447 1324 1451 1328
rect 1655 1324 1659 1328
rect 1863 1324 1867 1328
rect 2007 1321 2011 1325
rect 2047 1321 2051 1325
rect 2071 1324 2075 1328
rect 2207 1324 2211 1328
rect 2383 1324 2387 1328
rect 2567 1324 2571 1328
rect 2751 1324 2755 1328
rect 2935 1324 2939 1328
rect 3111 1324 3115 1328
rect 3279 1324 3283 1328
rect 3447 1324 3451 1328
rect 3623 1324 3627 1328
rect 3943 1321 3947 1325
rect 263 1315 267 1319
rect 387 1315 391 1319
rect 579 1315 583 1319
rect 739 1315 743 1319
rect 747 1315 751 1319
rect 1123 1315 1127 1319
rect 1323 1315 1327 1319
rect 1523 1315 1527 1319
rect 1743 1315 1747 1319
rect 2147 1315 2151 1319
rect 2283 1315 2287 1319
rect 2459 1315 2463 1319
rect 2643 1315 2647 1319
rect 2719 1315 2723 1319
rect 3011 1315 3015 1319
rect 3187 1315 3191 1319
rect 3355 1315 3359 1319
rect 3523 1315 3527 1319
rect 111 1304 115 1308
rect 159 1305 163 1309
rect 311 1305 315 1309
rect 479 1305 483 1309
rect 663 1305 667 1309
rect 855 1305 859 1309
rect 1047 1305 1051 1309
rect 1247 1305 1251 1309
rect 1447 1305 1451 1309
rect 1655 1305 1659 1309
rect 1863 1305 1867 1309
rect 2007 1304 2011 1308
rect 2047 1304 2051 1308
rect 2071 1305 2075 1309
rect 2207 1305 2211 1309
rect 2383 1305 2387 1309
rect 2567 1305 2571 1309
rect 2751 1305 2755 1309
rect 2935 1305 2939 1309
rect 3111 1305 3115 1309
rect 3279 1305 3283 1309
rect 3447 1305 3451 1309
rect 3623 1305 3627 1309
rect 3943 1304 3947 1308
rect 747 1295 751 1299
rect 263 1283 267 1287
rect 387 1287 391 1291
rect 619 1283 623 1287
rect 739 1287 743 1291
rect 1083 1287 1084 1291
rect 1084 1287 1087 1291
rect 1123 1287 1127 1291
rect 1323 1287 1327 1291
rect 2659 1295 2663 1299
rect 2147 1287 2151 1291
rect 2283 1287 2287 1291
rect 2459 1287 2463 1291
rect 2643 1287 2647 1291
rect 3199 1295 3203 1299
rect 3011 1287 3015 1291
rect 3187 1287 3191 1291
rect 2719 1279 2723 1283
rect 2983 1279 2987 1283
rect 3691 1283 3695 1287
rect 447 1267 448 1271
rect 448 1267 451 1271
rect 675 1267 679 1271
rect 771 1267 775 1271
rect 931 1267 935 1271
rect 1275 1267 1279 1271
rect 1455 1267 1459 1271
rect 1523 1267 1527 1271
rect 1771 1267 1775 1271
rect 1795 1267 1799 1271
rect 2227 1271 2231 1275
rect 2363 1271 2367 1275
rect 2507 1271 2511 1275
rect 2659 1271 2663 1275
rect 2971 1271 2975 1275
rect 2979 1271 2983 1275
rect 3331 1271 3335 1275
rect 3355 1271 3359 1275
rect 3699 1271 3703 1275
rect 3859 1271 3863 1275
rect 111 1248 115 1252
rect 407 1247 411 1251
rect 543 1247 547 1251
rect 695 1247 699 1251
rect 855 1247 859 1251
rect 1023 1247 1027 1251
rect 1191 1247 1195 1251
rect 1367 1247 1371 1251
rect 1543 1247 1547 1251
rect 1719 1247 1723 1251
rect 1895 1247 1899 1251
rect 2007 1248 2011 1252
rect 2047 1252 2051 1256
rect 2151 1251 2155 1255
rect 2287 1251 2291 1255
rect 2431 1251 2435 1255
rect 2583 1251 2587 1255
rect 2743 1251 2747 1255
rect 2903 1251 2907 1255
rect 3071 1251 3075 1255
rect 3247 1251 3251 1255
rect 3431 1251 3435 1255
rect 3615 1251 3619 1255
rect 3807 1251 3811 1255
rect 3943 1252 3947 1256
rect 619 1239 623 1243
rect 771 1239 775 1243
rect 931 1239 935 1243
rect 979 1239 983 1243
rect 111 1231 115 1235
rect 1267 1235 1271 1239
rect 1275 1239 1279 1243
rect 1455 1239 1459 1243
rect 1795 1239 1799 1243
rect 2227 1243 2231 1247
rect 2363 1243 2367 1247
rect 2507 1243 2511 1247
rect 2659 1243 2663 1247
rect 2667 1243 2671 1247
rect 2979 1243 2983 1247
rect 407 1228 411 1232
rect 543 1228 547 1232
rect 695 1228 699 1232
rect 855 1228 859 1232
rect 1023 1228 1027 1232
rect 1191 1228 1195 1232
rect 1367 1228 1371 1232
rect 1543 1228 1547 1232
rect 1719 1228 1723 1232
rect 1895 1228 1899 1232
rect 2007 1231 2011 1235
rect 2047 1235 2051 1239
rect 3331 1243 3335 1247
rect 3691 1243 3695 1247
rect 3883 1239 3887 1243
rect 2151 1232 2155 1236
rect 2287 1232 2291 1236
rect 2431 1232 2435 1236
rect 2583 1232 2587 1236
rect 2743 1232 2747 1236
rect 2903 1232 2907 1236
rect 3071 1232 3075 1236
rect 3247 1232 3251 1236
rect 3431 1232 3435 1236
rect 3615 1232 3619 1236
rect 3807 1232 3811 1236
rect 3943 1235 3947 1239
rect 2351 1211 2355 1215
rect 2667 1211 2671 1215
rect 111 1165 115 1169
rect 423 1168 427 1172
rect 591 1168 595 1172
rect 759 1168 763 1172
rect 927 1168 931 1172
rect 1095 1168 1099 1172
rect 1247 1168 1251 1172
rect 1399 1168 1403 1172
rect 1543 1168 1547 1172
rect 1687 1168 1691 1172
rect 1839 1168 1843 1172
rect 2007 1165 2011 1169
rect 2047 1169 2051 1173
rect 2311 1172 2315 1176
rect 2415 1172 2419 1176
rect 2527 1172 2531 1176
rect 2639 1172 2643 1176
rect 2767 1172 2771 1176
rect 2911 1172 2915 1176
rect 3071 1172 3075 1176
rect 3247 1172 3251 1176
rect 3439 1172 3443 1176
rect 3631 1172 3635 1176
rect 3831 1172 3835 1176
rect 3943 1169 3947 1173
rect 499 1159 503 1163
rect 675 1159 679 1163
rect 719 1159 723 1163
rect 879 1159 883 1163
rect 1323 1159 1327 1163
rect 1619 1159 1623 1163
rect 1763 1159 1767 1163
rect 1771 1159 1775 1163
rect 2387 1163 2391 1167
rect 2491 1163 2495 1167
rect 2603 1163 2607 1167
rect 2715 1163 2719 1167
rect 2723 1163 2727 1167
rect 2987 1163 2991 1167
rect 3139 1163 3143 1167
rect 3323 1163 3327 1167
rect 3379 1163 3383 1167
rect 3699 1163 3703 1167
rect 3899 1163 3903 1167
rect 111 1148 115 1152
rect 423 1149 427 1153
rect 591 1149 595 1153
rect 759 1149 763 1153
rect 927 1149 931 1153
rect 1095 1149 1099 1153
rect 1247 1149 1251 1153
rect 1399 1149 1403 1153
rect 1543 1149 1547 1153
rect 1687 1149 1691 1153
rect 1839 1149 1843 1153
rect 2007 1148 2011 1152
rect 2047 1152 2051 1156
rect 2311 1153 2315 1157
rect 2415 1153 2419 1157
rect 2527 1153 2531 1157
rect 2639 1153 2643 1157
rect 2767 1153 2771 1157
rect 2911 1153 2915 1157
rect 3071 1153 3075 1157
rect 3247 1153 3251 1157
rect 3439 1153 3443 1157
rect 3631 1153 3635 1157
rect 3831 1153 3835 1157
rect 3943 1152 3947 1156
rect 451 1127 455 1131
rect 499 1131 503 1135
rect 879 1131 883 1135
rect 1195 1127 1199 1131
rect 1267 1131 1271 1135
rect 1323 1131 1327 1135
rect 1583 1127 1584 1131
rect 1584 1127 1587 1131
rect 1619 1131 1623 1135
rect 1763 1131 1767 1135
rect 2351 1135 2352 1139
rect 2352 1135 2355 1139
rect 2387 1135 2391 1139
rect 2491 1135 2495 1139
rect 2603 1135 2607 1139
rect 2715 1135 2719 1139
rect 3379 1143 3383 1147
rect 2987 1135 2991 1139
rect 3323 1135 3327 1139
rect 3715 1131 3719 1135
rect 3883 1135 3887 1139
rect 719 1119 723 1123
rect 387 1111 391 1115
rect 563 1111 567 1115
rect 675 1111 679 1115
rect 907 1111 911 1115
rect 1043 1111 1047 1115
rect 1363 1111 1367 1115
rect 1499 1111 1503 1115
rect 2475 1115 2479 1119
rect 2483 1115 2487 1119
rect 2579 1115 2583 1119
rect 2675 1115 2679 1119
rect 2903 1115 2907 1119
rect 3135 1115 3136 1119
rect 3136 1115 3139 1119
rect 3171 1115 3175 1119
rect 3339 1115 3343 1119
rect 3579 1115 3583 1119
rect 3899 1115 3903 1119
rect 1239 1103 1243 1107
rect 3143 1107 3147 1111
rect 111 1092 115 1096
rect 375 1091 379 1095
rect 487 1091 491 1095
rect 599 1091 603 1095
rect 711 1091 715 1095
rect 831 1091 835 1095
rect 967 1091 971 1095
rect 1119 1091 1123 1095
rect 1279 1091 1283 1095
rect 1447 1091 1451 1095
rect 1623 1091 1627 1095
rect 2007 1092 2011 1096
rect 2047 1096 2051 1100
rect 2407 1095 2411 1099
rect 2503 1095 2507 1099
rect 2599 1095 2603 1099
rect 2695 1095 2699 1099
rect 2807 1095 2811 1099
rect 2943 1095 2947 1099
rect 3095 1095 3099 1099
rect 3263 1095 3267 1099
rect 3447 1095 3451 1099
rect 3639 1095 3643 1099
rect 3839 1095 3843 1099
rect 3943 1096 3947 1100
rect 451 1083 455 1087
rect 563 1083 567 1087
rect 675 1083 679 1087
rect 111 1075 115 1079
rect 787 1079 791 1083
rect 907 1083 911 1087
rect 1043 1083 1047 1087
rect 1195 1083 1199 1087
rect 1239 1083 1243 1087
rect 1363 1083 1367 1087
rect 1583 1083 1587 1087
rect 2483 1087 2487 1091
rect 2579 1087 2583 1091
rect 2675 1087 2679 1091
rect 2683 1087 2687 1091
rect 375 1072 379 1076
rect 487 1072 491 1076
rect 599 1072 603 1076
rect 711 1072 715 1076
rect 831 1072 835 1076
rect 967 1072 971 1076
rect 1119 1072 1123 1076
rect 1279 1072 1283 1076
rect 1447 1072 1451 1076
rect 1623 1072 1627 1076
rect 2007 1075 2011 1079
rect 2047 1079 2051 1083
rect 2895 1083 2899 1087
rect 2903 1087 2907 1091
rect 3171 1087 3175 1091
rect 3339 1087 3343 1091
rect 3383 1087 3387 1091
rect 3715 1087 3719 1091
rect 3915 1083 3919 1087
rect 2407 1076 2411 1080
rect 2503 1076 2507 1080
rect 2599 1076 2603 1080
rect 2695 1076 2699 1080
rect 2807 1076 2811 1080
rect 2943 1076 2947 1080
rect 3095 1076 3099 1080
rect 3263 1076 3267 1080
rect 3447 1076 3451 1080
rect 3639 1076 3643 1080
rect 3839 1076 3843 1080
rect 3943 1079 3947 1083
rect 111 1009 115 1013
rect 303 1012 307 1016
rect 447 1012 451 1016
rect 591 1012 595 1016
rect 727 1012 731 1016
rect 855 1012 859 1016
rect 975 1012 979 1016
rect 1087 1012 1091 1016
rect 1199 1012 1203 1016
rect 1311 1012 1315 1016
rect 1431 1012 1435 1016
rect 2007 1009 2011 1013
rect 2047 1009 2051 1013
rect 2455 1012 2459 1016
rect 2551 1012 2555 1016
rect 2647 1012 2651 1016
rect 2759 1012 2763 1016
rect 2887 1012 2891 1016
rect 3031 1012 3035 1016
rect 3183 1012 3187 1016
rect 3343 1012 3347 1016
rect 3503 1012 3507 1016
rect 3671 1012 3675 1016
rect 3839 1012 3843 1016
rect 3943 1009 3947 1013
rect 387 1003 391 1007
rect 395 1003 399 1007
rect 667 1003 671 1007
rect 803 1003 807 1007
rect 811 1003 815 1007
rect 1051 1003 1055 1007
rect 1163 1003 1167 1007
rect 1275 1003 1279 1007
rect 1387 1003 1391 1007
rect 1499 1003 1503 1007
rect 2543 1003 2547 1007
rect 2723 1003 2727 1007
rect 2835 1003 2839 1007
rect 2859 1003 2863 1007
rect 2991 1003 2995 1007
rect 3143 1003 3147 1007
rect 3295 1003 3299 1007
rect 3579 1003 3583 1007
rect 3907 1003 3911 1007
rect 111 992 115 996
rect 303 993 307 997
rect 447 993 451 997
rect 591 993 595 997
rect 727 993 731 997
rect 855 993 859 997
rect 975 993 979 997
rect 1087 993 1091 997
rect 1199 993 1203 997
rect 1311 993 1315 997
rect 1431 993 1435 997
rect 2007 992 2011 996
rect 2047 992 2051 996
rect 2455 993 2459 997
rect 2551 993 2555 997
rect 2647 993 2651 997
rect 2759 993 2763 997
rect 2887 993 2891 997
rect 3031 993 3035 997
rect 3183 993 3187 997
rect 3343 993 3347 997
rect 3503 993 3507 997
rect 3671 993 3675 997
rect 3839 993 3843 997
rect 3943 992 3947 996
rect 395 975 399 979
rect 523 971 527 975
rect 811 983 815 987
rect 787 975 791 979
rect 803 975 807 979
rect 1043 971 1047 975
rect 1051 975 1055 979
rect 1163 975 1167 979
rect 1275 975 1279 979
rect 1387 975 1391 979
rect 2543 975 2547 979
rect 2683 983 2687 987
rect 2859 979 2863 983
rect 2787 971 2791 975
rect 2895 975 2899 979
rect 2943 971 2947 975
rect 3295 975 3299 979
rect 3383 975 3384 979
rect 3384 975 3387 979
rect 3723 971 3727 975
rect 3915 975 3919 979
rect 323 959 327 963
rect 331 959 335 963
rect 667 959 668 963
rect 668 959 671 963
rect 707 959 711 963
rect 883 959 887 963
rect 1211 959 1215 963
rect 1355 959 1359 963
rect 1499 959 1503 963
rect 1635 959 1639 963
rect 1735 959 1736 963
rect 1736 959 1739 963
rect 2499 955 2503 959
rect 2595 955 2599 959
rect 2723 955 2727 959
rect 2835 955 2839 959
rect 2991 955 2992 959
rect 2992 955 2995 959
rect 3047 955 3051 959
rect 3687 955 3688 959
rect 3688 955 3691 959
rect 3907 955 3911 959
rect 111 940 115 944
rect 255 939 259 943
rect 447 939 451 943
rect 631 939 635 943
rect 807 939 811 943
rect 975 939 979 943
rect 331 931 335 935
rect 523 931 527 935
rect 707 931 711 935
rect 883 931 887 935
rect 1043 935 1047 939
rect 1127 939 1131 943
rect 1271 939 1275 943
rect 1415 939 1419 943
rect 1551 939 1555 943
rect 1695 939 1699 943
rect 2007 940 2011 944
rect 2047 936 2051 940
rect 111 923 115 927
rect 1051 927 1055 931
rect 1211 931 1215 935
rect 1355 931 1359 935
rect 1499 931 1503 935
rect 2423 935 2427 939
rect 1635 931 1639 935
rect 2519 935 2523 939
rect 2615 935 2619 939
rect 2711 935 2715 939
rect 2823 935 2827 939
rect 2951 935 2955 939
rect 3103 935 3107 939
rect 3271 935 3275 939
rect 3455 935 3459 939
rect 3647 935 3651 939
rect 3839 935 3843 939
rect 3943 936 3947 940
rect 255 920 259 924
rect 447 920 451 924
rect 631 920 635 924
rect 807 920 811 924
rect 975 920 979 924
rect 1127 920 1131 924
rect 1271 920 1275 924
rect 1415 920 1419 924
rect 1551 920 1555 924
rect 1695 920 1699 924
rect 2007 923 2011 927
rect 2499 927 2503 931
rect 2595 927 2599 931
rect 2047 919 2051 923
rect 2691 923 2695 927
rect 2787 927 2791 931
rect 2943 927 2947 931
rect 3047 927 3051 931
rect 3411 927 3415 931
rect 3723 927 3727 931
rect 3915 923 3919 927
rect 2423 916 2427 920
rect 2519 916 2523 920
rect 2615 916 2619 920
rect 2711 916 2715 920
rect 2823 916 2827 920
rect 2951 916 2955 920
rect 3103 916 3107 920
rect 3271 916 3275 920
rect 3455 916 3459 920
rect 3647 916 3651 920
rect 3839 916 3843 920
rect 3943 919 3947 923
rect 111 853 115 857
rect 255 856 259 860
rect 447 856 451 860
rect 639 856 643 860
rect 823 856 827 860
rect 999 856 1003 860
rect 1167 856 1171 860
rect 1327 856 1331 860
rect 1479 856 1483 860
rect 1631 856 1635 860
rect 1783 856 1787 860
rect 2007 853 2011 857
rect 2047 853 2051 857
rect 2343 856 2347 860
rect 2439 856 2443 860
rect 2535 856 2539 860
rect 2631 856 2635 860
rect 2735 856 2739 860
rect 2863 856 2867 860
rect 3015 856 3019 860
rect 3191 856 3195 860
rect 3391 856 3395 860
rect 3607 856 3611 860
rect 3823 856 3827 860
rect 3943 853 3947 857
rect 323 847 327 851
rect 515 847 519 851
rect 567 847 571 851
rect 771 847 775 851
rect 1243 847 1247 851
rect 1403 847 1407 851
rect 1555 847 1559 851
rect 1707 847 1711 851
rect 1735 847 1739 851
rect 2431 847 2435 851
rect 2527 847 2531 851
rect 2707 847 2711 851
rect 2715 847 2719 851
rect 2939 847 2943 851
rect 3091 847 3095 851
rect 3267 847 3271 851
rect 3467 847 3471 851
rect 3475 847 3479 851
rect 3891 847 3895 851
rect 111 836 115 840
rect 255 837 259 841
rect 447 837 451 841
rect 639 837 643 841
rect 823 837 827 841
rect 999 837 1003 841
rect 1167 837 1171 841
rect 1327 837 1331 841
rect 1479 837 1483 841
rect 1631 837 1635 841
rect 1783 837 1787 841
rect 2007 836 2011 840
rect 2047 836 2051 840
rect 2343 837 2347 841
rect 2439 837 2443 841
rect 2535 837 2539 841
rect 2631 837 2635 841
rect 2735 837 2739 841
rect 2863 837 2867 841
rect 3015 837 3019 841
rect 3191 837 3195 841
rect 3391 837 3395 841
rect 3607 837 3611 841
rect 3823 837 3827 841
rect 3943 836 3947 840
rect 235 815 239 819
rect 567 819 571 823
rect 771 819 775 823
rect 1051 819 1055 823
rect 1243 819 1247 823
rect 1403 819 1407 823
rect 1555 819 1559 823
rect 1707 819 1711 823
rect 2431 819 2435 823
rect 2527 819 2531 823
rect 2715 827 2719 831
rect 2691 819 2695 823
rect 2707 819 2711 823
rect 3411 827 3415 831
rect 2939 819 2943 823
rect 3091 819 3095 823
rect 3267 819 3271 823
rect 3467 819 3471 823
rect 3915 819 3919 823
rect 1519 811 1523 815
rect 3475 811 3479 815
rect 339 799 343 803
rect 511 799 512 803
rect 512 799 515 803
rect 547 799 551 803
rect 699 799 703 803
rect 975 799 976 803
rect 976 799 979 803
rect 1011 799 1015 803
rect 1231 799 1235 803
rect 1375 799 1379 803
rect 1491 799 1495 803
rect 1835 799 1839 803
rect 1987 799 1991 803
rect 2387 803 2391 807
rect 2571 803 2575 807
rect 2955 803 2959 807
rect 3155 803 3159 807
rect 3363 803 3367 807
rect 3771 803 3775 807
rect 111 780 115 784
rect 159 779 163 783
rect 311 779 315 783
rect 471 779 475 783
rect 623 779 627 783
rect 775 779 779 783
rect 935 779 939 783
rect 1095 779 1099 783
rect 1255 779 1259 783
rect 1415 779 1419 783
rect 1583 779 1587 783
rect 1751 779 1755 783
rect 1903 779 1907 783
rect 2007 780 2011 784
rect 2047 784 2051 788
rect 2311 783 2315 787
rect 2495 783 2499 787
rect 2687 783 2691 787
rect 2879 783 2883 787
rect 3079 783 3083 787
rect 3287 783 3291 787
rect 3503 783 3507 787
rect 3719 783 3723 787
rect 3943 784 3947 788
rect 235 771 239 775
rect 547 771 551 775
rect 699 771 703 775
rect 111 763 115 767
rect 851 767 855 771
rect 1011 771 1015 775
rect 1231 771 1235 775
rect 1375 771 1379 775
rect 1491 771 1495 775
rect 1519 771 1523 775
rect 1827 767 1831 771
rect 1835 771 1839 775
rect 2387 775 2391 779
rect 2571 775 2575 779
rect 2955 775 2959 779
rect 3155 775 3159 779
rect 3363 775 3367 779
rect 3447 775 3451 779
rect 3687 775 3691 779
rect 159 760 163 764
rect 311 760 315 764
rect 471 760 475 764
rect 623 760 627 764
rect 775 760 779 764
rect 935 760 939 764
rect 1095 760 1099 764
rect 1255 760 1259 764
rect 1415 760 1419 764
rect 1583 760 1587 764
rect 1751 760 1755 764
rect 1903 760 1907 764
rect 2007 763 2011 767
rect 2047 767 2051 771
rect 2311 764 2315 768
rect 2495 764 2499 768
rect 2687 764 2691 768
rect 2879 764 2883 768
rect 3079 764 3083 768
rect 3287 764 3291 768
rect 3503 764 3507 768
rect 3719 764 3723 768
rect 3943 767 3947 771
rect 111 697 115 701
rect 135 700 139 704
rect 263 700 267 704
rect 431 700 435 704
rect 623 700 627 704
rect 823 700 827 704
rect 1015 700 1019 704
rect 1207 700 1211 704
rect 1391 700 1395 704
rect 1567 700 1571 704
rect 1743 700 1747 704
rect 1903 700 1907 704
rect 2007 697 2011 701
rect 2047 697 2051 701
rect 2071 700 2075 704
rect 2255 700 2259 704
rect 2455 700 2459 704
rect 2655 700 2659 704
rect 2855 700 2859 704
rect 3047 700 3051 704
rect 3239 700 3243 704
rect 3439 700 3443 704
rect 3639 700 3643 704
rect 3839 700 3843 704
rect 3943 697 3947 701
rect 211 691 215 695
rect 339 691 343 695
rect 423 691 427 695
rect 543 691 547 695
rect 707 691 711 695
rect 975 691 979 695
rect 1467 691 1471 695
rect 1643 691 1647 695
rect 1651 691 1655 695
rect 111 680 115 684
rect 135 681 139 685
rect 263 681 267 685
rect 431 681 435 685
rect 623 681 627 685
rect 823 681 827 685
rect 1015 681 1019 685
rect 1207 681 1211 685
rect 1391 681 1395 685
rect 1567 681 1571 685
rect 1743 681 1747 685
rect 1811 683 1815 687
rect 1987 691 1991 695
rect 2339 691 2343 695
rect 2731 691 2735 695
rect 2931 691 2935 695
rect 3123 691 3127 695
rect 3315 691 3319 695
rect 3515 691 3519 695
rect 3559 691 3563 695
rect 3907 691 3911 695
rect 1903 681 1907 685
rect 2007 680 2011 684
rect 2047 680 2051 684
rect 2071 681 2075 685
rect 2255 681 2259 685
rect 2455 681 2459 685
rect 2655 681 2659 685
rect 2855 681 2859 685
rect 3047 681 3051 685
rect 3239 681 3243 685
rect 3439 681 3443 685
rect 3639 681 3643 685
rect 3839 681 3843 685
rect 3943 680 3947 684
rect 211 663 215 667
rect 543 663 547 667
rect 707 663 711 667
rect 851 663 855 667
rect 211 655 215 659
rect 1651 671 1655 675
rect 1467 663 1471 667
rect 1811 663 1815 667
rect 1827 663 1831 667
rect 2339 663 2343 667
rect 2507 659 2511 663
rect 3447 671 3451 675
rect 2931 663 2935 667
rect 3123 663 3127 667
rect 3315 663 3319 667
rect 3515 663 3519 667
rect 3891 663 3895 667
rect 3559 655 3563 659
rect 219 647 223 651
rect 287 647 288 651
rect 288 647 291 651
rect 423 647 424 651
rect 424 647 427 651
rect 459 647 463 651
rect 603 647 607 651
rect 911 647 912 651
rect 912 647 915 651
rect 947 647 951 651
rect 1155 647 1159 651
rect 1379 647 1383 651
rect 1643 647 1647 651
rect 2111 647 2112 651
rect 2112 647 2115 651
rect 2147 647 2151 651
rect 2307 647 2311 651
rect 2723 647 2727 651
rect 2731 647 2735 651
rect 3099 647 3103 651
rect 3283 647 3287 651
rect 3451 647 3455 651
rect 3779 647 3783 651
rect 3907 647 3911 651
rect 111 628 115 632
rect 135 627 139 631
rect 247 627 251 631
rect 383 627 387 631
rect 527 627 531 631
rect 687 627 691 631
rect 871 627 875 631
rect 1079 627 1083 631
rect 1303 627 1307 631
rect 1543 627 1547 631
rect 1783 627 1787 631
rect 2007 628 2011 632
rect 2047 628 2051 632
rect 2071 627 2075 631
rect 2231 627 2235 631
rect 2431 627 2435 631
rect 2631 627 2635 631
rect 2831 627 2835 631
rect 3023 627 3027 631
rect 3207 627 3211 631
rect 3375 627 3379 631
rect 3535 627 3539 631
rect 3695 627 3699 631
rect 3839 627 3843 631
rect 3943 628 3947 632
rect 211 619 215 623
rect 219 619 223 623
rect 459 619 463 623
rect 603 619 607 623
rect 111 611 115 615
rect 763 615 767 619
rect 947 619 951 623
rect 1155 619 1159 623
rect 1379 619 1383 623
rect 2147 619 2151 623
rect 2307 619 2311 623
rect 2507 619 2511 623
rect 2599 619 2603 623
rect 2723 619 2727 623
rect 3099 619 3103 623
rect 3283 619 3287 623
rect 3451 619 3455 623
rect 135 608 139 612
rect 247 608 251 612
rect 383 608 387 612
rect 527 608 531 612
rect 687 608 691 612
rect 871 608 875 612
rect 1079 608 1083 612
rect 1303 608 1307 612
rect 1543 608 1547 612
rect 1783 608 1787 612
rect 1851 611 1855 615
rect 2007 611 2011 615
rect 2047 611 2051 615
rect 3611 615 3615 619
rect 3771 619 3775 623
rect 3915 615 3919 619
rect 2071 608 2075 612
rect 2231 608 2235 612
rect 2431 608 2435 612
rect 2631 608 2635 612
rect 2831 608 2835 612
rect 3023 608 3027 612
rect 3207 608 3211 612
rect 3375 608 3379 612
rect 3535 608 3539 612
rect 3695 608 3699 612
rect 3839 608 3843 612
rect 3943 611 3947 615
rect 2111 551 2115 555
rect 111 541 115 545
rect 135 544 139 548
rect 295 544 299 548
rect 479 544 483 548
rect 663 544 667 548
rect 847 544 851 548
rect 1031 544 1035 548
rect 1215 544 1219 548
rect 1399 544 1403 548
rect 1591 544 1595 548
rect 1783 544 1787 548
rect 2007 541 2011 545
rect 2047 541 2051 545
rect 2071 544 2075 548
rect 2215 544 2219 548
rect 231 535 235 539
rect 287 535 291 539
rect 915 535 919 539
rect 1107 535 1111 539
rect 1115 535 1119 539
rect 1467 535 1471 539
rect 1727 535 1731 539
rect 2139 535 2143 539
rect 2399 544 2403 548
rect 2583 544 2587 548
rect 2775 544 2779 548
rect 2959 544 2963 548
rect 3143 544 3147 548
rect 3319 544 3323 548
rect 3495 544 3499 548
rect 3679 544 3683 548
rect 3839 544 3843 548
rect 3943 541 3947 545
rect 2531 535 2535 539
rect 3035 535 3039 539
rect 3231 535 3235 539
rect 3239 535 3243 539
rect 3907 535 3911 539
rect 111 524 115 528
rect 135 525 139 529
rect 295 525 299 529
rect 479 525 483 529
rect 663 525 667 529
rect 847 525 851 529
rect 1031 525 1035 529
rect 1215 525 1219 529
rect 1399 525 1403 529
rect 1591 525 1595 529
rect 1783 525 1787 529
rect 2007 524 2011 528
rect 2047 524 2051 528
rect 2071 525 2075 529
rect 2215 525 2219 529
rect 2399 525 2403 529
rect 2583 525 2587 529
rect 2775 525 2779 529
rect 2959 525 2963 529
rect 3143 525 3147 529
rect 3319 525 3323 529
rect 3495 525 3499 529
rect 3679 525 3683 529
rect 3839 525 3843 529
rect 3943 524 3947 528
rect 211 503 215 507
rect 231 507 235 511
rect 763 507 767 511
rect 1115 515 1119 519
rect 979 503 983 507
rect 1107 507 1111 511
rect 1727 507 1731 511
rect 1851 507 1855 511
rect 2599 515 2603 519
rect 2531 507 2535 511
rect 2803 503 2807 507
rect 3239 515 3243 519
rect 3035 507 3039 511
rect 3611 507 3615 511
rect 3915 507 3919 511
rect 247 491 251 495
rect 355 491 359 495
rect 531 491 535 495
rect 691 491 695 495
rect 971 491 975 495
rect 1107 491 1111 495
rect 1235 491 1239 495
rect 1467 491 1471 495
rect 1407 483 1411 487
rect 2139 487 2143 491
rect 2263 487 2264 491
rect 2264 487 2267 491
rect 2299 487 2303 491
rect 2467 487 2471 491
rect 2635 487 2639 491
rect 2979 487 2983 491
rect 3119 487 3123 491
rect 3231 487 3235 491
rect 3299 487 3303 491
rect 3619 487 3623 491
rect 3907 487 3911 491
rect 3799 479 3803 483
rect 111 472 115 476
rect 135 471 139 475
rect 287 471 291 475
rect 455 471 459 475
rect 615 471 619 475
rect 767 471 771 475
rect 903 471 907 475
rect 1031 471 1035 475
rect 1159 471 1163 475
rect 1287 471 1291 475
rect 1415 471 1419 475
rect 2007 472 2011 476
rect 2047 468 2051 472
rect 211 463 215 467
rect 247 463 251 467
rect 531 463 535 467
rect 691 463 695 467
rect 111 455 115 459
rect 843 459 847 463
rect 979 463 983 467
rect 1107 463 1111 467
rect 1235 463 1239 467
rect 2071 467 2075 471
rect 1399 459 1403 463
rect 1407 463 1411 467
rect 2223 467 2227 471
rect 2391 467 2395 471
rect 2559 467 2563 471
rect 2727 467 2731 471
rect 2895 467 2899 471
rect 3063 467 3067 471
rect 3223 467 3227 471
rect 3383 467 3387 471
rect 3543 467 3547 471
rect 3703 467 3707 471
rect 3839 467 3843 471
rect 3943 468 3947 472
rect 135 452 139 456
rect 287 452 291 456
rect 455 452 459 456
rect 615 452 619 456
rect 767 452 771 456
rect 903 452 907 456
rect 1031 452 1035 456
rect 1159 452 1163 456
rect 1287 452 1291 456
rect 1415 452 1419 456
rect 2007 455 2011 459
rect 2035 459 2039 463
rect 2299 459 2303 463
rect 2467 459 2471 463
rect 2635 459 2639 463
rect 2803 459 2807 463
rect 2887 459 2891 463
rect 2979 459 2983 463
rect 3299 459 3303 463
rect 3319 459 3323 463
rect 3619 459 3623 463
rect 3779 459 3783 463
rect 3799 459 3803 463
rect 2047 451 2051 455
rect 2071 448 2075 452
rect 2223 448 2227 452
rect 2391 448 2395 452
rect 2559 448 2563 452
rect 2727 448 2731 452
rect 2895 448 2899 452
rect 3063 448 3067 452
rect 3223 448 3227 452
rect 3383 448 3387 452
rect 3543 448 3547 452
rect 3703 448 3707 452
rect 3839 448 3843 452
rect 3943 451 3947 455
rect 111 389 115 393
rect 135 392 139 396
rect 287 392 291 396
rect 447 392 451 396
rect 599 392 603 396
rect 751 392 755 396
rect 903 392 907 396
rect 1079 392 1083 396
rect 1271 392 1275 396
rect 1479 392 1483 396
rect 1703 392 1707 396
rect 1903 392 1907 396
rect 2007 389 2011 393
rect 211 383 215 387
rect 355 383 359 387
rect 523 383 527 387
rect 531 383 535 387
rect 683 383 687 387
rect 971 383 975 387
rect 1211 383 1215 387
rect 1555 383 1559 387
rect 1639 383 1643 387
rect 1971 383 1975 387
rect 2047 385 2051 389
rect 2463 388 2467 392
rect 2559 388 2563 392
rect 2655 388 2659 392
rect 2751 388 2755 392
rect 2847 388 2851 392
rect 2943 388 2947 392
rect 3039 388 3043 392
rect 3135 388 3139 392
rect 3231 388 3235 392
rect 3943 385 3947 389
rect 2263 379 2267 383
rect 2551 379 2555 383
rect 2647 379 2651 383
rect 2743 379 2747 383
rect 2923 379 2927 383
rect 3019 379 3023 383
rect 3115 379 3119 383
rect 3211 379 3215 383
rect 3299 379 3303 383
rect 111 372 115 376
rect 135 373 139 377
rect 287 373 291 377
rect 447 373 451 377
rect 599 373 603 377
rect 751 373 755 377
rect 903 373 907 377
rect 1079 373 1083 377
rect 1271 373 1275 377
rect 1479 373 1483 377
rect 1703 373 1707 377
rect 1903 373 1907 377
rect 2007 372 2011 376
rect 2047 368 2051 372
rect 2463 369 2467 373
rect 2559 369 2563 373
rect 2655 369 2659 373
rect 2751 369 2755 373
rect 2847 369 2851 373
rect 2943 369 2947 373
rect 3039 369 3043 373
rect 3135 369 3139 373
rect 3231 369 3235 373
rect 3943 368 3947 372
rect 211 355 215 359
rect 531 355 535 359
rect 683 355 687 359
rect 843 355 847 359
rect 1211 355 1215 359
rect 1235 351 1239 355
rect 1399 355 1403 359
rect 1555 355 1559 359
rect 2035 355 2039 359
rect 2551 351 2555 355
rect 2647 351 2651 355
rect 2743 351 2747 355
rect 1639 343 1643 347
rect 2859 347 2863 351
rect 2887 351 2888 355
rect 2888 351 2891 355
rect 2923 351 2927 355
rect 3019 351 3023 355
rect 3115 351 3119 355
rect 3211 351 3215 355
rect 243 335 247 339
rect 523 335 527 339
rect 627 335 631 339
rect 835 335 839 339
rect 1419 335 1423 339
rect 1603 335 1607 339
rect 1971 335 1975 339
rect 2439 335 2440 339
rect 2440 335 2443 339
rect 2475 335 2479 339
rect 2579 335 2583 339
rect 2699 335 2703 339
rect 2835 335 2839 339
rect 3155 335 3159 339
rect 3299 335 3303 339
rect 3559 335 3563 339
rect 3683 335 3687 339
rect 1819 327 1823 331
rect 3499 327 3503 331
rect 111 316 115 320
rect 159 315 163 319
rect 351 315 355 319
rect 551 315 555 319
rect 759 315 763 319
rect 959 315 963 319
rect 1159 315 1163 319
rect 1343 315 1347 319
rect 1527 315 1531 319
rect 1711 315 1715 319
rect 1895 315 1899 319
rect 2007 316 2011 320
rect 2047 316 2051 320
rect 2399 315 2403 319
rect 2503 315 2507 319
rect 2623 315 2627 319
rect 2759 315 2763 319
rect 2911 315 2915 319
rect 3071 315 3075 319
rect 3247 315 3251 319
rect 3423 315 3427 319
rect 3607 315 3611 319
rect 3791 315 3795 319
rect 3943 316 3947 320
rect 243 307 247 311
rect 627 307 631 311
rect 835 307 839 311
rect 903 307 907 311
rect 1235 307 1239 311
rect 1419 307 1423 311
rect 1603 307 1607 311
rect 111 299 115 303
rect 1787 303 1791 307
rect 1819 307 1823 311
rect 2475 307 2479 311
rect 2579 307 2583 311
rect 2699 307 2703 311
rect 2835 307 2839 311
rect 2859 307 2863 311
rect 3003 307 3007 311
rect 3155 307 3159 311
rect 3499 307 3503 311
rect 3683 307 3687 311
rect 159 296 163 300
rect 351 296 355 300
rect 551 296 555 300
rect 759 296 763 300
rect 959 296 963 300
rect 1159 296 1163 300
rect 1343 296 1347 300
rect 1527 296 1531 300
rect 1711 296 1715 300
rect 1895 296 1899 300
rect 2007 299 2011 303
rect 2047 299 2051 303
rect 3867 303 3871 307
rect 2399 296 2403 300
rect 2503 296 2507 300
rect 2623 296 2627 300
rect 2759 296 2763 300
rect 2911 296 2915 300
rect 3071 296 3075 300
rect 3247 296 3251 300
rect 3423 296 3427 300
rect 3607 296 3611 300
rect 3791 296 3795 300
rect 3943 299 3947 303
rect 2439 243 2443 247
rect 2047 233 2051 237
rect 2191 236 2195 240
rect 2351 236 2355 240
rect 2519 236 2523 240
rect 111 225 115 229
rect 223 228 227 232
rect 383 228 387 232
rect 543 228 547 232
rect 703 228 707 232
rect 863 228 867 232
rect 1031 228 1035 232
rect 1199 228 1203 232
rect 1367 228 1371 232
rect 1543 228 1547 232
rect 1727 228 1731 232
rect 1903 228 1907 232
rect 2007 225 2011 229
rect 2267 227 2271 231
rect 2427 227 2431 231
rect 2595 227 2599 231
rect 2687 236 2691 240
rect 2855 236 2859 240
rect 3031 236 3035 240
rect 3215 236 3219 240
rect 3407 236 3411 240
rect 3607 236 3611 240
rect 3807 236 3811 240
rect 3943 233 3947 237
rect 2931 227 2935 231
rect 3107 227 3111 231
rect 3291 227 3295 231
rect 3379 227 3383 231
rect 3559 227 3563 231
rect 3783 227 3787 231
rect 299 219 303 223
rect 619 219 623 223
rect 799 219 803 223
rect 1099 219 1103 223
rect 1115 219 1119 223
rect 1627 219 1631 223
rect 1971 219 1975 223
rect 2047 216 2051 220
rect 2191 217 2195 221
rect 2351 217 2355 221
rect 2519 217 2523 221
rect 2687 217 2691 221
rect 2855 217 2859 221
rect 3031 217 3035 221
rect 3215 217 3219 221
rect 3407 217 3411 221
rect 3607 217 3611 221
rect 3807 217 3811 221
rect 3943 216 3947 220
rect 111 208 115 212
rect 223 209 227 213
rect 383 209 387 213
rect 543 209 547 213
rect 703 209 707 213
rect 863 209 867 213
rect 1031 209 1035 213
rect 1199 209 1203 213
rect 1367 209 1371 213
rect 1543 209 1547 213
rect 1727 209 1731 213
rect 1903 209 1907 213
rect 2007 208 2011 212
rect 299 191 303 195
rect 799 191 803 195
rect 903 191 904 195
rect 904 191 907 195
rect 1115 191 1119 195
rect 1627 191 1631 195
rect 1787 191 1791 195
rect 2267 199 2271 203
rect 2427 199 2431 203
rect 2595 199 2599 203
rect 3003 207 3007 211
rect 2931 199 2935 203
rect 3107 199 3111 203
rect 3291 199 3295 203
rect 307 183 311 187
rect 1883 187 1887 191
rect 3867 199 3871 203
rect 2727 187 2731 191
rect 211 155 215 159
rect 411 155 415 159
rect 507 155 511 159
rect 619 155 623 159
rect 723 155 727 159
rect 851 155 855 159
rect 1099 155 1103 159
rect 1107 155 1111 159
rect 1227 155 1231 159
rect 1347 155 1351 159
rect 1459 155 1463 159
rect 1563 155 1567 159
rect 1667 155 1671 159
rect 1779 155 1783 159
rect 1971 155 1975 159
rect 3379 159 3383 163
rect 315 147 319 151
rect 859 147 863 151
rect 1979 151 1983 155
rect 2147 151 2151 155
rect 2243 151 2247 155
rect 2339 151 2343 155
rect 2443 151 2447 155
rect 2563 151 2567 155
rect 2719 151 2723 155
rect 2947 151 2951 155
rect 3067 151 3071 155
rect 3187 151 3191 155
rect 3299 151 3303 155
rect 3507 151 3511 155
rect 3783 151 3784 155
rect 3784 151 3787 155
rect 3819 151 3823 155
rect 111 136 115 140
rect 135 135 139 139
rect 231 135 235 139
rect 327 135 331 139
rect 423 135 427 139
rect 527 135 531 139
rect 647 135 651 139
rect 775 135 779 139
rect 903 135 907 139
rect 1031 135 1035 139
rect 1151 135 1155 139
rect 1271 135 1275 139
rect 1383 135 1387 139
rect 1487 135 1491 139
rect 1591 135 1595 139
rect 1703 135 1707 139
rect 1807 135 1811 139
rect 1903 135 1907 139
rect 2007 136 2011 140
rect 2047 132 2051 136
rect 211 127 215 131
rect 307 127 311 131
rect 315 127 319 131
rect 411 127 415 131
rect 507 127 511 131
rect 723 127 727 131
rect 851 127 855 131
rect 859 127 863 131
rect 1107 127 1111 131
rect 1227 127 1231 131
rect 1347 127 1351 131
rect 1459 127 1463 131
rect 1563 127 1567 131
rect 1667 127 1671 131
rect 1779 127 1783 131
rect 1883 127 1887 131
rect 2071 131 2075 135
rect 1979 127 1983 131
rect 2167 131 2171 135
rect 2263 131 2267 135
rect 2367 131 2371 135
rect 2487 131 2491 135
rect 2615 131 2619 135
rect 2743 131 2747 135
rect 2871 131 2875 135
rect 2991 131 2995 135
rect 3111 131 3115 135
rect 3223 131 3227 135
rect 3327 131 3331 135
rect 3431 131 3435 135
rect 3535 131 3539 135
rect 3639 131 3643 135
rect 3743 131 3747 135
rect 3839 131 3843 135
rect 3943 132 3947 136
rect 111 119 115 123
rect 135 116 139 120
rect 231 116 235 120
rect 327 116 331 120
rect 423 116 427 120
rect 527 116 531 120
rect 647 116 651 120
rect 775 116 779 120
rect 903 116 907 120
rect 1031 116 1035 120
rect 1151 116 1155 120
rect 1271 116 1275 120
rect 1383 116 1387 120
rect 1487 116 1491 120
rect 1591 116 1595 120
rect 1703 116 1707 120
rect 1807 116 1811 120
rect 1903 116 1907 120
rect 2007 119 2011 123
rect 2147 123 2151 127
rect 2243 123 2247 127
rect 2339 123 2343 127
rect 2443 123 2447 127
rect 2563 123 2567 127
rect 2719 123 2723 127
rect 2727 123 2731 127
rect 2947 123 2951 127
rect 3067 123 3071 127
rect 3187 123 3191 127
rect 3299 123 3303 127
rect 3507 123 3511 127
rect 3819 123 3823 127
rect 2047 115 2051 119
rect 2071 112 2075 116
rect 2167 112 2171 116
rect 2263 112 2267 116
rect 2367 112 2371 116
rect 2487 112 2491 116
rect 2615 112 2619 116
rect 2743 112 2747 116
rect 2871 112 2875 116
rect 2991 112 2995 116
rect 3111 112 3115 116
rect 3223 112 3227 116
rect 3327 112 3331 116
rect 3431 112 3435 116
rect 3535 112 3539 116
rect 3639 112 3643 116
rect 3743 112 3747 116
rect 3839 112 3843 116
rect 3943 115 3947 119
<< m3 >>
rect 2047 4030 2051 4031
rect 2047 4025 2051 4026
rect 2071 4030 2075 4031
rect 2071 4025 2075 4026
rect 3943 4030 3947 4031
rect 3943 4025 3947 4026
rect 1978 4023 1984 4024
rect 1978 4019 1979 4023
rect 1983 4019 1984 4023
rect 1978 4018 1984 4019
rect 111 4010 115 4011
rect 111 4005 115 4006
rect 151 4010 155 4011
rect 151 4005 155 4006
rect 279 4010 283 4011
rect 279 4005 283 4006
rect 431 4010 435 4011
rect 431 4005 435 4006
rect 607 4010 611 4011
rect 607 4005 611 4006
rect 791 4010 795 4011
rect 791 4005 795 4006
rect 975 4010 979 4011
rect 975 4005 979 4006
rect 1151 4010 1155 4011
rect 1151 4005 1155 4006
rect 1311 4010 1315 4011
rect 1311 4005 1315 4006
rect 1471 4010 1475 4011
rect 1471 4005 1475 4006
rect 1623 4010 1627 4011
rect 1623 4005 1627 4006
rect 1775 4010 1779 4011
rect 1775 4005 1779 4006
rect 1903 4010 1907 4011
rect 1903 4005 1907 4006
rect 112 3985 114 4005
rect 110 3984 116 3985
rect 152 3984 154 4005
rect 226 4003 232 4004
rect 226 3999 227 4003
rect 231 3999 232 4003
rect 226 3998 232 3999
rect 110 3980 111 3984
rect 115 3980 116 3984
rect 110 3979 116 3980
rect 150 3983 156 3984
rect 150 3979 151 3983
rect 155 3979 156 3983
rect 150 3978 156 3979
rect 228 3976 230 3998
rect 280 3984 282 4005
rect 354 4003 360 4004
rect 354 3999 355 4003
rect 359 3999 360 4003
rect 354 3998 360 3999
rect 278 3983 284 3984
rect 278 3979 279 3983
rect 283 3979 284 3983
rect 278 3978 284 3979
rect 356 3976 358 3998
rect 432 3984 434 4005
rect 506 4003 512 4004
rect 506 3999 507 4003
rect 511 3999 512 4003
rect 506 3998 512 3999
rect 430 3983 436 3984
rect 430 3979 431 3983
rect 435 3979 436 3983
rect 430 3978 436 3979
rect 508 3976 510 3998
rect 608 3984 610 4005
rect 682 4003 688 4004
rect 682 3999 683 4003
rect 687 3999 688 4003
rect 682 3998 688 3999
rect 606 3983 612 3984
rect 606 3979 607 3983
rect 611 3979 612 3983
rect 606 3978 612 3979
rect 684 3976 686 3998
rect 792 3984 794 4005
rect 866 4003 872 4004
rect 866 3999 867 4003
rect 871 3999 872 4003
rect 866 3998 872 3999
rect 790 3983 796 3984
rect 790 3979 791 3983
rect 795 3979 796 3983
rect 790 3978 796 3979
rect 868 3976 870 3998
rect 976 3984 978 4005
rect 1152 3984 1154 4005
rect 1226 4003 1232 4004
rect 1226 3999 1227 4003
rect 1231 3999 1232 4003
rect 1226 3998 1232 3999
rect 974 3983 980 3984
rect 974 3979 975 3983
rect 979 3979 980 3983
rect 974 3978 980 3979
rect 1150 3983 1156 3984
rect 1150 3979 1151 3983
rect 1155 3979 1156 3983
rect 1150 3978 1156 3979
rect 1228 3976 1230 3998
rect 1312 3984 1314 4005
rect 1386 4003 1392 4004
rect 1386 3999 1387 4003
rect 1391 3999 1392 4003
rect 1386 3998 1392 3999
rect 1310 3983 1316 3984
rect 1310 3979 1311 3983
rect 1315 3979 1316 3983
rect 1310 3978 1316 3979
rect 1388 3976 1390 3998
rect 1410 3995 1416 3996
rect 1410 3991 1411 3995
rect 1415 3991 1416 3995
rect 1410 3990 1416 3991
rect 226 3975 232 3976
rect 226 3971 227 3975
rect 231 3971 232 3975
rect 226 3970 232 3971
rect 354 3975 360 3976
rect 354 3971 355 3975
rect 359 3971 360 3975
rect 354 3970 360 3971
rect 506 3975 512 3976
rect 506 3971 507 3975
rect 511 3971 512 3975
rect 506 3970 512 3971
rect 682 3975 688 3976
rect 682 3971 683 3975
rect 687 3971 688 3975
rect 682 3970 688 3971
rect 866 3975 872 3976
rect 866 3971 867 3975
rect 871 3971 872 3975
rect 866 3970 872 3971
rect 918 3975 924 3976
rect 918 3971 919 3975
rect 923 3971 924 3975
rect 918 3970 924 3971
rect 1226 3975 1232 3976
rect 1226 3971 1227 3975
rect 1231 3971 1232 3975
rect 1226 3970 1232 3971
rect 1386 3975 1392 3976
rect 1386 3971 1387 3975
rect 1391 3971 1392 3975
rect 1386 3970 1392 3971
rect 110 3967 116 3968
rect 110 3963 111 3967
rect 115 3963 116 3967
rect 110 3962 116 3963
rect 150 3964 156 3965
rect 112 3935 114 3962
rect 150 3960 151 3964
rect 155 3960 156 3964
rect 150 3959 156 3960
rect 278 3964 284 3965
rect 278 3960 279 3964
rect 283 3960 284 3964
rect 278 3959 284 3960
rect 430 3964 436 3965
rect 430 3960 431 3964
rect 435 3960 436 3964
rect 430 3959 436 3960
rect 606 3964 612 3965
rect 606 3960 607 3964
rect 611 3960 612 3964
rect 606 3959 612 3960
rect 790 3964 796 3965
rect 790 3960 791 3964
rect 795 3960 796 3964
rect 790 3959 796 3960
rect 152 3935 154 3959
rect 280 3935 282 3959
rect 432 3935 434 3959
rect 608 3935 610 3959
rect 792 3935 794 3959
rect 111 3934 115 3935
rect 111 3929 115 3930
rect 151 3934 155 3935
rect 151 3929 155 3930
rect 279 3934 283 3935
rect 279 3929 283 3930
rect 303 3934 307 3935
rect 303 3929 307 3930
rect 423 3934 427 3935
rect 423 3929 427 3930
rect 431 3934 435 3935
rect 431 3929 435 3930
rect 551 3934 555 3935
rect 551 3929 555 3930
rect 607 3934 611 3935
rect 607 3929 611 3930
rect 687 3934 691 3935
rect 687 3929 691 3930
rect 791 3934 795 3935
rect 791 3929 795 3930
rect 815 3934 819 3935
rect 815 3929 819 3930
rect 112 3902 114 3929
rect 304 3905 306 3929
rect 424 3905 426 3929
rect 552 3905 554 3929
rect 688 3905 690 3929
rect 816 3905 818 3929
rect 302 3904 308 3905
rect 110 3901 116 3902
rect 110 3897 111 3901
rect 115 3897 116 3901
rect 302 3900 303 3904
rect 307 3900 308 3904
rect 302 3899 308 3900
rect 422 3904 428 3905
rect 422 3900 423 3904
rect 427 3900 428 3904
rect 422 3899 428 3900
rect 550 3904 556 3905
rect 550 3900 551 3904
rect 555 3900 556 3904
rect 550 3899 556 3900
rect 686 3904 692 3905
rect 686 3900 687 3904
rect 691 3900 692 3904
rect 686 3899 692 3900
rect 814 3904 820 3905
rect 814 3900 815 3904
rect 819 3900 820 3904
rect 814 3899 820 3900
rect 110 3896 116 3897
rect 378 3895 384 3896
rect 378 3891 379 3895
rect 383 3891 384 3895
rect 378 3890 384 3891
rect 498 3895 504 3896
rect 498 3891 499 3895
rect 503 3891 504 3895
rect 498 3890 504 3891
rect 626 3895 632 3896
rect 626 3891 627 3895
rect 631 3891 632 3895
rect 626 3890 632 3891
rect 762 3895 768 3896
rect 762 3891 763 3895
rect 767 3891 768 3895
rect 762 3890 768 3891
rect 770 3895 776 3896
rect 770 3891 771 3895
rect 775 3891 776 3895
rect 770 3890 776 3891
rect 302 3885 308 3886
rect 110 3884 116 3885
rect 110 3880 111 3884
rect 115 3880 116 3884
rect 302 3881 303 3885
rect 307 3881 308 3885
rect 302 3880 308 3881
rect 110 3879 116 3880
rect 112 3855 114 3879
rect 304 3855 306 3880
rect 380 3868 382 3890
rect 422 3885 428 3886
rect 422 3881 423 3885
rect 427 3881 428 3885
rect 422 3880 428 3881
rect 378 3867 384 3868
rect 378 3863 379 3867
rect 383 3863 384 3867
rect 378 3862 384 3863
rect 424 3855 426 3880
rect 500 3868 502 3890
rect 550 3885 556 3886
rect 550 3881 551 3885
rect 555 3881 556 3885
rect 550 3880 556 3881
rect 498 3867 504 3868
rect 498 3863 499 3867
rect 503 3863 504 3867
rect 498 3862 504 3863
rect 552 3855 554 3880
rect 628 3868 630 3890
rect 686 3885 692 3886
rect 686 3881 687 3885
rect 691 3881 692 3885
rect 686 3880 692 3881
rect 626 3867 632 3868
rect 626 3863 627 3867
rect 631 3863 632 3867
rect 626 3862 632 3863
rect 688 3855 690 3880
rect 764 3868 766 3890
rect 762 3867 768 3868
rect 762 3863 763 3867
rect 767 3863 768 3867
rect 762 3862 768 3863
rect 772 3856 774 3890
rect 814 3885 820 3886
rect 814 3881 815 3885
rect 819 3881 820 3885
rect 814 3880 820 3881
rect 770 3855 776 3856
rect 816 3855 818 3880
rect 920 3876 922 3970
rect 974 3964 980 3965
rect 974 3960 975 3964
rect 979 3960 980 3964
rect 974 3959 980 3960
rect 1150 3964 1156 3965
rect 1150 3960 1151 3964
rect 1155 3960 1156 3964
rect 1150 3959 1156 3960
rect 1310 3964 1316 3965
rect 1310 3960 1311 3964
rect 1315 3960 1316 3964
rect 1310 3959 1316 3960
rect 976 3935 978 3959
rect 1152 3935 1154 3959
rect 1312 3935 1314 3959
rect 943 3934 947 3935
rect 943 3929 947 3930
rect 975 3934 979 3935
rect 975 3929 979 3930
rect 1071 3934 1075 3935
rect 1071 3929 1075 3930
rect 1151 3934 1155 3935
rect 1151 3929 1155 3930
rect 1199 3934 1203 3935
rect 1199 3929 1203 3930
rect 1311 3934 1315 3935
rect 1311 3929 1315 3930
rect 1327 3934 1331 3935
rect 1327 3929 1331 3930
rect 944 3905 946 3929
rect 1072 3905 1074 3929
rect 1200 3905 1202 3929
rect 1328 3905 1330 3929
rect 942 3904 948 3905
rect 942 3900 943 3904
rect 947 3900 948 3904
rect 942 3899 948 3900
rect 1070 3904 1076 3905
rect 1070 3900 1071 3904
rect 1075 3900 1076 3904
rect 1070 3899 1076 3900
rect 1198 3904 1204 3905
rect 1198 3900 1199 3904
rect 1203 3900 1204 3904
rect 1198 3899 1204 3900
rect 1326 3904 1332 3905
rect 1326 3900 1327 3904
rect 1331 3900 1332 3904
rect 1326 3899 1332 3900
rect 1412 3896 1414 3990
rect 1472 3984 1474 4005
rect 1546 4003 1552 4004
rect 1546 3999 1547 4003
rect 1551 3999 1552 4003
rect 1546 3998 1552 3999
rect 1470 3983 1476 3984
rect 1470 3979 1471 3983
rect 1475 3979 1476 3983
rect 1470 3978 1476 3979
rect 1548 3976 1550 3998
rect 1624 3984 1626 4005
rect 1698 4003 1704 4004
rect 1698 3999 1699 4003
rect 1703 3999 1704 4003
rect 1698 3998 1704 3999
rect 1622 3983 1628 3984
rect 1622 3979 1623 3983
rect 1627 3979 1628 3983
rect 1622 3978 1628 3979
rect 1700 3976 1702 3998
rect 1776 3984 1778 4005
rect 1850 4003 1856 4004
rect 1850 3999 1851 4003
rect 1855 3999 1856 4003
rect 1850 3998 1856 3999
rect 1774 3983 1780 3984
rect 1774 3979 1775 3983
rect 1779 3979 1780 3983
rect 1774 3978 1780 3979
rect 1852 3976 1854 3998
rect 1904 3984 1906 4005
rect 1902 3983 1908 3984
rect 1902 3979 1903 3983
rect 1907 3979 1908 3983
rect 1902 3978 1908 3979
rect 1980 3976 1982 4018
rect 2007 4010 2011 4011
rect 2007 4005 2011 4006
rect 2048 4005 2050 4025
rect 2008 3985 2010 4005
rect 2046 4004 2052 4005
rect 2072 4004 2074 4025
rect 3944 4005 3946 4025
rect 3942 4004 3948 4005
rect 2046 4000 2047 4004
rect 2051 4000 2052 4004
rect 2046 3999 2052 4000
rect 2070 4003 2076 4004
rect 2070 3999 2071 4003
rect 2075 3999 2076 4003
rect 3942 4000 3943 4004
rect 3947 4000 3948 4004
rect 3942 3999 3948 4000
rect 2070 3998 2076 3999
rect 2146 3991 2152 3992
rect 2046 3987 2052 3988
rect 2006 3984 2012 3985
rect 2006 3980 2007 3984
rect 2011 3980 2012 3984
rect 2046 3983 2047 3987
rect 2051 3983 2052 3987
rect 2146 3987 2147 3991
rect 2151 3987 2152 3991
rect 2146 3986 2152 3987
rect 3942 3987 3948 3988
rect 2046 3982 2052 3983
rect 2070 3984 2076 3985
rect 2006 3979 2012 3980
rect 1546 3975 1552 3976
rect 1546 3971 1547 3975
rect 1551 3971 1552 3975
rect 1546 3970 1552 3971
rect 1698 3975 1704 3976
rect 1698 3971 1699 3975
rect 1703 3971 1704 3975
rect 1698 3970 1704 3971
rect 1850 3975 1856 3976
rect 1850 3971 1851 3975
rect 1855 3971 1856 3975
rect 1850 3970 1856 3971
rect 1978 3975 1984 3976
rect 1978 3971 1979 3975
rect 1983 3971 1984 3975
rect 1978 3970 1984 3971
rect 2006 3967 2012 3968
rect 1470 3964 1476 3965
rect 1470 3960 1471 3964
rect 1475 3960 1476 3964
rect 1470 3959 1476 3960
rect 1622 3964 1628 3965
rect 1622 3960 1623 3964
rect 1627 3960 1628 3964
rect 1622 3959 1628 3960
rect 1774 3964 1780 3965
rect 1774 3960 1775 3964
rect 1779 3960 1780 3964
rect 1774 3959 1780 3960
rect 1902 3964 1908 3965
rect 1902 3960 1903 3964
rect 1907 3960 1908 3964
rect 2006 3963 2007 3967
rect 2011 3963 2012 3967
rect 2006 3962 2012 3963
rect 1902 3959 1908 3960
rect 1472 3935 1474 3959
rect 1624 3935 1626 3959
rect 1776 3935 1778 3959
rect 1904 3935 1906 3959
rect 2008 3935 2010 3962
rect 2048 3955 2050 3982
rect 2070 3980 2071 3984
rect 2075 3980 2076 3984
rect 2070 3979 2076 3980
rect 2072 3955 2074 3979
rect 2047 3954 2051 3955
rect 2047 3949 2051 3950
rect 2071 3954 2075 3955
rect 2071 3949 2075 3950
rect 2079 3954 2083 3955
rect 2079 3949 2083 3950
rect 1463 3934 1467 3935
rect 1463 3929 1467 3930
rect 1471 3934 1475 3935
rect 1471 3929 1475 3930
rect 1623 3934 1627 3935
rect 1623 3929 1627 3930
rect 1775 3934 1779 3935
rect 1775 3929 1779 3930
rect 1903 3934 1907 3935
rect 1903 3929 1907 3930
rect 2007 3934 2011 3935
rect 2007 3929 2011 3930
rect 1464 3905 1466 3929
rect 1462 3904 1468 3905
rect 1462 3900 1463 3904
rect 1467 3900 1468 3904
rect 2008 3902 2010 3929
rect 2048 3922 2050 3949
rect 2080 3925 2082 3949
rect 2078 3924 2084 3925
rect 2046 3921 2052 3922
rect 2046 3917 2047 3921
rect 2051 3917 2052 3921
rect 2078 3920 2079 3924
rect 2083 3920 2084 3924
rect 2078 3919 2084 3920
rect 2046 3916 2052 3917
rect 2078 3905 2084 3906
rect 2046 3904 2052 3905
rect 1462 3899 1468 3900
rect 2006 3901 2012 3902
rect 2006 3897 2007 3901
rect 2011 3897 2012 3901
rect 2046 3900 2047 3904
rect 2051 3900 2052 3904
rect 2078 3901 2079 3905
rect 2083 3901 2084 3905
rect 2078 3900 2084 3901
rect 2046 3899 2052 3900
rect 2006 3896 2012 3897
rect 1018 3895 1024 3896
rect 1018 3891 1019 3895
rect 1023 3891 1024 3895
rect 1018 3890 1024 3891
rect 1146 3895 1152 3896
rect 1146 3891 1147 3895
rect 1151 3891 1152 3895
rect 1146 3890 1152 3891
rect 1274 3895 1280 3896
rect 1274 3891 1275 3895
rect 1279 3891 1280 3895
rect 1274 3890 1280 3891
rect 1402 3895 1408 3896
rect 1402 3891 1403 3895
rect 1407 3891 1408 3895
rect 1402 3890 1408 3891
rect 1410 3895 1416 3896
rect 1410 3891 1411 3895
rect 1415 3891 1416 3895
rect 1410 3890 1416 3891
rect 942 3885 948 3886
rect 942 3881 943 3885
rect 947 3881 948 3885
rect 942 3880 948 3881
rect 918 3875 924 3876
rect 918 3871 919 3875
rect 923 3871 924 3875
rect 918 3870 924 3871
rect 944 3855 946 3880
rect 1020 3868 1022 3890
rect 1070 3885 1076 3886
rect 1070 3881 1071 3885
rect 1075 3881 1076 3885
rect 1070 3880 1076 3881
rect 1018 3867 1024 3868
rect 982 3863 988 3864
rect 982 3859 983 3863
rect 987 3859 988 3863
rect 1018 3863 1019 3867
rect 1023 3863 1024 3867
rect 1018 3862 1024 3863
rect 982 3858 988 3859
rect 111 3854 115 3855
rect 111 3849 115 3850
rect 303 3854 307 3855
rect 303 3849 307 3850
rect 415 3854 419 3855
rect 415 3849 419 3850
rect 423 3854 427 3855
rect 423 3849 427 3850
rect 551 3854 555 3855
rect 551 3849 555 3850
rect 567 3854 571 3855
rect 567 3849 571 3850
rect 687 3854 691 3855
rect 687 3849 691 3850
rect 727 3854 731 3855
rect 770 3851 771 3855
rect 775 3851 776 3855
rect 770 3850 776 3851
rect 815 3854 819 3855
rect 727 3849 731 3850
rect 815 3849 819 3850
rect 887 3854 891 3855
rect 887 3849 891 3850
rect 943 3854 947 3855
rect 943 3849 947 3850
rect 112 3829 114 3849
rect 110 3828 116 3829
rect 416 3828 418 3849
rect 490 3847 496 3848
rect 490 3843 491 3847
rect 495 3843 496 3847
rect 490 3842 496 3843
rect 110 3824 111 3828
rect 115 3824 116 3828
rect 110 3823 116 3824
rect 414 3827 420 3828
rect 414 3823 415 3827
rect 419 3823 420 3827
rect 414 3822 420 3823
rect 492 3820 494 3842
rect 568 3828 570 3849
rect 642 3847 648 3848
rect 642 3843 643 3847
rect 647 3843 648 3847
rect 642 3842 648 3843
rect 566 3827 572 3828
rect 566 3823 567 3827
rect 571 3823 572 3827
rect 566 3822 572 3823
rect 644 3820 646 3842
rect 728 3828 730 3849
rect 802 3847 808 3848
rect 802 3843 803 3847
rect 807 3843 808 3847
rect 802 3842 808 3843
rect 726 3827 732 3828
rect 726 3823 727 3827
rect 731 3823 732 3827
rect 726 3822 732 3823
rect 804 3820 806 3842
rect 888 3828 890 3849
rect 886 3827 892 3828
rect 886 3823 887 3827
rect 891 3823 892 3827
rect 886 3822 892 3823
rect 984 3820 986 3858
rect 1072 3855 1074 3880
rect 1148 3868 1150 3890
rect 1198 3885 1204 3886
rect 1198 3881 1199 3885
rect 1203 3881 1204 3885
rect 1198 3880 1204 3881
rect 1146 3867 1152 3868
rect 1146 3863 1147 3867
rect 1151 3863 1152 3867
rect 1146 3862 1152 3863
rect 1200 3855 1202 3880
rect 1276 3868 1278 3890
rect 1326 3885 1332 3886
rect 1326 3881 1327 3885
rect 1331 3881 1332 3885
rect 1326 3880 1332 3881
rect 1274 3867 1280 3868
rect 1274 3863 1275 3867
rect 1279 3863 1280 3867
rect 1274 3862 1280 3863
rect 1328 3855 1330 3880
rect 1404 3868 1406 3890
rect 1462 3885 1468 3886
rect 1462 3881 1463 3885
rect 1467 3881 1468 3885
rect 1462 3880 1468 3881
rect 2006 3884 2012 3885
rect 2006 3880 2007 3884
rect 2011 3880 2012 3884
rect 1402 3867 1408 3868
rect 1402 3863 1403 3867
rect 1407 3863 1408 3867
rect 1402 3862 1408 3863
rect 1464 3855 1466 3880
rect 2006 3879 2012 3880
rect 2048 3879 2050 3899
rect 2080 3879 2082 3900
rect 2148 3888 2150 3986
rect 3942 3983 3943 3987
rect 3947 3983 3948 3987
rect 3942 3982 3948 3983
rect 3944 3955 3946 3982
rect 2215 3954 2219 3955
rect 2215 3949 2219 3950
rect 2359 3954 2363 3955
rect 2359 3949 2363 3950
rect 2503 3954 2507 3955
rect 2503 3949 2507 3950
rect 2647 3954 2651 3955
rect 2647 3949 2651 3950
rect 2791 3954 2795 3955
rect 2791 3949 2795 3950
rect 2927 3954 2931 3955
rect 2927 3949 2931 3950
rect 3055 3954 3059 3955
rect 3055 3949 3059 3950
rect 3175 3954 3179 3955
rect 3175 3949 3179 3950
rect 3295 3954 3299 3955
rect 3295 3949 3299 3950
rect 3415 3954 3419 3955
rect 3415 3949 3419 3950
rect 3535 3954 3539 3955
rect 3535 3949 3539 3950
rect 3943 3954 3947 3955
rect 3943 3949 3947 3950
rect 2216 3925 2218 3949
rect 2360 3925 2362 3949
rect 2504 3925 2506 3949
rect 2648 3925 2650 3949
rect 2792 3925 2794 3949
rect 2928 3925 2930 3949
rect 3056 3925 3058 3949
rect 3176 3925 3178 3949
rect 3296 3925 3298 3949
rect 3416 3925 3418 3949
rect 3536 3925 3538 3949
rect 2214 3924 2220 3925
rect 2214 3920 2215 3924
rect 2219 3920 2220 3924
rect 2214 3919 2220 3920
rect 2358 3924 2364 3925
rect 2358 3920 2359 3924
rect 2363 3920 2364 3924
rect 2358 3919 2364 3920
rect 2502 3924 2508 3925
rect 2502 3920 2503 3924
rect 2507 3920 2508 3924
rect 2502 3919 2508 3920
rect 2646 3924 2652 3925
rect 2646 3920 2647 3924
rect 2651 3920 2652 3924
rect 2646 3919 2652 3920
rect 2790 3924 2796 3925
rect 2790 3920 2791 3924
rect 2795 3920 2796 3924
rect 2790 3919 2796 3920
rect 2926 3924 2932 3925
rect 2926 3920 2927 3924
rect 2931 3920 2932 3924
rect 2926 3919 2932 3920
rect 3054 3924 3060 3925
rect 3054 3920 3055 3924
rect 3059 3920 3060 3924
rect 3054 3919 3060 3920
rect 3174 3924 3180 3925
rect 3174 3920 3175 3924
rect 3179 3920 3180 3924
rect 3174 3919 3180 3920
rect 3294 3924 3300 3925
rect 3294 3920 3295 3924
rect 3299 3920 3300 3924
rect 3294 3919 3300 3920
rect 3414 3924 3420 3925
rect 3414 3920 3415 3924
rect 3419 3920 3420 3924
rect 3414 3919 3420 3920
rect 3534 3924 3540 3925
rect 3534 3920 3535 3924
rect 3539 3920 3540 3924
rect 3944 3922 3946 3949
rect 3534 3919 3540 3920
rect 3942 3921 3948 3922
rect 3942 3917 3943 3921
rect 3947 3917 3948 3921
rect 3942 3916 3948 3917
rect 2154 3915 2160 3916
rect 2154 3911 2155 3915
rect 2159 3911 2160 3915
rect 2154 3910 2160 3911
rect 2290 3915 2296 3916
rect 2290 3911 2291 3915
rect 2295 3911 2296 3915
rect 2290 3910 2296 3911
rect 2434 3915 2440 3916
rect 2434 3911 2435 3915
rect 2439 3911 2440 3915
rect 2434 3910 2440 3911
rect 2578 3915 2584 3916
rect 2578 3911 2579 3915
rect 2583 3911 2584 3915
rect 2578 3910 2584 3911
rect 2714 3915 2720 3916
rect 2714 3911 2715 3915
rect 2719 3911 2720 3915
rect 2714 3910 2720 3911
rect 2866 3915 2872 3916
rect 2866 3911 2867 3915
rect 2871 3911 2872 3915
rect 2866 3910 2872 3911
rect 3002 3915 3008 3916
rect 3002 3911 3003 3915
rect 3007 3911 3008 3915
rect 3002 3910 3008 3911
rect 3130 3915 3136 3916
rect 3130 3911 3131 3915
rect 3135 3911 3136 3915
rect 3130 3910 3136 3911
rect 3250 3915 3256 3916
rect 3250 3911 3251 3915
rect 3255 3911 3256 3915
rect 3250 3910 3256 3911
rect 3370 3915 3376 3916
rect 3370 3911 3371 3915
rect 3375 3911 3376 3915
rect 3370 3910 3376 3911
rect 3490 3915 3496 3916
rect 3490 3911 3491 3915
rect 3495 3911 3496 3915
rect 3490 3910 3496 3911
rect 3610 3915 3616 3916
rect 3610 3911 3611 3915
rect 3615 3911 3616 3915
rect 3610 3910 3616 3911
rect 2156 3888 2158 3910
rect 2214 3905 2220 3906
rect 2214 3901 2215 3905
rect 2219 3901 2220 3905
rect 2214 3900 2220 3901
rect 2146 3887 2152 3888
rect 2146 3883 2147 3887
rect 2151 3883 2152 3887
rect 2146 3882 2152 3883
rect 2154 3887 2160 3888
rect 2154 3883 2155 3887
rect 2159 3883 2160 3887
rect 2154 3882 2160 3883
rect 2216 3879 2218 3900
rect 2292 3888 2294 3910
rect 2358 3905 2364 3906
rect 2358 3901 2359 3905
rect 2363 3901 2364 3905
rect 2358 3900 2364 3901
rect 2290 3887 2296 3888
rect 2290 3883 2291 3887
rect 2295 3883 2296 3887
rect 2290 3882 2296 3883
rect 2360 3879 2362 3900
rect 2436 3888 2438 3910
rect 2502 3905 2508 3906
rect 2502 3901 2503 3905
rect 2507 3901 2508 3905
rect 2502 3900 2508 3901
rect 2434 3887 2440 3888
rect 2434 3883 2435 3887
rect 2439 3883 2440 3887
rect 2434 3882 2440 3883
rect 2504 3879 2506 3900
rect 2580 3888 2582 3910
rect 2646 3905 2652 3906
rect 2646 3901 2647 3905
rect 2651 3901 2652 3905
rect 2646 3900 2652 3901
rect 2578 3887 2584 3888
rect 2578 3883 2579 3887
rect 2583 3883 2584 3887
rect 2578 3882 2584 3883
rect 2648 3879 2650 3900
rect 2008 3855 2010 3879
rect 2047 3878 2051 3879
rect 2047 3873 2051 3874
rect 2079 3878 2083 3879
rect 2079 3873 2083 3874
rect 2215 3878 2219 3879
rect 2215 3873 2219 3874
rect 2255 3878 2259 3879
rect 2255 3873 2259 3874
rect 2359 3878 2363 3879
rect 2359 3873 2363 3874
rect 2383 3878 2387 3879
rect 2383 3873 2387 3874
rect 2503 3878 2507 3879
rect 2503 3873 2507 3874
rect 2519 3878 2523 3879
rect 2519 3873 2523 3874
rect 2647 3878 2651 3879
rect 2647 3873 2651 3874
rect 2671 3878 2675 3879
rect 2671 3873 2675 3874
rect 1039 3854 1043 3855
rect 1039 3849 1043 3850
rect 1071 3854 1075 3855
rect 1071 3849 1075 3850
rect 1191 3854 1195 3855
rect 1191 3849 1195 3850
rect 1199 3854 1203 3855
rect 1199 3849 1203 3850
rect 1327 3854 1331 3855
rect 1327 3849 1331 3850
rect 1343 3854 1347 3855
rect 1343 3849 1347 3850
rect 1463 3854 1467 3855
rect 1463 3849 1467 3850
rect 1495 3854 1499 3855
rect 1495 3849 1499 3850
rect 1647 3854 1651 3855
rect 1647 3849 1651 3850
rect 2007 3854 2011 3855
rect 2048 3853 2050 3873
rect 2007 3849 2011 3850
rect 2046 3852 2052 3853
rect 2256 3852 2258 3873
rect 2330 3871 2336 3872
rect 2330 3867 2331 3871
rect 2335 3867 2336 3871
rect 2330 3866 2336 3867
rect 1040 3828 1042 3849
rect 1138 3847 1144 3848
rect 1138 3843 1139 3847
rect 1143 3843 1144 3847
rect 1138 3842 1144 3843
rect 1038 3827 1044 3828
rect 1038 3823 1039 3827
rect 1043 3823 1044 3827
rect 1038 3822 1044 3823
rect 1140 3820 1142 3842
rect 1192 3828 1194 3849
rect 1274 3847 1280 3848
rect 1274 3843 1275 3847
rect 1279 3843 1280 3847
rect 1274 3842 1280 3843
rect 1190 3827 1196 3828
rect 1190 3823 1191 3827
rect 1195 3823 1196 3827
rect 1190 3822 1196 3823
rect 1276 3820 1278 3842
rect 1344 3828 1346 3849
rect 1426 3847 1432 3848
rect 1426 3843 1427 3847
rect 1431 3843 1432 3847
rect 1426 3842 1432 3843
rect 1342 3827 1348 3828
rect 1342 3823 1343 3827
rect 1347 3823 1348 3827
rect 1342 3822 1348 3823
rect 1428 3820 1430 3842
rect 1496 3828 1498 3849
rect 1562 3847 1568 3848
rect 1562 3843 1563 3847
rect 1567 3843 1568 3847
rect 1562 3842 1568 3843
rect 1578 3847 1584 3848
rect 1578 3843 1579 3847
rect 1583 3843 1584 3847
rect 1578 3842 1584 3843
rect 1494 3827 1500 3828
rect 1494 3823 1495 3827
rect 1499 3823 1500 3827
rect 1564 3824 1566 3842
rect 1494 3822 1500 3823
rect 1562 3823 1568 3824
rect 490 3819 496 3820
rect 490 3815 491 3819
rect 495 3815 496 3819
rect 490 3814 496 3815
rect 642 3819 648 3820
rect 642 3815 643 3819
rect 647 3815 648 3819
rect 642 3814 648 3815
rect 802 3819 808 3820
rect 802 3815 803 3819
rect 807 3815 808 3819
rect 802 3814 808 3815
rect 858 3819 864 3820
rect 858 3815 859 3819
rect 863 3815 864 3819
rect 858 3814 864 3815
rect 982 3819 988 3820
rect 982 3815 983 3819
rect 987 3815 988 3819
rect 982 3814 988 3815
rect 1138 3819 1144 3820
rect 1138 3815 1139 3819
rect 1143 3815 1144 3819
rect 1138 3814 1144 3815
rect 1274 3819 1280 3820
rect 1274 3815 1275 3819
rect 1279 3815 1280 3819
rect 1274 3814 1280 3815
rect 1426 3819 1432 3820
rect 1426 3815 1427 3819
rect 1431 3815 1432 3819
rect 1562 3819 1563 3823
rect 1567 3819 1568 3823
rect 1562 3818 1568 3819
rect 1426 3814 1432 3815
rect 110 3811 116 3812
rect 110 3807 111 3811
rect 115 3807 116 3811
rect 110 3806 116 3807
rect 414 3808 420 3809
rect 112 3775 114 3806
rect 414 3804 415 3808
rect 419 3804 420 3808
rect 414 3803 420 3804
rect 566 3808 572 3809
rect 566 3804 567 3808
rect 571 3804 572 3808
rect 566 3803 572 3804
rect 726 3808 732 3809
rect 726 3804 727 3808
rect 731 3804 732 3808
rect 726 3803 732 3804
rect 416 3775 418 3803
rect 568 3775 570 3803
rect 728 3775 730 3803
rect 111 3774 115 3775
rect 111 3769 115 3770
rect 399 3774 403 3775
rect 399 3769 403 3770
rect 415 3774 419 3775
rect 415 3769 419 3770
rect 567 3774 571 3775
rect 567 3769 571 3770
rect 727 3774 731 3775
rect 727 3769 731 3770
rect 751 3774 755 3775
rect 751 3769 755 3770
rect 112 3742 114 3769
rect 400 3745 402 3769
rect 438 3755 444 3756
rect 438 3751 439 3755
rect 443 3751 444 3755
rect 438 3750 444 3751
rect 398 3744 404 3745
rect 110 3741 116 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 398 3740 399 3744
rect 403 3740 404 3744
rect 398 3739 404 3740
rect 110 3736 116 3737
rect 398 3725 404 3726
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 398 3721 399 3725
rect 403 3721 404 3725
rect 398 3720 404 3721
rect 110 3719 116 3720
rect 112 3687 114 3719
rect 400 3687 402 3720
rect 440 3708 442 3750
rect 568 3745 570 3769
rect 752 3745 754 3769
rect 860 3756 862 3814
rect 886 3808 892 3809
rect 886 3804 887 3808
rect 891 3804 892 3808
rect 886 3803 892 3804
rect 1038 3808 1044 3809
rect 1038 3804 1039 3808
rect 1043 3804 1044 3808
rect 1038 3803 1044 3804
rect 1190 3808 1196 3809
rect 1190 3804 1191 3808
rect 1195 3804 1196 3808
rect 1190 3803 1196 3804
rect 1342 3808 1348 3809
rect 1342 3804 1343 3808
rect 1347 3804 1348 3808
rect 1342 3803 1348 3804
rect 1494 3808 1500 3809
rect 1494 3804 1495 3808
rect 1499 3804 1500 3808
rect 1494 3803 1500 3804
rect 888 3775 890 3803
rect 1040 3775 1042 3803
rect 1192 3775 1194 3803
rect 1344 3775 1346 3803
rect 1496 3775 1498 3803
rect 887 3774 891 3775
rect 887 3769 891 3770
rect 935 3774 939 3775
rect 935 3769 939 3770
rect 1039 3774 1043 3775
rect 1039 3769 1043 3770
rect 1127 3774 1131 3775
rect 1127 3769 1131 3770
rect 1191 3774 1195 3775
rect 1191 3769 1195 3770
rect 1311 3774 1315 3775
rect 1311 3769 1315 3770
rect 1343 3774 1347 3775
rect 1343 3769 1347 3770
rect 1495 3774 1499 3775
rect 1495 3769 1499 3770
rect 1503 3774 1507 3775
rect 1503 3769 1507 3770
rect 858 3755 864 3756
rect 858 3751 859 3755
rect 863 3751 864 3755
rect 858 3750 864 3751
rect 936 3745 938 3769
rect 1128 3745 1130 3769
rect 1312 3745 1314 3769
rect 1504 3745 1506 3769
rect 566 3744 572 3745
rect 566 3740 567 3744
rect 571 3740 572 3744
rect 566 3739 572 3740
rect 750 3744 756 3745
rect 750 3740 751 3744
rect 755 3740 756 3744
rect 750 3739 756 3740
rect 934 3744 940 3745
rect 934 3740 935 3744
rect 939 3740 940 3744
rect 934 3739 940 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1310 3744 1316 3745
rect 1310 3740 1311 3744
rect 1315 3740 1316 3744
rect 1310 3739 1316 3740
rect 1502 3744 1508 3745
rect 1502 3740 1503 3744
rect 1507 3740 1508 3744
rect 1502 3739 1508 3740
rect 1580 3736 1582 3842
rect 1648 3828 1650 3849
rect 2008 3829 2010 3849
rect 2046 3848 2047 3852
rect 2051 3848 2052 3852
rect 2046 3847 2052 3848
rect 2254 3851 2260 3852
rect 2254 3847 2255 3851
rect 2259 3847 2260 3851
rect 2254 3846 2260 3847
rect 2332 3844 2334 3866
rect 2384 3852 2386 3873
rect 2458 3871 2464 3872
rect 2458 3867 2459 3871
rect 2463 3867 2464 3871
rect 2458 3866 2464 3867
rect 2382 3851 2388 3852
rect 2382 3847 2383 3851
rect 2387 3847 2388 3851
rect 2382 3846 2388 3847
rect 2460 3844 2462 3866
rect 2520 3852 2522 3873
rect 2672 3852 2674 3873
rect 2716 3872 2718 3910
rect 2790 3905 2796 3906
rect 2790 3901 2791 3905
rect 2795 3901 2796 3905
rect 2790 3900 2796 3901
rect 2792 3879 2794 3900
rect 2868 3888 2870 3910
rect 2926 3905 2932 3906
rect 2926 3901 2927 3905
rect 2931 3901 2932 3905
rect 2926 3900 2932 3901
rect 2866 3887 2872 3888
rect 2866 3883 2867 3887
rect 2871 3883 2872 3887
rect 2866 3882 2872 3883
rect 2928 3879 2930 3900
rect 3004 3888 3006 3910
rect 3054 3905 3060 3906
rect 3054 3901 3055 3905
rect 3059 3901 3060 3905
rect 3054 3900 3060 3901
rect 3002 3887 3008 3888
rect 3002 3883 3003 3887
rect 3007 3883 3008 3887
rect 3002 3882 3008 3883
rect 3056 3879 3058 3900
rect 3132 3888 3134 3910
rect 3174 3905 3180 3906
rect 3174 3901 3175 3905
rect 3179 3901 3180 3905
rect 3174 3900 3180 3901
rect 3130 3887 3136 3888
rect 3130 3883 3131 3887
rect 3135 3883 3136 3887
rect 3130 3882 3136 3883
rect 3078 3879 3084 3880
rect 3176 3879 3178 3900
rect 3252 3888 3254 3910
rect 3294 3905 3300 3906
rect 3294 3901 3295 3905
rect 3299 3901 3300 3905
rect 3294 3900 3300 3901
rect 3250 3887 3256 3888
rect 3250 3883 3251 3887
rect 3255 3883 3256 3887
rect 3250 3882 3256 3883
rect 3296 3879 3298 3900
rect 3372 3888 3374 3910
rect 3414 3905 3420 3906
rect 3414 3901 3415 3905
rect 3419 3901 3420 3905
rect 3414 3900 3420 3901
rect 3370 3887 3376 3888
rect 3370 3883 3371 3887
rect 3375 3883 3376 3887
rect 3370 3882 3376 3883
rect 3416 3879 3418 3900
rect 3492 3888 3494 3910
rect 3534 3905 3540 3906
rect 3534 3901 3535 3905
rect 3539 3901 3540 3905
rect 3534 3900 3540 3901
rect 3490 3887 3496 3888
rect 3490 3883 3491 3887
rect 3495 3883 3496 3887
rect 3490 3882 3496 3883
rect 3536 3879 3538 3900
rect 2791 3878 2795 3879
rect 2791 3873 2795 3874
rect 2831 3878 2835 3879
rect 2831 3873 2835 3874
rect 2927 3878 2931 3879
rect 2927 3873 2931 3874
rect 2991 3878 2995 3879
rect 2991 3873 2995 3874
rect 3055 3878 3059 3879
rect 3078 3875 3079 3879
rect 3083 3875 3084 3879
rect 3078 3874 3084 3875
rect 3159 3878 3163 3879
rect 3055 3873 3059 3874
rect 2710 3871 2718 3872
rect 2710 3867 2711 3871
rect 2715 3868 2718 3871
rect 2746 3871 2752 3872
rect 2715 3867 2716 3868
rect 2710 3866 2716 3867
rect 2746 3867 2747 3871
rect 2751 3867 2752 3871
rect 2746 3866 2752 3867
rect 2518 3851 2524 3852
rect 2518 3847 2519 3851
rect 2523 3847 2524 3851
rect 2518 3846 2524 3847
rect 2670 3851 2676 3852
rect 2670 3847 2671 3851
rect 2675 3847 2676 3851
rect 2670 3846 2676 3847
rect 2748 3844 2750 3866
rect 2778 3863 2784 3864
rect 2778 3859 2779 3863
rect 2783 3859 2784 3863
rect 2778 3858 2784 3859
rect 2780 3844 2782 3858
rect 2832 3852 2834 3873
rect 2992 3852 2994 3873
rect 3026 3871 3032 3872
rect 3026 3867 3027 3871
rect 3031 3867 3032 3871
rect 3026 3866 3032 3867
rect 3066 3871 3072 3872
rect 3066 3867 3067 3871
rect 3071 3867 3072 3871
rect 3066 3866 3072 3867
rect 2830 3851 2836 3852
rect 2830 3847 2831 3851
rect 2835 3847 2836 3851
rect 2830 3846 2836 3847
rect 2990 3851 2996 3852
rect 2990 3847 2991 3851
rect 2995 3847 2996 3851
rect 2990 3846 2996 3847
rect 2330 3843 2336 3844
rect 2330 3839 2331 3843
rect 2335 3839 2336 3843
rect 2330 3838 2336 3839
rect 2458 3843 2464 3844
rect 2458 3839 2459 3843
rect 2463 3839 2464 3843
rect 2746 3843 2752 3844
rect 2458 3838 2464 3839
rect 2594 3839 2600 3840
rect 2046 3835 2052 3836
rect 2046 3831 2047 3835
rect 2051 3831 2052 3835
rect 2594 3835 2595 3839
rect 2599 3835 2600 3839
rect 2746 3839 2747 3843
rect 2751 3839 2752 3843
rect 2746 3838 2752 3839
rect 2778 3843 2784 3844
rect 2778 3839 2779 3843
rect 2783 3839 2784 3843
rect 2778 3838 2784 3839
rect 2594 3834 2600 3835
rect 2046 3830 2052 3831
rect 2254 3832 2260 3833
rect 2006 3828 2012 3829
rect 1646 3827 1652 3828
rect 1646 3823 1647 3827
rect 1651 3823 1652 3827
rect 2006 3824 2007 3828
rect 2011 3824 2012 3828
rect 2006 3823 2012 3824
rect 1646 3822 1652 3823
rect 2006 3811 2012 3812
rect 1646 3808 1652 3809
rect 1646 3804 1647 3808
rect 1651 3804 1652 3808
rect 2006 3807 2007 3811
rect 2011 3807 2012 3811
rect 2006 3806 2012 3807
rect 1646 3803 1652 3804
rect 1648 3775 1650 3803
rect 2008 3775 2010 3806
rect 2048 3803 2050 3830
rect 2254 3828 2255 3832
rect 2259 3828 2260 3832
rect 2254 3827 2260 3828
rect 2382 3832 2388 3833
rect 2382 3828 2383 3832
rect 2387 3828 2388 3832
rect 2382 3827 2388 3828
rect 2518 3832 2524 3833
rect 2518 3828 2519 3832
rect 2523 3828 2524 3832
rect 2518 3827 2524 3828
rect 2256 3803 2258 3827
rect 2384 3803 2386 3827
rect 2520 3803 2522 3827
rect 2047 3802 2051 3803
rect 2047 3797 2051 3798
rect 2071 3802 2075 3803
rect 2071 3797 2075 3798
rect 2199 3802 2203 3803
rect 2199 3797 2203 3798
rect 2255 3802 2259 3803
rect 2255 3797 2259 3798
rect 2375 3802 2379 3803
rect 2375 3797 2379 3798
rect 2383 3802 2387 3803
rect 2383 3797 2387 3798
rect 2519 3802 2523 3803
rect 2519 3797 2523 3798
rect 2559 3802 2563 3803
rect 2559 3797 2563 3798
rect 1647 3774 1651 3775
rect 1647 3769 1651 3770
rect 1695 3774 1699 3775
rect 1695 3769 1699 3770
rect 1887 3774 1891 3775
rect 1887 3769 1891 3770
rect 2007 3774 2011 3775
rect 2048 3770 2050 3797
rect 2072 3773 2074 3797
rect 2200 3773 2202 3797
rect 2376 3773 2378 3797
rect 2560 3773 2562 3797
rect 2070 3772 2076 3773
rect 2007 3769 2011 3770
rect 2046 3769 2052 3770
rect 1696 3745 1698 3769
rect 1888 3745 1890 3769
rect 1694 3744 1700 3745
rect 1694 3740 1695 3744
rect 1699 3740 1700 3744
rect 1694 3739 1700 3740
rect 1886 3744 1892 3745
rect 1886 3740 1887 3744
rect 1891 3740 1892 3744
rect 2008 3742 2010 3769
rect 2046 3765 2047 3769
rect 2051 3765 2052 3769
rect 2070 3768 2071 3772
rect 2075 3768 2076 3772
rect 2070 3767 2076 3768
rect 2198 3772 2204 3773
rect 2198 3768 2199 3772
rect 2203 3768 2204 3772
rect 2198 3767 2204 3768
rect 2374 3772 2380 3773
rect 2374 3768 2375 3772
rect 2379 3768 2380 3772
rect 2374 3767 2380 3768
rect 2558 3772 2564 3773
rect 2558 3768 2559 3772
rect 2563 3768 2564 3772
rect 2558 3767 2564 3768
rect 2046 3764 2052 3765
rect 2138 3763 2144 3764
rect 2138 3759 2139 3763
rect 2143 3759 2144 3763
rect 2138 3758 2144 3759
rect 2302 3763 2308 3764
rect 2302 3759 2303 3763
rect 2307 3759 2308 3763
rect 2302 3758 2308 3759
rect 2070 3753 2076 3754
rect 2046 3752 2052 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2070 3749 2071 3753
rect 2075 3749 2076 3753
rect 2070 3748 2076 3749
rect 2046 3747 2052 3748
rect 1886 3739 1892 3740
rect 2006 3741 2012 3742
rect 2006 3737 2007 3741
rect 2011 3737 2012 3741
rect 2006 3736 2012 3737
rect 474 3735 480 3736
rect 474 3731 475 3735
rect 479 3731 480 3735
rect 474 3730 480 3731
rect 642 3735 648 3736
rect 642 3731 643 3735
rect 647 3731 648 3735
rect 642 3730 648 3731
rect 826 3735 832 3736
rect 826 3731 827 3735
rect 831 3731 832 3735
rect 826 3730 832 3731
rect 1010 3735 1016 3736
rect 1010 3731 1011 3735
rect 1015 3731 1016 3735
rect 1010 3730 1016 3731
rect 1386 3735 1392 3736
rect 1386 3731 1387 3735
rect 1391 3731 1392 3735
rect 1386 3730 1392 3731
rect 1578 3735 1584 3736
rect 1578 3731 1579 3735
rect 1583 3731 1584 3735
rect 1578 3730 1584 3731
rect 1586 3735 1592 3736
rect 1586 3731 1587 3735
rect 1591 3731 1592 3735
rect 1586 3730 1592 3731
rect 1798 3735 1804 3736
rect 1798 3731 1799 3735
rect 1803 3731 1804 3735
rect 1798 3730 1804 3731
rect 476 3708 478 3730
rect 566 3725 572 3726
rect 566 3721 567 3725
rect 571 3721 572 3725
rect 566 3720 572 3721
rect 438 3707 444 3708
rect 438 3703 439 3707
rect 443 3703 444 3707
rect 438 3702 444 3703
rect 474 3707 480 3708
rect 474 3703 475 3707
rect 479 3703 480 3707
rect 474 3702 480 3703
rect 568 3687 570 3720
rect 644 3708 646 3730
rect 750 3725 756 3726
rect 750 3721 751 3725
rect 755 3721 756 3725
rect 750 3720 756 3721
rect 642 3707 648 3708
rect 642 3703 643 3707
rect 647 3703 648 3707
rect 642 3702 648 3703
rect 618 3687 624 3688
rect 752 3687 754 3720
rect 828 3708 830 3730
rect 934 3725 940 3726
rect 934 3721 935 3725
rect 939 3721 940 3725
rect 934 3720 940 3721
rect 826 3707 832 3708
rect 826 3703 827 3707
rect 831 3703 832 3707
rect 826 3702 832 3703
rect 936 3687 938 3720
rect 1012 3708 1014 3730
rect 1126 3725 1132 3726
rect 1126 3721 1127 3725
rect 1131 3721 1132 3725
rect 1126 3720 1132 3721
rect 1310 3725 1316 3726
rect 1310 3721 1311 3725
rect 1315 3721 1316 3725
rect 1310 3720 1316 3721
rect 1010 3707 1016 3708
rect 1010 3703 1011 3707
rect 1015 3703 1016 3707
rect 1010 3702 1016 3703
rect 1128 3687 1130 3720
rect 1312 3687 1314 3720
rect 1388 3708 1390 3730
rect 1502 3725 1508 3726
rect 1502 3721 1503 3725
rect 1507 3721 1508 3725
rect 1502 3720 1508 3721
rect 1386 3707 1392 3708
rect 1386 3703 1387 3707
rect 1391 3703 1392 3707
rect 1386 3702 1392 3703
rect 1458 3687 1464 3688
rect 1504 3687 1506 3720
rect 1588 3716 1590 3730
rect 1694 3725 1700 3726
rect 1694 3721 1695 3725
rect 1699 3721 1700 3725
rect 1694 3720 1700 3721
rect 1586 3715 1592 3716
rect 1586 3711 1587 3715
rect 1591 3711 1592 3715
rect 1586 3710 1592 3711
rect 1696 3687 1698 3720
rect 1800 3708 1802 3730
rect 1886 3725 1892 3726
rect 1886 3721 1887 3725
rect 1891 3721 1892 3725
rect 1886 3720 1892 3721
rect 2006 3724 2012 3725
rect 2006 3720 2007 3724
rect 2011 3720 2012 3724
rect 1798 3707 1804 3708
rect 1798 3703 1799 3707
rect 1803 3703 1804 3707
rect 1798 3702 1804 3703
rect 1866 3703 1872 3704
rect 1866 3699 1867 3703
rect 1871 3699 1872 3703
rect 1866 3698 1872 3699
rect 111 3686 115 3687
rect 111 3681 115 3682
rect 367 3686 371 3687
rect 367 3681 371 3682
rect 399 3686 403 3687
rect 399 3681 403 3682
rect 519 3686 523 3687
rect 519 3681 523 3682
rect 567 3686 571 3687
rect 618 3683 619 3687
rect 623 3683 624 3687
rect 618 3682 624 3683
rect 679 3686 683 3687
rect 567 3681 571 3682
rect 112 3661 114 3681
rect 110 3660 116 3661
rect 368 3660 370 3681
rect 442 3679 448 3680
rect 442 3675 443 3679
rect 447 3675 448 3679
rect 442 3674 448 3675
rect 110 3656 111 3660
rect 115 3656 116 3660
rect 110 3655 116 3656
rect 366 3659 372 3660
rect 366 3655 367 3659
rect 371 3655 372 3659
rect 366 3654 372 3655
rect 444 3652 446 3674
rect 520 3660 522 3681
rect 518 3659 524 3660
rect 518 3655 519 3659
rect 523 3655 524 3659
rect 518 3654 524 3655
rect 620 3652 622 3682
rect 679 3681 683 3682
rect 751 3686 755 3687
rect 751 3681 755 3682
rect 847 3686 851 3687
rect 847 3681 851 3682
rect 935 3686 939 3687
rect 935 3681 939 3682
rect 1015 3686 1019 3687
rect 1015 3681 1019 3682
rect 1127 3686 1131 3687
rect 1127 3681 1131 3682
rect 1175 3686 1179 3687
rect 1175 3681 1179 3682
rect 1311 3686 1315 3687
rect 1311 3681 1315 3682
rect 1327 3686 1331 3687
rect 1458 3683 1459 3687
rect 1463 3683 1464 3687
rect 1458 3682 1464 3683
rect 1479 3686 1483 3687
rect 1327 3681 1331 3682
rect 680 3660 682 3681
rect 762 3679 768 3680
rect 762 3675 763 3679
rect 767 3675 768 3679
rect 762 3674 768 3675
rect 678 3659 684 3660
rect 678 3655 679 3659
rect 683 3655 684 3659
rect 678 3654 684 3655
rect 764 3652 766 3674
rect 848 3660 850 3681
rect 1016 3660 1018 3681
rect 1176 3660 1178 3681
rect 1250 3679 1256 3680
rect 1250 3675 1251 3679
rect 1255 3675 1256 3679
rect 1250 3674 1256 3675
rect 846 3659 852 3660
rect 846 3655 847 3659
rect 851 3655 852 3659
rect 846 3654 852 3655
rect 1014 3659 1020 3660
rect 1014 3655 1015 3659
rect 1019 3655 1020 3659
rect 1014 3654 1020 3655
rect 1174 3659 1180 3660
rect 1174 3655 1175 3659
rect 1179 3655 1180 3659
rect 1174 3654 1180 3655
rect 1252 3652 1254 3674
rect 1328 3660 1330 3681
rect 1402 3679 1408 3680
rect 1402 3675 1403 3679
rect 1407 3675 1408 3679
rect 1402 3674 1408 3675
rect 1326 3659 1332 3660
rect 1326 3655 1327 3659
rect 1331 3655 1332 3659
rect 1326 3654 1332 3655
rect 1404 3652 1406 3674
rect 442 3651 448 3652
rect 442 3647 443 3651
rect 447 3647 448 3651
rect 618 3651 624 3652
rect 442 3646 448 3647
rect 594 3647 600 3648
rect 110 3643 116 3644
rect 110 3639 111 3643
rect 115 3639 116 3643
rect 594 3643 595 3647
rect 599 3643 600 3647
rect 618 3647 619 3651
rect 623 3647 624 3651
rect 618 3646 624 3647
rect 762 3651 768 3652
rect 762 3647 763 3651
rect 767 3647 768 3651
rect 762 3646 768 3647
rect 1250 3651 1256 3652
rect 1250 3647 1251 3651
rect 1255 3647 1256 3651
rect 1250 3646 1256 3647
rect 1402 3651 1408 3652
rect 1402 3647 1403 3651
rect 1407 3647 1408 3651
rect 1402 3646 1408 3647
rect 594 3642 600 3643
rect 110 3638 116 3639
rect 366 3640 372 3641
rect 112 3603 114 3638
rect 366 3636 367 3640
rect 371 3636 372 3640
rect 366 3635 372 3636
rect 518 3640 524 3641
rect 518 3636 519 3640
rect 523 3636 524 3640
rect 518 3635 524 3636
rect 368 3603 370 3635
rect 520 3603 522 3635
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 271 3602 275 3603
rect 271 3597 275 3598
rect 367 3602 371 3603
rect 367 3597 371 3598
rect 415 3602 419 3603
rect 415 3597 419 3598
rect 519 3602 523 3603
rect 519 3597 523 3598
rect 575 3602 579 3603
rect 575 3597 579 3598
rect 112 3570 114 3597
rect 272 3573 274 3597
rect 416 3573 418 3597
rect 576 3573 578 3597
rect 270 3572 276 3573
rect 110 3569 116 3570
rect 110 3565 111 3569
rect 115 3565 116 3569
rect 270 3568 271 3572
rect 275 3568 276 3572
rect 270 3567 276 3568
rect 414 3572 420 3573
rect 414 3568 415 3572
rect 419 3568 420 3572
rect 414 3567 420 3568
rect 574 3572 580 3573
rect 574 3568 575 3572
rect 579 3568 580 3572
rect 574 3567 580 3568
rect 110 3564 116 3565
rect 346 3563 352 3564
rect 346 3559 347 3563
rect 351 3559 352 3563
rect 346 3558 352 3559
rect 482 3563 488 3564
rect 482 3559 483 3563
rect 487 3559 488 3563
rect 482 3558 488 3559
rect 270 3553 276 3554
rect 110 3552 116 3553
rect 110 3548 111 3552
rect 115 3548 116 3552
rect 270 3549 271 3553
rect 275 3549 276 3553
rect 270 3548 276 3549
rect 110 3547 116 3548
rect 112 3519 114 3547
rect 272 3519 274 3548
rect 348 3536 350 3558
rect 414 3553 420 3554
rect 414 3549 415 3553
rect 419 3549 420 3553
rect 414 3548 420 3549
rect 346 3535 352 3536
rect 346 3531 347 3535
rect 351 3531 352 3535
rect 346 3530 352 3531
rect 416 3519 418 3548
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 159 3518 163 3519
rect 159 3513 163 3514
rect 271 3518 275 3519
rect 271 3513 275 3514
rect 287 3518 291 3519
rect 287 3513 291 3514
rect 415 3518 419 3519
rect 415 3513 419 3514
rect 423 3518 427 3519
rect 423 3513 427 3514
rect 112 3493 114 3513
rect 110 3492 116 3493
rect 160 3492 162 3513
rect 234 3511 240 3512
rect 234 3507 235 3511
rect 239 3507 240 3511
rect 234 3506 240 3507
rect 110 3488 111 3492
rect 115 3488 116 3492
rect 110 3487 116 3488
rect 158 3491 164 3492
rect 158 3487 159 3491
rect 163 3487 164 3491
rect 158 3486 164 3487
rect 236 3484 238 3506
rect 288 3492 290 3513
rect 424 3492 426 3513
rect 484 3512 486 3558
rect 574 3553 580 3554
rect 574 3549 575 3553
rect 579 3549 580 3553
rect 574 3548 580 3549
rect 576 3519 578 3548
rect 596 3536 598 3642
rect 678 3640 684 3641
rect 678 3636 679 3640
rect 683 3636 684 3640
rect 678 3635 684 3636
rect 846 3640 852 3641
rect 846 3636 847 3640
rect 851 3636 852 3640
rect 846 3635 852 3636
rect 1014 3640 1020 3641
rect 1014 3636 1015 3640
rect 1019 3636 1020 3640
rect 1014 3635 1020 3636
rect 1174 3640 1180 3641
rect 1174 3636 1175 3640
rect 1179 3636 1180 3640
rect 1174 3635 1180 3636
rect 1326 3640 1332 3641
rect 1326 3636 1327 3640
rect 1331 3636 1332 3640
rect 1326 3635 1332 3636
rect 680 3603 682 3635
rect 848 3603 850 3635
rect 1016 3603 1018 3635
rect 1176 3603 1178 3635
rect 1328 3603 1330 3635
rect 679 3602 683 3603
rect 679 3597 683 3598
rect 735 3602 739 3603
rect 735 3597 739 3598
rect 847 3602 851 3603
rect 847 3597 851 3598
rect 895 3602 899 3603
rect 895 3597 899 3598
rect 1015 3602 1019 3603
rect 1015 3597 1019 3598
rect 1055 3602 1059 3603
rect 1055 3597 1059 3598
rect 1175 3602 1179 3603
rect 1175 3597 1179 3598
rect 1215 3602 1219 3603
rect 1215 3597 1219 3598
rect 1327 3602 1331 3603
rect 1327 3597 1331 3598
rect 1375 3602 1379 3603
rect 1375 3597 1379 3598
rect 736 3573 738 3597
rect 896 3573 898 3597
rect 1056 3573 1058 3597
rect 1216 3573 1218 3597
rect 1376 3573 1378 3597
rect 734 3572 740 3573
rect 734 3568 735 3572
rect 739 3568 740 3572
rect 734 3567 740 3568
rect 894 3572 900 3573
rect 894 3568 895 3572
rect 899 3568 900 3572
rect 894 3567 900 3568
rect 1054 3572 1060 3573
rect 1054 3568 1055 3572
rect 1059 3568 1060 3572
rect 1054 3567 1060 3568
rect 1214 3572 1220 3573
rect 1214 3568 1215 3572
rect 1219 3568 1220 3572
rect 1214 3567 1220 3568
rect 1374 3572 1380 3573
rect 1374 3568 1375 3572
rect 1379 3568 1380 3572
rect 1374 3567 1380 3568
rect 1460 3564 1462 3682
rect 1479 3681 1483 3682
rect 1503 3686 1507 3687
rect 1503 3681 1507 3682
rect 1631 3686 1635 3687
rect 1631 3681 1635 3682
rect 1695 3686 1699 3687
rect 1695 3681 1699 3682
rect 1791 3686 1795 3687
rect 1791 3681 1795 3682
rect 1480 3660 1482 3681
rect 1554 3679 1560 3680
rect 1554 3675 1555 3679
rect 1559 3675 1560 3679
rect 1554 3674 1560 3675
rect 1478 3659 1484 3660
rect 1478 3655 1479 3659
rect 1483 3655 1484 3659
rect 1478 3654 1484 3655
rect 1556 3652 1558 3674
rect 1632 3660 1634 3681
rect 1706 3679 1712 3680
rect 1706 3675 1707 3679
rect 1711 3675 1712 3679
rect 1706 3674 1712 3675
rect 1630 3659 1636 3660
rect 1630 3655 1631 3659
rect 1635 3655 1636 3659
rect 1630 3654 1636 3655
rect 1708 3652 1710 3674
rect 1792 3660 1794 3681
rect 1790 3659 1796 3660
rect 1790 3655 1791 3659
rect 1795 3655 1796 3659
rect 1790 3654 1796 3655
rect 1868 3652 1870 3698
rect 1888 3687 1890 3720
rect 2006 3719 2012 3720
rect 2008 3687 2010 3719
rect 2048 3715 2050 3747
rect 2072 3715 2074 3748
rect 2047 3714 2051 3715
rect 2047 3709 2051 3710
rect 2071 3714 2075 3715
rect 2071 3709 2075 3710
rect 2048 3689 2050 3709
rect 2046 3688 2052 3689
rect 2072 3688 2074 3709
rect 2140 3708 2142 3758
rect 2198 3753 2204 3754
rect 2198 3749 2199 3753
rect 2203 3749 2204 3753
rect 2198 3748 2204 3749
rect 2200 3715 2202 3748
rect 2304 3736 2306 3758
rect 2374 3753 2380 3754
rect 2374 3749 2375 3753
rect 2379 3749 2380 3753
rect 2374 3748 2380 3749
rect 2558 3753 2564 3754
rect 2558 3749 2559 3753
rect 2563 3749 2564 3753
rect 2558 3748 2564 3749
rect 2302 3735 2308 3736
rect 2302 3731 2303 3735
rect 2307 3731 2308 3735
rect 2302 3730 2308 3731
rect 2376 3715 2378 3748
rect 2560 3715 2562 3748
rect 2596 3736 2598 3834
rect 2670 3832 2676 3833
rect 2670 3828 2671 3832
rect 2675 3828 2676 3832
rect 2670 3827 2676 3828
rect 2830 3832 2836 3833
rect 2830 3828 2831 3832
rect 2835 3828 2836 3832
rect 2830 3827 2836 3828
rect 2990 3832 2996 3833
rect 2990 3828 2991 3832
rect 2995 3828 2996 3832
rect 2990 3827 2996 3828
rect 2672 3803 2674 3827
rect 2832 3803 2834 3827
rect 2992 3803 2994 3827
rect 2671 3802 2675 3803
rect 2671 3797 2675 3798
rect 2751 3802 2755 3803
rect 2751 3797 2755 3798
rect 2831 3802 2835 3803
rect 2831 3797 2835 3798
rect 2951 3802 2955 3803
rect 2951 3797 2955 3798
rect 2991 3802 2995 3803
rect 2991 3797 2995 3798
rect 2752 3773 2754 3797
rect 2952 3773 2954 3797
rect 2750 3772 2756 3773
rect 2750 3768 2751 3772
rect 2755 3768 2756 3772
rect 2750 3767 2756 3768
rect 2950 3772 2956 3773
rect 2950 3768 2951 3772
rect 2955 3768 2956 3772
rect 2950 3767 2956 3768
rect 3028 3764 3030 3866
rect 3068 3844 3070 3866
rect 3080 3844 3082 3874
rect 3159 3873 3163 3874
rect 3175 3878 3179 3879
rect 3175 3873 3179 3874
rect 3295 3878 3299 3879
rect 3295 3873 3299 3874
rect 3327 3878 3331 3879
rect 3327 3873 3331 3874
rect 3415 3878 3419 3879
rect 3415 3873 3419 3874
rect 3495 3878 3499 3879
rect 3495 3873 3499 3874
rect 3535 3878 3539 3879
rect 3535 3873 3539 3874
rect 3160 3852 3162 3873
rect 3328 3852 3330 3873
rect 3496 3852 3498 3873
rect 3612 3872 3614 3910
rect 3942 3904 3948 3905
rect 3942 3900 3943 3904
rect 3947 3900 3948 3904
rect 3942 3899 3948 3900
rect 3944 3879 3946 3899
rect 3663 3878 3667 3879
rect 3663 3873 3667 3874
rect 3943 3878 3947 3879
rect 3943 3873 3947 3874
rect 3602 3871 3608 3872
rect 3602 3867 3603 3871
rect 3607 3867 3608 3871
rect 3602 3866 3608 3867
rect 3610 3871 3616 3872
rect 3610 3867 3611 3871
rect 3615 3867 3616 3871
rect 3610 3866 3616 3867
rect 3158 3851 3164 3852
rect 3158 3847 3159 3851
rect 3163 3847 3164 3851
rect 3158 3846 3164 3847
rect 3326 3851 3332 3852
rect 3326 3847 3327 3851
rect 3331 3847 3332 3851
rect 3326 3846 3332 3847
rect 3494 3851 3500 3852
rect 3494 3847 3495 3851
rect 3499 3847 3500 3851
rect 3494 3846 3500 3847
rect 3604 3844 3606 3866
rect 3664 3852 3666 3873
rect 3944 3853 3946 3873
rect 3942 3852 3948 3853
rect 3662 3851 3668 3852
rect 3662 3847 3663 3851
rect 3667 3847 3668 3851
rect 3942 3848 3943 3852
rect 3947 3848 3948 3852
rect 3942 3847 3948 3848
rect 3662 3846 3668 3847
rect 3066 3843 3072 3844
rect 3066 3839 3067 3843
rect 3071 3839 3072 3843
rect 3066 3838 3072 3839
rect 3078 3843 3084 3844
rect 3078 3839 3079 3843
rect 3083 3839 3084 3843
rect 3602 3843 3608 3844
rect 3078 3838 3084 3839
rect 3402 3839 3408 3840
rect 3402 3835 3403 3839
rect 3407 3835 3408 3839
rect 3602 3839 3603 3843
rect 3607 3839 3608 3843
rect 3602 3838 3608 3839
rect 3402 3834 3408 3835
rect 3942 3835 3948 3836
rect 3158 3832 3164 3833
rect 3158 3828 3159 3832
rect 3163 3828 3164 3832
rect 3158 3827 3164 3828
rect 3326 3832 3332 3833
rect 3326 3828 3327 3832
rect 3331 3828 3332 3832
rect 3326 3827 3332 3828
rect 3160 3803 3162 3827
rect 3328 3803 3330 3827
rect 3143 3802 3147 3803
rect 3143 3797 3147 3798
rect 3159 3802 3163 3803
rect 3159 3797 3163 3798
rect 3327 3802 3331 3803
rect 3327 3797 3331 3798
rect 3335 3802 3339 3803
rect 3335 3797 3339 3798
rect 3144 3773 3146 3797
rect 3336 3773 3338 3797
rect 3142 3772 3148 3773
rect 3142 3768 3143 3772
rect 3147 3768 3148 3772
rect 3142 3767 3148 3768
rect 3334 3772 3340 3773
rect 3334 3768 3335 3772
rect 3339 3768 3340 3772
rect 3334 3767 3340 3768
rect 2634 3763 2640 3764
rect 2634 3759 2635 3763
rect 2639 3759 2640 3763
rect 2634 3758 2640 3759
rect 2642 3763 2648 3764
rect 2642 3759 2643 3763
rect 2647 3759 2648 3763
rect 2642 3758 2648 3759
rect 3026 3763 3032 3764
rect 3026 3759 3027 3763
rect 3031 3759 3032 3763
rect 3026 3758 3032 3759
rect 3046 3763 3052 3764
rect 3046 3759 3047 3763
rect 3051 3759 3052 3763
rect 3046 3758 3052 3759
rect 2636 3736 2638 3758
rect 2644 3744 2646 3758
rect 2750 3753 2756 3754
rect 2750 3749 2751 3753
rect 2755 3749 2756 3753
rect 2750 3748 2756 3749
rect 2950 3753 2956 3754
rect 2950 3749 2951 3753
rect 2955 3749 2956 3753
rect 2950 3748 2956 3749
rect 2642 3743 2648 3744
rect 2642 3739 2643 3743
rect 2647 3739 2648 3743
rect 2642 3738 2648 3739
rect 2594 3735 2600 3736
rect 2594 3731 2595 3735
rect 2599 3731 2600 3735
rect 2594 3730 2600 3731
rect 2634 3735 2640 3736
rect 2634 3731 2635 3735
rect 2639 3731 2640 3735
rect 2634 3730 2640 3731
rect 2752 3715 2754 3748
rect 2952 3715 2954 3748
rect 3048 3736 3050 3758
rect 3142 3753 3148 3754
rect 3142 3749 3143 3753
rect 3147 3749 3148 3753
rect 3142 3748 3148 3749
rect 3334 3753 3340 3754
rect 3334 3749 3335 3753
rect 3339 3749 3340 3753
rect 3334 3748 3340 3749
rect 3046 3735 3052 3736
rect 3046 3731 3047 3735
rect 3051 3731 3052 3735
rect 3046 3730 3052 3731
rect 3144 3715 3146 3748
rect 3194 3731 3200 3732
rect 3194 3727 3195 3731
rect 3199 3727 3200 3731
rect 3194 3726 3200 3727
rect 2199 3714 2203 3715
rect 2199 3709 2203 3710
rect 2263 3714 2267 3715
rect 2263 3709 2267 3710
rect 2375 3714 2379 3715
rect 2375 3709 2379 3710
rect 2479 3714 2483 3715
rect 2479 3709 2483 3710
rect 2559 3714 2563 3715
rect 2559 3709 2563 3710
rect 2695 3714 2699 3715
rect 2695 3709 2699 3710
rect 2751 3714 2755 3715
rect 2751 3709 2755 3710
rect 2911 3714 2915 3715
rect 2911 3709 2915 3710
rect 2951 3714 2955 3715
rect 2951 3709 2955 3710
rect 3119 3714 3123 3715
rect 3119 3709 3123 3710
rect 3143 3714 3147 3715
rect 3143 3709 3147 3710
rect 2138 3707 2144 3708
rect 2138 3703 2139 3707
rect 2143 3703 2144 3707
rect 2138 3702 2144 3703
rect 2146 3707 2152 3708
rect 2146 3703 2147 3707
rect 2151 3703 2152 3707
rect 2146 3702 2152 3703
rect 1887 3686 1891 3687
rect 1887 3681 1891 3682
rect 2007 3686 2011 3687
rect 2046 3684 2047 3688
rect 2051 3684 2052 3688
rect 2046 3683 2052 3684
rect 2070 3687 2076 3688
rect 2070 3683 2071 3687
rect 2075 3683 2076 3687
rect 2070 3682 2076 3683
rect 2007 3681 2011 3682
rect 2008 3661 2010 3681
rect 2148 3680 2150 3702
rect 2264 3688 2266 3709
rect 2338 3707 2344 3708
rect 2338 3703 2339 3707
rect 2343 3703 2344 3707
rect 2338 3702 2344 3703
rect 2262 3687 2268 3688
rect 2262 3683 2263 3687
rect 2267 3683 2268 3687
rect 2262 3682 2268 3683
rect 2340 3680 2342 3702
rect 2480 3688 2482 3709
rect 2696 3688 2698 3709
rect 2912 3688 2914 3709
rect 2986 3707 2992 3708
rect 2986 3703 2987 3707
rect 2991 3703 2992 3707
rect 2986 3702 2992 3703
rect 2478 3687 2484 3688
rect 2478 3683 2479 3687
rect 2483 3683 2484 3687
rect 2478 3682 2484 3683
rect 2694 3687 2700 3688
rect 2694 3683 2695 3687
rect 2699 3683 2700 3687
rect 2694 3682 2700 3683
rect 2910 3687 2916 3688
rect 2910 3683 2911 3687
rect 2915 3683 2916 3687
rect 2910 3682 2916 3683
rect 2988 3680 2990 3702
rect 3018 3699 3024 3700
rect 3018 3695 3019 3699
rect 3023 3695 3024 3699
rect 3018 3694 3024 3695
rect 2146 3679 2152 3680
rect 2146 3675 2147 3679
rect 2151 3675 2152 3679
rect 2146 3674 2152 3675
rect 2338 3679 2344 3680
rect 2338 3675 2339 3679
rect 2343 3675 2344 3679
rect 2338 3674 2344 3675
rect 2662 3679 2668 3680
rect 2662 3675 2663 3679
rect 2667 3675 2668 3679
rect 2662 3674 2668 3675
rect 2986 3679 2992 3680
rect 2986 3675 2987 3679
rect 2991 3675 2992 3679
rect 2986 3674 2992 3675
rect 2046 3671 2052 3672
rect 2046 3667 2047 3671
rect 2051 3667 2052 3671
rect 2046 3666 2052 3667
rect 2070 3668 2076 3669
rect 2006 3660 2012 3661
rect 2006 3656 2007 3660
rect 2011 3656 2012 3660
rect 2006 3655 2012 3656
rect 1554 3651 1560 3652
rect 1554 3647 1555 3651
rect 1559 3647 1560 3651
rect 1554 3646 1560 3647
rect 1706 3651 1712 3652
rect 1706 3647 1707 3651
rect 1711 3647 1712 3651
rect 1706 3646 1712 3647
rect 1866 3651 1872 3652
rect 1866 3647 1867 3651
rect 1871 3647 1872 3651
rect 1866 3646 1872 3647
rect 2006 3643 2012 3644
rect 1478 3640 1484 3641
rect 1478 3636 1479 3640
rect 1483 3636 1484 3640
rect 1478 3635 1484 3636
rect 1630 3640 1636 3641
rect 1630 3636 1631 3640
rect 1635 3636 1636 3640
rect 1630 3635 1636 3636
rect 1790 3640 1796 3641
rect 1790 3636 1791 3640
rect 1795 3636 1796 3640
rect 2006 3639 2007 3643
rect 2011 3639 2012 3643
rect 2006 3638 2012 3639
rect 1790 3635 1796 3636
rect 1480 3603 1482 3635
rect 1632 3603 1634 3635
rect 1792 3603 1794 3635
rect 2008 3603 2010 3638
rect 2048 3635 2050 3666
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 2262 3668 2268 3669
rect 2262 3664 2263 3668
rect 2267 3664 2268 3668
rect 2262 3663 2268 3664
rect 2478 3668 2484 3669
rect 2478 3664 2479 3668
rect 2483 3664 2484 3668
rect 2478 3663 2484 3664
rect 2072 3635 2074 3663
rect 2264 3635 2266 3663
rect 2480 3635 2482 3663
rect 2047 3634 2051 3635
rect 2047 3629 2051 3630
rect 2071 3634 2075 3635
rect 2071 3629 2075 3630
rect 2111 3634 2115 3635
rect 2111 3629 2115 3630
rect 2263 3634 2267 3635
rect 2263 3629 2267 3630
rect 2271 3634 2275 3635
rect 2271 3629 2275 3630
rect 2455 3634 2459 3635
rect 2455 3629 2459 3630
rect 2479 3634 2483 3635
rect 2479 3629 2483 3630
rect 2655 3634 2659 3635
rect 2655 3629 2659 3630
rect 1479 3602 1483 3603
rect 1479 3597 1483 3598
rect 1543 3602 1547 3603
rect 1543 3597 1547 3598
rect 1631 3602 1635 3603
rect 1631 3597 1635 3598
rect 1791 3602 1795 3603
rect 1791 3597 1795 3598
rect 2007 3602 2011 3603
rect 2048 3602 2050 3629
rect 2112 3605 2114 3629
rect 2272 3605 2274 3629
rect 2456 3605 2458 3629
rect 2656 3605 2658 3629
rect 2110 3604 2116 3605
rect 2007 3597 2011 3598
rect 2046 3601 2052 3602
rect 2046 3597 2047 3601
rect 2051 3597 2052 3601
rect 2110 3600 2111 3604
rect 2115 3600 2116 3604
rect 2110 3599 2116 3600
rect 2270 3604 2276 3605
rect 2270 3600 2271 3604
rect 2275 3600 2276 3604
rect 2270 3599 2276 3600
rect 2454 3604 2460 3605
rect 2454 3600 2455 3604
rect 2459 3600 2460 3604
rect 2454 3599 2460 3600
rect 2654 3604 2660 3605
rect 2654 3600 2655 3604
rect 2659 3600 2660 3604
rect 2654 3599 2660 3600
rect 1544 3573 1546 3597
rect 1542 3572 1548 3573
rect 1542 3568 1543 3572
rect 1547 3568 1548 3572
rect 2008 3570 2010 3597
rect 2046 3596 2052 3597
rect 2186 3595 2192 3596
rect 2186 3591 2187 3595
rect 2191 3591 2192 3595
rect 2186 3590 2192 3591
rect 2346 3595 2352 3596
rect 2346 3591 2347 3595
rect 2351 3591 2352 3595
rect 2346 3590 2352 3591
rect 2530 3595 2536 3596
rect 2530 3591 2531 3595
rect 2535 3591 2536 3595
rect 2530 3590 2536 3591
rect 2110 3585 2116 3586
rect 2046 3584 2052 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2110 3581 2111 3585
rect 2115 3581 2116 3585
rect 2110 3580 2116 3581
rect 2046 3579 2052 3580
rect 1542 3567 1548 3568
rect 2006 3569 2012 3570
rect 2006 3565 2007 3569
rect 2011 3565 2012 3569
rect 2006 3564 2012 3565
rect 650 3563 656 3564
rect 650 3559 651 3563
rect 655 3559 656 3563
rect 650 3558 656 3559
rect 810 3563 816 3564
rect 810 3559 811 3563
rect 815 3559 816 3563
rect 810 3558 816 3559
rect 818 3563 824 3564
rect 818 3559 819 3563
rect 823 3559 824 3563
rect 818 3558 824 3559
rect 1130 3563 1136 3564
rect 1130 3559 1131 3563
rect 1135 3559 1136 3563
rect 1130 3558 1136 3559
rect 1290 3563 1296 3564
rect 1290 3559 1291 3563
rect 1295 3559 1296 3563
rect 1290 3558 1296 3559
rect 1450 3563 1456 3564
rect 1450 3559 1451 3563
rect 1455 3559 1456 3563
rect 1450 3558 1456 3559
rect 1458 3563 1464 3564
rect 1458 3559 1459 3563
rect 1463 3559 1464 3563
rect 1458 3558 1464 3559
rect 652 3536 654 3558
rect 734 3553 740 3554
rect 734 3549 735 3553
rect 739 3549 740 3553
rect 734 3548 740 3549
rect 594 3535 600 3536
rect 594 3531 595 3535
rect 599 3531 600 3535
rect 594 3530 600 3531
rect 650 3535 656 3536
rect 650 3531 651 3535
rect 655 3531 656 3535
rect 650 3530 656 3531
rect 736 3519 738 3548
rect 812 3536 814 3558
rect 820 3544 822 3558
rect 894 3553 900 3554
rect 894 3549 895 3553
rect 899 3549 900 3553
rect 894 3548 900 3549
rect 1054 3553 1060 3554
rect 1054 3549 1055 3553
rect 1059 3549 1060 3553
rect 1054 3548 1060 3549
rect 818 3543 824 3544
rect 818 3539 819 3543
rect 823 3539 824 3543
rect 818 3538 824 3539
rect 810 3535 816 3536
rect 810 3531 811 3535
rect 815 3531 816 3535
rect 810 3530 816 3531
rect 896 3519 898 3548
rect 1056 3519 1058 3548
rect 1132 3540 1134 3558
rect 1214 3553 1220 3554
rect 1214 3549 1215 3553
rect 1219 3549 1220 3553
rect 1214 3548 1220 3549
rect 1130 3539 1136 3540
rect 1130 3535 1131 3539
rect 1135 3535 1136 3539
rect 1130 3534 1136 3535
rect 1216 3519 1218 3548
rect 1292 3536 1294 3558
rect 1374 3553 1380 3554
rect 1374 3549 1375 3553
rect 1379 3549 1380 3553
rect 1374 3548 1380 3549
rect 1290 3535 1296 3536
rect 1290 3531 1291 3535
rect 1295 3531 1296 3535
rect 1290 3530 1296 3531
rect 1338 3527 1344 3528
rect 1338 3523 1339 3527
rect 1343 3523 1344 3527
rect 1338 3522 1344 3523
rect 559 3518 563 3519
rect 559 3513 563 3514
rect 575 3518 579 3519
rect 575 3513 579 3514
rect 695 3518 699 3519
rect 695 3513 699 3514
rect 735 3518 739 3519
rect 735 3513 739 3514
rect 831 3518 835 3519
rect 831 3513 835 3514
rect 895 3518 899 3519
rect 895 3513 899 3514
rect 967 3518 971 3519
rect 967 3513 971 3514
rect 1055 3518 1059 3519
rect 1055 3513 1059 3514
rect 1095 3518 1099 3519
rect 1095 3513 1099 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1231 3518 1235 3519
rect 1231 3513 1235 3514
rect 482 3511 488 3512
rect 482 3507 483 3511
rect 487 3507 488 3511
rect 482 3506 488 3507
rect 498 3511 504 3512
rect 498 3507 499 3511
rect 503 3507 504 3511
rect 498 3506 504 3507
rect 286 3491 292 3492
rect 286 3487 287 3491
rect 291 3487 292 3491
rect 286 3486 292 3487
rect 422 3491 428 3492
rect 422 3487 423 3491
rect 427 3487 428 3491
rect 422 3486 428 3487
rect 500 3484 502 3506
rect 560 3492 562 3513
rect 634 3511 640 3512
rect 634 3507 635 3511
rect 639 3507 640 3511
rect 634 3506 640 3507
rect 558 3491 564 3492
rect 558 3487 559 3491
rect 563 3487 564 3491
rect 558 3486 564 3487
rect 636 3484 638 3506
rect 642 3503 648 3504
rect 642 3499 643 3503
rect 647 3499 648 3503
rect 642 3498 648 3499
rect 644 3484 646 3498
rect 696 3492 698 3513
rect 832 3492 834 3513
rect 882 3511 888 3512
rect 882 3507 883 3511
rect 887 3507 888 3511
rect 882 3506 888 3507
rect 906 3511 912 3512
rect 906 3507 907 3511
rect 911 3507 912 3511
rect 906 3506 912 3507
rect 694 3491 700 3492
rect 694 3487 695 3491
rect 699 3487 700 3491
rect 694 3486 700 3487
rect 830 3491 836 3492
rect 830 3487 831 3491
rect 835 3487 836 3491
rect 830 3486 836 3487
rect 234 3483 240 3484
rect 234 3479 235 3483
rect 239 3479 240 3483
rect 498 3483 504 3484
rect 234 3478 240 3479
rect 362 3479 368 3480
rect 110 3475 116 3476
rect 110 3471 111 3475
rect 115 3471 116 3475
rect 362 3475 363 3479
rect 367 3475 368 3479
rect 498 3479 499 3483
rect 503 3479 504 3483
rect 498 3478 504 3479
rect 634 3483 640 3484
rect 634 3479 635 3483
rect 639 3479 640 3483
rect 634 3478 640 3479
rect 642 3483 648 3484
rect 642 3479 643 3483
rect 647 3479 648 3483
rect 642 3478 648 3479
rect 362 3474 368 3475
rect 110 3470 116 3471
rect 158 3472 164 3473
rect 112 3435 114 3470
rect 158 3468 159 3472
rect 163 3468 164 3472
rect 158 3467 164 3468
rect 286 3472 292 3473
rect 286 3468 287 3472
rect 291 3468 292 3472
rect 286 3467 292 3468
rect 160 3435 162 3467
rect 288 3435 290 3467
rect 111 3434 115 3435
rect 111 3429 115 3430
rect 135 3434 139 3435
rect 135 3429 139 3430
rect 159 3434 163 3435
rect 159 3429 163 3430
rect 247 3434 251 3435
rect 247 3429 251 3430
rect 287 3434 291 3435
rect 287 3429 291 3430
rect 112 3402 114 3429
rect 136 3405 138 3429
rect 248 3405 250 3429
rect 134 3404 140 3405
rect 110 3401 116 3402
rect 110 3397 111 3401
rect 115 3397 116 3401
rect 134 3400 135 3404
rect 139 3400 140 3404
rect 134 3399 140 3400
rect 246 3404 252 3405
rect 246 3400 247 3404
rect 251 3400 252 3404
rect 246 3399 252 3400
rect 110 3396 116 3397
rect 202 3395 208 3396
rect 202 3391 203 3395
rect 207 3391 208 3395
rect 202 3390 208 3391
rect 218 3395 224 3396
rect 218 3391 219 3395
rect 223 3391 224 3395
rect 218 3390 224 3391
rect 134 3385 140 3386
rect 110 3384 116 3385
rect 110 3380 111 3384
rect 115 3380 116 3384
rect 134 3381 135 3385
rect 139 3381 140 3385
rect 134 3380 140 3381
rect 110 3379 116 3380
rect 112 3351 114 3379
rect 136 3351 138 3380
rect 111 3350 115 3351
rect 111 3345 115 3346
rect 135 3350 139 3351
rect 135 3345 139 3346
rect 112 3325 114 3345
rect 110 3324 116 3325
rect 136 3324 138 3345
rect 204 3344 206 3390
rect 220 3368 222 3390
rect 246 3385 252 3386
rect 246 3381 247 3385
rect 251 3381 252 3385
rect 246 3380 252 3381
rect 218 3367 224 3368
rect 218 3363 219 3367
rect 223 3363 224 3367
rect 218 3362 224 3363
rect 248 3351 250 3380
rect 364 3368 366 3474
rect 422 3472 428 3473
rect 422 3468 423 3472
rect 427 3468 428 3472
rect 422 3467 428 3468
rect 558 3472 564 3473
rect 558 3468 559 3472
rect 563 3468 564 3472
rect 558 3467 564 3468
rect 694 3472 700 3473
rect 694 3468 695 3472
rect 699 3468 700 3472
rect 694 3467 700 3468
rect 830 3472 836 3473
rect 830 3468 831 3472
rect 835 3468 836 3472
rect 830 3467 836 3468
rect 424 3435 426 3467
rect 560 3435 562 3467
rect 696 3435 698 3467
rect 832 3435 834 3467
rect 383 3434 387 3435
rect 383 3429 387 3430
rect 423 3434 427 3435
rect 423 3429 427 3430
rect 527 3434 531 3435
rect 527 3429 531 3430
rect 559 3434 563 3435
rect 559 3429 563 3430
rect 671 3434 675 3435
rect 671 3429 675 3430
rect 695 3434 699 3435
rect 695 3429 699 3430
rect 815 3434 819 3435
rect 815 3429 819 3430
rect 831 3434 835 3435
rect 831 3429 835 3430
rect 384 3405 386 3429
rect 528 3405 530 3429
rect 672 3405 674 3429
rect 816 3405 818 3429
rect 382 3404 388 3405
rect 382 3400 383 3404
rect 387 3400 388 3404
rect 382 3399 388 3400
rect 526 3404 532 3405
rect 526 3400 527 3404
rect 531 3400 532 3404
rect 526 3399 532 3400
rect 670 3404 676 3405
rect 670 3400 671 3404
rect 675 3400 676 3404
rect 670 3399 676 3400
rect 814 3404 820 3405
rect 814 3400 815 3404
rect 819 3400 820 3404
rect 814 3399 820 3400
rect 884 3396 886 3506
rect 908 3484 910 3506
rect 968 3492 970 3513
rect 1042 3511 1048 3512
rect 1042 3507 1043 3511
rect 1047 3507 1048 3511
rect 1042 3506 1048 3507
rect 966 3491 972 3492
rect 966 3487 967 3491
rect 971 3487 972 3491
rect 966 3486 972 3487
rect 1044 3484 1046 3506
rect 1096 3492 1098 3513
rect 1170 3511 1176 3512
rect 1170 3507 1171 3511
rect 1175 3507 1176 3511
rect 1170 3506 1176 3507
rect 1094 3491 1100 3492
rect 1094 3487 1095 3491
rect 1099 3487 1100 3491
rect 1094 3486 1100 3487
rect 1172 3484 1174 3506
rect 1232 3492 1234 3513
rect 1306 3511 1312 3512
rect 1306 3507 1307 3511
rect 1311 3507 1312 3511
rect 1306 3506 1312 3507
rect 1230 3491 1236 3492
rect 1230 3487 1231 3491
rect 1235 3487 1236 3491
rect 1230 3486 1236 3487
rect 1308 3484 1310 3506
rect 1340 3484 1342 3522
rect 1376 3519 1378 3548
rect 1452 3536 1454 3558
rect 1542 3553 1548 3554
rect 1542 3549 1543 3553
rect 1547 3549 1548 3553
rect 1542 3548 1548 3549
rect 2006 3552 2012 3553
rect 2006 3548 2007 3552
rect 2011 3548 2012 3552
rect 1450 3535 1456 3536
rect 1450 3531 1451 3535
rect 1455 3531 1456 3535
rect 1450 3530 1456 3531
rect 1544 3519 1546 3548
rect 2006 3547 2012 3548
rect 2008 3519 2010 3547
rect 2048 3543 2050 3579
rect 2112 3543 2114 3580
rect 2188 3568 2190 3590
rect 2270 3585 2276 3586
rect 2270 3581 2271 3585
rect 2275 3581 2276 3585
rect 2270 3580 2276 3581
rect 2186 3567 2192 3568
rect 2186 3563 2187 3567
rect 2191 3563 2192 3567
rect 2186 3562 2192 3563
rect 2272 3543 2274 3580
rect 2348 3568 2350 3590
rect 2454 3585 2460 3586
rect 2454 3581 2455 3585
rect 2459 3581 2460 3585
rect 2454 3580 2460 3581
rect 2346 3567 2352 3568
rect 2346 3563 2347 3567
rect 2351 3563 2352 3567
rect 2346 3562 2352 3563
rect 2456 3543 2458 3580
rect 2532 3568 2534 3590
rect 2654 3585 2660 3586
rect 2654 3581 2655 3585
rect 2659 3581 2660 3585
rect 2654 3580 2660 3581
rect 2530 3567 2536 3568
rect 2530 3563 2531 3567
rect 2535 3563 2536 3567
rect 2530 3562 2536 3563
rect 2656 3543 2658 3580
rect 2664 3576 2666 3674
rect 2694 3668 2700 3669
rect 2694 3664 2695 3668
rect 2699 3664 2700 3668
rect 2694 3663 2700 3664
rect 2910 3668 2916 3669
rect 2910 3664 2911 3668
rect 2915 3664 2916 3668
rect 2910 3663 2916 3664
rect 2696 3635 2698 3663
rect 2912 3635 2914 3663
rect 2695 3634 2699 3635
rect 2695 3629 2699 3630
rect 2871 3634 2875 3635
rect 2871 3629 2875 3630
rect 2911 3634 2915 3635
rect 2911 3629 2915 3630
rect 2872 3605 2874 3629
rect 2870 3604 2876 3605
rect 2870 3600 2871 3604
rect 2875 3600 2876 3604
rect 2870 3599 2876 3600
rect 3020 3596 3022 3694
rect 3120 3688 3122 3709
rect 3118 3687 3124 3688
rect 3118 3683 3119 3687
rect 3123 3683 3124 3687
rect 3118 3682 3124 3683
rect 3196 3680 3198 3726
rect 3336 3715 3338 3748
rect 3404 3736 3406 3834
rect 3494 3832 3500 3833
rect 3494 3828 3495 3832
rect 3499 3828 3500 3832
rect 3494 3827 3500 3828
rect 3662 3832 3668 3833
rect 3662 3828 3663 3832
rect 3667 3828 3668 3832
rect 3942 3831 3943 3835
rect 3947 3831 3948 3835
rect 3942 3830 3948 3831
rect 3662 3827 3668 3828
rect 3496 3803 3498 3827
rect 3664 3803 3666 3827
rect 3944 3803 3946 3830
rect 3495 3802 3499 3803
rect 3495 3797 3499 3798
rect 3535 3802 3539 3803
rect 3535 3797 3539 3798
rect 3663 3802 3667 3803
rect 3663 3797 3667 3798
rect 3735 3802 3739 3803
rect 3735 3797 3739 3798
rect 3943 3802 3947 3803
rect 3943 3797 3947 3798
rect 3536 3773 3538 3797
rect 3736 3773 3738 3797
rect 3534 3772 3540 3773
rect 3534 3768 3535 3772
rect 3539 3768 3540 3772
rect 3534 3767 3540 3768
rect 3734 3772 3740 3773
rect 3734 3768 3735 3772
rect 3739 3768 3740 3772
rect 3944 3770 3946 3797
rect 3734 3767 3740 3768
rect 3942 3769 3948 3770
rect 3942 3765 3943 3769
rect 3947 3765 3948 3769
rect 3942 3764 3948 3765
rect 3410 3763 3416 3764
rect 3410 3759 3411 3763
rect 3415 3759 3416 3763
rect 3410 3758 3416 3759
rect 3610 3763 3616 3764
rect 3610 3759 3611 3763
rect 3615 3759 3616 3763
rect 3610 3758 3616 3759
rect 3802 3763 3808 3764
rect 3802 3759 3803 3763
rect 3807 3759 3808 3763
rect 3802 3758 3808 3759
rect 3412 3736 3414 3758
rect 3534 3753 3540 3754
rect 3534 3749 3535 3753
rect 3539 3749 3540 3753
rect 3534 3748 3540 3749
rect 3402 3735 3408 3736
rect 3402 3731 3403 3735
rect 3407 3731 3408 3735
rect 3402 3730 3408 3731
rect 3410 3735 3416 3736
rect 3410 3731 3411 3735
rect 3415 3731 3416 3735
rect 3410 3730 3416 3731
rect 3536 3715 3538 3748
rect 3612 3736 3614 3758
rect 3734 3753 3740 3754
rect 3734 3749 3735 3753
rect 3739 3749 3740 3753
rect 3734 3748 3740 3749
rect 3610 3735 3616 3736
rect 3610 3731 3611 3735
rect 3615 3731 3616 3735
rect 3610 3730 3616 3731
rect 3736 3715 3738 3748
rect 3319 3714 3323 3715
rect 3319 3709 3323 3710
rect 3335 3714 3339 3715
rect 3335 3709 3339 3710
rect 3519 3714 3523 3715
rect 3519 3709 3523 3710
rect 3535 3714 3539 3715
rect 3535 3709 3539 3710
rect 3727 3714 3731 3715
rect 3727 3709 3731 3710
rect 3735 3714 3739 3715
rect 3735 3709 3739 3710
rect 3320 3688 3322 3709
rect 3394 3707 3400 3708
rect 3394 3703 3395 3707
rect 3399 3703 3400 3707
rect 3394 3702 3400 3703
rect 3318 3687 3324 3688
rect 3318 3683 3319 3687
rect 3323 3683 3324 3687
rect 3318 3682 3324 3683
rect 3396 3680 3398 3702
rect 3520 3688 3522 3709
rect 3618 3699 3624 3700
rect 3618 3695 3619 3699
rect 3623 3695 3624 3699
rect 3618 3694 3624 3695
rect 3518 3687 3524 3688
rect 3518 3683 3519 3687
rect 3523 3683 3524 3687
rect 3518 3682 3524 3683
rect 3620 3680 3622 3694
rect 3728 3688 3730 3709
rect 3804 3708 3806 3758
rect 3942 3752 3948 3753
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 3942 3747 3948 3748
rect 3944 3715 3946 3747
rect 3943 3714 3947 3715
rect 3943 3709 3947 3710
rect 3802 3707 3808 3708
rect 3802 3703 3803 3707
rect 3807 3703 3808 3707
rect 3802 3702 3808 3703
rect 3944 3689 3946 3709
rect 3942 3688 3948 3689
rect 3726 3687 3732 3688
rect 3726 3683 3727 3687
rect 3731 3683 3732 3687
rect 3942 3684 3943 3688
rect 3947 3684 3948 3688
rect 3942 3683 3948 3684
rect 3726 3682 3732 3683
rect 3194 3679 3200 3680
rect 3194 3675 3195 3679
rect 3199 3675 3200 3679
rect 3194 3674 3200 3675
rect 3394 3679 3400 3680
rect 3394 3675 3395 3679
rect 3399 3675 3400 3679
rect 3618 3679 3624 3680
rect 3394 3674 3400 3675
rect 3594 3675 3600 3676
rect 3594 3671 3595 3675
rect 3599 3671 3600 3675
rect 3618 3675 3619 3679
rect 3623 3675 3624 3679
rect 3618 3674 3624 3675
rect 3594 3670 3600 3671
rect 3942 3671 3948 3672
rect 3118 3668 3124 3669
rect 3118 3664 3119 3668
rect 3123 3664 3124 3668
rect 3118 3663 3124 3664
rect 3318 3668 3324 3669
rect 3318 3664 3319 3668
rect 3323 3664 3324 3668
rect 3318 3663 3324 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3120 3635 3122 3663
rect 3320 3635 3322 3663
rect 3520 3635 3522 3663
rect 3095 3634 3099 3635
rect 3095 3629 3099 3630
rect 3119 3634 3123 3635
rect 3119 3629 3123 3630
rect 3319 3634 3323 3635
rect 3319 3629 3323 3630
rect 3327 3634 3331 3635
rect 3327 3629 3331 3630
rect 3519 3634 3523 3635
rect 3519 3629 3523 3630
rect 3567 3634 3571 3635
rect 3567 3629 3571 3630
rect 3096 3605 3098 3629
rect 3328 3605 3330 3629
rect 3568 3605 3570 3629
rect 3094 3604 3100 3605
rect 3094 3600 3095 3604
rect 3099 3600 3100 3604
rect 3094 3599 3100 3600
rect 3326 3604 3332 3605
rect 3326 3600 3327 3604
rect 3331 3600 3332 3604
rect 3326 3599 3332 3600
rect 3566 3604 3572 3605
rect 3566 3600 3567 3604
rect 3571 3600 3572 3604
rect 3566 3599 3572 3600
rect 2730 3595 2736 3596
rect 2730 3591 2731 3595
rect 2735 3591 2736 3595
rect 2730 3590 2736 3591
rect 2862 3595 2868 3596
rect 2862 3591 2863 3595
rect 2867 3591 2868 3595
rect 2862 3590 2868 3591
rect 3018 3595 3024 3596
rect 3018 3591 3019 3595
rect 3023 3591 3024 3595
rect 3018 3590 3024 3591
rect 3394 3595 3400 3596
rect 3394 3591 3395 3595
rect 3399 3591 3400 3595
rect 3394 3590 3400 3591
rect 2662 3575 2668 3576
rect 2662 3571 2663 3575
rect 2667 3571 2668 3575
rect 2662 3570 2668 3571
rect 2732 3568 2734 3590
rect 2730 3567 2736 3568
rect 2730 3563 2731 3567
rect 2735 3563 2736 3567
rect 2730 3562 2736 3563
rect 2047 3542 2051 3543
rect 2047 3537 2051 3538
rect 2111 3542 2115 3543
rect 2111 3537 2115 3538
rect 2271 3542 2275 3543
rect 2271 3537 2275 3538
rect 2287 3542 2291 3543
rect 2287 3537 2291 3538
rect 2383 3542 2387 3543
rect 2383 3537 2387 3538
rect 2455 3542 2459 3543
rect 2455 3537 2459 3538
rect 2479 3542 2483 3543
rect 2479 3537 2483 3538
rect 2575 3542 2579 3543
rect 2575 3537 2579 3538
rect 2655 3542 2659 3543
rect 2655 3537 2659 3538
rect 2671 3542 2675 3543
rect 2671 3537 2675 3538
rect 2767 3542 2771 3543
rect 2767 3537 2771 3538
rect 1367 3518 1371 3519
rect 1367 3513 1371 3514
rect 1375 3518 1379 3519
rect 1375 3513 1379 3514
rect 1543 3518 1547 3519
rect 1543 3513 1547 3514
rect 2007 3518 2011 3519
rect 2048 3517 2050 3537
rect 2007 3513 2011 3514
rect 2046 3516 2052 3517
rect 2288 3516 2290 3537
rect 2354 3535 2360 3536
rect 2354 3531 2355 3535
rect 2359 3531 2360 3535
rect 2354 3530 2360 3531
rect 2362 3535 2368 3536
rect 2362 3531 2363 3535
rect 2367 3531 2368 3535
rect 2362 3530 2368 3531
rect 1368 3492 1370 3513
rect 2008 3493 2010 3513
rect 2046 3512 2047 3516
rect 2051 3512 2052 3516
rect 2046 3511 2052 3512
rect 2286 3515 2292 3516
rect 2286 3511 2287 3515
rect 2291 3511 2292 3515
rect 2286 3510 2292 3511
rect 2356 3501 2358 3530
rect 2364 3508 2366 3530
rect 2384 3516 2386 3537
rect 2466 3535 2472 3536
rect 2466 3531 2467 3535
rect 2471 3531 2472 3535
rect 2466 3530 2472 3531
rect 2382 3515 2388 3516
rect 2382 3511 2383 3515
rect 2387 3511 2388 3515
rect 2382 3510 2388 3511
rect 2468 3508 2470 3530
rect 2480 3516 2482 3537
rect 2554 3535 2560 3536
rect 2554 3531 2555 3535
rect 2559 3531 2560 3535
rect 2554 3530 2560 3531
rect 2478 3515 2484 3516
rect 2478 3511 2479 3515
rect 2483 3511 2484 3515
rect 2478 3510 2484 3511
rect 2556 3508 2558 3530
rect 2576 3516 2578 3537
rect 2672 3516 2674 3537
rect 2738 3535 2744 3536
rect 2738 3531 2739 3535
rect 2743 3531 2744 3535
rect 2738 3530 2744 3531
rect 2746 3535 2752 3536
rect 2746 3531 2747 3535
rect 2751 3531 2752 3535
rect 2746 3530 2752 3531
rect 2574 3515 2580 3516
rect 2574 3511 2575 3515
rect 2579 3511 2580 3515
rect 2574 3510 2580 3511
rect 2670 3515 2676 3516
rect 2670 3511 2671 3515
rect 2675 3511 2676 3515
rect 2670 3510 2676 3511
rect 2362 3507 2368 3508
rect 2362 3503 2363 3507
rect 2367 3503 2368 3507
rect 2362 3502 2368 3503
rect 2466 3507 2472 3508
rect 2466 3503 2467 3507
rect 2471 3503 2472 3507
rect 2466 3502 2472 3503
rect 2554 3507 2560 3508
rect 2554 3503 2555 3507
rect 2559 3503 2560 3507
rect 2554 3502 2560 3503
rect 2355 3500 2359 3501
rect 2046 3499 2052 3500
rect 2046 3495 2047 3499
rect 2051 3495 2052 3499
rect 2046 3494 2052 3495
rect 2286 3496 2292 3497
rect 2006 3492 2012 3493
rect 1366 3491 1372 3492
rect 1366 3487 1367 3491
rect 1371 3487 1372 3491
rect 2006 3488 2007 3492
rect 2011 3488 2012 3492
rect 2006 3487 2012 3488
rect 1366 3486 1372 3487
rect 906 3483 912 3484
rect 906 3479 907 3483
rect 911 3479 912 3483
rect 906 3478 912 3479
rect 1042 3483 1048 3484
rect 1042 3479 1043 3483
rect 1047 3479 1048 3483
rect 1042 3478 1048 3479
rect 1170 3483 1176 3484
rect 1170 3479 1171 3483
rect 1175 3479 1176 3483
rect 1170 3478 1176 3479
rect 1306 3483 1312 3484
rect 1306 3479 1307 3483
rect 1311 3479 1312 3483
rect 1306 3478 1312 3479
rect 1338 3483 1344 3484
rect 1338 3479 1339 3483
rect 1343 3479 1344 3483
rect 1338 3478 1344 3479
rect 2006 3475 2012 3476
rect 966 3472 972 3473
rect 966 3468 967 3472
rect 971 3468 972 3472
rect 966 3467 972 3468
rect 1094 3472 1100 3473
rect 1094 3468 1095 3472
rect 1099 3468 1100 3472
rect 1094 3467 1100 3468
rect 1230 3472 1236 3473
rect 1230 3468 1231 3472
rect 1235 3468 1236 3472
rect 1230 3467 1236 3468
rect 1366 3472 1372 3473
rect 1366 3468 1367 3472
rect 1371 3468 1372 3472
rect 2006 3471 2007 3475
rect 2011 3471 2012 3475
rect 2006 3470 2012 3471
rect 1366 3467 1372 3468
rect 968 3435 970 3467
rect 1096 3435 1098 3467
rect 1232 3435 1234 3467
rect 1368 3435 1370 3467
rect 2008 3435 2010 3470
rect 2048 3467 2050 3494
rect 2286 3492 2287 3496
rect 2291 3492 2292 3496
rect 2546 3499 2552 3500
rect 2355 3495 2359 3496
rect 2382 3496 2388 3497
rect 2286 3491 2292 3492
rect 2382 3492 2383 3496
rect 2387 3492 2388 3496
rect 2382 3491 2388 3492
rect 2478 3496 2484 3497
rect 2478 3492 2479 3496
rect 2483 3492 2484 3496
rect 2546 3495 2547 3499
rect 2551 3495 2552 3499
rect 2740 3499 2742 3530
rect 2748 3508 2750 3530
rect 2768 3516 2770 3537
rect 2842 3535 2848 3536
rect 2842 3531 2843 3535
rect 2847 3531 2848 3535
rect 2842 3530 2848 3531
rect 2766 3515 2772 3516
rect 2766 3511 2767 3515
rect 2771 3511 2772 3515
rect 2766 3510 2772 3511
rect 2844 3508 2846 3530
rect 2746 3507 2752 3508
rect 2746 3503 2747 3507
rect 2751 3503 2752 3507
rect 2746 3502 2752 3503
rect 2842 3507 2848 3508
rect 2842 3503 2843 3507
rect 2847 3503 2848 3507
rect 2842 3502 2848 3503
rect 2864 3501 2866 3590
rect 2870 3585 2876 3586
rect 2870 3581 2871 3585
rect 2875 3581 2876 3585
rect 2870 3580 2876 3581
rect 3094 3585 3100 3586
rect 3094 3581 3095 3585
rect 3099 3581 3100 3585
rect 3094 3580 3100 3581
rect 3326 3585 3332 3586
rect 3326 3581 3327 3585
rect 3331 3581 3332 3585
rect 3326 3580 3332 3581
rect 2872 3543 2874 3580
rect 3096 3543 3098 3580
rect 3190 3563 3196 3564
rect 3190 3559 3191 3563
rect 3195 3559 3196 3563
rect 3190 3558 3196 3559
rect 2871 3542 2875 3543
rect 2871 3537 2875 3538
rect 2983 3542 2987 3543
rect 2983 3537 2987 3538
rect 3095 3542 3099 3543
rect 3095 3537 3099 3538
rect 3103 3542 3107 3543
rect 3103 3537 3107 3538
rect 2872 3516 2874 3537
rect 2946 3535 2952 3536
rect 2946 3531 2947 3535
rect 2951 3531 2952 3535
rect 2946 3530 2952 3531
rect 2870 3515 2876 3516
rect 2870 3511 2871 3515
rect 2875 3511 2876 3515
rect 2870 3510 2876 3511
rect 2948 3508 2950 3530
rect 2984 3516 2986 3537
rect 3058 3535 3064 3536
rect 3058 3531 3059 3535
rect 3063 3531 3064 3535
rect 3058 3530 3064 3531
rect 2982 3515 2988 3516
rect 2982 3511 2983 3515
rect 2987 3511 2988 3515
rect 2982 3510 2988 3511
rect 3060 3508 3062 3530
rect 3104 3516 3106 3537
rect 3102 3515 3108 3516
rect 3102 3511 3103 3515
rect 3107 3511 3108 3515
rect 3102 3510 3108 3511
rect 3192 3508 3194 3558
rect 3328 3543 3330 3580
rect 3223 3542 3227 3543
rect 3223 3537 3227 3538
rect 3327 3542 3331 3543
rect 3327 3537 3331 3538
rect 3351 3542 3355 3543
rect 3351 3537 3355 3538
rect 3224 3516 3226 3537
rect 3230 3535 3236 3536
rect 3230 3531 3231 3535
rect 3235 3531 3236 3535
rect 3230 3530 3236 3531
rect 3222 3515 3228 3516
rect 3222 3511 3223 3515
rect 3227 3511 3228 3515
rect 3222 3510 3228 3511
rect 2946 3507 2952 3508
rect 2946 3503 2947 3507
rect 2951 3503 2952 3507
rect 2946 3502 2952 3503
rect 3058 3507 3064 3508
rect 3058 3503 3059 3507
rect 3063 3503 3064 3507
rect 3058 3502 3064 3503
rect 3066 3507 3072 3508
rect 3066 3503 3067 3507
rect 3071 3503 3072 3507
rect 3066 3502 3072 3503
rect 3190 3507 3196 3508
rect 3190 3503 3191 3507
rect 3195 3503 3196 3507
rect 3190 3502 3196 3503
rect 2863 3500 2867 3501
rect 2740 3497 2750 3499
rect 2546 3494 2552 3495
rect 2574 3496 2580 3497
rect 2478 3491 2484 3492
rect 2288 3467 2290 3491
rect 2384 3467 2386 3491
rect 2480 3467 2482 3491
rect 2047 3466 2051 3467
rect 2047 3461 2051 3462
rect 2287 3466 2291 3467
rect 2287 3461 2291 3462
rect 2383 3466 2387 3467
rect 2383 3461 2387 3462
rect 2479 3466 2483 3467
rect 2479 3461 2483 3462
rect 2487 3466 2491 3467
rect 2487 3461 2491 3462
rect 967 3434 971 3435
rect 967 3429 971 3430
rect 1095 3434 1099 3435
rect 1095 3429 1099 3430
rect 1119 3434 1123 3435
rect 1119 3429 1123 3430
rect 1231 3434 1235 3435
rect 1231 3429 1235 3430
rect 1271 3434 1275 3435
rect 1271 3429 1275 3430
rect 1367 3434 1371 3435
rect 1367 3429 1371 3430
rect 2007 3434 2011 3435
rect 2048 3434 2050 3461
rect 2488 3437 2490 3461
rect 2486 3436 2492 3437
rect 2007 3429 2011 3430
rect 2046 3433 2052 3434
rect 2046 3429 2047 3433
rect 2051 3429 2052 3433
rect 2486 3432 2487 3436
rect 2491 3432 2492 3436
rect 2486 3431 2492 3432
rect 968 3405 970 3429
rect 1120 3405 1122 3429
rect 1272 3405 1274 3429
rect 966 3404 972 3405
rect 966 3400 967 3404
rect 971 3400 972 3404
rect 966 3399 972 3400
rect 1118 3404 1124 3405
rect 1118 3400 1119 3404
rect 1123 3400 1124 3404
rect 1118 3399 1124 3400
rect 1270 3404 1276 3405
rect 1270 3400 1271 3404
rect 1275 3400 1276 3404
rect 2008 3402 2010 3429
rect 2046 3428 2052 3429
rect 2486 3417 2492 3418
rect 2046 3416 2052 3417
rect 2046 3412 2047 3416
rect 2051 3412 2052 3416
rect 2486 3413 2487 3417
rect 2491 3413 2492 3417
rect 2486 3412 2492 3413
rect 2046 3411 2052 3412
rect 1270 3399 1276 3400
rect 2006 3401 2012 3402
rect 2006 3397 2007 3401
rect 2011 3397 2012 3401
rect 2006 3396 2012 3397
rect 458 3395 464 3396
rect 458 3391 459 3395
rect 463 3391 464 3395
rect 458 3390 464 3391
rect 602 3395 608 3396
rect 602 3391 603 3395
rect 607 3391 608 3395
rect 602 3390 608 3391
rect 610 3395 616 3396
rect 610 3391 611 3395
rect 615 3391 616 3395
rect 610 3390 616 3391
rect 882 3395 888 3396
rect 882 3391 883 3395
rect 887 3391 888 3395
rect 882 3390 888 3391
rect 902 3395 908 3396
rect 902 3391 903 3395
rect 907 3391 908 3395
rect 902 3390 908 3391
rect 1194 3395 1200 3396
rect 1194 3391 1195 3395
rect 1199 3391 1200 3395
rect 1194 3390 1200 3391
rect 1234 3395 1240 3396
rect 1234 3391 1235 3395
rect 1239 3391 1240 3395
rect 1234 3390 1240 3391
rect 382 3385 388 3386
rect 382 3381 383 3385
rect 387 3381 388 3385
rect 382 3380 388 3381
rect 362 3367 368 3368
rect 362 3363 363 3367
rect 367 3363 368 3367
rect 362 3362 368 3363
rect 384 3351 386 3380
rect 460 3368 462 3390
rect 526 3385 532 3386
rect 526 3381 527 3385
rect 531 3381 532 3385
rect 526 3380 532 3381
rect 458 3367 464 3368
rect 458 3363 459 3367
rect 463 3363 464 3367
rect 458 3362 464 3363
rect 528 3351 530 3380
rect 604 3368 606 3390
rect 612 3376 614 3390
rect 670 3385 676 3386
rect 670 3381 671 3385
rect 675 3381 676 3385
rect 670 3380 676 3381
rect 814 3385 820 3386
rect 814 3381 815 3385
rect 819 3381 820 3385
rect 814 3380 820 3381
rect 610 3375 616 3376
rect 610 3371 611 3375
rect 615 3371 616 3375
rect 610 3370 616 3371
rect 602 3367 608 3368
rect 602 3363 603 3367
rect 607 3363 608 3367
rect 602 3362 608 3363
rect 672 3351 674 3380
rect 816 3351 818 3380
rect 904 3368 906 3390
rect 966 3385 972 3386
rect 966 3381 967 3385
rect 971 3381 972 3385
rect 966 3380 972 3381
rect 1118 3385 1124 3386
rect 1118 3381 1119 3385
rect 1123 3381 1124 3385
rect 1118 3380 1124 3381
rect 902 3367 908 3368
rect 902 3363 903 3367
rect 907 3363 908 3367
rect 902 3362 908 3363
rect 968 3351 970 3380
rect 1120 3351 1122 3380
rect 1196 3368 1198 3390
rect 1236 3376 1238 3390
rect 1270 3385 1276 3386
rect 1270 3381 1271 3385
rect 1275 3381 1276 3385
rect 1270 3380 1276 3381
rect 2006 3384 2012 3385
rect 2006 3380 2007 3384
rect 2011 3380 2012 3384
rect 2048 3383 2050 3411
rect 2488 3383 2490 3412
rect 2548 3400 2550 3494
rect 2574 3492 2575 3496
rect 2579 3492 2580 3496
rect 2574 3491 2580 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2576 3467 2578 3491
rect 2672 3467 2674 3491
rect 2575 3466 2579 3467
rect 2575 3461 2579 3462
rect 2583 3466 2587 3467
rect 2583 3461 2587 3462
rect 2671 3466 2675 3467
rect 2671 3461 2675 3462
rect 2679 3466 2683 3467
rect 2679 3461 2683 3462
rect 2584 3437 2586 3461
rect 2680 3437 2682 3461
rect 2582 3436 2588 3437
rect 2582 3432 2583 3436
rect 2587 3432 2588 3436
rect 2582 3431 2588 3432
rect 2678 3436 2684 3437
rect 2678 3432 2679 3436
rect 2683 3432 2684 3436
rect 2678 3431 2684 3432
rect 2748 3428 2750 3497
rect 2766 3496 2772 3497
rect 2766 3492 2767 3496
rect 2771 3492 2772 3496
rect 2863 3495 2867 3496
rect 2870 3496 2876 3497
rect 2766 3491 2772 3492
rect 2870 3492 2871 3496
rect 2875 3492 2876 3496
rect 2870 3491 2876 3492
rect 2982 3496 2988 3497
rect 2982 3492 2983 3496
rect 2987 3492 2988 3496
rect 2982 3491 2988 3492
rect 2768 3467 2770 3491
rect 2872 3467 2874 3491
rect 2984 3467 2986 3491
rect 2767 3466 2771 3467
rect 2767 3461 2771 3462
rect 2783 3466 2787 3467
rect 2783 3461 2787 3462
rect 2871 3466 2875 3467
rect 2871 3461 2875 3462
rect 2895 3466 2899 3467
rect 2895 3461 2899 3462
rect 2983 3466 2987 3467
rect 2983 3461 2987 3462
rect 3015 3466 3019 3467
rect 3015 3461 3019 3462
rect 2784 3437 2786 3461
rect 2896 3437 2898 3461
rect 3016 3437 3018 3461
rect 2782 3436 2788 3437
rect 2782 3432 2783 3436
rect 2787 3432 2788 3436
rect 2782 3431 2788 3432
rect 2894 3436 2900 3437
rect 2894 3432 2895 3436
rect 2899 3432 2900 3436
rect 2894 3431 2900 3432
rect 3014 3436 3020 3437
rect 3014 3432 3015 3436
rect 3019 3432 3020 3436
rect 3014 3431 3020 3432
rect 2562 3427 2568 3428
rect 2562 3423 2563 3427
rect 2567 3423 2568 3427
rect 2562 3422 2568 3423
rect 2658 3427 2664 3428
rect 2658 3423 2659 3427
rect 2663 3423 2664 3427
rect 2658 3422 2664 3423
rect 2746 3427 2752 3428
rect 2746 3423 2747 3427
rect 2751 3423 2752 3427
rect 2746 3422 2752 3423
rect 2886 3427 2892 3428
rect 2886 3423 2887 3427
rect 2891 3423 2892 3427
rect 2886 3422 2892 3423
rect 2990 3427 2996 3428
rect 2990 3423 2991 3427
rect 2995 3423 2996 3427
rect 2990 3422 2996 3423
rect 2564 3400 2566 3422
rect 2582 3417 2588 3418
rect 2582 3413 2583 3417
rect 2587 3413 2588 3417
rect 2582 3412 2588 3413
rect 2546 3399 2552 3400
rect 2546 3395 2547 3399
rect 2551 3395 2552 3399
rect 2546 3394 2552 3395
rect 2562 3399 2568 3400
rect 2562 3395 2563 3399
rect 2567 3395 2568 3399
rect 2562 3394 2568 3395
rect 2584 3383 2586 3412
rect 2660 3400 2662 3422
rect 2678 3417 2684 3418
rect 2678 3413 2679 3417
rect 2683 3413 2684 3417
rect 2678 3412 2684 3413
rect 2782 3417 2788 3418
rect 2782 3413 2783 3417
rect 2787 3413 2788 3417
rect 2782 3412 2788 3413
rect 2658 3399 2664 3400
rect 2658 3395 2659 3399
rect 2663 3395 2664 3399
rect 2658 3394 2664 3395
rect 2680 3383 2682 3412
rect 2784 3383 2786 3412
rect 2888 3400 2890 3422
rect 2894 3417 2900 3418
rect 2894 3413 2895 3417
rect 2899 3413 2900 3417
rect 2894 3412 2900 3413
rect 2886 3399 2892 3400
rect 2886 3395 2887 3399
rect 2891 3395 2892 3399
rect 2886 3394 2892 3395
rect 2896 3383 2898 3412
rect 2992 3400 2994 3422
rect 3014 3417 3020 3418
rect 3014 3413 3015 3417
rect 3019 3413 3020 3417
rect 3014 3412 3020 3413
rect 2990 3399 2996 3400
rect 2990 3395 2991 3399
rect 2995 3395 2996 3399
rect 2990 3394 2996 3395
rect 3016 3383 3018 3412
rect 3068 3400 3070 3502
rect 3102 3496 3108 3497
rect 3102 3492 3103 3496
rect 3107 3492 3108 3496
rect 3102 3491 3108 3492
rect 3222 3496 3228 3497
rect 3222 3492 3223 3496
rect 3227 3492 3228 3496
rect 3222 3491 3228 3492
rect 3104 3467 3106 3491
rect 3224 3467 3226 3491
rect 3103 3466 3107 3467
rect 3103 3461 3107 3462
rect 3143 3466 3147 3467
rect 3143 3461 3147 3462
rect 3223 3466 3227 3467
rect 3223 3461 3227 3462
rect 3144 3437 3146 3461
rect 3142 3436 3148 3437
rect 3142 3432 3143 3436
rect 3147 3432 3148 3436
rect 3142 3431 3148 3432
rect 3232 3428 3234 3530
rect 3352 3516 3354 3537
rect 3396 3536 3398 3590
rect 3566 3585 3572 3586
rect 3566 3581 3567 3585
rect 3571 3581 3572 3585
rect 3566 3580 3572 3581
rect 3568 3543 3570 3580
rect 3596 3568 3598 3670
rect 3726 3668 3732 3669
rect 3726 3664 3727 3668
rect 3731 3664 3732 3668
rect 3942 3667 3943 3671
rect 3947 3667 3948 3671
rect 3942 3666 3948 3667
rect 3726 3663 3732 3664
rect 3728 3635 3730 3663
rect 3944 3635 3946 3666
rect 3727 3634 3731 3635
rect 3727 3629 3731 3630
rect 3943 3634 3947 3635
rect 3943 3629 3947 3630
rect 3944 3602 3946 3629
rect 3942 3601 3948 3602
rect 3942 3597 3943 3601
rect 3947 3597 3948 3601
rect 3942 3596 3948 3597
rect 3942 3584 3948 3585
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 3942 3579 3948 3580
rect 3594 3567 3600 3568
rect 3594 3563 3595 3567
rect 3599 3563 3600 3567
rect 3594 3562 3600 3563
rect 3944 3543 3946 3579
rect 3487 3542 3491 3543
rect 3487 3537 3491 3538
rect 3567 3542 3571 3543
rect 3567 3537 3571 3538
rect 3943 3542 3947 3543
rect 3943 3537 3947 3538
rect 3390 3535 3398 3536
rect 3390 3531 3391 3535
rect 3395 3532 3398 3535
rect 3426 3535 3432 3536
rect 3395 3531 3396 3532
rect 3390 3530 3396 3531
rect 3426 3531 3427 3535
rect 3431 3531 3432 3535
rect 3426 3530 3432 3531
rect 3350 3515 3356 3516
rect 3350 3511 3351 3515
rect 3355 3511 3356 3515
rect 3350 3510 3356 3511
rect 3428 3508 3430 3530
rect 3488 3516 3490 3537
rect 3944 3517 3946 3537
rect 3942 3516 3948 3517
rect 3486 3515 3492 3516
rect 3486 3511 3487 3515
rect 3491 3511 3492 3515
rect 3942 3512 3943 3516
rect 3947 3512 3948 3516
rect 3942 3511 3948 3512
rect 3486 3510 3492 3511
rect 3426 3507 3432 3508
rect 3426 3503 3427 3507
rect 3431 3503 3432 3507
rect 3426 3502 3432 3503
rect 3466 3507 3472 3508
rect 3466 3503 3467 3507
rect 3471 3503 3472 3507
rect 3466 3502 3472 3503
rect 3350 3496 3356 3497
rect 3350 3492 3351 3496
rect 3355 3492 3356 3496
rect 3350 3491 3356 3492
rect 3352 3467 3354 3491
rect 3271 3466 3275 3467
rect 3271 3461 3275 3462
rect 3351 3466 3355 3467
rect 3351 3461 3355 3462
rect 3407 3466 3411 3467
rect 3407 3461 3411 3462
rect 3272 3437 3274 3461
rect 3408 3437 3410 3461
rect 3270 3436 3276 3437
rect 3270 3432 3271 3436
rect 3275 3432 3276 3436
rect 3270 3431 3276 3432
rect 3406 3436 3412 3437
rect 3406 3432 3407 3436
rect 3411 3432 3412 3436
rect 3406 3431 3412 3432
rect 3230 3427 3236 3428
rect 3230 3423 3231 3427
rect 3235 3423 3236 3427
rect 3230 3422 3236 3423
rect 3338 3427 3344 3428
rect 3338 3423 3339 3427
rect 3343 3423 3344 3427
rect 3338 3422 3344 3423
rect 3378 3427 3384 3428
rect 3378 3423 3379 3427
rect 3383 3423 3384 3427
rect 3378 3422 3384 3423
rect 3142 3417 3148 3418
rect 3142 3413 3143 3417
rect 3147 3413 3148 3417
rect 3142 3412 3148 3413
rect 3270 3417 3276 3418
rect 3270 3413 3271 3417
rect 3275 3413 3276 3417
rect 3270 3412 3276 3413
rect 3066 3399 3072 3400
rect 3066 3395 3067 3399
rect 3071 3395 3072 3399
rect 3066 3394 3072 3395
rect 3098 3395 3104 3396
rect 3098 3391 3099 3395
rect 3103 3391 3104 3395
rect 3098 3390 3104 3391
rect 1234 3375 1240 3376
rect 1234 3371 1235 3375
rect 1239 3371 1240 3375
rect 1234 3370 1240 3371
rect 1194 3367 1200 3368
rect 1158 3363 1164 3364
rect 1158 3359 1159 3363
rect 1163 3359 1164 3363
rect 1194 3363 1195 3367
rect 1199 3363 1200 3367
rect 1194 3362 1200 3363
rect 1158 3358 1164 3359
rect 1160 3355 1162 3358
rect 1160 3353 1166 3355
rect 247 3350 251 3351
rect 247 3345 251 3346
rect 263 3350 267 3351
rect 263 3345 267 3346
rect 383 3350 387 3351
rect 383 3345 387 3346
rect 431 3350 435 3351
rect 431 3345 435 3346
rect 527 3350 531 3351
rect 527 3345 531 3346
rect 599 3350 603 3351
rect 599 3345 603 3346
rect 671 3350 675 3351
rect 671 3345 675 3346
rect 767 3350 771 3351
rect 767 3345 771 3346
rect 815 3350 819 3351
rect 815 3345 819 3346
rect 927 3350 931 3351
rect 927 3345 931 3346
rect 967 3350 971 3351
rect 967 3345 971 3346
rect 1087 3350 1091 3351
rect 1087 3345 1091 3346
rect 1119 3350 1123 3351
rect 1119 3345 1123 3346
rect 202 3343 208 3344
rect 202 3339 203 3343
rect 207 3339 208 3343
rect 202 3338 208 3339
rect 210 3343 216 3344
rect 210 3339 211 3343
rect 215 3339 216 3343
rect 210 3338 216 3339
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 134 3323 140 3324
rect 134 3319 135 3323
rect 139 3319 140 3323
rect 134 3318 140 3319
rect 212 3316 214 3338
rect 264 3324 266 3345
rect 338 3343 344 3344
rect 338 3339 339 3343
rect 343 3339 344 3343
rect 338 3338 344 3339
rect 262 3323 268 3324
rect 262 3319 263 3323
rect 267 3319 268 3323
rect 262 3318 268 3319
rect 340 3316 342 3338
rect 432 3324 434 3345
rect 506 3343 512 3344
rect 506 3339 507 3343
rect 511 3339 512 3343
rect 506 3338 512 3339
rect 430 3323 436 3324
rect 430 3319 431 3323
rect 435 3319 436 3323
rect 430 3318 436 3319
rect 508 3316 510 3338
rect 600 3324 602 3345
rect 768 3324 770 3345
rect 928 3324 930 3345
rect 1002 3343 1008 3344
rect 1002 3339 1003 3343
rect 1007 3339 1008 3343
rect 1002 3338 1008 3339
rect 598 3323 604 3324
rect 598 3319 599 3323
rect 603 3319 604 3323
rect 598 3318 604 3319
rect 766 3323 772 3324
rect 766 3319 767 3323
rect 771 3319 772 3323
rect 766 3318 772 3319
rect 926 3323 932 3324
rect 926 3319 927 3323
rect 931 3319 932 3323
rect 926 3318 932 3319
rect 1004 3316 1006 3338
rect 1088 3324 1090 3345
rect 1086 3323 1092 3324
rect 1086 3319 1087 3323
rect 1091 3319 1092 3323
rect 1086 3318 1092 3319
rect 1164 3316 1166 3353
rect 1272 3351 1274 3380
rect 2006 3379 2012 3380
rect 2047 3382 2051 3383
rect 2008 3351 2010 3379
rect 2047 3377 2051 3378
rect 2351 3382 2355 3383
rect 2351 3377 2355 3378
rect 2479 3382 2483 3383
rect 2479 3377 2483 3378
rect 2487 3382 2491 3383
rect 2487 3377 2491 3378
rect 2583 3382 2587 3383
rect 2583 3377 2587 3378
rect 2615 3382 2619 3383
rect 2615 3377 2619 3378
rect 2679 3382 2683 3383
rect 2679 3377 2683 3378
rect 2751 3382 2755 3383
rect 2751 3377 2755 3378
rect 2783 3382 2787 3383
rect 2783 3377 2787 3378
rect 2887 3382 2891 3383
rect 2887 3377 2891 3378
rect 2895 3382 2899 3383
rect 2895 3377 2899 3378
rect 3015 3382 3019 3383
rect 3015 3377 3019 3378
rect 3023 3382 3027 3383
rect 3023 3377 3027 3378
rect 2048 3357 2050 3377
rect 2046 3356 2052 3357
rect 2352 3356 2354 3377
rect 2426 3375 2432 3376
rect 2426 3371 2427 3375
rect 2431 3371 2432 3375
rect 2426 3370 2432 3371
rect 2046 3352 2047 3356
rect 2051 3352 2052 3356
rect 2046 3351 2052 3352
rect 2350 3355 2356 3356
rect 2350 3351 2351 3355
rect 2355 3351 2356 3355
rect 1239 3350 1243 3351
rect 1239 3345 1243 3346
rect 1271 3350 1275 3351
rect 1271 3345 1275 3346
rect 1391 3350 1395 3351
rect 1391 3345 1395 3346
rect 1551 3350 1555 3351
rect 1551 3345 1555 3346
rect 2007 3350 2011 3351
rect 2350 3350 2356 3351
rect 2428 3348 2430 3370
rect 2480 3356 2482 3377
rect 2554 3375 2560 3376
rect 2554 3371 2555 3375
rect 2559 3371 2560 3375
rect 2554 3370 2560 3371
rect 2478 3355 2484 3356
rect 2478 3351 2479 3355
rect 2483 3351 2484 3355
rect 2478 3350 2484 3351
rect 2556 3348 2558 3370
rect 2616 3356 2618 3377
rect 2718 3367 2724 3368
rect 2718 3363 2719 3367
rect 2723 3363 2724 3367
rect 2718 3362 2724 3363
rect 2614 3355 2620 3356
rect 2614 3351 2615 3355
rect 2619 3351 2620 3355
rect 2614 3350 2620 3351
rect 2720 3348 2722 3362
rect 2752 3356 2754 3377
rect 2850 3375 2856 3376
rect 2850 3371 2851 3375
rect 2855 3371 2856 3375
rect 2850 3370 2856 3371
rect 2750 3355 2756 3356
rect 2750 3351 2751 3355
rect 2755 3351 2756 3355
rect 2750 3350 2756 3351
rect 2007 3345 2011 3346
rect 2426 3347 2432 3348
rect 1218 3335 1224 3336
rect 1218 3331 1219 3335
rect 1223 3331 1224 3335
rect 1218 3330 1224 3331
rect 1220 3316 1222 3330
rect 1240 3324 1242 3345
rect 1322 3343 1328 3344
rect 1322 3339 1323 3343
rect 1327 3339 1328 3343
rect 1322 3338 1328 3339
rect 1238 3323 1244 3324
rect 1238 3319 1239 3323
rect 1243 3319 1244 3323
rect 1238 3318 1244 3319
rect 1324 3316 1326 3338
rect 1392 3324 1394 3345
rect 1474 3343 1480 3344
rect 1474 3339 1475 3343
rect 1479 3339 1480 3343
rect 1474 3338 1480 3339
rect 1390 3323 1396 3324
rect 1390 3319 1391 3323
rect 1395 3319 1396 3323
rect 1390 3318 1396 3319
rect 1476 3316 1478 3338
rect 1552 3324 1554 3345
rect 1562 3343 1568 3344
rect 1562 3339 1563 3343
rect 1567 3339 1568 3343
rect 1562 3338 1568 3339
rect 1550 3323 1556 3324
rect 1550 3319 1551 3323
rect 1555 3319 1556 3323
rect 1550 3318 1556 3319
rect 210 3315 216 3316
rect 210 3311 211 3315
rect 215 3311 216 3315
rect 210 3310 216 3311
rect 338 3315 344 3316
rect 338 3311 339 3315
rect 343 3311 344 3315
rect 338 3310 344 3311
rect 506 3315 512 3316
rect 506 3311 507 3315
rect 511 3311 512 3315
rect 506 3310 512 3311
rect 738 3315 744 3316
rect 738 3311 739 3315
rect 743 3311 744 3315
rect 738 3310 744 3311
rect 1002 3315 1008 3316
rect 1002 3311 1003 3315
rect 1007 3311 1008 3315
rect 1002 3310 1008 3311
rect 1162 3315 1168 3316
rect 1162 3311 1163 3315
rect 1167 3311 1168 3315
rect 1162 3310 1168 3311
rect 1218 3315 1224 3316
rect 1218 3311 1219 3315
rect 1223 3311 1224 3315
rect 1218 3310 1224 3311
rect 1322 3315 1328 3316
rect 1322 3311 1323 3315
rect 1327 3311 1328 3315
rect 1322 3310 1328 3311
rect 1474 3315 1480 3316
rect 1474 3311 1475 3315
rect 1479 3311 1480 3315
rect 1474 3310 1480 3311
rect 110 3307 116 3308
rect 110 3303 111 3307
rect 115 3303 116 3307
rect 110 3302 116 3303
rect 134 3304 140 3305
rect 112 3267 114 3302
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 262 3304 268 3305
rect 262 3300 263 3304
rect 267 3300 268 3304
rect 262 3299 268 3300
rect 430 3304 436 3305
rect 430 3300 431 3304
rect 435 3300 436 3304
rect 430 3299 436 3300
rect 598 3304 604 3305
rect 598 3300 599 3304
rect 603 3300 604 3304
rect 598 3299 604 3300
rect 136 3267 138 3299
rect 264 3267 266 3299
rect 432 3267 434 3299
rect 600 3267 602 3299
rect 111 3266 115 3267
rect 111 3261 115 3262
rect 135 3266 139 3267
rect 135 3261 139 3262
rect 143 3266 147 3267
rect 143 3261 147 3262
rect 263 3266 267 3267
rect 263 3261 267 3262
rect 295 3266 299 3267
rect 295 3261 299 3262
rect 431 3266 435 3267
rect 431 3261 435 3262
rect 455 3266 459 3267
rect 455 3261 459 3262
rect 599 3266 603 3267
rect 599 3261 603 3262
rect 623 3266 627 3267
rect 623 3261 627 3262
rect 112 3234 114 3261
rect 144 3237 146 3261
rect 296 3237 298 3261
rect 456 3237 458 3261
rect 624 3237 626 3261
rect 142 3236 148 3237
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 142 3232 143 3236
rect 147 3232 148 3236
rect 142 3231 148 3232
rect 294 3236 300 3237
rect 294 3232 295 3236
rect 299 3232 300 3236
rect 294 3231 300 3232
rect 454 3236 460 3237
rect 454 3232 455 3236
rect 459 3232 460 3236
rect 454 3231 460 3232
rect 622 3236 628 3237
rect 622 3232 623 3236
rect 627 3232 628 3236
rect 622 3231 628 3232
rect 110 3228 116 3229
rect 218 3227 224 3228
rect 218 3223 219 3227
rect 223 3223 224 3227
rect 218 3222 224 3223
rect 370 3227 376 3228
rect 370 3223 371 3227
rect 375 3223 376 3227
rect 370 3222 376 3223
rect 530 3227 536 3228
rect 530 3223 531 3227
rect 535 3223 536 3227
rect 530 3222 536 3223
rect 698 3227 704 3228
rect 698 3223 699 3227
rect 703 3223 704 3227
rect 698 3222 704 3223
rect 142 3217 148 3218
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 142 3213 143 3217
rect 147 3213 148 3217
rect 142 3212 148 3213
rect 110 3211 116 3212
rect 112 3191 114 3211
rect 144 3191 146 3212
rect 183 3204 187 3205
rect 220 3200 222 3222
rect 294 3217 300 3218
rect 294 3213 295 3217
rect 299 3213 300 3217
rect 294 3212 300 3213
rect 182 3199 188 3200
rect 182 3195 183 3199
rect 187 3195 188 3199
rect 182 3194 188 3195
rect 218 3199 224 3200
rect 218 3195 219 3199
rect 223 3195 224 3199
rect 218 3194 224 3195
rect 296 3191 298 3212
rect 372 3200 374 3222
rect 454 3217 460 3218
rect 454 3213 455 3217
rect 459 3213 460 3217
rect 454 3212 460 3213
rect 370 3199 376 3200
rect 370 3195 371 3199
rect 375 3195 376 3199
rect 370 3194 376 3195
rect 456 3191 458 3212
rect 532 3200 534 3222
rect 622 3217 628 3218
rect 622 3213 623 3217
rect 627 3213 628 3217
rect 622 3212 628 3213
rect 530 3199 536 3200
rect 530 3195 531 3199
rect 535 3195 536 3199
rect 530 3194 536 3195
rect 624 3191 626 3212
rect 700 3200 702 3222
rect 740 3205 742 3310
rect 766 3304 772 3305
rect 766 3300 767 3304
rect 771 3300 772 3304
rect 766 3299 772 3300
rect 926 3304 932 3305
rect 926 3300 927 3304
rect 931 3300 932 3304
rect 926 3299 932 3300
rect 1086 3304 1092 3305
rect 1086 3300 1087 3304
rect 1091 3300 1092 3304
rect 1086 3299 1092 3300
rect 1238 3304 1244 3305
rect 1238 3300 1239 3304
rect 1243 3300 1244 3304
rect 1238 3299 1244 3300
rect 1390 3304 1396 3305
rect 1390 3300 1391 3304
rect 1395 3300 1396 3304
rect 1390 3299 1396 3300
rect 1550 3304 1556 3305
rect 1550 3300 1551 3304
rect 1555 3300 1556 3304
rect 1550 3299 1556 3300
rect 768 3267 770 3299
rect 928 3267 930 3299
rect 1088 3267 1090 3299
rect 1240 3267 1242 3299
rect 1392 3267 1394 3299
rect 1552 3267 1554 3299
rect 767 3266 771 3267
rect 767 3261 771 3262
rect 791 3266 795 3267
rect 791 3261 795 3262
rect 927 3266 931 3267
rect 927 3261 931 3262
rect 959 3266 963 3267
rect 959 3261 963 3262
rect 1087 3266 1091 3267
rect 1087 3261 1091 3262
rect 1127 3266 1131 3267
rect 1127 3261 1131 3262
rect 1239 3266 1243 3267
rect 1239 3261 1243 3262
rect 1303 3266 1307 3267
rect 1303 3261 1307 3262
rect 1391 3266 1395 3267
rect 1391 3261 1395 3262
rect 1479 3266 1483 3267
rect 1479 3261 1483 3262
rect 1551 3266 1555 3267
rect 1551 3261 1555 3262
rect 792 3237 794 3261
rect 960 3237 962 3261
rect 1128 3237 1130 3261
rect 1304 3237 1306 3261
rect 1480 3237 1482 3261
rect 790 3236 796 3237
rect 790 3232 791 3236
rect 795 3232 796 3236
rect 790 3231 796 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 958 3231 964 3232
rect 1126 3236 1132 3237
rect 1126 3232 1127 3236
rect 1131 3232 1132 3236
rect 1126 3231 1132 3232
rect 1302 3236 1308 3237
rect 1302 3232 1303 3236
rect 1307 3232 1308 3236
rect 1302 3231 1308 3232
rect 1478 3236 1484 3237
rect 1478 3232 1479 3236
rect 1483 3232 1484 3236
rect 1478 3231 1484 3232
rect 1564 3228 1566 3338
rect 2008 3325 2010 3345
rect 2426 3343 2427 3347
rect 2431 3343 2432 3347
rect 2426 3342 2432 3343
rect 2554 3347 2560 3348
rect 2554 3343 2555 3347
rect 2559 3343 2560 3347
rect 2554 3342 2560 3343
rect 2718 3347 2724 3348
rect 2718 3343 2719 3347
rect 2723 3343 2724 3347
rect 2718 3342 2724 3343
rect 2046 3339 2052 3340
rect 2046 3335 2047 3339
rect 2051 3335 2052 3339
rect 2682 3339 2688 3340
rect 2046 3334 2052 3335
rect 2350 3336 2356 3337
rect 2006 3324 2012 3325
rect 2006 3320 2007 3324
rect 2011 3320 2012 3324
rect 2006 3319 2012 3320
rect 2006 3307 2012 3308
rect 2006 3303 2007 3307
rect 2011 3303 2012 3307
rect 2048 3303 2050 3334
rect 2350 3332 2351 3336
rect 2355 3332 2356 3336
rect 2350 3331 2356 3332
rect 2478 3336 2484 3337
rect 2478 3332 2479 3336
rect 2483 3332 2484 3336
rect 2478 3331 2484 3332
rect 2614 3336 2620 3337
rect 2614 3332 2615 3336
rect 2619 3332 2620 3336
rect 2682 3335 2683 3339
rect 2687 3335 2688 3339
rect 2682 3334 2688 3335
rect 2750 3336 2756 3337
rect 2614 3331 2620 3332
rect 2352 3303 2354 3331
rect 2480 3303 2482 3331
rect 2616 3303 2618 3331
rect 2006 3302 2012 3303
rect 2047 3302 2051 3303
rect 2008 3267 2010 3302
rect 2047 3297 2051 3298
rect 2127 3302 2131 3303
rect 2127 3297 2131 3298
rect 2295 3302 2299 3303
rect 2295 3297 2299 3298
rect 2351 3302 2355 3303
rect 2351 3297 2355 3298
rect 2455 3302 2459 3303
rect 2455 3297 2459 3298
rect 2479 3302 2483 3303
rect 2479 3297 2483 3298
rect 2615 3302 2619 3303
rect 2615 3297 2619 3298
rect 2048 3270 2050 3297
rect 2128 3273 2130 3297
rect 2296 3273 2298 3297
rect 2456 3273 2458 3297
rect 2616 3273 2618 3297
rect 2126 3272 2132 3273
rect 2046 3269 2052 3270
rect 2007 3266 2011 3267
rect 2046 3265 2047 3269
rect 2051 3265 2052 3269
rect 2126 3268 2127 3272
rect 2131 3268 2132 3272
rect 2126 3267 2132 3268
rect 2294 3272 2300 3273
rect 2294 3268 2295 3272
rect 2299 3268 2300 3272
rect 2294 3267 2300 3268
rect 2454 3272 2460 3273
rect 2454 3268 2455 3272
rect 2459 3268 2460 3272
rect 2454 3267 2460 3268
rect 2614 3272 2620 3273
rect 2614 3268 2615 3272
rect 2619 3268 2620 3272
rect 2614 3267 2620 3268
rect 2046 3264 2052 3265
rect 2007 3261 2011 3262
rect 2214 3263 2220 3264
rect 2008 3234 2010 3261
rect 2214 3259 2215 3263
rect 2219 3259 2220 3263
rect 2214 3258 2220 3259
rect 2222 3263 2228 3264
rect 2222 3259 2223 3263
rect 2227 3259 2228 3263
rect 2222 3258 2228 3259
rect 2398 3263 2404 3264
rect 2398 3259 2399 3263
rect 2403 3259 2404 3263
rect 2398 3258 2404 3259
rect 2126 3253 2132 3254
rect 2046 3252 2052 3253
rect 2046 3248 2047 3252
rect 2051 3248 2052 3252
rect 2126 3249 2127 3253
rect 2131 3249 2132 3253
rect 2126 3248 2132 3249
rect 2046 3247 2052 3248
rect 2006 3233 2012 3234
rect 2006 3229 2007 3233
rect 2011 3229 2012 3233
rect 2006 3228 2012 3229
rect 1034 3227 1040 3228
rect 1034 3223 1035 3227
rect 1039 3223 1040 3227
rect 1034 3222 1040 3223
rect 1202 3227 1208 3228
rect 1202 3223 1203 3227
rect 1207 3223 1208 3227
rect 1202 3222 1208 3223
rect 1378 3227 1384 3228
rect 1378 3223 1379 3227
rect 1383 3223 1384 3227
rect 1378 3222 1384 3223
rect 1562 3227 1568 3228
rect 2048 3227 2050 3247
rect 2128 3227 2130 3248
rect 1562 3223 1563 3227
rect 1567 3223 1568 3227
rect 1562 3222 1568 3223
rect 2047 3226 2051 3227
rect 790 3217 796 3218
rect 790 3213 791 3217
rect 795 3213 796 3217
rect 790 3212 796 3213
rect 958 3217 964 3218
rect 958 3213 959 3217
rect 963 3213 964 3217
rect 958 3212 964 3213
rect 739 3204 743 3205
rect 698 3199 704 3200
rect 739 3199 743 3200
rect 698 3195 699 3199
rect 703 3195 704 3199
rect 698 3194 704 3195
rect 792 3191 794 3212
rect 960 3191 962 3212
rect 1036 3204 1038 3222
rect 1126 3217 1132 3218
rect 1126 3213 1127 3217
rect 1131 3213 1132 3217
rect 1126 3212 1132 3213
rect 1034 3203 1040 3204
rect 1034 3199 1035 3203
rect 1039 3199 1040 3203
rect 1034 3198 1040 3199
rect 1128 3191 1130 3212
rect 1204 3200 1206 3222
rect 1302 3217 1308 3218
rect 1302 3213 1303 3217
rect 1307 3213 1308 3217
rect 1302 3212 1308 3213
rect 1202 3199 1208 3200
rect 1202 3195 1203 3199
rect 1207 3195 1208 3199
rect 1202 3194 1208 3195
rect 1304 3191 1306 3212
rect 1380 3200 1382 3222
rect 2047 3221 2051 3222
rect 2071 3226 2075 3227
rect 2071 3221 2075 3222
rect 2127 3226 2131 3227
rect 2127 3221 2131 3222
rect 2207 3226 2211 3227
rect 2207 3221 2211 3222
rect 1478 3217 1484 3218
rect 1478 3213 1479 3217
rect 1483 3213 1484 3217
rect 1478 3212 1484 3213
rect 2006 3216 2012 3217
rect 2006 3212 2007 3216
rect 2011 3212 2012 3216
rect 1378 3199 1384 3200
rect 1378 3195 1379 3199
rect 1383 3195 1384 3199
rect 1378 3194 1384 3195
rect 1480 3191 1482 3212
rect 2006 3211 2012 3212
rect 1638 3191 1644 3192
rect 2008 3191 2010 3211
rect 2048 3201 2050 3221
rect 2046 3200 2052 3201
rect 2072 3200 2074 3221
rect 2208 3200 2210 3221
rect 2216 3220 2218 3258
rect 2224 3236 2226 3258
rect 2294 3253 2300 3254
rect 2294 3249 2295 3253
rect 2299 3249 2300 3253
rect 2294 3248 2300 3249
rect 2222 3235 2228 3236
rect 2222 3231 2223 3235
rect 2227 3231 2228 3235
rect 2222 3230 2228 3231
rect 2296 3227 2298 3248
rect 2400 3236 2402 3258
rect 2454 3253 2460 3254
rect 2454 3249 2455 3253
rect 2459 3249 2460 3253
rect 2454 3248 2460 3249
rect 2614 3253 2620 3254
rect 2614 3249 2615 3253
rect 2619 3249 2620 3253
rect 2614 3248 2620 3249
rect 2398 3235 2404 3236
rect 2398 3231 2399 3235
rect 2403 3231 2404 3235
rect 2398 3230 2404 3231
rect 2456 3227 2458 3248
rect 2616 3227 2618 3248
rect 2684 3236 2686 3334
rect 2750 3332 2751 3336
rect 2755 3332 2756 3336
rect 2750 3331 2756 3332
rect 2752 3303 2754 3331
rect 2751 3302 2755 3303
rect 2751 3297 2755 3298
rect 2775 3302 2779 3303
rect 2775 3297 2779 3298
rect 2776 3273 2778 3297
rect 2774 3272 2780 3273
rect 2774 3268 2775 3272
rect 2779 3268 2780 3272
rect 2774 3267 2780 3268
rect 2852 3264 2854 3370
rect 2888 3356 2890 3377
rect 2962 3375 2968 3376
rect 2962 3371 2963 3375
rect 2967 3371 2968 3375
rect 2962 3370 2968 3371
rect 2886 3355 2892 3356
rect 2886 3351 2887 3355
rect 2891 3351 2892 3355
rect 2886 3350 2892 3351
rect 2964 3348 2966 3370
rect 3024 3356 3026 3377
rect 3022 3355 3028 3356
rect 3022 3351 3023 3355
rect 3027 3351 3028 3355
rect 3022 3350 3028 3351
rect 3100 3348 3102 3390
rect 3144 3383 3146 3412
rect 3272 3383 3274 3412
rect 3143 3382 3147 3383
rect 3143 3377 3147 3378
rect 3159 3382 3163 3383
rect 3159 3377 3163 3378
rect 3271 3382 3275 3383
rect 3271 3377 3275 3378
rect 3303 3382 3307 3383
rect 3303 3377 3307 3378
rect 3160 3356 3162 3377
rect 3242 3375 3248 3376
rect 3242 3371 3243 3375
rect 3247 3371 3248 3375
rect 3242 3370 3248 3371
rect 3158 3355 3164 3356
rect 3158 3351 3159 3355
rect 3163 3351 3164 3355
rect 3158 3350 3164 3351
rect 3244 3348 3246 3370
rect 3304 3356 3306 3377
rect 3340 3376 3342 3422
rect 3380 3400 3382 3422
rect 3406 3417 3412 3418
rect 3406 3413 3407 3417
rect 3411 3413 3412 3417
rect 3406 3412 3412 3413
rect 3378 3399 3384 3400
rect 3378 3395 3379 3399
rect 3383 3395 3384 3399
rect 3378 3394 3384 3395
rect 3408 3383 3410 3412
rect 3468 3400 3470 3502
rect 3942 3499 3948 3500
rect 3486 3496 3492 3497
rect 3486 3492 3487 3496
rect 3491 3492 3492 3496
rect 3942 3495 3943 3499
rect 3947 3495 3948 3499
rect 3942 3494 3948 3495
rect 3486 3491 3492 3492
rect 3488 3467 3490 3491
rect 3944 3467 3946 3494
rect 3487 3466 3491 3467
rect 3487 3461 3491 3462
rect 3943 3466 3947 3467
rect 3943 3461 3947 3462
rect 3944 3434 3946 3461
rect 3942 3433 3948 3434
rect 3942 3429 3943 3433
rect 3947 3429 3948 3433
rect 3942 3428 3948 3429
rect 3942 3416 3948 3417
rect 3942 3412 3943 3416
rect 3947 3412 3948 3416
rect 3942 3411 3948 3412
rect 3466 3399 3472 3400
rect 3466 3395 3467 3399
rect 3471 3395 3472 3399
rect 3466 3394 3472 3395
rect 3944 3383 3946 3411
rect 3407 3382 3411 3383
rect 3407 3377 3411 3378
rect 3943 3382 3947 3383
rect 3943 3377 3947 3378
rect 3338 3375 3344 3376
rect 3338 3371 3339 3375
rect 3343 3371 3344 3375
rect 3338 3370 3344 3371
rect 3944 3357 3946 3377
rect 3942 3356 3948 3357
rect 3302 3355 3308 3356
rect 3302 3351 3303 3355
rect 3307 3351 3308 3355
rect 3942 3352 3943 3356
rect 3947 3352 3948 3356
rect 3942 3351 3948 3352
rect 3302 3350 3308 3351
rect 2962 3347 2968 3348
rect 2962 3343 2963 3347
rect 2967 3343 2968 3347
rect 2962 3342 2968 3343
rect 3098 3347 3104 3348
rect 3098 3343 3099 3347
rect 3103 3343 3104 3347
rect 3242 3347 3248 3348
rect 3098 3342 3104 3343
rect 3234 3343 3240 3344
rect 3234 3339 3235 3343
rect 3239 3339 3240 3343
rect 3242 3343 3243 3347
rect 3247 3343 3248 3347
rect 3242 3342 3248 3343
rect 3234 3338 3240 3339
rect 3942 3339 3948 3340
rect 2886 3336 2892 3337
rect 2886 3332 2887 3336
rect 2891 3332 2892 3336
rect 2886 3331 2892 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3158 3336 3164 3337
rect 3158 3332 3159 3336
rect 3163 3332 3164 3336
rect 3158 3331 3164 3332
rect 2888 3303 2890 3331
rect 3024 3303 3026 3331
rect 3160 3303 3162 3331
rect 2887 3302 2891 3303
rect 2887 3297 2891 3298
rect 2935 3302 2939 3303
rect 2935 3297 2939 3298
rect 3023 3302 3027 3303
rect 3023 3297 3027 3298
rect 3095 3302 3099 3303
rect 3095 3297 3099 3298
rect 3159 3302 3163 3303
rect 3159 3297 3163 3298
rect 2936 3273 2938 3297
rect 3096 3273 3098 3297
rect 2934 3272 2940 3273
rect 2934 3268 2935 3272
rect 2939 3268 2940 3272
rect 2934 3267 2940 3268
rect 3094 3272 3100 3273
rect 3094 3268 3095 3272
rect 3099 3268 3100 3272
rect 3094 3267 3100 3268
rect 2850 3263 2856 3264
rect 2850 3259 2851 3263
rect 2855 3259 2856 3263
rect 2850 3258 2856 3259
rect 3022 3263 3028 3264
rect 3022 3259 3023 3263
rect 3027 3259 3028 3263
rect 3022 3258 3028 3259
rect 3030 3263 3036 3264
rect 3030 3259 3031 3263
rect 3035 3259 3036 3263
rect 3030 3258 3036 3259
rect 3178 3263 3184 3264
rect 3178 3259 3179 3263
rect 3183 3259 3184 3263
rect 3178 3258 3184 3259
rect 2774 3253 2780 3254
rect 2774 3249 2775 3253
rect 2779 3249 2780 3253
rect 2774 3248 2780 3249
rect 2934 3253 2940 3254
rect 2934 3249 2935 3253
rect 2939 3249 2940 3253
rect 2934 3248 2940 3249
rect 2682 3235 2688 3236
rect 2682 3231 2683 3235
rect 2687 3231 2688 3235
rect 2682 3230 2688 3231
rect 2776 3227 2778 3248
rect 2936 3227 2938 3248
rect 2295 3226 2299 3227
rect 2295 3221 2299 3222
rect 2375 3226 2379 3227
rect 2375 3221 2379 3222
rect 2455 3226 2459 3227
rect 2455 3221 2459 3222
rect 2543 3226 2547 3227
rect 2543 3221 2547 3222
rect 2615 3226 2619 3227
rect 2615 3221 2619 3222
rect 2703 3226 2707 3227
rect 2703 3221 2707 3222
rect 2775 3226 2779 3227
rect 2775 3221 2779 3222
rect 2863 3226 2867 3227
rect 2863 3221 2867 3222
rect 2935 3226 2939 3227
rect 2935 3221 2939 3222
rect 3015 3226 3019 3227
rect 3015 3221 3019 3222
rect 2214 3219 2220 3220
rect 2214 3215 2215 3219
rect 2219 3215 2220 3219
rect 2214 3214 2220 3215
rect 2282 3219 2288 3220
rect 2282 3215 2283 3219
rect 2287 3215 2288 3219
rect 2282 3214 2288 3215
rect 2046 3196 2047 3200
rect 2051 3196 2052 3200
rect 2046 3195 2052 3196
rect 2070 3199 2076 3200
rect 2070 3195 2071 3199
rect 2075 3195 2076 3199
rect 2070 3194 2076 3195
rect 2206 3199 2212 3200
rect 2206 3195 2207 3199
rect 2211 3195 2212 3199
rect 2206 3194 2212 3195
rect 2284 3192 2286 3214
rect 2376 3200 2378 3221
rect 2494 3219 2500 3220
rect 2494 3215 2495 3219
rect 2499 3215 2500 3219
rect 2494 3214 2500 3215
rect 2374 3199 2380 3200
rect 2374 3195 2375 3199
rect 2379 3195 2380 3199
rect 2374 3194 2380 3195
rect 2496 3192 2498 3214
rect 2502 3211 2508 3212
rect 2502 3207 2503 3211
rect 2507 3207 2508 3211
rect 2502 3206 2508 3207
rect 2504 3192 2506 3206
rect 2544 3200 2546 3221
rect 2704 3200 2706 3221
rect 2714 3219 2720 3220
rect 2714 3215 2715 3219
rect 2719 3215 2720 3219
rect 2714 3214 2720 3215
rect 2790 3219 2796 3220
rect 2790 3215 2791 3219
rect 2795 3215 2796 3219
rect 2790 3214 2796 3215
rect 2542 3199 2548 3200
rect 2542 3195 2543 3199
rect 2547 3195 2548 3199
rect 2542 3194 2548 3195
rect 2702 3199 2708 3200
rect 2702 3195 2703 3199
rect 2707 3195 2708 3199
rect 2702 3194 2708 3195
rect 2282 3191 2288 3192
rect 111 3190 115 3191
rect 111 3185 115 3186
rect 143 3190 147 3191
rect 143 3185 147 3186
rect 295 3190 299 3191
rect 295 3185 299 3186
rect 431 3190 435 3191
rect 431 3185 435 3186
rect 455 3190 459 3191
rect 455 3185 459 3186
rect 567 3190 571 3191
rect 567 3185 571 3186
rect 623 3190 627 3191
rect 623 3185 627 3186
rect 703 3190 707 3191
rect 703 3185 707 3186
rect 791 3190 795 3191
rect 791 3185 795 3186
rect 855 3190 859 3191
rect 855 3185 859 3186
rect 959 3190 963 3191
rect 959 3185 963 3186
rect 1031 3190 1035 3191
rect 1031 3185 1035 3186
rect 1127 3190 1131 3191
rect 1127 3185 1131 3186
rect 1231 3190 1235 3191
rect 1231 3185 1235 3186
rect 1303 3190 1307 3191
rect 1303 3185 1307 3186
rect 1455 3190 1459 3191
rect 1455 3185 1459 3186
rect 1479 3190 1483 3191
rect 1638 3187 1639 3191
rect 1643 3187 1644 3191
rect 1638 3186 1644 3187
rect 1687 3190 1691 3191
rect 1479 3185 1483 3186
rect 112 3165 114 3185
rect 110 3164 116 3165
rect 296 3164 298 3185
rect 370 3183 376 3184
rect 370 3179 371 3183
rect 375 3179 376 3183
rect 370 3178 376 3179
rect 110 3160 111 3164
rect 115 3160 116 3164
rect 110 3159 116 3160
rect 294 3163 300 3164
rect 294 3159 295 3163
rect 299 3159 300 3163
rect 294 3158 300 3159
rect 372 3156 374 3178
rect 432 3164 434 3185
rect 506 3183 512 3184
rect 506 3179 507 3183
rect 511 3179 512 3183
rect 506 3178 512 3179
rect 430 3163 436 3164
rect 430 3159 431 3163
rect 435 3159 436 3163
rect 430 3158 436 3159
rect 508 3156 510 3178
rect 568 3164 570 3185
rect 642 3183 648 3184
rect 642 3179 643 3183
rect 647 3179 648 3183
rect 642 3178 648 3179
rect 566 3163 572 3164
rect 566 3159 567 3163
rect 571 3159 572 3163
rect 566 3158 572 3159
rect 644 3156 646 3178
rect 704 3164 706 3185
rect 856 3164 858 3185
rect 922 3183 928 3184
rect 922 3179 923 3183
rect 927 3179 928 3183
rect 922 3178 928 3179
rect 930 3183 936 3184
rect 930 3179 931 3183
rect 935 3179 936 3183
rect 930 3178 936 3179
rect 702 3163 708 3164
rect 702 3159 703 3163
rect 707 3159 708 3163
rect 702 3158 708 3159
rect 854 3163 860 3164
rect 854 3159 855 3163
rect 859 3159 860 3163
rect 854 3158 860 3159
rect 370 3155 376 3156
rect 370 3151 371 3155
rect 375 3151 376 3155
rect 370 3150 376 3151
rect 506 3155 512 3156
rect 506 3151 507 3155
rect 511 3151 512 3155
rect 506 3150 512 3151
rect 642 3155 648 3156
rect 642 3151 643 3155
rect 647 3151 648 3155
rect 642 3150 648 3151
rect 650 3155 656 3156
rect 650 3151 651 3155
rect 655 3151 656 3155
rect 650 3150 656 3151
rect 110 3147 116 3148
rect 110 3143 111 3147
rect 115 3143 116 3147
rect 110 3142 116 3143
rect 294 3144 300 3145
rect 112 3115 114 3142
rect 294 3140 295 3144
rect 299 3140 300 3144
rect 294 3139 300 3140
rect 430 3144 436 3145
rect 430 3140 431 3144
rect 435 3140 436 3144
rect 430 3139 436 3140
rect 566 3144 572 3145
rect 566 3140 567 3144
rect 571 3140 572 3144
rect 566 3139 572 3140
rect 296 3115 298 3139
rect 432 3115 434 3139
rect 568 3115 570 3139
rect 111 3114 115 3115
rect 111 3109 115 3110
rect 295 3114 299 3115
rect 295 3109 299 3110
rect 311 3114 315 3115
rect 311 3109 315 3110
rect 407 3114 411 3115
rect 407 3109 411 3110
rect 431 3114 435 3115
rect 431 3109 435 3110
rect 503 3114 507 3115
rect 503 3109 507 3110
rect 567 3114 571 3115
rect 567 3109 571 3110
rect 599 3114 603 3115
rect 599 3109 603 3110
rect 112 3082 114 3109
rect 312 3085 314 3109
rect 350 3103 356 3104
rect 350 3099 351 3103
rect 355 3099 356 3103
rect 350 3098 356 3099
rect 310 3084 316 3085
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 310 3080 311 3084
rect 315 3080 316 3084
rect 310 3079 316 3080
rect 110 3076 116 3077
rect 310 3065 316 3066
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 310 3061 311 3065
rect 315 3061 316 3065
rect 310 3060 316 3061
rect 110 3059 116 3060
rect 112 3039 114 3059
rect 312 3039 314 3060
rect 352 3048 354 3098
rect 408 3085 410 3109
rect 504 3085 506 3109
rect 600 3085 602 3109
rect 652 3104 654 3150
rect 702 3144 708 3145
rect 702 3140 703 3144
rect 707 3140 708 3144
rect 702 3139 708 3140
rect 854 3144 860 3145
rect 854 3140 855 3144
rect 859 3140 860 3144
rect 854 3139 860 3140
rect 704 3115 706 3139
rect 856 3115 858 3139
rect 695 3114 699 3115
rect 695 3109 699 3110
rect 703 3114 707 3115
rect 703 3109 707 3110
rect 807 3114 811 3115
rect 807 3109 811 3110
rect 855 3114 859 3115
rect 855 3109 859 3110
rect 650 3103 656 3104
rect 650 3099 651 3103
rect 655 3099 656 3103
rect 650 3098 656 3099
rect 696 3085 698 3109
rect 808 3085 810 3109
rect 924 3092 926 3178
rect 932 3156 934 3178
rect 1032 3164 1034 3185
rect 1106 3183 1112 3184
rect 1106 3179 1107 3183
rect 1111 3179 1112 3183
rect 1106 3178 1112 3179
rect 1030 3163 1036 3164
rect 1030 3159 1031 3163
rect 1035 3159 1036 3163
rect 1030 3158 1036 3159
rect 1108 3156 1110 3178
rect 1232 3164 1234 3185
rect 1382 3183 1388 3184
rect 1382 3179 1383 3183
rect 1387 3179 1388 3183
rect 1382 3178 1388 3179
rect 1230 3163 1236 3164
rect 1230 3159 1231 3163
rect 1235 3159 1236 3163
rect 1230 3158 1236 3159
rect 1384 3156 1386 3178
rect 1456 3164 1458 3185
rect 1530 3183 1536 3184
rect 1530 3179 1531 3183
rect 1535 3179 1536 3183
rect 1530 3178 1536 3179
rect 1454 3163 1460 3164
rect 1454 3159 1455 3163
rect 1459 3159 1460 3163
rect 1454 3158 1460 3159
rect 1532 3156 1534 3178
rect 1640 3156 1642 3186
rect 1687 3185 1691 3186
rect 1903 3190 1907 3191
rect 1903 3185 1907 3186
rect 2007 3190 2011 3191
rect 2007 3185 2011 3186
rect 2146 3187 2152 3188
rect 1688 3164 1690 3185
rect 1904 3164 1906 3185
rect 1962 3183 1968 3184
rect 1962 3179 1963 3183
rect 1967 3179 1968 3183
rect 1962 3178 1968 3179
rect 1686 3163 1692 3164
rect 1686 3159 1687 3163
rect 1691 3159 1692 3163
rect 1686 3158 1692 3159
rect 1902 3163 1908 3164
rect 1902 3159 1903 3163
rect 1907 3159 1908 3163
rect 1902 3158 1908 3159
rect 930 3155 936 3156
rect 930 3151 931 3155
rect 935 3151 936 3155
rect 930 3150 936 3151
rect 1106 3155 1112 3156
rect 1106 3151 1107 3155
rect 1111 3151 1112 3155
rect 1106 3150 1112 3151
rect 1382 3155 1388 3156
rect 1382 3151 1383 3155
rect 1387 3151 1388 3155
rect 1382 3150 1388 3151
rect 1530 3155 1536 3156
rect 1530 3151 1531 3155
rect 1535 3151 1536 3155
rect 1530 3150 1536 3151
rect 1638 3155 1644 3156
rect 1638 3151 1639 3155
rect 1643 3151 1644 3155
rect 1638 3150 1644 3151
rect 1030 3144 1036 3145
rect 1030 3140 1031 3144
rect 1035 3140 1036 3144
rect 1030 3139 1036 3140
rect 1230 3144 1236 3145
rect 1230 3140 1231 3144
rect 1235 3140 1236 3144
rect 1230 3139 1236 3140
rect 1454 3144 1460 3145
rect 1454 3140 1455 3144
rect 1459 3140 1460 3144
rect 1454 3139 1460 3140
rect 1686 3144 1692 3145
rect 1686 3140 1687 3144
rect 1691 3140 1692 3144
rect 1686 3139 1692 3140
rect 1902 3144 1908 3145
rect 1902 3140 1903 3144
rect 1907 3140 1908 3144
rect 1902 3139 1908 3140
rect 1032 3115 1034 3139
rect 1232 3115 1234 3139
rect 1456 3115 1458 3139
rect 1688 3115 1690 3139
rect 1904 3115 1906 3139
rect 943 3114 947 3115
rect 943 3109 947 3110
rect 1031 3114 1035 3115
rect 1031 3109 1035 3110
rect 1087 3114 1091 3115
rect 1087 3109 1091 3110
rect 1231 3114 1235 3115
rect 1231 3109 1235 3110
rect 1247 3114 1251 3115
rect 1247 3109 1251 3110
rect 1407 3114 1411 3115
rect 1407 3109 1411 3110
rect 1455 3114 1459 3115
rect 1455 3109 1459 3110
rect 1575 3114 1579 3115
rect 1575 3109 1579 3110
rect 1687 3114 1691 3115
rect 1687 3109 1691 3110
rect 1751 3114 1755 3115
rect 1751 3109 1755 3110
rect 1903 3114 1907 3115
rect 1903 3109 1907 3110
rect 922 3091 928 3092
rect 922 3087 923 3091
rect 927 3087 928 3091
rect 922 3086 928 3087
rect 944 3085 946 3109
rect 1088 3085 1090 3109
rect 1248 3085 1250 3109
rect 1408 3085 1410 3109
rect 1576 3085 1578 3109
rect 1752 3085 1754 3109
rect 1904 3085 1906 3109
rect 1964 3108 1966 3178
rect 2008 3165 2010 3185
rect 2046 3183 2052 3184
rect 2046 3179 2047 3183
rect 2051 3179 2052 3183
rect 2146 3183 2147 3187
rect 2151 3183 2152 3187
rect 2282 3187 2283 3191
rect 2287 3187 2288 3191
rect 2282 3186 2288 3187
rect 2494 3191 2500 3192
rect 2494 3187 2495 3191
rect 2499 3187 2500 3191
rect 2494 3186 2500 3187
rect 2502 3191 2508 3192
rect 2502 3187 2503 3191
rect 2507 3187 2508 3191
rect 2502 3186 2508 3187
rect 2146 3182 2152 3183
rect 2046 3178 2052 3179
rect 2070 3180 2076 3181
rect 2006 3164 2012 3165
rect 2006 3160 2007 3164
rect 2011 3160 2012 3164
rect 2006 3159 2012 3160
rect 1970 3147 1976 3148
rect 1970 3143 1971 3147
rect 1975 3143 1976 3147
rect 1970 3142 1976 3143
rect 2006 3147 2012 3148
rect 2048 3147 2050 3178
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2072 3147 2074 3175
rect 2006 3143 2007 3147
rect 2011 3143 2012 3147
rect 2006 3142 2012 3143
rect 2047 3146 2051 3147
rect 1962 3107 1968 3108
rect 1962 3103 1963 3107
rect 1967 3103 1968 3107
rect 1962 3102 1968 3103
rect 406 3084 412 3085
rect 406 3080 407 3084
rect 411 3080 412 3084
rect 406 3079 412 3080
rect 502 3084 508 3085
rect 502 3080 503 3084
rect 507 3080 508 3084
rect 502 3079 508 3080
rect 598 3084 604 3085
rect 598 3080 599 3084
rect 603 3080 604 3084
rect 598 3079 604 3080
rect 694 3084 700 3085
rect 694 3080 695 3084
rect 699 3080 700 3084
rect 694 3079 700 3080
rect 806 3084 812 3085
rect 806 3080 807 3084
rect 811 3080 812 3084
rect 806 3079 812 3080
rect 942 3084 948 3085
rect 942 3080 943 3084
rect 947 3080 948 3084
rect 942 3079 948 3080
rect 1086 3084 1092 3085
rect 1086 3080 1087 3084
rect 1091 3080 1092 3084
rect 1086 3079 1092 3080
rect 1246 3084 1252 3085
rect 1246 3080 1247 3084
rect 1251 3080 1252 3084
rect 1246 3079 1252 3080
rect 1406 3084 1412 3085
rect 1406 3080 1407 3084
rect 1411 3080 1412 3084
rect 1406 3079 1412 3080
rect 1574 3084 1580 3085
rect 1574 3080 1575 3084
rect 1579 3080 1580 3084
rect 1574 3079 1580 3080
rect 1750 3084 1756 3085
rect 1750 3080 1751 3084
rect 1755 3080 1756 3084
rect 1750 3079 1756 3080
rect 1902 3084 1908 3085
rect 1902 3080 1903 3084
rect 1907 3080 1908 3084
rect 1902 3079 1908 3080
rect 386 3075 392 3076
rect 386 3071 387 3075
rect 391 3071 392 3075
rect 386 3070 392 3071
rect 482 3075 488 3076
rect 482 3071 483 3075
rect 487 3071 488 3075
rect 482 3070 488 3071
rect 578 3075 584 3076
rect 578 3071 579 3075
rect 583 3071 584 3075
rect 578 3070 584 3071
rect 674 3075 680 3076
rect 674 3071 675 3075
rect 679 3071 680 3075
rect 674 3070 680 3071
rect 770 3075 776 3076
rect 770 3071 771 3075
rect 775 3071 776 3075
rect 770 3070 776 3071
rect 778 3075 784 3076
rect 778 3071 779 3075
rect 783 3071 784 3075
rect 778 3070 784 3071
rect 1018 3075 1024 3076
rect 1018 3071 1019 3075
rect 1023 3071 1024 3075
rect 1018 3070 1024 3071
rect 1162 3075 1168 3076
rect 1162 3071 1163 3075
rect 1167 3071 1168 3075
rect 1162 3070 1168 3071
rect 1322 3075 1328 3076
rect 1322 3071 1323 3075
rect 1327 3071 1328 3075
rect 1322 3070 1328 3071
rect 1650 3075 1656 3076
rect 1650 3071 1651 3075
rect 1655 3071 1656 3075
rect 1650 3070 1656 3071
rect 1826 3075 1832 3076
rect 1826 3071 1827 3075
rect 1831 3071 1832 3075
rect 1826 3070 1832 3071
rect 1834 3075 1840 3076
rect 1834 3071 1835 3075
rect 1839 3071 1840 3075
rect 1834 3070 1840 3071
rect 388 3048 390 3070
rect 406 3065 412 3066
rect 406 3061 407 3065
rect 411 3061 412 3065
rect 406 3060 412 3061
rect 350 3047 356 3048
rect 350 3043 351 3047
rect 355 3043 356 3047
rect 350 3042 356 3043
rect 386 3047 392 3048
rect 386 3043 387 3047
rect 391 3043 392 3047
rect 386 3042 392 3043
rect 408 3039 410 3060
rect 463 3052 467 3053
rect 484 3048 486 3070
rect 502 3065 508 3066
rect 502 3061 503 3065
rect 507 3061 508 3065
rect 502 3060 508 3061
rect 463 3047 467 3048
rect 482 3047 488 3048
rect 111 3038 115 3039
rect 111 3033 115 3034
rect 311 3038 315 3039
rect 311 3033 315 3034
rect 407 3038 411 3039
rect 407 3033 411 3034
rect 423 3038 427 3039
rect 423 3033 427 3034
rect 112 3013 114 3033
rect 110 3012 116 3013
rect 424 3012 426 3033
rect 464 3032 466 3047
rect 482 3043 483 3047
rect 487 3043 488 3047
rect 482 3042 488 3043
rect 504 3039 506 3060
rect 580 3048 582 3070
rect 598 3065 604 3066
rect 598 3061 599 3065
rect 603 3061 604 3065
rect 598 3060 604 3061
rect 578 3047 584 3048
rect 578 3043 579 3047
rect 583 3043 584 3047
rect 578 3042 584 3043
rect 600 3039 602 3060
rect 676 3048 678 3070
rect 694 3065 700 3066
rect 694 3061 695 3065
rect 699 3061 700 3065
rect 694 3060 700 3061
rect 674 3047 680 3048
rect 674 3043 675 3047
rect 679 3043 680 3047
rect 674 3042 680 3043
rect 696 3039 698 3060
rect 772 3048 774 3070
rect 780 3053 782 3070
rect 806 3065 812 3066
rect 806 3061 807 3065
rect 811 3061 812 3065
rect 806 3060 812 3061
rect 942 3065 948 3066
rect 942 3061 943 3065
rect 947 3061 948 3065
rect 942 3060 948 3061
rect 779 3052 783 3053
rect 770 3047 776 3048
rect 779 3047 783 3048
rect 770 3043 771 3047
rect 775 3043 776 3047
rect 770 3042 776 3043
rect 808 3039 810 3060
rect 944 3039 946 3060
rect 1020 3048 1022 3070
rect 1086 3065 1092 3066
rect 1086 3061 1087 3065
rect 1091 3061 1092 3065
rect 1086 3060 1092 3061
rect 1018 3047 1024 3048
rect 1018 3043 1019 3047
rect 1023 3043 1024 3047
rect 1018 3042 1024 3043
rect 1088 3039 1090 3060
rect 1164 3048 1166 3070
rect 1246 3065 1252 3066
rect 1246 3061 1247 3065
rect 1251 3061 1252 3065
rect 1246 3060 1252 3061
rect 1162 3047 1168 3048
rect 1162 3043 1163 3047
rect 1167 3043 1168 3047
rect 1162 3042 1168 3043
rect 1248 3039 1250 3060
rect 1324 3048 1326 3070
rect 1406 3065 1412 3066
rect 1406 3061 1407 3065
rect 1411 3061 1412 3065
rect 1406 3060 1412 3061
rect 1574 3065 1580 3066
rect 1574 3061 1575 3065
rect 1579 3061 1580 3065
rect 1574 3060 1580 3061
rect 1322 3047 1328 3048
rect 1322 3043 1323 3047
rect 1327 3043 1328 3047
rect 1322 3042 1328 3043
rect 1278 3039 1284 3040
rect 1408 3039 1410 3060
rect 1576 3039 1578 3060
rect 1652 3048 1654 3070
rect 1750 3065 1756 3066
rect 1750 3061 1751 3065
rect 1755 3061 1756 3065
rect 1750 3060 1756 3061
rect 1650 3047 1656 3048
rect 1650 3043 1651 3047
rect 1655 3043 1656 3047
rect 1650 3042 1656 3043
rect 1752 3039 1754 3060
rect 503 3038 507 3039
rect 503 3033 507 3034
rect 519 3038 523 3039
rect 519 3033 523 3034
rect 599 3038 603 3039
rect 599 3033 603 3034
rect 615 3038 619 3039
rect 615 3033 619 3034
rect 695 3038 699 3039
rect 695 3033 699 3034
rect 711 3038 715 3039
rect 711 3033 715 3034
rect 807 3038 811 3039
rect 807 3033 811 3034
rect 815 3038 819 3039
rect 815 3033 819 3034
rect 935 3038 939 3039
rect 935 3033 939 3034
rect 943 3038 947 3039
rect 943 3033 947 3034
rect 1055 3038 1059 3039
rect 1055 3033 1059 3034
rect 1087 3038 1091 3039
rect 1087 3033 1091 3034
rect 1183 3038 1187 3039
rect 1183 3033 1187 3034
rect 1247 3038 1251 3039
rect 1278 3035 1279 3039
rect 1283 3035 1284 3039
rect 1278 3034 1284 3035
rect 1311 3038 1315 3039
rect 1247 3033 1251 3034
rect 462 3031 468 3032
rect 462 3027 463 3031
rect 467 3027 468 3031
rect 462 3026 468 3027
rect 510 3031 516 3032
rect 510 3027 511 3031
rect 515 3027 516 3031
rect 510 3026 516 3027
rect 110 3008 111 3012
rect 115 3008 116 3012
rect 110 3007 116 3008
rect 422 3011 428 3012
rect 422 3007 423 3011
rect 427 3007 428 3011
rect 422 3006 428 3007
rect 512 3004 514 3026
rect 520 3012 522 3033
rect 606 3031 612 3032
rect 606 3027 607 3031
rect 611 3027 612 3031
rect 606 3026 612 3027
rect 518 3011 524 3012
rect 518 3007 519 3011
rect 523 3007 524 3011
rect 518 3006 524 3007
rect 608 3004 610 3026
rect 616 3012 618 3033
rect 702 3031 708 3032
rect 702 3027 703 3031
rect 707 3027 708 3031
rect 702 3026 708 3027
rect 614 3011 620 3012
rect 614 3007 615 3011
rect 619 3007 620 3011
rect 614 3006 620 3007
rect 704 3004 706 3026
rect 712 3012 714 3033
rect 786 3031 792 3032
rect 786 3027 787 3031
rect 791 3027 792 3031
rect 786 3026 792 3027
rect 710 3011 716 3012
rect 710 3007 711 3011
rect 715 3007 716 3011
rect 710 3006 716 3007
rect 788 3004 790 3026
rect 816 3012 818 3033
rect 890 3031 896 3032
rect 890 3027 891 3031
rect 895 3027 896 3031
rect 890 3026 896 3027
rect 814 3011 820 3012
rect 814 3007 815 3011
rect 819 3007 820 3011
rect 814 3006 820 3007
rect 892 3004 894 3026
rect 936 3012 938 3033
rect 1010 3031 1016 3032
rect 1010 3027 1011 3031
rect 1015 3027 1016 3031
rect 1010 3026 1016 3027
rect 934 3011 940 3012
rect 934 3007 935 3011
rect 939 3007 940 3011
rect 934 3006 940 3007
rect 1012 3004 1014 3026
rect 1056 3012 1058 3033
rect 1130 3031 1136 3032
rect 1130 3027 1131 3031
rect 1135 3027 1136 3031
rect 1130 3026 1136 3027
rect 1054 3011 1060 3012
rect 1054 3007 1055 3011
rect 1059 3007 1060 3011
rect 1054 3006 1060 3007
rect 1132 3004 1134 3026
rect 1184 3012 1186 3033
rect 1258 3031 1264 3032
rect 1258 3027 1259 3031
rect 1263 3027 1264 3031
rect 1258 3026 1264 3027
rect 1182 3011 1188 3012
rect 1182 3007 1183 3011
rect 1187 3007 1188 3011
rect 1182 3006 1188 3007
rect 1260 3004 1262 3026
rect 1280 3004 1282 3034
rect 1311 3033 1315 3034
rect 1407 3038 1411 3039
rect 1407 3033 1411 3034
rect 1431 3038 1435 3039
rect 1431 3033 1435 3034
rect 1551 3038 1555 3039
rect 1551 3033 1555 3034
rect 1575 3038 1579 3039
rect 1575 3033 1579 3034
rect 1671 3038 1675 3039
rect 1671 3033 1675 3034
rect 1751 3038 1755 3039
rect 1751 3033 1755 3034
rect 1799 3038 1803 3039
rect 1799 3033 1803 3034
rect 1312 3012 1314 3033
rect 1432 3012 1434 3033
rect 1514 3031 1520 3032
rect 1514 3027 1515 3031
rect 1519 3027 1520 3031
rect 1514 3026 1520 3027
rect 1310 3011 1316 3012
rect 1310 3007 1311 3011
rect 1315 3007 1316 3011
rect 1310 3006 1316 3007
rect 1430 3011 1436 3012
rect 1430 3007 1431 3011
rect 1435 3007 1436 3011
rect 1430 3006 1436 3007
rect 1516 3004 1518 3026
rect 1552 3012 1554 3033
rect 1634 3031 1640 3032
rect 1634 3027 1635 3031
rect 1639 3027 1640 3031
rect 1634 3026 1640 3027
rect 1550 3011 1556 3012
rect 1550 3007 1551 3011
rect 1555 3007 1556 3011
rect 1550 3006 1556 3007
rect 1636 3004 1638 3026
rect 1672 3012 1674 3033
rect 1800 3012 1802 3033
rect 1828 3032 1830 3070
rect 1836 3056 1838 3070
rect 1902 3065 1908 3066
rect 1902 3061 1903 3065
rect 1907 3061 1908 3065
rect 1902 3060 1908 3061
rect 1834 3055 1840 3056
rect 1834 3051 1835 3055
rect 1839 3051 1840 3055
rect 1834 3050 1840 3051
rect 1904 3039 1906 3060
rect 1972 3048 1974 3142
rect 2008 3115 2010 3142
rect 2047 3141 2051 3142
rect 2071 3146 2075 3147
rect 2071 3141 2075 3142
rect 2007 3114 2011 3115
rect 2048 3114 2050 3141
rect 2072 3117 2074 3141
rect 2070 3116 2076 3117
rect 2007 3109 2011 3110
rect 2046 3113 2052 3114
rect 2046 3109 2047 3113
rect 2051 3109 2052 3113
rect 2070 3112 2071 3116
rect 2075 3112 2076 3116
rect 2070 3111 2076 3112
rect 2008 3082 2010 3109
rect 2046 3108 2052 3109
rect 2070 3097 2076 3098
rect 2046 3096 2052 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2070 3093 2071 3097
rect 2075 3093 2076 3097
rect 2070 3092 2076 3093
rect 2046 3091 2052 3092
rect 2006 3081 2012 3082
rect 2006 3077 2007 3081
rect 2011 3077 2012 3081
rect 2006 3076 2012 3077
rect 2048 3067 2050 3091
rect 2072 3067 2074 3092
rect 2148 3080 2150 3182
rect 2206 3180 2212 3181
rect 2206 3176 2207 3180
rect 2211 3176 2212 3180
rect 2206 3175 2212 3176
rect 2374 3180 2380 3181
rect 2374 3176 2375 3180
rect 2379 3176 2380 3180
rect 2374 3175 2380 3176
rect 2542 3180 2548 3181
rect 2542 3176 2543 3180
rect 2547 3176 2548 3180
rect 2542 3175 2548 3176
rect 2702 3180 2708 3181
rect 2702 3176 2703 3180
rect 2707 3176 2708 3180
rect 2702 3175 2708 3176
rect 2208 3147 2210 3175
rect 2376 3147 2378 3175
rect 2544 3147 2546 3175
rect 2704 3147 2706 3175
rect 2207 3146 2211 3147
rect 2207 3141 2211 3142
rect 2343 3146 2347 3147
rect 2343 3141 2347 3142
rect 2375 3146 2379 3147
rect 2375 3141 2379 3142
rect 2543 3146 2547 3147
rect 2543 3141 2547 3142
rect 2631 3146 2635 3147
rect 2631 3141 2635 3142
rect 2703 3146 2707 3147
rect 2703 3141 2707 3142
rect 2344 3117 2346 3141
rect 2632 3117 2634 3141
rect 2342 3116 2348 3117
rect 2342 3112 2343 3116
rect 2347 3112 2348 3116
rect 2342 3111 2348 3112
rect 2630 3116 2636 3117
rect 2630 3112 2631 3116
rect 2635 3112 2636 3116
rect 2630 3111 2636 3112
rect 2716 3108 2718 3214
rect 2792 3192 2794 3214
rect 2864 3200 2866 3221
rect 3016 3200 3018 3221
rect 3024 3220 3026 3258
rect 3032 3236 3034 3258
rect 3094 3253 3100 3254
rect 3094 3249 3095 3253
rect 3099 3249 3100 3253
rect 3094 3248 3100 3249
rect 3030 3235 3036 3236
rect 3030 3231 3031 3235
rect 3035 3231 3036 3235
rect 3030 3230 3036 3231
rect 3096 3227 3098 3248
rect 3180 3236 3182 3258
rect 3236 3236 3238 3338
rect 3302 3336 3308 3337
rect 3302 3332 3303 3336
rect 3307 3332 3308 3336
rect 3942 3335 3943 3339
rect 3947 3335 3948 3339
rect 3942 3334 3948 3335
rect 3302 3331 3308 3332
rect 3304 3303 3306 3331
rect 3944 3303 3946 3334
rect 3263 3302 3267 3303
rect 3263 3297 3267 3298
rect 3303 3302 3307 3303
rect 3303 3297 3307 3298
rect 3943 3302 3947 3303
rect 3943 3297 3947 3298
rect 3264 3273 3266 3297
rect 3262 3272 3268 3273
rect 3262 3268 3263 3272
rect 3267 3268 3268 3272
rect 3944 3270 3946 3297
rect 3262 3267 3268 3268
rect 3942 3269 3948 3270
rect 3942 3265 3943 3269
rect 3947 3265 3948 3269
rect 3942 3264 3948 3265
rect 3262 3253 3268 3254
rect 3262 3249 3263 3253
rect 3267 3249 3268 3253
rect 3262 3248 3268 3249
rect 3942 3252 3948 3253
rect 3942 3248 3943 3252
rect 3947 3248 3948 3252
rect 3178 3235 3184 3236
rect 3178 3231 3179 3235
rect 3183 3231 3184 3235
rect 3178 3230 3184 3231
rect 3234 3235 3240 3236
rect 3234 3231 3235 3235
rect 3239 3231 3240 3235
rect 3234 3230 3240 3231
rect 3264 3227 3266 3248
rect 3942 3247 3948 3248
rect 3944 3227 3946 3247
rect 3095 3226 3099 3227
rect 3095 3221 3099 3222
rect 3167 3226 3171 3227
rect 3167 3221 3171 3222
rect 3263 3226 3267 3227
rect 3263 3221 3267 3222
rect 3327 3226 3331 3227
rect 3327 3221 3331 3222
rect 3943 3226 3947 3227
rect 3943 3221 3947 3222
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3215 3028 3219
rect 3022 3214 3028 3215
rect 3168 3200 3170 3221
rect 3242 3219 3248 3220
rect 3242 3215 3243 3219
rect 3247 3215 3248 3219
rect 3242 3214 3248 3215
rect 2862 3199 2868 3200
rect 2862 3195 2863 3199
rect 2867 3195 2868 3199
rect 2862 3194 2868 3195
rect 3014 3199 3020 3200
rect 3014 3195 3015 3199
rect 3019 3195 3020 3199
rect 3014 3194 3020 3195
rect 3166 3199 3172 3200
rect 3166 3195 3167 3199
rect 3171 3195 3172 3199
rect 3166 3194 3172 3195
rect 3244 3192 3246 3214
rect 3328 3200 3330 3221
rect 3944 3201 3946 3221
rect 3942 3200 3948 3201
rect 3326 3199 3332 3200
rect 3326 3195 3327 3199
rect 3331 3195 3332 3199
rect 3942 3196 3943 3200
rect 3947 3196 3948 3200
rect 3942 3195 3948 3196
rect 3326 3194 3332 3195
rect 2790 3191 2796 3192
rect 2790 3187 2791 3191
rect 2795 3187 2796 3191
rect 2790 3186 2796 3187
rect 3242 3191 3248 3192
rect 3242 3187 3243 3191
rect 3247 3187 3248 3191
rect 3242 3186 3248 3187
rect 3402 3187 3408 3188
rect 3402 3183 3403 3187
rect 3407 3183 3408 3187
rect 3402 3182 3408 3183
rect 3942 3183 3948 3184
rect 2862 3180 2868 3181
rect 2862 3176 2863 3180
rect 2867 3176 2868 3180
rect 2862 3175 2868 3176
rect 3014 3180 3020 3181
rect 3014 3176 3015 3180
rect 3019 3176 3020 3180
rect 3014 3175 3020 3176
rect 3166 3180 3172 3181
rect 3166 3176 3167 3180
rect 3171 3176 3172 3180
rect 3166 3175 3172 3176
rect 3326 3180 3332 3181
rect 3326 3176 3327 3180
rect 3331 3176 3332 3180
rect 3326 3175 3332 3176
rect 2864 3147 2866 3175
rect 3016 3147 3018 3175
rect 3168 3147 3170 3175
rect 3328 3147 3330 3175
rect 2863 3146 2867 3147
rect 2863 3141 2867 3142
rect 2903 3146 2907 3147
rect 2903 3141 2907 3142
rect 3015 3146 3019 3147
rect 3015 3141 3019 3142
rect 3167 3146 3171 3147
rect 3167 3141 3171 3142
rect 3175 3146 3179 3147
rect 3175 3141 3179 3142
rect 3327 3146 3331 3147
rect 3327 3141 3331 3142
rect 2904 3117 2906 3141
rect 3176 3117 3178 3141
rect 2902 3116 2908 3117
rect 2902 3112 2903 3116
rect 2907 3112 2908 3116
rect 2902 3111 2908 3112
rect 3174 3116 3180 3117
rect 3174 3112 3175 3116
rect 3179 3112 3180 3116
rect 3174 3111 3180 3112
rect 2418 3107 2424 3108
rect 2418 3103 2419 3107
rect 2423 3103 2424 3107
rect 2418 3102 2424 3103
rect 2714 3107 2720 3108
rect 2714 3103 2715 3107
rect 2719 3103 2720 3107
rect 2714 3102 2720 3103
rect 2990 3107 2996 3108
rect 2990 3103 2991 3107
rect 2995 3103 2996 3107
rect 2990 3102 2996 3103
rect 3006 3107 3012 3108
rect 3006 3103 3007 3107
rect 3011 3103 3012 3107
rect 3006 3102 3012 3103
rect 3258 3107 3264 3108
rect 3258 3103 3259 3107
rect 3263 3103 3264 3107
rect 3258 3102 3264 3103
rect 2342 3097 2348 3098
rect 2342 3093 2343 3097
rect 2347 3093 2348 3097
rect 2342 3092 2348 3093
rect 2146 3079 2152 3080
rect 2146 3075 2147 3079
rect 2151 3075 2152 3079
rect 2146 3074 2152 3075
rect 2344 3067 2346 3092
rect 2420 3080 2422 3102
rect 2630 3097 2636 3098
rect 2630 3093 2631 3097
rect 2635 3093 2636 3097
rect 2630 3092 2636 3093
rect 2902 3097 2908 3098
rect 2902 3093 2903 3097
rect 2907 3093 2908 3097
rect 2902 3092 2908 3093
rect 2418 3079 2424 3080
rect 2418 3075 2419 3079
rect 2423 3075 2424 3079
rect 2418 3074 2424 3075
rect 2632 3067 2634 3092
rect 2826 3071 2832 3072
rect 2826 3067 2827 3071
rect 2831 3067 2832 3071
rect 2904 3067 2906 3092
rect 2047 3066 2051 3067
rect 2006 3064 2012 3065
rect 2006 3060 2007 3064
rect 2011 3060 2012 3064
rect 2047 3061 2051 3062
rect 2071 3066 2075 3067
rect 2071 3061 2075 3062
rect 2343 3066 2347 3067
rect 2343 3061 2347 3062
rect 2487 3066 2491 3067
rect 2487 3061 2491 3062
rect 2615 3066 2619 3067
rect 2615 3061 2619 3062
rect 2631 3066 2635 3067
rect 2631 3061 2635 3062
rect 2743 3066 2747 3067
rect 2826 3066 2832 3067
rect 2863 3066 2867 3067
rect 2743 3061 2747 3062
rect 2006 3059 2012 3060
rect 1970 3047 1976 3048
rect 1970 3043 1971 3047
rect 1975 3043 1976 3047
rect 1970 3042 1976 3043
rect 2008 3039 2010 3059
rect 2048 3041 2050 3061
rect 2046 3040 2052 3041
rect 2488 3040 2490 3061
rect 2494 3059 2500 3060
rect 2494 3055 2495 3059
rect 2499 3055 2500 3059
rect 2494 3054 2500 3055
rect 2562 3059 2568 3060
rect 2562 3055 2563 3059
rect 2567 3055 2568 3059
rect 2562 3054 2568 3055
rect 1903 3038 1907 3039
rect 1903 3033 1907 3034
rect 2007 3038 2011 3039
rect 2046 3036 2047 3040
rect 2051 3036 2052 3040
rect 2046 3035 2052 3036
rect 2486 3039 2492 3040
rect 2486 3035 2487 3039
rect 2491 3035 2492 3039
rect 2486 3034 2492 3035
rect 2007 3033 2011 3034
rect 1826 3031 1832 3032
rect 1826 3027 1827 3031
rect 1831 3027 1832 3031
rect 1826 3026 1832 3027
rect 1874 3031 1880 3032
rect 1874 3027 1875 3031
rect 1879 3027 1880 3031
rect 1874 3026 1880 3027
rect 1670 3011 1676 3012
rect 1670 3007 1671 3011
rect 1675 3007 1676 3011
rect 1670 3006 1676 3007
rect 1798 3011 1804 3012
rect 1798 3007 1799 3011
rect 1803 3007 1804 3011
rect 1798 3006 1804 3007
rect 1876 3004 1878 3026
rect 1882 3023 1888 3024
rect 1882 3019 1883 3023
rect 1887 3019 1888 3023
rect 1882 3018 1888 3019
rect 1884 3004 1886 3018
rect 1904 3012 1906 3033
rect 2008 3013 2010 3033
rect 2046 3023 2052 3024
rect 2046 3019 2047 3023
rect 2051 3019 2052 3023
rect 2046 3018 2052 3019
rect 2486 3020 2492 3021
rect 2006 3012 2012 3013
rect 1902 3011 1908 3012
rect 1902 3007 1903 3011
rect 1907 3007 1908 3011
rect 2006 3008 2007 3012
rect 2011 3008 2012 3012
rect 2006 3007 2012 3008
rect 1902 3006 1908 3007
rect 510 3003 516 3004
rect 510 2999 511 3003
rect 515 2999 516 3003
rect 510 2998 516 2999
rect 606 3003 612 3004
rect 606 2999 607 3003
rect 611 2999 612 3003
rect 606 2998 612 2999
rect 702 3003 708 3004
rect 702 2999 703 3003
rect 707 2999 708 3003
rect 702 2998 708 2999
rect 786 3003 792 3004
rect 786 2999 787 3003
rect 791 2999 792 3003
rect 786 2998 792 2999
rect 890 3003 896 3004
rect 890 2999 891 3003
rect 895 2999 896 3003
rect 890 2998 896 2999
rect 1010 3003 1016 3004
rect 1010 2999 1011 3003
rect 1015 2999 1016 3003
rect 1010 2998 1016 2999
rect 1130 3003 1136 3004
rect 1130 2999 1131 3003
rect 1135 2999 1136 3003
rect 1130 2998 1136 2999
rect 1258 3003 1264 3004
rect 1258 2999 1259 3003
rect 1263 2999 1264 3003
rect 1258 2998 1264 2999
rect 1278 3003 1284 3004
rect 1278 2999 1279 3003
rect 1283 2999 1284 3003
rect 1514 3003 1520 3004
rect 1278 2998 1284 2999
rect 1506 2999 1512 3000
rect 110 2995 116 2996
rect 110 2991 111 2995
rect 115 2991 116 2995
rect 1506 2995 1507 2999
rect 1511 2995 1512 2999
rect 1514 2999 1515 3003
rect 1519 2999 1520 3003
rect 1514 2998 1520 2999
rect 1634 3003 1640 3004
rect 1634 2999 1635 3003
rect 1639 2999 1640 3003
rect 1634 2998 1640 2999
rect 1874 3003 1880 3004
rect 1874 2999 1875 3003
rect 1879 2999 1880 3003
rect 1874 2998 1880 2999
rect 1882 3003 1888 3004
rect 1882 2999 1883 3003
rect 1887 2999 1888 3003
rect 1882 2998 1888 2999
rect 1506 2994 1512 2995
rect 2006 2995 2012 2996
rect 110 2990 116 2991
rect 422 2992 428 2993
rect 112 2939 114 2990
rect 422 2988 423 2992
rect 427 2988 428 2992
rect 422 2987 428 2988
rect 518 2992 524 2993
rect 518 2988 519 2992
rect 523 2988 524 2992
rect 518 2987 524 2988
rect 614 2992 620 2993
rect 614 2988 615 2992
rect 619 2988 620 2992
rect 614 2987 620 2988
rect 710 2992 716 2993
rect 710 2988 711 2992
rect 715 2988 716 2992
rect 710 2987 716 2988
rect 814 2992 820 2993
rect 814 2988 815 2992
rect 819 2988 820 2992
rect 814 2987 820 2988
rect 934 2992 940 2993
rect 934 2988 935 2992
rect 939 2988 940 2992
rect 934 2987 940 2988
rect 1054 2992 1060 2993
rect 1054 2988 1055 2992
rect 1059 2988 1060 2992
rect 1054 2987 1060 2988
rect 1182 2992 1188 2993
rect 1182 2988 1183 2992
rect 1187 2988 1188 2992
rect 1182 2987 1188 2988
rect 1310 2992 1316 2993
rect 1310 2988 1311 2992
rect 1315 2988 1316 2992
rect 1310 2987 1316 2988
rect 1430 2992 1436 2993
rect 1430 2988 1431 2992
rect 1435 2988 1436 2992
rect 1430 2987 1436 2988
rect 424 2939 426 2987
rect 520 2939 522 2987
rect 616 2939 618 2987
rect 712 2939 714 2987
rect 816 2939 818 2987
rect 936 2939 938 2987
rect 1056 2939 1058 2987
rect 1184 2939 1186 2987
rect 1312 2939 1314 2987
rect 1432 2939 1434 2987
rect 111 2938 115 2939
rect 111 2933 115 2934
rect 423 2938 427 2939
rect 423 2933 427 2934
rect 519 2938 523 2939
rect 519 2933 523 2934
rect 615 2938 619 2939
rect 615 2933 619 2934
rect 711 2938 715 2939
rect 711 2933 715 2934
rect 815 2938 819 2939
rect 815 2933 819 2934
rect 935 2938 939 2939
rect 935 2933 939 2934
rect 1055 2938 1059 2939
rect 1055 2933 1059 2934
rect 1183 2938 1187 2939
rect 1183 2933 1187 2934
rect 1311 2938 1315 2939
rect 1311 2933 1315 2934
rect 1431 2938 1435 2939
rect 1431 2933 1435 2934
rect 1479 2938 1483 2939
rect 1479 2933 1483 2934
rect 112 2906 114 2933
rect 1480 2909 1482 2933
rect 1478 2908 1484 2909
rect 110 2905 116 2906
rect 110 2901 111 2905
rect 115 2901 116 2905
rect 1478 2904 1479 2908
rect 1483 2904 1484 2908
rect 1478 2903 1484 2904
rect 110 2900 116 2901
rect 1478 2889 1484 2890
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 1478 2885 1479 2889
rect 1483 2885 1484 2889
rect 1478 2884 1484 2885
rect 110 2883 116 2884
rect 112 2855 114 2883
rect 1480 2855 1482 2884
rect 1508 2872 1510 2994
rect 1550 2992 1556 2993
rect 1550 2988 1551 2992
rect 1555 2988 1556 2992
rect 1550 2987 1556 2988
rect 1670 2992 1676 2993
rect 1670 2988 1671 2992
rect 1675 2988 1676 2992
rect 1670 2987 1676 2988
rect 1798 2992 1804 2993
rect 1798 2988 1799 2992
rect 1803 2988 1804 2992
rect 1798 2987 1804 2988
rect 1902 2992 1908 2993
rect 1902 2988 1903 2992
rect 1907 2988 1908 2992
rect 2006 2991 2007 2995
rect 2011 2991 2012 2995
rect 2006 2990 2012 2991
rect 1902 2987 1908 2988
rect 1552 2939 1554 2987
rect 1672 2939 1674 2987
rect 1800 2939 1802 2987
rect 1904 2939 1906 2987
rect 2008 2939 2010 2990
rect 2048 2987 2050 3018
rect 2486 3016 2487 3020
rect 2491 3016 2492 3020
rect 2486 3015 2492 3016
rect 2488 2987 2490 3015
rect 2047 2986 2051 2987
rect 2047 2981 2051 2982
rect 2407 2986 2411 2987
rect 2407 2981 2411 2982
rect 2487 2986 2491 2987
rect 2487 2981 2491 2982
rect 2048 2954 2050 2981
rect 2408 2957 2410 2981
rect 2406 2956 2412 2957
rect 2046 2953 2052 2954
rect 2046 2949 2047 2953
rect 2051 2949 2052 2953
rect 2406 2952 2407 2956
rect 2411 2952 2412 2956
rect 2406 2951 2412 2952
rect 2046 2948 2052 2949
rect 2496 2948 2498 3054
rect 2564 3032 2566 3054
rect 2616 3040 2618 3061
rect 2690 3059 2696 3060
rect 2690 3055 2691 3059
rect 2695 3055 2696 3059
rect 2690 3054 2696 3055
rect 2614 3039 2620 3040
rect 2614 3035 2615 3039
rect 2619 3035 2620 3039
rect 2614 3034 2620 3035
rect 2692 3032 2694 3054
rect 2744 3040 2746 3061
rect 2818 3059 2824 3060
rect 2818 3055 2819 3059
rect 2823 3055 2824 3059
rect 2818 3054 2824 3055
rect 2742 3039 2748 3040
rect 2742 3035 2743 3039
rect 2747 3035 2748 3039
rect 2742 3034 2748 3035
rect 2820 3032 2822 3054
rect 2828 3032 2830 3066
rect 2863 3061 2867 3062
rect 2903 3066 2907 3067
rect 2903 3061 2907 3062
rect 2983 3066 2987 3067
rect 2983 3061 2987 3062
rect 2864 3040 2866 3061
rect 2984 3040 2986 3061
rect 2992 3060 2994 3102
rect 3008 3080 3010 3102
rect 3174 3097 3180 3098
rect 3174 3093 3175 3097
rect 3179 3093 3180 3097
rect 3174 3092 3180 3093
rect 3006 3079 3012 3080
rect 3006 3075 3007 3079
rect 3011 3075 3012 3079
rect 3006 3074 3012 3075
rect 3176 3067 3178 3092
rect 3260 3080 3262 3102
rect 3404 3080 3406 3182
rect 3942 3179 3943 3183
rect 3947 3179 3948 3183
rect 3942 3178 3948 3179
rect 3944 3147 3946 3178
rect 3447 3146 3451 3147
rect 3447 3141 3451 3142
rect 3943 3146 3947 3147
rect 3943 3141 3947 3142
rect 3448 3117 3450 3141
rect 3446 3116 3452 3117
rect 3446 3112 3447 3116
rect 3451 3112 3452 3116
rect 3944 3114 3946 3141
rect 3446 3111 3452 3112
rect 3942 3113 3948 3114
rect 3942 3109 3943 3113
rect 3947 3109 3948 3113
rect 3942 3108 3948 3109
rect 3446 3097 3452 3098
rect 3446 3093 3447 3097
rect 3451 3093 3452 3097
rect 3446 3092 3452 3093
rect 3942 3096 3948 3097
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 3258 3079 3264 3080
rect 3258 3075 3259 3079
rect 3263 3075 3264 3079
rect 3258 3074 3264 3075
rect 3402 3079 3408 3080
rect 3402 3075 3403 3079
rect 3407 3075 3408 3079
rect 3402 3074 3408 3075
rect 3448 3067 3450 3092
rect 3942 3091 3948 3092
rect 3944 3067 3946 3091
rect 3103 3066 3107 3067
rect 3103 3061 3107 3062
rect 3175 3066 3179 3067
rect 3175 3061 3179 3062
rect 3215 3066 3219 3067
rect 3215 3061 3219 3062
rect 3327 3066 3331 3067
rect 3327 3061 3331 3062
rect 3431 3066 3435 3067
rect 3431 3061 3435 3062
rect 3447 3066 3451 3067
rect 3447 3061 3451 3062
rect 3535 3066 3539 3067
rect 3535 3061 3539 3062
rect 3639 3066 3643 3067
rect 3639 3061 3643 3062
rect 3743 3066 3747 3067
rect 3743 3061 3747 3062
rect 3839 3066 3843 3067
rect 3839 3061 3843 3062
rect 3943 3066 3947 3067
rect 3943 3061 3947 3062
rect 2990 3059 2996 3060
rect 2990 3055 2991 3059
rect 2995 3055 2996 3059
rect 2990 3054 2996 3055
rect 3058 3059 3064 3060
rect 3058 3055 3059 3059
rect 3063 3055 3064 3059
rect 3058 3054 3064 3055
rect 2862 3039 2868 3040
rect 2862 3035 2863 3039
rect 2867 3035 2868 3039
rect 2862 3034 2868 3035
rect 2982 3039 2988 3040
rect 2982 3035 2983 3039
rect 2987 3035 2988 3039
rect 2982 3034 2988 3035
rect 3060 3032 3062 3054
rect 3104 3040 3106 3061
rect 3198 3059 3204 3060
rect 3198 3055 3199 3059
rect 3203 3055 3204 3059
rect 3198 3054 3204 3055
rect 3102 3039 3108 3040
rect 3102 3035 3103 3039
rect 3107 3035 3108 3039
rect 3102 3034 3108 3035
rect 3200 3032 3202 3054
rect 3216 3040 3218 3061
rect 3290 3059 3296 3060
rect 3290 3055 3291 3059
rect 3295 3055 3296 3059
rect 3290 3054 3296 3055
rect 3214 3039 3220 3040
rect 3214 3035 3215 3039
rect 3219 3035 3220 3039
rect 3214 3034 3220 3035
rect 3292 3032 3294 3054
rect 3328 3040 3330 3061
rect 3402 3059 3408 3060
rect 3402 3055 3403 3059
rect 3407 3055 3408 3059
rect 3402 3054 3408 3055
rect 3326 3039 3332 3040
rect 3326 3035 3327 3039
rect 3331 3035 3332 3039
rect 3326 3034 3332 3035
rect 3404 3032 3406 3054
rect 3432 3040 3434 3061
rect 3536 3040 3538 3061
rect 3602 3059 3608 3060
rect 3602 3055 3603 3059
rect 3607 3055 3608 3059
rect 3602 3054 3608 3055
rect 3610 3059 3616 3060
rect 3610 3055 3611 3059
rect 3615 3055 3616 3059
rect 3610 3054 3616 3055
rect 3430 3039 3436 3040
rect 3430 3035 3431 3039
rect 3435 3035 3436 3039
rect 3430 3034 3436 3035
rect 3534 3039 3540 3040
rect 3534 3035 3535 3039
rect 3539 3035 3540 3039
rect 3534 3034 3540 3035
rect 2562 3031 2568 3032
rect 2562 3027 2563 3031
rect 2567 3027 2568 3031
rect 2562 3026 2568 3027
rect 2690 3031 2696 3032
rect 2690 3027 2691 3031
rect 2695 3027 2696 3031
rect 2690 3026 2696 3027
rect 2818 3031 2824 3032
rect 2818 3027 2819 3031
rect 2823 3027 2824 3031
rect 2818 3026 2824 3027
rect 2826 3031 2832 3032
rect 2826 3027 2827 3031
rect 2831 3027 2832 3031
rect 2826 3026 2832 3027
rect 3058 3031 3064 3032
rect 3058 3027 3059 3031
rect 3063 3027 3064 3031
rect 3058 3026 3064 3027
rect 3198 3031 3204 3032
rect 3198 3027 3199 3031
rect 3203 3027 3204 3031
rect 3198 3026 3204 3027
rect 3290 3031 3296 3032
rect 3290 3027 3291 3031
rect 3295 3027 3296 3031
rect 3290 3026 3296 3027
rect 3402 3031 3408 3032
rect 3402 3027 3403 3031
rect 3407 3027 3408 3031
rect 3402 3026 3408 3027
rect 2614 3020 2620 3021
rect 2614 3016 2615 3020
rect 2619 3016 2620 3020
rect 2614 3015 2620 3016
rect 2742 3020 2748 3021
rect 2742 3016 2743 3020
rect 2747 3016 2748 3020
rect 2742 3015 2748 3016
rect 2862 3020 2868 3021
rect 2862 3016 2863 3020
rect 2867 3016 2868 3020
rect 2862 3015 2868 3016
rect 2982 3020 2988 3021
rect 2982 3016 2983 3020
rect 2987 3016 2988 3020
rect 2982 3015 2988 3016
rect 3102 3020 3108 3021
rect 3102 3016 3103 3020
rect 3107 3016 3108 3020
rect 3102 3015 3108 3016
rect 3214 3020 3220 3021
rect 3214 3016 3215 3020
rect 3219 3016 3220 3020
rect 3214 3015 3220 3016
rect 3326 3020 3332 3021
rect 3326 3016 3327 3020
rect 3331 3016 3332 3020
rect 3326 3015 3332 3016
rect 3430 3020 3436 3021
rect 3430 3016 3431 3020
rect 3435 3016 3436 3020
rect 3430 3015 3436 3016
rect 3534 3020 3540 3021
rect 3534 3016 3535 3020
rect 3539 3016 3540 3020
rect 3534 3015 3540 3016
rect 2616 2987 2618 3015
rect 2744 2987 2746 3015
rect 2864 2987 2866 3015
rect 2984 2987 2986 3015
rect 3104 2987 3106 3015
rect 3216 2987 3218 3015
rect 3328 2987 3330 3015
rect 3432 2987 3434 3015
rect 3536 2987 3538 3015
rect 2575 2986 2579 2987
rect 2575 2981 2579 2982
rect 2615 2986 2619 2987
rect 2615 2981 2619 2982
rect 2743 2986 2747 2987
rect 2743 2981 2747 2982
rect 2767 2986 2771 2987
rect 2767 2981 2771 2982
rect 2863 2986 2867 2987
rect 2863 2981 2867 2982
rect 2967 2986 2971 2987
rect 2967 2981 2971 2982
rect 2983 2986 2987 2987
rect 2983 2981 2987 2982
rect 3103 2986 3107 2987
rect 3103 2981 3107 2982
rect 3183 2986 3187 2987
rect 3183 2981 3187 2982
rect 3215 2986 3219 2987
rect 3215 2981 3219 2982
rect 3327 2986 3331 2987
rect 3327 2981 3331 2982
rect 3399 2986 3403 2987
rect 3399 2981 3403 2982
rect 3431 2986 3435 2987
rect 3431 2981 3435 2982
rect 3535 2986 3539 2987
rect 3535 2981 3539 2982
rect 2576 2957 2578 2981
rect 2768 2957 2770 2981
rect 2968 2957 2970 2981
rect 3184 2957 3186 2981
rect 3400 2957 3402 2981
rect 2574 2956 2580 2957
rect 2574 2952 2575 2956
rect 2579 2952 2580 2956
rect 2574 2951 2580 2952
rect 2766 2956 2772 2957
rect 2766 2952 2767 2956
rect 2771 2952 2772 2956
rect 2766 2951 2772 2952
rect 2966 2956 2972 2957
rect 2966 2952 2967 2956
rect 2971 2952 2972 2956
rect 2966 2951 2972 2952
rect 3182 2956 3188 2957
rect 3182 2952 3183 2956
rect 3187 2952 3188 2956
rect 3182 2951 3188 2952
rect 3398 2956 3404 2957
rect 3398 2952 3399 2956
rect 3403 2952 3404 2956
rect 3398 2951 3404 2952
rect 3604 2948 3606 3054
rect 3612 3032 3614 3054
rect 3640 3040 3642 3061
rect 3714 3059 3720 3060
rect 3714 3055 3715 3059
rect 3719 3055 3720 3059
rect 3714 3054 3720 3055
rect 3638 3039 3644 3040
rect 3638 3035 3639 3039
rect 3643 3035 3644 3039
rect 3638 3034 3644 3035
rect 3716 3032 3718 3054
rect 3744 3040 3746 3061
rect 3818 3059 3824 3060
rect 3818 3055 3819 3059
rect 3823 3055 3824 3059
rect 3818 3054 3824 3055
rect 3742 3039 3748 3040
rect 3742 3035 3743 3039
rect 3747 3035 3748 3039
rect 3742 3034 3748 3035
rect 3820 3032 3822 3054
rect 3840 3040 3842 3061
rect 3944 3041 3946 3061
rect 3942 3040 3948 3041
rect 3838 3039 3844 3040
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3942 3036 3943 3040
rect 3947 3036 3948 3040
rect 3942 3035 3948 3036
rect 3838 3034 3844 3035
rect 3610 3031 3616 3032
rect 3610 3027 3611 3031
rect 3615 3027 3616 3031
rect 3610 3026 3616 3027
rect 3714 3031 3720 3032
rect 3714 3027 3715 3031
rect 3719 3027 3720 3031
rect 3714 3026 3720 3027
rect 3818 3031 3824 3032
rect 3818 3027 3819 3031
rect 3823 3027 3824 3031
rect 3818 3026 3824 3027
rect 3906 3023 3912 3024
rect 3638 3020 3644 3021
rect 3638 3016 3639 3020
rect 3643 3016 3644 3020
rect 3638 3015 3644 3016
rect 3742 3020 3748 3021
rect 3742 3016 3743 3020
rect 3747 3016 3748 3020
rect 3742 3015 3748 3016
rect 3838 3020 3844 3021
rect 3838 3016 3839 3020
rect 3843 3016 3844 3020
rect 3906 3019 3907 3023
rect 3911 3019 3912 3023
rect 3906 3018 3912 3019
rect 3942 3023 3948 3024
rect 3942 3019 3943 3023
rect 3947 3019 3948 3023
rect 3942 3018 3948 3019
rect 3838 3015 3844 3016
rect 3640 2987 3642 3015
rect 3744 2987 3746 3015
rect 3840 2987 3842 3015
rect 3623 2986 3627 2987
rect 3623 2981 3627 2982
rect 3639 2986 3643 2987
rect 3639 2981 3643 2982
rect 3743 2986 3747 2987
rect 3743 2981 3747 2982
rect 3839 2986 3843 2987
rect 3839 2981 3843 2982
rect 3624 2957 3626 2981
rect 3840 2957 3842 2981
rect 3622 2956 3628 2957
rect 3622 2952 3623 2956
rect 3627 2952 3628 2956
rect 3622 2951 3628 2952
rect 3838 2956 3844 2957
rect 3838 2952 3839 2956
rect 3843 2952 3844 2956
rect 3838 2951 3844 2952
rect 2494 2947 2500 2948
rect 2494 2943 2495 2947
rect 2499 2943 2500 2947
rect 2494 2942 2500 2943
rect 2502 2947 2508 2948
rect 2502 2943 2503 2947
rect 2507 2943 2508 2947
rect 2502 2942 2508 2943
rect 2694 2947 2700 2948
rect 2694 2943 2695 2947
rect 2699 2943 2700 2947
rect 2694 2942 2700 2943
rect 2922 2947 2928 2948
rect 2922 2943 2923 2947
rect 2927 2943 2928 2947
rect 2922 2942 2928 2943
rect 3114 2947 3120 2948
rect 3114 2943 3115 2947
rect 3119 2943 3120 2947
rect 3114 2942 3120 2943
rect 3474 2947 3480 2948
rect 3474 2943 3475 2947
rect 3479 2943 3480 2947
rect 3474 2942 3480 2943
rect 3602 2947 3608 2948
rect 3602 2943 3603 2947
rect 3607 2943 3608 2947
rect 3602 2942 3608 2943
rect 1551 2938 1555 2939
rect 1551 2933 1555 2934
rect 1575 2938 1579 2939
rect 1575 2933 1579 2934
rect 1671 2938 1675 2939
rect 1671 2933 1675 2934
rect 1767 2938 1771 2939
rect 1767 2933 1771 2934
rect 1799 2938 1803 2939
rect 1799 2933 1803 2934
rect 1863 2938 1867 2939
rect 1863 2933 1867 2934
rect 1903 2938 1907 2939
rect 1903 2933 1907 2934
rect 2007 2938 2011 2939
rect 2406 2937 2412 2938
rect 2007 2933 2011 2934
rect 2046 2936 2052 2937
rect 1576 2909 1578 2933
rect 1672 2909 1674 2933
rect 1768 2909 1770 2933
rect 1864 2909 1866 2933
rect 1574 2908 1580 2909
rect 1574 2904 1575 2908
rect 1579 2904 1580 2908
rect 1574 2903 1580 2904
rect 1670 2908 1676 2909
rect 1670 2904 1671 2908
rect 1675 2904 1676 2908
rect 1670 2903 1676 2904
rect 1766 2908 1772 2909
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1862 2908 1868 2909
rect 1862 2904 1863 2908
rect 1867 2904 1868 2908
rect 2008 2906 2010 2933
rect 2046 2932 2047 2936
rect 2051 2932 2052 2936
rect 2406 2933 2407 2937
rect 2411 2933 2412 2937
rect 2406 2932 2412 2933
rect 2046 2931 2052 2932
rect 1862 2903 1868 2904
rect 2006 2905 2012 2906
rect 2006 2901 2007 2905
rect 2011 2901 2012 2905
rect 2006 2900 2012 2901
rect 1554 2899 1560 2900
rect 1554 2895 1555 2899
rect 1559 2895 1560 2899
rect 1554 2894 1560 2895
rect 1650 2899 1656 2900
rect 1650 2895 1651 2899
rect 1655 2895 1656 2899
rect 1650 2894 1656 2895
rect 1746 2899 1752 2900
rect 1746 2895 1747 2899
rect 1751 2895 1752 2899
rect 1746 2894 1752 2895
rect 1842 2899 1848 2900
rect 1842 2895 1843 2899
rect 1847 2895 1848 2899
rect 1842 2894 1848 2895
rect 1930 2899 1936 2900
rect 1930 2895 1931 2899
rect 1935 2895 1936 2899
rect 2048 2895 2050 2931
rect 2408 2895 2410 2932
rect 2504 2920 2506 2942
rect 2574 2937 2580 2938
rect 2574 2933 2575 2937
rect 2579 2933 2580 2937
rect 2574 2932 2580 2933
rect 2502 2919 2508 2920
rect 2502 2915 2503 2919
rect 2507 2915 2508 2919
rect 2502 2914 2508 2915
rect 2576 2895 2578 2932
rect 2696 2920 2698 2942
rect 2766 2937 2772 2938
rect 2766 2933 2767 2937
rect 2771 2933 2772 2937
rect 2766 2932 2772 2933
rect 2694 2919 2700 2920
rect 2694 2915 2695 2919
rect 2699 2915 2700 2919
rect 2694 2914 2700 2915
rect 2768 2895 2770 2932
rect 2924 2920 2926 2942
rect 2966 2937 2972 2938
rect 2966 2933 2967 2937
rect 2971 2933 2972 2937
rect 2966 2932 2972 2933
rect 2922 2919 2928 2920
rect 2922 2915 2923 2919
rect 2927 2915 2928 2919
rect 2922 2914 2928 2915
rect 2968 2895 2970 2932
rect 3116 2920 3118 2942
rect 3182 2937 3188 2938
rect 3182 2933 3183 2937
rect 3187 2933 3188 2937
rect 3182 2932 3188 2933
rect 3398 2937 3404 2938
rect 3398 2933 3399 2937
rect 3403 2933 3404 2937
rect 3398 2932 3404 2933
rect 3114 2919 3120 2920
rect 3114 2915 3115 2919
rect 3119 2915 3120 2919
rect 3114 2914 3120 2915
rect 3130 2915 3136 2916
rect 3130 2911 3131 2915
rect 3135 2911 3136 2915
rect 3130 2910 3136 2911
rect 1930 2894 1936 2895
rect 2047 2894 2051 2895
rect 1556 2872 1558 2894
rect 1574 2889 1580 2890
rect 1574 2885 1575 2889
rect 1579 2885 1580 2889
rect 1574 2884 1580 2885
rect 1506 2871 1512 2872
rect 1506 2867 1507 2871
rect 1511 2867 1512 2871
rect 1506 2866 1512 2867
rect 1554 2871 1560 2872
rect 1554 2867 1555 2871
rect 1559 2867 1560 2871
rect 1554 2866 1560 2867
rect 1576 2855 1578 2884
rect 1652 2872 1654 2894
rect 1670 2889 1676 2890
rect 1670 2885 1671 2889
rect 1675 2885 1676 2889
rect 1670 2884 1676 2885
rect 1650 2871 1656 2872
rect 1650 2867 1651 2871
rect 1655 2867 1656 2871
rect 1650 2866 1656 2867
rect 1672 2855 1674 2884
rect 1748 2872 1750 2894
rect 1766 2889 1772 2890
rect 1766 2885 1767 2889
rect 1771 2885 1772 2889
rect 1766 2884 1772 2885
rect 1746 2871 1752 2872
rect 1746 2867 1747 2871
rect 1751 2867 1752 2871
rect 1746 2866 1752 2867
rect 1768 2855 1770 2884
rect 1844 2872 1846 2894
rect 1862 2889 1868 2890
rect 1862 2885 1863 2889
rect 1867 2885 1868 2889
rect 1862 2884 1868 2885
rect 1842 2871 1848 2872
rect 1842 2867 1843 2871
rect 1847 2867 1848 2871
rect 1842 2866 1848 2867
rect 1864 2855 1866 2884
rect 111 2854 115 2855
rect 111 2849 115 2850
rect 279 2854 283 2855
rect 447 2854 451 2855
rect 279 2849 283 2850
rect 354 2851 360 2852
rect 112 2829 114 2849
rect 110 2828 116 2829
rect 280 2828 282 2849
rect 354 2847 355 2851
rect 359 2847 360 2851
rect 447 2849 451 2850
rect 631 2854 635 2855
rect 631 2849 635 2850
rect 815 2854 819 2855
rect 815 2849 819 2850
rect 999 2854 1003 2855
rect 999 2849 1003 2850
rect 1183 2854 1187 2855
rect 1183 2849 1187 2850
rect 1359 2854 1363 2855
rect 1359 2849 1363 2850
rect 1479 2854 1483 2855
rect 1479 2849 1483 2850
rect 1527 2854 1531 2855
rect 1527 2849 1531 2850
rect 1575 2854 1579 2855
rect 1575 2849 1579 2850
rect 1671 2854 1675 2855
rect 1671 2849 1675 2850
rect 1695 2854 1699 2855
rect 1695 2849 1699 2850
rect 1767 2854 1771 2855
rect 1767 2849 1771 2850
rect 1863 2854 1867 2855
rect 1863 2849 1867 2850
rect 354 2846 360 2847
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 110 2823 116 2824
rect 278 2827 284 2828
rect 278 2823 279 2827
rect 283 2823 284 2827
rect 278 2822 284 2823
rect 356 2820 358 2846
rect 438 2843 444 2844
rect 438 2839 439 2843
rect 443 2839 444 2843
rect 438 2838 444 2839
rect 354 2819 360 2820
rect 354 2815 355 2819
rect 359 2815 360 2819
rect 354 2814 360 2815
rect 110 2811 116 2812
rect 110 2807 111 2811
rect 115 2807 116 2811
rect 110 2806 116 2807
rect 278 2808 284 2809
rect 112 2779 114 2806
rect 278 2804 279 2808
rect 283 2804 284 2808
rect 278 2803 284 2804
rect 280 2779 282 2803
rect 111 2778 115 2779
rect 111 2773 115 2774
rect 239 2778 243 2779
rect 239 2773 243 2774
rect 279 2778 283 2779
rect 279 2773 283 2774
rect 351 2778 355 2779
rect 351 2773 355 2774
rect 112 2746 114 2773
rect 240 2749 242 2773
rect 352 2749 354 2773
rect 238 2748 244 2749
rect 110 2745 116 2746
rect 110 2741 111 2745
rect 115 2741 116 2745
rect 238 2744 239 2748
rect 243 2744 244 2748
rect 238 2743 244 2744
rect 350 2748 356 2749
rect 350 2744 351 2748
rect 355 2744 356 2748
rect 350 2743 356 2744
rect 110 2740 116 2741
rect 440 2740 442 2838
rect 448 2828 450 2849
rect 522 2847 528 2848
rect 522 2843 523 2847
rect 527 2843 528 2847
rect 522 2842 528 2843
rect 446 2827 452 2828
rect 446 2823 447 2827
rect 451 2823 452 2827
rect 446 2822 452 2823
rect 524 2820 526 2842
rect 632 2828 634 2849
rect 706 2847 712 2848
rect 706 2843 707 2847
rect 711 2843 712 2847
rect 706 2842 712 2843
rect 630 2827 636 2828
rect 630 2823 631 2827
rect 635 2823 636 2827
rect 630 2822 636 2823
rect 708 2820 710 2842
rect 816 2828 818 2849
rect 890 2847 896 2848
rect 890 2843 891 2847
rect 895 2843 896 2847
rect 890 2842 896 2843
rect 814 2827 820 2828
rect 814 2823 815 2827
rect 819 2823 820 2827
rect 814 2822 820 2823
rect 892 2820 894 2842
rect 1000 2828 1002 2849
rect 1184 2828 1186 2849
rect 1258 2847 1264 2848
rect 1258 2843 1259 2847
rect 1263 2843 1264 2847
rect 1258 2842 1264 2843
rect 998 2827 1004 2828
rect 998 2823 999 2827
rect 1003 2823 1004 2827
rect 998 2822 1004 2823
rect 1182 2827 1188 2828
rect 1182 2823 1183 2827
rect 1187 2823 1188 2827
rect 1182 2822 1188 2823
rect 1260 2820 1262 2842
rect 1360 2828 1362 2849
rect 1458 2839 1464 2840
rect 1458 2835 1459 2839
rect 1463 2835 1464 2839
rect 1458 2834 1464 2835
rect 1358 2827 1364 2828
rect 1358 2823 1359 2827
rect 1363 2823 1364 2827
rect 1358 2822 1364 2823
rect 1460 2820 1462 2834
rect 1528 2828 1530 2849
rect 1610 2847 1616 2848
rect 1610 2843 1611 2847
rect 1615 2843 1616 2847
rect 1610 2842 1616 2843
rect 1526 2827 1532 2828
rect 1526 2823 1527 2827
rect 1531 2823 1532 2827
rect 1526 2822 1532 2823
rect 1612 2820 1614 2842
rect 1696 2828 1698 2849
rect 1778 2847 1784 2848
rect 1778 2843 1779 2847
rect 1783 2843 1784 2847
rect 1778 2842 1784 2843
rect 1694 2827 1700 2828
rect 1694 2823 1695 2827
rect 1699 2823 1700 2827
rect 1694 2822 1700 2823
rect 1780 2820 1782 2842
rect 1864 2828 1866 2849
rect 1932 2848 1934 2894
rect 2047 2889 2051 2890
rect 2407 2894 2411 2895
rect 2407 2889 2411 2890
rect 2551 2894 2555 2895
rect 2551 2889 2555 2890
rect 2575 2894 2579 2895
rect 2575 2889 2579 2890
rect 2671 2894 2675 2895
rect 2671 2889 2675 2890
rect 2767 2894 2771 2895
rect 2767 2889 2771 2890
rect 2799 2894 2803 2895
rect 2799 2889 2803 2890
rect 2927 2894 2931 2895
rect 2927 2889 2931 2890
rect 2967 2894 2971 2895
rect 2967 2889 2971 2890
rect 3055 2894 3059 2895
rect 3055 2889 3059 2890
rect 2006 2888 2012 2889
rect 2006 2884 2007 2888
rect 2011 2884 2012 2888
rect 2006 2883 2012 2884
rect 2008 2855 2010 2883
rect 2048 2869 2050 2889
rect 2046 2868 2052 2869
rect 2552 2868 2554 2889
rect 2626 2887 2632 2888
rect 2626 2883 2627 2887
rect 2631 2883 2632 2887
rect 2626 2882 2632 2883
rect 2046 2864 2047 2868
rect 2051 2864 2052 2868
rect 2046 2863 2052 2864
rect 2550 2867 2556 2868
rect 2550 2863 2551 2867
rect 2555 2863 2556 2867
rect 2550 2862 2556 2863
rect 2628 2860 2630 2882
rect 2672 2868 2674 2889
rect 2746 2887 2752 2888
rect 2746 2883 2747 2887
rect 2751 2883 2752 2887
rect 2746 2882 2752 2883
rect 2670 2867 2676 2868
rect 2670 2863 2671 2867
rect 2675 2863 2676 2867
rect 2670 2862 2676 2863
rect 2748 2860 2750 2882
rect 2800 2868 2802 2889
rect 2874 2887 2880 2888
rect 2874 2883 2875 2887
rect 2879 2883 2880 2887
rect 2874 2882 2880 2883
rect 2798 2867 2804 2868
rect 2798 2863 2799 2867
rect 2803 2863 2804 2867
rect 2798 2862 2804 2863
rect 2876 2860 2878 2882
rect 2914 2879 2920 2880
rect 2914 2875 2915 2879
rect 2919 2875 2920 2879
rect 2914 2874 2920 2875
rect 2626 2859 2632 2860
rect 2626 2855 2627 2859
rect 2631 2855 2632 2859
rect 2007 2854 2011 2855
rect 2626 2854 2632 2855
rect 2746 2859 2752 2860
rect 2746 2855 2747 2859
rect 2751 2855 2752 2859
rect 2746 2854 2752 2855
rect 2874 2859 2880 2860
rect 2874 2855 2875 2859
rect 2879 2855 2880 2859
rect 2874 2854 2880 2855
rect 2007 2849 2011 2850
rect 2046 2851 2052 2852
rect 1930 2847 1936 2848
rect 1930 2843 1931 2847
rect 1935 2843 1936 2847
rect 1930 2842 1936 2843
rect 2008 2829 2010 2849
rect 2046 2847 2047 2851
rect 2051 2847 2052 2851
rect 2046 2846 2052 2847
rect 2550 2848 2556 2849
rect 2006 2828 2012 2829
rect 1862 2827 1868 2828
rect 1862 2823 1863 2827
rect 1867 2823 1868 2827
rect 2006 2824 2007 2828
rect 2011 2824 2012 2828
rect 2006 2823 2012 2824
rect 1862 2822 1868 2823
rect 522 2819 528 2820
rect 522 2815 523 2819
rect 527 2815 528 2819
rect 522 2814 528 2815
rect 706 2819 712 2820
rect 706 2815 707 2819
rect 711 2815 712 2819
rect 706 2814 712 2815
rect 890 2819 896 2820
rect 890 2815 891 2819
rect 895 2815 896 2819
rect 890 2814 896 2815
rect 966 2819 972 2820
rect 966 2815 967 2819
rect 971 2815 972 2819
rect 966 2814 972 2815
rect 1258 2819 1264 2820
rect 1258 2815 1259 2819
rect 1263 2815 1264 2819
rect 1458 2819 1464 2820
rect 1258 2814 1264 2815
rect 1434 2815 1440 2816
rect 446 2808 452 2809
rect 446 2804 447 2808
rect 451 2804 452 2808
rect 446 2803 452 2804
rect 630 2808 636 2809
rect 630 2804 631 2808
rect 635 2804 636 2808
rect 630 2803 636 2804
rect 814 2808 820 2809
rect 814 2804 815 2808
rect 819 2804 820 2808
rect 814 2803 820 2804
rect 448 2779 450 2803
rect 632 2779 634 2803
rect 816 2779 818 2803
rect 447 2778 451 2779
rect 447 2773 451 2774
rect 471 2778 475 2779
rect 471 2773 475 2774
rect 607 2778 611 2779
rect 607 2773 611 2774
rect 631 2778 635 2779
rect 631 2773 635 2774
rect 743 2778 747 2779
rect 743 2773 747 2774
rect 815 2778 819 2779
rect 815 2773 819 2774
rect 879 2778 883 2779
rect 879 2773 883 2774
rect 472 2749 474 2773
rect 608 2749 610 2773
rect 744 2749 746 2773
rect 880 2749 882 2773
rect 470 2748 476 2749
rect 470 2744 471 2748
rect 475 2744 476 2748
rect 470 2743 476 2744
rect 606 2748 612 2749
rect 606 2744 607 2748
rect 611 2744 612 2748
rect 606 2743 612 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 878 2748 884 2749
rect 878 2744 879 2748
rect 883 2744 884 2748
rect 878 2743 884 2744
rect 314 2739 320 2740
rect 314 2735 315 2739
rect 319 2735 320 2739
rect 314 2734 320 2735
rect 426 2739 432 2740
rect 426 2735 427 2739
rect 431 2735 432 2739
rect 426 2734 432 2735
rect 438 2739 444 2740
rect 438 2735 439 2739
rect 443 2735 444 2739
rect 438 2734 444 2735
rect 554 2739 560 2740
rect 554 2735 555 2739
rect 559 2735 560 2739
rect 554 2734 560 2735
rect 726 2739 732 2740
rect 726 2735 727 2739
rect 731 2735 732 2739
rect 726 2734 732 2735
rect 850 2739 856 2740
rect 850 2735 851 2739
rect 855 2735 856 2739
rect 850 2734 856 2735
rect 238 2729 244 2730
rect 110 2728 116 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 238 2725 239 2729
rect 243 2725 244 2729
rect 238 2724 244 2725
rect 110 2723 116 2724
rect 112 2703 114 2723
rect 240 2703 242 2724
rect 316 2712 318 2734
rect 350 2729 356 2730
rect 350 2725 351 2729
rect 355 2725 356 2729
rect 350 2724 356 2725
rect 314 2711 320 2712
rect 298 2707 304 2708
rect 298 2703 299 2707
rect 303 2703 304 2707
rect 314 2707 315 2711
rect 319 2707 320 2711
rect 314 2706 320 2707
rect 352 2703 354 2724
rect 428 2712 430 2734
rect 470 2729 476 2730
rect 470 2725 471 2729
rect 475 2725 476 2729
rect 470 2724 476 2725
rect 426 2711 432 2712
rect 426 2707 427 2711
rect 431 2707 432 2711
rect 426 2706 432 2707
rect 472 2703 474 2724
rect 111 2702 115 2703
rect 111 2697 115 2698
rect 223 2702 227 2703
rect 223 2697 227 2698
rect 239 2702 243 2703
rect 298 2702 304 2703
rect 351 2702 355 2703
rect 239 2697 243 2698
rect 112 2677 114 2697
rect 110 2676 116 2677
rect 224 2676 226 2697
rect 110 2672 111 2676
rect 115 2672 116 2676
rect 110 2671 116 2672
rect 222 2675 228 2676
rect 222 2671 223 2675
rect 227 2671 228 2675
rect 222 2670 228 2671
rect 300 2668 302 2702
rect 351 2697 355 2698
rect 367 2702 371 2703
rect 367 2697 371 2698
rect 471 2702 475 2703
rect 471 2697 475 2698
rect 503 2702 507 2703
rect 503 2697 507 2698
rect 306 2695 312 2696
rect 306 2691 307 2695
rect 311 2691 312 2695
rect 306 2690 312 2691
rect 308 2668 310 2690
rect 368 2676 370 2697
rect 434 2695 440 2696
rect 434 2691 435 2695
rect 439 2691 440 2695
rect 434 2690 440 2691
rect 366 2675 372 2676
rect 366 2671 367 2675
rect 371 2671 372 2675
rect 366 2670 372 2671
rect 298 2667 304 2668
rect 298 2663 299 2667
rect 303 2663 304 2667
rect 298 2662 304 2663
rect 306 2667 312 2668
rect 306 2663 307 2667
rect 311 2663 312 2667
rect 306 2662 312 2663
rect 110 2659 116 2660
rect 110 2655 111 2659
rect 115 2655 116 2659
rect 110 2654 116 2655
rect 222 2656 228 2657
rect 112 2627 114 2654
rect 222 2652 223 2656
rect 227 2652 228 2656
rect 222 2651 228 2652
rect 366 2656 372 2657
rect 366 2652 367 2656
rect 371 2652 372 2656
rect 366 2651 372 2652
rect 224 2627 226 2651
rect 368 2627 370 2651
rect 111 2626 115 2627
rect 111 2621 115 2622
rect 175 2626 179 2627
rect 175 2621 179 2622
rect 223 2626 227 2627
rect 223 2621 227 2622
rect 367 2626 371 2627
rect 367 2621 371 2622
rect 112 2594 114 2621
rect 176 2597 178 2621
rect 368 2597 370 2621
rect 174 2596 180 2597
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 174 2592 175 2596
rect 179 2592 180 2596
rect 174 2591 180 2592
rect 366 2596 372 2597
rect 366 2592 367 2596
rect 371 2592 372 2596
rect 366 2591 372 2592
rect 110 2588 116 2589
rect 436 2588 438 2690
rect 504 2676 506 2697
rect 556 2696 558 2734
rect 606 2729 612 2730
rect 606 2725 607 2729
rect 611 2725 612 2729
rect 606 2724 612 2725
rect 608 2703 610 2724
rect 728 2712 730 2734
rect 742 2729 748 2730
rect 742 2725 743 2729
rect 747 2725 748 2729
rect 742 2724 748 2725
rect 726 2711 732 2712
rect 726 2707 727 2711
rect 731 2707 732 2711
rect 726 2706 732 2707
rect 744 2703 746 2724
rect 852 2712 854 2734
rect 878 2729 884 2730
rect 878 2725 879 2729
rect 883 2725 884 2729
rect 878 2724 884 2725
rect 850 2711 856 2712
rect 850 2707 851 2711
rect 855 2707 856 2711
rect 850 2706 856 2707
rect 880 2703 882 2724
rect 968 2712 970 2814
rect 1434 2811 1435 2815
rect 1439 2811 1440 2815
rect 1458 2815 1459 2819
rect 1463 2815 1464 2819
rect 1458 2814 1464 2815
rect 1610 2819 1616 2820
rect 1610 2815 1611 2819
rect 1615 2815 1616 2819
rect 1610 2814 1616 2815
rect 1778 2819 1784 2820
rect 2048 2819 2050 2846
rect 2550 2844 2551 2848
rect 2555 2844 2556 2848
rect 2550 2843 2556 2844
rect 2670 2848 2676 2849
rect 2670 2844 2671 2848
rect 2675 2844 2676 2848
rect 2670 2843 2676 2844
rect 2798 2848 2804 2849
rect 2798 2844 2799 2848
rect 2803 2844 2804 2848
rect 2798 2843 2804 2844
rect 2552 2819 2554 2843
rect 2672 2819 2674 2843
rect 2800 2819 2802 2843
rect 1778 2815 1779 2819
rect 1783 2815 1784 2819
rect 1778 2814 1784 2815
rect 2047 2818 2051 2819
rect 2047 2813 2051 2814
rect 2439 2818 2443 2819
rect 2439 2813 2443 2814
rect 2551 2818 2555 2819
rect 2551 2813 2555 2814
rect 2567 2818 2571 2819
rect 2567 2813 2571 2814
rect 2671 2818 2675 2819
rect 2671 2813 2675 2814
rect 2695 2818 2699 2819
rect 2695 2813 2699 2814
rect 2799 2818 2803 2819
rect 2799 2813 2803 2814
rect 2831 2818 2835 2819
rect 2831 2813 2835 2814
rect 1434 2810 1440 2811
rect 2006 2811 2012 2812
rect 998 2808 1004 2809
rect 998 2804 999 2808
rect 1003 2804 1004 2808
rect 998 2803 1004 2804
rect 1182 2808 1188 2809
rect 1182 2804 1183 2808
rect 1187 2804 1188 2808
rect 1182 2803 1188 2804
rect 1358 2808 1364 2809
rect 1358 2804 1359 2808
rect 1363 2804 1364 2808
rect 1358 2803 1364 2804
rect 1000 2779 1002 2803
rect 1184 2779 1186 2803
rect 1360 2779 1362 2803
rect 999 2778 1003 2779
rect 999 2773 1003 2774
rect 1015 2778 1019 2779
rect 1015 2773 1019 2774
rect 1151 2778 1155 2779
rect 1151 2773 1155 2774
rect 1183 2778 1187 2779
rect 1183 2773 1187 2774
rect 1287 2778 1291 2779
rect 1287 2773 1291 2774
rect 1359 2778 1363 2779
rect 1359 2773 1363 2774
rect 1423 2778 1427 2779
rect 1423 2773 1427 2774
rect 1016 2749 1018 2773
rect 1152 2749 1154 2773
rect 1288 2749 1290 2773
rect 1424 2749 1426 2773
rect 1014 2748 1020 2749
rect 1014 2744 1015 2748
rect 1019 2744 1020 2748
rect 1014 2743 1020 2744
rect 1150 2748 1156 2749
rect 1150 2744 1151 2748
rect 1155 2744 1156 2748
rect 1150 2743 1156 2744
rect 1286 2748 1292 2749
rect 1286 2744 1287 2748
rect 1291 2744 1292 2748
rect 1286 2743 1292 2744
rect 1422 2748 1428 2749
rect 1422 2744 1423 2748
rect 1427 2744 1428 2748
rect 1422 2743 1428 2744
rect 1090 2739 1096 2740
rect 1090 2735 1091 2739
rect 1095 2735 1096 2739
rect 1090 2734 1096 2735
rect 1238 2739 1244 2740
rect 1238 2735 1239 2739
rect 1243 2735 1244 2739
rect 1238 2734 1244 2735
rect 1246 2739 1252 2740
rect 1246 2735 1247 2739
rect 1251 2735 1252 2739
rect 1246 2734 1252 2735
rect 1014 2729 1020 2730
rect 1014 2725 1015 2729
rect 1019 2725 1020 2729
rect 1014 2724 1020 2725
rect 966 2711 972 2712
rect 966 2707 967 2711
rect 971 2707 972 2711
rect 966 2706 972 2707
rect 1016 2703 1018 2724
rect 1092 2712 1094 2734
rect 1150 2729 1156 2730
rect 1150 2725 1151 2729
rect 1155 2725 1156 2729
rect 1150 2724 1156 2725
rect 1090 2711 1096 2712
rect 1090 2707 1091 2711
rect 1095 2707 1096 2711
rect 1090 2706 1096 2707
rect 1152 2703 1154 2724
rect 607 2702 611 2703
rect 607 2697 611 2698
rect 639 2702 643 2703
rect 639 2697 643 2698
rect 743 2702 747 2703
rect 743 2697 747 2698
rect 767 2702 771 2703
rect 767 2697 771 2698
rect 879 2702 883 2703
rect 879 2697 883 2698
rect 887 2702 891 2703
rect 887 2697 891 2698
rect 999 2702 1003 2703
rect 999 2697 1003 2698
rect 1015 2702 1019 2703
rect 1015 2697 1019 2698
rect 1111 2702 1115 2703
rect 1111 2697 1115 2698
rect 1151 2702 1155 2703
rect 1151 2697 1155 2698
rect 1231 2702 1235 2703
rect 1231 2697 1235 2698
rect 554 2695 560 2696
rect 554 2691 555 2695
rect 559 2691 560 2695
rect 554 2690 560 2691
rect 578 2695 584 2696
rect 578 2691 579 2695
rect 583 2691 584 2695
rect 578 2690 584 2691
rect 502 2675 508 2676
rect 502 2671 503 2675
rect 507 2671 508 2675
rect 502 2670 508 2671
rect 580 2668 582 2690
rect 640 2676 642 2697
rect 714 2695 720 2696
rect 714 2691 715 2695
rect 719 2691 720 2695
rect 714 2690 720 2691
rect 638 2675 644 2676
rect 638 2671 639 2675
rect 643 2671 644 2675
rect 638 2670 644 2671
rect 716 2668 718 2690
rect 768 2676 770 2697
rect 888 2676 890 2697
rect 970 2695 976 2696
rect 970 2691 971 2695
rect 975 2691 976 2695
rect 970 2690 976 2691
rect 766 2675 772 2676
rect 766 2671 767 2675
rect 771 2671 772 2675
rect 766 2670 772 2671
rect 886 2675 892 2676
rect 886 2671 887 2675
rect 891 2671 892 2675
rect 886 2670 892 2671
rect 972 2668 974 2690
rect 1000 2676 1002 2697
rect 1082 2695 1088 2696
rect 1082 2691 1083 2695
rect 1087 2691 1088 2695
rect 1082 2690 1088 2691
rect 998 2675 1004 2676
rect 998 2671 999 2675
rect 1003 2671 1004 2675
rect 998 2670 1004 2671
rect 1084 2668 1086 2690
rect 1112 2676 1114 2697
rect 1232 2676 1234 2697
rect 1240 2696 1242 2734
rect 1248 2720 1250 2734
rect 1286 2729 1292 2730
rect 1286 2725 1287 2729
rect 1291 2725 1292 2729
rect 1286 2724 1292 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1246 2719 1252 2720
rect 1246 2715 1247 2719
rect 1251 2715 1252 2719
rect 1246 2714 1252 2715
rect 1288 2703 1290 2724
rect 1424 2703 1426 2724
rect 1436 2712 1438 2810
rect 1526 2808 1532 2809
rect 1526 2804 1527 2808
rect 1531 2804 1532 2808
rect 1526 2803 1532 2804
rect 1694 2808 1700 2809
rect 1694 2804 1695 2808
rect 1699 2804 1700 2808
rect 1694 2803 1700 2804
rect 1862 2808 1868 2809
rect 1862 2804 1863 2808
rect 1867 2804 1868 2808
rect 2006 2807 2007 2811
rect 2011 2807 2012 2811
rect 2006 2806 2012 2807
rect 1862 2803 1868 2804
rect 1528 2779 1530 2803
rect 1696 2779 1698 2803
rect 1864 2779 1866 2803
rect 2008 2779 2010 2806
rect 2048 2786 2050 2813
rect 2440 2789 2442 2813
rect 2568 2789 2570 2813
rect 2696 2789 2698 2813
rect 2832 2789 2834 2813
rect 2438 2788 2444 2789
rect 2046 2785 2052 2786
rect 2046 2781 2047 2785
rect 2051 2781 2052 2785
rect 2438 2784 2439 2788
rect 2443 2784 2444 2788
rect 2438 2783 2444 2784
rect 2566 2788 2572 2789
rect 2566 2784 2567 2788
rect 2571 2784 2572 2788
rect 2566 2783 2572 2784
rect 2694 2788 2700 2789
rect 2694 2784 2695 2788
rect 2699 2784 2700 2788
rect 2694 2783 2700 2784
rect 2830 2788 2836 2789
rect 2830 2784 2831 2788
rect 2835 2784 2836 2788
rect 2830 2783 2836 2784
rect 2046 2780 2052 2781
rect 2916 2780 2918 2874
rect 2928 2868 2930 2889
rect 3002 2887 3008 2888
rect 3002 2883 3003 2887
rect 3007 2883 3008 2887
rect 3002 2882 3008 2883
rect 2926 2867 2932 2868
rect 2926 2863 2927 2867
rect 2931 2863 2932 2867
rect 2926 2862 2932 2863
rect 3004 2860 3006 2882
rect 3056 2868 3058 2889
rect 3054 2867 3060 2868
rect 3054 2863 3055 2867
rect 3059 2863 3060 2867
rect 3054 2862 3060 2863
rect 3132 2860 3134 2910
rect 3184 2895 3186 2932
rect 3400 2895 3402 2932
rect 3476 2920 3478 2942
rect 3622 2937 3628 2938
rect 3622 2933 3623 2937
rect 3627 2933 3628 2937
rect 3622 2932 3628 2933
rect 3838 2937 3844 2938
rect 3838 2933 3839 2937
rect 3843 2933 3844 2937
rect 3838 2932 3844 2933
rect 3474 2919 3480 2920
rect 3474 2915 3475 2919
rect 3479 2915 3480 2919
rect 3474 2914 3480 2915
rect 3624 2895 3626 2932
rect 3840 2895 3842 2932
rect 3908 2920 3910 3018
rect 3944 2987 3946 3018
rect 3943 2986 3947 2987
rect 3943 2981 3947 2982
rect 3944 2954 3946 2981
rect 3942 2953 3948 2954
rect 3942 2949 3943 2953
rect 3947 2949 3948 2953
rect 3942 2948 3948 2949
rect 3914 2947 3920 2948
rect 3914 2943 3915 2947
rect 3919 2943 3920 2947
rect 3914 2942 3920 2943
rect 3906 2919 3912 2920
rect 3906 2915 3907 2919
rect 3911 2915 3912 2919
rect 3906 2914 3912 2915
rect 3183 2894 3187 2895
rect 3183 2889 3187 2890
rect 3311 2894 3315 2895
rect 3311 2889 3315 2890
rect 3399 2894 3403 2895
rect 3399 2889 3403 2890
rect 3439 2894 3443 2895
rect 3439 2889 3443 2890
rect 3575 2894 3579 2895
rect 3575 2889 3579 2890
rect 3623 2894 3627 2895
rect 3623 2889 3627 2890
rect 3839 2894 3843 2895
rect 3839 2889 3843 2890
rect 3184 2868 3186 2889
rect 3266 2887 3272 2888
rect 3266 2883 3267 2887
rect 3271 2883 3272 2887
rect 3266 2882 3272 2883
rect 3182 2867 3188 2868
rect 3182 2863 3183 2867
rect 3187 2863 3188 2867
rect 3182 2862 3188 2863
rect 3268 2860 3270 2882
rect 3312 2868 3314 2889
rect 3440 2868 3442 2889
rect 3466 2887 3472 2888
rect 3466 2883 3467 2887
rect 3471 2883 3472 2887
rect 3466 2882 3472 2883
rect 3514 2887 3520 2888
rect 3514 2883 3515 2887
rect 3519 2883 3520 2887
rect 3514 2882 3520 2883
rect 3310 2867 3316 2868
rect 3310 2863 3311 2867
rect 3315 2863 3316 2867
rect 3310 2862 3316 2863
rect 3438 2867 3444 2868
rect 3438 2863 3439 2867
rect 3443 2863 3444 2867
rect 3438 2862 3444 2863
rect 3002 2859 3008 2860
rect 3002 2855 3003 2859
rect 3007 2855 3008 2859
rect 3002 2854 3008 2855
rect 3130 2859 3136 2860
rect 3130 2855 3131 2859
rect 3135 2855 3136 2859
rect 3130 2854 3136 2855
rect 3142 2859 3148 2860
rect 3142 2855 3143 2859
rect 3147 2855 3148 2859
rect 3142 2854 3148 2855
rect 3266 2859 3272 2860
rect 3266 2855 3267 2859
rect 3271 2855 3272 2859
rect 3266 2854 3272 2855
rect 2926 2848 2932 2849
rect 2926 2844 2927 2848
rect 2931 2844 2932 2848
rect 2926 2843 2932 2844
rect 3054 2848 3060 2849
rect 3054 2844 3055 2848
rect 3059 2844 3060 2848
rect 3054 2843 3060 2844
rect 2928 2819 2930 2843
rect 3056 2819 3058 2843
rect 2927 2818 2931 2819
rect 2927 2813 2931 2814
rect 2967 2818 2971 2819
rect 2967 2813 2971 2814
rect 3055 2818 3059 2819
rect 3055 2813 3059 2814
rect 3103 2818 3107 2819
rect 3103 2813 3107 2814
rect 2968 2789 2970 2813
rect 3104 2789 3106 2813
rect 2966 2788 2972 2789
rect 2966 2784 2967 2788
rect 2971 2784 2972 2788
rect 2966 2783 2972 2784
rect 3102 2788 3108 2789
rect 3102 2784 3103 2788
rect 3107 2784 3108 2788
rect 3102 2783 3108 2784
rect 2514 2779 2520 2780
rect 1527 2778 1531 2779
rect 1527 2773 1531 2774
rect 1567 2778 1571 2779
rect 1567 2773 1571 2774
rect 1695 2778 1699 2779
rect 1695 2773 1699 2774
rect 1863 2778 1867 2779
rect 1863 2773 1867 2774
rect 2007 2778 2011 2779
rect 2514 2775 2515 2779
rect 2519 2775 2520 2779
rect 2514 2774 2520 2775
rect 2642 2779 2648 2780
rect 2642 2775 2643 2779
rect 2647 2775 2648 2779
rect 2642 2774 2648 2775
rect 2770 2779 2776 2780
rect 2770 2775 2771 2779
rect 2775 2775 2776 2779
rect 2770 2774 2776 2775
rect 2906 2779 2912 2780
rect 2906 2775 2907 2779
rect 2911 2775 2912 2779
rect 2906 2774 2912 2775
rect 2914 2779 2920 2780
rect 2914 2775 2915 2779
rect 2919 2775 2920 2779
rect 2914 2774 2920 2775
rect 2007 2773 2011 2774
rect 1568 2749 1570 2773
rect 1566 2748 1572 2749
rect 1566 2744 1567 2748
rect 1571 2744 1572 2748
rect 2008 2746 2010 2773
rect 2438 2769 2444 2770
rect 2046 2768 2052 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2438 2765 2439 2769
rect 2443 2765 2444 2769
rect 2438 2764 2444 2765
rect 2046 2763 2052 2764
rect 1566 2743 1572 2744
rect 2006 2745 2012 2746
rect 2006 2741 2007 2745
rect 2011 2741 2012 2745
rect 2006 2740 2012 2741
rect 1498 2739 1504 2740
rect 1498 2735 1499 2739
rect 1503 2735 1504 2739
rect 1498 2734 1504 2735
rect 1506 2739 1512 2740
rect 1506 2735 1507 2739
rect 1511 2735 1512 2739
rect 2048 2735 2050 2763
rect 2440 2735 2442 2764
rect 2516 2752 2518 2774
rect 2566 2769 2572 2770
rect 2566 2765 2567 2769
rect 2571 2765 2572 2769
rect 2566 2764 2572 2765
rect 2514 2751 2520 2752
rect 2514 2747 2515 2751
rect 2519 2747 2520 2751
rect 2514 2746 2520 2747
rect 2568 2735 2570 2764
rect 2644 2752 2646 2774
rect 2694 2769 2700 2770
rect 2694 2765 2695 2769
rect 2699 2765 2700 2769
rect 2694 2764 2700 2765
rect 2642 2751 2648 2752
rect 2642 2747 2643 2751
rect 2647 2747 2648 2751
rect 2642 2746 2648 2747
rect 2696 2735 2698 2764
rect 2772 2752 2774 2774
rect 2830 2769 2836 2770
rect 2830 2765 2831 2769
rect 2835 2765 2836 2769
rect 2830 2764 2836 2765
rect 2770 2751 2776 2752
rect 2770 2747 2771 2751
rect 2775 2747 2776 2751
rect 2770 2746 2776 2747
rect 2832 2735 2834 2764
rect 2908 2752 2910 2774
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2966 2764 2972 2765
rect 3102 2769 3108 2770
rect 3102 2765 3103 2769
rect 3107 2765 3108 2769
rect 3102 2764 3108 2765
rect 2906 2751 2912 2752
rect 2906 2747 2907 2751
rect 2911 2747 2912 2751
rect 2906 2746 2912 2747
rect 2968 2735 2970 2764
rect 3104 2735 3106 2764
rect 3144 2752 3146 2854
rect 3182 2848 3188 2849
rect 3182 2844 3183 2848
rect 3187 2844 3188 2848
rect 3182 2843 3188 2844
rect 3310 2848 3316 2849
rect 3310 2844 3311 2848
rect 3315 2844 3316 2848
rect 3310 2843 3316 2844
rect 3438 2848 3444 2849
rect 3438 2844 3439 2848
rect 3443 2844 3444 2848
rect 3438 2843 3444 2844
rect 3184 2819 3186 2843
rect 3312 2819 3314 2843
rect 3440 2819 3442 2843
rect 3183 2818 3187 2819
rect 3183 2813 3187 2814
rect 3247 2818 3251 2819
rect 3247 2813 3251 2814
rect 3311 2818 3315 2819
rect 3311 2813 3315 2814
rect 3391 2818 3395 2819
rect 3391 2813 3395 2814
rect 3439 2818 3443 2819
rect 3439 2813 3443 2814
rect 3248 2789 3250 2813
rect 3392 2789 3394 2813
rect 3246 2788 3252 2789
rect 3246 2784 3247 2788
rect 3251 2784 3252 2788
rect 3246 2783 3252 2784
rect 3390 2788 3396 2789
rect 3390 2784 3391 2788
rect 3395 2784 3396 2788
rect 3390 2783 3396 2784
rect 3468 2780 3470 2882
rect 3516 2860 3518 2882
rect 3522 2879 3528 2880
rect 3522 2875 3523 2879
rect 3527 2875 3528 2879
rect 3522 2874 3528 2875
rect 3524 2860 3526 2874
rect 3576 2868 3578 2889
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3574 2862 3580 2863
rect 3514 2859 3520 2860
rect 3514 2855 3515 2859
rect 3519 2855 3520 2859
rect 3514 2854 3520 2855
rect 3522 2859 3528 2860
rect 3522 2855 3523 2859
rect 3527 2855 3528 2859
rect 3522 2854 3528 2855
rect 3574 2848 3580 2849
rect 3574 2844 3575 2848
rect 3579 2844 3580 2848
rect 3574 2843 3580 2844
rect 3576 2819 3578 2843
rect 3543 2818 3547 2819
rect 3543 2813 3547 2814
rect 3575 2818 3579 2819
rect 3575 2813 3579 2814
rect 3703 2818 3707 2819
rect 3703 2813 3707 2814
rect 3839 2818 3843 2819
rect 3839 2813 3843 2814
rect 3544 2789 3546 2813
rect 3704 2789 3706 2813
rect 3840 2789 3842 2813
rect 3542 2788 3548 2789
rect 3542 2784 3543 2788
rect 3547 2784 3548 2788
rect 3542 2783 3548 2784
rect 3702 2788 3708 2789
rect 3702 2784 3703 2788
rect 3707 2784 3708 2788
rect 3702 2783 3708 2784
rect 3838 2788 3844 2789
rect 3838 2784 3839 2788
rect 3843 2784 3844 2788
rect 3838 2783 3844 2784
rect 3178 2779 3184 2780
rect 3178 2775 3179 2779
rect 3183 2775 3184 2779
rect 3178 2774 3184 2775
rect 3322 2779 3328 2780
rect 3322 2775 3323 2779
rect 3327 2775 3328 2779
rect 3322 2774 3328 2775
rect 3466 2779 3472 2780
rect 3466 2775 3467 2779
rect 3471 2775 3472 2779
rect 3466 2774 3472 2775
rect 3474 2779 3480 2780
rect 3474 2775 3475 2779
rect 3479 2775 3480 2779
rect 3474 2774 3480 2775
rect 3630 2779 3636 2780
rect 3630 2775 3631 2779
rect 3635 2775 3636 2779
rect 3630 2774 3636 2775
rect 3906 2779 3912 2780
rect 3906 2775 3907 2779
rect 3911 2775 3912 2779
rect 3906 2774 3912 2775
rect 3180 2752 3182 2774
rect 3246 2769 3252 2770
rect 3246 2765 3247 2769
rect 3251 2765 3252 2769
rect 3246 2764 3252 2765
rect 3142 2751 3148 2752
rect 3142 2747 3143 2751
rect 3147 2747 3148 2751
rect 3142 2746 3148 2747
rect 3178 2751 3184 2752
rect 3178 2747 3179 2751
rect 3183 2747 3184 2751
rect 3178 2746 3184 2747
rect 3248 2735 3250 2764
rect 1506 2734 1512 2735
rect 2047 2734 2051 2735
rect 1500 2712 1502 2734
rect 1508 2720 1510 2734
rect 1566 2729 1572 2730
rect 2047 2729 2051 2730
rect 2335 2734 2339 2735
rect 2335 2729 2339 2730
rect 2439 2734 2443 2735
rect 2439 2729 2443 2730
rect 2495 2734 2499 2735
rect 2495 2729 2499 2730
rect 2567 2734 2571 2735
rect 2567 2729 2571 2730
rect 2663 2734 2667 2735
rect 2663 2729 2667 2730
rect 2695 2734 2699 2735
rect 2695 2729 2699 2730
rect 2831 2734 2835 2735
rect 2831 2729 2835 2730
rect 2967 2734 2971 2735
rect 2967 2729 2971 2730
rect 2999 2734 3003 2735
rect 2999 2729 3003 2730
rect 3103 2734 3107 2735
rect 3103 2729 3107 2730
rect 3167 2734 3171 2735
rect 3167 2729 3171 2730
rect 3247 2734 3251 2735
rect 3247 2729 3251 2730
rect 1566 2725 1567 2729
rect 1571 2725 1572 2729
rect 1566 2724 1572 2725
rect 2006 2728 2012 2729
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 1506 2719 1512 2720
rect 1506 2715 1507 2719
rect 1511 2715 1512 2719
rect 1506 2714 1512 2715
rect 1434 2711 1440 2712
rect 1434 2707 1435 2711
rect 1439 2707 1440 2711
rect 1434 2706 1440 2707
rect 1498 2711 1504 2712
rect 1498 2707 1499 2711
rect 1503 2707 1504 2711
rect 1498 2706 1504 2707
rect 1568 2703 1570 2724
rect 2006 2723 2012 2724
rect 2008 2703 2010 2723
rect 2048 2709 2050 2729
rect 2046 2708 2052 2709
rect 2336 2708 2338 2729
rect 2402 2727 2408 2728
rect 2402 2723 2403 2727
rect 2407 2723 2408 2727
rect 2402 2722 2408 2723
rect 2410 2727 2416 2728
rect 2410 2723 2411 2727
rect 2415 2723 2416 2727
rect 2410 2722 2416 2723
rect 2046 2704 2047 2708
rect 2051 2704 2052 2708
rect 2046 2703 2052 2704
rect 2334 2707 2340 2708
rect 2334 2703 2335 2707
rect 2339 2703 2340 2707
rect 1287 2702 1291 2703
rect 1287 2697 1291 2698
rect 1351 2702 1355 2703
rect 1351 2697 1355 2698
rect 1423 2702 1427 2703
rect 1423 2697 1427 2698
rect 1567 2702 1571 2703
rect 1567 2697 1571 2698
rect 2007 2702 2011 2703
rect 2334 2702 2340 2703
rect 2007 2697 2011 2698
rect 1238 2695 1244 2696
rect 1238 2691 1239 2695
rect 1243 2691 1244 2695
rect 1238 2690 1244 2691
rect 1306 2695 1312 2696
rect 1306 2691 1307 2695
rect 1311 2691 1312 2695
rect 1306 2690 1312 2691
rect 1110 2675 1116 2676
rect 1110 2671 1111 2675
rect 1115 2671 1116 2675
rect 1110 2670 1116 2671
rect 1230 2675 1236 2676
rect 1230 2671 1231 2675
rect 1235 2671 1236 2675
rect 1230 2670 1236 2671
rect 1308 2668 1310 2690
rect 1314 2687 1320 2688
rect 1314 2683 1315 2687
rect 1319 2683 1320 2687
rect 1314 2682 1320 2683
rect 1316 2668 1318 2682
rect 1352 2676 1354 2697
rect 2008 2677 2010 2697
rect 2046 2691 2052 2692
rect 2046 2687 2047 2691
rect 2051 2687 2052 2691
rect 2046 2686 2052 2687
rect 2334 2688 2340 2689
rect 2006 2676 2012 2677
rect 1350 2675 1356 2676
rect 1350 2671 1351 2675
rect 1355 2671 1356 2675
rect 2006 2672 2007 2676
rect 2011 2672 2012 2676
rect 2006 2671 2012 2672
rect 1350 2670 1356 2671
rect 578 2667 584 2668
rect 578 2663 579 2667
rect 583 2663 584 2667
rect 578 2662 584 2663
rect 714 2667 720 2668
rect 714 2663 715 2667
rect 719 2663 720 2667
rect 714 2662 720 2663
rect 750 2667 756 2668
rect 750 2663 751 2667
rect 755 2663 756 2667
rect 750 2662 756 2663
rect 878 2667 884 2668
rect 878 2663 879 2667
rect 883 2663 884 2667
rect 878 2662 884 2663
rect 970 2667 976 2668
rect 970 2663 971 2667
rect 975 2663 976 2667
rect 970 2662 976 2663
rect 1082 2667 1088 2668
rect 1082 2663 1083 2667
rect 1087 2663 1088 2667
rect 1082 2662 1088 2663
rect 1306 2667 1312 2668
rect 1306 2663 1307 2667
rect 1311 2663 1312 2667
rect 1306 2662 1312 2663
rect 1314 2667 1320 2668
rect 1314 2663 1315 2667
rect 1319 2663 1320 2667
rect 1314 2662 1320 2663
rect 502 2656 508 2657
rect 502 2652 503 2656
rect 507 2652 508 2656
rect 502 2651 508 2652
rect 638 2656 644 2657
rect 638 2652 639 2656
rect 643 2652 644 2656
rect 638 2651 644 2652
rect 504 2627 506 2651
rect 640 2627 642 2651
rect 503 2626 507 2627
rect 503 2621 507 2622
rect 543 2626 547 2627
rect 543 2621 547 2622
rect 639 2626 643 2627
rect 639 2621 643 2622
rect 711 2626 715 2627
rect 711 2621 715 2622
rect 544 2597 546 2621
rect 712 2597 714 2621
rect 542 2596 548 2597
rect 542 2592 543 2596
rect 547 2592 548 2596
rect 542 2591 548 2592
rect 710 2596 716 2597
rect 710 2592 711 2596
rect 715 2592 716 2596
rect 710 2591 716 2592
rect 250 2587 256 2588
rect 250 2583 251 2587
rect 255 2583 256 2587
rect 250 2582 256 2583
rect 434 2587 440 2588
rect 434 2583 435 2587
rect 439 2583 440 2587
rect 434 2582 440 2583
rect 618 2587 624 2588
rect 618 2583 619 2587
rect 623 2583 624 2587
rect 618 2582 624 2583
rect 630 2587 636 2588
rect 630 2583 631 2587
rect 635 2583 636 2587
rect 630 2582 636 2583
rect 174 2577 180 2578
rect 110 2576 116 2577
rect 110 2572 111 2576
rect 115 2572 116 2576
rect 174 2573 175 2577
rect 179 2573 180 2577
rect 174 2572 180 2573
rect 110 2571 116 2572
rect 112 2547 114 2571
rect 176 2547 178 2572
rect 252 2560 254 2582
rect 366 2577 372 2578
rect 366 2573 367 2577
rect 371 2573 372 2577
rect 366 2572 372 2573
rect 542 2577 548 2578
rect 542 2573 543 2577
rect 547 2573 548 2577
rect 542 2572 548 2573
rect 250 2559 256 2560
rect 210 2555 216 2556
rect 210 2551 211 2555
rect 215 2551 216 2555
rect 250 2555 251 2559
rect 255 2555 256 2559
rect 250 2554 256 2555
rect 210 2550 216 2551
rect 111 2546 115 2547
rect 111 2541 115 2542
rect 135 2546 139 2547
rect 135 2541 139 2542
rect 175 2546 179 2547
rect 175 2541 179 2542
rect 112 2521 114 2541
rect 110 2520 116 2521
rect 136 2520 138 2541
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 134 2519 140 2520
rect 134 2515 135 2519
rect 139 2515 140 2519
rect 134 2514 140 2515
rect 212 2512 214 2550
rect 368 2547 370 2572
rect 544 2547 546 2572
rect 271 2546 275 2547
rect 271 2541 275 2542
rect 367 2546 371 2547
rect 367 2541 371 2542
rect 439 2546 443 2547
rect 439 2541 443 2542
rect 543 2546 547 2547
rect 543 2541 547 2542
rect 607 2546 611 2547
rect 607 2541 611 2542
rect 218 2539 224 2540
rect 218 2535 219 2539
rect 223 2535 224 2539
rect 218 2534 224 2535
rect 220 2512 222 2534
rect 272 2520 274 2541
rect 354 2539 360 2540
rect 354 2535 355 2539
rect 359 2535 360 2539
rect 354 2534 360 2535
rect 270 2519 276 2520
rect 270 2515 271 2519
rect 275 2515 276 2519
rect 270 2514 276 2515
rect 356 2512 358 2534
rect 440 2520 442 2541
rect 478 2539 484 2540
rect 478 2535 479 2539
rect 483 2535 484 2539
rect 478 2534 484 2535
rect 438 2519 444 2520
rect 438 2515 439 2519
rect 443 2515 444 2519
rect 438 2514 444 2515
rect 210 2511 216 2512
rect 210 2507 211 2511
rect 215 2507 216 2511
rect 210 2506 216 2507
rect 218 2511 224 2512
rect 218 2507 219 2511
rect 223 2507 224 2511
rect 218 2506 224 2507
rect 354 2511 360 2512
rect 354 2507 355 2511
rect 359 2507 360 2511
rect 354 2506 360 2507
rect 110 2503 116 2504
rect 110 2499 111 2503
rect 115 2499 116 2503
rect 110 2498 116 2499
rect 134 2500 140 2501
rect 112 2467 114 2498
rect 134 2496 135 2500
rect 139 2496 140 2500
rect 134 2495 140 2496
rect 270 2500 276 2501
rect 270 2496 271 2500
rect 275 2496 276 2500
rect 270 2495 276 2496
rect 438 2500 444 2501
rect 438 2496 439 2500
rect 443 2496 444 2500
rect 438 2495 444 2496
rect 136 2467 138 2495
rect 272 2467 274 2495
rect 440 2467 442 2495
rect 111 2466 115 2467
rect 111 2461 115 2462
rect 135 2466 139 2467
rect 135 2461 139 2462
rect 271 2466 275 2467
rect 271 2461 275 2462
rect 311 2466 315 2467
rect 311 2461 315 2462
rect 439 2466 443 2467
rect 439 2461 443 2462
rect 112 2434 114 2461
rect 136 2437 138 2461
rect 312 2437 314 2461
rect 134 2436 140 2437
rect 110 2433 116 2434
rect 110 2429 111 2433
rect 115 2429 116 2433
rect 134 2432 135 2436
rect 139 2432 140 2436
rect 134 2431 140 2432
rect 310 2436 316 2437
rect 310 2432 311 2436
rect 315 2432 316 2436
rect 310 2431 316 2432
rect 110 2428 116 2429
rect 480 2428 482 2534
rect 608 2520 610 2541
rect 620 2540 622 2582
rect 632 2560 634 2582
rect 710 2577 716 2578
rect 710 2573 711 2577
rect 715 2573 716 2577
rect 710 2572 716 2573
rect 630 2559 636 2560
rect 630 2555 631 2559
rect 635 2555 636 2559
rect 630 2554 636 2555
rect 712 2547 714 2572
rect 752 2560 754 2662
rect 766 2656 772 2657
rect 766 2652 767 2656
rect 771 2652 772 2656
rect 766 2651 772 2652
rect 768 2627 770 2651
rect 767 2626 771 2627
rect 767 2621 771 2622
rect 863 2626 867 2627
rect 863 2621 867 2622
rect 864 2597 866 2621
rect 862 2596 868 2597
rect 862 2592 863 2596
rect 867 2592 868 2596
rect 862 2591 868 2592
rect 862 2577 868 2578
rect 862 2573 863 2577
rect 867 2573 868 2577
rect 862 2572 868 2573
rect 750 2559 756 2560
rect 750 2555 751 2559
rect 755 2555 756 2559
rect 750 2554 756 2555
rect 864 2547 866 2572
rect 880 2560 882 2662
rect 2006 2659 2012 2660
rect 886 2656 892 2657
rect 886 2652 887 2656
rect 891 2652 892 2656
rect 886 2651 892 2652
rect 998 2656 1004 2657
rect 998 2652 999 2656
rect 1003 2652 1004 2656
rect 998 2651 1004 2652
rect 1110 2656 1116 2657
rect 1110 2652 1111 2656
rect 1115 2652 1116 2656
rect 1110 2651 1116 2652
rect 1230 2656 1236 2657
rect 1230 2652 1231 2656
rect 1235 2652 1236 2656
rect 1230 2651 1236 2652
rect 1350 2656 1356 2657
rect 1350 2652 1351 2656
rect 1355 2652 1356 2656
rect 2006 2655 2007 2659
rect 2011 2655 2012 2659
rect 2048 2655 2050 2686
rect 2334 2684 2335 2688
rect 2339 2684 2340 2688
rect 2334 2683 2340 2684
rect 2336 2655 2338 2683
rect 2006 2654 2012 2655
rect 2047 2654 2051 2655
rect 1350 2651 1356 2652
rect 888 2627 890 2651
rect 1000 2627 1002 2651
rect 1112 2627 1114 2651
rect 1232 2627 1234 2651
rect 1352 2627 1354 2651
rect 2008 2627 2010 2654
rect 2047 2649 2051 2650
rect 2127 2654 2131 2655
rect 2127 2649 2131 2650
rect 2279 2654 2283 2655
rect 2279 2649 2283 2650
rect 2335 2654 2339 2655
rect 2335 2649 2339 2650
rect 887 2626 891 2627
rect 887 2621 891 2622
rect 999 2626 1003 2627
rect 999 2621 1003 2622
rect 1007 2626 1011 2627
rect 1007 2621 1011 2622
rect 1111 2626 1115 2627
rect 1111 2621 1115 2622
rect 1143 2626 1147 2627
rect 1143 2621 1147 2622
rect 1231 2626 1235 2627
rect 1231 2621 1235 2622
rect 1279 2626 1283 2627
rect 1279 2621 1283 2622
rect 1351 2626 1355 2627
rect 1351 2621 1355 2622
rect 1423 2626 1427 2627
rect 1423 2621 1427 2622
rect 2007 2626 2011 2627
rect 2048 2622 2050 2649
rect 2128 2625 2130 2649
rect 2280 2625 2282 2649
rect 2404 2632 2406 2722
rect 2412 2700 2414 2722
rect 2496 2708 2498 2729
rect 2664 2708 2666 2729
rect 2738 2727 2744 2728
rect 2738 2723 2739 2727
rect 2743 2723 2744 2727
rect 2738 2722 2744 2723
rect 2494 2707 2500 2708
rect 2494 2703 2495 2707
rect 2499 2703 2500 2707
rect 2494 2702 2500 2703
rect 2662 2707 2668 2708
rect 2662 2703 2663 2707
rect 2667 2703 2668 2707
rect 2662 2702 2668 2703
rect 2740 2700 2742 2722
rect 2832 2708 2834 2729
rect 3000 2708 3002 2729
rect 3074 2727 3080 2728
rect 3074 2723 3075 2727
rect 3079 2723 3080 2727
rect 3074 2722 3080 2723
rect 2830 2707 2836 2708
rect 2830 2703 2831 2707
rect 2835 2703 2836 2707
rect 2830 2702 2836 2703
rect 2998 2707 3004 2708
rect 2998 2703 2999 2707
rect 3003 2703 3004 2707
rect 2998 2702 3004 2703
rect 3076 2700 3078 2722
rect 3168 2708 3170 2729
rect 3324 2728 3326 2774
rect 3390 2769 3396 2770
rect 3390 2765 3391 2769
rect 3395 2765 3396 2769
rect 3390 2764 3396 2765
rect 3392 2735 3394 2764
rect 3476 2752 3478 2774
rect 3542 2769 3548 2770
rect 3542 2765 3543 2769
rect 3547 2765 3548 2769
rect 3542 2764 3548 2765
rect 3474 2751 3480 2752
rect 3474 2747 3475 2751
rect 3479 2747 3480 2751
rect 3474 2746 3480 2747
rect 3544 2735 3546 2764
rect 3632 2752 3634 2774
rect 3702 2769 3708 2770
rect 3702 2765 3703 2769
rect 3707 2765 3708 2769
rect 3702 2764 3708 2765
rect 3838 2769 3844 2770
rect 3838 2765 3839 2769
rect 3843 2765 3844 2769
rect 3838 2764 3844 2765
rect 3630 2751 3636 2752
rect 3630 2747 3631 2751
rect 3635 2747 3636 2751
rect 3630 2746 3636 2747
rect 3704 2735 3706 2764
rect 3762 2747 3768 2748
rect 3762 2743 3763 2747
rect 3767 2743 3768 2747
rect 3762 2742 3768 2743
rect 3335 2734 3339 2735
rect 3335 2729 3339 2730
rect 3391 2734 3395 2735
rect 3391 2729 3395 2730
rect 3511 2734 3515 2735
rect 3511 2729 3515 2730
rect 3543 2734 3547 2735
rect 3543 2729 3547 2730
rect 3687 2734 3691 2735
rect 3687 2729 3691 2730
rect 3703 2734 3707 2735
rect 3703 2729 3707 2730
rect 3322 2727 3328 2728
rect 3322 2723 3323 2727
rect 3327 2723 3328 2727
rect 3322 2722 3328 2723
rect 3258 2719 3264 2720
rect 3258 2715 3259 2719
rect 3263 2715 3264 2719
rect 3258 2714 3264 2715
rect 3166 2707 3172 2708
rect 3166 2703 3167 2707
rect 3171 2703 3172 2707
rect 3166 2702 3172 2703
rect 3260 2700 3262 2714
rect 3336 2708 3338 2729
rect 3512 2708 3514 2729
rect 3578 2727 3584 2728
rect 3578 2723 3579 2727
rect 3583 2723 3584 2727
rect 3578 2722 3584 2723
rect 3586 2727 3592 2728
rect 3586 2723 3587 2727
rect 3591 2723 3592 2727
rect 3586 2722 3592 2723
rect 3334 2707 3340 2708
rect 3334 2703 3335 2707
rect 3339 2703 3340 2707
rect 3334 2702 3340 2703
rect 3510 2707 3516 2708
rect 3510 2703 3511 2707
rect 3515 2703 3516 2707
rect 3510 2702 3516 2703
rect 2410 2699 2416 2700
rect 2410 2695 2411 2699
rect 2415 2695 2416 2699
rect 2410 2694 2416 2695
rect 2738 2699 2744 2700
rect 2738 2695 2739 2699
rect 2743 2695 2744 2699
rect 2738 2694 2744 2695
rect 3074 2699 3080 2700
rect 3074 2695 3075 2699
rect 3079 2695 3080 2699
rect 3258 2699 3264 2700
rect 3074 2694 3080 2695
rect 3242 2695 3248 2696
rect 3242 2691 3243 2695
rect 3247 2691 3248 2695
rect 3258 2695 3259 2699
rect 3263 2695 3264 2699
rect 3258 2694 3264 2695
rect 3242 2690 3248 2691
rect 3580 2691 3582 2722
rect 3588 2700 3590 2722
rect 3688 2708 3690 2729
rect 3686 2707 3692 2708
rect 3686 2703 3687 2707
rect 3691 2703 3692 2707
rect 3686 2702 3692 2703
rect 3764 2700 3766 2742
rect 3840 2735 3842 2764
rect 3839 2734 3843 2735
rect 3839 2729 3843 2730
rect 3840 2708 3842 2729
rect 3908 2728 3910 2774
rect 3916 2752 3918 2942
rect 3942 2936 3948 2937
rect 3942 2932 3943 2936
rect 3947 2932 3948 2936
rect 3942 2931 3948 2932
rect 3944 2895 3946 2931
rect 3943 2894 3947 2895
rect 3943 2889 3947 2890
rect 3944 2869 3946 2889
rect 3942 2868 3948 2869
rect 3942 2864 3943 2868
rect 3947 2864 3948 2868
rect 3942 2863 3948 2864
rect 3942 2851 3948 2852
rect 3942 2847 3943 2851
rect 3947 2847 3948 2851
rect 3942 2846 3948 2847
rect 3944 2819 3946 2846
rect 3943 2818 3947 2819
rect 3943 2813 3947 2814
rect 3944 2786 3946 2813
rect 3942 2785 3948 2786
rect 3942 2781 3943 2785
rect 3947 2781 3948 2785
rect 3942 2780 3948 2781
rect 3942 2768 3948 2769
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 3942 2763 3948 2764
rect 3914 2751 3920 2752
rect 3914 2747 3915 2751
rect 3919 2747 3920 2751
rect 3914 2746 3920 2747
rect 3944 2735 3946 2763
rect 3943 2734 3947 2735
rect 3943 2729 3947 2730
rect 3906 2727 3912 2728
rect 3906 2723 3907 2727
rect 3911 2723 3912 2727
rect 3906 2722 3912 2723
rect 3944 2709 3946 2729
rect 3942 2708 3948 2709
rect 3838 2707 3844 2708
rect 3838 2703 3839 2707
rect 3843 2703 3844 2707
rect 3942 2704 3943 2708
rect 3947 2704 3948 2708
rect 3942 2703 3948 2704
rect 3838 2702 3844 2703
rect 3586 2699 3592 2700
rect 3586 2695 3587 2699
rect 3591 2695 3592 2699
rect 3586 2694 3592 2695
rect 3762 2699 3768 2700
rect 3762 2695 3763 2699
rect 3767 2695 3768 2699
rect 3762 2694 3768 2695
rect 3906 2691 3912 2692
rect 2494 2688 2500 2689
rect 2494 2684 2495 2688
rect 2499 2684 2500 2688
rect 2494 2683 2500 2684
rect 2662 2688 2668 2689
rect 2662 2684 2663 2688
rect 2667 2684 2668 2688
rect 2662 2683 2668 2684
rect 2830 2688 2836 2689
rect 2830 2684 2831 2688
rect 2835 2684 2836 2688
rect 2830 2683 2836 2684
rect 2998 2688 3004 2689
rect 2998 2684 2999 2688
rect 3003 2684 3004 2688
rect 2998 2683 3004 2684
rect 3166 2688 3172 2689
rect 3166 2684 3167 2688
rect 3171 2684 3172 2688
rect 3166 2683 3172 2684
rect 2496 2655 2498 2683
rect 2664 2655 2666 2683
rect 2832 2655 2834 2683
rect 3000 2655 3002 2683
rect 3168 2655 3170 2683
rect 2447 2654 2451 2655
rect 2447 2649 2451 2650
rect 2495 2654 2499 2655
rect 2495 2649 2499 2650
rect 2623 2654 2627 2655
rect 2623 2649 2627 2650
rect 2663 2654 2667 2655
rect 2663 2649 2667 2650
rect 2807 2654 2811 2655
rect 2807 2649 2811 2650
rect 2831 2654 2835 2655
rect 2831 2649 2835 2650
rect 2991 2654 2995 2655
rect 2991 2649 2995 2650
rect 2999 2654 3003 2655
rect 2999 2649 3003 2650
rect 3167 2654 3171 2655
rect 3167 2649 3171 2650
rect 3175 2654 3179 2655
rect 3175 2649 3179 2650
rect 2402 2631 2408 2632
rect 2402 2627 2403 2631
rect 2407 2627 2408 2631
rect 2402 2626 2408 2627
rect 2448 2625 2450 2649
rect 2624 2625 2626 2649
rect 2808 2625 2810 2649
rect 2992 2625 2994 2649
rect 3176 2625 3178 2649
rect 2126 2624 2132 2625
rect 2007 2621 2011 2622
rect 2046 2621 2052 2622
rect 1008 2597 1010 2621
rect 1144 2597 1146 2621
rect 1280 2597 1282 2621
rect 1424 2597 1426 2621
rect 1006 2596 1012 2597
rect 1006 2592 1007 2596
rect 1011 2592 1012 2596
rect 1006 2591 1012 2592
rect 1142 2596 1148 2597
rect 1142 2592 1143 2596
rect 1147 2592 1148 2596
rect 1142 2591 1148 2592
rect 1278 2596 1284 2597
rect 1278 2592 1279 2596
rect 1283 2592 1284 2596
rect 1278 2591 1284 2592
rect 1422 2596 1428 2597
rect 1422 2592 1423 2596
rect 1427 2592 1428 2596
rect 2008 2594 2010 2621
rect 2046 2617 2047 2621
rect 2051 2617 2052 2621
rect 2126 2620 2127 2624
rect 2131 2620 2132 2624
rect 2126 2619 2132 2620
rect 2278 2624 2284 2625
rect 2278 2620 2279 2624
rect 2283 2620 2284 2624
rect 2278 2619 2284 2620
rect 2446 2624 2452 2625
rect 2446 2620 2447 2624
rect 2451 2620 2452 2624
rect 2446 2619 2452 2620
rect 2622 2624 2628 2625
rect 2622 2620 2623 2624
rect 2627 2620 2628 2624
rect 2622 2619 2628 2620
rect 2806 2624 2812 2625
rect 2806 2620 2807 2624
rect 2811 2620 2812 2624
rect 2806 2619 2812 2620
rect 2990 2624 2996 2625
rect 2990 2620 2991 2624
rect 2995 2620 2996 2624
rect 2990 2619 2996 2620
rect 3174 2624 3180 2625
rect 3174 2620 3175 2624
rect 3179 2620 3180 2624
rect 3174 2619 3180 2620
rect 2046 2616 2052 2617
rect 2202 2615 2208 2616
rect 2202 2611 2203 2615
rect 2207 2611 2208 2615
rect 2202 2610 2208 2611
rect 2354 2615 2360 2616
rect 2354 2611 2355 2615
rect 2359 2611 2360 2615
rect 2354 2610 2360 2611
rect 2522 2615 2528 2616
rect 2522 2611 2523 2615
rect 2527 2611 2528 2615
rect 2522 2610 2528 2611
rect 2698 2615 2704 2616
rect 2698 2611 2699 2615
rect 2703 2611 2704 2615
rect 2698 2610 2704 2611
rect 2890 2615 2896 2616
rect 2890 2611 2891 2615
rect 2895 2611 2896 2615
rect 2890 2610 2896 2611
rect 3102 2615 3108 2616
rect 3102 2611 3103 2615
rect 3107 2611 3108 2615
rect 3102 2610 3108 2611
rect 2126 2605 2132 2606
rect 2046 2604 2052 2605
rect 2046 2600 2047 2604
rect 2051 2600 2052 2604
rect 2126 2601 2127 2605
rect 2131 2601 2132 2605
rect 2126 2600 2132 2601
rect 2046 2599 2052 2600
rect 1422 2591 1428 2592
rect 2006 2593 2012 2594
rect 2006 2589 2007 2593
rect 2011 2589 2012 2593
rect 2006 2588 2012 2589
rect 938 2587 944 2588
rect 938 2583 939 2587
rect 943 2583 944 2587
rect 938 2582 944 2583
rect 1082 2587 1088 2588
rect 1082 2583 1083 2587
rect 1087 2583 1088 2587
rect 1082 2582 1088 2583
rect 1218 2587 1224 2588
rect 1218 2583 1219 2587
rect 1223 2583 1224 2587
rect 1218 2582 1224 2583
rect 1354 2587 1360 2588
rect 1354 2583 1355 2587
rect 1359 2583 1360 2587
rect 1354 2582 1360 2583
rect 1366 2587 1372 2588
rect 1366 2583 1367 2587
rect 1371 2583 1372 2587
rect 1366 2582 1372 2583
rect 940 2560 942 2582
rect 1006 2577 1012 2578
rect 1006 2573 1007 2577
rect 1011 2573 1012 2577
rect 1006 2572 1012 2573
rect 878 2559 884 2560
rect 878 2555 879 2559
rect 883 2555 884 2559
rect 878 2554 884 2555
rect 938 2559 944 2560
rect 938 2555 939 2559
rect 943 2555 944 2559
rect 938 2554 944 2555
rect 1008 2547 1010 2572
rect 1084 2560 1086 2582
rect 1142 2577 1148 2578
rect 1142 2573 1143 2577
rect 1147 2573 1148 2577
rect 1142 2572 1148 2573
rect 1082 2559 1088 2560
rect 1082 2555 1083 2559
rect 1087 2555 1088 2559
rect 1082 2554 1088 2555
rect 1144 2547 1146 2572
rect 1220 2560 1222 2582
rect 1278 2577 1284 2578
rect 1278 2573 1279 2577
rect 1283 2573 1284 2577
rect 1278 2572 1284 2573
rect 1218 2559 1224 2560
rect 1218 2555 1219 2559
rect 1223 2555 1224 2559
rect 1218 2554 1224 2555
rect 1280 2547 1282 2572
rect 1356 2560 1358 2582
rect 1354 2559 1360 2560
rect 1354 2555 1355 2559
rect 1359 2555 1360 2559
rect 1354 2554 1360 2555
rect 1368 2548 1370 2582
rect 1422 2577 1428 2578
rect 1422 2573 1423 2577
rect 1427 2573 1428 2577
rect 1422 2572 1428 2573
rect 2006 2576 2012 2577
rect 2006 2572 2007 2576
rect 2011 2572 2012 2576
rect 1366 2547 1372 2548
rect 1424 2547 1426 2572
rect 2006 2571 2012 2572
rect 2048 2571 2050 2599
rect 2128 2571 2130 2600
rect 2204 2588 2206 2610
rect 2278 2605 2284 2606
rect 2278 2601 2279 2605
rect 2283 2601 2284 2605
rect 2278 2600 2284 2601
rect 2202 2587 2208 2588
rect 2166 2583 2172 2584
rect 2166 2578 2167 2583
rect 2171 2578 2172 2583
rect 2202 2583 2203 2587
rect 2207 2583 2208 2587
rect 2202 2582 2208 2583
rect 2167 2575 2171 2576
rect 2280 2571 2282 2600
rect 2356 2588 2358 2610
rect 2446 2605 2452 2606
rect 2446 2601 2447 2605
rect 2451 2601 2452 2605
rect 2446 2600 2452 2601
rect 2354 2587 2360 2588
rect 2354 2583 2355 2587
rect 2359 2583 2360 2587
rect 2354 2582 2360 2583
rect 2448 2571 2450 2600
rect 2524 2588 2526 2610
rect 2622 2605 2628 2606
rect 2622 2601 2623 2605
rect 2627 2601 2628 2605
rect 2622 2600 2628 2601
rect 2522 2587 2528 2588
rect 2522 2583 2523 2587
rect 2527 2583 2528 2587
rect 2522 2582 2528 2583
rect 2599 2580 2603 2581
rect 2599 2575 2603 2576
rect 2008 2547 2010 2571
rect 2047 2570 2051 2571
rect 2047 2565 2051 2566
rect 2071 2570 2075 2571
rect 2071 2565 2075 2566
rect 2127 2570 2131 2571
rect 2127 2565 2131 2566
rect 2183 2570 2187 2571
rect 2183 2565 2187 2566
rect 2279 2570 2283 2571
rect 2279 2565 2283 2566
rect 2319 2570 2323 2571
rect 2319 2565 2323 2566
rect 2447 2570 2451 2571
rect 2447 2565 2451 2566
rect 2471 2570 2475 2571
rect 2471 2565 2475 2566
rect 711 2546 715 2547
rect 711 2541 715 2542
rect 775 2546 779 2547
rect 775 2541 779 2542
rect 863 2546 867 2547
rect 863 2541 867 2542
rect 927 2546 931 2547
rect 927 2541 931 2542
rect 1007 2546 1011 2547
rect 1007 2541 1011 2542
rect 1079 2546 1083 2547
rect 1079 2541 1083 2542
rect 1143 2546 1147 2547
rect 1143 2541 1147 2542
rect 1223 2546 1227 2547
rect 1223 2541 1227 2542
rect 1279 2546 1283 2547
rect 1279 2541 1283 2542
rect 1359 2546 1363 2547
rect 1366 2543 1367 2547
rect 1371 2543 1372 2547
rect 1366 2542 1372 2543
rect 1423 2546 1427 2547
rect 1359 2541 1363 2542
rect 1423 2541 1427 2542
rect 1495 2546 1499 2547
rect 1495 2541 1499 2542
rect 1639 2546 1643 2547
rect 1639 2541 1643 2542
rect 2007 2546 2011 2547
rect 2048 2545 2050 2565
rect 2007 2541 2011 2542
rect 2046 2544 2052 2545
rect 2072 2544 2074 2565
rect 2146 2563 2152 2564
rect 2146 2559 2147 2563
rect 2151 2559 2152 2563
rect 2146 2558 2152 2559
rect 618 2539 624 2540
rect 618 2535 619 2539
rect 623 2535 624 2539
rect 618 2534 624 2535
rect 682 2539 688 2540
rect 682 2535 683 2539
rect 687 2535 688 2539
rect 682 2534 688 2535
rect 606 2519 612 2520
rect 606 2515 607 2519
rect 611 2515 612 2519
rect 606 2514 612 2515
rect 684 2512 686 2534
rect 776 2520 778 2541
rect 850 2539 856 2540
rect 850 2535 851 2539
rect 855 2535 856 2539
rect 850 2534 856 2535
rect 774 2519 780 2520
rect 774 2515 775 2519
rect 779 2515 780 2519
rect 774 2514 780 2515
rect 852 2512 854 2534
rect 928 2520 930 2541
rect 1080 2520 1082 2541
rect 1154 2539 1160 2540
rect 1154 2535 1155 2539
rect 1159 2535 1160 2539
rect 1154 2534 1160 2535
rect 926 2519 932 2520
rect 926 2515 927 2519
rect 931 2515 932 2519
rect 926 2514 932 2515
rect 1078 2519 1084 2520
rect 1078 2515 1079 2519
rect 1083 2515 1084 2519
rect 1078 2514 1084 2515
rect 1156 2512 1158 2534
rect 1224 2520 1226 2541
rect 1298 2539 1304 2540
rect 1298 2535 1299 2539
rect 1303 2535 1304 2539
rect 1298 2534 1304 2535
rect 1222 2519 1228 2520
rect 1222 2515 1223 2519
rect 1227 2515 1228 2519
rect 1222 2514 1228 2515
rect 1300 2512 1302 2534
rect 1360 2520 1362 2541
rect 1434 2539 1440 2540
rect 1434 2535 1435 2539
rect 1439 2535 1440 2539
rect 1434 2534 1440 2535
rect 1358 2519 1364 2520
rect 1358 2515 1359 2519
rect 1363 2515 1364 2519
rect 1358 2514 1364 2515
rect 1436 2512 1438 2534
rect 1496 2520 1498 2541
rect 1570 2539 1576 2540
rect 1570 2535 1571 2539
rect 1575 2535 1576 2539
rect 1570 2534 1576 2535
rect 1494 2519 1500 2520
rect 1494 2515 1495 2519
rect 1499 2515 1500 2519
rect 1494 2514 1500 2515
rect 1572 2512 1574 2534
rect 1640 2520 1642 2541
rect 2008 2521 2010 2541
rect 2046 2540 2047 2544
rect 2051 2540 2052 2544
rect 2046 2539 2052 2540
rect 2070 2543 2076 2544
rect 2070 2539 2071 2543
rect 2075 2539 2076 2543
rect 2070 2538 2076 2539
rect 2148 2536 2150 2558
rect 2184 2544 2186 2565
rect 2258 2563 2264 2564
rect 2258 2559 2259 2563
rect 2263 2559 2264 2563
rect 2258 2558 2264 2559
rect 2182 2543 2188 2544
rect 2182 2539 2183 2543
rect 2187 2539 2188 2543
rect 2182 2538 2188 2539
rect 2260 2536 2262 2558
rect 2298 2555 2304 2556
rect 2298 2551 2299 2555
rect 2303 2551 2304 2555
rect 2298 2550 2304 2551
rect 2146 2535 2152 2536
rect 2146 2531 2147 2535
rect 2151 2531 2152 2535
rect 2146 2530 2152 2531
rect 2258 2535 2264 2536
rect 2258 2531 2259 2535
rect 2263 2531 2264 2535
rect 2258 2530 2264 2531
rect 2046 2527 2052 2528
rect 2046 2523 2047 2527
rect 2051 2523 2052 2527
rect 2046 2522 2052 2523
rect 2070 2524 2076 2525
rect 2006 2520 2012 2521
rect 1638 2519 1644 2520
rect 1638 2515 1639 2519
rect 1643 2515 1644 2519
rect 2006 2516 2007 2520
rect 2011 2516 2012 2520
rect 2006 2515 2012 2516
rect 1638 2514 1644 2515
rect 682 2511 688 2512
rect 682 2507 683 2511
rect 687 2507 688 2511
rect 682 2506 688 2507
rect 850 2511 856 2512
rect 850 2507 851 2511
rect 855 2507 856 2511
rect 1154 2511 1160 2512
rect 850 2506 856 2507
rect 1002 2507 1008 2508
rect 1002 2503 1003 2507
rect 1007 2503 1008 2507
rect 1154 2507 1155 2511
rect 1159 2507 1160 2511
rect 1154 2506 1160 2507
rect 1298 2511 1304 2512
rect 1298 2507 1299 2511
rect 1303 2507 1304 2511
rect 1298 2506 1304 2507
rect 1434 2511 1440 2512
rect 1434 2507 1435 2511
rect 1439 2507 1440 2511
rect 1434 2506 1440 2507
rect 1570 2511 1576 2512
rect 1570 2507 1571 2511
rect 1575 2507 1576 2511
rect 1570 2506 1576 2507
rect 1578 2511 1584 2512
rect 1578 2507 1579 2511
rect 1583 2507 1584 2511
rect 1578 2506 1584 2507
rect 1002 2502 1008 2503
rect 606 2500 612 2501
rect 606 2496 607 2500
rect 611 2496 612 2500
rect 606 2495 612 2496
rect 774 2500 780 2501
rect 774 2496 775 2500
rect 779 2496 780 2500
rect 774 2495 780 2496
rect 926 2500 932 2501
rect 926 2496 927 2500
rect 931 2496 932 2500
rect 926 2495 932 2496
rect 608 2467 610 2495
rect 776 2467 778 2495
rect 928 2467 930 2495
rect 511 2466 515 2467
rect 511 2461 515 2462
rect 607 2466 611 2467
rect 607 2461 611 2462
rect 711 2466 715 2467
rect 711 2461 715 2462
rect 775 2466 779 2467
rect 775 2461 779 2462
rect 903 2466 907 2467
rect 903 2461 907 2462
rect 927 2466 931 2467
rect 927 2461 931 2462
rect 512 2437 514 2461
rect 712 2437 714 2461
rect 904 2437 906 2461
rect 510 2436 516 2437
rect 510 2432 511 2436
rect 515 2432 516 2436
rect 510 2431 516 2432
rect 710 2436 716 2437
rect 710 2432 711 2436
rect 715 2432 716 2436
rect 710 2431 716 2432
rect 902 2436 908 2437
rect 902 2432 903 2436
rect 907 2432 908 2436
rect 902 2431 908 2432
rect 210 2427 216 2428
rect 210 2423 211 2427
rect 215 2423 216 2427
rect 210 2422 216 2423
rect 386 2427 392 2428
rect 386 2423 387 2427
rect 391 2423 392 2427
rect 386 2422 392 2423
rect 478 2427 484 2428
rect 478 2423 479 2427
rect 483 2423 484 2427
rect 478 2422 484 2423
rect 618 2427 624 2428
rect 618 2423 619 2427
rect 623 2423 624 2427
rect 618 2422 624 2423
rect 846 2427 852 2428
rect 846 2423 847 2427
rect 851 2423 852 2427
rect 846 2422 852 2423
rect 134 2417 140 2418
rect 110 2416 116 2417
rect 110 2412 111 2416
rect 115 2412 116 2416
rect 134 2413 135 2417
rect 139 2413 140 2417
rect 134 2412 140 2413
rect 110 2411 116 2412
rect 112 2391 114 2411
rect 136 2391 138 2412
rect 212 2400 214 2422
rect 310 2417 316 2418
rect 310 2413 311 2417
rect 315 2413 316 2417
rect 310 2412 316 2413
rect 210 2399 216 2400
rect 210 2395 211 2399
rect 215 2395 216 2399
rect 210 2394 216 2395
rect 210 2391 216 2392
rect 312 2391 314 2412
rect 388 2400 390 2422
rect 510 2417 516 2418
rect 510 2413 511 2417
rect 515 2413 516 2417
rect 510 2412 516 2413
rect 386 2399 392 2400
rect 386 2395 387 2399
rect 391 2395 392 2399
rect 386 2394 392 2395
rect 512 2391 514 2412
rect 111 2390 115 2391
rect 111 2385 115 2386
rect 135 2390 139 2391
rect 210 2387 211 2391
rect 215 2387 216 2391
rect 210 2386 216 2387
rect 311 2390 315 2391
rect 135 2385 139 2386
rect 112 2365 114 2385
rect 110 2364 116 2365
rect 136 2364 138 2385
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 110 2359 116 2360
rect 134 2363 140 2364
rect 134 2359 135 2363
rect 139 2359 140 2363
rect 134 2358 140 2359
rect 212 2356 214 2386
rect 311 2385 315 2386
rect 327 2390 331 2391
rect 327 2385 331 2386
rect 511 2390 515 2391
rect 511 2385 515 2386
rect 551 2390 555 2391
rect 551 2385 555 2386
rect 246 2383 252 2384
rect 246 2379 247 2383
rect 251 2379 252 2383
rect 246 2378 252 2379
rect 248 2356 250 2378
rect 328 2364 330 2385
rect 346 2383 352 2384
rect 346 2379 347 2383
rect 351 2379 352 2383
rect 346 2378 352 2379
rect 326 2363 332 2364
rect 326 2359 327 2363
rect 331 2359 332 2363
rect 326 2358 332 2359
rect 210 2355 216 2356
rect 210 2351 211 2355
rect 215 2351 216 2355
rect 210 2350 216 2351
rect 246 2355 252 2356
rect 246 2351 247 2355
rect 251 2351 252 2355
rect 246 2350 252 2351
rect 110 2347 116 2348
rect 110 2343 111 2347
rect 115 2343 116 2347
rect 110 2342 116 2343
rect 134 2344 140 2345
rect 112 2307 114 2342
rect 134 2340 135 2344
rect 139 2340 140 2344
rect 134 2339 140 2340
rect 326 2344 332 2345
rect 326 2340 327 2344
rect 331 2340 332 2344
rect 326 2339 332 2340
rect 136 2307 138 2339
rect 328 2307 330 2339
rect 111 2306 115 2307
rect 111 2301 115 2302
rect 135 2306 139 2307
rect 135 2301 139 2302
rect 271 2306 275 2307
rect 271 2301 275 2302
rect 327 2306 331 2307
rect 327 2301 331 2302
rect 112 2274 114 2301
rect 136 2277 138 2301
rect 272 2277 274 2301
rect 134 2276 140 2277
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 134 2272 135 2276
rect 139 2272 140 2276
rect 134 2271 140 2272
rect 270 2276 276 2277
rect 270 2272 271 2276
rect 275 2272 276 2276
rect 270 2271 276 2272
rect 110 2268 116 2269
rect 348 2268 350 2378
rect 552 2364 554 2385
rect 620 2384 622 2422
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 712 2391 714 2412
rect 848 2400 850 2422
rect 902 2417 908 2418
rect 902 2413 903 2417
rect 907 2413 908 2417
rect 902 2412 908 2413
rect 846 2399 852 2400
rect 846 2395 847 2399
rect 851 2395 852 2399
rect 846 2394 852 2395
rect 904 2391 906 2412
rect 1004 2400 1006 2502
rect 1078 2500 1084 2501
rect 1078 2496 1079 2500
rect 1083 2496 1084 2500
rect 1078 2495 1084 2496
rect 1222 2500 1228 2501
rect 1222 2496 1223 2500
rect 1227 2496 1228 2500
rect 1222 2495 1228 2496
rect 1358 2500 1364 2501
rect 1358 2496 1359 2500
rect 1363 2496 1364 2500
rect 1358 2495 1364 2496
rect 1494 2500 1500 2501
rect 1494 2496 1495 2500
rect 1499 2496 1500 2500
rect 1494 2495 1500 2496
rect 1080 2467 1082 2495
rect 1224 2467 1226 2495
rect 1360 2467 1362 2495
rect 1496 2467 1498 2495
rect 1079 2466 1083 2467
rect 1079 2461 1083 2462
rect 1223 2466 1227 2467
rect 1223 2461 1227 2462
rect 1239 2466 1243 2467
rect 1239 2461 1243 2462
rect 1359 2466 1363 2467
rect 1359 2461 1363 2462
rect 1391 2466 1395 2467
rect 1391 2461 1395 2462
rect 1495 2466 1499 2467
rect 1495 2461 1499 2462
rect 1527 2466 1531 2467
rect 1527 2461 1531 2462
rect 1080 2437 1082 2461
rect 1240 2437 1242 2461
rect 1392 2437 1394 2461
rect 1528 2437 1530 2461
rect 1078 2436 1084 2437
rect 1078 2432 1079 2436
rect 1083 2432 1084 2436
rect 1078 2431 1084 2432
rect 1238 2436 1244 2437
rect 1238 2432 1239 2436
rect 1243 2432 1244 2436
rect 1238 2431 1244 2432
rect 1390 2436 1396 2437
rect 1390 2432 1391 2436
rect 1395 2432 1396 2436
rect 1390 2431 1396 2432
rect 1526 2436 1532 2437
rect 1526 2432 1527 2436
rect 1531 2432 1532 2436
rect 1526 2431 1532 2432
rect 1154 2427 1160 2428
rect 1154 2423 1155 2427
rect 1159 2423 1160 2427
rect 1154 2422 1160 2423
rect 1314 2427 1320 2428
rect 1314 2423 1315 2427
rect 1319 2423 1320 2427
rect 1314 2422 1320 2423
rect 1466 2427 1472 2428
rect 1466 2423 1467 2427
rect 1471 2423 1472 2427
rect 1466 2422 1472 2423
rect 1474 2427 1480 2428
rect 1474 2423 1475 2427
rect 1479 2423 1480 2427
rect 1474 2422 1480 2423
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1002 2399 1008 2400
rect 1002 2395 1003 2399
rect 1007 2395 1008 2399
rect 1002 2394 1008 2395
rect 1080 2391 1082 2412
rect 1156 2400 1158 2422
rect 1238 2417 1244 2418
rect 1238 2413 1239 2417
rect 1243 2413 1244 2417
rect 1238 2412 1244 2413
rect 1154 2399 1160 2400
rect 1154 2395 1155 2399
rect 1159 2395 1160 2399
rect 1154 2394 1160 2395
rect 1240 2391 1242 2412
rect 1316 2400 1318 2422
rect 1390 2417 1396 2418
rect 1390 2413 1391 2417
rect 1395 2413 1396 2417
rect 1390 2412 1396 2413
rect 1314 2399 1320 2400
rect 1314 2395 1315 2399
rect 1319 2395 1320 2399
rect 1314 2394 1320 2395
rect 1392 2391 1394 2412
rect 1468 2400 1470 2422
rect 1466 2399 1472 2400
rect 1466 2395 1467 2399
rect 1471 2395 1472 2399
rect 1466 2394 1472 2395
rect 1476 2392 1478 2422
rect 1526 2417 1532 2418
rect 1526 2413 1527 2417
rect 1531 2413 1532 2417
rect 1526 2412 1532 2413
rect 1474 2391 1480 2392
rect 1528 2391 1530 2412
rect 1580 2408 1582 2506
rect 2006 2503 2012 2504
rect 1638 2500 1644 2501
rect 1638 2496 1639 2500
rect 1643 2496 1644 2500
rect 2006 2499 2007 2503
rect 2011 2499 2012 2503
rect 2006 2498 2012 2499
rect 1638 2495 1644 2496
rect 1640 2467 1642 2495
rect 2008 2467 2010 2498
rect 2048 2491 2050 2522
rect 2070 2520 2071 2524
rect 2075 2520 2076 2524
rect 2070 2519 2076 2520
rect 2182 2524 2188 2525
rect 2182 2520 2183 2524
rect 2187 2520 2188 2524
rect 2182 2519 2188 2520
rect 2072 2491 2074 2519
rect 2184 2491 2186 2519
rect 2047 2490 2051 2491
rect 2047 2485 2051 2486
rect 2071 2490 2075 2491
rect 2071 2485 2075 2486
rect 2183 2490 2187 2491
rect 2183 2485 2187 2486
rect 2215 2490 2219 2491
rect 2215 2485 2219 2486
rect 1639 2466 1643 2467
rect 1639 2461 1643 2462
rect 1663 2466 1667 2467
rect 1663 2461 1667 2462
rect 1791 2466 1795 2467
rect 1791 2461 1795 2462
rect 1903 2466 1907 2467
rect 1903 2461 1907 2462
rect 2007 2466 2011 2467
rect 2007 2461 2011 2462
rect 1664 2437 1666 2461
rect 1792 2437 1794 2461
rect 1904 2437 1906 2461
rect 1662 2436 1668 2437
rect 1662 2432 1663 2436
rect 1667 2432 1668 2436
rect 1662 2431 1668 2432
rect 1790 2436 1796 2437
rect 1790 2432 1791 2436
rect 1795 2432 1796 2436
rect 1790 2431 1796 2432
rect 1902 2436 1908 2437
rect 1902 2432 1903 2436
rect 1907 2432 1908 2436
rect 2008 2434 2010 2461
rect 2048 2458 2050 2485
rect 2072 2461 2074 2485
rect 2216 2461 2218 2485
rect 2070 2460 2076 2461
rect 2046 2457 2052 2458
rect 2046 2453 2047 2457
rect 2051 2453 2052 2457
rect 2070 2456 2071 2460
rect 2075 2456 2076 2460
rect 2070 2455 2076 2456
rect 2214 2460 2220 2461
rect 2214 2456 2215 2460
rect 2219 2456 2220 2460
rect 2214 2455 2220 2456
rect 2046 2452 2052 2453
rect 2300 2452 2302 2550
rect 2320 2544 2322 2565
rect 2394 2563 2400 2564
rect 2394 2559 2395 2563
rect 2399 2559 2400 2563
rect 2394 2558 2400 2559
rect 2318 2543 2324 2544
rect 2318 2539 2319 2543
rect 2323 2539 2324 2543
rect 2318 2538 2324 2539
rect 2396 2536 2398 2558
rect 2472 2544 2474 2565
rect 2546 2563 2552 2564
rect 2546 2559 2547 2563
rect 2551 2559 2552 2563
rect 2546 2558 2552 2559
rect 2470 2543 2476 2544
rect 2470 2539 2471 2543
rect 2475 2539 2476 2543
rect 2470 2538 2476 2539
rect 2548 2536 2550 2558
rect 2600 2536 2602 2575
rect 2624 2571 2626 2600
rect 2700 2588 2702 2610
rect 2806 2605 2812 2606
rect 2806 2601 2807 2605
rect 2811 2601 2812 2605
rect 2806 2600 2812 2601
rect 2698 2587 2704 2588
rect 2698 2583 2699 2587
rect 2703 2583 2704 2587
rect 2698 2582 2704 2583
rect 2808 2571 2810 2600
rect 2623 2570 2627 2571
rect 2623 2565 2627 2566
rect 2639 2570 2643 2571
rect 2639 2565 2643 2566
rect 2807 2570 2811 2571
rect 2807 2565 2811 2566
rect 2823 2570 2827 2571
rect 2823 2565 2827 2566
rect 2640 2544 2642 2565
rect 2824 2544 2826 2565
rect 2892 2564 2894 2610
rect 2990 2605 2996 2606
rect 2990 2601 2991 2605
rect 2995 2601 2996 2605
rect 2990 2600 2996 2601
rect 2992 2571 2994 2600
rect 3104 2588 3106 2610
rect 3174 2605 3180 2606
rect 3174 2601 3175 2605
rect 3179 2601 3180 2605
rect 3174 2600 3180 2601
rect 3102 2587 3108 2588
rect 3102 2583 3103 2587
rect 3107 2583 3108 2587
rect 3102 2582 3108 2583
rect 3176 2571 3178 2600
rect 3244 2588 3246 2690
rect 3580 2689 3590 2691
rect 3334 2688 3340 2689
rect 3334 2684 3335 2688
rect 3339 2684 3340 2688
rect 3334 2683 3340 2684
rect 3510 2688 3516 2689
rect 3510 2684 3511 2688
rect 3515 2684 3516 2688
rect 3510 2683 3516 2684
rect 3336 2655 3338 2683
rect 3512 2655 3514 2683
rect 3335 2654 3339 2655
rect 3335 2649 3339 2650
rect 3351 2654 3355 2655
rect 3351 2649 3355 2650
rect 3511 2654 3515 2655
rect 3511 2649 3515 2650
rect 3519 2654 3523 2655
rect 3519 2649 3523 2650
rect 3352 2625 3354 2649
rect 3520 2625 3522 2649
rect 3350 2624 3356 2625
rect 3350 2620 3351 2624
rect 3355 2620 3356 2624
rect 3350 2619 3356 2620
rect 3518 2624 3524 2625
rect 3518 2620 3519 2624
rect 3523 2620 3524 2624
rect 3518 2619 3524 2620
rect 3588 2616 3590 2689
rect 3686 2688 3692 2689
rect 3686 2684 3687 2688
rect 3691 2684 3692 2688
rect 3686 2683 3692 2684
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3906 2687 3907 2691
rect 3911 2687 3912 2691
rect 3906 2686 3912 2687
rect 3942 2691 3948 2692
rect 3942 2687 3943 2691
rect 3947 2687 3948 2691
rect 3942 2686 3948 2687
rect 3838 2683 3844 2684
rect 3688 2655 3690 2683
rect 3840 2655 3842 2683
rect 3687 2654 3691 2655
rect 3687 2649 3691 2650
rect 3839 2654 3843 2655
rect 3839 2649 3843 2650
rect 3688 2625 3690 2649
rect 3840 2625 3842 2649
rect 3686 2624 3692 2625
rect 3686 2620 3687 2624
rect 3691 2620 3692 2624
rect 3686 2619 3692 2620
rect 3838 2624 3844 2625
rect 3838 2620 3839 2624
rect 3843 2620 3844 2624
rect 3838 2619 3844 2620
rect 3426 2615 3432 2616
rect 3426 2611 3427 2615
rect 3431 2611 3432 2615
rect 3426 2610 3432 2611
rect 3586 2615 3592 2616
rect 3586 2611 3587 2615
rect 3591 2611 3592 2615
rect 3586 2610 3592 2611
rect 3618 2615 3624 2616
rect 3618 2611 3619 2615
rect 3623 2611 3624 2615
rect 3618 2610 3624 2611
rect 3350 2605 3356 2606
rect 3350 2601 3351 2605
rect 3355 2601 3356 2605
rect 3350 2600 3356 2601
rect 3242 2587 3248 2588
rect 3242 2583 3243 2587
rect 3247 2583 3248 2587
rect 3242 2582 3248 2583
rect 3352 2571 3354 2600
rect 3428 2588 3430 2610
rect 3518 2605 3524 2606
rect 3518 2601 3519 2605
rect 3523 2601 3524 2605
rect 3518 2600 3524 2601
rect 3426 2587 3432 2588
rect 3426 2583 3427 2587
rect 3431 2583 3432 2587
rect 3426 2582 3432 2583
rect 3520 2571 3522 2600
rect 3620 2596 3622 2610
rect 3686 2605 3692 2606
rect 3686 2601 3687 2605
rect 3691 2601 3692 2605
rect 3686 2600 3692 2601
rect 3838 2605 3844 2606
rect 3838 2601 3839 2605
rect 3843 2601 3844 2605
rect 3838 2600 3844 2601
rect 3618 2595 3624 2596
rect 3618 2591 3619 2595
rect 3623 2591 3624 2595
rect 3618 2590 3624 2591
rect 3688 2571 3690 2600
rect 3726 2583 3732 2584
rect 3726 2579 3727 2583
rect 3731 2579 3732 2583
rect 3726 2578 3732 2579
rect 2991 2570 2995 2571
rect 2991 2565 2995 2566
rect 3031 2570 3035 2571
rect 3031 2565 3035 2566
rect 3175 2570 3179 2571
rect 3175 2565 3179 2566
rect 3263 2570 3267 2571
rect 3263 2565 3267 2566
rect 3351 2570 3355 2571
rect 3351 2565 3355 2566
rect 3503 2570 3507 2571
rect 3503 2565 3507 2566
rect 3519 2570 3523 2571
rect 3519 2565 3523 2566
rect 3687 2570 3691 2571
rect 3687 2565 3691 2566
rect 2890 2563 2896 2564
rect 2890 2559 2891 2563
rect 2895 2559 2896 2563
rect 2890 2558 2896 2559
rect 2898 2563 2904 2564
rect 2898 2559 2899 2563
rect 2903 2559 2904 2563
rect 2898 2558 2904 2559
rect 2638 2543 2644 2544
rect 2638 2539 2639 2543
rect 2643 2539 2644 2543
rect 2638 2538 2644 2539
rect 2822 2543 2828 2544
rect 2822 2539 2823 2543
rect 2827 2539 2828 2543
rect 2822 2538 2828 2539
rect 2900 2536 2902 2558
rect 3032 2544 3034 2565
rect 3106 2563 3112 2564
rect 3106 2559 3107 2563
rect 3111 2559 3112 2563
rect 3106 2558 3112 2559
rect 3030 2543 3036 2544
rect 3030 2539 3031 2543
rect 3035 2539 3036 2543
rect 3030 2538 3036 2539
rect 3108 2536 3110 2558
rect 3264 2544 3266 2565
rect 3338 2563 3344 2564
rect 3338 2559 3339 2563
rect 3343 2559 3344 2563
rect 3338 2558 3344 2559
rect 3262 2543 3268 2544
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3340 2536 3342 2558
rect 3504 2544 3506 2565
rect 3698 2563 3704 2564
rect 3698 2559 3699 2563
rect 3703 2559 3704 2563
rect 3698 2558 3704 2559
rect 3502 2543 3508 2544
rect 3502 2539 3503 2543
rect 3507 2539 3508 2543
rect 3502 2538 3508 2539
rect 2394 2535 2400 2536
rect 2394 2531 2395 2535
rect 2399 2531 2400 2535
rect 2394 2530 2400 2531
rect 2546 2535 2552 2536
rect 2546 2531 2547 2535
rect 2551 2531 2552 2535
rect 2546 2530 2552 2531
rect 2598 2535 2604 2536
rect 2598 2531 2599 2535
rect 2603 2531 2604 2535
rect 2598 2530 2604 2531
rect 2898 2535 2904 2536
rect 2898 2531 2899 2535
rect 2903 2531 2904 2535
rect 2898 2530 2904 2531
rect 3106 2535 3112 2536
rect 3106 2531 3107 2535
rect 3111 2531 3112 2535
rect 3106 2530 3112 2531
rect 3338 2535 3344 2536
rect 3338 2531 3339 2535
rect 3343 2531 3344 2535
rect 3338 2530 3344 2531
rect 3450 2535 3456 2536
rect 3450 2531 3451 2535
rect 3455 2531 3456 2535
rect 3450 2530 3456 2531
rect 2318 2524 2324 2525
rect 2318 2520 2319 2524
rect 2323 2520 2324 2524
rect 2318 2519 2324 2520
rect 2470 2524 2476 2525
rect 2470 2520 2471 2524
rect 2475 2520 2476 2524
rect 2470 2519 2476 2520
rect 2638 2524 2644 2525
rect 2638 2520 2639 2524
rect 2643 2520 2644 2524
rect 2638 2519 2644 2520
rect 2822 2524 2828 2525
rect 2822 2520 2823 2524
rect 2827 2520 2828 2524
rect 2822 2519 2828 2520
rect 3030 2524 3036 2525
rect 3030 2520 3031 2524
rect 3035 2520 3036 2524
rect 3030 2519 3036 2520
rect 3262 2524 3268 2525
rect 3262 2520 3263 2524
rect 3267 2520 3268 2524
rect 3262 2519 3268 2520
rect 2320 2491 2322 2519
rect 2472 2491 2474 2519
rect 2640 2491 2642 2519
rect 2824 2491 2826 2519
rect 3032 2491 3034 2519
rect 3264 2491 3266 2519
rect 2319 2490 2323 2491
rect 2319 2485 2323 2486
rect 2383 2490 2387 2491
rect 2383 2485 2387 2486
rect 2471 2490 2475 2491
rect 2471 2485 2475 2486
rect 2559 2490 2563 2491
rect 2559 2485 2563 2486
rect 2639 2490 2643 2491
rect 2639 2485 2643 2486
rect 2751 2490 2755 2491
rect 2751 2485 2755 2486
rect 2823 2490 2827 2491
rect 2823 2485 2827 2486
rect 2951 2490 2955 2491
rect 2951 2485 2955 2486
rect 3031 2490 3035 2491
rect 3031 2485 3035 2486
rect 3167 2490 3171 2491
rect 3167 2485 3171 2486
rect 3263 2490 3267 2491
rect 3263 2485 3267 2486
rect 3391 2490 3395 2491
rect 3391 2485 3395 2486
rect 2384 2461 2386 2485
rect 2560 2461 2562 2485
rect 2752 2461 2754 2485
rect 2952 2461 2954 2485
rect 3168 2461 3170 2485
rect 3392 2461 3394 2485
rect 2382 2460 2388 2461
rect 2382 2456 2383 2460
rect 2387 2456 2388 2460
rect 2382 2455 2388 2456
rect 2558 2460 2564 2461
rect 2558 2456 2559 2460
rect 2563 2456 2564 2460
rect 2558 2455 2564 2456
rect 2750 2460 2756 2461
rect 2750 2456 2751 2460
rect 2755 2456 2756 2460
rect 2750 2455 2756 2456
rect 2950 2460 2956 2461
rect 2950 2456 2951 2460
rect 2955 2456 2956 2460
rect 2950 2455 2956 2456
rect 3166 2460 3172 2461
rect 3166 2456 3167 2460
rect 3171 2456 3172 2460
rect 3166 2455 3172 2456
rect 3390 2460 3396 2461
rect 3390 2456 3391 2460
rect 3395 2456 3396 2460
rect 3390 2455 3396 2456
rect 2146 2451 2152 2452
rect 2146 2447 2147 2451
rect 2151 2447 2152 2451
rect 2146 2446 2152 2447
rect 2290 2451 2296 2452
rect 2290 2447 2291 2451
rect 2295 2447 2296 2451
rect 2290 2446 2296 2447
rect 2298 2451 2304 2452
rect 2298 2447 2299 2451
rect 2303 2447 2304 2451
rect 2298 2446 2304 2447
rect 2470 2451 2476 2452
rect 2470 2447 2471 2451
rect 2475 2447 2476 2451
rect 2470 2446 2476 2447
rect 2642 2451 2648 2452
rect 2642 2447 2643 2451
rect 2647 2447 2648 2451
rect 2642 2446 2648 2447
rect 2898 2451 2904 2452
rect 2898 2447 2899 2451
rect 2903 2447 2904 2451
rect 2898 2446 2904 2447
rect 3034 2451 3040 2452
rect 3034 2447 3035 2451
rect 3039 2447 3040 2451
rect 3034 2446 3040 2447
rect 2070 2441 2076 2442
rect 2046 2440 2052 2441
rect 2046 2436 2047 2440
rect 2051 2436 2052 2440
rect 2070 2437 2071 2441
rect 2075 2437 2076 2441
rect 2070 2436 2076 2437
rect 2046 2435 2052 2436
rect 1902 2431 1908 2432
rect 2006 2433 2012 2434
rect 2006 2429 2007 2433
rect 2011 2429 2012 2433
rect 2006 2428 2012 2429
rect 1738 2427 1744 2428
rect 1738 2423 1739 2427
rect 1743 2423 1744 2427
rect 1738 2422 1744 2423
rect 1866 2427 1872 2428
rect 1866 2423 1867 2427
rect 1871 2423 1872 2427
rect 1866 2422 1872 2423
rect 1662 2417 1668 2418
rect 1662 2413 1663 2417
rect 1667 2413 1668 2417
rect 1662 2412 1668 2413
rect 1578 2407 1584 2408
rect 1578 2403 1579 2407
rect 1583 2403 1584 2407
rect 1578 2402 1584 2403
rect 1664 2391 1666 2412
rect 1740 2400 1742 2422
rect 1790 2417 1796 2418
rect 1790 2413 1791 2417
rect 1795 2413 1796 2417
rect 1790 2412 1796 2413
rect 1738 2399 1744 2400
rect 1738 2395 1739 2399
rect 1743 2395 1744 2399
rect 1738 2394 1744 2395
rect 1792 2391 1794 2412
rect 1868 2400 1870 2422
rect 1902 2417 1908 2418
rect 1902 2413 1903 2417
rect 1907 2413 1908 2417
rect 1902 2412 1908 2413
rect 2006 2416 2012 2417
rect 2006 2412 2007 2416
rect 2011 2412 2012 2416
rect 1866 2399 1872 2400
rect 1866 2395 1867 2399
rect 1871 2395 1872 2399
rect 1866 2394 1872 2395
rect 1818 2391 1824 2392
rect 1904 2391 1906 2412
rect 2006 2411 2012 2412
rect 2008 2391 2010 2411
rect 2048 2399 2050 2435
rect 2072 2399 2074 2436
rect 2148 2424 2150 2446
rect 2214 2441 2220 2442
rect 2214 2437 2215 2441
rect 2219 2437 2220 2441
rect 2214 2436 2220 2437
rect 2146 2423 2152 2424
rect 2146 2419 2147 2423
rect 2151 2419 2152 2423
rect 2146 2418 2152 2419
rect 2216 2399 2218 2436
rect 2292 2424 2294 2446
rect 2382 2441 2388 2442
rect 2382 2437 2383 2441
rect 2387 2437 2388 2441
rect 2382 2436 2388 2437
rect 2290 2423 2296 2424
rect 2290 2419 2291 2423
rect 2295 2419 2296 2423
rect 2290 2418 2296 2419
rect 2384 2399 2386 2436
rect 2047 2398 2051 2399
rect 2047 2393 2051 2394
rect 2071 2398 2075 2399
rect 2071 2393 2075 2394
rect 2215 2398 2219 2399
rect 2215 2393 2219 2394
rect 2247 2398 2251 2399
rect 2247 2393 2251 2394
rect 2383 2398 2387 2399
rect 2383 2393 2387 2394
rect 2431 2398 2435 2399
rect 2431 2393 2435 2394
rect 711 2390 715 2391
rect 711 2385 715 2386
rect 767 2390 771 2391
rect 767 2385 771 2386
rect 903 2390 907 2391
rect 903 2385 907 2386
rect 975 2390 979 2391
rect 975 2385 979 2386
rect 1079 2390 1083 2391
rect 1079 2385 1083 2386
rect 1175 2390 1179 2391
rect 1175 2385 1179 2386
rect 1239 2390 1243 2391
rect 1239 2385 1243 2386
rect 1367 2390 1371 2391
rect 1367 2385 1371 2386
rect 1391 2390 1395 2391
rect 1474 2387 1475 2391
rect 1479 2387 1480 2391
rect 1474 2386 1480 2387
rect 1527 2390 1531 2391
rect 1391 2385 1395 2386
rect 1527 2385 1531 2386
rect 1551 2390 1555 2391
rect 1551 2385 1555 2386
rect 1663 2390 1667 2391
rect 1663 2385 1667 2386
rect 1735 2390 1739 2391
rect 1735 2385 1739 2386
rect 1791 2390 1795 2391
rect 1818 2387 1819 2391
rect 1823 2387 1824 2391
rect 1818 2386 1824 2387
rect 1903 2390 1907 2391
rect 1791 2385 1795 2386
rect 618 2383 624 2384
rect 618 2379 619 2383
rect 623 2379 624 2383
rect 618 2378 624 2379
rect 626 2383 632 2384
rect 626 2379 627 2383
rect 631 2379 632 2383
rect 626 2378 632 2379
rect 550 2363 556 2364
rect 550 2359 551 2363
rect 555 2359 556 2363
rect 550 2358 556 2359
rect 628 2356 630 2378
rect 768 2364 770 2385
rect 842 2383 848 2384
rect 842 2379 843 2383
rect 847 2379 848 2383
rect 842 2378 848 2379
rect 766 2363 772 2364
rect 766 2359 767 2363
rect 771 2359 772 2363
rect 766 2358 772 2359
rect 844 2356 846 2378
rect 976 2364 978 2385
rect 1176 2364 1178 2385
rect 1250 2383 1256 2384
rect 1250 2379 1251 2383
rect 1255 2379 1256 2383
rect 1250 2378 1256 2379
rect 974 2363 980 2364
rect 974 2359 975 2363
rect 979 2359 980 2363
rect 974 2358 980 2359
rect 1174 2363 1180 2364
rect 1174 2359 1175 2363
rect 1179 2359 1180 2363
rect 1174 2358 1180 2359
rect 1252 2356 1254 2378
rect 1368 2364 1370 2385
rect 1442 2383 1448 2384
rect 1442 2379 1443 2383
rect 1447 2379 1448 2383
rect 1442 2378 1448 2379
rect 1366 2363 1372 2364
rect 1366 2359 1367 2363
rect 1371 2359 1372 2363
rect 1366 2358 1372 2359
rect 1444 2356 1446 2378
rect 1552 2364 1554 2385
rect 1626 2383 1632 2384
rect 1626 2379 1627 2383
rect 1631 2379 1632 2383
rect 1626 2378 1632 2379
rect 1550 2363 1556 2364
rect 1550 2359 1551 2363
rect 1555 2359 1556 2363
rect 1550 2358 1556 2359
rect 1628 2356 1630 2378
rect 1736 2364 1738 2385
rect 1734 2363 1740 2364
rect 1734 2359 1735 2363
rect 1739 2359 1740 2363
rect 1734 2358 1740 2359
rect 1820 2356 1822 2386
rect 1903 2385 1907 2386
rect 2007 2390 2011 2391
rect 2007 2385 2011 2386
rect 1904 2364 1906 2385
rect 2008 2365 2010 2385
rect 2048 2373 2050 2393
rect 2054 2383 2060 2384
rect 2054 2379 2055 2383
rect 2059 2379 2060 2383
rect 2054 2378 2060 2379
rect 2046 2372 2052 2373
rect 2046 2368 2047 2372
rect 2051 2368 2052 2372
rect 2046 2367 2052 2368
rect 2006 2364 2012 2365
rect 2056 2364 2058 2378
rect 2072 2372 2074 2393
rect 2154 2391 2160 2392
rect 2154 2387 2155 2391
rect 2159 2387 2160 2391
rect 2154 2386 2160 2387
rect 2070 2371 2076 2372
rect 2070 2367 2071 2371
rect 2075 2367 2076 2371
rect 2070 2366 2076 2367
rect 2156 2364 2158 2386
rect 2248 2372 2250 2393
rect 2258 2391 2264 2392
rect 2258 2387 2259 2391
rect 2263 2387 2264 2391
rect 2258 2386 2264 2387
rect 2246 2371 2252 2372
rect 2246 2367 2247 2371
rect 2251 2367 2252 2371
rect 2246 2366 2252 2367
rect 1902 2363 1908 2364
rect 1902 2359 1903 2363
rect 1907 2359 1908 2363
rect 2006 2360 2007 2364
rect 2011 2360 2012 2364
rect 2006 2359 2012 2360
rect 2054 2363 2060 2364
rect 2054 2359 2055 2363
rect 2059 2359 2060 2363
rect 1902 2358 1908 2359
rect 2054 2358 2060 2359
rect 2154 2363 2160 2364
rect 2154 2359 2155 2363
rect 2159 2359 2160 2363
rect 2154 2358 2160 2359
rect 626 2355 632 2356
rect 626 2351 627 2355
rect 631 2351 632 2355
rect 626 2350 632 2351
rect 842 2355 848 2356
rect 842 2351 843 2355
rect 847 2351 848 2355
rect 842 2350 848 2351
rect 966 2355 972 2356
rect 966 2351 967 2355
rect 971 2351 972 2355
rect 966 2350 972 2351
rect 1250 2355 1256 2356
rect 1250 2351 1251 2355
rect 1255 2351 1256 2355
rect 1250 2350 1256 2351
rect 1442 2355 1448 2356
rect 1442 2351 1443 2355
rect 1447 2351 1448 2355
rect 1442 2350 1448 2351
rect 1626 2355 1632 2356
rect 1626 2351 1627 2355
rect 1631 2351 1632 2355
rect 1626 2350 1632 2351
rect 1670 2355 1676 2356
rect 1670 2351 1671 2355
rect 1675 2351 1676 2355
rect 1670 2350 1676 2351
rect 1818 2355 1824 2356
rect 1818 2351 1819 2355
rect 1823 2351 1824 2355
rect 1818 2350 1824 2351
rect 2046 2355 2052 2356
rect 2046 2351 2047 2355
rect 2051 2351 2052 2355
rect 2046 2350 2052 2351
rect 2070 2352 2076 2353
rect 550 2344 556 2345
rect 550 2340 551 2344
rect 555 2340 556 2344
rect 550 2339 556 2340
rect 766 2344 772 2345
rect 766 2340 767 2344
rect 771 2340 772 2344
rect 766 2339 772 2340
rect 552 2307 554 2339
rect 768 2307 770 2339
rect 431 2306 435 2307
rect 431 2301 435 2302
rect 551 2306 555 2307
rect 551 2301 555 2302
rect 591 2306 595 2307
rect 591 2301 595 2302
rect 751 2306 755 2307
rect 751 2301 755 2302
rect 767 2306 771 2307
rect 767 2301 771 2302
rect 919 2306 923 2307
rect 919 2301 923 2302
rect 432 2277 434 2301
rect 592 2277 594 2301
rect 752 2277 754 2301
rect 920 2277 922 2301
rect 430 2276 436 2277
rect 430 2272 431 2276
rect 435 2272 436 2276
rect 430 2271 436 2272
rect 590 2276 596 2277
rect 590 2272 591 2276
rect 595 2272 596 2276
rect 590 2271 596 2272
rect 750 2276 756 2277
rect 750 2272 751 2276
rect 755 2272 756 2276
rect 750 2271 756 2272
rect 918 2276 924 2277
rect 918 2272 919 2276
rect 923 2272 924 2276
rect 918 2271 924 2272
rect 210 2267 216 2268
rect 210 2263 211 2267
rect 215 2263 216 2267
rect 210 2262 216 2263
rect 346 2267 352 2268
rect 346 2263 347 2267
rect 351 2263 352 2267
rect 346 2262 352 2263
rect 378 2267 384 2268
rect 378 2263 379 2267
rect 383 2263 384 2267
rect 378 2262 384 2263
rect 666 2267 672 2268
rect 666 2263 667 2267
rect 671 2263 672 2267
rect 666 2262 672 2263
rect 734 2267 740 2268
rect 734 2263 735 2267
rect 739 2263 740 2267
rect 734 2262 740 2263
rect 134 2257 140 2258
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 134 2253 135 2257
rect 139 2253 140 2257
rect 134 2252 140 2253
rect 110 2251 116 2252
rect 112 2231 114 2251
rect 136 2231 138 2252
rect 212 2240 214 2262
rect 270 2257 276 2258
rect 270 2253 271 2257
rect 275 2253 276 2257
rect 270 2252 276 2253
rect 210 2239 216 2240
rect 210 2235 211 2239
rect 215 2235 216 2239
rect 210 2234 216 2235
rect 272 2231 274 2252
rect 380 2248 382 2262
rect 430 2257 436 2258
rect 430 2253 431 2257
rect 435 2253 436 2257
rect 430 2252 436 2253
rect 590 2257 596 2258
rect 590 2253 591 2257
rect 595 2253 596 2257
rect 590 2252 596 2253
rect 378 2247 384 2248
rect 378 2243 379 2247
rect 383 2243 384 2247
rect 378 2242 384 2243
rect 402 2235 408 2236
rect 402 2231 403 2235
rect 407 2231 408 2235
rect 432 2231 434 2252
rect 592 2231 594 2252
rect 111 2230 115 2231
rect 111 2225 115 2226
rect 135 2230 139 2231
rect 135 2225 139 2226
rect 159 2230 163 2231
rect 159 2225 163 2226
rect 271 2230 275 2231
rect 271 2225 275 2226
rect 327 2230 331 2231
rect 402 2230 408 2231
rect 431 2230 435 2231
rect 327 2225 331 2226
rect 112 2205 114 2225
rect 110 2204 116 2205
rect 160 2204 162 2225
rect 234 2223 240 2224
rect 234 2219 235 2223
rect 239 2219 240 2223
rect 234 2218 240 2219
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 110 2199 116 2200
rect 158 2203 164 2204
rect 158 2199 159 2203
rect 163 2199 164 2203
rect 158 2198 164 2199
rect 236 2196 238 2218
rect 328 2204 330 2225
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 404 2196 406 2230
rect 431 2225 435 2226
rect 495 2230 499 2231
rect 495 2225 499 2226
rect 591 2230 595 2231
rect 591 2225 595 2226
rect 410 2215 416 2216
rect 410 2211 411 2215
rect 415 2211 416 2215
rect 410 2210 416 2211
rect 412 2196 414 2210
rect 496 2204 498 2225
rect 668 2224 670 2262
rect 736 2240 738 2262
rect 750 2257 756 2258
rect 750 2253 751 2257
rect 755 2253 756 2257
rect 750 2252 756 2253
rect 918 2257 924 2258
rect 918 2253 919 2257
rect 923 2253 924 2257
rect 918 2252 924 2253
rect 734 2239 740 2240
rect 734 2235 735 2239
rect 739 2235 740 2239
rect 734 2234 740 2235
rect 752 2231 754 2252
rect 920 2231 922 2252
rect 968 2244 970 2350
rect 974 2344 980 2345
rect 974 2340 975 2344
rect 979 2340 980 2344
rect 974 2339 980 2340
rect 1174 2344 1180 2345
rect 1174 2340 1175 2344
rect 1179 2340 1180 2344
rect 1174 2339 1180 2340
rect 1366 2344 1372 2345
rect 1366 2340 1367 2344
rect 1371 2340 1372 2344
rect 1366 2339 1372 2340
rect 1550 2344 1556 2345
rect 1550 2340 1551 2344
rect 1555 2340 1556 2344
rect 1550 2339 1556 2340
rect 976 2307 978 2339
rect 1176 2307 1178 2339
rect 1368 2307 1370 2339
rect 1552 2307 1554 2339
rect 975 2306 979 2307
rect 975 2301 979 2302
rect 1087 2306 1091 2307
rect 1087 2301 1091 2302
rect 1175 2306 1179 2307
rect 1175 2301 1179 2302
rect 1263 2306 1267 2307
rect 1263 2301 1267 2302
rect 1367 2306 1371 2307
rect 1367 2301 1371 2302
rect 1447 2306 1451 2307
rect 1447 2301 1451 2302
rect 1551 2306 1555 2307
rect 1551 2301 1555 2302
rect 1631 2306 1635 2307
rect 1631 2301 1635 2302
rect 1088 2277 1090 2301
rect 1264 2277 1266 2301
rect 1448 2277 1450 2301
rect 1632 2277 1634 2301
rect 1086 2276 1092 2277
rect 1086 2272 1087 2276
rect 1091 2272 1092 2276
rect 1086 2271 1092 2272
rect 1262 2276 1268 2277
rect 1262 2272 1263 2276
rect 1267 2272 1268 2276
rect 1262 2271 1268 2272
rect 1446 2276 1452 2277
rect 1446 2272 1447 2276
rect 1451 2272 1452 2276
rect 1446 2271 1452 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 994 2267 1000 2268
rect 994 2263 995 2267
rect 999 2263 1000 2267
rect 994 2262 1000 2263
rect 1162 2267 1168 2268
rect 1162 2263 1163 2267
rect 1167 2263 1168 2267
rect 1162 2262 1168 2263
rect 1338 2267 1344 2268
rect 1338 2263 1339 2267
rect 1343 2263 1344 2267
rect 1338 2262 1344 2263
rect 1522 2267 1528 2268
rect 1522 2263 1523 2267
rect 1527 2263 1528 2267
rect 1522 2262 1528 2263
rect 966 2243 972 2244
rect 966 2239 967 2243
rect 971 2239 972 2243
rect 996 2240 998 2262
rect 1086 2257 1092 2258
rect 1086 2253 1087 2257
rect 1091 2253 1092 2257
rect 1086 2252 1092 2253
rect 966 2238 972 2239
rect 994 2239 1000 2240
rect 986 2235 992 2236
rect 986 2231 987 2235
rect 991 2231 992 2235
rect 994 2235 995 2239
rect 999 2235 1000 2239
rect 994 2234 1000 2235
rect 1088 2231 1090 2252
rect 1164 2240 1166 2262
rect 1262 2257 1268 2258
rect 1262 2253 1263 2257
rect 1267 2253 1268 2257
rect 1262 2252 1268 2253
rect 1162 2239 1168 2240
rect 1162 2235 1163 2239
rect 1167 2235 1168 2239
rect 1162 2234 1168 2235
rect 1264 2231 1266 2252
rect 1340 2240 1342 2262
rect 1446 2257 1452 2258
rect 1446 2253 1447 2257
rect 1451 2253 1452 2257
rect 1446 2252 1452 2253
rect 1338 2239 1344 2240
rect 1338 2235 1339 2239
rect 1343 2235 1344 2239
rect 1338 2234 1344 2235
rect 1448 2231 1450 2252
rect 679 2230 683 2231
rect 679 2225 683 2226
rect 751 2230 755 2231
rect 751 2225 755 2226
rect 879 2230 883 2231
rect 879 2225 883 2226
rect 919 2230 923 2231
rect 986 2230 992 2231
rect 1087 2230 1091 2231
rect 919 2225 923 2226
rect 562 2223 568 2224
rect 562 2219 563 2223
rect 567 2219 568 2223
rect 562 2218 568 2219
rect 666 2223 672 2224
rect 666 2219 667 2223
rect 671 2219 672 2223
rect 666 2218 672 2219
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 234 2195 240 2196
rect 234 2191 235 2195
rect 239 2191 240 2195
rect 234 2190 240 2191
rect 402 2195 408 2196
rect 402 2191 403 2195
rect 407 2191 408 2195
rect 402 2190 408 2191
rect 410 2195 416 2196
rect 410 2191 411 2195
rect 415 2191 416 2195
rect 410 2190 416 2191
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 110 2182 116 2183
rect 158 2184 164 2185
rect 112 2155 114 2182
rect 158 2180 159 2184
rect 163 2180 164 2184
rect 158 2179 164 2180
rect 326 2184 332 2185
rect 326 2180 327 2184
rect 331 2180 332 2184
rect 326 2179 332 2180
rect 494 2184 500 2185
rect 494 2180 495 2184
rect 499 2180 500 2184
rect 494 2179 500 2180
rect 160 2155 162 2179
rect 328 2155 330 2179
rect 496 2155 498 2179
rect 111 2154 115 2155
rect 111 2149 115 2150
rect 159 2154 163 2155
rect 159 2149 163 2150
rect 223 2154 227 2155
rect 223 2149 227 2150
rect 327 2154 331 2155
rect 327 2149 331 2150
rect 359 2154 363 2155
rect 359 2149 363 2150
rect 495 2154 499 2155
rect 495 2149 499 2150
rect 112 2122 114 2149
rect 224 2125 226 2149
rect 360 2125 362 2149
rect 496 2125 498 2149
rect 222 2124 228 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 222 2120 223 2124
rect 227 2120 228 2124
rect 222 2119 228 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 494 2124 500 2125
rect 494 2120 495 2124
rect 499 2120 500 2124
rect 494 2119 500 2120
rect 110 2116 116 2117
rect 564 2116 566 2218
rect 680 2204 682 2225
rect 880 2204 882 2225
rect 678 2203 684 2204
rect 678 2199 679 2203
rect 683 2199 684 2203
rect 678 2198 684 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 988 2196 990 2230
rect 1087 2225 1091 2226
rect 1095 2230 1099 2231
rect 1095 2225 1099 2226
rect 1263 2230 1267 2231
rect 1263 2225 1267 2226
rect 1327 2230 1331 2231
rect 1327 2225 1331 2226
rect 1447 2230 1451 2231
rect 1447 2225 1451 2226
rect 1096 2204 1098 2225
rect 1162 2223 1168 2224
rect 1162 2219 1163 2223
rect 1167 2219 1168 2223
rect 1162 2218 1168 2219
rect 1094 2203 1100 2204
rect 1094 2199 1095 2203
rect 1099 2199 1100 2203
rect 1094 2198 1100 2199
rect 826 2195 832 2196
rect 826 2191 827 2195
rect 831 2191 832 2195
rect 826 2190 832 2191
rect 986 2195 992 2196
rect 986 2191 987 2195
rect 991 2191 992 2195
rect 986 2190 992 2191
rect 678 2184 684 2185
rect 678 2180 679 2184
rect 683 2180 684 2184
rect 678 2179 684 2180
rect 680 2155 682 2179
rect 639 2154 643 2155
rect 639 2149 643 2150
rect 679 2154 683 2155
rect 679 2149 683 2150
rect 783 2154 787 2155
rect 783 2149 787 2150
rect 640 2125 642 2149
rect 784 2125 786 2149
rect 638 2124 644 2125
rect 638 2120 639 2124
rect 643 2120 644 2124
rect 638 2119 644 2120
rect 782 2124 788 2125
rect 782 2120 783 2124
rect 787 2120 788 2124
rect 782 2119 788 2120
rect 298 2115 304 2116
rect 298 2111 299 2115
rect 303 2111 304 2115
rect 298 2110 304 2111
rect 434 2115 440 2116
rect 434 2111 435 2115
rect 439 2111 440 2115
rect 434 2110 440 2111
rect 562 2115 568 2116
rect 562 2111 563 2115
rect 567 2111 568 2115
rect 562 2110 568 2111
rect 578 2115 584 2116
rect 578 2111 579 2115
rect 583 2111 584 2115
rect 578 2110 584 2111
rect 222 2105 228 2106
rect 110 2104 116 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 222 2101 223 2105
rect 227 2101 228 2105
rect 222 2100 228 2101
rect 110 2099 116 2100
rect 112 2071 114 2099
rect 224 2071 226 2100
rect 300 2084 302 2110
rect 358 2105 364 2106
rect 358 2101 359 2105
rect 363 2101 364 2105
rect 358 2100 364 2101
rect 298 2083 304 2084
rect 298 2079 299 2083
rect 303 2079 304 2083
rect 298 2078 304 2079
rect 360 2071 362 2100
rect 436 2088 438 2110
rect 494 2105 500 2106
rect 494 2101 495 2105
rect 499 2101 500 2105
rect 494 2100 500 2101
rect 434 2087 440 2088
rect 434 2083 435 2087
rect 439 2083 440 2087
rect 434 2082 440 2083
rect 496 2071 498 2100
rect 580 2096 582 2110
rect 638 2105 644 2106
rect 638 2101 639 2105
rect 643 2101 644 2105
rect 638 2100 644 2101
rect 782 2105 788 2106
rect 782 2101 783 2105
rect 787 2101 788 2105
rect 782 2100 788 2101
rect 578 2095 584 2096
rect 578 2091 579 2095
rect 583 2091 584 2095
rect 578 2090 584 2091
rect 640 2071 642 2100
rect 690 2083 696 2084
rect 690 2079 691 2083
rect 695 2079 696 2083
rect 690 2078 696 2079
rect 111 2070 115 2071
rect 111 2065 115 2066
rect 223 2070 227 2071
rect 223 2065 227 2066
rect 359 2070 363 2071
rect 359 2065 363 2066
rect 375 2070 379 2071
rect 375 2065 379 2066
rect 495 2070 499 2071
rect 495 2065 499 2066
rect 615 2070 619 2071
rect 615 2065 619 2066
rect 639 2070 643 2071
rect 639 2065 643 2066
rect 112 2045 114 2065
rect 110 2044 116 2045
rect 376 2044 378 2065
rect 414 2063 420 2064
rect 414 2059 415 2063
rect 419 2059 420 2063
rect 414 2058 420 2059
rect 450 2063 456 2064
rect 450 2059 451 2063
rect 455 2059 456 2063
rect 450 2058 456 2059
rect 110 2040 111 2044
rect 115 2040 116 2044
rect 110 2039 116 2040
rect 374 2043 380 2044
rect 374 2039 375 2043
rect 379 2039 380 2043
rect 374 2038 380 2039
rect 110 2027 116 2028
rect 110 2023 111 2027
rect 115 2023 116 2027
rect 110 2022 116 2023
rect 374 2024 380 2025
rect 112 1987 114 2022
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 376 1987 378 2019
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 375 1986 379 1987
rect 375 1981 379 1982
rect 112 1954 114 1981
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 110 1948 116 1949
rect 416 1948 418 2058
rect 452 2036 454 2058
rect 496 2044 498 2065
rect 570 2063 576 2064
rect 570 2059 571 2063
rect 575 2059 576 2063
rect 570 2058 576 2059
rect 494 2043 500 2044
rect 494 2039 495 2043
rect 499 2039 500 2043
rect 494 2038 500 2039
rect 572 2036 574 2058
rect 616 2044 618 2065
rect 614 2043 620 2044
rect 614 2039 615 2043
rect 619 2039 620 2043
rect 614 2038 620 2039
rect 692 2036 694 2078
rect 784 2071 786 2100
rect 828 2088 830 2190
rect 878 2184 884 2185
rect 878 2180 879 2184
rect 883 2180 884 2184
rect 878 2179 884 2180
rect 1094 2184 1100 2185
rect 1094 2180 1095 2184
rect 1099 2180 1100 2184
rect 1094 2179 1100 2180
rect 880 2155 882 2179
rect 1096 2155 1098 2179
rect 879 2154 883 2155
rect 879 2149 883 2150
rect 935 2154 939 2155
rect 935 2149 939 2150
rect 1095 2154 1099 2155
rect 1095 2149 1099 2150
rect 936 2125 938 2149
rect 1096 2125 1098 2149
rect 934 2124 940 2125
rect 934 2120 935 2124
rect 939 2120 940 2124
rect 934 2119 940 2120
rect 1094 2124 1100 2125
rect 1094 2120 1095 2124
rect 1099 2120 1100 2124
rect 1094 2119 1100 2120
rect 1164 2116 1166 2218
rect 1328 2204 1330 2225
rect 1524 2224 1526 2262
rect 1630 2257 1636 2258
rect 1630 2253 1631 2257
rect 1635 2253 1636 2257
rect 1630 2252 1636 2253
rect 1632 2231 1634 2252
rect 1672 2240 1674 2350
rect 2006 2347 2012 2348
rect 1734 2344 1740 2345
rect 1734 2340 1735 2344
rect 1739 2340 1740 2344
rect 1734 2339 1740 2340
rect 1902 2344 1908 2345
rect 1902 2340 1903 2344
rect 1907 2340 1908 2344
rect 2006 2343 2007 2347
rect 2011 2343 2012 2347
rect 2006 2342 2012 2343
rect 1902 2339 1908 2340
rect 1736 2307 1738 2339
rect 1904 2307 1906 2339
rect 2008 2307 2010 2342
rect 2048 2323 2050 2350
rect 2070 2348 2071 2352
rect 2075 2348 2076 2352
rect 2070 2347 2076 2348
rect 2246 2352 2252 2353
rect 2246 2348 2247 2352
rect 2251 2348 2252 2352
rect 2246 2347 2252 2348
rect 2072 2323 2074 2347
rect 2248 2323 2250 2347
rect 2047 2322 2051 2323
rect 2047 2317 2051 2318
rect 2071 2322 2075 2323
rect 2071 2317 2075 2318
rect 2175 2322 2179 2323
rect 2175 2317 2179 2318
rect 2247 2322 2251 2323
rect 2247 2317 2251 2318
rect 1735 2306 1739 2307
rect 1735 2301 1739 2302
rect 1815 2306 1819 2307
rect 1815 2301 1819 2302
rect 1903 2306 1907 2307
rect 1903 2301 1907 2302
rect 2007 2306 2011 2307
rect 2007 2301 2011 2302
rect 1816 2277 1818 2301
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 2008 2274 2010 2301
rect 2048 2290 2050 2317
rect 2072 2293 2074 2317
rect 2176 2293 2178 2317
rect 2070 2292 2076 2293
rect 2046 2289 2052 2290
rect 2046 2285 2047 2289
rect 2051 2285 2052 2289
rect 2070 2288 2071 2292
rect 2075 2288 2076 2292
rect 2070 2287 2076 2288
rect 2174 2292 2180 2293
rect 2174 2288 2175 2292
rect 2179 2288 2180 2292
rect 2174 2287 2180 2288
rect 2046 2284 2052 2285
rect 2260 2284 2262 2386
rect 2432 2372 2434 2393
rect 2472 2392 2474 2446
rect 2558 2441 2564 2442
rect 2558 2437 2559 2441
rect 2563 2437 2564 2441
rect 2558 2436 2564 2437
rect 2560 2399 2562 2436
rect 2644 2424 2646 2446
rect 2750 2441 2756 2442
rect 2750 2437 2751 2441
rect 2755 2437 2756 2441
rect 2750 2436 2756 2437
rect 2642 2423 2648 2424
rect 2642 2419 2643 2423
rect 2647 2419 2648 2423
rect 2642 2418 2648 2419
rect 2752 2399 2754 2436
rect 2900 2424 2902 2446
rect 2950 2441 2956 2442
rect 2950 2437 2951 2441
rect 2955 2437 2956 2441
rect 2950 2436 2956 2437
rect 2898 2423 2904 2424
rect 2898 2419 2899 2423
rect 2903 2419 2904 2423
rect 2898 2418 2904 2419
rect 2952 2399 2954 2436
rect 3036 2424 3038 2446
rect 3166 2441 3172 2442
rect 3166 2437 3167 2441
rect 3171 2437 3172 2441
rect 3166 2436 3172 2437
rect 3390 2441 3396 2442
rect 3390 2437 3391 2441
rect 3395 2437 3396 2441
rect 3390 2436 3396 2437
rect 3034 2423 3040 2424
rect 3034 2419 3035 2423
rect 3039 2419 3040 2423
rect 3034 2418 3040 2419
rect 3168 2399 3170 2436
rect 3392 2399 3394 2436
rect 3452 2424 3454 2530
rect 3502 2524 3508 2525
rect 3502 2520 3503 2524
rect 3507 2520 3508 2524
rect 3502 2519 3508 2520
rect 3504 2491 3506 2519
rect 3503 2490 3507 2491
rect 3503 2485 3507 2486
rect 3623 2490 3627 2491
rect 3623 2485 3627 2486
rect 3624 2461 3626 2485
rect 3622 2460 3628 2461
rect 3622 2456 3623 2460
rect 3627 2456 3628 2460
rect 3622 2455 3628 2456
rect 3700 2452 3702 2558
rect 3728 2536 3730 2578
rect 3840 2571 3842 2600
rect 3908 2588 3910 2686
rect 3944 2655 3946 2686
rect 3943 2654 3947 2655
rect 3943 2649 3947 2650
rect 3944 2622 3946 2649
rect 3942 2621 3948 2622
rect 3942 2617 3943 2621
rect 3947 2617 3948 2621
rect 3942 2616 3948 2617
rect 3922 2615 3928 2616
rect 3922 2611 3923 2615
rect 3927 2611 3928 2615
rect 3922 2610 3928 2611
rect 3906 2587 3912 2588
rect 3906 2583 3907 2587
rect 3911 2583 3912 2587
rect 3906 2582 3912 2583
rect 3743 2570 3747 2571
rect 3743 2565 3747 2566
rect 3839 2570 3843 2571
rect 3839 2565 3843 2566
rect 3744 2544 3746 2565
rect 3742 2543 3748 2544
rect 3742 2539 3743 2543
rect 3747 2539 3748 2543
rect 3742 2538 3748 2539
rect 3726 2535 3732 2536
rect 3726 2531 3727 2535
rect 3731 2531 3732 2535
rect 3726 2530 3732 2531
rect 3742 2524 3748 2525
rect 3742 2520 3743 2524
rect 3747 2520 3748 2524
rect 3742 2519 3748 2520
rect 3744 2491 3746 2519
rect 3743 2490 3747 2491
rect 3743 2485 3747 2486
rect 3839 2490 3843 2491
rect 3839 2485 3843 2486
rect 3840 2461 3842 2485
rect 3838 2460 3844 2461
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3838 2455 3844 2456
rect 3698 2451 3704 2452
rect 3698 2447 3699 2451
rect 3703 2447 3704 2451
rect 3698 2446 3704 2447
rect 3906 2451 3912 2452
rect 3906 2447 3907 2451
rect 3911 2447 3912 2451
rect 3906 2446 3912 2447
rect 3622 2441 3628 2442
rect 3622 2437 3623 2441
rect 3627 2437 3628 2441
rect 3622 2436 3628 2437
rect 3838 2441 3844 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3450 2423 3456 2424
rect 3450 2419 3451 2423
rect 3455 2419 3456 2423
rect 3450 2418 3456 2419
rect 3624 2399 3626 2436
rect 3746 2419 3752 2420
rect 3746 2415 3747 2419
rect 3751 2415 3752 2419
rect 3746 2414 3752 2415
rect 2559 2398 2563 2399
rect 2559 2393 2563 2394
rect 2607 2398 2611 2399
rect 2607 2393 2611 2394
rect 2751 2398 2755 2399
rect 2751 2393 2755 2394
rect 2775 2398 2779 2399
rect 2775 2393 2779 2394
rect 2935 2398 2939 2399
rect 2935 2393 2939 2394
rect 2951 2398 2955 2399
rect 2951 2393 2955 2394
rect 3103 2398 3107 2399
rect 3103 2393 3107 2394
rect 3167 2398 3171 2399
rect 3167 2393 3171 2394
rect 3391 2398 3395 2399
rect 3391 2393 3395 2394
rect 3623 2398 3627 2399
rect 3623 2393 3627 2394
rect 2470 2391 2476 2392
rect 2470 2387 2471 2391
rect 2475 2387 2476 2391
rect 2470 2386 2476 2387
rect 2506 2391 2512 2392
rect 2506 2387 2507 2391
rect 2511 2387 2512 2391
rect 2506 2386 2512 2387
rect 2430 2371 2436 2372
rect 2430 2367 2431 2371
rect 2435 2367 2436 2371
rect 2430 2366 2436 2367
rect 2508 2364 2510 2386
rect 2608 2372 2610 2393
rect 2682 2391 2688 2392
rect 2682 2387 2683 2391
rect 2687 2387 2688 2391
rect 2682 2386 2688 2387
rect 2606 2371 2612 2372
rect 2606 2367 2607 2371
rect 2611 2367 2612 2371
rect 2606 2366 2612 2367
rect 2684 2364 2686 2386
rect 2776 2372 2778 2393
rect 2850 2391 2856 2392
rect 2850 2387 2851 2391
rect 2855 2387 2856 2391
rect 2850 2386 2856 2387
rect 2774 2371 2780 2372
rect 2774 2367 2775 2371
rect 2779 2367 2780 2371
rect 2774 2366 2780 2367
rect 2852 2364 2854 2386
rect 2936 2372 2938 2393
rect 3010 2391 3016 2392
rect 3010 2387 3011 2391
rect 3015 2387 3016 2391
rect 3010 2386 3016 2387
rect 2934 2371 2940 2372
rect 2934 2367 2935 2371
rect 2939 2367 2940 2371
rect 2934 2366 2940 2367
rect 3012 2364 3014 2386
rect 3104 2372 3106 2393
rect 3102 2371 3108 2372
rect 3102 2367 3103 2371
rect 3107 2367 3108 2371
rect 3102 2366 3108 2367
rect 2506 2363 2512 2364
rect 2506 2359 2507 2363
rect 2511 2359 2512 2363
rect 2506 2358 2512 2359
rect 2682 2363 2688 2364
rect 2682 2359 2683 2363
rect 2687 2359 2688 2363
rect 2682 2358 2688 2359
rect 2850 2363 2856 2364
rect 2850 2359 2851 2363
rect 2855 2359 2856 2363
rect 2850 2358 2856 2359
rect 3010 2363 3016 2364
rect 3010 2359 3011 2363
rect 3015 2359 3016 2363
rect 3010 2358 3016 2359
rect 3018 2363 3024 2364
rect 3018 2359 3019 2363
rect 3023 2359 3024 2363
rect 3018 2358 3024 2359
rect 2430 2352 2436 2353
rect 2430 2348 2431 2352
rect 2435 2348 2436 2352
rect 2430 2347 2436 2348
rect 2606 2352 2612 2353
rect 2606 2348 2607 2352
rect 2611 2348 2612 2352
rect 2606 2347 2612 2348
rect 2774 2352 2780 2353
rect 2774 2348 2775 2352
rect 2779 2348 2780 2352
rect 2774 2347 2780 2348
rect 2934 2352 2940 2353
rect 2934 2348 2935 2352
rect 2939 2348 2940 2352
rect 2934 2347 2940 2348
rect 2432 2323 2434 2347
rect 2608 2323 2610 2347
rect 2776 2323 2778 2347
rect 2936 2323 2938 2347
rect 2311 2322 2315 2323
rect 2311 2317 2315 2318
rect 2431 2322 2435 2323
rect 2431 2317 2435 2318
rect 2447 2322 2451 2323
rect 2447 2317 2451 2318
rect 2591 2322 2595 2323
rect 2591 2317 2595 2318
rect 2607 2322 2611 2323
rect 2607 2317 2611 2318
rect 2751 2322 2755 2323
rect 2751 2317 2755 2318
rect 2775 2322 2779 2323
rect 2775 2317 2779 2318
rect 2935 2322 2939 2323
rect 2935 2317 2939 2318
rect 2312 2293 2314 2317
rect 2448 2293 2450 2317
rect 2592 2293 2594 2317
rect 2752 2293 2754 2317
rect 2936 2293 2938 2317
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2446 2292 2452 2293
rect 2446 2288 2447 2292
rect 2451 2288 2452 2292
rect 2446 2287 2452 2288
rect 2590 2292 2596 2293
rect 2590 2288 2591 2292
rect 2595 2288 2596 2292
rect 2590 2287 2596 2288
rect 2750 2292 2756 2293
rect 2750 2288 2751 2292
rect 2755 2288 2756 2292
rect 2750 2287 2756 2288
rect 2934 2292 2940 2293
rect 2934 2288 2935 2292
rect 2939 2288 2940 2292
rect 2934 2287 2940 2288
rect 2146 2283 2152 2284
rect 2146 2279 2147 2283
rect 2151 2279 2152 2283
rect 2146 2278 2152 2279
rect 2258 2283 2264 2284
rect 2258 2279 2259 2283
rect 2263 2279 2264 2283
rect 2258 2278 2264 2279
rect 2266 2283 2272 2284
rect 2266 2279 2267 2283
rect 2271 2279 2272 2283
rect 2266 2278 2272 2279
rect 2522 2283 2528 2284
rect 2522 2279 2523 2283
rect 2527 2279 2528 2283
rect 2522 2278 2528 2279
rect 2530 2283 2536 2284
rect 2530 2279 2531 2283
rect 2535 2279 2536 2283
rect 2530 2278 2536 2279
rect 2826 2283 2832 2284
rect 2826 2279 2827 2283
rect 2831 2279 2832 2283
rect 2826 2278 2832 2279
rect 3010 2283 3016 2284
rect 3010 2279 3011 2283
rect 3015 2279 3016 2283
rect 3010 2278 3016 2279
rect 1814 2271 1820 2272
rect 2006 2273 2012 2274
rect 2070 2273 2076 2274
rect 2006 2269 2007 2273
rect 2011 2269 2012 2273
rect 2006 2268 2012 2269
rect 2046 2272 2052 2273
rect 2046 2268 2047 2272
rect 2051 2268 2052 2272
rect 2070 2269 2071 2273
rect 2075 2269 2076 2273
rect 2070 2268 2076 2269
rect 1706 2267 1712 2268
rect 1706 2263 1707 2267
rect 1711 2263 1712 2267
rect 1706 2262 1712 2263
rect 1882 2267 1888 2268
rect 2046 2267 2052 2268
rect 1882 2263 1883 2267
rect 1887 2263 1888 2267
rect 1882 2262 1888 2263
rect 1708 2240 1710 2262
rect 1814 2257 1820 2258
rect 1814 2253 1815 2257
rect 1819 2253 1820 2257
rect 1814 2252 1820 2253
rect 1670 2239 1676 2240
rect 1670 2235 1671 2239
rect 1675 2235 1676 2239
rect 1670 2234 1676 2235
rect 1706 2239 1712 2240
rect 1706 2235 1707 2239
rect 1711 2235 1712 2239
rect 1706 2234 1712 2235
rect 1816 2231 1818 2252
rect 1567 2230 1571 2231
rect 1567 2225 1571 2226
rect 1631 2230 1635 2231
rect 1631 2225 1635 2226
rect 1815 2230 1819 2231
rect 1815 2225 1819 2226
rect 1410 2223 1416 2224
rect 1410 2219 1411 2223
rect 1415 2219 1416 2223
rect 1410 2218 1416 2219
rect 1522 2223 1528 2224
rect 1522 2219 1523 2223
rect 1527 2219 1528 2223
rect 1522 2218 1528 2219
rect 1326 2203 1332 2204
rect 1326 2199 1327 2203
rect 1331 2199 1332 2203
rect 1326 2198 1332 2199
rect 1412 2196 1414 2218
rect 1568 2204 1570 2225
rect 1816 2204 1818 2225
rect 1884 2224 1886 2262
rect 2006 2256 2012 2257
rect 2006 2252 2007 2256
rect 2011 2252 2012 2256
rect 2006 2251 2012 2252
rect 2008 2231 2010 2251
rect 2048 2239 2050 2267
rect 2072 2239 2074 2268
rect 2148 2256 2150 2278
rect 2174 2273 2180 2274
rect 2174 2269 2175 2273
rect 2179 2269 2180 2273
rect 2174 2268 2180 2269
rect 2146 2255 2152 2256
rect 2146 2251 2147 2255
rect 2151 2251 2152 2255
rect 2146 2250 2152 2251
rect 2176 2239 2178 2268
rect 2268 2264 2270 2278
rect 2310 2273 2316 2274
rect 2310 2269 2311 2273
rect 2315 2269 2316 2273
rect 2310 2268 2316 2269
rect 2446 2273 2452 2274
rect 2446 2269 2447 2273
rect 2451 2269 2452 2273
rect 2446 2268 2452 2269
rect 2266 2263 2272 2264
rect 2266 2259 2267 2263
rect 2271 2259 2272 2263
rect 2266 2258 2272 2259
rect 2312 2239 2314 2268
rect 2448 2239 2450 2268
rect 2524 2256 2526 2278
rect 2532 2264 2534 2278
rect 2590 2273 2596 2274
rect 2590 2269 2591 2273
rect 2595 2269 2596 2273
rect 2590 2268 2596 2269
rect 2750 2273 2756 2274
rect 2750 2269 2751 2273
rect 2755 2269 2756 2273
rect 2750 2268 2756 2269
rect 2530 2263 2536 2264
rect 2530 2259 2531 2263
rect 2535 2259 2536 2263
rect 2530 2258 2536 2259
rect 2522 2255 2528 2256
rect 2482 2251 2488 2252
rect 2482 2247 2483 2251
rect 2487 2247 2488 2251
rect 2522 2251 2523 2255
rect 2527 2251 2528 2255
rect 2522 2250 2528 2251
rect 2482 2246 2488 2247
rect 2047 2238 2051 2239
rect 2047 2233 2051 2234
rect 2071 2238 2075 2239
rect 2071 2233 2075 2234
rect 2111 2238 2115 2239
rect 2111 2233 2115 2234
rect 2175 2238 2179 2239
rect 2175 2233 2179 2234
rect 2255 2238 2259 2239
rect 2255 2233 2259 2234
rect 2311 2238 2315 2239
rect 2311 2233 2315 2234
rect 2407 2238 2411 2239
rect 2407 2233 2411 2234
rect 2447 2238 2451 2239
rect 2447 2233 2451 2234
rect 2007 2230 2011 2231
rect 2007 2225 2011 2226
rect 1882 2223 1888 2224
rect 1882 2219 1883 2223
rect 1887 2219 1888 2223
rect 1882 2218 1888 2219
rect 2008 2205 2010 2225
rect 2048 2213 2050 2233
rect 2046 2212 2052 2213
rect 2112 2212 2114 2233
rect 2186 2231 2192 2232
rect 2186 2227 2187 2231
rect 2191 2227 2192 2231
rect 2186 2226 2192 2227
rect 2046 2208 2047 2212
rect 2051 2208 2052 2212
rect 2046 2207 2052 2208
rect 2110 2211 2116 2212
rect 2110 2207 2111 2211
rect 2115 2207 2116 2211
rect 2110 2206 2116 2207
rect 2006 2204 2012 2205
rect 2188 2204 2190 2226
rect 2256 2212 2258 2233
rect 2330 2231 2336 2232
rect 2330 2227 2331 2231
rect 2335 2227 2336 2231
rect 2330 2226 2336 2227
rect 2254 2211 2260 2212
rect 2254 2207 2255 2211
rect 2259 2207 2260 2211
rect 2254 2206 2260 2207
rect 2332 2204 2334 2226
rect 2408 2212 2410 2233
rect 2406 2211 2412 2212
rect 2406 2207 2407 2211
rect 2411 2207 2412 2211
rect 2406 2206 2412 2207
rect 2484 2204 2486 2246
rect 2592 2239 2594 2268
rect 2752 2239 2754 2268
rect 2828 2252 2830 2278
rect 2934 2273 2940 2274
rect 2934 2269 2935 2273
rect 2939 2269 2940 2273
rect 2934 2268 2940 2269
rect 2826 2251 2832 2252
rect 2826 2247 2827 2251
rect 2831 2247 2832 2251
rect 2826 2246 2832 2247
rect 2936 2239 2938 2268
rect 3012 2256 3014 2278
rect 3020 2264 3022 2358
rect 3102 2352 3108 2353
rect 3102 2348 3103 2352
rect 3107 2348 3108 2352
rect 3102 2347 3108 2348
rect 3104 2323 3106 2347
rect 3103 2322 3107 2323
rect 3103 2317 3107 2318
rect 3143 2322 3147 2323
rect 3143 2317 3147 2318
rect 3375 2322 3379 2323
rect 3375 2317 3379 2318
rect 3615 2322 3619 2323
rect 3615 2317 3619 2318
rect 3144 2293 3146 2317
rect 3376 2293 3378 2317
rect 3616 2293 3618 2317
rect 3142 2292 3148 2293
rect 3142 2288 3143 2292
rect 3147 2288 3148 2292
rect 3142 2287 3148 2288
rect 3374 2292 3380 2293
rect 3374 2288 3375 2292
rect 3379 2288 3380 2292
rect 3374 2287 3380 2288
rect 3614 2292 3620 2293
rect 3614 2288 3615 2292
rect 3619 2288 3620 2292
rect 3614 2287 3620 2288
rect 3218 2283 3224 2284
rect 3218 2279 3219 2283
rect 3223 2279 3224 2283
rect 3218 2278 3224 2279
rect 3450 2283 3456 2284
rect 3450 2279 3451 2283
rect 3455 2279 3456 2283
rect 3450 2278 3456 2279
rect 3506 2283 3512 2284
rect 3506 2279 3507 2283
rect 3511 2279 3512 2283
rect 3506 2278 3512 2279
rect 3142 2273 3148 2274
rect 3142 2269 3143 2273
rect 3147 2269 3148 2273
rect 3142 2268 3148 2269
rect 3018 2263 3024 2264
rect 3018 2259 3019 2263
rect 3023 2259 3024 2263
rect 3018 2258 3024 2259
rect 3010 2255 3016 2256
rect 3010 2251 3011 2255
rect 3015 2251 3016 2255
rect 3010 2250 3016 2251
rect 3144 2239 3146 2268
rect 3220 2256 3222 2278
rect 3374 2273 3380 2274
rect 3374 2269 3375 2273
rect 3379 2269 3380 2273
rect 3374 2268 3380 2269
rect 3218 2255 3224 2256
rect 3218 2251 3219 2255
rect 3223 2251 3224 2255
rect 3218 2250 3224 2251
rect 3376 2239 3378 2268
rect 3452 2256 3454 2278
rect 3450 2255 3456 2256
rect 3450 2251 3451 2255
rect 3455 2251 3456 2255
rect 3450 2250 3456 2251
rect 3508 2240 3510 2278
rect 3614 2273 3620 2274
rect 3614 2269 3615 2273
rect 3619 2269 3620 2273
rect 3614 2268 3620 2269
rect 3506 2239 3512 2240
rect 3616 2239 3618 2268
rect 2559 2238 2563 2239
rect 2559 2233 2563 2234
rect 2591 2238 2595 2239
rect 2591 2233 2595 2234
rect 2719 2238 2723 2239
rect 2719 2233 2723 2234
rect 2751 2238 2755 2239
rect 2751 2233 2755 2234
rect 2879 2238 2883 2239
rect 2879 2233 2883 2234
rect 2935 2238 2939 2239
rect 2935 2233 2939 2234
rect 3047 2238 3051 2239
rect 3047 2233 3051 2234
rect 3143 2238 3147 2239
rect 3143 2233 3147 2234
rect 3223 2238 3227 2239
rect 3223 2233 3227 2234
rect 3375 2238 3379 2239
rect 3375 2233 3379 2234
rect 3407 2238 3411 2239
rect 3506 2235 3507 2239
rect 3511 2235 3512 2239
rect 3506 2234 3512 2235
rect 3591 2238 3595 2239
rect 3407 2233 3411 2234
rect 3591 2233 3595 2234
rect 3615 2238 3619 2239
rect 3615 2233 3619 2234
rect 2490 2223 2496 2224
rect 2490 2219 2491 2223
rect 2495 2219 2496 2223
rect 2490 2218 2496 2219
rect 2492 2204 2494 2218
rect 2560 2212 2562 2233
rect 2642 2231 2648 2232
rect 2642 2227 2643 2231
rect 2647 2227 2648 2231
rect 2642 2226 2648 2227
rect 2658 2231 2664 2232
rect 2658 2227 2659 2231
rect 2663 2227 2664 2231
rect 2658 2226 2664 2227
rect 2558 2211 2564 2212
rect 2558 2207 2559 2211
rect 2563 2207 2564 2211
rect 2558 2206 2564 2207
rect 2644 2204 2646 2226
rect 1566 2203 1572 2204
rect 1566 2199 1567 2203
rect 1571 2199 1572 2203
rect 1566 2198 1572 2199
rect 1814 2203 1820 2204
rect 1814 2199 1815 2203
rect 1819 2199 1820 2203
rect 2006 2200 2007 2204
rect 2011 2200 2012 2204
rect 2006 2199 2012 2200
rect 2186 2203 2192 2204
rect 2186 2199 2187 2203
rect 2191 2199 2192 2203
rect 1814 2198 1820 2199
rect 2186 2198 2192 2199
rect 2330 2203 2336 2204
rect 2330 2199 2331 2203
rect 2335 2199 2336 2203
rect 2330 2198 2336 2199
rect 2482 2203 2488 2204
rect 2482 2199 2483 2203
rect 2487 2199 2488 2203
rect 2482 2198 2488 2199
rect 2490 2203 2496 2204
rect 2490 2199 2491 2203
rect 2495 2199 2496 2203
rect 2490 2198 2496 2199
rect 2642 2203 2648 2204
rect 2642 2199 2643 2203
rect 2647 2199 2648 2203
rect 2642 2198 2648 2199
rect 1302 2195 1308 2196
rect 1302 2191 1303 2195
rect 1307 2191 1308 2195
rect 1302 2190 1308 2191
rect 1410 2195 1416 2196
rect 1410 2191 1411 2195
rect 1415 2191 1416 2195
rect 2046 2195 2052 2196
rect 1410 2190 1416 2191
rect 1890 2191 1896 2192
rect 1263 2154 1267 2155
rect 1263 2149 1267 2150
rect 1264 2125 1266 2149
rect 1262 2124 1268 2125
rect 1262 2120 1263 2124
rect 1267 2120 1268 2124
rect 1262 2119 1268 2120
rect 1010 2115 1016 2116
rect 1010 2111 1011 2115
rect 1015 2111 1016 2115
rect 1010 2110 1016 2111
rect 1162 2115 1168 2116
rect 1162 2111 1163 2115
rect 1167 2111 1168 2115
rect 1162 2110 1168 2111
rect 934 2105 940 2106
rect 934 2101 935 2105
rect 939 2101 940 2105
rect 934 2100 940 2101
rect 822 2087 830 2088
rect 822 2083 823 2087
rect 827 2084 830 2087
rect 827 2083 828 2084
rect 822 2082 828 2083
rect 936 2071 938 2100
rect 1012 2088 1014 2110
rect 1094 2105 1100 2106
rect 1094 2101 1095 2105
rect 1099 2101 1100 2105
rect 1094 2100 1100 2101
rect 1262 2105 1268 2106
rect 1262 2101 1263 2105
rect 1267 2101 1268 2105
rect 1262 2100 1268 2101
rect 1010 2087 1016 2088
rect 1002 2083 1008 2084
rect 1002 2079 1003 2083
rect 1007 2079 1008 2083
rect 1010 2083 1011 2087
rect 1015 2083 1016 2087
rect 1010 2082 1016 2083
rect 1002 2078 1008 2079
rect 751 2070 755 2071
rect 751 2065 755 2066
rect 783 2070 787 2071
rect 783 2065 787 2066
rect 895 2070 899 2071
rect 895 2065 899 2066
rect 935 2070 939 2071
rect 935 2065 939 2066
rect 752 2044 754 2065
rect 826 2063 832 2064
rect 826 2059 827 2063
rect 831 2059 832 2063
rect 826 2058 832 2059
rect 750 2043 756 2044
rect 750 2039 751 2043
rect 755 2039 756 2043
rect 750 2038 756 2039
rect 828 2036 830 2058
rect 896 2044 898 2065
rect 894 2043 900 2044
rect 894 2039 895 2043
rect 899 2039 900 2043
rect 894 2038 900 2039
rect 1004 2036 1006 2078
rect 1096 2071 1098 2100
rect 1264 2071 1266 2100
rect 1304 2088 1306 2190
rect 1890 2187 1891 2191
rect 1895 2187 1896 2191
rect 2046 2191 2047 2195
rect 2051 2191 2052 2195
rect 2046 2190 2052 2191
rect 2110 2192 2116 2193
rect 1890 2186 1896 2187
rect 2006 2187 2012 2188
rect 1326 2184 1332 2185
rect 1326 2180 1327 2184
rect 1331 2180 1332 2184
rect 1326 2179 1332 2180
rect 1566 2184 1572 2185
rect 1566 2180 1567 2184
rect 1571 2180 1572 2184
rect 1566 2179 1572 2180
rect 1814 2184 1820 2185
rect 1814 2180 1815 2184
rect 1819 2180 1820 2184
rect 1814 2179 1820 2180
rect 1328 2155 1330 2179
rect 1568 2155 1570 2179
rect 1816 2155 1818 2179
rect 1327 2154 1331 2155
rect 1327 2149 1331 2150
rect 1447 2154 1451 2155
rect 1447 2149 1451 2150
rect 1567 2154 1571 2155
rect 1567 2149 1571 2150
rect 1631 2154 1635 2155
rect 1631 2149 1635 2150
rect 1815 2154 1819 2155
rect 1815 2149 1819 2150
rect 1823 2154 1827 2155
rect 1823 2149 1827 2150
rect 1448 2125 1450 2149
rect 1632 2125 1634 2149
rect 1824 2125 1826 2149
rect 1446 2124 1452 2125
rect 1446 2120 1447 2124
rect 1451 2120 1452 2124
rect 1446 2119 1452 2120
rect 1630 2124 1636 2125
rect 1630 2120 1631 2124
rect 1635 2120 1636 2124
rect 1630 2119 1636 2120
rect 1822 2124 1828 2125
rect 1822 2120 1823 2124
rect 1827 2120 1828 2124
rect 1822 2119 1828 2120
rect 1338 2115 1344 2116
rect 1338 2111 1339 2115
rect 1343 2111 1344 2115
rect 1338 2110 1344 2111
rect 1522 2115 1528 2116
rect 1522 2111 1523 2115
rect 1527 2111 1528 2115
rect 1522 2110 1528 2111
rect 1622 2115 1628 2116
rect 1622 2111 1623 2115
rect 1627 2111 1628 2115
rect 1622 2110 1628 2111
rect 1814 2115 1820 2116
rect 1814 2111 1815 2115
rect 1819 2111 1820 2115
rect 1814 2110 1820 2111
rect 1340 2088 1342 2110
rect 1446 2105 1452 2106
rect 1446 2101 1447 2105
rect 1451 2101 1452 2105
rect 1446 2100 1452 2101
rect 1302 2087 1308 2088
rect 1302 2083 1303 2087
rect 1307 2083 1308 2087
rect 1302 2082 1308 2083
rect 1338 2087 1344 2088
rect 1338 2083 1339 2087
rect 1343 2083 1344 2087
rect 1338 2082 1344 2083
rect 1448 2071 1450 2100
rect 1524 2088 1526 2110
rect 1522 2087 1528 2088
rect 1522 2083 1523 2087
rect 1527 2083 1528 2087
rect 1522 2082 1528 2083
rect 1047 2070 1051 2071
rect 1047 2065 1051 2066
rect 1095 2070 1099 2071
rect 1095 2065 1099 2066
rect 1215 2070 1219 2071
rect 1215 2065 1219 2066
rect 1263 2070 1267 2071
rect 1263 2065 1267 2066
rect 1399 2070 1403 2071
rect 1399 2065 1403 2066
rect 1447 2070 1451 2071
rect 1447 2065 1451 2066
rect 1583 2070 1587 2071
rect 1583 2065 1587 2066
rect 1048 2044 1050 2065
rect 1130 2063 1136 2064
rect 1130 2059 1131 2063
rect 1135 2059 1136 2063
rect 1130 2058 1136 2059
rect 1046 2043 1052 2044
rect 1046 2039 1047 2043
rect 1051 2039 1052 2043
rect 1046 2038 1052 2039
rect 1132 2036 1134 2058
rect 1216 2044 1218 2065
rect 1226 2063 1232 2064
rect 1226 2059 1227 2063
rect 1231 2059 1232 2063
rect 1226 2058 1232 2059
rect 1214 2043 1220 2044
rect 1214 2039 1215 2043
rect 1219 2039 1220 2043
rect 1214 2038 1220 2039
rect 450 2035 456 2036
rect 450 2031 451 2035
rect 455 2031 456 2035
rect 450 2030 456 2031
rect 570 2035 576 2036
rect 570 2031 571 2035
rect 575 2031 576 2035
rect 570 2030 576 2031
rect 690 2035 696 2036
rect 690 2031 691 2035
rect 695 2031 696 2035
rect 690 2030 696 2031
rect 826 2035 832 2036
rect 826 2031 827 2035
rect 831 2031 832 2035
rect 826 2030 832 2031
rect 886 2035 892 2036
rect 886 2031 887 2035
rect 891 2031 892 2035
rect 886 2030 892 2031
rect 1002 2035 1008 2036
rect 1002 2031 1003 2035
rect 1007 2031 1008 2035
rect 1002 2030 1008 2031
rect 1130 2035 1136 2036
rect 1130 2031 1131 2035
rect 1135 2031 1136 2035
rect 1130 2030 1136 2031
rect 494 2024 500 2025
rect 494 2020 495 2024
rect 499 2020 500 2024
rect 494 2019 500 2020
rect 614 2024 620 2025
rect 614 2020 615 2024
rect 619 2020 620 2024
rect 614 2019 620 2020
rect 750 2024 756 2025
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 496 1987 498 2019
rect 616 1987 618 2019
rect 752 1987 754 2019
rect 495 1986 499 1987
rect 495 1981 499 1982
rect 511 1986 515 1987
rect 511 1981 515 1982
rect 615 1986 619 1987
rect 615 1981 619 1982
rect 623 1986 627 1987
rect 623 1981 627 1982
rect 743 1986 747 1987
rect 743 1981 747 1982
rect 751 1986 755 1987
rect 751 1981 755 1982
rect 871 1986 875 1987
rect 871 1981 875 1982
rect 512 1957 514 1981
rect 624 1957 626 1981
rect 744 1957 746 1981
rect 872 1957 874 1981
rect 510 1956 516 1957
rect 510 1952 511 1956
rect 515 1952 516 1956
rect 510 1951 516 1952
rect 622 1956 628 1957
rect 622 1952 623 1956
rect 627 1952 628 1956
rect 622 1951 628 1952
rect 742 1956 748 1957
rect 742 1952 743 1956
rect 747 1952 748 1956
rect 742 1951 748 1952
rect 870 1956 876 1957
rect 870 1952 871 1956
rect 875 1952 876 1956
rect 870 1951 876 1952
rect 414 1947 420 1948
rect 414 1943 415 1947
rect 419 1943 420 1947
rect 414 1942 420 1943
rect 594 1947 600 1948
rect 594 1943 595 1947
rect 599 1943 600 1947
rect 594 1942 600 1943
rect 718 1947 724 1948
rect 718 1943 719 1947
rect 723 1943 724 1947
rect 718 1942 724 1943
rect 510 1937 516 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 510 1933 511 1937
rect 515 1933 516 1937
rect 510 1932 516 1933
rect 110 1931 116 1932
rect 112 1903 114 1931
rect 512 1903 514 1932
rect 596 1920 598 1942
rect 622 1937 628 1938
rect 622 1933 623 1937
rect 627 1933 628 1937
rect 622 1932 628 1933
rect 594 1919 600 1920
rect 594 1915 595 1919
rect 599 1915 600 1919
rect 594 1914 600 1915
rect 624 1903 626 1932
rect 720 1920 722 1942
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 870 1937 876 1938
rect 870 1933 871 1937
rect 875 1933 876 1937
rect 870 1932 876 1933
rect 718 1919 724 1920
rect 718 1915 719 1919
rect 723 1915 724 1919
rect 718 1914 724 1915
rect 744 1903 746 1932
rect 872 1903 874 1932
rect 888 1920 890 2030
rect 894 2024 900 2025
rect 894 2020 895 2024
rect 899 2020 900 2024
rect 894 2019 900 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1214 2024 1220 2025
rect 1214 2020 1215 2024
rect 1219 2020 1220 2024
rect 1214 2019 1220 2020
rect 896 1987 898 2019
rect 1048 1987 1050 2019
rect 1216 1987 1218 2019
rect 895 1986 899 1987
rect 895 1981 899 1982
rect 1007 1986 1011 1987
rect 1007 1981 1011 1982
rect 1047 1986 1051 1987
rect 1047 1981 1051 1982
rect 1143 1986 1147 1987
rect 1143 1981 1147 1982
rect 1215 1986 1219 1987
rect 1215 1981 1219 1982
rect 1008 1957 1010 1981
rect 1144 1957 1146 1981
rect 1006 1956 1012 1957
rect 1006 1952 1007 1956
rect 1011 1952 1012 1956
rect 1006 1951 1012 1952
rect 1142 1956 1148 1957
rect 1142 1952 1143 1956
rect 1147 1952 1148 1956
rect 1142 1951 1148 1952
rect 1228 1948 1230 2058
rect 1400 2044 1402 2065
rect 1482 2063 1488 2064
rect 1482 2059 1483 2063
rect 1487 2059 1488 2063
rect 1482 2058 1488 2059
rect 1398 2043 1404 2044
rect 1398 2039 1399 2043
rect 1403 2039 1404 2043
rect 1398 2038 1404 2039
rect 1484 2036 1486 2058
rect 1584 2044 1586 2065
rect 1624 2064 1626 2110
rect 1630 2105 1636 2106
rect 1630 2101 1631 2105
rect 1635 2101 1636 2105
rect 1630 2100 1636 2101
rect 1632 2071 1634 2100
rect 1631 2070 1635 2071
rect 1631 2065 1635 2066
rect 1775 2070 1779 2071
rect 1775 2065 1779 2066
rect 1622 2063 1628 2064
rect 1622 2059 1623 2063
rect 1627 2059 1628 2063
rect 1622 2058 1628 2059
rect 1776 2044 1778 2065
rect 1816 2064 1818 2110
rect 1822 2105 1828 2106
rect 1822 2101 1823 2105
rect 1827 2101 1828 2105
rect 1822 2100 1828 2101
rect 1824 2071 1826 2100
rect 1892 2088 1894 2186
rect 2006 2183 2007 2187
rect 2011 2183 2012 2187
rect 2006 2182 2012 2183
rect 2008 2155 2010 2182
rect 2007 2154 2011 2155
rect 2048 2151 2050 2190
rect 2110 2188 2111 2192
rect 2115 2188 2116 2192
rect 2110 2187 2116 2188
rect 2254 2192 2260 2193
rect 2254 2188 2255 2192
rect 2259 2188 2260 2192
rect 2254 2187 2260 2188
rect 2406 2192 2412 2193
rect 2406 2188 2407 2192
rect 2411 2188 2412 2192
rect 2406 2187 2412 2188
rect 2558 2192 2564 2193
rect 2558 2188 2559 2192
rect 2563 2188 2564 2192
rect 2558 2187 2564 2188
rect 2112 2151 2114 2187
rect 2256 2151 2258 2187
rect 2408 2151 2410 2187
rect 2560 2151 2562 2187
rect 2007 2149 2011 2150
rect 2047 2150 2051 2151
rect 2008 2122 2010 2149
rect 2047 2145 2051 2146
rect 2111 2150 2115 2151
rect 2111 2145 2115 2146
rect 2255 2150 2259 2151
rect 2255 2145 2259 2146
rect 2287 2150 2291 2151
rect 2287 2145 2291 2146
rect 2407 2150 2411 2151
rect 2407 2145 2411 2146
rect 2431 2150 2435 2151
rect 2431 2145 2435 2146
rect 2559 2150 2563 2151
rect 2559 2145 2563 2146
rect 2583 2150 2587 2151
rect 2583 2145 2587 2146
rect 2006 2121 2012 2122
rect 2006 2117 2007 2121
rect 2011 2117 2012 2121
rect 2048 2118 2050 2145
rect 2288 2121 2290 2145
rect 2432 2121 2434 2145
rect 2584 2121 2586 2145
rect 2286 2120 2292 2121
rect 2006 2116 2012 2117
rect 2046 2117 2052 2118
rect 2046 2113 2047 2117
rect 2051 2113 2052 2117
rect 2286 2116 2287 2120
rect 2291 2116 2292 2120
rect 2286 2115 2292 2116
rect 2430 2120 2436 2121
rect 2430 2116 2431 2120
rect 2435 2116 2436 2120
rect 2430 2115 2436 2116
rect 2582 2120 2588 2121
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2046 2112 2052 2113
rect 2660 2112 2662 2226
rect 2720 2212 2722 2233
rect 2880 2212 2882 2233
rect 2954 2231 2960 2232
rect 2954 2227 2955 2231
rect 2959 2227 2960 2231
rect 2954 2226 2960 2227
rect 2718 2211 2724 2212
rect 2718 2207 2719 2211
rect 2723 2207 2724 2211
rect 2718 2206 2724 2207
rect 2878 2211 2884 2212
rect 2878 2207 2879 2211
rect 2883 2207 2884 2211
rect 2878 2206 2884 2207
rect 2956 2204 2958 2226
rect 3048 2212 3050 2233
rect 3122 2231 3128 2232
rect 3122 2227 3123 2231
rect 3127 2227 3128 2231
rect 3122 2226 3128 2227
rect 3046 2211 3052 2212
rect 3046 2207 3047 2211
rect 3051 2207 3052 2211
rect 3046 2206 3052 2207
rect 3124 2204 3126 2226
rect 3224 2212 3226 2233
rect 3298 2231 3304 2232
rect 3298 2227 3299 2231
rect 3303 2227 3304 2231
rect 3298 2226 3304 2227
rect 3222 2211 3228 2212
rect 3222 2207 3223 2211
rect 3227 2207 3228 2211
rect 3222 2206 3228 2207
rect 3300 2204 3302 2226
rect 3408 2212 3410 2233
rect 3482 2231 3488 2232
rect 3482 2227 3483 2231
rect 3487 2227 3488 2231
rect 3482 2226 3488 2227
rect 3406 2211 3412 2212
rect 3406 2207 3407 2211
rect 3411 2207 3412 2211
rect 3406 2206 3412 2207
rect 3484 2204 3486 2226
rect 3592 2212 3594 2233
rect 3590 2211 3596 2212
rect 3590 2207 3591 2211
rect 3595 2207 3596 2211
rect 3590 2206 3596 2207
rect 3748 2204 3750 2414
rect 3840 2399 3842 2436
rect 3839 2398 3843 2399
rect 3839 2393 3843 2394
rect 3839 2322 3843 2323
rect 3839 2317 3843 2318
rect 3840 2293 3842 2317
rect 3838 2292 3844 2293
rect 3838 2288 3839 2292
rect 3843 2288 3844 2292
rect 3838 2287 3844 2288
rect 3838 2273 3844 2274
rect 3838 2269 3839 2273
rect 3843 2269 3844 2273
rect 3838 2268 3844 2269
rect 3840 2239 3842 2268
rect 3908 2256 3910 2446
rect 3924 2424 3926 2610
rect 3942 2604 3948 2605
rect 3942 2600 3943 2604
rect 3947 2600 3948 2604
rect 3942 2599 3948 2600
rect 3944 2571 3946 2599
rect 3943 2570 3947 2571
rect 3943 2565 3947 2566
rect 3944 2545 3946 2565
rect 3942 2544 3948 2545
rect 3942 2540 3943 2544
rect 3947 2540 3948 2544
rect 3942 2539 3948 2540
rect 3942 2527 3948 2528
rect 3942 2523 3943 2527
rect 3947 2523 3948 2527
rect 3942 2522 3948 2523
rect 3944 2491 3946 2522
rect 3943 2490 3947 2491
rect 3943 2485 3947 2486
rect 3944 2458 3946 2485
rect 3942 2457 3948 2458
rect 3942 2453 3943 2457
rect 3947 2453 3948 2457
rect 3942 2452 3948 2453
rect 3942 2440 3948 2441
rect 3942 2436 3943 2440
rect 3947 2436 3948 2440
rect 3942 2435 3948 2436
rect 3922 2423 3928 2424
rect 3922 2419 3923 2423
rect 3927 2419 3928 2423
rect 3922 2418 3928 2419
rect 3944 2399 3946 2435
rect 3943 2398 3947 2399
rect 3943 2393 3947 2394
rect 3944 2373 3946 2393
rect 3942 2372 3948 2373
rect 3942 2368 3943 2372
rect 3947 2368 3948 2372
rect 3942 2367 3948 2368
rect 3942 2355 3948 2356
rect 3942 2351 3943 2355
rect 3947 2351 3948 2355
rect 3942 2350 3948 2351
rect 3944 2323 3946 2350
rect 3943 2322 3947 2323
rect 3943 2317 3947 2318
rect 3944 2290 3946 2317
rect 3942 2289 3948 2290
rect 3942 2285 3943 2289
rect 3947 2285 3948 2289
rect 3942 2284 3948 2285
rect 3914 2283 3920 2284
rect 3914 2279 3915 2283
rect 3919 2279 3920 2283
rect 3914 2278 3920 2279
rect 3906 2255 3912 2256
rect 3906 2251 3907 2255
rect 3911 2251 3912 2255
rect 3906 2250 3912 2251
rect 3783 2238 3787 2239
rect 3783 2233 3787 2234
rect 3839 2238 3843 2239
rect 3839 2233 3843 2234
rect 3784 2212 3786 2233
rect 3866 2231 3872 2232
rect 3866 2227 3867 2231
rect 3871 2227 3872 2231
rect 3866 2226 3872 2227
rect 3782 2211 3788 2212
rect 3782 2207 3783 2211
rect 3787 2207 3788 2211
rect 3782 2206 3788 2207
rect 2954 2203 2960 2204
rect 2954 2199 2955 2203
rect 2959 2199 2960 2203
rect 2954 2198 2960 2199
rect 3122 2203 3128 2204
rect 3122 2199 3123 2203
rect 3127 2199 3128 2203
rect 3122 2198 3128 2199
rect 3298 2203 3304 2204
rect 3298 2199 3299 2203
rect 3303 2199 3304 2203
rect 3298 2198 3304 2199
rect 3482 2203 3488 2204
rect 3482 2199 3483 2203
rect 3487 2199 3488 2203
rect 3482 2198 3488 2199
rect 3558 2203 3564 2204
rect 3558 2199 3559 2203
rect 3563 2199 3564 2203
rect 3558 2198 3564 2199
rect 3746 2203 3752 2204
rect 3746 2199 3747 2203
rect 3751 2199 3752 2203
rect 3746 2198 3752 2199
rect 2718 2192 2724 2193
rect 2718 2188 2719 2192
rect 2723 2188 2724 2192
rect 2718 2187 2724 2188
rect 2878 2192 2884 2193
rect 2878 2188 2879 2192
rect 2883 2188 2884 2192
rect 2878 2187 2884 2188
rect 3046 2192 3052 2193
rect 3046 2188 3047 2192
rect 3051 2188 3052 2192
rect 3046 2187 3052 2188
rect 3222 2192 3228 2193
rect 3222 2188 3223 2192
rect 3227 2188 3228 2192
rect 3222 2187 3228 2188
rect 3406 2192 3412 2193
rect 3406 2188 3407 2192
rect 3411 2188 3412 2192
rect 3406 2187 3412 2188
rect 2720 2151 2722 2187
rect 2880 2151 2882 2187
rect 3048 2151 3050 2187
rect 3224 2151 3226 2187
rect 3408 2151 3410 2187
rect 2719 2150 2723 2151
rect 2719 2145 2723 2146
rect 2735 2150 2739 2151
rect 2735 2145 2739 2146
rect 2879 2150 2883 2151
rect 2879 2145 2883 2146
rect 2887 2150 2891 2151
rect 2887 2145 2891 2146
rect 3047 2150 3051 2151
rect 3047 2145 3051 2146
rect 3207 2150 3211 2151
rect 3207 2145 3211 2146
rect 3223 2150 3227 2151
rect 3223 2145 3227 2146
rect 3367 2150 3371 2151
rect 3367 2145 3371 2146
rect 3407 2150 3411 2151
rect 3407 2145 3411 2146
rect 3527 2150 3531 2151
rect 3527 2145 3531 2146
rect 2736 2121 2738 2145
rect 2888 2121 2890 2145
rect 3048 2121 3050 2145
rect 3086 2143 3092 2144
rect 3086 2139 3087 2143
rect 3091 2139 3092 2143
rect 3086 2138 3092 2139
rect 2734 2120 2740 2121
rect 2734 2116 2735 2120
rect 2739 2116 2740 2120
rect 2734 2115 2740 2116
rect 2886 2120 2892 2121
rect 2886 2116 2887 2120
rect 2891 2116 2892 2120
rect 2886 2115 2892 2116
rect 3046 2120 3052 2121
rect 3046 2116 3047 2120
rect 3051 2116 3052 2120
rect 3046 2115 3052 2116
rect 2362 2111 2368 2112
rect 2362 2107 2363 2111
rect 2367 2107 2368 2111
rect 2362 2106 2368 2107
rect 2506 2111 2512 2112
rect 2506 2107 2507 2111
rect 2511 2107 2512 2111
rect 2506 2106 2512 2107
rect 2658 2111 2664 2112
rect 2658 2107 2659 2111
rect 2663 2107 2664 2111
rect 2658 2106 2664 2107
rect 2666 2111 2672 2112
rect 2666 2107 2667 2111
rect 2671 2107 2672 2111
rect 2666 2106 2672 2107
rect 2818 2111 2824 2112
rect 2818 2107 2819 2111
rect 2823 2107 2824 2111
rect 2818 2106 2824 2107
rect 2006 2104 2012 2105
rect 2006 2100 2007 2104
rect 2011 2100 2012 2104
rect 2286 2101 2292 2102
rect 2006 2099 2012 2100
rect 2046 2100 2052 2101
rect 1890 2087 1896 2088
rect 1890 2083 1891 2087
rect 1895 2083 1896 2087
rect 1890 2082 1896 2083
rect 2008 2071 2010 2099
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2286 2097 2287 2101
rect 2291 2097 2292 2101
rect 2286 2096 2292 2097
rect 2046 2095 2052 2096
rect 1823 2070 1827 2071
rect 1823 2065 1827 2066
rect 2007 2070 2011 2071
rect 2048 2067 2050 2095
rect 2288 2067 2290 2096
rect 2364 2084 2366 2106
rect 2430 2101 2436 2102
rect 2430 2097 2431 2101
rect 2435 2097 2436 2101
rect 2430 2096 2436 2097
rect 2362 2083 2368 2084
rect 2362 2079 2363 2083
rect 2367 2079 2368 2083
rect 2362 2078 2368 2079
rect 2432 2067 2434 2096
rect 2508 2084 2510 2106
rect 2582 2101 2588 2102
rect 2582 2097 2583 2101
rect 2587 2097 2588 2101
rect 2582 2096 2588 2097
rect 2506 2083 2512 2084
rect 2506 2079 2507 2083
rect 2511 2079 2512 2083
rect 2506 2078 2512 2079
rect 2584 2067 2586 2096
rect 2668 2092 2670 2106
rect 2734 2101 2740 2102
rect 2734 2097 2735 2101
rect 2739 2097 2740 2101
rect 2734 2096 2740 2097
rect 2666 2091 2672 2092
rect 2666 2087 2667 2091
rect 2671 2087 2672 2091
rect 2666 2086 2672 2087
rect 2736 2067 2738 2096
rect 2820 2084 2822 2106
rect 2886 2101 2892 2102
rect 2886 2097 2887 2101
rect 2891 2097 2892 2101
rect 2886 2096 2892 2097
rect 3046 2101 3052 2102
rect 3046 2097 3047 2101
rect 3051 2097 3052 2101
rect 3046 2096 3052 2097
rect 2818 2083 2824 2084
rect 2818 2079 2819 2083
rect 2823 2079 2824 2083
rect 2818 2078 2824 2079
rect 2888 2067 2890 2096
rect 2926 2079 2932 2080
rect 2926 2075 2927 2079
rect 2931 2075 2932 2079
rect 2926 2074 2932 2075
rect 2007 2065 2011 2066
rect 2047 2066 2051 2067
rect 1814 2063 1820 2064
rect 1814 2059 1815 2063
rect 1819 2059 1820 2063
rect 1814 2058 1820 2059
rect 2008 2045 2010 2065
rect 2047 2061 2051 2062
rect 2287 2066 2291 2067
rect 2287 2061 2291 2062
rect 2431 2066 2435 2067
rect 2431 2061 2435 2062
rect 2503 2066 2507 2067
rect 2503 2061 2507 2062
rect 2583 2066 2587 2067
rect 2583 2061 2587 2062
rect 2671 2066 2675 2067
rect 2671 2061 2675 2062
rect 2735 2066 2739 2067
rect 2735 2061 2739 2062
rect 2839 2066 2843 2067
rect 2839 2061 2843 2062
rect 2887 2066 2891 2067
rect 2887 2061 2891 2062
rect 2006 2044 2012 2045
rect 1582 2043 1588 2044
rect 1582 2039 1583 2043
rect 1587 2039 1588 2043
rect 1582 2038 1588 2039
rect 1774 2043 1780 2044
rect 1774 2039 1775 2043
rect 1779 2039 1780 2043
rect 2006 2040 2007 2044
rect 2011 2040 2012 2044
rect 2048 2041 2050 2061
rect 2006 2039 2012 2040
rect 2046 2040 2052 2041
rect 2504 2040 2506 2061
rect 2562 2059 2568 2060
rect 2562 2055 2563 2059
rect 2567 2055 2568 2059
rect 2562 2054 2568 2055
rect 1774 2038 1780 2039
rect 2046 2036 2047 2040
rect 2051 2036 2052 2040
rect 1482 2035 1488 2036
rect 1474 2031 1480 2032
rect 1474 2027 1475 2031
rect 1479 2027 1480 2031
rect 1482 2031 1483 2035
rect 1487 2031 1488 2035
rect 1482 2030 1488 2031
rect 1754 2035 1760 2036
rect 2046 2035 2052 2036
rect 2502 2039 2508 2040
rect 2502 2035 2503 2039
rect 2507 2035 2508 2039
rect 1754 2031 1755 2035
rect 1759 2031 1760 2035
rect 2502 2034 2508 2035
rect 1754 2030 1760 2031
rect 1474 2026 1480 2027
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1400 1987 1402 2019
rect 1279 1986 1283 1987
rect 1279 1981 1283 1982
rect 1399 1986 1403 1987
rect 1399 1981 1403 1982
rect 1415 1986 1419 1987
rect 1415 1981 1419 1982
rect 1280 1957 1282 1981
rect 1416 1957 1418 1981
rect 1278 1956 1284 1957
rect 1278 1952 1279 1956
rect 1283 1952 1284 1956
rect 1278 1951 1284 1952
rect 1414 1956 1420 1957
rect 1414 1952 1415 1956
rect 1419 1952 1420 1956
rect 1414 1951 1420 1952
rect 946 1947 952 1948
rect 946 1943 947 1947
rect 951 1943 952 1947
rect 946 1942 952 1943
rect 1082 1947 1088 1948
rect 1082 1943 1083 1947
rect 1087 1943 1088 1947
rect 1082 1942 1088 1943
rect 1226 1947 1232 1948
rect 1226 1943 1227 1947
rect 1231 1943 1232 1947
rect 1226 1942 1232 1943
rect 1346 1947 1352 1948
rect 1346 1943 1347 1947
rect 1351 1943 1352 1947
rect 1346 1942 1352 1943
rect 948 1920 950 1942
rect 1006 1937 1012 1938
rect 1006 1933 1007 1937
rect 1011 1933 1012 1937
rect 1006 1932 1012 1933
rect 886 1919 892 1920
rect 886 1915 887 1919
rect 891 1915 892 1919
rect 886 1914 892 1915
rect 946 1919 952 1920
rect 946 1915 947 1919
rect 951 1915 952 1919
rect 946 1914 952 1915
rect 1008 1903 1010 1932
rect 111 1902 115 1903
rect 111 1897 115 1898
rect 511 1902 515 1903
rect 511 1897 515 1898
rect 551 1902 555 1903
rect 551 1897 555 1898
rect 623 1902 627 1903
rect 623 1897 627 1898
rect 663 1902 667 1903
rect 663 1897 667 1898
rect 743 1902 747 1903
rect 743 1897 747 1898
rect 783 1902 787 1903
rect 783 1897 787 1898
rect 871 1902 875 1903
rect 871 1897 875 1898
rect 911 1902 915 1903
rect 911 1897 915 1898
rect 1007 1902 1011 1903
rect 1007 1897 1011 1898
rect 1047 1902 1051 1903
rect 1047 1897 1051 1898
rect 112 1877 114 1897
rect 110 1876 116 1877
rect 552 1876 554 1897
rect 578 1895 584 1896
rect 578 1891 579 1895
rect 583 1891 584 1895
rect 578 1890 584 1891
rect 646 1895 652 1896
rect 646 1891 647 1895
rect 651 1891 652 1895
rect 646 1890 652 1891
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 550 1875 556 1876
rect 550 1871 551 1875
rect 555 1871 556 1875
rect 550 1870 556 1871
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 110 1854 116 1855
rect 550 1856 556 1857
rect 112 1827 114 1854
rect 550 1852 551 1856
rect 555 1852 556 1856
rect 550 1851 556 1852
rect 552 1827 554 1851
rect 111 1826 115 1827
rect 111 1821 115 1822
rect 503 1826 507 1827
rect 503 1821 507 1822
rect 551 1826 555 1827
rect 551 1821 555 1822
rect 112 1794 114 1821
rect 504 1797 506 1821
rect 502 1796 508 1797
rect 110 1793 116 1794
rect 110 1789 111 1793
rect 115 1789 116 1793
rect 502 1792 503 1796
rect 507 1792 508 1796
rect 502 1791 508 1792
rect 110 1788 116 1789
rect 580 1788 582 1890
rect 648 1868 650 1890
rect 664 1876 666 1897
rect 784 1876 786 1897
rect 858 1895 864 1896
rect 858 1891 859 1895
rect 863 1891 864 1895
rect 858 1890 864 1891
rect 662 1875 668 1876
rect 662 1871 663 1875
rect 667 1871 668 1875
rect 662 1870 668 1871
rect 782 1875 788 1876
rect 782 1871 783 1875
rect 787 1871 788 1875
rect 782 1870 788 1871
rect 860 1868 862 1890
rect 912 1876 914 1897
rect 1048 1876 1050 1897
rect 1084 1896 1086 1942
rect 1142 1937 1148 1938
rect 1142 1933 1143 1937
rect 1147 1933 1148 1937
rect 1142 1932 1148 1933
rect 1278 1937 1284 1938
rect 1278 1933 1279 1937
rect 1283 1933 1284 1937
rect 1278 1932 1284 1933
rect 1144 1903 1146 1932
rect 1280 1903 1282 1932
rect 1143 1902 1147 1903
rect 1143 1897 1147 1898
rect 1175 1902 1179 1903
rect 1175 1897 1179 1898
rect 1279 1902 1283 1903
rect 1279 1897 1283 1898
rect 1311 1902 1315 1903
rect 1311 1897 1315 1898
rect 1082 1895 1088 1896
rect 1082 1891 1083 1895
rect 1087 1891 1088 1895
rect 1082 1890 1088 1891
rect 1176 1876 1178 1897
rect 1214 1895 1220 1896
rect 1214 1891 1215 1895
rect 1219 1894 1220 1895
rect 1219 1891 1222 1894
rect 1214 1890 1222 1891
rect 910 1875 916 1876
rect 910 1871 911 1875
rect 915 1871 916 1875
rect 910 1870 916 1871
rect 1046 1875 1052 1876
rect 1046 1871 1047 1875
rect 1051 1871 1052 1875
rect 1046 1870 1052 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1174 1870 1180 1871
rect 646 1867 652 1868
rect 646 1863 647 1867
rect 651 1863 652 1867
rect 646 1862 652 1863
rect 858 1867 864 1868
rect 858 1863 859 1867
rect 863 1863 864 1867
rect 858 1862 864 1863
rect 1038 1867 1044 1868
rect 1038 1863 1039 1867
rect 1043 1863 1044 1867
rect 1038 1862 1044 1863
rect 662 1856 668 1857
rect 662 1852 663 1856
rect 667 1852 668 1856
rect 662 1851 668 1852
rect 782 1856 788 1857
rect 782 1852 783 1856
rect 787 1852 788 1856
rect 782 1851 788 1852
rect 910 1856 916 1857
rect 910 1852 911 1856
rect 915 1852 916 1856
rect 910 1851 916 1852
rect 664 1827 666 1851
rect 784 1827 786 1851
rect 912 1827 914 1851
rect 615 1826 619 1827
rect 615 1821 619 1822
rect 663 1826 667 1827
rect 663 1821 667 1822
rect 735 1826 739 1827
rect 735 1821 739 1822
rect 783 1826 787 1827
rect 783 1821 787 1822
rect 863 1826 867 1827
rect 863 1821 867 1822
rect 911 1826 915 1827
rect 911 1821 915 1822
rect 999 1826 1003 1827
rect 999 1821 1003 1822
rect 616 1797 618 1821
rect 736 1797 738 1821
rect 864 1797 866 1821
rect 1000 1797 1002 1821
rect 614 1796 620 1797
rect 614 1792 615 1796
rect 619 1792 620 1796
rect 614 1791 620 1792
rect 734 1796 740 1797
rect 734 1792 735 1796
rect 739 1792 740 1796
rect 734 1791 740 1792
rect 862 1796 868 1797
rect 862 1792 863 1796
rect 867 1792 868 1796
rect 862 1791 868 1792
rect 998 1796 1004 1797
rect 998 1792 999 1796
rect 1003 1792 1004 1796
rect 998 1791 1004 1792
rect 578 1787 584 1788
rect 578 1783 579 1787
rect 583 1783 584 1787
rect 578 1782 584 1783
rect 590 1787 596 1788
rect 590 1783 591 1787
rect 595 1783 596 1787
rect 590 1782 596 1783
rect 710 1787 716 1788
rect 710 1783 711 1787
rect 715 1783 716 1787
rect 710 1782 716 1783
rect 930 1787 936 1788
rect 930 1783 931 1787
rect 935 1783 936 1787
rect 930 1782 936 1783
rect 970 1787 976 1788
rect 970 1783 971 1787
rect 975 1783 976 1787
rect 970 1782 976 1783
rect 502 1777 508 1778
rect 110 1776 116 1777
rect 110 1772 111 1776
rect 115 1772 116 1776
rect 502 1773 503 1777
rect 507 1773 508 1777
rect 502 1772 508 1773
rect 110 1771 116 1772
rect 112 1751 114 1771
rect 504 1751 506 1772
rect 592 1760 594 1782
rect 614 1777 620 1778
rect 614 1773 615 1777
rect 619 1773 620 1777
rect 614 1772 620 1773
rect 590 1759 596 1760
rect 590 1755 591 1759
rect 595 1755 596 1759
rect 590 1754 596 1755
rect 616 1751 618 1772
rect 712 1760 714 1782
rect 734 1777 740 1778
rect 734 1773 735 1777
rect 739 1773 740 1777
rect 734 1772 740 1773
rect 862 1777 868 1778
rect 862 1773 863 1777
rect 867 1773 868 1777
rect 862 1772 868 1773
rect 710 1759 716 1760
rect 710 1755 711 1759
rect 715 1755 716 1759
rect 710 1754 716 1755
rect 736 1751 738 1772
rect 794 1755 800 1756
rect 794 1751 795 1755
rect 799 1751 800 1755
rect 864 1751 866 1772
rect 932 1752 934 1782
rect 972 1760 974 1782
rect 998 1777 1004 1778
rect 998 1773 999 1777
rect 1003 1773 1004 1777
rect 998 1772 1004 1773
rect 970 1759 976 1760
rect 970 1755 971 1759
rect 975 1755 976 1759
rect 970 1754 976 1755
rect 930 1751 936 1752
rect 1000 1751 1002 1772
rect 1040 1760 1042 1862
rect 1046 1856 1052 1857
rect 1046 1852 1047 1856
rect 1051 1852 1052 1856
rect 1046 1851 1052 1852
rect 1174 1856 1180 1857
rect 1174 1852 1175 1856
rect 1179 1852 1180 1856
rect 1174 1851 1180 1852
rect 1048 1827 1050 1851
rect 1176 1827 1178 1851
rect 1047 1826 1051 1827
rect 1047 1821 1051 1822
rect 1151 1826 1155 1827
rect 1151 1821 1155 1822
rect 1175 1826 1179 1827
rect 1175 1821 1179 1822
rect 1152 1797 1154 1821
rect 1150 1796 1156 1797
rect 1150 1792 1151 1796
rect 1155 1792 1156 1796
rect 1150 1791 1156 1792
rect 1220 1788 1222 1890
rect 1312 1876 1314 1897
rect 1348 1896 1350 1942
rect 1414 1937 1420 1938
rect 1414 1933 1415 1937
rect 1419 1933 1420 1937
rect 1414 1932 1420 1933
rect 1416 1903 1418 1932
rect 1476 1920 1478 2026
rect 1582 2024 1588 2025
rect 1582 2020 1583 2024
rect 1587 2020 1588 2024
rect 1582 2019 1588 2020
rect 1584 1987 1586 2019
rect 1559 1986 1563 1987
rect 1559 1981 1563 1982
rect 1583 1986 1587 1987
rect 1583 1981 1587 1982
rect 1703 1986 1707 1987
rect 1703 1981 1707 1982
rect 1560 1957 1562 1981
rect 1704 1957 1706 1981
rect 1558 1956 1564 1957
rect 1558 1952 1559 1956
rect 1563 1952 1564 1956
rect 1558 1951 1564 1952
rect 1702 1956 1708 1957
rect 1702 1952 1703 1956
rect 1707 1952 1708 1956
rect 1702 1951 1708 1952
rect 1490 1947 1496 1948
rect 1490 1943 1491 1947
rect 1495 1943 1496 1947
rect 1490 1942 1496 1943
rect 1518 1947 1524 1948
rect 1518 1943 1519 1947
rect 1523 1943 1524 1947
rect 1518 1942 1524 1943
rect 1492 1920 1494 1942
rect 1520 1928 1522 1942
rect 1558 1937 1564 1938
rect 1558 1933 1559 1937
rect 1563 1933 1564 1937
rect 1558 1932 1564 1933
rect 1702 1937 1708 1938
rect 1702 1933 1703 1937
rect 1707 1933 1708 1937
rect 1702 1932 1708 1933
rect 1518 1927 1524 1928
rect 1518 1923 1519 1927
rect 1523 1923 1524 1927
rect 1518 1922 1524 1923
rect 1474 1919 1480 1920
rect 1474 1915 1475 1919
rect 1479 1915 1480 1919
rect 1474 1914 1480 1915
rect 1490 1919 1496 1920
rect 1490 1915 1491 1919
rect 1495 1915 1496 1919
rect 1490 1914 1496 1915
rect 1560 1903 1562 1932
rect 1704 1903 1706 1932
rect 1756 1920 1758 2030
rect 2006 2027 2012 2028
rect 1774 2024 1780 2025
rect 1774 2020 1775 2024
rect 1779 2020 1780 2024
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2006 2022 2012 2023
rect 2046 2023 2052 2024
rect 1774 2019 1780 2020
rect 1776 1987 1778 2019
rect 2008 1987 2010 2022
rect 2046 2019 2047 2023
rect 2051 2019 2052 2023
rect 2046 2018 2052 2019
rect 2502 2020 2508 2021
rect 2048 1987 2050 2018
rect 2502 2016 2503 2020
rect 2507 2016 2508 2020
rect 2502 2015 2508 2016
rect 2504 1987 2506 2015
rect 1775 1986 1779 1987
rect 1775 1981 1779 1982
rect 2007 1986 2011 1987
rect 2007 1981 2011 1982
rect 2047 1986 2051 1987
rect 2047 1981 2051 1982
rect 2495 1986 2499 1987
rect 2495 1981 2499 1982
rect 2503 1986 2507 1987
rect 2503 1981 2507 1982
rect 2008 1954 2010 1981
rect 2048 1954 2050 1981
rect 2496 1957 2498 1981
rect 2494 1956 2500 1957
rect 2006 1953 2012 1954
rect 2006 1949 2007 1953
rect 2011 1949 2012 1953
rect 2006 1948 2012 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2494 1952 2495 1956
rect 2499 1952 2500 1956
rect 2494 1951 2500 1952
rect 2046 1948 2052 1949
rect 2564 1948 2566 2054
rect 2672 2040 2674 2061
rect 2746 2059 2752 2060
rect 2746 2055 2747 2059
rect 2751 2055 2752 2059
rect 2746 2054 2752 2055
rect 2670 2039 2676 2040
rect 2670 2035 2671 2039
rect 2675 2035 2676 2039
rect 2670 2034 2676 2035
rect 2748 2032 2750 2054
rect 2840 2040 2842 2061
rect 2914 2059 2920 2060
rect 2914 2055 2915 2059
rect 2919 2055 2920 2059
rect 2914 2054 2920 2055
rect 2838 2039 2844 2040
rect 2838 2035 2839 2039
rect 2843 2035 2844 2039
rect 2838 2034 2844 2035
rect 2916 2032 2918 2054
rect 2928 2032 2930 2074
rect 3048 2067 3050 2096
rect 3088 2084 3090 2138
rect 3208 2121 3210 2145
rect 3368 2121 3370 2145
rect 3528 2121 3530 2145
rect 3560 2144 3562 2198
rect 3590 2192 3596 2193
rect 3590 2188 3591 2192
rect 3595 2188 3596 2192
rect 3590 2187 3596 2188
rect 3782 2192 3788 2193
rect 3782 2188 3783 2192
rect 3787 2188 3788 2192
rect 3782 2187 3788 2188
rect 3592 2151 3594 2187
rect 3784 2151 3786 2187
rect 3591 2150 3595 2151
rect 3591 2145 3595 2146
rect 3695 2150 3699 2151
rect 3695 2145 3699 2146
rect 3783 2150 3787 2151
rect 3783 2145 3787 2146
rect 3839 2150 3843 2151
rect 3839 2145 3843 2146
rect 3558 2143 3564 2144
rect 3558 2139 3559 2143
rect 3563 2139 3564 2143
rect 3558 2138 3564 2139
rect 3696 2121 3698 2145
rect 3840 2121 3842 2145
rect 3206 2120 3212 2121
rect 3206 2116 3207 2120
rect 3211 2116 3212 2120
rect 3206 2115 3212 2116
rect 3366 2120 3372 2121
rect 3366 2116 3367 2120
rect 3371 2116 3372 2120
rect 3366 2115 3372 2116
rect 3526 2120 3532 2121
rect 3526 2116 3527 2120
rect 3531 2116 3532 2120
rect 3526 2115 3532 2116
rect 3694 2120 3700 2121
rect 3694 2116 3695 2120
rect 3699 2116 3700 2120
rect 3694 2115 3700 2116
rect 3838 2120 3844 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3838 2115 3844 2116
rect 3122 2111 3128 2112
rect 3122 2107 3123 2111
rect 3127 2107 3128 2111
rect 3122 2106 3128 2107
rect 3282 2111 3288 2112
rect 3282 2107 3283 2111
rect 3287 2107 3288 2111
rect 3282 2106 3288 2107
rect 3442 2111 3448 2112
rect 3442 2107 3443 2111
rect 3447 2107 3448 2111
rect 3442 2106 3448 2107
rect 3602 2111 3608 2112
rect 3602 2107 3603 2111
rect 3607 2107 3608 2111
rect 3602 2106 3608 2107
rect 3618 2111 3624 2112
rect 3618 2107 3619 2111
rect 3623 2107 3624 2111
rect 3618 2106 3624 2107
rect 3124 2084 3126 2106
rect 3206 2101 3212 2102
rect 3206 2097 3207 2101
rect 3211 2097 3212 2101
rect 3206 2096 3212 2097
rect 3086 2083 3092 2084
rect 3086 2079 3087 2083
rect 3091 2079 3092 2083
rect 3086 2078 3092 2079
rect 3122 2083 3128 2084
rect 3122 2079 3123 2083
rect 3127 2079 3128 2083
rect 3122 2078 3128 2079
rect 3208 2067 3210 2096
rect 3284 2084 3286 2106
rect 3366 2101 3372 2102
rect 3366 2097 3367 2101
rect 3371 2097 3372 2101
rect 3366 2096 3372 2097
rect 3282 2083 3288 2084
rect 3282 2079 3283 2083
rect 3287 2079 3288 2083
rect 3282 2078 3288 2079
rect 3368 2067 3370 2096
rect 3444 2084 3446 2106
rect 3526 2101 3532 2102
rect 3526 2097 3527 2101
rect 3531 2097 3532 2101
rect 3526 2096 3532 2097
rect 3442 2083 3448 2084
rect 3442 2079 3443 2083
rect 3447 2079 3448 2083
rect 3442 2078 3448 2079
rect 3528 2067 3530 2096
rect 3604 2084 3606 2106
rect 3602 2083 3608 2084
rect 3602 2079 3603 2083
rect 3607 2079 3608 2083
rect 3602 2078 3608 2079
rect 3620 2068 3622 2106
rect 3694 2101 3700 2102
rect 3694 2097 3695 2101
rect 3699 2097 3700 2101
rect 3694 2096 3700 2097
rect 3838 2101 3844 2102
rect 3838 2097 3839 2101
rect 3843 2097 3844 2101
rect 3838 2096 3844 2097
rect 3618 2067 3624 2068
rect 3696 2067 3698 2096
rect 3840 2067 3842 2096
rect 3007 2066 3011 2067
rect 3007 2061 3011 2062
rect 3047 2066 3051 2067
rect 3047 2061 3051 2062
rect 3167 2066 3171 2067
rect 3167 2061 3171 2062
rect 3207 2066 3211 2067
rect 3207 2061 3211 2062
rect 3311 2066 3315 2067
rect 3311 2061 3315 2062
rect 3367 2066 3371 2067
rect 3367 2061 3371 2062
rect 3455 2066 3459 2067
rect 3455 2061 3459 2062
rect 3527 2066 3531 2067
rect 3527 2061 3531 2062
rect 3591 2066 3595 2067
rect 3618 2063 3619 2067
rect 3623 2063 3624 2067
rect 3618 2062 3624 2063
rect 3695 2066 3699 2067
rect 3591 2061 3595 2062
rect 3695 2061 3699 2062
rect 3727 2066 3731 2067
rect 3727 2061 3731 2062
rect 3839 2066 3843 2067
rect 3839 2061 3843 2062
rect 3008 2040 3010 2061
rect 3168 2040 3170 2061
rect 3242 2059 3248 2060
rect 3242 2055 3243 2059
rect 3247 2055 3248 2059
rect 3242 2054 3248 2055
rect 3006 2039 3012 2040
rect 3006 2035 3007 2039
rect 3011 2035 3012 2039
rect 3006 2034 3012 2035
rect 3166 2039 3172 2040
rect 3166 2035 3167 2039
rect 3171 2035 3172 2039
rect 3166 2034 3172 2035
rect 3244 2032 3246 2054
rect 3312 2040 3314 2061
rect 3386 2059 3392 2060
rect 3386 2055 3387 2059
rect 3391 2055 3392 2059
rect 3386 2054 3392 2055
rect 3310 2039 3316 2040
rect 3310 2035 3311 2039
rect 3315 2035 3316 2039
rect 3310 2034 3316 2035
rect 3388 2032 3390 2054
rect 3456 2040 3458 2061
rect 3592 2040 3594 2061
rect 3666 2059 3672 2060
rect 3666 2055 3667 2059
rect 3671 2055 3672 2059
rect 3666 2054 3672 2055
rect 3454 2039 3460 2040
rect 3454 2035 3455 2039
rect 3459 2035 3460 2039
rect 3454 2034 3460 2035
rect 3590 2039 3596 2040
rect 3590 2035 3591 2039
rect 3595 2035 3596 2039
rect 3590 2034 3596 2035
rect 3668 2032 3670 2054
rect 3728 2040 3730 2061
rect 3840 2040 3842 2061
rect 3726 2039 3732 2040
rect 3726 2035 3727 2039
rect 3731 2035 3732 2039
rect 3726 2034 3732 2035
rect 3838 2039 3844 2040
rect 3838 2035 3839 2039
rect 3843 2035 3844 2039
rect 3838 2034 3844 2035
rect 2746 2031 2752 2032
rect 2746 2027 2747 2031
rect 2751 2027 2752 2031
rect 2746 2026 2752 2027
rect 2914 2031 2920 2032
rect 2914 2027 2915 2031
rect 2919 2027 2920 2031
rect 2914 2026 2920 2027
rect 2926 2031 2932 2032
rect 2926 2027 2927 2031
rect 2931 2027 2932 2031
rect 2926 2026 2932 2027
rect 3242 2031 3248 2032
rect 3242 2027 3243 2031
rect 3247 2027 3248 2031
rect 3242 2026 3248 2027
rect 3386 2031 3392 2032
rect 3386 2027 3387 2031
rect 3391 2027 3392 2031
rect 3386 2026 3392 2027
rect 3666 2031 3672 2032
rect 3666 2027 3667 2031
rect 3671 2027 3672 2031
rect 3666 2026 3672 2027
rect 3710 2031 3716 2032
rect 3710 2027 3711 2031
rect 3715 2027 3716 2031
rect 3710 2026 3716 2027
rect 2670 2020 2676 2021
rect 2670 2016 2671 2020
rect 2675 2016 2676 2020
rect 2670 2015 2676 2016
rect 2838 2020 2844 2021
rect 2838 2016 2839 2020
rect 2843 2016 2844 2020
rect 2838 2015 2844 2016
rect 3006 2020 3012 2021
rect 3006 2016 3007 2020
rect 3011 2016 3012 2020
rect 3006 2015 3012 2016
rect 3166 2020 3172 2021
rect 3166 2016 3167 2020
rect 3171 2016 3172 2020
rect 3166 2015 3172 2016
rect 3310 2020 3316 2021
rect 3310 2016 3311 2020
rect 3315 2016 3316 2020
rect 3310 2015 3316 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3590 2020 3596 2021
rect 3590 2016 3591 2020
rect 3595 2016 3596 2020
rect 3590 2015 3596 2016
rect 2672 1987 2674 2015
rect 2840 1987 2842 2015
rect 3008 1987 3010 2015
rect 3168 1987 3170 2015
rect 3312 1987 3314 2015
rect 3456 1987 3458 2015
rect 3592 1987 3594 2015
rect 2591 1986 2595 1987
rect 2591 1981 2595 1982
rect 2671 1986 2675 1987
rect 2671 1981 2675 1982
rect 2695 1986 2699 1987
rect 2695 1981 2699 1982
rect 2807 1986 2811 1987
rect 2807 1981 2811 1982
rect 2839 1986 2843 1987
rect 2839 1981 2843 1982
rect 2927 1986 2931 1987
rect 2927 1981 2931 1982
rect 3007 1986 3011 1987
rect 3007 1981 3011 1982
rect 3047 1986 3051 1987
rect 3047 1981 3051 1982
rect 3167 1986 3171 1987
rect 3167 1981 3171 1982
rect 3175 1986 3179 1987
rect 3175 1981 3179 1982
rect 3295 1986 3299 1987
rect 3295 1981 3299 1982
rect 3311 1986 3315 1987
rect 3311 1981 3315 1982
rect 3415 1986 3419 1987
rect 3415 1981 3419 1982
rect 3455 1986 3459 1987
rect 3455 1981 3459 1982
rect 3543 1986 3547 1987
rect 3543 1981 3547 1982
rect 3591 1986 3595 1987
rect 3591 1981 3595 1982
rect 3671 1986 3675 1987
rect 3671 1981 3675 1982
rect 2592 1957 2594 1981
rect 2696 1957 2698 1981
rect 2808 1957 2810 1981
rect 2928 1957 2930 1981
rect 3048 1957 3050 1981
rect 3176 1957 3178 1981
rect 3296 1957 3298 1981
rect 3416 1957 3418 1981
rect 3544 1957 3546 1981
rect 3672 1957 3674 1981
rect 2590 1956 2596 1957
rect 2590 1952 2591 1956
rect 2595 1952 2596 1956
rect 2590 1951 2596 1952
rect 2694 1956 2700 1957
rect 2694 1952 2695 1956
rect 2699 1952 2700 1956
rect 2694 1951 2700 1952
rect 2806 1956 2812 1957
rect 2806 1952 2807 1956
rect 2811 1952 2812 1956
rect 2806 1951 2812 1952
rect 2926 1956 2932 1957
rect 2926 1952 2927 1956
rect 2931 1952 2932 1956
rect 2926 1951 2932 1952
rect 3046 1956 3052 1957
rect 3046 1952 3047 1956
rect 3051 1952 3052 1956
rect 3046 1951 3052 1952
rect 3174 1956 3180 1957
rect 3174 1952 3175 1956
rect 3179 1952 3180 1956
rect 3174 1951 3180 1952
rect 3294 1956 3300 1957
rect 3294 1952 3295 1956
rect 3299 1952 3300 1956
rect 3294 1951 3300 1952
rect 3414 1956 3420 1957
rect 3414 1952 3415 1956
rect 3419 1952 3420 1956
rect 3414 1951 3420 1952
rect 3542 1956 3548 1957
rect 3542 1952 3543 1956
rect 3547 1952 3548 1956
rect 3542 1951 3548 1952
rect 3670 1956 3676 1957
rect 3670 1952 3671 1956
rect 3675 1952 3676 1956
rect 3670 1951 3676 1952
rect 1770 1947 1776 1948
rect 1770 1943 1771 1947
rect 1775 1943 1776 1947
rect 1770 1942 1776 1943
rect 2562 1947 2568 1948
rect 2562 1943 2563 1947
rect 2567 1943 2568 1947
rect 2562 1942 2568 1943
rect 2578 1947 2584 1948
rect 2578 1943 2579 1947
rect 2583 1943 2584 1947
rect 2578 1942 2584 1943
rect 2682 1947 2688 1948
rect 2682 1943 2683 1947
rect 2687 1943 2688 1947
rect 2682 1942 2688 1943
rect 2778 1947 2784 1948
rect 2778 1943 2779 1947
rect 2783 1943 2784 1947
rect 2778 1942 2784 1943
rect 3002 1947 3008 1948
rect 3002 1943 3003 1947
rect 3007 1943 3008 1947
rect 3002 1942 3008 1943
rect 3122 1947 3128 1948
rect 3122 1943 3123 1947
rect 3127 1943 3128 1947
rect 3122 1942 3128 1943
rect 3130 1947 3136 1948
rect 3130 1943 3131 1947
rect 3135 1943 3136 1947
rect 3130 1942 3136 1943
rect 3258 1947 3264 1948
rect 3258 1943 3259 1947
rect 3263 1943 3264 1947
rect 3258 1942 3264 1943
rect 3386 1947 3392 1948
rect 3386 1943 3387 1947
rect 3391 1943 3392 1947
rect 3386 1942 3392 1943
rect 3630 1947 3636 1948
rect 3630 1943 3631 1947
rect 3635 1943 3636 1947
rect 3630 1942 3636 1943
rect 1754 1919 1760 1920
rect 1754 1915 1755 1919
rect 1759 1915 1760 1919
rect 1754 1914 1760 1915
rect 1415 1902 1419 1903
rect 1415 1897 1419 1898
rect 1447 1902 1451 1903
rect 1447 1897 1451 1898
rect 1559 1902 1563 1903
rect 1559 1897 1563 1898
rect 1583 1902 1587 1903
rect 1583 1897 1587 1898
rect 1703 1902 1707 1903
rect 1703 1897 1707 1898
rect 1719 1902 1723 1903
rect 1719 1897 1723 1898
rect 1346 1895 1352 1896
rect 1346 1891 1347 1895
rect 1351 1891 1352 1895
rect 1346 1890 1352 1891
rect 1386 1895 1392 1896
rect 1386 1891 1387 1895
rect 1391 1891 1392 1895
rect 1386 1890 1392 1891
rect 1310 1875 1316 1876
rect 1310 1871 1311 1875
rect 1315 1871 1316 1875
rect 1310 1870 1316 1871
rect 1388 1868 1390 1890
rect 1448 1876 1450 1897
rect 1522 1895 1528 1896
rect 1522 1891 1523 1895
rect 1527 1891 1528 1895
rect 1522 1890 1528 1891
rect 1446 1875 1452 1876
rect 1446 1871 1447 1875
rect 1451 1871 1452 1875
rect 1446 1870 1452 1871
rect 1524 1868 1526 1890
rect 1584 1876 1586 1897
rect 1720 1876 1722 1897
rect 1772 1896 1774 1942
rect 2494 1937 2500 1938
rect 2006 1936 2012 1937
rect 2006 1932 2007 1936
rect 2011 1932 2012 1936
rect 2006 1931 2012 1932
rect 2046 1936 2052 1937
rect 2046 1932 2047 1936
rect 2051 1932 2052 1936
rect 2494 1933 2495 1937
rect 2499 1933 2500 1937
rect 2494 1932 2500 1933
rect 2046 1931 2052 1932
rect 2008 1903 2010 1931
rect 2048 1907 2050 1931
rect 2496 1907 2498 1932
rect 2580 1920 2582 1942
rect 2590 1937 2596 1938
rect 2590 1933 2591 1937
rect 2595 1933 2596 1937
rect 2590 1932 2596 1933
rect 2578 1919 2584 1920
rect 2578 1915 2579 1919
rect 2583 1915 2584 1919
rect 2578 1914 2584 1915
rect 2592 1907 2594 1932
rect 2684 1920 2686 1942
rect 2694 1937 2700 1938
rect 2694 1933 2695 1937
rect 2699 1933 2700 1937
rect 2694 1932 2700 1933
rect 2682 1919 2688 1920
rect 2682 1915 2683 1919
rect 2687 1915 2688 1919
rect 2682 1914 2688 1915
rect 2696 1907 2698 1932
rect 2780 1920 2782 1942
rect 2806 1937 2812 1938
rect 2806 1933 2807 1937
rect 2811 1933 2812 1937
rect 2806 1932 2812 1933
rect 2926 1937 2932 1938
rect 2926 1933 2927 1937
rect 2931 1933 2932 1937
rect 2926 1932 2932 1933
rect 2778 1919 2784 1920
rect 2778 1915 2779 1919
rect 2783 1915 2784 1919
rect 2778 1914 2784 1915
rect 2808 1907 2810 1932
rect 2866 1915 2872 1916
rect 2866 1911 2867 1915
rect 2871 1911 2872 1915
rect 2866 1910 2872 1911
rect 2047 1906 2051 1907
rect 2007 1902 2011 1903
rect 1922 1899 1928 1900
rect 1770 1895 1776 1896
rect 1770 1891 1771 1895
rect 1775 1891 1776 1895
rect 1922 1895 1923 1899
rect 1927 1895 1928 1899
rect 2047 1901 2051 1902
rect 2071 1906 2075 1907
rect 2071 1901 2075 1902
rect 2247 1906 2251 1907
rect 2247 1901 2251 1902
rect 2439 1906 2443 1907
rect 2439 1901 2443 1902
rect 2495 1906 2499 1907
rect 2495 1901 2499 1902
rect 2591 1906 2595 1907
rect 2591 1901 2595 1902
rect 2623 1906 2627 1907
rect 2623 1901 2627 1902
rect 2695 1906 2699 1907
rect 2695 1901 2699 1902
rect 2791 1906 2795 1907
rect 2791 1901 2795 1902
rect 2807 1906 2811 1907
rect 2807 1901 2811 1902
rect 2007 1897 2011 1898
rect 1922 1894 1928 1895
rect 1770 1890 1776 1891
rect 1582 1875 1588 1876
rect 1582 1871 1583 1875
rect 1587 1871 1588 1875
rect 1582 1870 1588 1871
rect 1718 1875 1724 1876
rect 1718 1871 1719 1875
rect 1723 1871 1724 1875
rect 1718 1870 1724 1871
rect 1386 1867 1392 1868
rect 1386 1863 1387 1867
rect 1391 1863 1392 1867
rect 1386 1862 1392 1863
rect 1522 1867 1528 1868
rect 1522 1863 1523 1867
rect 1527 1863 1528 1867
rect 1522 1862 1528 1863
rect 1702 1867 1708 1868
rect 1702 1863 1703 1867
rect 1707 1863 1708 1867
rect 1702 1862 1708 1863
rect 1310 1856 1316 1857
rect 1310 1852 1311 1856
rect 1315 1852 1316 1856
rect 1310 1851 1316 1852
rect 1446 1856 1452 1857
rect 1446 1852 1447 1856
rect 1451 1852 1452 1856
rect 1446 1851 1452 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1312 1827 1314 1851
rect 1448 1827 1450 1851
rect 1584 1827 1586 1851
rect 1311 1826 1315 1827
rect 1311 1821 1315 1822
rect 1319 1826 1323 1827
rect 1319 1821 1323 1822
rect 1447 1826 1451 1827
rect 1447 1821 1451 1822
rect 1487 1826 1491 1827
rect 1487 1821 1491 1822
rect 1583 1826 1587 1827
rect 1583 1821 1587 1822
rect 1663 1826 1667 1827
rect 1663 1821 1667 1822
rect 1320 1797 1322 1821
rect 1488 1797 1490 1821
rect 1664 1797 1666 1821
rect 1318 1796 1324 1797
rect 1318 1792 1319 1796
rect 1323 1792 1324 1796
rect 1318 1791 1324 1792
rect 1486 1796 1492 1797
rect 1486 1792 1487 1796
rect 1491 1792 1492 1796
rect 1486 1791 1492 1792
rect 1662 1796 1668 1797
rect 1662 1792 1663 1796
rect 1667 1792 1668 1796
rect 1662 1791 1668 1792
rect 1218 1787 1224 1788
rect 1218 1783 1219 1787
rect 1223 1783 1224 1787
rect 1218 1782 1224 1783
rect 1262 1787 1268 1788
rect 1262 1783 1263 1787
rect 1267 1783 1268 1787
rect 1262 1782 1268 1783
rect 1562 1787 1568 1788
rect 1562 1783 1563 1787
rect 1567 1783 1568 1787
rect 1562 1782 1568 1783
rect 1150 1777 1156 1778
rect 1150 1773 1151 1777
rect 1155 1773 1156 1777
rect 1150 1772 1156 1773
rect 1038 1759 1044 1760
rect 1038 1755 1039 1759
rect 1043 1755 1044 1759
rect 1038 1754 1044 1755
rect 1152 1751 1154 1772
rect 1264 1760 1266 1782
rect 1318 1777 1324 1778
rect 1318 1773 1319 1777
rect 1323 1773 1324 1777
rect 1318 1772 1324 1773
rect 1486 1777 1492 1778
rect 1486 1773 1487 1777
rect 1491 1773 1492 1777
rect 1486 1772 1492 1773
rect 1262 1759 1268 1760
rect 1262 1755 1263 1759
rect 1267 1755 1268 1759
rect 1262 1754 1268 1755
rect 1320 1751 1322 1772
rect 1358 1755 1364 1756
rect 1358 1751 1359 1755
rect 1363 1751 1366 1755
rect 1488 1751 1490 1772
rect 111 1750 115 1751
rect 111 1745 115 1746
rect 343 1750 347 1751
rect 343 1745 347 1746
rect 463 1750 467 1751
rect 463 1745 467 1746
rect 503 1750 507 1751
rect 503 1745 507 1746
rect 591 1750 595 1751
rect 591 1745 595 1746
rect 615 1750 619 1751
rect 615 1745 619 1746
rect 719 1750 723 1751
rect 719 1745 723 1746
rect 735 1750 739 1751
rect 794 1750 800 1751
rect 847 1750 851 1751
rect 735 1745 739 1746
rect 112 1725 114 1745
rect 110 1724 116 1725
rect 344 1724 346 1745
rect 418 1743 424 1744
rect 418 1739 419 1743
rect 423 1739 424 1743
rect 418 1738 424 1739
rect 110 1720 111 1724
rect 115 1720 116 1724
rect 110 1719 116 1720
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1719 348 1723
rect 342 1718 348 1719
rect 420 1716 422 1738
rect 464 1724 466 1745
rect 538 1743 544 1744
rect 538 1739 539 1743
rect 543 1739 544 1743
rect 538 1738 544 1739
rect 462 1723 468 1724
rect 462 1719 463 1723
rect 467 1719 468 1723
rect 462 1718 468 1719
rect 540 1716 542 1738
rect 592 1724 594 1745
rect 666 1743 672 1744
rect 666 1739 667 1743
rect 671 1739 672 1743
rect 666 1738 672 1739
rect 590 1723 596 1724
rect 590 1719 591 1723
rect 595 1719 596 1723
rect 590 1718 596 1719
rect 668 1716 670 1738
rect 720 1724 722 1745
rect 738 1735 744 1736
rect 738 1731 739 1735
rect 743 1731 744 1735
rect 738 1730 744 1731
rect 718 1723 724 1724
rect 718 1719 719 1723
rect 723 1719 724 1723
rect 718 1718 724 1719
rect 418 1715 424 1716
rect 418 1711 419 1715
rect 423 1711 424 1715
rect 418 1710 424 1711
rect 538 1715 544 1716
rect 538 1711 539 1715
rect 543 1711 544 1715
rect 538 1710 544 1711
rect 666 1715 672 1716
rect 666 1711 667 1715
rect 671 1711 672 1715
rect 666 1710 672 1711
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 110 1702 116 1703
rect 342 1704 348 1705
rect 112 1671 114 1702
rect 342 1700 343 1704
rect 347 1700 348 1704
rect 342 1699 348 1700
rect 462 1704 468 1705
rect 462 1700 463 1704
rect 467 1700 468 1704
rect 462 1699 468 1700
rect 590 1704 596 1705
rect 590 1700 591 1704
rect 595 1700 596 1704
rect 590 1699 596 1700
rect 718 1704 724 1705
rect 718 1700 719 1704
rect 723 1700 724 1704
rect 718 1699 724 1700
rect 344 1671 346 1699
rect 464 1671 466 1699
rect 592 1671 594 1699
rect 720 1671 722 1699
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 159 1670 163 1671
rect 159 1665 163 1666
rect 295 1670 299 1671
rect 295 1665 299 1666
rect 343 1670 347 1671
rect 343 1665 347 1666
rect 455 1670 459 1671
rect 455 1665 459 1666
rect 463 1670 467 1671
rect 463 1665 467 1666
rect 591 1670 595 1671
rect 591 1665 595 1666
rect 623 1670 627 1671
rect 623 1665 627 1666
rect 719 1670 723 1671
rect 719 1665 723 1666
rect 112 1638 114 1665
rect 160 1641 162 1665
rect 296 1641 298 1665
rect 456 1641 458 1665
rect 624 1641 626 1665
rect 158 1640 164 1641
rect 110 1637 116 1638
rect 110 1633 111 1637
rect 115 1633 116 1637
rect 158 1636 159 1640
rect 163 1636 164 1640
rect 158 1635 164 1636
rect 294 1640 300 1641
rect 294 1636 295 1640
rect 299 1636 300 1640
rect 294 1635 300 1636
rect 454 1640 460 1641
rect 454 1636 455 1640
rect 459 1636 460 1640
rect 454 1635 460 1636
rect 622 1640 628 1641
rect 622 1636 623 1640
rect 627 1636 628 1640
rect 622 1635 628 1636
rect 110 1632 116 1633
rect 740 1632 742 1730
rect 796 1716 798 1750
rect 847 1745 851 1746
rect 863 1750 867 1751
rect 930 1747 931 1751
rect 935 1747 936 1751
rect 930 1746 936 1747
rect 983 1750 987 1751
rect 863 1745 867 1746
rect 983 1745 987 1746
rect 999 1750 1003 1751
rect 999 1745 1003 1746
rect 1127 1750 1131 1751
rect 1127 1745 1131 1746
rect 1151 1750 1155 1751
rect 1151 1745 1155 1746
rect 1279 1750 1283 1751
rect 1279 1745 1283 1746
rect 1319 1750 1323 1751
rect 1358 1750 1366 1751
rect 1319 1745 1323 1746
rect 848 1724 850 1745
rect 922 1743 928 1744
rect 922 1739 923 1743
rect 927 1739 928 1743
rect 922 1738 928 1739
rect 846 1723 852 1724
rect 846 1719 847 1723
rect 851 1719 852 1723
rect 846 1718 852 1719
rect 924 1716 926 1738
rect 984 1724 986 1745
rect 1128 1724 1130 1745
rect 1158 1743 1164 1744
rect 1158 1739 1159 1743
rect 1163 1739 1164 1743
rect 1158 1738 1164 1739
rect 1202 1743 1208 1744
rect 1202 1739 1203 1743
rect 1207 1739 1208 1743
rect 1202 1738 1208 1739
rect 982 1723 988 1724
rect 982 1719 983 1723
rect 987 1719 988 1723
rect 982 1718 988 1719
rect 1126 1723 1132 1724
rect 1126 1719 1127 1723
rect 1131 1719 1132 1723
rect 1126 1718 1132 1719
rect 794 1715 800 1716
rect 794 1711 795 1715
rect 799 1711 800 1715
rect 794 1710 800 1711
rect 922 1715 928 1716
rect 922 1711 923 1715
rect 927 1711 928 1715
rect 922 1710 928 1711
rect 1058 1711 1064 1712
rect 1058 1707 1059 1711
rect 1063 1707 1064 1711
rect 1058 1706 1064 1707
rect 846 1704 852 1705
rect 846 1700 847 1704
rect 851 1700 852 1704
rect 846 1699 852 1700
rect 982 1704 988 1705
rect 982 1700 983 1704
rect 987 1700 988 1704
rect 982 1699 988 1700
rect 848 1671 850 1699
rect 984 1671 986 1699
rect 799 1670 803 1671
rect 799 1665 803 1666
rect 847 1670 851 1671
rect 847 1665 851 1666
rect 983 1670 987 1671
rect 983 1665 987 1666
rect 800 1641 802 1665
rect 984 1641 986 1665
rect 798 1640 804 1641
rect 798 1636 799 1640
rect 803 1636 804 1640
rect 798 1635 804 1636
rect 982 1640 988 1641
rect 982 1636 983 1640
rect 987 1636 988 1640
rect 982 1635 988 1636
rect 234 1631 240 1632
rect 234 1627 235 1631
rect 239 1627 240 1631
rect 234 1626 240 1627
rect 370 1631 376 1632
rect 370 1627 371 1631
rect 375 1627 376 1631
rect 370 1626 376 1627
rect 530 1631 536 1632
rect 530 1627 531 1631
rect 535 1627 536 1631
rect 530 1626 536 1627
rect 698 1631 704 1632
rect 698 1627 699 1631
rect 703 1627 704 1631
rect 698 1626 704 1627
rect 738 1631 744 1632
rect 738 1627 739 1631
rect 743 1627 744 1631
rect 738 1626 744 1627
rect 1050 1631 1056 1632
rect 1050 1627 1051 1631
rect 1055 1627 1056 1631
rect 1050 1626 1056 1627
rect 158 1621 164 1622
rect 110 1620 116 1621
rect 110 1616 111 1620
rect 115 1616 116 1620
rect 158 1617 159 1621
rect 163 1617 164 1621
rect 158 1616 164 1617
rect 110 1615 116 1616
rect 112 1595 114 1615
rect 160 1595 162 1616
rect 236 1608 238 1626
rect 294 1621 300 1622
rect 294 1617 295 1621
rect 299 1617 300 1621
rect 294 1616 300 1617
rect 234 1607 240 1608
rect 234 1603 235 1607
rect 239 1603 240 1607
rect 234 1602 240 1603
rect 296 1595 298 1616
rect 372 1604 374 1626
rect 454 1621 460 1622
rect 454 1617 455 1621
rect 459 1617 460 1621
rect 454 1616 460 1617
rect 370 1603 376 1604
rect 370 1599 371 1603
rect 375 1599 376 1603
rect 370 1598 376 1599
rect 456 1595 458 1616
rect 532 1604 534 1626
rect 622 1621 628 1622
rect 622 1617 623 1621
rect 627 1617 628 1621
rect 622 1616 628 1617
rect 530 1603 536 1604
rect 530 1599 531 1603
rect 535 1599 536 1603
rect 530 1598 536 1599
rect 624 1595 626 1616
rect 700 1604 702 1626
rect 798 1621 804 1622
rect 798 1617 799 1621
rect 803 1617 804 1621
rect 798 1616 804 1617
rect 982 1621 988 1622
rect 982 1617 983 1621
rect 987 1617 988 1621
rect 982 1616 988 1617
rect 698 1603 704 1604
rect 698 1599 699 1603
rect 703 1599 704 1603
rect 698 1598 704 1599
rect 738 1595 744 1596
rect 800 1595 802 1616
rect 984 1595 986 1616
rect 111 1594 115 1595
rect 111 1589 115 1590
rect 135 1594 139 1595
rect 135 1589 139 1590
rect 159 1594 163 1595
rect 159 1589 163 1590
rect 255 1594 259 1595
rect 255 1589 259 1590
rect 295 1594 299 1595
rect 295 1589 299 1590
rect 423 1594 427 1595
rect 423 1589 427 1590
rect 455 1594 459 1595
rect 455 1589 459 1590
rect 607 1594 611 1595
rect 607 1589 611 1590
rect 623 1594 627 1595
rect 738 1591 739 1595
rect 743 1591 744 1595
rect 738 1590 744 1591
rect 799 1594 803 1595
rect 623 1589 627 1590
rect 112 1569 114 1589
rect 110 1568 116 1569
rect 136 1568 138 1589
rect 202 1587 208 1588
rect 202 1583 203 1587
rect 207 1583 208 1587
rect 202 1582 208 1583
rect 210 1587 216 1588
rect 210 1583 211 1587
rect 215 1583 216 1587
rect 210 1582 216 1583
rect 110 1564 111 1568
rect 115 1564 116 1568
rect 110 1563 116 1564
rect 134 1567 140 1568
rect 134 1563 135 1567
rect 139 1563 140 1567
rect 134 1562 140 1563
rect 110 1551 116 1552
rect 110 1547 111 1551
rect 115 1547 116 1551
rect 110 1546 116 1547
rect 134 1548 140 1549
rect 112 1515 114 1546
rect 134 1544 135 1548
rect 139 1544 140 1548
rect 134 1543 140 1544
rect 136 1515 138 1543
rect 111 1514 115 1515
rect 111 1509 115 1510
rect 135 1514 139 1515
rect 135 1509 139 1510
rect 112 1482 114 1509
rect 136 1485 138 1509
rect 204 1492 206 1582
rect 212 1560 214 1582
rect 256 1568 258 1589
rect 330 1587 336 1588
rect 330 1583 331 1587
rect 335 1583 336 1587
rect 330 1582 336 1583
rect 254 1567 260 1568
rect 254 1563 255 1567
rect 259 1563 260 1567
rect 254 1562 260 1563
rect 332 1560 334 1582
rect 424 1568 426 1589
rect 498 1587 504 1588
rect 498 1583 499 1587
rect 503 1583 504 1587
rect 498 1582 504 1583
rect 422 1567 428 1568
rect 422 1563 423 1567
rect 427 1563 428 1567
rect 422 1562 428 1563
rect 500 1560 502 1582
rect 608 1568 610 1589
rect 682 1587 688 1588
rect 682 1583 683 1587
rect 687 1583 688 1587
rect 682 1582 688 1583
rect 606 1567 612 1568
rect 606 1563 607 1567
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 684 1560 686 1582
rect 740 1560 742 1590
rect 799 1589 803 1590
rect 983 1594 987 1595
rect 983 1589 987 1590
rect 991 1594 995 1595
rect 991 1589 995 1590
rect 800 1568 802 1589
rect 992 1568 994 1589
rect 1052 1588 1054 1626
rect 1060 1604 1062 1706
rect 1126 1704 1132 1705
rect 1126 1700 1127 1704
rect 1131 1700 1132 1704
rect 1126 1699 1132 1700
rect 1128 1671 1130 1699
rect 1127 1670 1131 1671
rect 1127 1665 1131 1666
rect 1160 1632 1162 1738
rect 1204 1716 1206 1738
rect 1280 1724 1282 1745
rect 1354 1743 1360 1744
rect 1354 1739 1355 1743
rect 1359 1739 1360 1743
rect 1354 1738 1360 1739
rect 1278 1723 1284 1724
rect 1278 1719 1279 1723
rect 1283 1719 1284 1723
rect 1278 1718 1284 1719
rect 1356 1716 1358 1738
rect 1364 1716 1366 1750
rect 1439 1750 1443 1751
rect 1439 1745 1443 1746
rect 1487 1750 1491 1751
rect 1487 1745 1491 1746
rect 1440 1724 1442 1745
rect 1564 1744 1566 1782
rect 1662 1777 1668 1778
rect 1662 1773 1663 1777
rect 1667 1773 1668 1777
rect 1662 1772 1668 1773
rect 1664 1751 1666 1772
rect 1704 1760 1706 1862
rect 1710 1859 1716 1860
rect 1710 1855 1711 1859
rect 1715 1855 1716 1859
rect 1710 1854 1716 1855
rect 1718 1856 1724 1857
rect 1712 1760 1714 1854
rect 1718 1852 1719 1856
rect 1723 1852 1724 1856
rect 1718 1851 1724 1852
rect 1720 1827 1722 1851
rect 1719 1826 1723 1827
rect 1719 1821 1723 1822
rect 1847 1826 1851 1827
rect 1847 1821 1851 1822
rect 1848 1797 1850 1821
rect 1846 1796 1852 1797
rect 1846 1792 1847 1796
rect 1851 1792 1852 1796
rect 1846 1791 1852 1792
rect 1924 1788 1926 1894
rect 2008 1877 2010 1897
rect 2048 1881 2050 1901
rect 2046 1880 2052 1881
rect 2072 1880 2074 1901
rect 2248 1880 2250 1901
rect 2322 1899 2328 1900
rect 2322 1895 2323 1899
rect 2327 1895 2328 1899
rect 2322 1894 2328 1895
rect 2006 1876 2012 1877
rect 2006 1872 2007 1876
rect 2011 1872 2012 1876
rect 2046 1876 2047 1880
rect 2051 1876 2052 1880
rect 2046 1875 2052 1876
rect 2070 1879 2076 1880
rect 2070 1875 2071 1879
rect 2075 1875 2076 1879
rect 2070 1874 2076 1875
rect 2246 1879 2252 1880
rect 2246 1875 2247 1879
rect 2251 1875 2252 1879
rect 2246 1874 2252 1875
rect 2324 1872 2326 1894
rect 2440 1880 2442 1901
rect 2514 1899 2520 1900
rect 2514 1895 2515 1899
rect 2519 1895 2520 1899
rect 2514 1894 2520 1895
rect 2478 1891 2484 1892
rect 2478 1887 2479 1891
rect 2483 1887 2484 1891
rect 2478 1886 2484 1887
rect 2438 1879 2444 1880
rect 2438 1875 2439 1879
rect 2443 1875 2444 1879
rect 2438 1874 2444 1875
rect 2006 1871 2012 1872
rect 2322 1871 2328 1872
rect 2146 1867 2152 1868
rect 2046 1863 2052 1864
rect 2006 1859 2012 1860
rect 2006 1855 2007 1859
rect 2011 1855 2012 1859
rect 2046 1859 2047 1863
rect 2051 1859 2052 1863
rect 2146 1863 2147 1867
rect 2151 1863 2152 1867
rect 2322 1867 2323 1871
rect 2327 1867 2328 1871
rect 2322 1866 2328 1867
rect 2146 1862 2152 1863
rect 2046 1858 2052 1859
rect 2070 1860 2076 1861
rect 2006 1854 2012 1855
rect 2008 1827 2010 1854
rect 2048 1831 2050 1858
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2070 1855 2076 1856
rect 2072 1831 2074 1855
rect 2047 1830 2051 1831
rect 2007 1826 2011 1827
rect 2047 1825 2051 1826
rect 2071 1830 2075 1831
rect 2071 1825 2075 1826
rect 2095 1830 2099 1831
rect 2095 1825 2099 1826
rect 2007 1821 2011 1822
rect 2008 1794 2010 1821
rect 2048 1798 2050 1825
rect 2096 1801 2098 1825
rect 2094 1800 2100 1801
rect 2046 1797 2052 1798
rect 2006 1793 2012 1794
rect 2006 1789 2007 1793
rect 2011 1789 2012 1793
rect 2046 1793 2047 1797
rect 2051 1793 2052 1797
rect 2094 1796 2095 1800
rect 2099 1796 2100 1800
rect 2094 1795 2100 1796
rect 2046 1792 2052 1793
rect 2006 1788 2012 1789
rect 1922 1787 1928 1788
rect 1922 1783 1923 1787
rect 1927 1783 1928 1787
rect 1922 1782 1928 1783
rect 2094 1781 2100 1782
rect 2046 1780 2052 1781
rect 1846 1777 1852 1778
rect 1846 1773 1847 1777
rect 1851 1773 1852 1777
rect 1846 1772 1852 1773
rect 2006 1776 2012 1777
rect 2006 1772 2007 1776
rect 2011 1772 2012 1776
rect 2046 1776 2047 1780
rect 2051 1776 2052 1780
rect 2094 1777 2095 1781
rect 2099 1777 2100 1781
rect 2094 1776 2100 1777
rect 2046 1775 2052 1776
rect 1702 1759 1708 1760
rect 1702 1755 1703 1759
rect 1707 1755 1708 1759
rect 1702 1754 1708 1755
rect 1710 1759 1716 1760
rect 1710 1755 1711 1759
rect 1715 1755 1716 1759
rect 1710 1754 1716 1755
rect 1848 1751 1850 1772
rect 2006 1771 2012 1772
rect 2008 1751 2010 1771
rect 2048 1755 2050 1775
rect 2096 1755 2098 1776
rect 2148 1764 2150 1862
rect 2246 1860 2252 1861
rect 2246 1856 2247 1860
rect 2251 1856 2252 1860
rect 2246 1855 2252 1856
rect 2438 1860 2444 1861
rect 2438 1856 2439 1860
rect 2443 1856 2444 1860
rect 2438 1855 2444 1856
rect 2248 1831 2250 1855
rect 2440 1831 2442 1855
rect 2231 1830 2235 1831
rect 2231 1825 2235 1826
rect 2247 1830 2251 1831
rect 2247 1825 2251 1826
rect 2367 1830 2371 1831
rect 2367 1825 2371 1826
rect 2439 1830 2443 1831
rect 2439 1825 2443 1826
rect 2232 1801 2234 1825
rect 2368 1801 2370 1825
rect 2230 1800 2236 1801
rect 2230 1796 2231 1800
rect 2235 1796 2236 1800
rect 2230 1795 2236 1796
rect 2366 1800 2372 1801
rect 2366 1796 2367 1800
rect 2371 1796 2372 1800
rect 2366 1795 2372 1796
rect 2480 1792 2482 1886
rect 2516 1872 2518 1894
rect 2624 1880 2626 1901
rect 2792 1880 2794 1901
rect 2622 1879 2628 1880
rect 2622 1875 2623 1879
rect 2627 1875 2628 1879
rect 2622 1874 2628 1875
rect 2790 1879 2796 1880
rect 2790 1875 2791 1879
rect 2795 1875 2796 1879
rect 2790 1874 2796 1875
rect 2868 1872 2870 1910
rect 2928 1907 2930 1932
rect 3004 1920 3006 1942
rect 3046 1937 3052 1938
rect 3046 1933 3047 1937
rect 3051 1933 3052 1937
rect 3046 1932 3052 1933
rect 3002 1919 3008 1920
rect 3002 1915 3003 1919
rect 3007 1915 3008 1919
rect 3002 1914 3008 1915
rect 3048 1907 3050 1932
rect 3124 1920 3126 1942
rect 3132 1928 3134 1942
rect 3174 1937 3180 1938
rect 3174 1933 3175 1937
rect 3179 1933 3180 1937
rect 3174 1932 3180 1933
rect 3130 1927 3136 1928
rect 3130 1923 3131 1927
rect 3135 1923 3136 1927
rect 3130 1922 3136 1923
rect 3122 1919 3128 1920
rect 3122 1915 3123 1919
rect 3127 1915 3128 1919
rect 3122 1914 3128 1915
rect 3176 1907 3178 1932
rect 3260 1908 3262 1942
rect 3294 1937 3300 1938
rect 3294 1933 3295 1937
rect 3299 1933 3300 1937
rect 3294 1932 3300 1933
rect 3258 1907 3264 1908
rect 3296 1907 3298 1932
rect 3388 1920 3390 1942
rect 3414 1937 3420 1938
rect 3414 1933 3415 1937
rect 3419 1933 3420 1937
rect 3414 1932 3420 1933
rect 3542 1937 3548 1938
rect 3542 1933 3543 1937
rect 3547 1933 3548 1937
rect 3542 1932 3548 1933
rect 3386 1919 3392 1920
rect 3386 1915 3387 1919
rect 3391 1915 3392 1919
rect 3386 1914 3392 1915
rect 3416 1907 3418 1932
rect 3544 1907 3546 1932
rect 3632 1920 3634 1942
rect 3670 1937 3676 1938
rect 3670 1933 3671 1937
rect 3675 1933 3676 1937
rect 3670 1932 3676 1933
rect 3630 1919 3636 1920
rect 3630 1915 3631 1919
rect 3635 1915 3636 1919
rect 3630 1914 3636 1915
rect 3672 1907 3674 1932
rect 3712 1920 3714 2026
rect 3726 2020 3732 2021
rect 3726 2016 3727 2020
rect 3731 2016 3732 2020
rect 3726 2015 3732 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3838 2015 3844 2016
rect 3728 1987 3730 2015
rect 3840 1987 3842 2015
rect 3727 1986 3731 1987
rect 3727 1981 3731 1982
rect 3799 1986 3803 1987
rect 3799 1981 3803 1982
rect 3839 1986 3843 1987
rect 3839 1981 3843 1982
rect 3800 1957 3802 1981
rect 3798 1956 3804 1957
rect 3798 1952 3799 1956
rect 3803 1952 3804 1956
rect 3798 1951 3804 1952
rect 3868 1948 3870 2226
rect 3906 2111 3912 2112
rect 3906 2107 3907 2111
rect 3911 2107 3912 2111
rect 3906 2106 3912 2107
rect 3908 2060 3910 2106
rect 3916 2084 3918 2278
rect 3942 2272 3948 2273
rect 3942 2268 3943 2272
rect 3947 2268 3948 2272
rect 3942 2267 3948 2268
rect 3944 2239 3946 2267
rect 3943 2238 3947 2239
rect 3943 2233 3947 2234
rect 3944 2213 3946 2233
rect 3942 2212 3948 2213
rect 3942 2208 3943 2212
rect 3947 2208 3948 2212
rect 3942 2207 3948 2208
rect 3942 2195 3948 2196
rect 3942 2191 3943 2195
rect 3947 2191 3948 2195
rect 3942 2190 3948 2191
rect 3944 2151 3946 2190
rect 3943 2150 3947 2151
rect 3943 2145 3947 2146
rect 3944 2118 3946 2145
rect 3942 2117 3948 2118
rect 3942 2113 3943 2117
rect 3947 2113 3948 2117
rect 3942 2112 3948 2113
rect 3942 2100 3948 2101
rect 3942 2096 3943 2100
rect 3947 2096 3948 2100
rect 3942 2095 3948 2096
rect 3914 2083 3920 2084
rect 3914 2079 3915 2083
rect 3919 2079 3920 2083
rect 3914 2078 3920 2079
rect 3944 2067 3946 2095
rect 3943 2066 3947 2067
rect 3943 2061 3947 2062
rect 3906 2059 3912 2060
rect 3906 2055 3907 2059
rect 3911 2055 3912 2059
rect 3906 2054 3912 2055
rect 3944 2041 3946 2061
rect 3942 2040 3948 2041
rect 3942 2036 3943 2040
rect 3947 2036 3948 2040
rect 3942 2035 3948 2036
rect 3914 2027 3920 2028
rect 3914 2023 3915 2027
rect 3919 2023 3920 2027
rect 3914 2022 3920 2023
rect 3942 2023 3948 2024
rect 3866 1947 3872 1948
rect 3866 1943 3867 1947
rect 3871 1943 3872 1947
rect 3866 1942 3872 1943
rect 3798 1937 3804 1938
rect 3798 1933 3799 1937
rect 3803 1933 3804 1937
rect 3798 1932 3804 1933
rect 3710 1919 3716 1920
rect 3710 1915 3711 1919
rect 3715 1915 3716 1919
rect 3710 1914 3716 1915
rect 3800 1907 3802 1932
rect 3858 1915 3864 1916
rect 3858 1911 3859 1915
rect 3863 1911 3864 1915
rect 3858 1910 3864 1911
rect 2927 1906 2931 1907
rect 2927 1901 2931 1902
rect 2959 1906 2963 1907
rect 2959 1901 2963 1902
rect 3047 1906 3051 1907
rect 3047 1901 3051 1902
rect 3127 1906 3131 1907
rect 3127 1901 3131 1902
rect 3175 1906 3179 1907
rect 3258 1903 3259 1907
rect 3263 1903 3264 1907
rect 3258 1902 3264 1903
rect 3295 1906 3299 1907
rect 3175 1901 3179 1902
rect 3295 1901 3299 1902
rect 3303 1906 3307 1907
rect 3303 1901 3307 1902
rect 3415 1906 3419 1907
rect 3415 1901 3419 1902
rect 3487 1906 3491 1907
rect 3487 1901 3491 1902
rect 3543 1906 3547 1907
rect 3543 1901 3547 1902
rect 3671 1906 3675 1907
rect 3671 1901 3675 1902
rect 3799 1906 3803 1907
rect 3799 1901 3803 1902
rect 3839 1906 3843 1907
rect 3839 1901 3843 1902
rect 2960 1880 2962 1901
rect 3034 1899 3040 1900
rect 3034 1895 3035 1899
rect 3039 1895 3040 1899
rect 3034 1894 3040 1895
rect 2958 1879 2964 1880
rect 2958 1875 2959 1879
rect 2963 1875 2964 1879
rect 2958 1874 2964 1875
rect 3036 1872 3038 1894
rect 3128 1880 3130 1901
rect 3202 1899 3208 1900
rect 3202 1895 3203 1899
rect 3207 1895 3208 1899
rect 3202 1894 3208 1895
rect 3126 1879 3132 1880
rect 3126 1875 3127 1879
rect 3131 1875 3132 1879
rect 3126 1874 3132 1875
rect 3204 1872 3206 1894
rect 3304 1880 3306 1901
rect 3378 1899 3384 1900
rect 3378 1895 3379 1899
rect 3383 1895 3384 1899
rect 3378 1894 3384 1895
rect 3302 1879 3308 1880
rect 3302 1875 3303 1879
rect 3307 1875 3308 1879
rect 3302 1874 3308 1875
rect 3380 1872 3382 1894
rect 3488 1880 3490 1901
rect 3562 1899 3568 1900
rect 3562 1895 3563 1899
rect 3567 1895 3568 1899
rect 3562 1894 3568 1895
rect 3486 1879 3492 1880
rect 3486 1875 3487 1879
rect 3491 1875 3492 1879
rect 3486 1874 3492 1875
rect 3564 1872 3566 1894
rect 3672 1880 3674 1901
rect 3840 1880 3842 1901
rect 3670 1879 3676 1880
rect 3670 1875 3671 1879
rect 3675 1875 3676 1879
rect 3670 1874 3676 1875
rect 3838 1879 3844 1880
rect 3838 1875 3839 1879
rect 3843 1875 3844 1879
rect 3838 1874 3844 1875
rect 2514 1871 2520 1872
rect 2514 1867 2515 1871
rect 2519 1867 2520 1871
rect 2514 1866 2520 1867
rect 2866 1871 2872 1872
rect 2866 1867 2867 1871
rect 2871 1867 2872 1871
rect 2866 1866 2872 1867
rect 3034 1871 3040 1872
rect 3034 1867 3035 1871
rect 3039 1867 3040 1871
rect 3034 1866 3040 1867
rect 3202 1871 3208 1872
rect 3202 1867 3203 1871
rect 3207 1867 3208 1871
rect 3202 1866 3208 1867
rect 3378 1871 3384 1872
rect 3378 1867 3379 1871
rect 3383 1867 3384 1871
rect 3378 1866 3384 1867
rect 3562 1871 3568 1872
rect 3562 1867 3563 1871
rect 3567 1867 3568 1871
rect 3562 1866 3568 1867
rect 3606 1871 3612 1872
rect 3606 1867 3607 1871
rect 3611 1867 3612 1871
rect 3606 1866 3612 1867
rect 2622 1860 2628 1861
rect 2622 1856 2623 1860
rect 2627 1856 2628 1860
rect 2622 1855 2628 1856
rect 2790 1860 2796 1861
rect 2790 1856 2791 1860
rect 2795 1856 2796 1860
rect 2790 1855 2796 1856
rect 2958 1860 2964 1861
rect 2958 1856 2959 1860
rect 2963 1856 2964 1860
rect 2958 1855 2964 1856
rect 3126 1860 3132 1861
rect 3126 1856 3127 1860
rect 3131 1856 3132 1860
rect 3126 1855 3132 1856
rect 3302 1860 3308 1861
rect 3302 1856 3303 1860
rect 3307 1856 3308 1860
rect 3302 1855 3308 1856
rect 3486 1860 3492 1861
rect 3486 1856 3487 1860
rect 3491 1856 3492 1860
rect 3486 1855 3492 1856
rect 2624 1831 2626 1855
rect 2792 1831 2794 1855
rect 2960 1831 2962 1855
rect 3128 1831 3130 1855
rect 3304 1831 3306 1855
rect 3488 1831 3490 1855
rect 2511 1830 2515 1831
rect 2511 1825 2515 1826
rect 2623 1830 2627 1831
rect 2623 1825 2627 1826
rect 2671 1830 2675 1831
rect 2671 1825 2675 1826
rect 2791 1830 2795 1831
rect 2791 1825 2795 1826
rect 2855 1830 2859 1831
rect 2855 1825 2859 1826
rect 2959 1830 2963 1831
rect 2959 1825 2963 1826
rect 3071 1830 3075 1831
rect 3071 1825 3075 1826
rect 3127 1830 3131 1831
rect 3127 1825 3131 1826
rect 3303 1830 3307 1831
rect 3303 1825 3307 1826
rect 3487 1830 3491 1831
rect 3487 1825 3491 1826
rect 3543 1830 3547 1831
rect 3543 1825 3547 1826
rect 2512 1801 2514 1825
rect 2672 1801 2674 1825
rect 2856 1801 2858 1825
rect 3072 1801 3074 1825
rect 3304 1801 3306 1825
rect 3544 1801 3546 1825
rect 2510 1800 2516 1801
rect 2510 1796 2511 1800
rect 2515 1796 2516 1800
rect 2510 1795 2516 1796
rect 2670 1800 2676 1801
rect 2670 1796 2671 1800
rect 2675 1796 2676 1800
rect 2670 1795 2676 1796
rect 2854 1800 2860 1801
rect 2854 1796 2855 1800
rect 2859 1796 2860 1800
rect 2854 1795 2860 1796
rect 3070 1800 3076 1801
rect 3070 1796 3071 1800
rect 3075 1796 3076 1800
rect 3070 1795 3076 1796
rect 3302 1800 3308 1801
rect 3302 1796 3303 1800
rect 3307 1796 3308 1800
rect 3302 1795 3308 1796
rect 3542 1800 3548 1801
rect 3542 1796 3543 1800
rect 3547 1796 3548 1800
rect 3542 1795 3548 1796
rect 2170 1791 2176 1792
rect 2170 1787 2171 1791
rect 2175 1787 2176 1791
rect 2170 1786 2176 1787
rect 2306 1791 2312 1792
rect 2306 1787 2307 1791
rect 2311 1787 2312 1791
rect 2306 1786 2312 1787
rect 2434 1791 2440 1792
rect 2434 1787 2435 1791
rect 2439 1787 2440 1791
rect 2434 1786 2440 1787
rect 2478 1791 2484 1792
rect 2478 1787 2479 1791
rect 2483 1787 2484 1791
rect 2478 1786 2484 1787
rect 2770 1791 2776 1792
rect 2770 1787 2771 1791
rect 2775 1787 2776 1791
rect 2770 1786 2776 1787
rect 2938 1791 2944 1792
rect 2938 1787 2939 1791
rect 2943 1787 2944 1791
rect 2938 1786 2944 1787
rect 3166 1791 3172 1792
rect 3166 1787 3167 1791
rect 3171 1787 3172 1791
rect 3166 1786 3172 1787
rect 3422 1791 3428 1792
rect 3422 1787 3423 1791
rect 3427 1787 3428 1791
rect 3422 1786 3428 1787
rect 2172 1764 2174 1786
rect 2230 1781 2236 1782
rect 2230 1777 2231 1781
rect 2235 1777 2236 1781
rect 2230 1776 2236 1777
rect 2146 1763 2152 1764
rect 2146 1759 2147 1763
rect 2151 1759 2152 1763
rect 2146 1758 2152 1759
rect 2170 1763 2176 1764
rect 2170 1759 2171 1763
rect 2175 1759 2176 1763
rect 2170 1758 2176 1759
rect 2232 1755 2234 1776
rect 2308 1764 2310 1786
rect 2366 1781 2372 1782
rect 2366 1777 2367 1781
rect 2371 1777 2372 1781
rect 2366 1776 2372 1777
rect 2306 1763 2312 1764
rect 2306 1759 2307 1763
rect 2311 1759 2312 1763
rect 2306 1758 2312 1759
rect 2368 1755 2370 1776
rect 2047 1754 2051 1755
rect 1599 1750 1603 1751
rect 1599 1745 1603 1746
rect 1663 1750 1667 1751
rect 1663 1745 1667 1746
rect 1847 1750 1851 1751
rect 1847 1745 1851 1746
rect 2007 1750 2011 1751
rect 2047 1749 2051 1750
rect 2095 1754 2099 1755
rect 2095 1749 2099 1750
rect 2183 1754 2187 1755
rect 2183 1749 2187 1750
rect 2231 1754 2235 1755
rect 2231 1749 2235 1750
rect 2287 1754 2291 1755
rect 2287 1749 2291 1750
rect 2367 1754 2371 1755
rect 2367 1749 2371 1750
rect 2391 1754 2395 1755
rect 2436 1753 2438 1786
rect 2510 1781 2516 1782
rect 2510 1777 2511 1781
rect 2515 1777 2516 1781
rect 2510 1776 2516 1777
rect 2670 1781 2676 1782
rect 2670 1777 2671 1781
rect 2675 1777 2676 1781
rect 2670 1776 2676 1777
rect 2512 1755 2514 1776
rect 2672 1755 2674 1776
rect 2682 1759 2688 1760
rect 2682 1755 2683 1759
rect 2687 1755 2688 1759
rect 2428 1752 2438 1753
rect 2391 1749 2395 1750
rect 2426 1751 2438 1752
rect 2495 1754 2499 1755
rect 2007 1745 2011 1746
rect 1562 1743 1568 1744
rect 1562 1739 1563 1743
rect 1567 1739 1568 1743
rect 1562 1738 1568 1739
rect 1600 1724 1602 1745
rect 2008 1725 2010 1745
rect 2048 1729 2050 1749
rect 2046 1728 2052 1729
rect 2184 1728 2186 1749
rect 2266 1747 2272 1748
rect 2266 1743 2267 1747
rect 2271 1743 2272 1747
rect 2266 1742 2272 1743
rect 2006 1724 2012 1725
rect 1438 1723 1444 1724
rect 1438 1719 1439 1723
rect 1443 1719 1444 1723
rect 1438 1718 1444 1719
rect 1598 1723 1604 1724
rect 1598 1719 1599 1723
rect 1603 1719 1604 1723
rect 2006 1720 2007 1724
rect 2011 1720 2012 1724
rect 2046 1724 2047 1728
rect 2051 1724 2052 1728
rect 2046 1723 2052 1724
rect 2182 1727 2188 1728
rect 2182 1723 2183 1727
rect 2187 1723 2188 1727
rect 2182 1722 2188 1723
rect 2268 1720 2270 1742
rect 2288 1728 2290 1749
rect 2374 1747 2380 1748
rect 2374 1743 2375 1747
rect 2379 1743 2380 1747
rect 2374 1742 2380 1743
rect 2286 1727 2292 1728
rect 2286 1723 2287 1727
rect 2291 1723 2292 1727
rect 2286 1722 2292 1723
rect 2376 1720 2378 1742
rect 2392 1728 2394 1749
rect 2426 1747 2427 1751
rect 2431 1747 2432 1751
rect 2495 1749 2499 1750
rect 2511 1754 2515 1755
rect 2511 1749 2515 1750
rect 2599 1754 2603 1755
rect 2599 1749 2603 1750
rect 2671 1754 2675 1755
rect 2682 1754 2688 1755
rect 2703 1754 2707 1755
rect 2671 1749 2675 1750
rect 2426 1746 2432 1747
rect 2496 1728 2498 1749
rect 2570 1747 2576 1748
rect 2570 1743 2571 1747
rect 2575 1743 2576 1747
rect 2570 1742 2576 1743
rect 2390 1727 2396 1728
rect 2390 1723 2391 1727
rect 2395 1723 2396 1727
rect 2390 1722 2396 1723
rect 2494 1727 2500 1728
rect 2494 1723 2495 1727
rect 2499 1723 2500 1727
rect 2494 1722 2500 1723
rect 2572 1720 2574 1742
rect 2600 1728 2602 1749
rect 2626 1739 2632 1740
rect 2626 1735 2627 1739
rect 2631 1735 2632 1739
rect 2626 1734 2632 1735
rect 2598 1727 2604 1728
rect 2598 1723 2599 1727
rect 2603 1723 2604 1727
rect 2598 1722 2604 1723
rect 2006 1719 2012 1720
rect 2266 1719 2272 1720
rect 1598 1718 1604 1719
rect 1202 1715 1208 1716
rect 1202 1711 1203 1715
rect 1207 1711 1208 1715
rect 1202 1710 1208 1711
rect 1354 1715 1360 1716
rect 1354 1711 1355 1715
rect 1359 1711 1360 1715
rect 1354 1710 1360 1711
rect 1362 1715 1368 1716
rect 1362 1711 1363 1715
rect 1367 1711 1368 1715
rect 1362 1710 1368 1711
rect 1582 1715 1588 1716
rect 1582 1711 1583 1715
rect 1587 1711 1588 1715
rect 2258 1715 2264 1716
rect 1582 1710 1588 1711
rect 2046 1711 2052 1712
rect 1278 1704 1284 1705
rect 1278 1700 1279 1704
rect 1283 1700 1284 1704
rect 1278 1699 1284 1700
rect 1438 1704 1444 1705
rect 1438 1700 1439 1704
rect 1443 1700 1444 1704
rect 1438 1699 1444 1700
rect 1280 1671 1282 1699
rect 1440 1671 1442 1699
rect 1167 1670 1171 1671
rect 1167 1665 1171 1666
rect 1279 1670 1283 1671
rect 1279 1665 1283 1666
rect 1351 1670 1355 1671
rect 1351 1665 1355 1666
rect 1439 1670 1443 1671
rect 1439 1665 1443 1666
rect 1543 1670 1547 1671
rect 1543 1665 1547 1666
rect 1168 1641 1170 1665
rect 1352 1641 1354 1665
rect 1544 1641 1546 1665
rect 1166 1640 1172 1641
rect 1166 1636 1167 1640
rect 1171 1636 1172 1640
rect 1166 1635 1172 1636
rect 1350 1640 1356 1641
rect 1350 1636 1351 1640
rect 1355 1636 1356 1640
rect 1350 1635 1356 1636
rect 1542 1640 1548 1641
rect 1542 1636 1543 1640
rect 1547 1636 1548 1640
rect 1542 1635 1548 1636
rect 1158 1631 1164 1632
rect 1158 1627 1159 1631
rect 1163 1627 1164 1631
rect 1158 1626 1164 1627
rect 1166 1621 1172 1622
rect 1166 1617 1167 1621
rect 1171 1617 1172 1621
rect 1166 1616 1172 1617
rect 1350 1621 1356 1622
rect 1350 1617 1351 1621
rect 1355 1617 1356 1621
rect 1350 1616 1356 1617
rect 1542 1621 1548 1622
rect 1542 1617 1543 1621
rect 1547 1617 1548 1621
rect 1542 1616 1548 1617
rect 1058 1603 1064 1604
rect 1058 1599 1059 1603
rect 1063 1599 1064 1603
rect 1058 1598 1064 1599
rect 1168 1595 1170 1616
rect 1352 1595 1354 1616
rect 1442 1599 1448 1600
rect 1442 1595 1443 1599
rect 1447 1595 1448 1599
rect 1544 1595 1546 1616
rect 1584 1604 1586 1710
rect 2006 1707 2012 1708
rect 1598 1704 1604 1705
rect 1598 1700 1599 1704
rect 1603 1700 1604 1704
rect 2006 1703 2007 1707
rect 2011 1703 2012 1707
rect 2046 1707 2047 1711
rect 2051 1707 2052 1711
rect 2258 1711 2259 1715
rect 2263 1711 2264 1715
rect 2266 1715 2267 1719
rect 2271 1715 2272 1719
rect 2266 1714 2272 1715
rect 2374 1719 2380 1720
rect 2374 1715 2375 1719
rect 2379 1715 2380 1719
rect 2374 1714 2380 1715
rect 2570 1719 2576 1720
rect 2570 1715 2571 1719
rect 2575 1715 2576 1719
rect 2570 1714 2576 1715
rect 2258 1710 2264 1711
rect 2046 1706 2052 1707
rect 2182 1708 2188 1709
rect 2006 1702 2012 1703
rect 1598 1699 1604 1700
rect 1600 1671 1602 1699
rect 2008 1671 2010 1702
rect 2048 1679 2050 1706
rect 2182 1704 2183 1708
rect 2187 1704 2188 1708
rect 2182 1703 2188 1704
rect 2184 1679 2186 1703
rect 2047 1678 2051 1679
rect 2047 1673 2051 1674
rect 2183 1678 2187 1679
rect 2183 1673 2187 1674
rect 2231 1678 2235 1679
rect 2231 1673 2235 1674
rect 1599 1670 1603 1671
rect 1599 1665 1603 1666
rect 1735 1670 1739 1671
rect 1735 1665 1739 1666
rect 2007 1670 2011 1671
rect 2007 1665 2011 1666
rect 1736 1641 1738 1665
rect 1734 1640 1740 1641
rect 1734 1636 1735 1640
rect 1739 1636 1740 1640
rect 2008 1638 2010 1665
rect 2048 1646 2050 1673
rect 2232 1649 2234 1673
rect 2230 1648 2236 1649
rect 2046 1645 2052 1646
rect 2046 1641 2047 1645
rect 2051 1641 2052 1645
rect 2230 1644 2231 1648
rect 2235 1644 2236 1648
rect 2230 1643 2236 1644
rect 2046 1640 2052 1641
rect 1734 1635 1740 1636
rect 2006 1637 2012 1638
rect 2006 1633 2007 1637
rect 2011 1633 2012 1637
rect 2006 1632 2012 1633
rect 1618 1631 1624 1632
rect 1618 1627 1619 1631
rect 1623 1627 1624 1631
rect 1618 1626 1624 1627
rect 1802 1631 1808 1632
rect 1802 1627 1803 1631
rect 1807 1627 1808 1631
rect 2230 1629 2236 1630
rect 1802 1626 1808 1627
rect 2046 1628 2052 1629
rect 1620 1604 1622 1626
rect 1734 1621 1740 1622
rect 1734 1617 1735 1621
rect 1739 1617 1740 1621
rect 1734 1616 1740 1617
rect 1582 1603 1588 1604
rect 1582 1599 1583 1603
rect 1587 1599 1588 1603
rect 1582 1598 1588 1599
rect 1618 1603 1624 1604
rect 1618 1599 1619 1603
rect 1623 1599 1624 1603
rect 1618 1598 1624 1599
rect 1736 1595 1738 1616
rect 1167 1594 1171 1595
rect 1167 1589 1171 1590
rect 1183 1594 1187 1595
rect 1183 1589 1187 1590
rect 1351 1594 1355 1595
rect 1351 1589 1355 1590
rect 1367 1594 1371 1595
rect 1442 1594 1448 1595
rect 1543 1594 1547 1595
rect 1367 1589 1371 1590
rect 1050 1587 1056 1588
rect 1050 1583 1051 1587
rect 1055 1583 1056 1587
rect 1050 1582 1056 1583
rect 1184 1568 1186 1589
rect 1250 1587 1256 1588
rect 1250 1583 1251 1587
rect 1255 1583 1256 1587
rect 1250 1582 1256 1583
rect 1258 1587 1264 1588
rect 1258 1583 1259 1587
rect 1263 1583 1264 1587
rect 1258 1582 1264 1583
rect 798 1567 804 1568
rect 798 1563 799 1567
rect 803 1563 804 1567
rect 798 1562 804 1563
rect 990 1567 996 1568
rect 990 1563 991 1567
rect 995 1563 996 1567
rect 990 1562 996 1563
rect 1182 1567 1188 1568
rect 1182 1563 1183 1567
rect 1187 1563 1188 1567
rect 1182 1562 1188 1563
rect 210 1559 216 1560
rect 210 1555 211 1559
rect 215 1555 216 1559
rect 210 1554 216 1555
rect 330 1559 336 1560
rect 330 1555 331 1559
rect 335 1555 336 1559
rect 330 1554 336 1555
rect 498 1559 504 1560
rect 498 1555 499 1559
rect 503 1555 504 1559
rect 498 1554 504 1555
rect 682 1559 688 1560
rect 682 1555 683 1559
rect 687 1555 688 1559
rect 682 1554 688 1555
rect 738 1559 744 1560
rect 738 1555 739 1559
rect 743 1555 744 1559
rect 738 1554 744 1555
rect 1066 1555 1072 1556
rect 1066 1551 1067 1555
rect 1071 1551 1072 1555
rect 1066 1550 1072 1551
rect 254 1548 260 1549
rect 254 1544 255 1548
rect 259 1544 260 1548
rect 254 1543 260 1544
rect 422 1548 428 1549
rect 422 1544 423 1548
rect 427 1544 428 1548
rect 422 1543 428 1544
rect 606 1548 612 1549
rect 606 1544 607 1548
rect 611 1544 612 1548
rect 606 1543 612 1544
rect 798 1548 804 1549
rect 798 1544 799 1548
rect 803 1544 804 1548
rect 798 1543 804 1544
rect 990 1548 996 1549
rect 990 1544 991 1548
rect 995 1544 996 1548
rect 990 1543 996 1544
rect 256 1515 258 1543
rect 424 1515 426 1543
rect 608 1515 610 1543
rect 800 1515 802 1543
rect 992 1515 994 1543
rect 247 1514 251 1515
rect 247 1509 251 1510
rect 255 1514 259 1515
rect 255 1509 259 1510
rect 399 1514 403 1515
rect 399 1509 403 1510
rect 423 1514 427 1515
rect 423 1509 427 1510
rect 559 1514 563 1515
rect 559 1509 563 1510
rect 607 1514 611 1515
rect 607 1509 611 1510
rect 719 1514 723 1515
rect 719 1509 723 1510
rect 799 1514 803 1515
rect 799 1509 803 1510
rect 879 1514 883 1515
rect 879 1509 883 1510
rect 991 1514 995 1515
rect 991 1509 995 1510
rect 1039 1514 1043 1515
rect 1039 1509 1043 1510
rect 202 1491 208 1492
rect 202 1487 203 1491
rect 207 1487 208 1491
rect 202 1486 208 1487
rect 248 1485 250 1509
rect 400 1485 402 1509
rect 560 1485 562 1509
rect 720 1485 722 1509
rect 880 1485 882 1509
rect 1040 1485 1042 1509
rect 134 1484 140 1485
rect 110 1481 116 1482
rect 110 1477 111 1481
rect 115 1477 116 1481
rect 134 1480 135 1484
rect 139 1480 140 1484
rect 134 1479 140 1480
rect 246 1484 252 1485
rect 246 1480 247 1484
rect 251 1480 252 1484
rect 246 1479 252 1480
rect 398 1484 404 1485
rect 398 1480 399 1484
rect 403 1480 404 1484
rect 398 1479 404 1480
rect 558 1484 564 1485
rect 558 1480 559 1484
rect 563 1480 564 1484
rect 558 1479 564 1480
rect 718 1484 724 1485
rect 718 1480 719 1484
rect 723 1480 724 1484
rect 718 1479 724 1480
rect 878 1484 884 1485
rect 878 1480 879 1484
rect 883 1480 884 1484
rect 878 1479 884 1480
rect 1038 1484 1044 1485
rect 1038 1480 1039 1484
rect 1043 1480 1044 1484
rect 1038 1479 1044 1480
rect 110 1476 116 1477
rect 210 1475 216 1476
rect 210 1471 211 1475
rect 215 1471 216 1475
rect 210 1470 216 1471
rect 322 1475 328 1476
rect 322 1471 323 1475
rect 327 1471 328 1475
rect 322 1470 328 1471
rect 474 1475 480 1476
rect 474 1471 475 1475
rect 479 1471 480 1475
rect 474 1470 480 1471
rect 634 1475 640 1476
rect 634 1471 635 1475
rect 639 1471 640 1475
rect 634 1470 640 1471
rect 954 1475 960 1476
rect 954 1471 955 1475
rect 959 1471 960 1475
rect 954 1470 960 1471
rect 134 1465 140 1466
rect 110 1464 116 1465
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 134 1461 135 1465
rect 139 1461 140 1465
rect 134 1460 140 1461
rect 110 1459 116 1460
rect 112 1439 114 1459
rect 136 1439 138 1460
rect 212 1448 214 1470
rect 246 1465 252 1466
rect 246 1461 247 1465
rect 251 1461 252 1465
rect 246 1460 252 1461
rect 210 1447 216 1448
rect 210 1443 211 1447
rect 215 1443 216 1447
rect 210 1442 216 1443
rect 210 1439 216 1440
rect 248 1439 250 1460
rect 324 1448 326 1470
rect 398 1465 404 1466
rect 398 1461 399 1465
rect 403 1461 404 1465
rect 398 1460 404 1461
rect 322 1447 328 1448
rect 322 1443 323 1447
rect 327 1443 328 1447
rect 322 1442 328 1443
rect 400 1439 402 1460
rect 476 1448 478 1470
rect 558 1465 564 1466
rect 558 1461 559 1465
rect 563 1461 564 1465
rect 558 1460 564 1461
rect 474 1447 480 1448
rect 474 1443 475 1447
rect 479 1443 480 1447
rect 474 1442 480 1443
rect 560 1439 562 1460
rect 636 1448 638 1470
rect 718 1465 724 1466
rect 718 1461 719 1465
rect 723 1461 724 1465
rect 718 1460 724 1461
rect 878 1465 884 1466
rect 878 1461 879 1465
rect 883 1461 884 1465
rect 878 1460 884 1461
rect 634 1447 640 1448
rect 634 1443 635 1447
rect 639 1443 640 1447
rect 634 1442 640 1443
rect 720 1439 722 1460
rect 880 1439 882 1460
rect 111 1438 115 1439
rect 111 1433 115 1434
rect 135 1438 139 1439
rect 210 1435 211 1439
rect 215 1435 216 1439
rect 210 1434 216 1435
rect 247 1438 251 1439
rect 135 1433 139 1434
rect 112 1413 114 1433
rect 110 1412 116 1413
rect 136 1412 138 1433
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 110 1407 116 1408
rect 134 1411 140 1412
rect 134 1407 135 1411
rect 139 1407 140 1411
rect 134 1406 140 1407
rect 212 1404 214 1434
rect 247 1433 251 1434
rect 263 1438 267 1439
rect 263 1433 267 1434
rect 399 1438 403 1439
rect 399 1433 403 1434
rect 431 1438 435 1439
rect 431 1433 435 1434
rect 559 1438 563 1439
rect 559 1433 563 1434
rect 607 1438 611 1439
rect 607 1433 611 1434
rect 719 1438 723 1439
rect 719 1433 723 1434
rect 791 1438 795 1439
rect 791 1433 795 1434
rect 879 1438 883 1439
rect 879 1433 883 1434
rect 218 1431 224 1432
rect 218 1427 219 1431
rect 223 1427 224 1431
rect 218 1426 224 1427
rect 220 1404 222 1426
rect 264 1412 266 1433
rect 366 1431 372 1432
rect 366 1427 367 1431
rect 371 1427 372 1431
rect 366 1426 372 1427
rect 262 1411 268 1412
rect 262 1407 263 1411
rect 267 1407 268 1411
rect 262 1406 268 1407
rect 368 1404 370 1426
rect 432 1412 434 1433
rect 578 1431 584 1432
rect 578 1427 579 1431
rect 583 1427 584 1431
rect 578 1426 584 1427
rect 430 1411 436 1412
rect 430 1407 431 1411
rect 435 1407 436 1411
rect 430 1406 436 1407
rect 210 1403 216 1404
rect 210 1399 211 1403
rect 215 1399 216 1403
rect 210 1398 216 1399
rect 218 1403 224 1404
rect 218 1399 219 1403
rect 223 1399 224 1403
rect 218 1398 224 1399
rect 366 1403 372 1404
rect 366 1399 367 1403
rect 371 1399 372 1403
rect 366 1398 372 1399
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 110 1390 116 1391
rect 134 1392 140 1393
rect 112 1359 114 1390
rect 134 1388 135 1392
rect 139 1388 140 1392
rect 134 1387 140 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 430 1392 436 1393
rect 430 1388 431 1392
rect 435 1388 436 1392
rect 430 1387 436 1388
rect 136 1359 138 1387
rect 264 1359 266 1387
rect 432 1359 434 1387
rect 111 1358 115 1359
rect 111 1353 115 1354
rect 135 1358 139 1359
rect 135 1353 139 1354
rect 159 1358 163 1359
rect 159 1353 163 1354
rect 263 1358 267 1359
rect 263 1353 267 1354
rect 311 1358 315 1359
rect 311 1353 315 1354
rect 431 1358 435 1359
rect 431 1353 435 1354
rect 479 1358 483 1359
rect 479 1353 483 1354
rect 112 1326 114 1353
rect 160 1329 162 1353
rect 312 1329 314 1353
rect 480 1329 482 1353
rect 158 1328 164 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 158 1324 159 1328
rect 163 1324 164 1328
rect 158 1323 164 1324
rect 310 1328 316 1329
rect 310 1324 311 1328
rect 315 1324 316 1328
rect 310 1323 316 1324
rect 478 1328 484 1329
rect 478 1324 479 1328
rect 483 1324 484 1328
rect 478 1323 484 1324
rect 110 1320 116 1321
rect 580 1320 582 1426
rect 608 1412 610 1433
rect 682 1431 688 1432
rect 682 1427 683 1431
rect 687 1427 688 1431
rect 682 1426 688 1427
rect 606 1411 612 1412
rect 606 1407 607 1411
rect 611 1407 612 1411
rect 606 1406 612 1407
rect 684 1404 686 1426
rect 690 1423 696 1424
rect 690 1419 691 1423
rect 695 1419 696 1423
rect 690 1418 696 1419
rect 692 1404 694 1418
rect 792 1412 794 1433
rect 956 1432 958 1470
rect 1038 1465 1044 1466
rect 1038 1461 1039 1465
rect 1043 1461 1044 1465
rect 1038 1460 1044 1461
rect 1040 1439 1042 1460
rect 1068 1448 1070 1550
rect 1182 1548 1188 1549
rect 1182 1544 1183 1548
rect 1187 1544 1188 1548
rect 1182 1543 1188 1544
rect 1184 1515 1186 1543
rect 1183 1514 1187 1515
rect 1183 1509 1187 1510
rect 1184 1485 1186 1509
rect 1182 1484 1188 1485
rect 1182 1480 1183 1484
rect 1187 1480 1188 1484
rect 1182 1479 1188 1480
rect 1252 1476 1254 1582
rect 1260 1560 1262 1582
rect 1368 1568 1370 1589
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 1444 1560 1446 1594
rect 1543 1589 1547 1590
rect 1551 1594 1555 1595
rect 1551 1589 1555 1590
rect 1735 1594 1739 1595
rect 1735 1589 1739 1590
rect 1552 1568 1554 1589
rect 1634 1587 1640 1588
rect 1634 1583 1635 1587
rect 1639 1583 1640 1587
rect 1634 1582 1640 1583
rect 1550 1567 1556 1568
rect 1550 1563 1551 1567
rect 1555 1563 1556 1567
rect 1550 1562 1556 1563
rect 1636 1560 1638 1582
rect 1736 1568 1738 1589
rect 1804 1588 1806 1626
rect 2046 1624 2047 1628
rect 2051 1624 2052 1628
rect 2230 1625 2231 1629
rect 2235 1625 2236 1629
rect 2230 1624 2236 1625
rect 2046 1623 2052 1624
rect 2006 1620 2012 1621
rect 2006 1616 2007 1620
rect 2011 1616 2012 1620
rect 2006 1615 2012 1616
rect 2008 1595 2010 1615
rect 2048 1595 2050 1623
rect 2232 1595 2234 1624
rect 2260 1612 2262 1710
rect 2286 1708 2292 1709
rect 2286 1704 2287 1708
rect 2291 1704 2292 1708
rect 2286 1703 2292 1704
rect 2390 1708 2396 1709
rect 2390 1704 2391 1708
rect 2395 1704 2396 1708
rect 2390 1703 2396 1704
rect 2494 1708 2500 1709
rect 2494 1704 2495 1708
rect 2499 1704 2500 1708
rect 2494 1703 2500 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2288 1679 2290 1703
rect 2392 1679 2394 1703
rect 2496 1679 2498 1703
rect 2600 1679 2602 1703
rect 2287 1678 2291 1679
rect 2287 1673 2291 1674
rect 2367 1678 2371 1679
rect 2367 1673 2371 1674
rect 2391 1678 2395 1679
rect 2391 1673 2395 1674
rect 2495 1678 2499 1679
rect 2495 1673 2499 1674
rect 2519 1678 2523 1679
rect 2519 1673 2523 1674
rect 2599 1678 2603 1679
rect 2599 1673 2603 1674
rect 2368 1649 2370 1673
rect 2520 1649 2522 1673
rect 2366 1648 2372 1649
rect 2366 1644 2367 1648
rect 2371 1644 2372 1648
rect 2366 1643 2372 1644
rect 2518 1648 2524 1649
rect 2518 1644 2519 1648
rect 2523 1644 2524 1648
rect 2518 1643 2524 1644
rect 2628 1640 2630 1734
rect 2684 1720 2686 1754
rect 2703 1749 2707 1750
rect 2704 1728 2706 1749
rect 2772 1748 2774 1786
rect 2854 1781 2860 1782
rect 2854 1777 2855 1781
rect 2859 1777 2860 1781
rect 2854 1776 2860 1777
rect 2856 1755 2858 1776
rect 2940 1764 2942 1786
rect 3070 1781 3076 1782
rect 3070 1777 3071 1781
rect 3075 1777 3076 1781
rect 3070 1776 3076 1777
rect 2938 1763 2944 1764
rect 2938 1759 2939 1763
rect 2943 1759 2944 1763
rect 2938 1758 2944 1759
rect 3072 1755 3074 1776
rect 3168 1764 3170 1786
rect 3302 1781 3308 1782
rect 3302 1777 3303 1781
rect 3307 1777 3308 1781
rect 3302 1776 3308 1777
rect 3166 1763 3172 1764
rect 3166 1759 3167 1763
rect 3171 1759 3172 1763
rect 3166 1758 3172 1759
rect 3304 1755 3306 1776
rect 3424 1764 3426 1786
rect 3542 1781 3548 1782
rect 3542 1777 3543 1781
rect 3547 1777 3548 1781
rect 3542 1776 3548 1777
rect 3422 1763 3428 1764
rect 3422 1759 3423 1763
rect 3427 1759 3428 1763
rect 3422 1758 3428 1759
rect 3544 1755 3546 1776
rect 3608 1764 3610 1866
rect 3670 1860 3676 1861
rect 3670 1856 3671 1860
rect 3675 1856 3676 1860
rect 3670 1855 3676 1856
rect 3838 1860 3844 1861
rect 3838 1856 3839 1860
rect 3843 1856 3844 1860
rect 3838 1855 3844 1856
rect 3672 1831 3674 1855
rect 3840 1831 3842 1855
rect 3671 1830 3675 1831
rect 3671 1825 3675 1826
rect 3791 1830 3795 1831
rect 3791 1825 3795 1826
rect 3839 1830 3843 1831
rect 3839 1825 3843 1826
rect 3792 1801 3794 1825
rect 3790 1800 3796 1801
rect 3790 1796 3791 1800
rect 3795 1796 3796 1800
rect 3790 1795 3796 1796
rect 3860 1792 3862 1910
rect 3916 1900 3918 2022
rect 3942 2019 3943 2023
rect 3947 2019 3948 2023
rect 3942 2018 3948 2019
rect 3944 1987 3946 2018
rect 3943 1986 3947 1987
rect 3943 1981 3947 1982
rect 3944 1954 3946 1981
rect 3942 1953 3948 1954
rect 3942 1949 3943 1953
rect 3947 1949 3948 1953
rect 3942 1948 3948 1949
rect 3942 1936 3948 1937
rect 3942 1932 3943 1936
rect 3947 1932 3948 1936
rect 3942 1931 3948 1932
rect 3944 1907 3946 1931
rect 3943 1906 3947 1907
rect 3943 1901 3947 1902
rect 3914 1899 3920 1900
rect 3914 1895 3915 1899
rect 3919 1895 3920 1899
rect 3914 1894 3920 1895
rect 3944 1881 3946 1901
rect 3942 1880 3948 1881
rect 3942 1876 3943 1880
rect 3947 1876 3948 1880
rect 3942 1875 3948 1876
rect 3914 1867 3920 1868
rect 3914 1863 3915 1867
rect 3919 1863 3920 1867
rect 3914 1862 3920 1863
rect 3942 1863 3948 1864
rect 3858 1791 3864 1792
rect 3858 1787 3859 1791
rect 3863 1787 3864 1791
rect 3858 1786 3864 1787
rect 3790 1781 3796 1782
rect 3790 1777 3791 1781
rect 3795 1777 3796 1781
rect 3790 1776 3796 1777
rect 3606 1763 3612 1764
rect 3606 1759 3607 1763
rect 3611 1759 3612 1763
rect 3606 1758 3612 1759
rect 3792 1755 3794 1776
rect 3798 1759 3804 1760
rect 3798 1755 3799 1759
rect 3803 1755 3804 1759
rect 2807 1754 2811 1755
rect 2807 1749 2811 1750
rect 2855 1754 2859 1755
rect 2855 1749 2859 1750
rect 2911 1754 2915 1755
rect 2911 1749 2915 1750
rect 3015 1754 3019 1755
rect 3015 1749 3019 1750
rect 3071 1754 3075 1755
rect 3071 1749 3075 1750
rect 3127 1754 3131 1755
rect 3127 1749 3131 1750
rect 3303 1754 3307 1755
rect 3303 1749 3307 1750
rect 3543 1754 3547 1755
rect 3543 1749 3547 1750
rect 3791 1754 3795 1755
rect 3798 1754 3804 1755
rect 3791 1749 3795 1750
rect 2770 1747 2776 1748
rect 2770 1743 2771 1747
rect 2775 1743 2776 1747
rect 2770 1742 2776 1743
rect 2778 1747 2784 1748
rect 2778 1743 2779 1747
rect 2783 1743 2784 1747
rect 2778 1742 2784 1743
rect 2702 1727 2708 1728
rect 2702 1723 2703 1727
rect 2707 1723 2708 1727
rect 2702 1722 2708 1723
rect 2780 1720 2782 1742
rect 2808 1728 2810 1749
rect 2882 1747 2888 1748
rect 2882 1743 2883 1747
rect 2887 1743 2888 1747
rect 2882 1742 2888 1743
rect 2806 1727 2812 1728
rect 2806 1723 2807 1727
rect 2811 1723 2812 1727
rect 2806 1722 2812 1723
rect 2884 1720 2886 1742
rect 2912 1728 2914 1749
rect 2986 1747 2992 1748
rect 2986 1743 2987 1747
rect 2991 1743 2992 1747
rect 2986 1742 2992 1743
rect 2910 1727 2916 1728
rect 2910 1723 2911 1727
rect 2915 1723 2916 1727
rect 2910 1722 2916 1723
rect 2988 1720 2990 1742
rect 3016 1728 3018 1749
rect 3090 1747 3096 1748
rect 3090 1743 3091 1747
rect 3095 1743 3096 1747
rect 3090 1742 3096 1743
rect 3014 1727 3020 1728
rect 3014 1723 3015 1727
rect 3019 1723 3020 1727
rect 3014 1722 3020 1723
rect 3092 1720 3094 1742
rect 3128 1728 3130 1749
rect 3126 1727 3132 1728
rect 3126 1723 3127 1727
rect 3131 1723 3132 1727
rect 3126 1722 3132 1723
rect 2682 1719 2688 1720
rect 2682 1715 2683 1719
rect 2687 1715 2688 1719
rect 2682 1714 2688 1715
rect 2778 1719 2784 1720
rect 2778 1715 2779 1719
rect 2783 1715 2784 1719
rect 2778 1714 2784 1715
rect 2882 1719 2888 1720
rect 2882 1715 2883 1719
rect 2887 1715 2888 1719
rect 2882 1714 2888 1715
rect 2986 1719 2992 1720
rect 2986 1715 2987 1719
rect 2991 1715 2992 1719
rect 2986 1714 2992 1715
rect 3090 1719 3096 1720
rect 3090 1715 3091 1719
rect 3095 1715 3096 1719
rect 3090 1714 3096 1715
rect 3202 1715 3208 1716
rect 3202 1711 3203 1715
rect 3207 1711 3208 1715
rect 3202 1710 3208 1711
rect 2702 1708 2708 1709
rect 2702 1704 2703 1708
rect 2707 1704 2708 1708
rect 2702 1703 2708 1704
rect 2806 1708 2812 1709
rect 2806 1704 2807 1708
rect 2811 1704 2812 1708
rect 2806 1703 2812 1704
rect 2910 1708 2916 1709
rect 2910 1704 2911 1708
rect 2915 1704 2916 1708
rect 2910 1703 2916 1704
rect 3014 1708 3020 1709
rect 3014 1704 3015 1708
rect 3019 1704 3020 1708
rect 3014 1703 3020 1704
rect 3126 1708 3132 1709
rect 3126 1704 3127 1708
rect 3131 1704 3132 1708
rect 3126 1703 3132 1704
rect 2704 1679 2706 1703
rect 2808 1679 2810 1703
rect 2912 1679 2914 1703
rect 3016 1679 3018 1703
rect 3128 1679 3130 1703
rect 2679 1678 2683 1679
rect 2679 1673 2683 1674
rect 2703 1678 2707 1679
rect 2703 1673 2707 1674
rect 2807 1678 2811 1679
rect 2807 1673 2811 1674
rect 2847 1678 2851 1679
rect 2847 1673 2851 1674
rect 2911 1678 2915 1679
rect 2911 1673 2915 1674
rect 3015 1678 3019 1679
rect 3015 1673 3019 1674
rect 3023 1678 3027 1679
rect 3023 1673 3027 1674
rect 3127 1678 3131 1679
rect 3127 1673 3131 1674
rect 3191 1678 3195 1679
rect 3191 1673 3195 1674
rect 2680 1649 2682 1673
rect 2848 1649 2850 1673
rect 3024 1649 3026 1673
rect 3192 1649 3194 1673
rect 2678 1648 2684 1649
rect 2678 1644 2679 1648
rect 2683 1644 2684 1648
rect 2678 1643 2684 1644
rect 2846 1648 2852 1649
rect 2846 1644 2847 1648
rect 2851 1644 2852 1648
rect 2846 1643 2852 1644
rect 3022 1648 3028 1649
rect 3022 1644 3023 1648
rect 3027 1644 3028 1648
rect 3022 1643 3028 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 2306 1639 2312 1640
rect 2306 1635 2307 1639
rect 2311 1635 2312 1639
rect 2306 1634 2312 1635
rect 2442 1639 2448 1640
rect 2442 1635 2443 1639
rect 2447 1635 2448 1639
rect 2442 1634 2448 1635
rect 2594 1639 2600 1640
rect 2594 1635 2595 1639
rect 2599 1635 2600 1639
rect 2594 1634 2600 1635
rect 2626 1639 2632 1640
rect 2626 1635 2627 1639
rect 2631 1635 2632 1639
rect 2626 1634 2632 1635
rect 2762 1639 2768 1640
rect 2762 1635 2763 1639
rect 2767 1635 2768 1639
rect 2762 1634 2768 1635
rect 3106 1639 3112 1640
rect 3106 1635 3107 1639
rect 3111 1635 3112 1639
rect 3106 1634 3112 1635
rect 2308 1612 2310 1634
rect 2366 1629 2372 1630
rect 2366 1625 2367 1629
rect 2371 1625 2372 1629
rect 2366 1624 2372 1625
rect 2258 1611 2264 1612
rect 2258 1607 2259 1611
rect 2263 1607 2264 1611
rect 2258 1606 2264 1607
rect 2306 1611 2312 1612
rect 2306 1607 2307 1611
rect 2311 1607 2312 1611
rect 2306 1606 2312 1607
rect 2368 1595 2370 1624
rect 2444 1612 2446 1634
rect 2518 1629 2524 1630
rect 2518 1625 2519 1629
rect 2523 1625 2524 1629
rect 2518 1624 2524 1625
rect 2442 1611 2448 1612
rect 2442 1607 2443 1611
rect 2447 1607 2448 1611
rect 2442 1606 2448 1607
rect 2520 1595 2522 1624
rect 1903 1594 1907 1595
rect 1903 1589 1907 1590
rect 2007 1594 2011 1595
rect 2007 1589 2011 1590
rect 2047 1594 2051 1595
rect 2047 1589 2051 1590
rect 2071 1594 2075 1595
rect 2071 1589 2075 1590
rect 2231 1594 2235 1595
rect 2231 1589 2235 1590
rect 2271 1594 2275 1595
rect 2271 1589 2275 1590
rect 2367 1594 2371 1595
rect 2367 1589 2371 1590
rect 2495 1594 2499 1595
rect 2495 1589 2499 1590
rect 2519 1594 2523 1595
rect 2519 1589 2523 1590
rect 1802 1587 1808 1588
rect 1802 1583 1803 1587
rect 1807 1583 1808 1587
rect 1802 1582 1808 1583
rect 1762 1579 1768 1580
rect 1762 1575 1763 1579
rect 1767 1575 1768 1579
rect 1762 1574 1768 1575
rect 1734 1567 1740 1568
rect 1734 1563 1735 1567
rect 1739 1563 1740 1567
rect 1734 1562 1740 1563
rect 1258 1559 1264 1560
rect 1258 1555 1259 1559
rect 1263 1555 1264 1559
rect 1258 1554 1264 1555
rect 1442 1559 1448 1560
rect 1442 1555 1443 1559
rect 1447 1555 1448 1559
rect 1442 1554 1448 1555
rect 1454 1559 1460 1560
rect 1454 1555 1455 1559
rect 1459 1555 1460 1559
rect 1454 1554 1460 1555
rect 1634 1559 1640 1560
rect 1634 1555 1635 1559
rect 1639 1555 1640 1559
rect 1634 1554 1640 1555
rect 1366 1548 1372 1549
rect 1366 1544 1367 1548
rect 1371 1544 1372 1548
rect 1366 1543 1372 1544
rect 1368 1515 1370 1543
rect 1319 1514 1323 1515
rect 1319 1509 1323 1510
rect 1367 1514 1371 1515
rect 1367 1509 1371 1510
rect 1447 1514 1451 1515
rect 1447 1509 1451 1510
rect 1320 1485 1322 1509
rect 1448 1485 1450 1509
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1446 1484 1452 1485
rect 1446 1480 1447 1484
rect 1451 1480 1452 1484
rect 1446 1479 1452 1480
rect 1250 1475 1256 1476
rect 1250 1471 1251 1475
rect 1255 1471 1256 1475
rect 1250 1470 1256 1471
rect 1394 1475 1400 1476
rect 1394 1471 1395 1475
rect 1399 1471 1400 1475
rect 1394 1470 1400 1471
rect 1182 1465 1188 1466
rect 1182 1461 1183 1465
rect 1187 1461 1188 1465
rect 1182 1460 1188 1461
rect 1318 1465 1324 1466
rect 1318 1461 1319 1465
rect 1323 1461 1324 1465
rect 1318 1460 1324 1461
rect 1066 1447 1072 1448
rect 1066 1443 1067 1447
rect 1071 1443 1072 1447
rect 1066 1442 1072 1443
rect 1184 1439 1186 1460
rect 1242 1443 1248 1444
rect 1242 1439 1243 1443
rect 1247 1439 1248 1443
rect 1320 1439 1322 1460
rect 1396 1448 1398 1470
rect 1446 1465 1452 1466
rect 1446 1461 1447 1465
rect 1451 1461 1452 1465
rect 1446 1460 1452 1461
rect 1394 1447 1400 1448
rect 1394 1443 1395 1447
rect 1399 1443 1400 1447
rect 1394 1442 1400 1443
rect 1448 1439 1450 1460
rect 1456 1456 1458 1554
rect 1550 1548 1556 1549
rect 1550 1544 1551 1548
rect 1555 1544 1556 1548
rect 1550 1543 1556 1544
rect 1734 1548 1740 1549
rect 1734 1544 1735 1548
rect 1739 1544 1740 1548
rect 1734 1543 1740 1544
rect 1552 1515 1554 1543
rect 1736 1515 1738 1543
rect 1551 1514 1555 1515
rect 1551 1509 1555 1510
rect 1567 1514 1571 1515
rect 1567 1509 1571 1510
rect 1687 1514 1691 1515
rect 1687 1509 1691 1510
rect 1735 1514 1739 1515
rect 1735 1509 1739 1510
rect 1568 1485 1570 1509
rect 1688 1485 1690 1509
rect 1566 1484 1572 1485
rect 1566 1480 1567 1484
rect 1571 1480 1572 1484
rect 1566 1479 1572 1480
rect 1686 1484 1692 1485
rect 1686 1480 1687 1484
rect 1691 1480 1692 1484
rect 1686 1479 1692 1480
rect 1764 1476 1766 1574
rect 1904 1568 1906 1589
rect 1978 1587 1984 1588
rect 1978 1583 1979 1587
rect 1983 1583 1984 1587
rect 1978 1582 1984 1583
rect 1902 1567 1908 1568
rect 1902 1563 1903 1567
rect 1907 1563 1908 1567
rect 1902 1562 1908 1563
rect 1980 1560 1982 1582
rect 2008 1569 2010 1589
rect 2048 1569 2050 1589
rect 2006 1568 2012 1569
rect 2006 1564 2007 1568
rect 2011 1564 2012 1568
rect 2006 1563 2012 1564
rect 2046 1568 2052 1569
rect 2072 1568 2074 1589
rect 2146 1587 2152 1588
rect 2146 1583 2147 1587
rect 2151 1583 2152 1587
rect 2146 1582 2152 1583
rect 2046 1564 2047 1568
rect 2051 1564 2052 1568
rect 2046 1563 2052 1564
rect 2070 1567 2076 1568
rect 2070 1563 2071 1567
rect 2075 1563 2076 1567
rect 2070 1562 2076 1563
rect 2148 1560 2150 1582
rect 2272 1568 2274 1589
rect 2346 1587 2352 1588
rect 2346 1583 2347 1587
rect 2351 1583 2352 1587
rect 2346 1582 2352 1583
rect 2270 1567 2276 1568
rect 2270 1563 2271 1567
rect 2275 1563 2276 1567
rect 2270 1562 2276 1563
rect 2348 1560 2350 1582
rect 2496 1568 2498 1589
rect 2596 1588 2598 1634
rect 2678 1629 2684 1630
rect 2678 1625 2679 1629
rect 2683 1625 2684 1629
rect 2678 1624 2684 1625
rect 2680 1595 2682 1624
rect 2764 1612 2766 1634
rect 2846 1629 2852 1630
rect 2846 1625 2847 1629
rect 2851 1625 2852 1629
rect 2846 1624 2852 1625
rect 3022 1629 3028 1630
rect 3022 1625 3023 1629
rect 3027 1625 3028 1629
rect 3022 1624 3028 1625
rect 2762 1611 2768 1612
rect 2762 1607 2763 1611
rect 2767 1607 2768 1611
rect 2762 1606 2768 1607
rect 2786 1607 2792 1608
rect 2786 1603 2787 1607
rect 2791 1603 2792 1607
rect 2786 1602 2792 1603
rect 2679 1594 2683 1595
rect 2679 1589 2683 1590
rect 2711 1594 2715 1595
rect 2711 1589 2715 1590
rect 2594 1587 2600 1588
rect 2594 1583 2595 1587
rect 2599 1583 2600 1587
rect 2594 1582 2600 1583
rect 2712 1568 2714 1589
rect 2494 1567 2500 1568
rect 2494 1563 2495 1567
rect 2499 1563 2500 1567
rect 2494 1562 2500 1563
rect 2710 1567 2716 1568
rect 2710 1563 2711 1567
rect 2715 1563 2716 1567
rect 2710 1562 2716 1563
rect 2788 1560 2790 1602
rect 2848 1595 2850 1624
rect 3024 1595 3026 1624
rect 2847 1594 2851 1595
rect 2847 1589 2851 1590
rect 2911 1594 2915 1595
rect 2911 1589 2915 1590
rect 3023 1594 3027 1595
rect 3023 1589 3027 1590
rect 3095 1594 3099 1595
rect 3095 1589 3099 1590
rect 2912 1568 2914 1589
rect 2994 1587 3000 1588
rect 2994 1583 2995 1587
rect 2999 1583 3000 1587
rect 2994 1582 3000 1583
rect 2910 1567 2916 1568
rect 2910 1563 2911 1567
rect 2915 1563 2916 1567
rect 2910 1562 2916 1563
rect 2996 1560 2998 1582
rect 3096 1568 3098 1589
rect 3108 1588 3110 1634
rect 3190 1629 3196 1630
rect 3190 1625 3191 1629
rect 3195 1625 3196 1629
rect 3190 1624 3196 1625
rect 3192 1595 3194 1624
rect 3204 1612 3206 1710
rect 3359 1678 3363 1679
rect 3359 1673 3363 1674
rect 3527 1678 3531 1679
rect 3527 1673 3531 1674
rect 3695 1678 3699 1679
rect 3695 1673 3699 1674
rect 3360 1649 3362 1673
rect 3528 1649 3530 1673
rect 3696 1649 3698 1673
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3526 1648 3532 1649
rect 3526 1644 3527 1648
rect 3531 1644 3532 1648
rect 3526 1643 3532 1644
rect 3694 1648 3700 1649
rect 3694 1644 3695 1648
rect 3699 1644 3700 1648
rect 3694 1643 3700 1644
rect 3434 1639 3440 1640
rect 3434 1635 3435 1639
rect 3439 1635 3440 1639
rect 3434 1634 3440 1635
rect 3602 1639 3608 1640
rect 3602 1635 3603 1639
rect 3607 1635 3608 1639
rect 3602 1634 3608 1635
rect 3358 1629 3364 1630
rect 3358 1625 3359 1629
rect 3363 1625 3364 1629
rect 3358 1624 3364 1625
rect 3202 1611 3208 1612
rect 3202 1607 3203 1611
rect 3207 1607 3208 1611
rect 3202 1606 3208 1607
rect 3360 1595 3362 1624
rect 3436 1612 3438 1634
rect 3526 1629 3532 1630
rect 3526 1625 3527 1629
rect 3531 1625 3532 1629
rect 3526 1624 3532 1625
rect 3434 1611 3440 1612
rect 3398 1607 3404 1608
rect 3398 1603 3399 1607
rect 3403 1603 3404 1607
rect 3434 1607 3435 1611
rect 3439 1607 3440 1611
rect 3434 1606 3440 1607
rect 3398 1602 3404 1603
rect 3191 1594 3195 1595
rect 3191 1589 3195 1590
rect 3263 1594 3267 1595
rect 3263 1589 3267 1590
rect 3359 1594 3363 1595
rect 3359 1589 3363 1590
rect 3106 1587 3112 1588
rect 3106 1583 3107 1587
rect 3111 1583 3112 1587
rect 3106 1582 3112 1583
rect 3202 1587 3208 1588
rect 3202 1583 3203 1587
rect 3207 1583 3208 1587
rect 3202 1582 3208 1583
rect 3094 1567 3100 1568
rect 3094 1563 3095 1567
rect 3099 1563 3100 1567
rect 3094 1562 3100 1563
rect 1978 1559 1984 1560
rect 1978 1555 1979 1559
rect 1983 1555 1984 1559
rect 1978 1554 1984 1555
rect 2146 1559 2152 1560
rect 2146 1555 2147 1559
rect 2151 1555 2152 1559
rect 2146 1554 2152 1555
rect 2346 1559 2352 1560
rect 2346 1555 2347 1559
rect 2351 1555 2352 1559
rect 2346 1554 2352 1555
rect 2418 1559 2424 1560
rect 2418 1555 2419 1559
rect 2423 1555 2424 1559
rect 2418 1554 2424 1555
rect 2786 1559 2792 1560
rect 2786 1555 2787 1559
rect 2791 1555 2792 1559
rect 2786 1554 2792 1555
rect 2994 1559 3000 1560
rect 2994 1555 2995 1559
rect 2999 1555 3000 1559
rect 2994 1554 3000 1555
rect 2006 1551 2012 1552
rect 1902 1548 1908 1549
rect 1902 1544 1903 1548
rect 1907 1544 1908 1548
rect 2006 1547 2007 1551
rect 2011 1547 2012 1551
rect 2006 1546 2012 1547
rect 2046 1551 2052 1552
rect 2046 1547 2047 1551
rect 2051 1547 2052 1551
rect 2046 1546 2052 1547
rect 2070 1548 2076 1549
rect 1902 1543 1908 1544
rect 1904 1515 1906 1543
rect 2008 1515 2010 1546
rect 2048 1519 2050 1546
rect 2070 1544 2071 1548
rect 2075 1544 2076 1548
rect 2070 1543 2076 1544
rect 2270 1548 2276 1549
rect 2270 1544 2271 1548
rect 2275 1544 2276 1548
rect 2270 1543 2276 1544
rect 2072 1519 2074 1543
rect 2272 1519 2274 1543
rect 2047 1518 2051 1519
rect 1807 1514 1811 1515
rect 1807 1509 1811 1510
rect 1903 1514 1907 1515
rect 1903 1509 1907 1510
rect 2007 1514 2011 1515
rect 2047 1513 2051 1514
rect 2071 1518 2075 1519
rect 2071 1513 2075 1514
rect 2271 1518 2275 1519
rect 2271 1513 2275 1514
rect 2007 1509 2011 1510
rect 1808 1485 1810 1509
rect 1904 1485 1906 1509
rect 1806 1484 1812 1485
rect 1806 1480 1807 1484
rect 1811 1480 1812 1484
rect 1806 1479 1812 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 2008 1482 2010 1509
rect 2048 1486 2050 1513
rect 2072 1489 2074 1513
rect 2070 1488 2076 1489
rect 2046 1485 2052 1486
rect 1902 1479 1908 1480
rect 2006 1481 2012 1482
rect 2006 1477 2007 1481
rect 2011 1477 2012 1481
rect 2046 1481 2047 1485
rect 2051 1481 2052 1485
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 2046 1480 2052 1481
rect 2006 1476 2012 1477
rect 2054 1479 2060 1480
rect 1522 1475 1528 1476
rect 1522 1471 1523 1475
rect 1527 1471 1528 1475
rect 1522 1470 1528 1471
rect 1642 1475 1648 1476
rect 1642 1471 1643 1475
rect 1647 1471 1648 1475
rect 1642 1470 1648 1471
rect 1762 1475 1768 1476
rect 1762 1471 1763 1475
rect 1767 1471 1768 1475
rect 1762 1470 1768 1471
rect 1882 1475 1888 1476
rect 1882 1471 1883 1475
rect 1887 1471 1888 1475
rect 1882 1470 1888 1471
rect 1894 1475 1900 1476
rect 1894 1471 1895 1475
rect 1899 1471 1900 1475
rect 2054 1475 2055 1479
rect 2059 1475 2060 1479
rect 2054 1474 2060 1475
rect 1894 1470 1900 1471
rect 1454 1455 1460 1456
rect 1454 1451 1455 1455
rect 1459 1451 1460 1455
rect 1454 1450 1460 1451
rect 1524 1448 1526 1470
rect 1566 1465 1572 1466
rect 1566 1461 1567 1465
rect 1571 1461 1572 1465
rect 1566 1460 1572 1461
rect 1522 1447 1528 1448
rect 1522 1443 1523 1447
rect 1527 1443 1528 1447
rect 1522 1442 1528 1443
rect 1568 1439 1570 1460
rect 1644 1448 1646 1470
rect 1686 1465 1692 1466
rect 1686 1461 1687 1465
rect 1691 1461 1692 1465
rect 1686 1460 1692 1461
rect 1806 1465 1812 1466
rect 1806 1461 1807 1465
rect 1811 1461 1812 1465
rect 1806 1460 1812 1461
rect 1642 1447 1648 1448
rect 1642 1443 1643 1447
rect 1647 1443 1648 1447
rect 1642 1442 1648 1443
rect 1688 1439 1690 1460
rect 1808 1439 1810 1460
rect 975 1438 979 1439
rect 975 1433 979 1434
rect 1039 1438 1043 1439
rect 1039 1433 1043 1434
rect 1159 1438 1163 1439
rect 1159 1433 1163 1434
rect 1183 1438 1187 1439
rect 1242 1438 1248 1439
rect 1319 1438 1323 1439
rect 1183 1433 1187 1434
rect 954 1431 960 1432
rect 954 1427 955 1431
rect 959 1427 960 1431
rect 954 1426 960 1427
rect 976 1412 978 1433
rect 1050 1431 1056 1432
rect 1050 1427 1051 1431
rect 1055 1427 1056 1431
rect 1050 1426 1056 1427
rect 790 1411 796 1412
rect 790 1407 791 1411
rect 795 1407 796 1411
rect 790 1406 796 1407
rect 974 1411 980 1412
rect 974 1407 975 1411
rect 979 1407 980 1411
rect 974 1406 980 1407
rect 1052 1404 1054 1426
rect 1160 1412 1162 1433
rect 1158 1411 1164 1412
rect 1158 1407 1159 1411
rect 1163 1407 1164 1411
rect 1158 1406 1164 1407
rect 1244 1404 1246 1438
rect 1319 1433 1323 1434
rect 1351 1438 1355 1439
rect 1351 1433 1355 1434
rect 1447 1438 1451 1439
rect 1447 1433 1451 1434
rect 1543 1438 1547 1439
rect 1543 1433 1547 1434
rect 1567 1438 1571 1439
rect 1567 1433 1571 1434
rect 1687 1438 1691 1439
rect 1687 1433 1691 1434
rect 1735 1438 1739 1439
rect 1735 1433 1739 1434
rect 1807 1438 1811 1439
rect 1807 1433 1811 1434
rect 1352 1412 1354 1433
rect 1434 1431 1440 1432
rect 1434 1427 1435 1431
rect 1439 1427 1440 1431
rect 1434 1426 1440 1427
rect 1350 1411 1356 1412
rect 1350 1407 1351 1411
rect 1355 1407 1356 1411
rect 1350 1406 1356 1407
rect 1436 1404 1438 1426
rect 1544 1412 1546 1433
rect 1626 1431 1632 1432
rect 1626 1427 1627 1431
rect 1631 1427 1632 1431
rect 1626 1426 1632 1427
rect 1542 1411 1548 1412
rect 1542 1407 1543 1411
rect 1547 1407 1548 1411
rect 1542 1406 1548 1407
rect 1628 1404 1630 1426
rect 1736 1412 1738 1433
rect 1884 1432 1886 1470
rect 1896 1448 1898 1470
rect 2046 1468 2052 1469
rect 1902 1465 1908 1466
rect 1902 1461 1903 1465
rect 1907 1461 1908 1465
rect 1902 1460 1908 1461
rect 2006 1464 2012 1465
rect 2006 1460 2007 1464
rect 2011 1460 2012 1464
rect 2046 1464 2047 1468
rect 2051 1464 2052 1468
rect 2046 1463 2052 1464
rect 1894 1447 1900 1448
rect 1894 1443 1895 1447
rect 1899 1443 1900 1447
rect 1894 1442 1900 1443
rect 1904 1439 1906 1460
rect 2006 1459 2012 1460
rect 2008 1439 2010 1459
rect 1903 1438 1907 1439
rect 1903 1433 1907 1434
rect 2007 1438 2011 1439
rect 2048 1435 2050 1463
rect 2056 1448 2058 1474
rect 2070 1469 2076 1470
rect 2070 1465 2071 1469
rect 2075 1465 2076 1469
rect 2070 1464 2076 1465
rect 2054 1447 2060 1448
rect 2054 1443 2055 1447
rect 2059 1443 2060 1447
rect 2054 1442 2060 1443
rect 2072 1435 2074 1464
rect 2420 1452 2422 1554
rect 2494 1548 2500 1549
rect 2494 1544 2495 1548
rect 2499 1544 2500 1548
rect 2494 1543 2500 1544
rect 2710 1548 2716 1549
rect 2710 1544 2711 1548
rect 2715 1544 2716 1548
rect 2710 1543 2716 1544
rect 2910 1548 2916 1549
rect 2910 1544 2911 1548
rect 2915 1544 2916 1548
rect 2910 1543 2916 1544
rect 3094 1548 3100 1549
rect 3094 1544 3095 1548
rect 3099 1544 3100 1548
rect 3094 1543 3100 1544
rect 2496 1519 2498 1543
rect 2712 1519 2714 1543
rect 2912 1519 2914 1543
rect 3096 1519 3098 1543
rect 2431 1518 2435 1519
rect 2431 1513 2435 1514
rect 2495 1518 2499 1519
rect 2495 1513 2499 1514
rect 2711 1518 2715 1519
rect 2711 1513 2715 1514
rect 2791 1518 2795 1519
rect 2791 1513 2795 1514
rect 2911 1518 2915 1519
rect 2911 1513 2915 1514
rect 3095 1518 3099 1519
rect 3095 1513 3099 1514
rect 3127 1518 3131 1519
rect 3127 1513 3131 1514
rect 2432 1489 2434 1513
rect 2792 1489 2794 1513
rect 3128 1489 3130 1513
rect 2430 1488 2436 1489
rect 2430 1484 2431 1488
rect 2435 1484 2436 1488
rect 2430 1483 2436 1484
rect 2790 1488 2796 1489
rect 2790 1484 2791 1488
rect 2795 1484 2796 1488
rect 2790 1483 2796 1484
rect 3126 1488 3132 1489
rect 3126 1484 3127 1488
rect 3131 1484 3132 1488
rect 3126 1483 3132 1484
rect 3204 1480 3206 1582
rect 3264 1568 3266 1589
rect 3338 1587 3344 1588
rect 3338 1583 3339 1587
rect 3343 1583 3344 1587
rect 3338 1582 3344 1583
rect 3262 1567 3268 1568
rect 3262 1563 3263 1567
rect 3267 1563 3268 1567
rect 3262 1562 3268 1563
rect 3340 1560 3342 1582
rect 3400 1560 3402 1602
rect 3528 1595 3530 1624
rect 3604 1612 3606 1634
rect 3694 1629 3700 1630
rect 3694 1625 3695 1629
rect 3699 1625 3700 1629
rect 3694 1624 3700 1625
rect 3602 1611 3608 1612
rect 3602 1607 3603 1611
rect 3607 1607 3608 1611
rect 3602 1606 3608 1607
rect 3696 1595 3698 1624
rect 3423 1594 3427 1595
rect 3423 1589 3427 1590
rect 3527 1594 3531 1595
rect 3527 1589 3531 1590
rect 3567 1594 3571 1595
rect 3567 1589 3571 1590
rect 3695 1594 3699 1595
rect 3695 1589 3699 1590
rect 3711 1594 3715 1595
rect 3711 1589 3715 1590
rect 3424 1568 3426 1589
rect 3568 1568 3570 1589
rect 3712 1568 3714 1589
rect 3422 1567 3428 1568
rect 3422 1563 3423 1567
rect 3427 1563 3428 1567
rect 3422 1562 3428 1563
rect 3566 1567 3572 1568
rect 3566 1563 3567 1567
rect 3571 1563 3572 1567
rect 3566 1562 3572 1563
rect 3710 1567 3716 1568
rect 3710 1563 3711 1567
rect 3715 1563 3716 1567
rect 3710 1562 3716 1563
rect 3800 1560 3802 1754
rect 3839 1678 3843 1679
rect 3839 1673 3843 1674
rect 3840 1649 3842 1673
rect 3838 1648 3844 1649
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 3906 1639 3912 1640
rect 3906 1635 3907 1639
rect 3911 1635 3912 1639
rect 3906 1634 3912 1635
rect 3838 1629 3844 1630
rect 3838 1625 3839 1629
rect 3843 1625 3844 1629
rect 3838 1624 3844 1625
rect 3840 1595 3842 1624
rect 3839 1594 3843 1595
rect 3839 1589 3843 1590
rect 3806 1587 3812 1588
rect 3806 1583 3807 1587
rect 3811 1583 3812 1587
rect 3806 1582 3812 1583
rect 3808 1560 3810 1582
rect 3840 1568 3842 1589
rect 3908 1588 3910 1634
rect 3916 1612 3918 1862
rect 3942 1859 3943 1863
rect 3947 1859 3948 1863
rect 3942 1858 3948 1859
rect 3944 1831 3946 1858
rect 3943 1830 3947 1831
rect 3943 1825 3947 1826
rect 3944 1798 3946 1825
rect 3942 1797 3948 1798
rect 3942 1793 3943 1797
rect 3947 1793 3948 1797
rect 3942 1792 3948 1793
rect 3942 1780 3948 1781
rect 3942 1776 3943 1780
rect 3947 1776 3948 1780
rect 3942 1775 3948 1776
rect 3944 1755 3946 1775
rect 3943 1754 3947 1755
rect 3943 1749 3947 1750
rect 3944 1729 3946 1749
rect 3942 1728 3948 1729
rect 3942 1724 3943 1728
rect 3947 1724 3948 1728
rect 3942 1723 3948 1724
rect 3942 1711 3948 1712
rect 3942 1707 3943 1711
rect 3947 1707 3948 1711
rect 3942 1706 3948 1707
rect 3944 1679 3946 1706
rect 3943 1678 3947 1679
rect 3943 1673 3947 1674
rect 3944 1646 3946 1673
rect 3942 1645 3948 1646
rect 3942 1641 3943 1645
rect 3947 1641 3948 1645
rect 3942 1640 3948 1641
rect 3942 1628 3948 1629
rect 3942 1624 3943 1628
rect 3947 1624 3948 1628
rect 3942 1623 3948 1624
rect 3914 1611 3920 1612
rect 3914 1607 3915 1611
rect 3919 1607 3920 1611
rect 3914 1606 3920 1607
rect 3944 1595 3946 1623
rect 3943 1594 3947 1595
rect 3943 1589 3947 1590
rect 3906 1587 3912 1588
rect 3906 1583 3907 1587
rect 3911 1583 3912 1587
rect 3906 1582 3912 1583
rect 3944 1569 3946 1589
rect 3942 1568 3948 1569
rect 3838 1567 3844 1568
rect 3838 1563 3839 1567
rect 3843 1563 3844 1567
rect 3942 1564 3943 1568
rect 3947 1564 3948 1568
rect 3942 1563 3948 1564
rect 3838 1562 3844 1563
rect 3338 1559 3344 1560
rect 3338 1555 3339 1559
rect 3343 1555 3344 1559
rect 3338 1554 3344 1555
rect 3398 1559 3404 1560
rect 3398 1555 3399 1559
rect 3403 1555 3404 1559
rect 3398 1554 3404 1555
rect 3506 1559 3512 1560
rect 3506 1555 3507 1559
rect 3511 1555 3512 1559
rect 3506 1554 3512 1555
rect 3798 1559 3804 1560
rect 3798 1555 3799 1559
rect 3803 1555 3804 1559
rect 3798 1554 3804 1555
rect 3806 1559 3812 1560
rect 3806 1555 3807 1559
rect 3811 1555 3812 1559
rect 3806 1554 3812 1555
rect 3262 1548 3268 1549
rect 3262 1544 3263 1548
rect 3267 1544 3268 1548
rect 3262 1543 3268 1544
rect 3422 1548 3428 1549
rect 3422 1544 3423 1548
rect 3427 1544 3428 1548
rect 3422 1543 3428 1544
rect 3264 1519 3266 1543
rect 3424 1519 3426 1543
rect 3263 1518 3267 1519
rect 3263 1513 3267 1514
rect 3423 1518 3427 1519
rect 3423 1513 3427 1514
rect 3463 1518 3467 1519
rect 3463 1513 3467 1514
rect 3464 1489 3466 1513
rect 3508 1499 3510 1554
rect 3942 1551 3948 1552
rect 3566 1548 3572 1549
rect 3566 1544 3567 1548
rect 3571 1544 3572 1548
rect 3566 1543 3572 1544
rect 3710 1548 3716 1549
rect 3710 1544 3711 1548
rect 3715 1544 3716 1548
rect 3710 1543 3716 1544
rect 3838 1548 3844 1549
rect 3838 1544 3839 1548
rect 3843 1544 3844 1548
rect 3942 1547 3943 1551
rect 3947 1547 3948 1551
rect 3942 1546 3948 1547
rect 3838 1543 3844 1544
rect 3568 1519 3570 1543
rect 3712 1519 3714 1543
rect 3840 1519 3842 1543
rect 3944 1519 3946 1546
rect 3567 1518 3571 1519
rect 3567 1513 3571 1514
rect 3711 1518 3715 1519
rect 3711 1513 3715 1514
rect 3799 1518 3803 1519
rect 3799 1513 3803 1514
rect 3839 1518 3843 1519
rect 3839 1513 3843 1514
rect 3943 1518 3947 1519
rect 3943 1513 3947 1514
rect 3504 1497 3510 1499
rect 3462 1488 3468 1489
rect 3462 1484 3463 1488
rect 3467 1484 3468 1488
rect 3462 1483 3468 1484
rect 2718 1479 2724 1480
rect 2718 1475 2719 1479
rect 2723 1475 2724 1479
rect 2718 1474 2724 1475
rect 2866 1479 2872 1480
rect 2866 1475 2867 1479
rect 2871 1475 2872 1479
rect 2866 1474 2872 1475
rect 3202 1479 3208 1480
rect 3202 1475 3203 1479
rect 3207 1475 3208 1479
rect 3202 1474 3208 1475
rect 2430 1469 2436 1470
rect 2430 1465 2431 1469
rect 2435 1465 2436 1469
rect 2430 1464 2436 1465
rect 2418 1451 2424 1452
rect 2418 1447 2419 1451
rect 2423 1447 2424 1451
rect 2418 1446 2424 1447
rect 2432 1435 2434 1464
rect 2720 1452 2722 1474
rect 2790 1469 2796 1470
rect 2790 1465 2791 1469
rect 2795 1465 2796 1469
rect 2790 1464 2796 1465
rect 2718 1451 2724 1452
rect 2718 1447 2719 1451
rect 2723 1447 2724 1451
rect 2718 1446 2724 1447
rect 2792 1435 2794 1464
rect 2007 1433 2011 1434
rect 2047 1434 2051 1435
rect 1742 1431 1748 1432
rect 1742 1427 1743 1431
rect 1747 1427 1748 1431
rect 1742 1426 1748 1427
rect 1882 1431 1888 1432
rect 1882 1427 1883 1431
rect 1887 1427 1888 1431
rect 1882 1426 1888 1427
rect 1734 1411 1740 1412
rect 1734 1407 1735 1411
rect 1739 1407 1740 1411
rect 1734 1406 1740 1407
rect 682 1403 688 1404
rect 682 1399 683 1403
rect 687 1399 688 1403
rect 682 1398 688 1399
rect 690 1403 696 1404
rect 690 1399 691 1403
rect 695 1399 696 1403
rect 690 1398 696 1399
rect 1050 1403 1056 1404
rect 1050 1399 1051 1403
rect 1055 1399 1056 1403
rect 1050 1398 1056 1399
rect 1082 1403 1088 1404
rect 1082 1399 1083 1403
rect 1087 1399 1088 1403
rect 1082 1398 1088 1399
rect 1242 1403 1248 1404
rect 1242 1399 1243 1403
rect 1247 1399 1248 1403
rect 1242 1398 1248 1399
rect 1434 1403 1440 1404
rect 1434 1399 1435 1403
rect 1439 1399 1440 1403
rect 1434 1398 1440 1399
rect 1626 1403 1632 1404
rect 1626 1399 1627 1403
rect 1631 1399 1632 1403
rect 1626 1398 1632 1399
rect 606 1392 612 1393
rect 606 1388 607 1392
rect 611 1388 612 1392
rect 606 1387 612 1388
rect 790 1392 796 1393
rect 790 1388 791 1392
rect 795 1388 796 1392
rect 790 1387 796 1388
rect 974 1392 980 1393
rect 974 1388 975 1392
rect 979 1388 980 1392
rect 974 1387 980 1388
rect 608 1359 610 1387
rect 792 1359 794 1387
rect 976 1359 978 1387
rect 607 1358 611 1359
rect 607 1353 611 1354
rect 663 1358 667 1359
rect 663 1353 667 1354
rect 791 1358 795 1359
rect 791 1353 795 1354
rect 855 1358 859 1359
rect 855 1353 859 1354
rect 975 1358 979 1359
rect 975 1353 979 1354
rect 1047 1358 1051 1359
rect 1047 1353 1051 1354
rect 664 1329 666 1353
rect 856 1329 858 1353
rect 1048 1329 1050 1353
rect 662 1328 668 1329
rect 662 1324 663 1328
rect 667 1324 668 1328
rect 662 1323 668 1324
rect 854 1328 860 1329
rect 854 1324 855 1328
rect 859 1324 860 1328
rect 854 1323 860 1324
rect 1046 1328 1052 1329
rect 1046 1324 1047 1328
rect 1051 1324 1052 1328
rect 1046 1323 1052 1324
rect 262 1319 268 1320
rect 262 1315 263 1319
rect 267 1315 268 1319
rect 262 1314 268 1315
rect 386 1319 392 1320
rect 386 1315 387 1319
rect 391 1315 392 1319
rect 386 1314 392 1315
rect 578 1319 584 1320
rect 578 1315 579 1319
rect 583 1315 584 1319
rect 578 1314 584 1315
rect 738 1319 744 1320
rect 738 1315 739 1319
rect 743 1315 744 1319
rect 738 1314 744 1315
rect 746 1319 752 1320
rect 746 1315 747 1319
rect 751 1315 752 1319
rect 746 1314 752 1315
rect 158 1309 164 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 158 1305 159 1309
rect 163 1305 164 1309
rect 158 1304 164 1305
rect 110 1303 116 1304
rect 112 1279 114 1303
rect 160 1279 162 1304
rect 264 1288 266 1314
rect 310 1309 316 1310
rect 310 1305 311 1309
rect 315 1305 316 1309
rect 310 1304 316 1305
rect 262 1287 268 1288
rect 262 1283 263 1287
rect 267 1283 268 1287
rect 262 1282 268 1283
rect 312 1279 314 1304
rect 388 1292 390 1314
rect 478 1309 484 1310
rect 478 1305 479 1309
rect 483 1305 484 1309
rect 478 1304 484 1305
rect 662 1309 668 1310
rect 662 1305 663 1309
rect 667 1305 668 1309
rect 662 1304 668 1305
rect 386 1291 392 1292
rect 386 1287 387 1291
rect 391 1287 392 1291
rect 386 1286 392 1287
rect 480 1279 482 1304
rect 618 1287 624 1288
rect 618 1283 619 1287
rect 623 1283 624 1287
rect 618 1282 624 1283
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 159 1278 163 1279
rect 159 1273 163 1274
rect 311 1278 315 1279
rect 311 1273 315 1274
rect 407 1278 411 1279
rect 407 1273 411 1274
rect 479 1278 483 1279
rect 479 1273 483 1274
rect 543 1278 547 1279
rect 543 1273 547 1274
rect 112 1253 114 1273
rect 110 1252 116 1253
rect 408 1252 410 1273
rect 446 1271 452 1272
rect 446 1266 447 1271
rect 451 1266 452 1271
rect 447 1263 451 1264
rect 544 1252 546 1273
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 406 1251 412 1252
rect 406 1247 407 1251
rect 411 1247 412 1251
rect 406 1246 412 1247
rect 542 1251 548 1252
rect 542 1247 543 1251
rect 547 1247 548 1251
rect 542 1246 548 1247
rect 620 1244 622 1282
rect 664 1279 666 1304
rect 740 1292 742 1314
rect 748 1300 750 1314
rect 854 1309 860 1310
rect 854 1305 855 1309
rect 859 1305 860 1309
rect 854 1304 860 1305
rect 1046 1309 1052 1310
rect 1046 1305 1047 1309
rect 1051 1305 1052 1309
rect 1046 1304 1052 1305
rect 746 1299 752 1300
rect 746 1295 747 1299
rect 751 1295 752 1299
rect 746 1294 752 1295
rect 738 1291 744 1292
rect 738 1287 739 1291
rect 743 1287 744 1291
rect 738 1286 744 1287
rect 856 1279 858 1304
rect 1048 1279 1050 1304
rect 1084 1292 1086 1398
rect 1158 1392 1164 1393
rect 1158 1388 1159 1392
rect 1163 1388 1164 1392
rect 1158 1387 1164 1388
rect 1350 1392 1356 1393
rect 1350 1388 1351 1392
rect 1355 1388 1356 1392
rect 1350 1387 1356 1388
rect 1542 1392 1548 1393
rect 1542 1388 1543 1392
rect 1547 1388 1548 1392
rect 1542 1387 1548 1388
rect 1734 1392 1740 1393
rect 1734 1388 1735 1392
rect 1739 1388 1740 1392
rect 1734 1387 1740 1388
rect 1160 1359 1162 1387
rect 1352 1359 1354 1387
rect 1544 1359 1546 1387
rect 1736 1359 1738 1387
rect 1159 1358 1163 1359
rect 1159 1353 1163 1354
rect 1247 1358 1251 1359
rect 1247 1353 1251 1354
rect 1351 1358 1355 1359
rect 1351 1353 1355 1354
rect 1447 1358 1451 1359
rect 1447 1353 1451 1354
rect 1543 1358 1547 1359
rect 1543 1353 1547 1354
rect 1655 1358 1659 1359
rect 1655 1353 1659 1354
rect 1735 1358 1739 1359
rect 1735 1353 1739 1354
rect 1248 1329 1250 1353
rect 1448 1329 1450 1353
rect 1656 1329 1658 1353
rect 1246 1328 1252 1329
rect 1246 1324 1247 1328
rect 1251 1324 1252 1328
rect 1246 1323 1252 1324
rect 1446 1328 1452 1329
rect 1446 1324 1447 1328
rect 1451 1324 1452 1328
rect 1446 1323 1452 1324
rect 1654 1328 1660 1329
rect 1654 1324 1655 1328
rect 1659 1324 1660 1328
rect 1654 1323 1660 1324
rect 1744 1320 1746 1426
rect 1904 1412 1906 1433
rect 1978 1427 1984 1428
rect 1978 1423 1979 1427
rect 1983 1423 1984 1427
rect 1978 1422 1984 1423
rect 1902 1411 1908 1412
rect 1902 1407 1903 1411
rect 1907 1407 1908 1411
rect 1902 1406 1908 1407
rect 1980 1404 1982 1422
rect 2008 1413 2010 1433
rect 2047 1429 2051 1430
rect 2071 1434 2075 1435
rect 2071 1429 2075 1430
rect 2271 1434 2275 1435
rect 2271 1429 2275 1430
rect 2431 1434 2435 1435
rect 2431 1429 2435 1430
rect 2495 1434 2499 1435
rect 2495 1429 2499 1430
rect 2711 1434 2715 1435
rect 2711 1429 2715 1430
rect 2791 1434 2795 1435
rect 2791 1429 2795 1430
rect 2006 1412 2012 1413
rect 2006 1408 2007 1412
rect 2011 1408 2012 1412
rect 2048 1409 2050 1429
rect 2006 1407 2012 1408
rect 2046 1408 2052 1409
rect 2072 1408 2074 1429
rect 2146 1427 2152 1428
rect 2146 1423 2147 1427
rect 2151 1423 2152 1427
rect 2146 1422 2152 1423
rect 2046 1404 2047 1408
rect 2051 1404 2052 1408
rect 1978 1403 1984 1404
rect 2046 1403 2052 1404
rect 2070 1407 2076 1408
rect 2070 1403 2071 1407
rect 2075 1403 2076 1407
rect 1978 1399 1979 1403
rect 1983 1399 1984 1403
rect 2070 1402 2076 1403
rect 2148 1400 2150 1422
rect 2272 1408 2274 1429
rect 2346 1427 2352 1428
rect 2346 1423 2347 1427
rect 2351 1423 2352 1427
rect 2346 1422 2352 1423
rect 2270 1407 2276 1408
rect 2270 1403 2271 1407
rect 2275 1403 2276 1407
rect 2270 1402 2276 1403
rect 2348 1400 2350 1422
rect 2496 1408 2498 1429
rect 2570 1427 2576 1428
rect 2570 1423 2571 1427
rect 2575 1423 2576 1427
rect 2570 1422 2576 1423
rect 2494 1407 2500 1408
rect 2494 1403 2495 1407
rect 2499 1403 2500 1407
rect 2494 1402 2500 1403
rect 2572 1400 2574 1422
rect 2712 1408 2714 1429
rect 2868 1428 2870 1474
rect 3126 1469 3132 1470
rect 3126 1465 3127 1469
rect 3131 1465 3132 1469
rect 3126 1464 3132 1465
rect 3462 1469 3468 1470
rect 3462 1465 3463 1469
rect 3467 1465 3468 1469
rect 3462 1464 3468 1465
rect 3128 1435 3130 1464
rect 3166 1447 3172 1448
rect 3166 1443 3167 1447
rect 3171 1443 3172 1447
rect 3166 1442 3174 1443
rect 3168 1441 3174 1442
rect 2911 1434 2915 1435
rect 2911 1429 2915 1430
rect 3095 1434 3099 1435
rect 3095 1429 3099 1430
rect 3127 1434 3131 1435
rect 3127 1429 3131 1430
rect 2866 1427 2872 1428
rect 2866 1423 2867 1427
rect 2871 1423 2872 1427
rect 2866 1422 2872 1423
rect 2912 1408 2914 1429
rect 2986 1427 2992 1428
rect 2986 1423 2987 1427
rect 2991 1423 2992 1427
rect 2986 1422 2992 1423
rect 2710 1407 2716 1408
rect 2710 1403 2711 1407
rect 2715 1403 2716 1407
rect 2710 1402 2716 1403
rect 2910 1407 2916 1408
rect 2910 1403 2911 1407
rect 2915 1403 2916 1407
rect 2910 1402 2916 1403
rect 2988 1400 2990 1422
rect 3096 1408 3098 1429
rect 3094 1407 3100 1408
rect 3094 1403 3095 1407
rect 3099 1403 3100 1407
rect 3094 1402 3100 1403
rect 3172 1400 3174 1441
rect 3464 1435 3466 1464
rect 3504 1452 3506 1497
rect 3800 1489 3802 1513
rect 3798 1488 3804 1489
rect 3798 1484 3799 1488
rect 3803 1484 3804 1488
rect 3944 1486 3946 1513
rect 3798 1483 3804 1484
rect 3942 1485 3948 1486
rect 3942 1481 3943 1485
rect 3947 1481 3948 1485
rect 3942 1480 3948 1481
rect 3538 1479 3544 1480
rect 3538 1475 3539 1479
rect 3543 1475 3544 1479
rect 3538 1474 3544 1475
rect 3866 1479 3872 1480
rect 3866 1475 3867 1479
rect 3871 1475 3872 1479
rect 3866 1474 3872 1475
rect 3540 1452 3542 1474
rect 3798 1469 3804 1470
rect 3798 1465 3799 1469
rect 3803 1465 3804 1469
rect 3798 1464 3804 1465
rect 3502 1451 3508 1452
rect 3502 1447 3503 1451
rect 3507 1447 3508 1451
rect 3502 1446 3508 1447
rect 3538 1451 3544 1452
rect 3538 1447 3539 1451
rect 3543 1447 3544 1451
rect 3538 1446 3544 1447
rect 3800 1435 3802 1464
rect 3271 1434 3275 1435
rect 3271 1429 3275 1430
rect 3439 1434 3443 1435
rect 3439 1429 3443 1430
rect 3463 1434 3467 1435
rect 3463 1429 3467 1430
rect 3607 1434 3611 1435
rect 3607 1429 3611 1430
rect 3783 1434 3787 1435
rect 3783 1429 3787 1430
rect 3799 1434 3803 1435
rect 3799 1429 3803 1430
rect 3272 1408 3274 1429
rect 3354 1427 3360 1428
rect 3354 1423 3355 1427
rect 3359 1423 3360 1427
rect 3354 1422 3360 1423
rect 3270 1407 3276 1408
rect 3270 1403 3271 1407
rect 3275 1403 3276 1407
rect 3270 1402 3276 1403
rect 3356 1400 3358 1422
rect 3440 1408 3442 1429
rect 3506 1427 3512 1428
rect 3506 1423 3507 1427
rect 3511 1423 3512 1427
rect 3506 1422 3512 1423
rect 3522 1427 3528 1428
rect 3522 1423 3523 1427
rect 3527 1423 3528 1427
rect 3522 1422 3528 1423
rect 3438 1407 3444 1408
rect 3438 1403 3439 1407
rect 3443 1403 3444 1407
rect 3508 1404 3510 1422
rect 3438 1402 3444 1403
rect 3506 1403 3512 1404
rect 1978 1398 1984 1399
rect 2146 1399 2152 1400
rect 2006 1395 2012 1396
rect 1902 1392 1908 1393
rect 1902 1388 1903 1392
rect 1907 1388 1908 1392
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2146 1395 2147 1399
rect 2151 1395 2152 1399
rect 2146 1394 2152 1395
rect 2346 1399 2352 1400
rect 2346 1395 2347 1399
rect 2351 1395 2352 1399
rect 2346 1394 2352 1395
rect 2570 1399 2576 1400
rect 2570 1395 2571 1399
rect 2575 1395 2576 1399
rect 2570 1394 2576 1395
rect 2658 1399 2664 1400
rect 2658 1395 2659 1399
rect 2663 1395 2664 1399
rect 2658 1394 2664 1395
rect 2986 1399 2992 1400
rect 2986 1395 2987 1399
rect 2991 1395 2992 1399
rect 2986 1394 2992 1395
rect 3170 1399 3176 1400
rect 3170 1395 3171 1399
rect 3175 1395 3176 1399
rect 3170 1394 3176 1395
rect 3198 1399 3204 1400
rect 3198 1395 3199 1399
rect 3203 1395 3204 1399
rect 3198 1394 3204 1395
rect 3354 1399 3360 1400
rect 3354 1395 3355 1399
rect 3359 1395 3360 1399
rect 3506 1399 3507 1403
rect 3511 1399 3512 1403
rect 3506 1398 3512 1399
rect 3354 1394 3360 1395
rect 2006 1390 2012 1391
rect 2046 1391 2052 1392
rect 1902 1387 1908 1388
rect 1904 1359 1906 1387
rect 2008 1359 2010 1390
rect 2046 1387 2047 1391
rect 2051 1387 2052 1391
rect 2046 1386 2052 1387
rect 2070 1388 2076 1389
rect 2048 1359 2050 1386
rect 2070 1384 2071 1388
rect 2075 1384 2076 1388
rect 2070 1383 2076 1384
rect 2270 1388 2276 1389
rect 2270 1384 2271 1388
rect 2275 1384 2276 1388
rect 2270 1383 2276 1384
rect 2494 1388 2500 1389
rect 2494 1384 2495 1388
rect 2499 1384 2500 1388
rect 2494 1383 2500 1384
rect 2072 1359 2074 1383
rect 2272 1359 2274 1383
rect 2496 1359 2498 1383
rect 1863 1358 1867 1359
rect 1863 1353 1867 1354
rect 1903 1358 1907 1359
rect 1903 1353 1907 1354
rect 2007 1358 2011 1359
rect 2007 1353 2011 1354
rect 2047 1358 2051 1359
rect 2047 1353 2051 1354
rect 2071 1358 2075 1359
rect 2071 1353 2075 1354
rect 2207 1358 2211 1359
rect 2207 1353 2211 1354
rect 2271 1358 2275 1359
rect 2271 1353 2275 1354
rect 2383 1358 2387 1359
rect 2383 1353 2387 1354
rect 2495 1358 2499 1359
rect 2495 1353 2499 1354
rect 2567 1358 2571 1359
rect 2567 1353 2571 1354
rect 1864 1329 1866 1353
rect 1862 1328 1868 1329
rect 1862 1324 1863 1328
rect 1867 1324 1868 1328
rect 2008 1326 2010 1353
rect 2048 1326 2050 1353
rect 2072 1329 2074 1353
rect 2208 1329 2210 1353
rect 2384 1329 2386 1353
rect 2568 1329 2570 1353
rect 2070 1328 2076 1329
rect 1862 1323 1868 1324
rect 2006 1325 2012 1326
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2046 1325 2052 1326
rect 2046 1321 2047 1325
rect 2051 1321 2052 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2206 1328 2212 1329
rect 2206 1324 2207 1328
rect 2211 1324 2212 1328
rect 2206 1323 2212 1324
rect 2382 1328 2388 1329
rect 2382 1324 2383 1328
rect 2387 1324 2388 1328
rect 2382 1323 2388 1324
rect 2566 1328 2572 1329
rect 2566 1324 2567 1328
rect 2571 1324 2572 1328
rect 2566 1323 2572 1324
rect 2046 1320 2052 1321
rect 1122 1319 1128 1320
rect 1122 1315 1123 1319
rect 1127 1315 1128 1319
rect 1122 1314 1128 1315
rect 1322 1319 1328 1320
rect 1322 1315 1323 1319
rect 1327 1315 1328 1319
rect 1322 1314 1328 1315
rect 1522 1319 1528 1320
rect 1522 1315 1523 1319
rect 1527 1315 1528 1319
rect 1522 1314 1528 1315
rect 1742 1319 1748 1320
rect 1742 1315 1743 1319
rect 1747 1315 1748 1319
rect 1742 1314 1748 1315
rect 2146 1319 2152 1320
rect 2146 1315 2147 1319
rect 2151 1315 2152 1319
rect 2146 1314 2152 1315
rect 2282 1319 2288 1320
rect 2282 1315 2283 1319
rect 2287 1315 2288 1319
rect 2282 1314 2288 1315
rect 2458 1319 2464 1320
rect 2458 1315 2459 1319
rect 2463 1315 2464 1319
rect 2458 1314 2464 1315
rect 2642 1319 2648 1320
rect 2642 1315 2643 1319
rect 2647 1315 2648 1319
rect 2642 1314 2648 1315
rect 1124 1292 1126 1314
rect 1246 1309 1252 1310
rect 1246 1305 1247 1309
rect 1251 1305 1252 1309
rect 1246 1304 1252 1305
rect 1082 1291 1088 1292
rect 1082 1287 1083 1291
rect 1087 1287 1088 1291
rect 1082 1286 1088 1287
rect 1122 1291 1128 1292
rect 1122 1287 1123 1291
rect 1127 1287 1128 1291
rect 1122 1286 1128 1287
rect 1248 1279 1250 1304
rect 1324 1292 1326 1314
rect 1446 1309 1452 1310
rect 1446 1305 1447 1309
rect 1451 1305 1452 1309
rect 1446 1304 1452 1305
rect 1322 1291 1328 1292
rect 1322 1287 1323 1291
rect 1327 1287 1328 1291
rect 1322 1286 1328 1287
rect 1448 1279 1450 1304
rect 663 1278 667 1279
rect 663 1273 667 1274
rect 695 1278 699 1279
rect 695 1273 699 1274
rect 855 1278 859 1279
rect 855 1273 859 1274
rect 1023 1278 1027 1279
rect 1023 1273 1027 1274
rect 1047 1278 1051 1279
rect 1047 1273 1051 1274
rect 1191 1278 1195 1279
rect 1191 1273 1195 1274
rect 1247 1278 1251 1279
rect 1247 1273 1251 1274
rect 1367 1278 1371 1279
rect 1367 1273 1371 1274
rect 1447 1278 1451 1279
rect 1447 1273 1451 1274
rect 674 1271 680 1272
rect 674 1267 675 1271
rect 679 1267 680 1271
rect 674 1266 680 1267
rect 618 1243 624 1244
rect 618 1239 619 1243
rect 623 1239 624 1243
rect 618 1238 624 1239
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 406 1232 412 1233
rect 112 1203 114 1230
rect 406 1228 407 1232
rect 411 1228 412 1232
rect 406 1227 412 1228
rect 542 1232 548 1233
rect 542 1228 543 1232
rect 547 1228 548 1232
rect 542 1227 548 1228
rect 408 1203 410 1227
rect 544 1203 546 1227
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 407 1202 411 1203
rect 407 1197 411 1198
rect 423 1202 427 1203
rect 423 1197 427 1198
rect 543 1202 547 1203
rect 543 1197 547 1198
rect 591 1202 595 1203
rect 591 1197 595 1198
rect 112 1170 114 1197
rect 424 1173 426 1197
rect 592 1173 594 1197
rect 422 1172 428 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 422 1168 423 1172
rect 427 1168 428 1172
rect 422 1167 428 1168
rect 590 1172 596 1173
rect 590 1168 591 1172
rect 595 1168 596 1172
rect 590 1167 596 1168
rect 110 1164 116 1165
rect 676 1164 678 1266
rect 696 1252 698 1273
rect 770 1271 776 1272
rect 770 1267 771 1271
rect 775 1267 776 1271
rect 770 1266 776 1267
rect 694 1251 700 1252
rect 694 1247 695 1251
rect 699 1247 700 1251
rect 694 1246 700 1247
rect 772 1244 774 1266
rect 856 1252 858 1273
rect 930 1271 936 1272
rect 930 1267 931 1271
rect 935 1267 936 1271
rect 930 1266 936 1267
rect 979 1268 983 1269
rect 854 1251 860 1252
rect 854 1247 855 1251
rect 859 1247 860 1251
rect 854 1246 860 1247
rect 932 1244 934 1266
rect 979 1263 983 1264
rect 980 1244 982 1263
rect 1024 1252 1026 1273
rect 1192 1252 1194 1273
rect 1274 1271 1280 1272
rect 1274 1267 1275 1271
rect 1279 1267 1280 1271
rect 1274 1266 1280 1267
rect 1022 1251 1028 1252
rect 1022 1247 1023 1251
rect 1027 1247 1028 1251
rect 1022 1246 1028 1247
rect 1190 1251 1196 1252
rect 1190 1247 1191 1251
rect 1195 1247 1196 1251
rect 1190 1246 1196 1247
rect 1276 1244 1278 1266
rect 1368 1252 1370 1273
rect 1524 1272 1526 1314
rect 1654 1309 1660 1310
rect 1654 1305 1655 1309
rect 1659 1305 1660 1309
rect 1654 1304 1660 1305
rect 1862 1309 1868 1310
rect 2070 1309 2076 1310
rect 1862 1305 1863 1309
rect 1867 1305 1868 1309
rect 1862 1304 1868 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 1656 1279 1658 1304
rect 1864 1279 1866 1304
rect 2006 1303 2012 1304
rect 2046 1308 2052 1309
rect 2046 1304 2047 1308
rect 2051 1304 2052 1308
rect 2070 1305 2071 1309
rect 2075 1305 2076 1309
rect 2070 1304 2076 1305
rect 2046 1303 2052 1304
rect 2008 1279 2010 1303
rect 2048 1283 2050 1303
rect 2072 1283 2074 1304
rect 2148 1292 2150 1314
rect 2206 1309 2212 1310
rect 2206 1305 2207 1309
rect 2211 1305 2212 1309
rect 2206 1304 2212 1305
rect 2146 1291 2152 1292
rect 2146 1287 2147 1291
rect 2151 1287 2152 1291
rect 2146 1286 2152 1287
rect 2208 1283 2210 1304
rect 2284 1292 2286 1314
rect 2382 1309 2388 1310
rect 2382 1305 2383 1309
rect 2387 1305 2388 1309
rect 2382 1304 2388 1305
rect 2282 1291 2288 1292
rect 2282 1287 2283 1291
rect 2287 1287 2288 1291
rect 2282 1286 2288 1287
rect 2384 1283 2386 1304
rect 2460 1292 2462 1314
rect 2566 1309 2572 1310
rect 2566 1305 2567 1309
rect 2571 1305 2572 1309
rect 2566 1304 2572 1305
rect 2458 1291 2464 1292
rect 2458 1287 2459 1291
rect 2463 1287 2464 1291
rect 2458 1286 2464 1287
rect 2568 1283 2570 1304
rect 2644 1292 2646 1314
rect 2660 1300 2662 1394
rect 2710 1388 2716 1389
rect 2710 1384 2711 1388
rect 2715 1384 2716 1388
rect 2710 1383 2716 1384
rect 2910 1388 2916 1389
rect 2910 1384 2911 1388
rect 2915 1384 2916 1388
rect 2910 1383 2916 1384
rect 3094 1388 3100 1389
rect 3094 1384 3095 1388
rect 3099 1384 3100 1388
rect 3094 1383 3100 1384
rect 2712 1359 2714 1383
rect 2912 1359 2914 1383
rect 3096 1359 3098 1383
rect 2711 1358 2715 1359
rect 2711 1353 2715 1354
rect 2751 1358 2755 1359
rect 2751 1353 2755 1354
rect 2911 1358 2915 1359
rect 2911 1353 2915 1354
rect 2935 1358 2939 1359
rect 2935 1353 2939 1354
rect 3095 1358 3099 1359
rect 3095 1353 3099 1354
rect 3111 1358 3115 1359
rect 3111 1353 3115 1354
rect 2752 1329 2754 1353
rect 2936 1329 2938 1353
rect 3112 1329 3114 1353
rect 2750 1328 2756 1329
rect 2750 1324 2751 1328
rect 2755 1324 2756 1328
rect 2750 1323 2756 1324
rect 2934 1328 2940 1329
rect 2934 1324 2935 1328
rect 2939 1324 2940 1328
rect 2934 1323 2940 1324
rect 3110 1328 3116 1329
rect 3110 1324 3111 1328
rect 3115 1324 3116 1328
rect 3110 1323 3116 1324
rect 2718 1319 2724 1320
rect 2718 1315 2719 1319
rect 2723 1315 2724 1319
rect 2718 1314 2724 1315
rect 3010 1319 3016 1320
rect 3010 1315 3011 1319
rect 3015 1315 3016 1319
rect 3010 1314 3016 1315
rect 3186 1319 3192 1320
rect 3186 1315 3187 1319
rect 3191 1315 3192 1319
rect 3186 1314 3192 1315
rect 2658 1299 2664 1300
rect 2658 1295 2659 1299
rect 2663 1295 2664 1299
rect 2658 1294 2664 1295
rect 2642 1291 2648 1292
rect 2642 1287 2643 1291
rect 2647 1287 2648 1291
rect 2642 1286 2648 1287
rect 2720 1284 2722 1314
rect 2750 1309 2756 1310
rect 2750 1305 2751 1309
rect 2755 1305 2756 1309
rect 2750 1304 2756 1305
rect 2934 1309 2940 1310
rect 2934 1305 2935 1309
rect 2939 1305 2940 1309
rect 2934 1304 2940 1305
rect 2718 1283 2724 1284
rect 2752 1283 2754 1304
rect 2936 1283 2938 1304
rect 3012 1292 3014 1314
rect 3110 1309 3116 1310
rect 3110 1305 3111 1309
rect 3115 1305 3116 1309
rect 3110 1304 3116 1305
rect 3010 1291 3016 1292
rect 3010 1287 3011 1291
rect 3015 1287 3016 1291
rect 3010 1286 3016 1287
rect 2982 1283 2988 1284
rect 3112 1283 3114 1304
rect 3188 1292 3190 1314
rect 3200 1300 3202 1394
rect 3270 1388 3276 1389
rect 3270 1384 3271 1388
rect 3275 1384 3276 1388
rect 3270 1383 3276 1384
rect 3438 1388 3444 1389
rect 3438 1384 3439 1388
rect 3443 1384 3444 1388
rect 3438 1383 3444 1384
rect 3272 1359 3274 1383
rect 3440 1359 3442 1383
rect 3271 1358 3275 1359
rect 3271 1353 3275 1354
rect 3279 1358 3283 1359
rect 3279 1353 3283 1354
rect 3439 1358 3443 1359
rect 3439 1353 3443 1354
rect 3447 1358 3451 1359
rect 3447 1353 3451 1354
rect 3280 1329 3282 1353
rect 3448 1329 3450 1353
rect 3278 1328 3284 1329
rect 3278 1324 3279 1328
rect 3283 1324 3284 1328
rect 3278 1323 3284 1324
rect 3446 1328 3452 1329
rect 3446 1324 3447 1328
rect 3451 1324 3452 1328
rect 3446 1323 3452 1324
rect 3524 1320 3526 1422
rect 3608 1408 3610 1429
rect 3784 1408 3786 1429
rect 3868 1428 3870 1474
rect 3942 1468 3948 1469
rect 3942 1464 3943 1468
rect 3947 1464 3948 1468
rect 3942 1463 3948 1464
rect 3944 1435 3946 1463
rect 3943 1434 3947 1435
rect 3943 1429 3947 1430
rect 3866 1427 3872 1428
rect 3866 1423 3867 1427
rect 3871 1423 3872 1427
rect 3866 1422 3872 1423
rect 3944 1409 3946 1429
rect 3942 1408 3948 1409
rect 3606 1407 3612 1408
rect 3606 1403 3607 1407
rect 3611 1403 3612 1407
rect 3606 1402 3612 1403
rect 3782 1407 3788 1408
rect 3782 1403 3783 1407
rect 3787 1403 3788 1407
rect 3942 1404 3943 1408
rect 3947 1404 3948 1408
rect 3942 1403 3948 1404
rect 3782 1402 3788 1403
rect 3858 1395 3864 1396
rect 3858 1391 3859 1395
rect 3863 1391 3864 1395
rect 3858 1390 3864 1391
rect 3942 1391 3948 1392
rect 3606 1388 3612 1389
rect 3606 1384 3607 1388
rect 3611 1384 3612 1388
rect 3606 1383 3612 1384
rect 3782 1388 3788 1389
rect 3782 1384 3783 1388
rect 3787 1384 3788 1388
rect 3782 1383 3788 1384
rect 3608 1359 3610 1383
rect 3784 1359 3786 1383
rect 3607 1358 3611 1359
rect 3607 1353 3611 1354
rect 3623 1358 3627 1359
rect 3623 1353 3627 1354
rect 3783 1358 3787 1359
rect 3783 1353 3787 1354
rect 3624 1329 3626 1353
rect 3622 1328 3628 1329
rect 3622 1324 3623 1328
rect 3627 1324 3628 1328
rect 3622 1323 3628 1324
rect 3354 1319 3360 1320
rect 3354 1315 3355 1319
rect 3359 1315 3360 1319
rect 3354 1314 3360 1315
rect 3522 1319 3528 1320
rect 3522 1315 3523 1319
rect 3527 1315 3528 1319
rect 3522 1314 3528 1315
rect 3278 1309 3284 1310
rect 3278 1305 3279 1309
rect 3283 1305 3284 1309
rect 3278 1304 3284 1305
rect 3198 1299 3204 1300
rect 3198 1295 3199 1299
rect 3203 1295 3204 1299
rect 3198 1294 3204 1295
rect 3186 1291 3192 1292
rect 3186 1287 3187 1291
rect 3191 1287 3192 1291
rect 3186 1286 3192 1287
rect 3280 1283 3282 1304
rect 2047 1282 2051 1283
rect 1543 1278 1547 1279
rect 1543 1273 1547 1274
rect 1655 1278 1659 1279
rect 1655 1273 1659 1274
rect 1719 1278 1723 1279
rect 1719 1273 1723 1274
rect 1863 1278 1867 1279
rect 1863 1273 1867 1274
rect 1895 1278 1899 1279
rect 1895 1273 1899 1274
rect 2007 1278 2011 1279
rect 2047 1277 2051 1278
rect 2071 1282 2075 1283
rect 2071 1277 2075 1278
rect 2151 1282 2155 1283
rect 2151 1277 2155 1278
rect 2207 1282 2211 1283
rect 2207 1277 2211 1278
rect 2287 1282 2291 1283
rect 2287 1277 2291 1278
rect 2383 1282 2387 1283
rect 2383 1277 2387 1278
rect 2431 1282 2435 1283
rect 2431 1277 2435 1278
rect 2567 1282 2571 1283
rect 2567 1277 2571 1278
rect 2583 1282 2587 1283
rect 2718 1279 2719 1283
rect 2723 1279 2724 1283
rect 2718 1278 2724 1279
rect 2743 1282 2747 1283
rect 2583 1277 2587 1278
rect 2743 1277 2747 1278
rect 2751 1282 2755 1283
rect 2751 1277 2755 1278
rect 2903 1282 2907 1283
rect 2903 1277 2907 1278
rect 2935 1282 2939 1283
rect 2935 1277 2939 1278
rect 2972 1281 2983 1283
rect 2007 1273 2011 1274
rect 1454 1271 1460 1272
rect 1454 1267 1455 1271
rect 1459 1267 1460 1271
rect 1454 1266 1460 1267
rect 1522 1271 1528 1272
rect 1522 1267 1523 1271
rect 1527 1267 1528 1271
rect 1522 1266 1528 1267
rect 1366 1251 1372 1252
rect 1366 1247 1367 1251
rect 1371 1247 1372 1251
rect 1366 1246 1372 1247
rect 1456 1244 1458 1266
rect 1544 1252 1546 1273
rect 1720 1252 1722 1273
rect 1770 1271 1776 1272
rect 1770 1267 1771 1271
rect 1775 1267 1776 1271
rect 1770 1266 1776 1267
rect 1794 1271 1800 1272
rect 1794 1267 1795 1271
rect 1799 1267 1800 1271
rect 1794 1266 1800 1267
rect 1542 1251 1548 1252
rect 1542 1247 1543 1251
rect 1547 1247 1548 1251
rect 1542 1246 1548 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 1718 1246 1724 1247
rect 770 1243 776 1244
rect 770 1239 771 1243
rect 775 1239 776 1243
rect 770 1238 776 1239
rect 930 1243 936 1244
rect 930 1239 931 1243
rect 935 1239 936 1243
rect 930 1238 936 1239
rect 978 1243 984 1244
rect 978 1239 979 1243
rect 983 1239 984 1243
rect 1274 1243 1280 1244
rect 978 1238 984 1239
rect 1266 1239 1272 1240
rect 1266 1235 1267 1239
rect 1271 1235 1272 1239
rect 1274 1239 1275 1243
rect 1279 1239 1280 1243
rect 1274 1238 1280 1239
rect 1454 1243 1460 1244
rect 1454 1239 1455 1243
rect 1459 1239 1460 1243
rect 1454 1238 1460 1239
rect 1266 1234 1272 1235
rect 694 1232 700 1233
rect 694 1228 695 1232
rect 699 1228 700 1232
rect 694 1227 700 1228
rect 854 1232 860 1233
rect 854 1228 855 1232
rect 859 1228 860 1232
rect 854 1227 860 1228
rect 1022 1232 1028 1233
rect 1022 1228 1023 1232
rect 1027 1228 1028 1232
rect 1022 1227 1028 1228
rect 1190 1232 1196 1233
rect 1190 1228 1191 1232
rect 1195 1228 1196 1232
rect 1190 1227 1196 1228
rect 696 1203 698 1227
rect 856 1203 858 1227
rect 1024 1203 1026 1227
rect 1192 1203 1194 1227
rect 695 1202 699 1203
rect 695 1197 699 1198
rect 759 1202 763 1203
rect 759 1197 763 1198
rect 855 1202 859 1203
rect 855 1197 859 1198
rect 927 1202 931 1203
rect 927 1197 931 1198
rect 1023 1202 1027 1203
rect 1023 1197 1027 1198
rect 1095 1202 1099 1203
rect 1095 1197 1099 1198
rect 1191 1202 1195 1203
rect 1191 1197 1195 1198
rect 1247 1202 1251 1203
rect 1247 1197 1251 1198
rect 760 1173 762 1197
rect 928 1173 930 1197
rect 1096 1173 1098 1197
rect 1248 1173 1250 1197
rect 758 1172 764 1173
rect 758 1168 759 1172
rect 763 1168 764 1172
rect 758 1167 764 1168
rect 926 1172 932 1173
rect 926 1168 927 1172
rect 931 1168 932 1172
rect 926 1167 932 1168
rect 1094 1172 1100 1173
rect 1094 1168 1095 1172
rect 1099 1168 1100 1172
rect 1094 1167 1100 1168
rect 1246 1172 1252 1173
rect 1246 1168 1247 1172
rect 1251 1168 1252 1172
rect 1246 1167 1252 1168
rect 498 1163 504 1164
rect 498 1159 499 1163
rect 503 1159 504 1163
rect 498 1158 504 1159
rect 674 1163 680 1164
rect 674 1159 675 1163
rect 679 1159 680 1163
rect 674 1158 680 1159
rect 718 1163 724 1164
rect 718 1159 719 1163
rect 723 1159 724 1163
rect 718 1158 724 1159
rect 878 1163 884 1164
rect 878 1159 879 1163
rect 883 1159 884 1163
rect 878 1158 884 1159
rect 422 1153 428 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 422 1149 423 1153
rect 427 1149 428 1153
rect 422 1148 428 1149
rect 110 1147 116 1148
rect 112 1123 114 1147
rect 424 1123 426 1148
rect 500 1136 502 1158
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 498 1135 504 1136
rect 450 1131 456 1132
rect 450 1127 451 1131
rect 455 1127 456 1131
rect 498 1131 499 1135
rect 503 1131 504 1135
rect 498 1130 504 1131
rect 450 1126 456 1127
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 423 1122 427 1123
rect 423 1117 427 1118
rect 112 1097 114 1117
rect 110 1096 116 1097
rect 376 1096 378 1117
rect 386 1115 392 1116
rect 386 1111 387 1115
rect 391 1111 392 1115
rect 386 1110 392 1111
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 110 1074 116 1075
rect 374 1076 380 1077
rect 112 1047 114 1074
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 376 1047 378 1071
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 303 1046 307 1047
rect 303 1041 307 1042
rect 375 1046 379 1047
rect 375 1041 379 1042
rect 112 1014 114 1041
rect 304 1017 306 1041
rect 302 1016 308 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 302 1012 303 1016
rect 307 1012 308 1016
rect 302 1011 308 1012
rect 110 1008 116 1009
rect 388 1008 390 1110
rect 452 1088 454 1126
rect 592 1123 594 1148
rect 720 1124 722 1158
rect 758 1153 764 1154
rect 758 1149 759 1153
rect 763 1149 764 1153
rect 758 1148 764 1149
rect 718 1123 724 1124
rect 760 1123 762 1148
rect 880 1136 882 1158
rect 926 1153 932 1154
rect 926 1149 927 1153
rect 931 1149 932 1153
rect 926 1148 932 1149
rect 1094 1153 1100 1154
rect 1094 1149 1095 1153
rect 1099 1149 1100 1153
rect 1094 1148 1100 1149
rect 1246 1153 1252 1154
rect 1246 1149 1247 1153
rect 1251 1149 1252 1153
rect 1246 1148 1252 1149
rect 878 1135 884 1136
rect 878 1131 879 1135
rect 883 1131 884 1135
rect 878 1130 884 1131
rect 928 1123 930 1148
rect 1096 1123 1098 1148
rect 1194 1131 1200 1132
rect 1194 1127 1195 1131
rect 1199 1127 1200 1131
rect 1194 1126 1200 1127
rect 487 1122 491 1123
rect 487 1117 491 1118
rect 591 1122 595 1123
rect 591 1117 595 1118
rect 599 1122 603 1123
rect 599 1117 603 1118
rect 711 1122 715 1123
rect 718 1119 719 1123
rect 723 1119 724 1123
rect 718 1118 724 1119
rect 759 1122 763 1123
rect 711 1117 715 1118
rect 759 1117 763 1118
rect 831 1122 835 1123
rect 831 1117 835 1118
rect 927 1122 931 1123
rect 927 1117 931 1118
rect 967 1122 971 1123
rect 967 1117 971 1118
rect 1095 1122 1099 1123
rect 1095 1117 1099 1118
rect 1119 1122 1123 1123
rect 1119 1117 1123 1118
rect 488 1096 490 1117
rect 562 1115 568 1116
rect 562 1111 563 1115
rect 567 1111 568 1115
rect 562 1110 568 1111
rect 486 1095 492 1096
rect 486 1091 487 1095
rect 491 1091 492 1095
rect 486 1090 492 1091
rect 564 1088 566 1110
rect 600 1096 602 1117
rect 674 1115 680 1116
rect 674 1111 675 1115
rect 679 1111 680 1115
rect 674 1110 680 1111
rect 598 1095 604 1096
rect 598 1091 599 1095
rect 603 1091 604 1095
rect 598 1090 604 1091
rect 676 1088 678 1110
rect 712 1096 714 1117
rect 832 1096 834 1117
rect 906 1115 912 1116
rect 906 1111 907 1115
rect 911 1111 912 1115
rect 906 1110 912 1111
rect 710 1095 716 1096
rect 710 1091 711 1095
rect 715 1091 716 1095
rect 710 1090 716 1091
rect 830 1095 836 1096
rect 830 1091 831 1095
rect 835 1091 836 1095
rect 830 1090 836 1091
rect 908 1088 910 1110
rect 968 1096 970 1117
rect 1042 1115 1048 1116
rect 1042 1111 1043 1115
rect 1047 1111 1048 1115
rect 1042 1110 1048 1111
rect 966 1095 972 1096
rect 966 1091 967 1095
rect 971 1091 972 1095
rect 966 1090 972 1091
rect 1044 1088 1046 1110
rect 1120 1096 1122 1117
rect 1118 1095 1124 1096
rect 1118 1091 1119 1095
rect 1123 1091 1124 1095
rect 1118 1090 1124 1091
rect 1196 1088 1198 1126
rect 1248 1123 1250 1148
rect 1268 1136 1270 1234
rect 1366 1232 1372 1233
rect 1366 1228 1367 1232
rect 1371 1228 1372 1232
rect 1366 1227 1372 1228
rect 1542 1232 1548 1233
rect 1542 1228 1543 1232
rect 1547 1228 1548 1232
rect 1542 1227 1548 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 1718 1227 1724 1228
rect 1368 1203 1370 1227
rect 1544 1203 1546 1227
rect 1720 1203 1722 1227
rect 1367 1202 1371 1203
rect 1367 1197 1371 1198
rect 1399 1202 1403 1203
rect 1399 1197 1403 1198
rect 1543 1202 1547 1203
rect 1543 1197 1547 1198
rect 1687 1202 1691 1203
rect 1687 1197 1691 1198
rect 1719 1202 1723 1203
rect 1719 1197 1723 1198
rect 1400 1173 1402 1197
rect 1544 1173 1546 1197
rect 1688 1173 1690 1197
rect 1398 1172 1404 1173
rect 1398 1168 1399 1172
rect 1403 1168 1404 1172
rect 1398 1167 1404 1168
rect 1542 1172 1548 1173
rect 1542 1168 1543 1172
rect 1547 1168 1548 1172
rect 1542 1167 1548 1168
rect 1686 1172 1692 1173
rect 1686 1168 1687 1172
rect 1691 1168 1692 1172
rect 1686 1167 1692 1168
rect 1772 1164 1774 1266
rect 1796 1244 1798 1266
rect 1896 1252 1898 1273
rect 2008 1253 2010 1273
rect 2048 1257 2050 1277
rect 2046 1256 2052 1257
rect 2152 1256 2154 1277
rect 2226 1275 2232 1276
rect 2226 1271 2227 1275
rect 2231 1271 2232 1275
rect 2226 1270 2232 1271
rect 2006 1252 2012 1253
rect 1894 1251 1900 1252
rect 1894 1247 1895 1251
rect 1899 1247 1900 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2046 1252 2047 1256
rect 2051 1252 2052 1256
rect 2046 1251 2052 1252
rect 2150 1255 2156 1256
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2228 1248 2230 1270
rect 2288 1256 2290 1277
rect 2362 1275 2368 1276
rect 2362 1271 2363 1275
rect 2367 1271 2368 1275
rect 2362 1270 2368 1271
rect 2286 1255 2292 1256
rect 2286 1251 2287 1255
rect 2291 1251 2292 1255
rect 2286 1250 2292 1251
rect 2364 1248 2366 1270
rect 2432 1256 2434 1277
rect 2506 1275 2512 1276
rect 2506 1271 2507 1275
rect 2511 1271 2512 1275
rect 2506 1270 2512 1271
rect 2430 1255 2436 1256
rect 2430 1251 2431 1255
rect 2435 1251 2436 1255
rect 2430 1250 2436 1251
rect 2508 1248 2510 1270
rect 2584 1256 2586 1277
rect 2658 1275 2664 1276
rect 2658 1271 2659 1275
rect 2663 1271 2664 1275
rect 2658 1270 2664 1271
rect 2582 1255 2588 1256
rect 2582 1251 2583 1255
rect 2587 1251 2588 1255
rect 2582 1250 2588 1251
rect 2660 1248 2662 1270
rect 2744 1256 2746 1277
rect 2904 1256 2906 1277
rect 2972 1276 2974 1281
rect 2982 1279 2983 1281
rect 2987 1279 2988 1283
rect 2982 1278 2988 1279
rect 3071 1282 3075 1283
rect 3071 1277 3075 1278
rect 3111 1282 3115 1283
rect 3111 1277 3115 1278
rect 3247 1282 3251 1283
rect 3247 1277 3251 1278
rect 3279 1282 3283 1283
rect 3279 1277 3283 1278
rect 2970 1275 2976 1276
rect 2970 1271 2971 1275
rect 2975 1271 2976 1275
rect 2970 1270 2976 1271
rect 2978 1275 2984 1276
rect 2978 1271 2979 1275
rect 2983 1271 2984 1275
rect 2978 1270 2984 1271
rect 2742 1255 2748 1256
rect 2742 1251 2743 1255
rect 2747 1251 2748 1255
rect 2742 1250 2748 1251
rect 2902 1255 2908 1256
rect 2902 1251 2903 1255
rect 2907 1251 2908 1255
rect 2902 1250 2908 1251
rect 2980 1248 2982 1270
rect 3072 1256 3074 1277
rect 3248 1256 3250 1277
rect 3356 1276 3358 1314
rect 3446 1309 3452 1310
rect 3446 1305 3447 1309
rect 3451 1305 3452 1309
rect 3446 1304 3452 1305
rect 3622 1309 3628 1310
rect 3622 1305 3623 1309
rect 3627 1305 3628 1309
rect 3622 1304 3628 1305
rect 3448 1283 3450 1304
rect 3624 1283 3626 1304
rect 3690 1287 3696 1288
rect 3690 1283 3691 1287
rect 3695 1283 3696 1287
rect 3431 1282 3435 1283
rect 3431 1277 3435 1278
rect 3447 1282 3451 1283
rect 3447 1277 3451 1278
rect 3615 1282 3619 1283
rect 3615 1277 3619 1278
rect 3623 1282 3627 1283
rect 3690 1282 3696 1283
rect 3807 1282 3811 1283
rect 3623 1277 3627 1278
rect 3330 1275 3336 1276
rect 3330 1271 3331 1275
rect 3335 1271 3336 1275
rect 3330 1270 3336 1271
rect 3354 1275 3360 1276
rect 3354 1271 3355 1275
rect 3359 1271 3360 1275
rect 3354 1270 3360 1271
rect 3070 1255 3076 1256
rect 3070 1251 3071 1255
rect 3075 1251 3076 1255
rect 3070 1250 3076 1251
rect 3246 1255 3252 1256
rect 3246 1251 3247 1255
rect 3251 1251 3252 1255
rect 3246 1250 3252 1251
rect 3332 1248 3334 1270
rect 3432 1256 3434 1277
rect 3616 1256 3618 1277
rect 3430 1255 3436 1256
rect 3430 1251 3431 1255
rect 3435 1251 3436 1255
rect 3430 1250 3436 1251
rect 3614 1255 3620 1256
rect 3614 1251 3615 1255
rect 3619 1251 3620 1255
rect 3614 1250 3620 1251
rect 3692 1248 3694 1282
rect 3807 1277 3811 1278
rect 3698 1275 3704 1276
rect 3698 1271 3699 1275
rect 3703 1271 3704 1275
rect 3698 1270 3704 1271
rect 2006 1247 2012 1248
rect 2226 1247 2232 1248
rect 1894 1246 1900 1247
rect 1794 1243 1800 1244
rect 1794 1239 1795 1243
rect 1799 1239 1800 1243
rect 2226 1243 2227 1247
rect 2231 1243 2232 1247
rect 2226 1242 2232 1243
rect 2362 1247 2368 1248
rect 2362 1243 2363 1247
rect 2367 1243 2368 1247
rect 2362 1242 2368 1243
rect 2506 1247 2512 1248
rect 2506 1243 2507 1247
rect 2511 1243 2512 1247
rect 2506 1242 2512 1243
rect 2658 1247 2664 1248
rect 2658 1243 2659 1247
rect 2663 1243 2664 1247
rect 2658 1242 2664 1243
rect 2666 1247 2672 1248
rect 2666 1243 2667 1247
rect 2671 1243 2672 1247
rect 2666 1242 2672 1243
rect 2978 1247 2984 1248
rect 2978 1243 2979 1247
rect 2983 1243 2984 1247
rect 2978 1242 2984 1243
rect 3330 1247 3336 1248
rect 3330 1243 3331 1247
rect 3335 1243 3336 1247
rect 3330 1242 3336 1243
rect 3690 1247 3696 1248
rect 3690 1243 3691 1247
rect 3695 1243 3696 1247
rect 3690 1242 3696 1243
rect 1794 1238 1800 1239
rect 2046 1239 2052 1240
rect 2006 1235 2012 1236
rect 1894 1232 1900 1233
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2046 1235 2047 1239
rect 2051 1235 2052 1239
rect 2046 1234 2052 1235
rect 2150 1236 2156 1237
rect 2006 1230 2012 1231
rect 1894 1227 1900 1228
rect 1896 1203 1898 1227
rect 2008 1203 2010 1230
rect 2048 1207 2050 1234
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2286 1236 2292 1237
rect 2286 1232 2287 1236
rect 2291 1232 2292 1236
rect 2286 1231 2292 1232
rect 2430 1236 2436 1237
rect 2430 1232 2431 1236
rect 2435 1232 2436 1236
rect 2430 1231 2436 1232
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 2582 1231 2588 1232
rect 2152 1207 2154 1231
rect 2288 1207 2290 1231
rect 2350 1215 2356 1216
rect 2350 1211 2351 1215
rect 2355 1211 2356 1215
rect 2350 1210 2356 1211
rect 2047 1206 2051 1207
rect 1839 1202 1843 1203
rect 1839 1197 1843 1198
rect 1895 1202 1899 1203
rect 1895 1197 1899 1198
rect 2007 1202 2011 1203
rect 2047 1201 2051 1202
rect 2151 1206 2155 1207
rect 2151 1201 2155 1202
rect 2287 1206 2291 1207
rect 2287 1201 2291 1202
rect 2311 1206 2315 1207
rect 2311 1201 2315 1202
rect 2007 1197 2011 1198
rect 1840 1173 1842 1197
rect 1838 1172 1844 1173
rect 1838 1168 1839 1172
rect 1843 1168 1844 1172
rect 2008 1170 2010 1197
rect 2048 1174 2050 1201
rect 2312 1177 2314 1201
rect 2310 1176 2316 1177
rect 2046 1173 2052 1174
rect 1838 1167 1844 1168
rect 2006 1169 2012 1170
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2046 1169 2047 1173
rect 2051 1169 2052 1173
rect 2310 1172 2311 1176
rect 2315 1172 2316 1176
rect 2310 1171 2316 1172
rect 2046 1168 2052 1169
rect 2006 1164 2012 1165
rect 1322 1163 1328 1164
rect 1322 1159 1323 1163
rect 1327 1159 1328 1163
rect 1322 1158 1328 1159
rect 1618 1163 1624 1164
rect 1618 1159 1619 1163
rect 1623 1159 1624 1163
rect 1618 1158 1624 1159
rect 1762 1163 1768 1164
rect 1762 1159 1763 1163
rect 1767 1159 1768 1163
rect 1762 1158 1768 1159
rect 1770 1163 1776 1164
rect 1770 1159 1771 1163
rect 1775 1159 1776 1163
rect 1770 1158 1776 1159
rect 1324 1136 1326 1158
rect 1398 1153 1404 1154
rect 1398 1149 1399 1153
rect 1403 1149 1404 1153
rect 1398 1148 1404 1149
rect 1542 1153 1548 1154
rect 1542 1149 1543 1153
rect 1547 1149 1548 1153
rect 1542 1148 1548 1149
rect 1266 1135 1272 1136
rect 1266 1131 1267 1135
rect 1271 1131 1272 1135
rect 1266 1130 1272 1131
rect 1322 1135 1328 1136
rect 1322 1131 1323 1135
rect 1327 1131 1328 1135
rect 1322 1130 1328 1131
rect 1400 1123 1402 1148
rect 1544 1123 1546 1148
rect 1620 1136 1622 1158
rect 1686 1153 1692 1154
rect 1686 1149 1687 1153
rect 1691 1149 1692 1153
rect 1686 1148 1692 1149
rect 1618 1135 1624 1136
rect 1582 1131 1588 1132
rect 1582 1127 1583 1131
rect 1587 1127 1588 1131
rect 1618 1131 1619 1135
rect 1623 1131 1624 1135
rect 1618 1130 1624 1131
rect 1582 1126 1588 1127
rect 1247 1122 1251 1123
rect 1247 1117 1251 1118
rect 1279 1122 1283 1123
rect 1279 1117 1283 1118
rect 1399 1122 1403 1123
rect 1399 1117 1403 1118
rect 1447 1122 1451 1123
rect 1447 1117 1451 1118
rect 1543 1122 1547 1123
rect 1543 1117 1547 1118
rect 1238 1107 1244 1108
rect 1238 1103 1239 1107
rect 1243 1103 1244 1107
rect 1238 1102 1244 1103
rect 1240 1088 1242 1102
rect 1280 1096 1282 1117
rect 1362 1115 1368 1116
rect 1362 1111 1363 1115
rect 1367 1111 1368 1115
rect 1362 1110 1368 1111
rect 1278 1095 1284 1096
rect 1278 1091 1279 1095
rect 1283 1091 1284 1095
rect 1278 1090 1284 1091
rect 1364 1088 1366 1110
rect 1448 1096 1450 1117
rect 1498 1115 1504 1116
rect 1498 1111 1499 1115
rect 1503 1111 1504 1115
rect 1498 1110 1504 1111
rect 1446 1095 1452 1096
rect 1446 1091 1447 1095
rect 1451 1091 1452 1095
rect 1446 1090 1452 1091
rect 450 1087 456 1088
rect 450 1083 451 1087
rect 455 1083 456 1087
rect 450 1082 456 1083
rect 562 1087 568 1088
rect 562 1083 563 1087
rect 567 1083 568 1087
rect 562 1082 568 1083
rect 674 1087 680 1088
rect 674 1083 675 1087
rect 679 1083 680 1087
rect 906 1087 912 1088
rect 674 1082 680 1083
rect 786 1083 792 1084
rect 786 1079 787 1083
rect 791 1079 792 1083
rect 906 1083 907 1087
rect 911 1083 912 1087
rect 906 1082 912 1083
rect 1042 1087 1048 1088
rect 1042 1083 1043 1087
rect 1047 1083 1048 1087
rect 1042 1082 1048 1083
rect 1194 1087 1200 1088
rect 1194 1083 1195 1087
rect 1199 1083 1200 1087
rect 1194 1082 1200 1083
rect 1238 1087 1244 1088
rect 1238 1083 1239 1087
rect 1243 1083 1244 1087
rect 1238 1082 1244 1083
rect 1362 1087 1368 1088
rect 1362 1083 1363 1087
rect 1367 1083 1368 1087
rect 1362 1082 1368 1083
rect 786 1078 792 1079
rect 486 1076 492 1077
rect 486 1072 487 1076
rect 491 1072 492 1076
rect 486 1071 492 1072
rect 598 1076 604 1077
rect 598 1072 599 1076
rect 603 1072 604 1076
rect 598 1071 604 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 488 1047 490 1071
rect 600 1047 602 1071
rect 712 1047 714 1071
rect 447 1046 451 1047
rect 447 1041 451 1042
rect 487 1046 491 1047
rect 487 1041 491 1042
rect 591 1046 595 1047
rect 591 1041 595 1042
rect 599 1046 603 1047
rect 599 1041 603 1042
rect 711 1046 715 1047
rect 711 1041 715 1042
rect 727 1046 731 1047
rect 727 1041 731 1042
rect 448 1017 450 1041
rect 592 1017 594 1041
rect 728 1017 730 1041
rect 446 1016 452 1017
rect 446 1012 447 1016
rect 451 1012 452 1016
rect 446 1011 452 1012
rect 590 1016 596 1017
rect 590 1012 591 1016
rect 595 1012 596 1016
rect 590 1011 596 1012
rect 726 1016 732 1017
rect 726 1012 727 1016
rect 731 1012 732 1016
rect 726 1011 732 1012
rect 386 1007 392 1008
rect 386 1003 387 1007
rect 391 1003 392 1007
rect 386 1002 392 1003
rect 394 1007 400 1008
rect 394 1003 395 1007
rect 399 1003 400 1007
rect 394 1002 400 1003
rect 666 1007 672 1008
rect 666 1003 667 1007
rect 671 1003 672 1007
rect 666 1002 672 1003
rect 302 997 308 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 302 993 303 997
rect 307 993 308 997
rect 302 992 308 993
rect 110 991 116 992
rect 112 971 114 991
rect 304 971 306 992
rect 396 980 398 1002
rect 446 997 452 998
rect 446 993 447 997
rect 451 993 452 997
rect 446 992 452 993
rect 590 997 596 998
rect 590 993 591 997
rect 595 993 596 997
rect 590 992 596 993
rect 394 979 400 980
rect 394 975 395 979
rect 399 975 400 979
rect 394 974 400 975
rect 448 971 450 992
rect 522 975 528 976
rect 522 971 523 975
rect 527 971 528 975
rect 592 971 594 992
rect 111 970 115 971
rect 111 965 115 966
rect 255 970 259 971
rect 255 965 259 966
rect 303 970 307 971
rect 303 965 307 966
rect 447 970 451 971
rect 522 970 528 971
rect 591 970 595 971
rect 447 965 451 966
rect 112 945 114 965
rect 110 944 116 945
rect 256 944 258 965
rect 322 963 328 964
rect 322 959 323 963
rect 327 959 328 963
rect 322 958 328 959
rect 330 963 336 964
rect 330 959 331 963
rect 335 959 336 963
rect 330 958 336 959
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 254 943 260 944
rect 254 939 255 943
rect 259 939 260 943
rect 254 938 260 939
rect 110 927 116 928
rect 110 923 111 927
rect 115 923 116 927
rect 110 922 116 923
rect 254 924 260 925
rect 112 891 114 922
rect 254 920 255 924
rect 259 920 260 924
rect 254 919 260 920
rect 256 891 258 919
rect 111 890 115 891
rect 111 885 115 886
rect 255 890 259 891
rect 255 885 259 886
rect 112 858 114 885
rect 256 861 258 885
rect 254 860 260 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 254 856 255 860
rect 259 856 260 860
rect 254 855 260 856
rect 110 852 116 853
rect 324 852 326 958
rect 332 936 334 958
rect 448 944 450 965
rect 446 943 452 944
rect 446 939 447 943
rect 451 939 452 943
rect 446 938 452 939
rect 524 936 526 970
rect 591 965 595 966
rect 631 970 635 971
rect 631 965 635 966
rect 632 944 634 965
rect 668 964 670 1002
rect 726 997 732 998
rect 726 993 727 997
rect 731 993 732 997
rect 726 992 732 993
rect 728 971 730 992
rect 788 980 790 1078
rect 830 1076 836 1077
rect 830 1072 831 1076
rect 835 1072 836 1076
rect 830 1071 836 1072
rect 966 1076 972 1077
rect 966 1072 967 1076
rect 971 1072 972 1076
rect 966 1071 972 1072
rect 1118 1076 1124 1077
rect 1118 1072 1119 1076
rect 1123 1072 1124 1076
rect 1118 1071 1124 1072
rect 1278 1076 1284 1077
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 1446 1076 1452 1077
rect 1446 1072 1447 1076
rect 1451 1072 1452 1076
rect 1446 1071 1452 1072
rect 832 1047 834 1071
rect 968 1047 970 1071
rect 1120 1047 1122 1071
rect 1280 1047 1282 1071
rect 1448 1047 1450 1071
rect 831 1046 835 1047
rect 831 1041 835 1042
rect 855 1046 859 1047
rect 855 1041 859 1042
rect 967 1046 971 1047
rect 967 1041 971 1042
rect 975 1046 979 1047
rect 975 1041 979 1042
rect 1087 1046 1091 1047
rect 1087 1041 1091 1042
rect 1119 1046 1123 1047
rect 1119 1041 1123 1042
rect 1199 1046 1203 1047
rect 1199 1041 1203 1042
rect 1279 1046 1283 1047
rect 1279 1041 1283 1042
rect 1311 1046 1315 1047
rect 1311 1041 1315 1042
rect 1431 1046 1435 1047
rect 1431 1041 1435 1042
rect 1447 1046 1451 1047
rect 1447 1041 1451 1042
rect 856 1017 858 1041
rect 976 1017 978 1041
rect 1088 1017 1090 1041
rect 1200 1017 1202 1041
rect 1312 1017 1314 1041
rect 1432 1017 1434 1041
rect 854 1016 860 1017
rect 854 1012 855 1016
rect 859 1012 860 1016
rect 854 1011 860 1012
rect 974 1016 980 1017
rect 974 1012 975 1016
rect 979 1012 980 1016
rect 974 1011 980 1012
rect 1086 1016 1092 1017
rect 1086 1012 1087 1016
rect 1091 1012 1092 1016
rect 1086 1011 1092 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1310 1016 1316 1017
rect 1310 1012 1311 1016
rect 1315 1012 1316 1016
rect 1310 1011 1316 1012
rect 1430 1016 1436 1017
rect 1430 1012 1431 1016
rect 1435 1012 1436 1016
rect 1430 1011 1436 1012
rect 1500 1008 1502 1110
rect 1584 1088 1586 1126
rect 1688 1123 1690 1148
rect 1764 1136 1766 1158
rect 2310 1157 2316 1158
rect 2046 1156 2052 1157
rect 1838 1153 1844 1154
rect 1838 1149 1839 1153
rect 1843 1149 1844 1153
rect 1838 1148 1844 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2046 1152 2047 1156
rect 2051 1152 2052 1156
rect 2310 1153 2311 1157
rect 2315 1153 2316 1157
rect 2310 1152 2316 1153
rect 2046 1151 2052 1152
rect 1762 1135 1768 1136
rect 1762 1131 1763 1135
rect 1767 1131 1768 1135
rect 1762 1130 1768 1131
rect 1840 1123 1842 1148
rect 2006 1147 2012 1148
rect 2008 1123 2010 1147
rect 2048 1127 2050 1151
rect 2312 1127 2314 1152
rect 2352 1140 2354 1210
rect 2432 1207 2434 1231
rect 2584 1207 2586 1231
rect 2668 1216 2670 1242
rect 2742 1236 2748 1237
rect 2742 1232 2743 1236
rect 2747 1232 2748 1236
rect 2742 1231 2748 1232
rect 2902 1236 2908 1237
rect 2902 1232 2903 1236
rect 2907 1232 2908 1236
rect 2902 1231 2908 1232
rect 3070 1236 3076 1237
rect 3070 1232 3071 1236
rect 3075 1232 3076 1236
rect 3070 1231 3076 1232
rect 3246 1236 3252 1237
rect 3246 1232 3247 1236
rect 3251 1232 3252 1236
rect 3246 1231 3252 1232
rect 3430 1236 3436 1237
rect 3430 1232 3431 1236
rect 3435 1232 3436 1236
rect 3430 1231 3436 1232
rect 3614 1236 3620 1237
rect 3614 1232 3615 1236
rect 3619 1232 3620 1236
rect 3614 1231 3620 1232
rect 2666 1215 2672 1216
rect 2666 1211 2667 1215
rect 2671 1211 2672 1215
rect 2666 1210 2672 1211
rect 2744 1207 2746 1231
rect 2904 1207 2906 1231
rect 3072 1207 3074 1231
rect 3248 1207 3250 1231
rect 3432 1207 3434 1231
rect 3616 1207 3618 1231
rect 2415 1206 2419 1207
rect 2415 1201 2419 1202
rect 2431 1206 2435 1207
rect 2431 1201 2435 1202
rect 2527 1206 2531 1207
rect 2527 1201 2531 1202
rect 2583 1206 2587 1207
rect 2583 1201 2587 1202
rect 2639 1206 2643 1207
rect 2639 1201 2643 1202
rect 2743 1206 2747 1207
rect 2743 1201 2747 1202
rect 2767 1206 2771 1207
rect 2767 1201 2771 1202
rect 2903 1206 2907 1207
rect 2903 1201 2907 1202
rect 2911 1206 2915 1207
rect 2911 1201 2915 1202
rect 3071 1206 3075 1207
rect 3071 1201 3075 1202
rect 3247 1206 3251 1207
rect 3247 1201 3251 1202
rect 3431 1206 3435 1207
rect 3431 1201 3435 1202
rect 3439 1206 3443 1207
rect 3439 1201 3443 1202
rect 3615 1206 3619 1207
rect 3615 1201 3619 1202
rect 3631 1206 3635 1207
rect 3631 1201 3635 1202
rect 2416 1177 2418 1201
rect 2528 1177 2530 1201
rect 2640 1177 2642 1201
rect 2768 1177 2770 1201
rect 2912 1177 2914 1201
rect 3072 1177 3074 1201
rect 3248 1177 3250 1201
rect 3440 1177 3442 1201
rect 3632 1177 3634 1201
rect 2414 1176 2420 1177
rect 2414 1172 2415 1176
rect 2419 1172 2420 1176
rect 2414 1171 2420 1172
rect 2526 1176 2532 1177
rect 2526 1172 2527 1176
rect 2531 1172 2532 1176
rect 2526 1171 2532 1172
rect 2638 1176 2644 1177
rect 2638 1172 2639 1176
rect 2643 1172 2644 1176
rect 2638 1171 2644 1172
rect 2766 1176 2772 1177
rect 2766 1172 2767 1176
rect 2771 1172 2772 1176
rect 2766 1171 2772 1172
rect 2910 1176 2916 1177
rect 2910 1172 2911 1176
rect 2915 1172 2916 1176
rect 2910 1171 2916 1172
rect 3070 1176 3076 1177
rect 3070 1172 3071 1176
rect 3075 1172 3076 1176
rect 3070 1171 3076 1172
rect 3246 1176 3252 1177
rect 3246 1172 3247 1176
rect 3251 1172 3252 1176
rect 3246 1171 3252 1172
rect 3438 1176 3444 1177
rect 3438 1172 3439 1176
rect 3443 1172 3444 1176
rect 3438 1171 3444 1172
rect 3630 1176 3636 1177
rect 3630 1172 3631 1176
rect 3635 1172 3636 1176
rect 3630 1171 3636 1172
rect 3700 1168 3702 1270
rect 3808 1256 3810 1277
rect 3860 1276 3862 1390
rect 3942 1387 3943 1391
rect 3947 1387 3948 1391
rect 3942 1386 3948 1387
rect 3944 1359 3946 1386
rect 3943 1358 3947 1359
rect 3943 1353 3947 1354
rect 3944 1326 3946 1353
rect 3942 1325 3948 1326
rect 3942 1321 3943 1325
rect 3947 1321 3948 1325
rect 3942 1320 3948 1321
rect 3942 1308 3948 1309
rect 3942 1304 3943 1308
rect 3947 1304 3948 1308
rect 3942 1303 3948 1304
rect 3944 1283 3946 1303
rect 3943 1282 3947 1283
rect 3943 1277 3947 1278
rect 3858 1275 3864 1276
rect 3858 1271 3859 1275
rect 3863 1271 3864 1275
rect 3858 1270 3864 1271
rect 3944 1257 3946 1277
rect 3942 1256 3948 1257
rect 3806 1255 3812 1256
rect 3806 1251 3807 1255
rect 3811 1251 3812 1255
rect 3942 1252 3943 1256
rect 3947 1252 3948 1256
rect 3942 1251 3948 1252
rect 3806 1250 3812 1251
rect 3882 1243 3888 1244
rect 3882 1239 3883 1243
rect 3887 1239 3888 1243
rect 3882 1238 3888 1239
rect 3942 1239 3948 1240
rect 3806 1236 3812 1237
rect 3806 1232 3807 1236
rect 3811 1232 3812 1236
rect 3806 1231 3812 1232
rect 3808 1207 3810 1231
rect 3807 1206 3811 1207
rect 3807 1201 3811 1202
rect 3831 1206 3835 1207
rect 3831 1201 3835 1202
rect 3832 1177 3834 1201
rect 3830 1176 3836 1177
rect 3830 1172 3831 1176
rect 3835 1172 3836 1176
rect 3830 1171 3836 1172
rect 2386 1167 2392 1168
rect 2386 1163 2387 1167
rect 2391 1163 2392 1167
rect 2386 1162 2392 1163
rect 2490 1167 2496 1168
rect 2490 1163 2491 1167
rect 2495 1163 2496 1167
rect 2490 1162 2496 1163
rect 2602 1167 2608 1168
rect 2602 1163 2603 1167
rect 2607 1163 2608 1167
rect 2602 1162 2608 1163
rect 2714 1167 2720 1168
rect 2714 1163 2715 1167
rect 2719 1163 2720 1167
rect 2714 1162 2720 1163
rect 2722 1167 2728 1168
rect 2722 1163 2723 1167
rect 2727 1163 2728 1167
rect 2722 1162 2728 1163
rect 2986 1167 2992 1168
rect 2986 1163 2987 1167
rect 2991 1163 2992 1167
rect 2986 1162 2992 1163
rect 3138 1167 3144 1168
rect 3138 1163 3139 1167
rect 3143 1163 3144 1167
rect 3138 1162 3144 1163
rect 3322 1167 3328 1168
rect 3322 1163 3323 1167
rect 3327 1163 3328 1167
rect 3322 1162 3328 1163
rect 3378 1167 3384 1168
rect 3378 1163 3379 1167
rect 3383 1163 3384 1167
rect 3378 1162 3384 1163
rect 3698 1167 3704 1168
rect 3698 1163 3699 1167
rect 3703 1163 3704 1167
rect 3698 1162 3704 1163
rect 2388 1140 2390 1162
rect 2414 1157 2420 1158
rect 2414 1153 2415 1157
rect 2419 1153 2420 1157
rect 2414 1152 2420 1153
rect 2350 1139 2356 1140
rect 2350 1135 2351 1139
rect 2355 1135 2356 1139
rect 2350 1134 2356 1135
rect 2386 1139 2392 1140
rect 2386 1135 2387 1139
rect 2391 1135 2392 1139
rect 2386 1134 2392 1135
rect 2416 1127 2418 1152
rect 2475 1140 2479 1141
rect 2492 1140 2494 1162
rect 2526 1157 2532 1158
rect 2526 1153 2527 1157
rect 2531 1153 2532 1157
rect 2526 1152 2532 1153
rect 2475 1135 2479 1136
rect 2490 1139 2496 1140
rect 2490 1135 2491 1139
rect 2495 1135 2496 1139
rect 2047 1126 2051 1127
rect 1623 1122 1627 1123
rect 1623 1117 1627 1118
rect 1687 1122 1691 1123
rect 1687 1117 1691 1118
rect 1839 1122 1843 1123
rect 1839 1117 1843 1118
rect 2007 1122 2011 1123
rect 2047 1121 2051 1122
rect 2311 1126 2315 1127
rect 2311 1121 2315 1122
rect 2407 1126 2411 1127
rect 2407 1121 2411 1122
rect 2415 1126 2419 1127
rect 2415 1121 2419 1122
rect 2007 1117 2011 1118
rect 1624 1096 1626 1117
rect 2008 1097 2010 1117
rect 2048 1101 2050 1121
rect 2046 1100 2052 1101
rect 2408 1100 2410 1121
rect 2476 1120 2478 1135
rect 2490 1134 2496 1135
rect 2528 1127 2530 1152
rect 2604 1140 2606 1162
rect 2638 1157 2644 1158
rect 2638 1153 2639 1157
rect 2643 1153 2644 1157
rect 2638 1152 2644 1153
rect 2602 1139 2608 1140
rect 2602 1135 2603 1139
rect 2607 1135 2608 1139
rect 2602 1134 2608 1135
rect 2640 1127 2642 1152
rect 2716 1140 2718 1162
rect 2724 1141 2726 1162
rect 2766 1157 2772 1158
rect 2766 1153 2767 1157
rect 2771 1153 2772 1157
rect 2766 1152 2772 1153
rect 2910 1157 2916 1158
rect 2910 1153 2911 1157
rect 2915 1153 2916 1157
rect 2910 1152 2916 1153
rect 2723 1140 2727 1141
rect 2714 1139 2720 1140
rect 2714 1135 2715 1139
rect 2719 1135 2720 1139
rect 2723 1135 2727 1136
rect 2714 1134 2720 1135
rect 2768 1127 2770 1152
rect 2912 1127 2914 1152
rect 2988 1140 2990 1162
rect 3070 1157 3076 1158
rect 3070 1153 3071 1157
rect 3075 1153 3076 1157
rect 3070 1152 3076 1153
rect 2986 1139 2992 1140
rect 2986 1135 2987 1139
rect 2991 1135 2992 1139
rect 2986 1134 2992 1135
rect 3072 1127 3074 1152
rect 2503 1126 2507 1127
rect 2503 1121 2507 1122
rect 2527 1126 2531 1127
rect 2527 1121 2531 1122
rect 2599 1126 2603 1127
rect 2599 1121 2603 1122
rect 2639 1126 2643 1127
rect 2639 1121 2643 1122
rect 2695 1126 2699 1127
rect 2695 1121 2699 1122
rect 2767 1126 2771 1127
rect 2767 1121 2771 1122
rect 2807 1126 2811 1127
rect 2807 1121 2811 1122
rect 2911 1126 2915 1127
rect 2911 1121 2915 1122
rect 2943 1126 2947 1127
rect 2943 1121 2947 1122
rect 3071 1126 3075 1127
rect 3071 1121 3075 1122
rect 3095 1126 3099 1127
rect 3095 1121 3099 1122
rect 2474 1119 2480 1120
rect 2474 1115 2475 1119
rect 2479 1115 2480 1119
rect 2474 1114 2480 1115
rect 2482 1119 2488 1120
rect 2482 1115 2483 1119
rect 2487 1115 2488 1119
rect 2482 1114 2488 1115
rect 2006 1096 2012 1097
rect 1622 1095 1628 1096
rect 1622 1091 1623 1095
rect 1627 1091 1628 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2046 1096 2047 1100
rect 2051 1096 2052 1100
rect 2046 1095 2052 1096
rect 2406 1099 2412 1100
rect 2406 1095 2407 1099
rect 2411 1095 2412 1099
rect 2406 1094 2412 1095
rect 2484 1092 2486 1114
rect 2504 1100 2506 1121
rect 2578 1119 2584 1120
rect 2578 1115 2579 1119
rect 2583 1115 2584 1119
rect 2578 1114 2584 1115
rect 2502 1099 2508 1100
rect 2502 1095 2503 1099
rect 2507 1095 2508 1099
rect 2502 1094 2508 1095
rect 2580 1092 2582 1114
rect 2600 1100 2602 1121
rect 2674 1119 2680 1120
rect 2674 1115 2675 1119
rect 2679 1115 2680 1119
rect 2674 1114 2680 1115
rect 2598 1099 2604 1100
rect 2598 1095 2599 1099
rect 2603 1095 2604 1099
rect 2598 1094 2604 1095
rect 2676 1092 2678 1114
rect 2696 1100 2698 1121
rect 2808 1100 2810 1121
rect 2902 1119 2908 1120
rect 2902 1115 2903 1119
rect 2907 1115 2908 1119
rect 2902 1114 2908 1115
rect 2694 1099 2700 1100
rect 2694 1095 2695 1099
rect 2699 1095 2700 1099
rect 2694 1094 2700 1095
rect 2806 1099 2812 1100
rect 2806 1095 2807 1099
rect 2811 1095 2812 1099
rect 2806 1094 2812 1095
rect 2904 1092 2906 1114
rect 2944 1100 2946 1121
rect 3096 1100 3098 1121
rect 3140 1120 3142 1162
rect 3246 1157 3252 1158
rect 3246 1153 3247 1157
rect 3251 1153 3252 1157
rect 3246 1152 3252 1153
rect 3248 1127 3250 1152
rect 3324 1140 3326 1162
rect 3380 1148 3382 1162
rect 3438 1157 3444 1158
rect 3438 1153 3439 1157
rect 3443 1153 3444 1157
rect 3438 1152 3444 1153
rect 3630 1157 3636 1158
rect 3630 1153 3631 1157
rect 3635 1153 3636 1157
rect 3630 1152 3636 1153
rect 3830 1157 3836 1158
rect 3830 1153 3831 1157
rect 3835 1153 3836 1157
rect 3830 1152 3836 1153
rect 3378 1147 3384 1148
rect 3378 1143 3379 1147
rect 3383 1143 3384 1147
rect 3378 1142 3384 1143
rect 3322 1139 3328 1140
rect 3322 1135 3323 1139
rect 3327 1135 3328 1139
rect 3322 1134 3328 1135
rect 3440 1127 3442 1152
rect 3632 1127 3634 1152
rect 3714 1135 3720 1136
rect 3714 1131 3715 1135
rect 3719 1131 3720 1135
rect 3714 1130 3720 1131
rect 3247 1126 3251 1127
rect 3247 1121 3251 1122
rect 3263 1126 3267 1127
rect 3263 1121 3267 1122
rect 3439 1126 3443 1127
rect 3439 1121 3443 1122
rect 3447 1126 3451 1127
rect 3447 1121 3451 1122
rect 3631 1126 3635 1127
rect 3631 1121 3635 1122
rect 3639 1126 3643 1127
rect 3639 1121 3643 1122
rect 3134 1119 3142 1120
rect 3134 1115 3135 1119
rect 3139 1116 3142 1119
rect 3170 1119 3176 1120
rect 3139 1115 3140 1116
rect 3134 1114 3140 1115
rect 3170 1115 3171 1119
rect 3175 1115 3176 1119
rect 3170 1114 3176 1115
rect 3142 1111 3148 1112
rect 3142 1107 3143 1111
rect 3147 1107 3148 1111
rect 3142 1106 3148 1107
rect 2942 1099 2948 1100
rect 2942 1095 2943 1099
rect 2947 1095 2948 1099
rect 2942 1094 2948 1095
rect 3094 1099 3100 1100
rect 3094 1095 3095 1099
rect 3099 1095 3100 1099
rect 3094 1094 3100 1095
rect 2006 1091 2012 1092
rect 2482 1091 2488 1092
rect 1622 1090 1628 1091
rect 1582 1087 1588 1088
rect 1582 1083 1583 1087
rect 1587 1083 1588 1087
rect 2482 1087 2483 1091
rect 2487 1087 2488 1091
rect 2482 1086 2488 1087
rect 2578 1091 2584 1092
rect 2578 1087 2579 1091
rect 2583 1087 2584 1091
rect 2578 1086 2584 1087
rect 2674 1091 2680 1092
rect 2674 1087 2675 1091
rect 2679 1087 2680 1091
rect 2674 1086 2680 1087
rect 2682 1091 2688 1092
rect 2682 1087 2683 1091
rect 2687 1087 2688 1091
rect 2902 1091 2908 1092
rect 2682 1086 2688 1087
rect 2894 1087 2900 1088
rect 1582 1082 1588 1083
rect 2046 1083 2052 1084
rect 2006 1079 2012 1080
rect 1622 1076 1628 1077
rect 1622 1072 1623 1076
rect 1627 1072 1628 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2046 1079 2047 1083
rect 2051 1079 2052 1083
rect 2046 1078 2052 1079
rect 2406 1080 2412 1081
rect 2006 1074 2012 1075
rect 1622 1071 1628 1072
rect 1624 1047 1626 1071
rect 2008 1047 2010 1074
rect 2048 1047 2050 1078
rect 2406 1076 2407 1080
rect 2411 1076 2412 1080
rect 2406 1075 2412 1076
rect 2502 1080 2508 1081
rect 2502 1076 2503 1080
rect 2507 1076 2508 1080
rect 2502 1075 2508 1076
rect 2598 1080 2604 1081
rect 2598 1076 2599 1080
rect 2603 1076 2604 1080
rect 2598 1075 2604 1076
rect 2408 1047 2410 1075
rect 2504 1047 2506 1075
rect 2600 1047 2602 1075
rect 1623 1046 1627 1047
rect 1623 1041 1627 1042
rect 2007 1046 2011 1047
rect 2007 1041 2011 1042
rect 2047 1046 2051 1047
rect 2047 1041 2051 1042
rect 2407 1046 2411 1047
rect 2407 1041 2411 1042
rect 2455 1046 2459 1047
rect 2455 1041 2459 1042
rect 2503 1046 2507 1047
rect 2503 1041 2507 1042
rect 2551 1046 2555 1047
rect 2551 1041 2555 1042
rect 2599 1046 2603 1047
rect 2599 1041 2603 1042
rect 2647 1046 2651 1047
rect 2647 1041 2651 1042
rect 2008 1014 2010 1041
rect 2048 1014 2050 1041
rect 2456 1017 2458 1041
rect 2552 1017 2554 1041
rect 2648 1017 2650 1041
rect 2454 1016 2460 1017
rect 2006 1013 2012 1014
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1013 2052 1014
rect 2046 1009 2047 1013
rect 2051 1009 2052 1013
rect 2454 1012 2455 1016
rect 2459 1012 2460 1016
rect 2454 1011 2460 1012
rect 2550 1016 2556 1017
rect 2550 1012 2551 1016
rect 2555 1012 2556 1016
rect 2550 1011 2556 1012
rect 2646 1016 2652 1017
rect 2646 1012 2647 1016
rect 2651 1012 2652 1016
rect 2646 1011 2652 1012
rect 2046 1008 2052 1009
rect 802 1007 808 1008
rect 802 1003 803 1007
rect 807 1003 808 1007
rect 802 1002 808 1003
rect 810 1007 816 1008
rect 810 1003 811 1007
rect 815 1003 816 1007
rect 810 1002 816 1003
rect 1050 1007 1056 1008
rect 1050 1003 1051 1007
rect 1055 1003 1056 1007
rect 1050 1002 1056 1003
rect 1162 1007 1168 1008
rect 1162 1003 1163 1007
rect 1167 1003 1168 1007
rect 1162 1002 1168 1003
rect 1274 1007 1280 1008
rect 1274 1003 1275 1007
rect 1279 1003 1280 1007
rect 1274 1002 1280 1003
rect 1386 1007 1392 1008
rect 1386 1003 1387 1007
rect 1391 1003 1392 1007
rect 1386 1002 1392 1003
rect 1498 1007 1504 1008
rect 1498 1003 1499 1007
rect 1503 1003 1504 1007
rect 1498 1002 1504 1003
rect 2542 1007 2548 1008
rect 2542 1003 2543 1007
rect 2547 1003 2548 1007
rect 2542 1002 2548 1003
rect 804 980 806 1002
rect 812 988 814 1002
rect 854 997 860 998
rect 854 993 855 997
rect 859 993 860 997
rect 854 992 860 993
rect 974 997 980 998
rect 974 993 975 997
rect 979 993 980 997
rect 974 992 980 993
rect 810 987 816 988
rect 810 983 811 987
rect 815 983 816 987
rect 810 982 816 983
rect 786 979 792 980
rect 786 975 787 979
rect 791 975 792 979
rect 786 974 792 975
rect 802 979 808 980
rect 802 975 803 979
rect 807 975 808 979
rect 802 974 808 975
rect 856 971 858 992
rect 976 971 978 992
rect 1052 980 1054 1002
rect 1086 997 1092 998
rect 1086 993 1087 997
rect 1091 993 1092 997
rect 1086 992 1092 993
rect 1050 979 1056 980
rect 1042 975 1048 976
rect 1042 971 1043 975
rect 1047 971 1048 975
rect 1050 975 1051 979
rect 1055 975 1056 979
rect 1050 974 1056 975
rect 1088 971 1090 992
rect 1164 980 1166 1002
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1162 979 1168 980
rect 1162 975 1163 979
rect 1167 975 1168 979
rect 1162 974 1168 975
rect 1200 971 1202 992
rect 1276 980 1278 1002
rect 1310 997 1316 998
rect 1310 993 1311 997
rect 1315 993 1316 997
rect 1310 992 1316 993
rect 1274 979 1280 980
rect 1274 975 1275 979
rect 1279 975 1280 979
rect 1274 974 1280 975
rect 1312 971 1314 992
rect 1388 980 1390 1002
rect 1430 997 1436 998
rect 2454 997 2460 998
rect 1430 993 1431 997
rect 1435 993 1436 997
rect 1430 992 1436 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 1386 979 1392 980
rect 1386 975 1387 979
rect 1391 975 1392 979
rect 1386 974 1392 975
rect 1432 971 1434 992
rect 2006 991 2012 992
rect 2046 996 2052 997
rect 2046 992 2047 996
rect 2051 992 2052 996
rect 2454 993 2455 997
rect 2459 993 2460 997
rect 2454 992 2460 993
rect 2046 991 2052 992
rect 2008 971 2010 991
rect 727 970 731 971
rect 727 965 731 966
rect 807 970 811 971
rect 807 965 811 966
rect 855 970 859 971
rect 855 965 859 966
rect 975 970 979 971
rect 1042 970 1048 971
rect 1087 970 1091 971
rect 975 965 979 966
rect 666 963 672 964
rect 666 959 667 963
rect 671 959 672 963
rect 666 958 672 959
rect 706 963 712 964
rect 706 959 707 963
rect 711 959 712 963
rect 706 958 712 959
rect 630 943 636 944
rect 630 939 631 943
rect 635 939 636 943
rect 630 938 636 939
rect 708 936 710 958
rect 808 944 810 965
rect 882 963 888 964
rect 882 959 883 963
rect 887 959 888 963
rect 882 958 888 959
rect 806 943 812 944
rect 806 939 807 943
rect 811 939 812 943
rect 806 938 812 939
rect 884 936 886 958
rect 976 944 978 965
rect 974 943 980 944
rect 974 939 975 943
rect 979 939 980 943
rect 1044 940 1046 970
rect 1087 965 1091 966
rect 1127 970 1131 971
rect 1127 965 1131 966
rect 1199 970 1203 971
rect 1199 965 1203 966
rect 1271 970 1275 971
rect 1271 965 1275 966
rect 1311 970 1315 971
rect 1311 965 1315 966
rect 1415 970 1419 971
rect 1415 965 1419 966
rect 1431 970 1435 971
rect 1431 965 1435 966
rect 1551 970 1555 971
rect 1551 965 1555 966
rect 1695 970 1699 971
rect 1695 965 1699 966
rect 2007 970 2011 971
rect 2048 967 2050 991
rect 2456 967 2458 992
rect 2544 980 2546 1002
rect 2550 997 2556 998
rect 2550 993 2551 997
rect 2555 993 2556 997
rect 2550 992 2556 993
rect 2646 997 2652 998
rect 2646 993 2647 997
rect 2651 993 2652 997
rect 2646 992 2652 993
rect 2542 979 2548 980
rect 2542 975 2543 979
rect 2547 975 2548 979
rect 2542 974 2548 975
rect 2552 967 2554 992
rect 2648 967 2650 992
rect 2684 988 2686 1086
rect 2894 1083 2895 1087
rect 2899 1083 2900 1087
rect 2902 1087 2903 1091
rect 2907 1087 2908 1091
rect 2902 1086 2908 1087
rect 2894 1082 2900 1083
rect 2694 1080 2700 1081
rect 2694 1076 2695 1080
rect 2699 1076 2700 1080
rect 2694 1075 2700 1076
rect 2806 1080 2812 1081
rect 2806 1076 2807 1080
rect 2811 1076 2812 1080
rect 2806 1075 2812 1076
rect 2696 1047 2698 1075
rect 2808 1047 2810 1075
rect 2695 1046 2699 1047
rect 2695 1041 2699 1042
rect 2759 1046 2763 1047
rect 2759 1041 2763 1042
rect 2807 1046 2811 1047
rect 2807 1041 2811 1042
rect 2887 1046 2891 1047
rect 2887 1041 2891 1042
rect 2760 1017 2762 1041
rect 2888 1017 2890 1041
rect 2758 1016 2764 1017
rect 2758 1012 2759 1016
rect 2763 1012 2764 1016
rect 2758 1011 2764 1012
rect 2886 1016 2892 1017
rect 2886 1012 2887 1016
rect 2891 1012 2892 1016
rect 2886 1011 2892 1012
rect 2722 1007 2728 1008
rect 2722 1003 2723 1007
rect 2727 1003 2728 1007
rect 2722 1002 2728 1003
rect 2834 1007 2840 1008
rect 2834 1003 2835 1007
rect 2839 1003 2840 1007
rect 2834 1002 2840 1003
rect 2858 1007 2864 1008
rect 2858 1003 2859 1007
rect 2863 1003 2864 1007
rect 2858 1002 2864 1003
rect 2682 987 2688 988
rect 2682 983 2683 987
rect 2687 983 2688 987
rect 2682 982 2688 983
rect 2007 965 2011 966
rect 2047 966 2051 967
rect 1128 944 1130 965
rect 1210 963 1216 964
rect 1210 959 1211 963
rect 1215 959 1216 963
rect 1210 958 1216 959
rect 1126 943 1132 944
rect 974 938 980 939
rect 1042 939 1048 940
rect 330 935 336 936
rect 330 931 331 935
rect 335 931 336 935
rect 330 930 336 931
rect 522 935 528 936
rect 522 931 523 935
rect 527 931 528 935
rect 522 930 528 931
rect 706 935 712 936
rect 706 931 707 935
rect 711 931 712 935
rect 706 930 712 931
rect 882 935 888 936
rect 882 931 883 935
rect 887 931 888 935
rect 1042 935 1043 939
rect 1047 935 1048 939
rect 1126 939 1127 943
rect 1131 939 1132 943
rect 1126 938 1132 939
rect 1212 936 1214 958
rect 1272 944 1274 965
rect 1354 963 1360 964
rect 1354 959 1355 963
rect 1359 959 1360 963
rect 1354 958 1360 959
rect 1270 943 1276 944
rect 1270 939 1271 943
rect 1275 939 1276 943
rect 1270 938 1276 939
rect 1356 936 1358 958
rect 1416 944 1418 965
rect 1498 963 1504 964
rect 1498 959 1499 963
rect 1503 959 1504 963
rect 1498 958 1504 959
rect 1414 943 1420 944
rect 1414 939 1415 943
rect 1419 939 1420 943
rect 1414 938 1420 939
rect 1500 936 1502 958
rect 1552 944 1554 965
rect 1634 963 1640 964
rect 1634 959 1635 963
rect 1639 959 1640 963
rect 1634 958 1640 959
rect 1550 943 1556 944
rect 1550 939 1551 943
rect 1555 939 1556 943
rect 1550 938 1556 939
rect 1636 936 1638 958
rect 1696 944 1698 965
rect 1734 963 1740 964
rect 1734 959 1735 963
rect 1739 959 1740 963
rect 1734 958 1740 959
rect 1694 943 1700 944
rect 1694 939 1695 943
rect 1699 939 1700 943
rect 1694 938 1700 939
rect 1042 934 1048 935
rect 1210 935 1216 936
rect 882 930 888 931
rect 1050 931 1056 932
rect 1050 927 1051 931
rect 1055 927 1056 931
rect 1210 931 1211 935
rect 1215 931 1216 935
rect 1210 930 1216 931
rect 1354 935 1360 936
rect 1354 931 1355 935
rect 1359 931 1360 935
rect 1354 930 1360 931
rect 1498 935 1504 936
rect 1498 931 1499 935
rect 1503 931 1504 935
rect 1498 930 1504 931
rect 1634 935 1640 936
rect 1634 931 1635 935
rect 1639 931 1640 935
rect 1634 930 1640 931
rect 1050 926 1056 927
rect 446 924 452 925
rect 446 920 447 924
rect 451 920 452 924
rect 446 919 452 920
rect 630 924 636 925
rect 630 920 631 924
rect 635 920 636 924
rect 630 919 636 920
rect 806 924 812 925
rect 806 920 807 924
rect 811 920 812 924
rect 806 919 812 920
rect 974 924 980 925
rect 974 920 975 924
rect 979 920 980 924
rect 974 919 980 920
rect 448 891 450 919
rect 632 891 634 919
rect 808 891 810 919
rect 976 891 978 919
rect 447 890 451 891
rect 447 885 451 886
rect 631 890 635 891
rect 631 885 635 886
rect 639 890 643 891
rect 639 885 643 886
rect 807 890 811 891
rect 807 885 811 886
rect 823 890 827 891
rect 823 885 827 886
rect 975 890 979 891
rect 975 885 979 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 448 861 450 885
rect 640 861 642 885
rect 824 861 826 885
rect 1000 861 1002 885
rect 446 860 452 861
rect 446 856 447 860
rect 451 856 452 860
rect 446 855 452 856
rect 638 860 644 861
rect 638 856 639 860
rect 643 856 644 860
rect 638 855 644 856
rect 822 860 828 861
rect 822 856 823 860
rect 827 856 828 860
rect 822 855 828 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 322 851 328 852
rect 322 847 323 851
rect 327 847 328 851
rect 322 846 328 847
rect 514 851 520 852
rect 514 847 515 851
rect 519 847 520 851
rect 514 846 520 847
rect 566 851 572 852
rect 566 847 567 851
rect 571 847 572 851
rect 566 846 572 847
rect 770 851 776 852
rect 770 847 771 851
rect 775 847 776 851
rect 770 846 776 847
rect 254 841 260 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 254 837 255 841
rect 259 837 260 841
rect 254 836 260 837
rect 446 841 452 842
rect 446 837 447 841
rect 451 837 452 841
rect 446 836 452 837
rect 110 835 116 836
rect 112 811 114 835
rect 234 819 240 820
rect 234 815 235 819
rect 239 815 240 819
rect 234 814 240 815
rect 111 810 115 811
rect 111 805 115 806
rect 159 810 163 811
rect 159 805 163 806
rect 112 785 114 805
rect 110 784 116 785
rect 160 784 162 805
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 158 783 164 784
rect 158 779 159 783
rect 163 779 164 783
rect 158 778 164 779
rect 236 776 238 814
rect 256 811 258 836
rect 448 811 450 836
rect 255 810 259 811
rect 255 805 259 806
rect 311 810 315 811
rect 311 805 315 806
rect 447 810 451 811
rect 447 805 451 806
rect 471 810 475 811
rect 471 805 475 806
rect 312 784 314 805
rect 338 803 344 804
rect 338 799 339 803
rect 343 799 344 803
rect 338 798 344 799
rect 310 783 316 784
rect 310 779 311 783
rect 315 779 316 783
rect 310 778 316 779
rect 234 775 240 776
rect 234 771 235 775
rect 239 771 240 775
rect 234 770 240 771
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 110 762 116 763
rect 158 764 164 765
rect 112 735 114 762
rect 158 760 159 764
rect 163 760 164 764
rect 158 759 164 760
rect 310 764 316 765
rect 310 760 311 764
rect 315 760 316 764
rect 310 759 316 760
rect 160 735 162 759
rect 312 735 314 759
rect 111 734 115 735
rect 111 729 115 730
rect 135 734 139 735
rect 135 729 139 730
rect 159 734 163 735
rect 159 729 163 730
rect 263 734 267 735
rect 263 729 267 730
rect 311 734 315 735
rect 311 729 315 730
rect 112 702 114 729
rect 136 705 138 729
rect 264 705 266 729
rect 134 704 140 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 134 700 135 704
rect 139 700 140 704
rect 134 699 140 700
rect 262 704 268 705
rect 262 700 263 704
rect 267 700 268 704
rect 262 699 268 700
rect 110 696 116 697
rect 340 696 342 798
rect 472 784 474 805
rect 516 804 518 846
rect 568 824 570 846
rect 638 841 644 842
rect 638 837 639 841
rect 643 837 644 841
rect 638 836 644 837
rect 566 823 572 824
rect 566 819 567 823
rect 571 819 572 823
rect 566 818 572 819
rect 640 811 642 836
rect 772 824 774 846
rect 822 841 828 842
rect 822 837 823 841
rect 827 837 828 841
rect 822 836 828 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 770 823 776 824
rect 770 819 771 823
rect 775 819 776 823
rect 770 818 776 819
rect 824 811 826 836
rect 1000 811 1002 836
rect 1052 824 1054 926
rect 1126 924 1132 925
rect 1126 920 1127 924
rect 1131 920 1132 924
rect 1126 919 1132 920
rect 1270 924 1276 925
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1414 924 1420 925
rect 1414 920 1415 924
rect 1419 920 1420 924
rect 1414 919 1420 920
rect 1550 924 1556 925
rect 1550 920 1551 924
rect 1555 920 1556 924
rect 1550 919 1556 920
rect 1694 924 1700 925
rect 1694 920 1695 924
rect 1699 920 1700 924
rect 1694 919 1700 920
rect 1128 891 1130 919
rect 1272 891 1274 919
rect 1416 891 1418 919
rect 1552 891 1554 919
rect 1696 891 1698 919
rect 1127 890 1131 891
rect 1127 885 1131 886
rect 1167 890 1171 891
rect 1167 885 1171 886
rect 1271 890 1275 891
rect 1271 885 1275 886
rect 1327 890 1331 891
rect 1327 885 1331 886
rect 1415 890 1419 891
rect 1415 885 1419 886
rect 1479 890 1483 891
rect 1479 885 1483 886
rect 1551 890 1555 891
rect 1551 885 1555 886
rect 1631 890 1635 891
rect 1631 885 1635 886
rect 1695 890 1699 891
rect 1695 885 1699 886
rect 1168 861 1170 885
rect 1328 861 1330 885
rect 1480 861 1482 885
rect 1632 861 1634 885
rect 1166 860 1172 861
rect 1166 856 1167 860
rect 1171 856 1172 860
rect 1166 855 1172 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1478 860 1484 861
rect 1478 856 1479 860
rect 1483 856 1484 860
rect 1478 855 1484 856
rect 1630 860 1636 861
rect 1630 856 1631 860
rect 1635 856 1636 860
rect 1630 855 1636 856
rect 1736 852 1738 958
rect 2008 945 2010 965
rect 2047 961 2051 962
rect 2423 966 2427 967
rect 2423 961 2427 962
rect 2455 966 2459 967
rect 2455 961 2459 962
rect 2519 966 2523 967
rect 2519 961 2523 962
rect 2551 966 2555 967
rect 2551 961 2555 962
rect 2615 966 2619 967
rect 2615 961 2619 962
rect 2647 966 2651 967
rect 2647 961 2651 962
rect 2711 966 2715 967
rect 2711 961 2715 962
rect 2006 944 2012 945
rect 2006 940 2007 944
rect 2011 940 2012 944
rect 2048 941 2050 961
rect 2006 939 2012 940
rect 2046 940 2052 941
rect 2424 940 2426 961
rect 2498 959 2504 960
rect 2498 955 2499 959
rect 2503 955 2504 959
rect 2498 954 2504 955
rect 2046 936 2047 940
rect 2051 936 2052 940
rect 2046 935 2052 936
rect 2422 939 2428 940
rect 2422 935 2423 939
rect 2427 935 2428 939
rect 2422 934 2428 935
rect 2500 932 2502 954
rect 2520 940 2522 961
rect 2594 959 2600 960
rect 2594 955 2595 959
rect 2599 955 2600 959
rect 2594 954 2600 955
rect 2518 939 2524 940
rect 2518 935 2519 939
rect 2523 935 2524 939
rect 2518 934 2524 935
rect 2596 932 2598 954
rect 2616 940 2618 961
rect 2712 940 2714 961
rect 2724 960 2726 1002
rect 2758 997 2764 998
rect 2758 993 2759 997
rect 2763 993 2764 997
rect 2758 992 2764 993
rect 2760 967 2762 992
rect 2786 975 2792 976
rect 2786 971 2787 975
rect 2791 971 2792 975
rect 2786 970 2792 971
rect 2759 966 2763 967
rect 2759 961 2763 962
rect 2722 959 2728 960
rect 2722 955 2723 959
rect 2727 955 2728 959
rect 2722 954 2728 955
rect 2614 939 2620 940
rect 2614 935 2615 939
rect 2619 935 2620 939
rect 2614 934 2620 935
rect 2710 939 2716 940
rect 2710 935 2711 939
rect 2715 935 2716 939
rect 2710 934 2716 935
rect 2788 932 2790 970
rect 2823 966 2827 967
rect 2823 961 2827 962
rect 2824 940 2826 961
rect 2836 960 2838 1002
rect 2860 984 2862 1002
rect 2886 997 2892 998
rect 2886 993 2887 997
rect 2891 993 2892 997
rect 2886 992 2892 993
rect 2858 983 2864 984
rect 2858 979 2859 983
rect 2863 979 2864 983
rect 2858 978 2864 979
rect 2888 967 2890 992
rect 2896 980 2898 1082
rect 2942 1080 2948 1081
rect 2942 1076 2943 1080
rect 2947 1076 2948 1080
rect 2942 1075 2948 1076
rect 3094 1080 3100 1081
rect 3094 1076 3095 1080
rect 3099 1076 3100 1080
rect 3094 1075 3100 1076
rect 2944 1047 2946 1075
rect 3096 1047 3098 1075
rect 2943 1046 2947 1047
rect 2943 1041 2947 1042
rect 3031 1046 3035 1047
rect 3031 1041 3035 1042
rect 3095 1046 3099 1047
rect 3095 1041 3099 1042
rect 3032 1017 3034 1041
rect 3030 1016 3036 1017
rect 3030 1012 3031 1016
rect 3035 1012 3036 1016
rect 3030 1011 3036 1012
rect 3144 1008 3146 1106
rect 3172 1092 3174 1114
rect 3264 1100 3266 1121
rect 3338 1119 3344 1120
rect 3338 1115 3339 1119
rect 3343 1115 3344 1119
rect 3338 1114 3344 1115
rect 3262 1099 3268 1100
rect 3262 1095 3263 1099
rect 3267 1095 3268 1099
rect 3262 1094 3268 1095
rect 3340 1092 3342 1114
rect 3448 1100 3450 1121
rect 3578 1119 3584 1120
rect 3578 1115 3579 1119
rect 3583 1115 3584 1119
rect 3578 1114 3584 1115
rect 3446 1099 3452 1100
rect 3446 1095 3447 1099
rect 3451 1095 3452 1099
rect 3446 1094 3452 1095
rect 3170 1091 3176 1092
rect 3170 1087 3171 1091
rect 3175 1087 3176 1091
rect 3170 1086 3176 1087
rect 3338 1091 3344 1092
rect 3338 1087 3339 1091
rect 3343 1087 3344 1091
rect 3338 1086 3344 1087
rect 3382 1091 3388 1092
rect 3382 1087 3383 1091
rect 3387 1087 3388 1091
rect 3382 1086 3388 1087
rect 3262 1080 3268 1081
rect 3262 1076 3263 1080
rect 3267 1076 3268 1080
rect 3262 1075 3268 1076
rect 3264 1047 3266 1075
rect 3183 1046 3187 1047
rect 3183 1041 3187 1042
rect 3263 1046 3267 1047
rect 3263 1041 3267 1042
rect 3343 1046 3347 1047
rect 3343 1041 3347 1042
rect 3184 1017 3186 1041
rect 3344 1017 3346 1041
rect 3182 1016 3188 1017
rect 3182 1012 3183 1016
rect 3187 1012 3188 1016
rect 3182 1011 3188 1012
rect 3342 1016 3348 1017
rect 3342 1012 3343 1016
rect 3347 1012 3348 1016
rect 3342 1011 3348 1012
rect 2990 1007 2996 1008
rect 2990 1003 2991 1007
rect 2995 1003 2996 1007
rect 2990 1002 2996 1003
rect 3142 1007 3148 1008
rect 3142 1003 3143 1007
rect 3147 1003 3148 1007
rect 3142 1002 3148 1003
rect 3294 1007 3300 1008
rect 3294 1003 3295 1007
rect 3299 1003 3300 1007
rect 3294 1002 3300 1003
rect 2894 979 2900 980
rect 2894 975 2895 979
rect 2899 975 2900 979
rect 2894 974 2900 975
rect 2942 975 2948 976
rect 2942 971 2943 975
rect 2947 971 2948 975
rect 2942 970 2948 971
rect 2887 966 2891 967
rect 2887 961 2891 962
rect 2834 959 2840 960
rect 2834 955 2835 959
rect 2839 955 2840 959
rect 2834 954 2840 955
rect 2822 939 2828 940
rect 2822 935 2823 939
rect 2827 935 2828 939
rect 2822 934 2828 935
rect 2944 932 2946 970
rect 2951 966 2955 967
rect 2951 961 2955 962
rect 2952 940 2954 961
rect 2992 960 2994 1002
rect 3030 997 3036 998
rect 3030 993 3031 997
rect 3035 993 3036 997
rect 3030 992 3036 993
rect 3182 997 3188 998
rect 3182 993 3183 997
rect 3187 993 3188 997
rect 3182 992 3188 993
rect 3032 967 3034 992
rect 3184 967 3186 992
rect 3296 980 3298 1002
rect 3342 997 3348 998
rect 3342 993 3343 997
rect 3347 993 3348 997
rect 3342 992 3348 993
rect 3294 979 3300 980
rect 3294 975 3295 979
rect 3299 975 3300 979
rect 3294 974 3300 975
rect 3344 967 3346 992
rect 3384 980 3386 1086
rect 3446 1080 3452 1081
rect 3446 1076 3447 1080
rect 3451 1076 3452 1080
rect 3446 1075 3452 1076
rect 3448 1047 3450 1075
rect 3447 1046 3451 1047
rect 3447 1041 3451 1042
rect 3503 1046 3507 1047
rect 3503 1041 3507 1042
rect 3504 1017 3506 1041
rect 3502 1016 3508 1017
rect 3502 1012 3503 1016
rect 3507 1012 3508 1016
rect 3502 1011 3508 1012
rect 3580 1008 3582 1114
rect 3640 1100 3642 1121
rect 3638 1099 3644 1100
rect 3638 1095 3639 1099
rect 3643 1095 3644 1099
rect 3638 1094 3644 1095
rect 3716 1092 3718 1130
rect 3832 1127 3834 1152
rect 3884 1140 3886 1238
rect 3942 1235 3943 1239
rect 3947 1235 3948 1239
rect 3942 1234 3948 1235
rect 3944 1207 3946 1234
rect 3943 1206 3947 1207
rect 3943 1201 3947 1202
rect 3944 1174 3946 1201
rect 3942 1173 3948 1174
rect 3942 1169 3943 1173
rect 3947 1169 3948 1173
rect 3942 1168 3948 1169
rect 3898 1167 3904 1168
rect 3898 1163 3899 1167
rect 3903 1163 3904 1167
rect 3898 1162 3904 1163
rect 3882 1139 3888 1140
rect 3882 1135 3883 1139
rect 3887 1135 3888 1139
rect 3882 1134 3888 1135
rect 3831 1126 3835 1127
rect 3831 1121 3835 1122
rect 3839 1126 3843 1127
rect 3839 1121 3843 1122
rect 3840 1100 3842 1121
rect 3900 1120 3902 1162
rect 3942 1156 3948 1157
rect 3942 1152 3943 1156
rect 3947 1152 3948 1156
rect 3942 1151 3948 1152
rect 3944 1127 3946 1151
rect 3943 1126 3947 1127
rect 3943 1121 3947 1122
rect 3898 1119 3904 1120
rect 3898 1115 3899 1119
rect 3903 1115 3904 1119
rect 3898 1114 3904 1115
rect 3944 1101 3946 1121
rect 3942 1100 3948 1101
rect 3838 1099 3844 1100
rect 3838 1095 3839 1099
rect 3843 1095 3844 1099
rect 3942 1096 3943 1100
rect 3947 1096 3948 1100
rect 3942 1095 3948 1096
rect 3838 1094 3844 1095
rect 3714 1091 3720 1092
rect 3714 1087 3715 1091
rect 3719 1087 3720 1091
rect 3714 1086 3720 1087
rect 3914 1087 3920 1088
rect 3914 1083 3915 1087
rect 3919 1083 3920 1087
rect 3914 1082 3920 1083
rect 3942 1083 3948 1084
rect 3638 1080 3644 1081
rect 3638 1076 3639 1080
rect 3643 1076 3644 1080
rect 3638 1075 3644 1076
rect 3838 1080 3844 1081
rect 3838 1076 3839 1080
rect 3843 1076 3844 1080
rect 3838 1075 3844 1076
rect 3640 1047 3642 1075
rect 3840 1047 3842 1075
rect 3639 1046 3643 1047
rect 3639 1041 3643 1042
rect 3671 1046 3675 1047
rect 3671 1041 3675 1042
rect 3839 1046 3843 1047
rect 3839 1041 3843 1042
rect 3672 1017 3674 1041
rect 3840 1017 3842 1041
rect 3670 1016 3676 1017
rect 3670 1012 3671 1016
rect 3675 1012 3676 1016
rect 3670 1011 3676 1012
rect 3838 1016 3844 1017
rect 3838 1012 3839 1016
rect 3843 1012 3844 1016
rect 3838 1011 3844 1012
rect 3578 1007 3584 1008
rect 3578 1003 3579 1007
rect 3583 1003 3584 1007
rect 3578 1002 3584 1003
rect 3906 1007 3912 1008
rect 3906 1003 3907 1007
rect 3911 1003 3912 1007
rect 3906 1002 3912 1003
rect 3502 997 3508 998
rect 3502 993 3503 997
rect 3507 993 3508 997
rect 3502 992 3508 993
rect 3670 997 3676 998
rect 3670 993 3671 997
rect 3675 993 3676 997
rect 3670 992 3676 993
rect 3838 997 3844 998
rect 3838 993 3839 997
rect 3843 993 3844 997
rect 3838 992 3844 993
rect 3382 979 3388 980
rect 3382 975 3383 979
rect 3387 975 3388 979
rect 3382 974 3388 975
rect 3504 967 3506 992
rect 3672 967 3674 992
rect 3722 975 3728 976
rect 3722 971 3723 975
rect 3727 971 3728 975
rect 3722 970 3728 971
rect 3031 966 3035 967
rect 3031 961 3035 962
rect 3103 966 3107 967
rect 3103 961 3107 962
rect 3183 966 3187 967
rect 3183 961 3187 962
rect 3271 966 3275 967
rect 3271 961 3275 962
rect 3343 966 3347 967
rect 3343 961 3347 962
rect 3455 966 3459 967
rect 3455 961 3459 962
rect 3503 966 3507 967
rect 3503 961 3507 962
rect 3647 966 3651 967
rect 3647 961 3651 962
rect 3671 966 3675 967
rect 3671 961 3675 962
rect 2990 959 2996 960
rect 2990 955 2991 959
rect 2995 955 2996 959
rect 2990 954 2996 955
rect 3046 959 3052 960
rect 3046 955 3047 959
rect 3051 955 3052 959
rect 3046 954 3052 955
rect 2950 939 2956 940
rect 2950 935 2951 939
rect 2955 935 2956 939
rect 2950 934 2956 935
rect 3048 932 3050 954
rect 3104 940 3106 961
rect 3272 940 3274 961
rect 3456 940 3458 961
rect 3648 940 3650 961
rect 3686 959 3692 960
rect 3686 955 3687 959
rect 3691 955 3692 959
rect 3686 954 3692 955
rect 3102 939 3108 940
rect 3102 935 3103 939
rect 3107 935 3108 939
rect 3102 934 3108 935
rect 3270 939 3276 940
rect 3270 935 3271 939
rect 3275 935 3276 939
rect 3270 934 3276 935
rect 3454 939 3460 940
rect 3454 935 3455 939
rect 3459 935 3460 939
rect 3454 934 3460 935
rect 3646 939 3652 940
rect 3646 935 3647 939
rect 3651 935 3652 939
rect 3646 934 3652 935
rect 2498 931 2504 932
rect 2006 927 2012 928
rect 2006 923 2007 927
rect 2011 923 2012 927
rect 2498 927 2499 931
rect 2503 927 2504 931
rect 2498 926 2504 927
rect 2594 931 2600 932
rect 2594 927 2595 931
rect 2599 927 2600 931
rect 2786 931 2792 932
rect 2594 926 2600 927
rect 2690 927 2696 928
rect 2006 922 2012 923
rect 2046 923 2052 924
rect 2008 891 2010 922
rect 2046 919 2047 923
rect 2051 919 2052 923
rect 2690 923 2691 927
rect 2695 923 2696 927
rect 2786 927 2787 931
rect 2791 927 2792 931
rect 2786 926 2792 927
rect 2942 931 2948 932
rect 2942 927 2943 931
rect 2947 927 2948 931
rect 2942 926 2948 927
rect 3046 931 3052 932
rect 3046 927 3047 931
rect 3051 927 3052 931
rect 3046 926 3052 927
rect 3410 931 3416 932
rect 3410 927 3411 931
rect 3415 927 3416 931
rect 3410 926 3416 927
rect 2690 922 2696 923
rect 2046 918 2052 919
rect 2422 920 2428 921
rect 2048 891 2050 918
rect 2422 916 2423 920
rect 2427 916 2428 920
rect 2422 915 2428 916
rect 2518 920 2524 921
rect 2518 916 2519 920
rect 2523 916 2524 920
rect 2518 915 2524 916
rect 2614 920 2620 921
rect 2614 916 2615 920
rect 2619 916 2620 920
rect 2614 915 2620 916
rect 2424 891 2426 915
rect 2520 891 2522 915
rect 2616 891 2618 915
rect 1783 890 1787 891
rect 1783 885 1787 886
rect 2007 890 2011 891
rect 2007 885 2011 886
rect 2047 890 2051 891
rect 2047 885 2051 886
rect 2343 890 2347 891
rect 2343 885 2347 886
rect 2423 890 2427 891
rect 2423 885 2427 886
rect 2439 890 2443 891
rect 2439 885 2443 886
rect 2519 890 2523 891
rect 2519 885 2523 886
rect 2535 890 2539 891
rect 2535 885 2539 886
rect 2615 890 2619 891
rect 2615 885 2619 886
rect 2631 890 2635 891
rect 2631 885 2635 886
rect 1784 861 1786 885
rect 1782 860 1788 861
rect 1782 856 1783 860
rect 1787 856 1788 860
rect 2008 858 2010 885
rect 2048 858 2050 885
rect 2344 861 2346 885
rect 2440 861 2442 885
rect 2536 861 2538 885
rect 2632 861 2634 885
rect 2342 860 2348 861
rect 1782 855 1788 856
rect 2006 857 2012 858
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2006 852 2012 853
rect 2046 857 2052 858
rect 2046 853 2047 857
rect 2051 853 2052 857
rect 2342 856 2343 860
rect 2347 856 2348 860
rect 2342 855 2348 856
rect 2438 860 2444 861
rect 2438 856 2439 860
rect 2443 856 2444 860
rect 2438 855 2444 856
rect 2534 860 2540 861
rect 2534 856 2535 860
rect 2539 856 2540 860
rect 2534 855 2540 856
rect 2630 860 2636 861
rect 2630 856 2631 860
rect 2635 856 2636 860
rect 2630 855 2636 856
rect 2046 852 2052 853
rect 1242 851 1248 852
rect 1242 847 1243 851
rect 1247 847 1248 851
rect 1242 846 1248 847
rect 1402 851 1408 852
rect 1402 847 1403 851
rect 1407 847 1408 851
rect 1402 846 1408 847
rect 1554 851 1560 852
rect 1554 847 1555 851
rect 1559 847 1560 851
rect 1554 846 1560 847
rect 1706 851 1712 852
rect 1706 847 1707 851
rect 1711 847 1712 851
rect 1706 846 1712 847
rect 1734 851 1740 852
rect 1734 847 1735 851
rect 1739 847 1740 851
rect 1734 846 1740 847
rect 2430 851 2436 852
rect 2430 847 2431 851
rect 2435 847 2436 851
rect 2430 846 2436 847
rect 2526 851 2532 852
rect 2526 847 2527 851
rect 2531 847 2532 851
rect 2526 846 2532 847
rect 1166 841 1172 842
rect 1166 837 1167 841
rect 1171 837 1172 841
rect 1166 836 1172 837
rect 1050 823 1056 824
rect 1050 819 1051 823
rect 1055 819 1056 823
rect 1050 818 1056 819
rect 1168 811 1170 836
rect 1244 824 1246 846
rect 1326 841 1332 842
rect 1326 837 1327 841
rect 1331 837 1332 841
rect 1326 836 1332 837
rect 1242 823 1248 824
rect 1242 819 1243 823
rect 1247 819 1248 823
rect 1242 818 1248 819
rect 1328 811 1330 836
rect 1404 824 1406 846
rect 1478 841 1484 842
rect 1478 837 1479 841
rect 1483 837 1484 841
rect 1478 836 1484 837
rect 1402 823 1408 824
rect 1402 819 1403 823
rect 1407 819 1408 823
rect 1402 818 1408 819
rect 1480 811 1482 836
rect 1556 824 1558 846
rect 1630 841 1636 842
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1554 823 1560 824
rect 1554 819 1555 823
rect 1559 819 1560 823
rect 1554 818 1560 819
rect 1518 815 1524 816
rect 1518 811 1519 815
rect 1523 811 1524 815
rect 1632 811 1634 836
rect 1708 824 1710 846
rect 1782 841 1788 842
rect 2342 841 2348 842
rect 1782 837 1783 841
rect 1787 837 1788 841
rect 1782 836 1788 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 1706 823 1712 824
rect 1706 819 1707 823
rect 1711 819 1712 823
rect 1706 818 1712 819
rect 1784 811 1786 836
rect 2006 835 2012 836
rect 2046 840 2052 841
rect 2046 836 2047 840
rect 2051 836 2052 840
rect 2342 837 2343 841
rect 2347 837 2348 841
rect 2342 836 2348 837
rect 2046 835 2052 836
rect 2008 811 2010 835
rect 2048 815 2050 835
rect 2344 815 2346 836
rect 2432 824 2434 846
rect 2438 841 2444 842
rect 2438 837 2439 841
rect 2443 837 2444 841
rect 2438 836 2444 837
rect 2430 823 2436 824
rect 2430 819 2431 823
rect 2435 819 2436 823
rect 2430 818 2436 819
rect 2440 815 2442 836
rect 2528 824 2530 846
rect 2534 841 2540 842
rect 2534 837 2535 841
rect 2539 837 2540 841
rect 2534 836 2540 837
rect 2630 841 2636 842
rect 2630 837 2631 841
rect 2635 837 2636 841
rect 2630 836 2636 837
rect 2526 823 2532 824
rect 2526 819 2527 823
rect 2531 819 2532 823
rect 2526 818 2532 819
rect 2536 815 2538 836
rect 2632 815 2634 836
rect 2692 824 2694 922
rect 2710 920 2716 921
rect 2710 916 2711 920
rect 2715 916 2716 920
rect 2710 915 2716 916
rect 2822 920 2828 921
rect 2822 916 2823 920
rect 2827 916 2828 920
rect 2822 915 2828 916
rect 2950 920 2956 921
rect 2950 916 2951 920
rect 2955 916 2956 920
rect 2950 915 2956 916
rect 3102 920 3108 921
rect 3102 916 3103 920
rect 3107 916 3108 920
rect 3102 915 3108 916
rect 3270 920 3276 921
rect 3270 916 3271 920
rect 3275 916 3276 920
rect 3270 915 3276 916
rect 2712 891 2714 915
rect 2824 891 2826 915
rect 2952 891 2954 915
rect 3104 891 3106 915
rect 3272 891 3274 915
rect 2711 890 2715 891
rect 2711 885 2715 886
rect 2735 890 2739 891
rect 2735 885 2739 886
rect 2823 890 2827 891
rect 2823 885 2827 886
rect 2863 890 2867 891
rect 2863 885 2867 886
rect 2951 890 2955 891
rect 2951 885 2955 886
rect 3015 890 3019 891
rect 3015 885 3019 886
rect 3103 890 3107 891
rect 3103 885 3107 886
rect 3191 890 3195 891
rect 3191 885 3195 886
rect 3271 890 3275 891
rect 3271 885 3275 886
rect 3391 890 3395 891
rect 3391 885 3395 886
rect 2736 861 2738 885
rect 2864 861 2866 885
rect 3016 861 3018 885
rect 3192 861 3194 885
rect 3392 861 3394 885
rect 2734 860 2740 861
rect 2734 856 2735 860
rect 2739 856 2740 860
rect 2734 855 2740 856
rect 2862 860 2868 861
rect 2862 856 2863 860
rect 2867 856 2868 860
rect 2862 855 2868 856
rect 3014 860 3020 861
rect 3014 856 3015 860
rect 3019 856 3020 860
rect 3014 855 3020 856
rect 3190 860 3196 861
rect 3190 856 3191 860
rect 3195 856 3196 860
rect 3190 855 3196 856
rect 3390 860 3396 861
rect 3390 856 3391 860
rect 3395 856 3396 860
rect 3390 855 3396 856
rect 2706 851 2712 852
rect 2706 847 2707 851
rect 2711 847 2712 851
rect 2706 846 2712 847
rect 2714 851 2720 852
rect 2714 847 2715 851
rect 2719 847 2720 851
rect 2714 846 2720 847
rect 2938 851 2944 852
rect 2938 847 2939 851
rect 2943 847 2944 851
rect 2938 846 2944 847
rect 3090 851 3096 852
rect 3090 847 3091 851
rect 3095 847 3096 851
rect 3090 846 3096 847
rect 3266 851 3272 852
rect 3266 847 3267 851
rect 3271 847 3272 851
rect 3266 846 3272 847
rect 2708 824 2710 846
rect 2716 832 2718 846
rect 2734 841 2740 842
rect 2734 837 2735 841
rect 2739 837 2740 841
rect 2734 836 2740 837
rect 2862 841 2868 842
rect 2862 837 2863 841
rect 2867 837 2868 841
rect 2862 836 2868 837
rect 2714 831 2720 832
rect 2714 827 2715 831
rect 2719 827 2720 831
rect 2714 826 2720 827
rect 2690 823 2696 824
rect 2690 819 2691 823
rect 2695 819 2696 823
rect 2690 818 2696 819
rect 2706 823 2712 824
rect 2706 819 2707 823
rect 2711 819 2712 823
rect 2706 818 2712 819
rect 2736 815 2738 836
rect 2864 815 2866 836
rect 2940 824 2942 846
rect 3014 841 3020 842
rect 3014 837 3015 841
rect 3019 837 3020 841
rect 3014 836 3020 837
rect 2938 823 2944 824
rect 2938 819 2939 823
rect 2943 819 2944 823
rect 2938 818 2944 819
rect 3016 815 3018 836
rect 3092 824 3094 846
rect 3190 841 3196 842
rect 3190 837 3191 841
rect 3195 837 3196 841
rect 3190 836 3196 837
rect 3090 823 3096 824
rect 3090 819 3091 823
rect 3095 819 3096 823
rect 3090 818 3096 819
rect 3192 815 3194 836
rect 3268 824 3270 846
rect 3390 841 3396 842
rect 3390 837 3391 841
rect 3395 837 3396 841
rect 3390 836 3396 837
rect 3266 823 3272 824
rect 3266 819 3267 823
rect 3271 819 3272 823
rect 3266 818 3272 819
rect 3392 815 3394 836
rect 3412 832 3414 926
rect 3454 920 3460 921
rect 3454 916 3455 920
rect 3459 916 3460 920
rect 3454 915 3460 916
rect 3646 920 3652 921
rect 3646 916 3647 920
rect 3651 916 3652 920
rect 3646 915 3652 916
rect 3456 891 3458 915
rect 3648 891 3650 915
rect 3455 890 3459 891
rect 3455 885 3459 886
rect 3607 890 3611 891
rect 3607 885 3611 886
rect 3647 890 3651 891
rect 3647 885 3651 886
rect 3608 861 3610 885
rect 3606 860 3612 861
rect 3606 856 3607 860
rect 3611 856 3612 860
rect 3606 855 3612 856
rect 3466 851 3472 852
rect 3466 847 3467 851
rect 3471 847 3472 851
rect 3466 846 3472 847
rect 3474 851 3480 852
rect 3474 847 3475 851
rect 3479 847 3480 851
rect 3474 846 3480 847
rect 3410 831 3416 832
rect 3410 827 3411 831
rect 3415 827 3416 831
rect 3410 826 3416 827
rect 3468 824 3470 846
rect 3466 823 3472 824
rect 3466 819 3467 823
rect 3471 819 3472 823
rect 3466 818 3472 819
rect 3476 816 3478 846
rect 3606 841 3612 842
rect 3606 837 3607 841
rect 3611 837 3612 841
rect 3606 836 3612 837
rect 3474 815 3480 816
rect 3608 815 3610 836
rect 2047 814 2051 815
rect 623 810 627 811
rect 623 805 627 806
rect 639 810 643 811
rect 639 805 643 806
rect 775 810 779 811
rect 775 805 779 806
rect 823 810 827 811
rect 823 805 827 806
rect 935 810 939 811
rect 935 805 939 806
rect 999 810 1003 811
rect 999 805 1003 806
rect 1095 810 1099 811
rect 1095 805 1099 806
rect 1167 810 1171 811
rect 1167 805 1171 806
rect 1255 810 1259 811
rect 1255 805 1259 806
rect 1327 810 1331 811
rect 1327 805 1331 806
rect 1415 810 1419 811
rect 1415 805 1419 806
rect 1479 810 1483 811
rect 1518 810 1524 811
rect 1583 810 1587 811
rect 1479 805 1483 806
rect 510 803 518 804
rect 510 799 511 803
rect 515 800 518 803
rect 546 803 552 804
rect 515 799 516 800
rect 510 798 516 799
rect 546 799 547 803
rect 551 799 552 803
rect 546 798 552 799
rect 470 783 476 784
rect 470 779 471 783
rect 475 779 476 783
rect 470 778 476 779
rect 548 776 550 798
rect 624 784 626 805
rect 698 803 704 804
rect 698 799 699 803
rect 703 799 704 803
rect 698 798 704 799
rect 622 783 628 784
rect 622 779 623 783
rect 627 779 628 783
rect 622 778 628 779
rect 700 776 702 798
rect 776 784 778 805
rect 936 784 938 805
rect 974 803 980 804
rect 974 799 975 803
rect 979 799 980 803
rect 974 798 980 799
rect 1010 803 1016 804
rect 1010 799 1011 803
rect 1015 799 1016 803
rect 1010 798 1016 799
rect 774 783 780 784
rect 774 779 775 783
rect 779 779 780 783
rect 774 778 780 779
rect 934 783 940 784
rect 934 779 935 783
rect 939 779 940 783
rect 934 778 940 779
rect 546 775 552 776
rect 546 771 547 775
rect 551 771 552 775
rect 546 770 552 771
rect 698 775 704 776
rect 698 771 699 775
rect 703 771 704 775
rect 698 770 704 771
rect 850 771 856 772
rect 850 767 851 771
rect 855 767 856 771
rect 850 766 856 767
rect 470 764 476 765
rect 470 760 471 764
rect 475 760 476 764
rect 470 759 476 760
rect 622 764 628 765
rect 622 760 623 764
rect 627 760 628 764
rect 622 759 628 760
rect 774 764 780 765
rect 774 760 775 764
rect 779 760 780 764
rect 774 759 780 760
rect 472 735 474 759
rect 624 735 626 759
rect 776 735 778 759
rect 431 734 435 735
rect 431 729 435 730
rect 471 734 475 735
rect 471 729 475 730
rect 623 734 627 735
rect 623 729 627 730
rect 775 734 779 735
rect 775 729 779 730
rect 823 734 827 735
rect 823 729 827 730
rect 432 705 434 729
rect 624 705 626 729
rect 824 705 826 729
rect 430 704 436 705
rect 430 700 431 704
rect 435 700 436 704
rect 430 699 436 700
rect 622 704 628 705
rect 622 700 623 704
rect 627 700 628 704
rect 622 699 628 700
rect 822 704 828 705
rect 822 700 823 704
rect 827 700 828 704
rect 822 699 828 700
rect 210 695 216 696
rect 210 691 211 695
rect 215 691 216 695
rect 210 690 216 691
rect 338 695 344 696
rect 338 691 339 695
rect 343 691 344 695
rect 338 690 344 691
rect 422 695 428 696
rect 422 691 423 695
rect 427 691 428 695
rect 422 690 428 691
rect 542 695 548 696
rect 542 691 543 695
rect 547 691 548 695
rect 542 690 548 691
rect 706 695 712 696
rect 706 691 707 695
rect 711 691 712 695
rect 706 690 712 691
rect 134 685 140 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 134 681 135 685
rect 139 681 140 685
rect 134 680 140 681
rect 110 679 116 680
rect 112 659 114 679
rect 136 659 138 680
rect 212 668 214 690
rect 262 685 268 686
rect 262 681 263 685
rect 267 681 268 685
rect 262 680 268 681
rect 210 667 216 668
rect 210 663 211 667
rect 215 663 216 667
rect 210 662 216 663
rect 210 659 216 660
rect 264 659 266 680
rect 111 658 115 659
rect 111 653 115 654
rect 135 658 139 659
rect 210 655 211 659
rect 215 655 216 659
rect 210 654 216 655
rect 247 658 251 659
rect 135 653 139 654
rect 112 633 114 653
rect 110 632 116 633
rect 136 632 138 653
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 134 631 140 632
rect 134 627 135 631
rect 139 627 140 631
rect 134 626 140 627
rect 212 624 214 654
rect 247 653 251 654
rect 263 658 267 659
rect 263 653 267 654
rect 383 658 387 659
rect 383 653 387 654
rect 218 651 224 652
rect 218 647 219 651
rect 223 647 224 651
rect 218 646 224 647
rect 220 624 222 646
rect 248 632 250 653
rect 286 651 292 652
rect 286 647 287 651
rect 291 647 292 651
rect 286 646 292 647
rect 246 631 252 632
rect 246 627 247 631
rect 251 627 252 631
rect 246 626 252 627
rect 210 623 216 624
rect 210 619 211 623
rect 215 619 216 623
rect 210 618 216 619
rect 218 623 224 624
rect 218 619 219 623
rect 223 619 224 623
rect 218 618 224 619
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 110 610 116 611
rect 134 612 140 613
rect 112 579 114 610
rect 134 608 135 612
rect 139 608 140 612
rect 134 607 140 608
rect 246 612 252 613
rect 246 608 247 612
rect 251 608 252 612
rect 246 607 252 608
rect 136 579 138 607
rect 248 579 250 607
rect 111 578 115 579
rect 111 573 115 574
rect 135 578 139 579
rect 135 573 139 574
rect 247 578 251 579
rect 247 573 251 574
rect 112 546 114 573
rect 136 549 138 573
rect 134 548 140 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 134 544 135 548
rect 139 544 140 548
rect 134 543 140 544
rect 110 540 116 541
rect 288 540 290 646
rect 384 632 386 653
rect 424 652 426 690
rect 430 685 436 686
rect 430 681 431 685
rect 435 681 436 685
rect 430 680 436 681
rect 432 659 434 680
rect 544 668 546 690
rect 622 685 628 686
rect 622 681 623 685
rect 627 681 628 685
rect 622 680 628 681
rect 542 667 548 668
rect 542 663 543 667
rect 547 663 548 667
rect 542 662 548 663
rect 624 659 626 680
rect 708 668 710 690
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 706 667 712 668
rect 706 663 707 667
rect 711 663 712 667
rect 706 662 712 663
rect 824 659 826 680
rect 852 668 854 766
rect 934 764 940 765
rect 934 760 935 764
rect 939 760 940 764
rect 934 759 940 760
rect 936 735 938 759
rect 935 734 939 735
rect 935 729 939 730
rect 976 696 978 798
rect 1012 776 1014 798
rect 1096 784 1098 805
rect 1230 803 1236 804
rect 1230 799 1231 803
rect 1235 799 1236 803
rect 1230 798 1236 799
rect 1094 783 1100 784
rect 1094 779 1095 783
rect 1099 779 1100 783
rect 1094 778 1100 779
rect 1232 776 1234 798
rect 1256 784 1258 805
rect 1374 803 1380 804
rect 1374 799 1375 803
rect 1379 799 1380 803
rect 1374 798 1380 799
rect 1254 783 1260 784
rect 1254 779 1255 783
rect 1259 779 1260 783
rect 1254 778 1260 779
rect 1376 776 1378 798
rect 1416 784 1418 805
rect 1490 803 1496 804
rect 1490 799 1491 803
rect 1495 799 1496 803
rect 1490 798 1496 799
rect 1414 783 1420 784
rect 1414 779 1415 783
rect 1419 779 1420 783
rect 1414 778 1420 779
rect 1492 776 1494 798
rect 1520 776 1522 810
rect 1583 805 1587 806
rect 1631 810 1635 811
rect 1631 805 1635 806
rect 1751 810 1755 811
rect 1751 805 1755 806
rect 1783 810 1787 811
rect 1783 805 1787 806
rect 1903 810 1907 811
rect 1903 805 1907 806
rect 2007 810 2011 811
rect 2047 809 2051 810
rect 2311 814 2315 815
rect 2311 809 2315 810
rect 2343 814 2347 815
rect 2343 809 2347 810
rect 2439 814 2443 815
rect 2439 809 2443 810
rect 2495 814 2499 815
rect 2495 809 2499 810
rect 2535 814 2539 815
rect 2535 809 2539 810
rect 2631 814 2635 815
rect 2631 809 2635 810
rect 2687 814 2691 815
rect 2687 809 2691 810
rect 2735 814 2739 815
rect 2735 809 2739 810
rect 2863 814 2867 815
rect 2863 809 2867 810
rect 2879 814 2883 815
rect 2879 809 2883 810
rect 3015 814 3019 815
rect 3015 809 3019 810
rect 3079 814 3083 815
rect 3079 809 3083 810
rect 3191 814 3195 815
rect 3191 809 3195 810
rect 3287 814 3291 815
rect 3287 809 3291 810
rect 3391 814 3395 815
rect 3474 811 3475 815
rect 3479 811 3480 815
rect 3474 810 3480 811
rect 3503 814 3507 815
rect 3391 809 3395 810
rect 3503 809 3507 810
rect 3607 814 3611 815
rect 3607 809 3611 810
rect 2007 805 2011 806
rect 1584 784 1586 805
rect 1752 784 1754 805
rect 1834 803 1840 804
rect 1834 799 1835 803
rect 1839 799 1840 803
rect 1834 798 1840 799
rect 1582 783 1588 784
rect 1582 779 1583 783
rect 1587 779 1588 783
rect 1582 778 1588 779
rect 1750 783 1756 784
rect 1750 779 1751 783
rect 1755 779 1756 783
rect 1750 778 1756 779
rect 1836 776 1838 798
rect 1904 784 1906 805
rect 1986 803 1992 804
rect 1986 799 1987 803
rect 1991 799 1992 803
rect 1986 798 1992 799
rect 1902 783 1908 784
rect 1902 779 1903 783
rect 1907 779 1908 783
rect 1902 778 1908 779
rect 1010 775 1016 776
rect 1010 771 1011 775
rect 1015 771 1016 775
rect 1010 770 1016 771
rect 1230 775 1236 776
rect 1230 771 1231 775
rect 1235 771 1236 775
rect 1230 770 1236 771
rect 1374 775 1380 776
rect 1374 771 1375 775
rect 1379 771 1380 775
rect 1374 770 1380 771
rect 1490 775 1496 776
rect 1490 771 1491 775
rect 1495 771 1496 775
rect 1490 770 1496 771
rect 1518 775 1524 776
rect 1518 771 1519 775
rect 1523 771 1524 775
rect 1834 775 1840 776
rect 1518 770 1524 771
rect 1826 771 1832 772
rect 1826 767 1827 771
rect 1831 767 1832 771
rect 1834 771 1835 775
rect 1839 771 1840 775
rect 1834 770 1840 771
rect 1826 766 1832 767
rect 1094 764 1100 765
rect 1094 760 1095 764
rect 1099 760 1100 764
rect 1094 759 1100 760
rect 1254 764 1260 765
rect 1254 760 1255 764
rect 1259 760 1260 764
rect 1254 759 1260 760
rect 1414 764 1420 765
rect 1414 760 1415 764
rect 1419 760 1420 764
rect 1414 759 1420 760
rect 1582 764 1588 765
rect 1582 760 1583 764
rect 1587 760 1588 764
rect 1582 759 1588 760
rect 1750 764 1756 765
rect 1750 760 1751 764
rect 1755 760 1756 764
rect 1750 759 1756 760
rect 1096 735 1098 759
rect 1256 735 1258 759
rect 1416 735 1418 759
rect 1584 735 1586 759
rect 1752 735 1754 759
rect 1015 734 1019 735
rect 1015 729 1019 730
rect 1095 734 1099 735
rect 1095 729 1099 730
rect 1207 734 1211 735
rect 1207 729 1211 730
rect 1255 734 1259 735
rect 1255 729 1259 730
rect 1391 734 1395 735
rect 1391 729 1395 730
rect 1415 734 1419 735
rect 1415 729 1419 730
rect 1567 734 1571 735
rect 1567 729 1571 730
rect 1583 734 1587 735
rect 1583 729 1587 730
rect 1743 734 1747 735
rect 1743 729 1747 730
rect 1751 734 1755 735
rect 1751 729 1755 730
rect 1016 705 1018 729
rect 1208 705 1210 729
rect 1392 705 1394 729
rect 1568 705 1570 729
rect 1744 705 1746 729
rect 1014 704 1020 705
rect 1014 700 1015 704
rect 1019 700 1020 704
rect 1014 699 1020 700
rect 1206 704 1212 705
rect 1206 700 1207 704
rect 1211 700 1212 704
rect 1206 699 1212 700
rect 1390 704 1396 705
rect 1390 700 1391 704
rect 1395 700 1396 704
rect 1390 699 1396 700
rect 1566 704 1572 705
rect 1566 700 1567 704
rect 1571 700 1572 704
rect 1566 699 1572 700
rect 1742 704 1748 705
rect 1742 700 1743 704
rect 1747 700 1748 704
rect 1742 699 1748 700
rect 974 695 980 696
rect 974 691 975 695
rect 979 691 980 695
rect 974 690 980 691
rect 1466 695 1472 696
rect 1466 691 1467 695
rect 1471 691 1472 695
rect 1466 690 1472 691
rect 1642 695 1648 696
rect 1642 691 1643 695
rect 1647 691 1648 695
rect 1642 690 1648 691
rect 1650 695 1656 696
rect 1650 691 1651 695
rect 1655 691 1656 695
rect 1650 690 1656 691
rect 1014 685 1020 686
rect 1014 681 1015 685
rect 1019 681 1020 685
rect 1014 680 1020 681
rect 1206 685 1212 686
rect 1206 681 1207 685
rect 1211 681 1212 685
rect 1206 680 1212 681
rect 1390 685 1396 686
rect 1390 681 1391 685
rect 1395 681 1396 685
rect 1390 680 1396 681
rect 850 667 856 668
rect 850 663 851 667
rect 855 663 856 667
rect 850 662 856 663
rect 1016 659 1018 680
rect 1208 659 1210 680
rect 1392 659 1394 680
rect 1468 668 1470 690
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 1466 667 1472 668
rect 1466 663 1467 667
rect 1471 663 1472 667
rect 1466 662 1472 663
rect 1568 659 1570 680
rect 431 658 435 659
rect 431 653 435 654
rect 527 658 531 659
rect 527 653 531 654
rect 623 658 627 659
rect 623 653 627 654
rect 687 658 691 659
rect 687 653 691 654
rect 823 658 827 659
rect 823 653 827 654
rect 871 658 875 659
rect 871 653 875 654
rect 1015 658 1019 659
rect 1015 653 1019 654
rect 1079 658 1083 659
rect 1079 653 1083 654
rect 1207 658 1211 659
rect 1207 653 1211 654
rect 1303 658 1307 659
rect 1303 653 1307 654
rect 1391 658 1395 659
rect 1391 653 1395 654
rect 1543 658 1547 659
rect 1543 653 1547 654
rect 1567 658 1571 659
rect 1567 653 1571 654
rect 422 651 428 652
rect 422 647 423 651
rect 427 647 428 651
rect 422 646 428 647
rect 458 651 464 652
rect 458 647 459 651
rect 463 647 464 651
rect 458 646 464 647
rect 382 631 388 632
rect 382 627 383 631
rect 387 627 388 631
rect 382 626 388 627
rect 460 624 462 646
rect 528 632 530 653
rect 602 651 608 652
rect 602 647 603 651
rect 607 647 608 651
rect 602 646 608 647
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 604 624 606 646
rect 688 632 690 653
rect 872 632 874 653
rect 910 651 916 652
rect 910 647 911 651
rect 915 650 916 651
rect 946 651 952 652
rect 915 647 918 650
rect 910 646 918 647
rect 946 647 947 651
rect 951 647 952 651
rect 946 646 952 647
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 870 631 876 632
rect 870 627 871 631
rect 875 627 876 631
rect 870 626 876 627
rect 458 623 464 624
rect 458 619 459 623
rect 463 619 464 623
rect 458 618 464 619
rect 602 623 608 624
rect 602 619 603 623
rect 607 619 608 623
rect 602 618 608 619
rect 762 619 768 620
rect 762 615 763 619
rect 767 615 768 619
rect 762 614 768 615
rect 382 612 388 613
rect 382 608 383 612
rect 387 608 388 612
rect 382 607 388 608
rect 526 612 532 613
rect 526 608 527 612
rect 531 608 532 612
rect 526 607 532 608
rect 686 612 692 613
rect 686 608 687 612
rect 691 608 692 612
rect 686 607 692 608
rect 384 579 386 607
rect 528 579 530 607
rect 688 579 690 607
rect 295 578 299 579
rect 295 573 299 574
rect 383 578 387 579
rect 383 573 387 574
rect 479 578 483 579
rect 479 573 483 574
rect 527 578 531 579
rect 527 573 531 574
rect 663 578 667 579
rect 663 573 667 574
rect 687 578 691 579
rect 687 573 691 574
rect 296 549 298 573
rect 480 549 482 573
rect 664 549 666 573
rect 294 548 300 549
rect 294 544 295 548
rect 299 544 300 548
rect 294 543 300 544
rect 478 548 484 549
rect 478 544 479 548
rect 483 544 484 548
rect 478 543 484 544
rect 662 548 668 549
rect 662 544 663 548
rect 667 544 668 548
rect 662 543 668 544
rect 230 539 236 540
rect 230 535 231 539
rect 235 535 236 539
rect 230 534 236 535
rect 286 539 292 540
rect 286 535 287 539
rect 291 535 292 539
rect 286 534 292 535
rect 134 529 140 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 134 525 135 529
rect 139 525 140 529
rect 134 524 140 525
rect 110 523 116 524
rect 112 503 114 523
rect 136 503 138 524
rect 232 512 234 534
rect 294 529 300 530
rect 294 525 295 529
rect 299 525 300 529
rect 294 524 300 525
rect 478 529 484 530
rect 478 525 479 529
rect 483 525 484 529
rect 478 524 484 525
rect 662 529 668 530
rect 662 525 663 529
rect 667 525 668 529
rect 662 524 668 525
rect 230 511 236 512
rect 210 507 216 508
rect 210 503 211 507
rect 215 503 216 507
rect 230 507 231 511
rect 235 507 236 511
rect 230 506 236 507
rect 296 503 298 524
rect 480 503 482 524
rect 664 503 666 524
rect 764 512 766 614
rect 870 612 876 613
rect 870 608 871 612
rect 875 608 876 612
rect 870 607 876 608
rect 872 579 874 607
rect 847 578 851 579
rect 847 573 851 574
rect 871 578 875 579
rect 871 573 875 574
rect 848 549 850 573
rect 846 548 852 549
rect 846 544 847 548
rect 851 544 852 548
rect 846 543 852 544
rect 916 540 918 646
rect 948 624 950 646
rect 1080 632 1082 653
rect 1154 651 1160 652
rect 1154 647 1155 651
rect 1159 647 1160 651
rect 1154 646 1160 647
rect 1078 631 1084 632
rect 1078 627 1079 631
rect 1083 627 1084 631
rect 1078 626 1084 627
rect 1156 624 1158 646
rect 1304 632 1306 653
rect 1378 651 1384 652
rect 1378 647 1379 651
rect 1383 647 1384 651
rect 1378 646 1384 647
rect 1302 631 1308 632
rect 1302 627 1303 631
rect 1307 627 1308 631
rect 1302 626 1308 627
rect 1380 624 1382 646
rect 1544 632 1546 653
rect 1644 652 1646 690
rect 1652 676 1654 690
rect 1810 687 1816 688
rect 1742 685 1748 686
rect 1742 681 1743 685
rect 1747 681 1748 685
rect 1810 683 1811 687
rect 1815 683 1816 687
rect 1810 682 1816 683
rect 1742 680 1748 681
rect 1650 675 1656 676
rect 1650 671 1651 675
rect 1655 671 1656 675
rect 1650 670 1656 671
rect 1744 659 1746 680
rect 1812 668 1814 682
rect 1828 668 1830 766
rect 1902 764 1908 765
rect 1902 760 1903 764
rect 1907 760 1908 764
rect 1902 759 1908 760
rect 1904 735 1906 759
rect 1903 734 1907 735
rect 1903 729 1907 730
rect 1904 705 1906 729
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 1902 699 1908 700
rect 1988 696 1990 798
rect 2008 785 2010 805
rect 2048 789 2050 809
rect 2046 788 2052 789
rect 2312 788 2314 809
rect 2386 807 2392 808
rect 2386 803 2387 807
rect 2391 803 2392 807
rect 2386 802 2392 803
rect 2006 784 2012 785
rect 2006 780 2007 784
rect 2011 780 2012 784
rect 2046 784 2047 788
rect 2051 784 2052 788
rect 2046 783 2052 784
rect 2310 787 2316 788
rect 2310 783 2311 787
rect 2315 783 2316 787
rect 2310 782 2316 783
rect 2388 780 2390 802
rect 2496 788 2498 809
rect 2570 807 2576 808
rect 2570 803 2571 807
rect 2575 803 2576 807
rect 2570 802 2576 803
rect 2494 787 2500 788
rect 2494 783 2495 787
rect 2499 783 2500 787
rect 2494 782 2500 783
rect 2572 780 2574 802
rect 2688 788 2690 809
rect 2880 788 2882 809
rect 2954 807 2960 808
rect 2954 803 2955 807
rect 2959 803 2960 807
rect 2954 802 2960 803
rect 2686 787 2692 788
rect 2686 783 2687 787
rect 2691 783 2692 787
rect 2686 782 2692 783
rect 2878 787 2884 788
rect 2878 783 2879 787
rect 2883 783 2884 787
rect 2878 782 2884 783
rect 2956 780 2958 802
rect 3080 788 3082 809
rect 3154 807 3160 808
rect 3154 803 3155 807
rect 3159 803 3160 807
rect 3154 802 3160 803
rect 3078 787 3084 788
rect 3078 783 3079 787
rect 3083 783 3084 787
rect 3078 782 3084 783
rect 3156 780 3158 802
rect 3288 788 3290 809
rect 3362 807 3368 808
rect 3362 803 3363 807
rect 3367 803 3368 807
rect 3362 802 3368 803
rect 3286 787 3292 788
rect 3286 783 3287 787
rect 3291 783 3292 787
rect 3286 782 3292 783
rect 3364 780 3366 802
rect 3504 788 3506 809
rect 3502 787 3508 788
rect 3502 783 3503 787
rect 3507 783 3508 787
rect 3502 782 3508 783
rect 3688 780 3690 954
rect 3724 932 3726 970
rect 3840 967 3842 992
rect 3839 966 3843 967
rect 3839 961 3843 962
rect 3840 940 3842 961
rect 3908 960 3910 1002
rect 3916 980 3918 1082
rect 3942 1079 3943 1083
rect 3947 1079 3948 1083
rect 3942 1078 3948 1079
rect 3944 1047 3946 1078
rect 3943 1046 3947 1047
rect 3943 1041 3947 1042
rect 3944 1014 3946 1041
rect 3942 1013 3948 1014
rect 3942 1009 3943 1013
rect 3947 1009 3948 1013
rect 3942 1008 3948 1009
rect 3942 996 3948 997
rect 3942 992 3943 996
rect 3947 992 3948 996
rect 3942 991 3948 992
rect 3914 979 3920 980
rect 3914 975 3915 979
rect 3919 975 3920 979
rect 3914 974 3920 975
rect 3944 967 3946 991
rect 3943 966 3947 967
rect 3943 961 3947 962
rect 3906 959 3912 960
rect 3906 955 3907 959
rect 3911 955 3912 959
rect 3906 954 3912 955
rect 3944 941 3946 961
rect 3942 940 3948 941
rect 3838 939 3844 940
rect 3838 935 3839 939
rect 3843 935 3844 939
rect 3942 936 3943 940
rect 3947 936 3948 940
rect 3942 935 3948 936
rect 3838 934 3844 935
rect 3722 931 3728 932
rect 3722 927 3723 931
rect 3727 927 3728 931
rect 3722 926 3728 927
rect 3914 927 3920 928
rect 3914 923 3915 927
rect 3919 923 3920 927
rect 3914 922 3920 923
rect 3942 923 3948 924
rect 3838 920 3844 921
rect 3838 916 3839 920
rect 3843 916 3844 920
rect 3838 915 3844 916
rect 3840 891 3842 915
rect 3823 890 3827 891
rect 3823 885 3827 886
rect 3839 890 3843 891
rect 3839 885 3843 886
rect 3824 861 3826 885
rect 3822 860 3828 861
rect 3822 856 3823 860
rect 3827 856 3828 860
rect 3822 855 3828 856
rect 3890 851 3896 852
rect 3890 847 3891 851
rect 3895 847 3896 851
rect 3890 846 3896 847
rect 3822 841 3828 842
rect 3822 837 3823 841
rect 3827 837 3828 841
rect 3822 836 3828 837
rect 3824 815 3826 836
rect 3719 814 3723 815
rect 3719 809 3723 810
rect 3823 814 3827 815
rect 3823 809 3827 810
rect 3720 788 3722 809
rect 3770 807 3776 808
rect 3770 803 3771 807
rect 3775 803 3776 807
rect 3770 802 3776 803
rect 3718 787 3724 788
rect 3718 783 3719 787
rect 3723 783 3724 787
rect 3718 782 3724 783
rect 2006 779 2012 780
rect 2386 779 2392 780
rect 2386 775 2387 779
rect 2391 775 2392 779
rect 2386 774 2392 775
rect 2570 779 2576 780
rect 2570 775 2571 779
rect 2575 775 2576 779
rect 2570 774 2576 775
rect 2954 779 2960 780
rect 2954 775 2955 779
rect 2959 775 2960 779
rect 2954 774 2960 775
rect 3154 779 3160 780
rect 3154 775 3155 779
rect 3159 775 3160 779
rect 3154 774 3160 775
rect 3362 779 3368 780
rect 3362 775 3363 779
rect 3367 775 3368 779
rect 3362 774 3368 775
rect 3446 779 3452 780
rect 3446 775 3447 779
rect 3451 775 3452 779
rect 3446 774 3452 775
rect 3686 779 3692 780
rect 3686 775 3687 779
rect 3691 775 3692 779
rect 3686 774 3692 775
rect 2046 771 2052 772
rect 2006 767 2012 768
rect 2006 763 2007 767
rect 2011 763 2012 767
rect 2046 767 2047 771
rect 2051 767 2052 771
rect 2046 766 2052 767
rect 2310 768 2316 769
rect 2006 762 2012 763
rect 2008 735 2010 762
rect 2048 735 2050 766
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2494 768 2500 769
rect 2494 764 2495 768
rect 2499 764 2500 768
rect 2494 763 2500 764
rect 2686 768 2692 769
rect 2686 764 2687 768
rect 2691 764 2692 768
rect 2686 763 2692 764
rect 2878 768 2884 769
rect 2878 764 2879 768
rect 2883 764 2884 768
rect 2878 763 2884 764
rect 3078 768 3084 769
rect 3078 764 3079 768
rect 3083 764 3084 768
rect 3078 763 3084 764
rect 3286 768 3292 769
rect 3286 764 3287 768
rect 3291 764 3292 768
rect 3286 763 3292 764
rect 2312 735 2314 763
rect 2496 735 2498 763
rect 2688 735 2690 763
rect 2880 735 2882 763
rect 3080 735 3082 763
rect 3288 735 3290 763
rect 2007 734 2011 735
rect 2007 729 2011 730
rect 2047 734 2051 735
rect 2047 729 2051 730
rect 2071 734 2075 735
rect 2071 729 2075 730
rect 2255 734 2259 735
rect 2255 729 2259 730
rect 2311 734 2315 735
rect 2311 729 2315 730
rect 2455 734 2459 735
rect 2455 729 2459 730
rect 2495 734 2499 735
rect 2495 729 2499 730
rect 2655 734 2659 735
rect 2655 729 2659 730
rect 2687 734 2691 735
rect 2687 729 2691 730
rect 2855 734 2859 735
rect 2855 729 2859 730
rect 2879 734 2883 735
rect 2879 729 2883 730
rect 3047 734 3051 735
rect 3047 729 3051 730
rect 3079 734 3083 735
rect 3079 729 3083 730
rect 3239 734 3243 735
rect 3239 729 3243 730
rect 3287 734 3291 735
rect 3287 729 3291 730
rect 3439 734 3443 735
rect 3439 729 3443 730
rect 2008 702 2010 729
rect 2048 702 2050 729
rect 2072 705 2074 729
rect 2256 705 2258 729
rect 2456 705 2458 729
rect 2656 705 2658 729
rect 2856 705 2858 729
rect 3048 705 3050 729
rect 3240 705 3242 729
rect 3440 705 3442 729
rect 2070 704 2076 705
rect 2006 701 2012 702
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2046 701 2052 702
rect 2046 697 2047 701
rect 2051 697 2052 701
rect 2070 700 2071 704
rect 2075 700 2076 704
rect 2070 699 2076 700
rect 2254 704 2260 705
rect 2254 700 2255 704
rect 2259 700 2260 704
rect 2254 699 2260 700
rect 2454 704 2460 705
rect 2454 700 2455 704
rect 2459 700 2460 704
rect 2454 699 2460 700
rect 2654 704 2660 705
rect 2654 700 2655 704
rect 2659 700 2660 704
rect 2654 699 2660 700
rect 2854 704 2860 705
rect 2854 700 2855 704
rect 2859 700 2860 704
rect 2854 699 2860 700
rect 3046 704 3052 705
rect 3046 700 3047 704
rect 3051 700 3052 704
rect 3046 699 3052 700
rect 3238 704 3244 705
rect 3238 700 3239 704
rect 3243 700 3244 704
rect 3238 699 3244 700
rect 3438 704 3444 705
rect 3438 700 3439 704
rect 3443 700 3444 704
rect 3438 699 3444 700
rect 2046 696 2052 697
rect 1986 695 1992 696
rect 1986 691 1987 695
rect 1991 691 1992 695
rect 1986 690 1992 691
rect 2338 695 2344 696
rect 2338 691 2339 695
rect 2343 691 2344 695
rect 2338 690 2344 691
rect 2730 695 2736 696
rect 2730 691 2731 695
rect 2735 691 2736 695
rect 2730 690 2736 691
rect 2930 695 2936 696
rect 2930 691 2931 695
rect 2935 691 2936 695
rect 2930 690 2936 691
rect 3122 695 3128 696
rect 3122 691 3123 695
rect 3127 691 3128 695
rect 3122 690 3128 691
rect 3314 695 3320 696
rect 3314 691 3315 695
rect 3319 691 3320 695
rect 3314 690 3320 691
rect 1902 685 1908 686
rect 2070 685 2076 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 1810 667 1816 668
rect 1810 663 1811 667
rect 1815 663 1816 667
rect 1810 662 1816 663
rect 1826 667 1832 668
rect 1826 663 1827 667
rect 1831 663 1832 667
rect 1826 662 1832 663
rect 1904 659 1906 680
rect 2006 679 2012 680
rect 2046 684 2052 685
rect 2046 680 2047 684
rect 2051 680 2052 684
rect 2070 681 2071 685
rect 2075 681 2076 685
rect 2070 680 2076 681
rect 2254 685 2260 686
rect 2254 681 2255 685
rect 2259 681 2260 685
rect 2254 680 2260 681
rect 2046 679 2052 680
rect 2008 659 2010 679
rect 2048 659 2050 679
rect 2072 659 2074 680
rect 2256 659 2258 680
rect 2340 668 2342 690
rect 2454 685 2460 686
rect 2454 681 2455 685
rect 2459 681 2460 685
rect 2454 680 2460 681
rect 2654 685 2660 686
rect 2654 681 2655 685
rect 2659 681 2660 685
rect 2654 680 2660 681
rect 2338 667 2344 668
rect 2338 663 2339 667
rect 2343 663 2344 667
rect 2338 662 2344 663
rect 2456 659 2458 680
rect 2506 663 2512 664
rect 2506 659 2507 663
rect 2511 659 2512 663
rect 2656 659 2658 680
rect 1743 658 1747 659
rect 1743 653 1747 654
rect 1783 658 1787 659
rect 1783 653 1787 654
rect 1903 658 1907 659
rect 1903 653 1907 654
rect 2007 658 2011 659
rect 2007 653 2011 654
rect 2047 658 2051 659
rect 2047 653 2051 654
rect 2071 658 2075 659
rect 2071 653 2075 654
rect 2231 658 2235 659
rect 2231 653 2235 654
rect 2255 658 2259 659
rect 2255 653 2259 654
rect 2431 658 2435 659
rect 2431 653 2435 654
rect 2455 658 2459 659
rect 2506 658 2512 659
rect 2631 658 2635 659
rect 2455 653 2459 654
rect 1642 651 1648 652
rect 1642 647 1643 651
rect 1647 647 1648 651
rect 1642 646 1648 647
rect 1784 632 1786 653
rect 2008 633 2010 653
rect 2048 633 2050 653
rect 2006 632 2012 633
rect 1542 631 1548 632
rect 1542 627 1543 631
rect 1547 627 1548 631
rect 1542 626 1548 627
rect 1782 631 1788 632
rect 1782 627 1783 631
rect 1787 627 1788 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 632 2052 633
rect 2072 632 2074 653
rect 2110 651 2116 652
rect 2110 647 2111 651
rect 2115 647 2116 651
rect 2110 646 2116 647
rect 2146 651 2152 652
rect 2146 647 2147 651
rect 2151 647 2152 651
rect 2146 646 2152 647
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2070 631 2076 632
rect 2070 627 2071 631
rect 2075 627 2076 631
rect 1782 626 1788 627
rect 2070 626 2076 627
rect 946 623 952 624
rect 946 619 947 623
rect 951 619 952 623
rect 946 618 952 619
rect 1154 623 1160 624
rect 1154 619 1155 623
rect 1159 619 1160 623
rect 1154 618 1160 619
rect 1378 623 1384 624
rect 1378 619 1379 623
rect 1383 619 1384 623
rect 1378 618 1384 619
rect 1850 615 1856 616
rect 1078 612 1084 613
rect 1078 608 1079 612
rect 1083 608 1084 612
rect 1078 607 1084 608
rect 1302 612 1308 613
rect 1302 608 1303 612
rect 1307 608 1308 612
rect 1302 607 1308 608
rect 1542 612 1548 613
rect 1542 608 1543 612
rect 1547 608 1548 612
rect 1542 607 1548 608
rect 1782 612 1788 613
rect 1782 608 1783 612
rect 1787 608 1788 612
rect 1850 611 1851 615
rect 1855 611 1856 615
rect 1850 610 1856 611
rect 2006 615 2012 616
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 615 2052 616
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 2046 610 2052 611
rect 2070 612 2076 613
rect 1782 607 1788 608
rect 1080 579 1082 607
rect 1304 579 1306 607
rect 1544 579 1546 607
rect 1784 579 1786 607
rect 1031 578 1035 579
rect 1031 573 1035 574
rect 1079 578 1083 579
rect 1079 573 1083 574
rect 1215 578 1219 579
rect 1215 573 1219 574
rect 1303 578 1307 579
rect 1303 573 1307 574
rect 1399 578 1403 579
rect 1399 573 1403 574
rect 1543 578 1547 579
rect 1543 573 1547 574
rect 1591 578 1595 579
rect 1591 573 1595 574
rect 1783 578 1787 579
rect 1783 573 1787 574
rect 1032 549 1034 573
rect 1216 549 1218 573
rect 1400 549 1402 573
rect 1592 549 1594 573
rect 1784 549 1786 573
rect 1030 548 1036 549
rect 1030 544 1031 548
rect 1035 544 1036 548
rect 1030 543 1036 544
rect 1214 548 1220 549
rect 1214 544 1215 548
rect 1219 544 1220 548
rect 1214 543 1220 544
rect 1398 548 1404 549
rect 1398 544 1399 548
rect 1403 544 1404 548
rect 1398 543 1404 544
rect 1590 548 1596 549
rect 1590 544 1591 548
rect 1595 544 1596 548
rect 1590 543 1596 544
rect 1782 548 1788 549
rect 1782 544 1783 548
rect 1787 544 1788 548
rect 1782 543 1788 544
rect 914 539 920 540
rect 914 535 915 539
rect 919 535 920 539
rect 914 534 920 535
rect 1106 539 1112 540
rect 1106 535 1107 539
rect 1111 535 1112 539
rect 1106 534 1112 535
rect 1114 539 1120 540
rect 1114 535 1115 539
rect 1119 535 1120 539
rect 1114 534 1120 535
rect 1466 539 1472 540
rect 1466 535 1467 539
rect 1471 535 1472 539
rect 1466 534 1472 535
rect 1726 539 1732 540
rect 1726 535 1727 539
rect 1731 535 1732 539
rect 1726 534 1732 535
rect 846 529 852 530
rect 846 525 847 529
rect 851 525 852 529
rect 846 524 852 525
rect 1030 529 1036 530
rect 1030 525 1031 529
rect 1035 525 1036 529
rect 1030 524 1036 525
rect 762 511 768 512
rect 762 507 763 511
rect 767 507 768 511
rect 762 506 768 507
rect 848 503 850 524
rect 978 507 984 508
rect 978 503 979 507
rect 983 503 984 507
rect 1032 503 1034 524
rect 1108 512 1110 534
rect 1116 520 1118 534
rect 1214 529 1220 530
rect 1214 525 1215 529
rect 1219 525 1220 529
rect 1214 524 1220 525
rect 1398 529 1404 530
rect 1398 525 1399 529
rect 1403 525 1404 529
rect 1398 524 1404 525
rect 1114 519 1120 520
rect 1114 515 1115 519
rect 1119 515 1120 519
rect 1114 514 1120 515
rect 1106 511 1112 512
rect 1106 507 1107 511
rect 1111 507 1112 511
rect 1106 506 1112 507
rect 1216 503 1218 524
rect 1400 503 1402 524
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 210 502 216 503
rect 287 502 291 503
rect 135 497 139 498
rect 112 477 114 497
rect 110 476 116 477
rect 136 476 138 497
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 212 468 214 502
rect 287 497 291 498
rect 295 502 299 503
rect 295 497 299 498
rect 455 502 459 503
rect 455 497 459 498
rect 479 502 483 503
rect 479 497 483 498
rect 615 502 619 503
rect 615 497 619 498
rect 663 502 667 503
rect 663 497 667 498
rect 767 502 771 503
rect 767 497 771 498
rect 847 502 851 503
rect 847 497 851 498
rect 903 502 907 503
rect 978 502 984 503
rect 1031 502 1035 503
rect 903 497 907 498
rect 246 495 252 496
rect 246 491 247 495
rect 251 491 252 495
rect 246 490 252 491
rect 248 468 250 490
rect 288 476 290 497
rect 354 495 360 496
rect 354 491 355 495
rect 359 491 360 495
rect 354 490 360 491
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 210 467 216 468
rect 210 463 211 467
rect 215 463 216 467
rect 210 462 216 463
rect 246 467 252 468
rect 246 463 247 467
rect 251 463 252 467
rect 246 462 252 463
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 110 454 116 455
rect 134 456 140 457
rect 112 427 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 136 427 138 451
rect 288 427 290 451
rect 111 426 115 427
rect 111 421 115 422
rect 135 426 139 427
rect 135 421 139 422
rect 287 426 291 427
rect 287 421 291 422
rect 112 394 114 421
rect 136 397 138 421
rect 288 397 290 421
rect 134 396 140 397
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 134 392 135 396
rect 139 392 140 396
rect 134 391 140 392
rect 286 396 292 397
rect 286 392 287 396
rect 291 392 292 396
rect 286 391 292 392
rect 110 388 116 389
rect 356 388 358 490
rect 456 476 458 497
rect 530 495 536 496
rect 530 491 531 495
rect 535 491 536 495
rect 530 490 536 491
rect 454 475 460 476
rect 454 471 455 475
rect 459 471 460 475
rect 454 470 460 471
rect 532 468 534 490
rect 616 476 618 497
rect 690 495 696 496
rect 690 491 691 495
rect 695 491 696 495
rect 690 490 696 491
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 692 468 694 490
rect 768 476 770 497
rect 904 476 906 497
rect 970 495 976 496
rect 970 491 971 495
rect 975 491 976 495
rect 970 490 976 491
rect 766 475 772 476
rect 766 471 767 475
rect 771 471 772 475
rect 766 470 772 471
rect 902 475 908 476
rect 902 471 903 475
rect 907 471 908 475
rect 902 470 908 471
rect 530 467 536 468
rect 530 463 531 467
rect 535 463 536 467
rect 530 462 536 463
rect 690 467 696 468
rect 690 463 691 467
rect 695 463 696 467
rect 690 462 696 463
rect 842 463 848 464
rect 842 459 843 463
rect 847 459 848 463
rect 842 458 848 459
rect 454 456 460 457
rect 454 452 455 456
rect 459 452 460 456
rect 454 451 460 452
rect 614 456 620 457
rect 614 452 615 456
rect 619 452 620 456
rect 614 451 620 452
rect 766 456 772 457
rect 766 452 767 456
rect 771 452 772 456
rect 766 451 772 452
rect 456 427 458 451
rect 616 427 618 451
rect 768 427 770 451
rect 447 426 451 427
rect 447 421 451 422
rect 455 426 459 427
rect 455 421 459 422
rect 599 426 603 427
rect 599 421 603 422
rect 615 426 619 427
rect 615 421 619 422
rect 751 426 755 427
rect 751 421 755 422
rect 767 426 771 427
rect 767 421 771 422
rect 448 397 450 421
rect 600 397 602 421
rect 752 397 754 421
rect 446 396 452 397
rect 446 392 447 396
rect 451 392 452 396
rect 446 391 452 392
rect 598 396 604 397
rect 598 392 599 396
rect 603 392 604 396
rect 598 391 604 392
rect 750 396 756 397
rect 750 392 751 396
rect 755 392 756 396
rect 750 391 756 392
rect 210 387 216 388
rect 210 383 211 387
rect 215 383 216 387
rect 210 382 216 383
rect 354 387 360 388
rect 354 383 355 387
rect 359 383 360 387
rect 354 382 360 383
rect 522 387 528 388
rect 522 383 523 387
rect 527 383 528 387
rect 522 382 528 383
rect 530 387 536 388
rect 530 383 531 387
rect 535 383 536 387
rect 530 382 536 383
rect 682 387 688 388
rect 682 383 683 387
rect 687 383 688 387
rect 682 382 688 383
rect 134 377 140 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 134 373 135 377
rect 139 373 140 377
rect 134 372 140 373
rect 110 371 116 372
rect 112 347 114 371
rect 136 347 138 372
rect 212 360 214 382
rect 286 377 292 378
rect 286 373 287 377
rect 291 373 292 377
rect 286 372 292 373
rect 446 377 452 378
rect 446 373 447 377
rect 451 373 452 377
rect 446 372 452 373
rect 210 359 216 360
rect 210 355 211 359
rect 215 355 216 359
rect 210 354 216 355
rect 288 347 290 372
rect 448 347 450 372
rect 111 346 115 347
rect 111 341 115 342
rect 135 346 139 347
rect 135 341 139 342
rect 159 346 163 347
rect 159 341 163 342
rect 287 346 291 347
rect 287 341 291 342
rect 351 346 355 347
rect 351 341 355 342
rect 447 346 451 347
rect 447 341 451 342
rect 112 321 114 341
rect 110 320 116 321
rect 160 320 162 341
rect 242 339 248 340
rect 242 335 243 339
rect 247 335 248 339
rect 242 334 248 335
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 158 319 164 320
rect 158 315 159 319
rect 163 315 164 319
rect 158 314 164 315
rect 244 312 246 334
rect 352 320 354 341
rect 524 340 526 382
rect 532 360 534 382
rect 598 377 604 378
rect 598 373 599 377
rect 603 373 604 377
rect 598 372 604 373
rect 530 359 536 360
rect 530 355 531 359
rect 535 355 536 359
rect 530 354 536 355
rect 600 347 602 372
rect 684 360 686 382
rect 750 377 756 378
rect 750 373 751 377
rect 755 373 756 377
rect 750 372 756 373
rect 682 359 688 360
rect 682 355 683 359
rect 687 355 688 359
rect 682 354 688 355
rect 752 347 754 372
rect 844 360 846 458
rect 902 456 908 457
rect 902 452 903 456
rect 907 452 908 456
rect 902 451 908 452
rect 904 427 906 451
rect 903 426 907 427
rect 903 421 907 422
rect 904 397 906 421
rect 902 396 908 397
rect 902 392 903 396
rect 907 392 908 396
rect 902 391 908 392
rect 972 388 974 490
rect 980 468 982 502
rect 1031 497 1035 498
rect 1159 502 1163 503
rect 1159 497 1163 498
rect 1215 502 1219 503
rect 1215 497 1219 498
rect 1287 502 1291 503
rect 1287 497 1291 498
rect 1399 502 1403 503
rect 1399 497 1403 498
rect 1415 502 1419 503
rect 1415 497 1419 498
rect 1032 476 1034 497
rect 1106 495 1112 496
rect 1106 491 1107 495
rect 1111 491 1112 495
rect 1106 490 1112 491
rect 1030 475 1036 476
rect 1030 471 1031 475
rect 1035 471 1036 475
rect 1030 470 1036 471
rect 1108 468 1110 490
rect 1160 476 1162 497
rect 1234 495 1240 496
rect 1234 491 1235 495
rect 1239 491 1240 495
rect 1234 490 1240 491
rect 1158 475 1164 476
rect 1158 471 1159 475
rect 1163 471 1164 475
rect 1158 470 1164 471
rect 1236 468 1238 490
rect 1288 476 1290 497
rect 1406 487 1412 488
rect 1406 483 1407 487
rect 1411 483 1412 487
rect 1406 482 1412 483
rect 1286 475 1292 476
rect 1286 471 1287 475
rect 1291 471 1292 475
rect 1286 470 1292 471
rect 1408 468 1410 482
rect 1416 476 1418 497
rect 1468 496 1470 534
rect 1590 529 1596 530
rect 1590 525 1591 529
rect 1595 525 1596 529
rect 1590 524 1596 525
rect 1592 503 1594 524
rect 1728 512 1730 534
rect 1782 529 1788 530
rect 1782 525 1783 529
rect 1787 525 1788 529
rect 1782 524 1788 525
rect 1726 511 1732 512
rect 1726 507 1727 511
rect 1731 507 1732 511
rect 1726 506 1732 507
rect 1784 503 1786 524
rect 1852 512 1854 610
rect 2008 579 2010 610
rect 2048 579 2050 610
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 2072 579 2074 607
rect 2007 578 2011 579
rect 2007 573 2011 574
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2008 546 2010 573
rect 2048 546 2050 573
rect 2072 549 2074 573
rect 2112 556 2114 646
rect 2148 624 2150 646
rect 2232 632 2234 653
rect 2306 651 2312 652
rect 2306 647 2307 651
rect 2311 647 2312 651
rect 2306 646 2312 647
rect 2230 631 2236 632
rect 2230 627 2231 631
rect 2235 627 2236 631
rect 2230 626 2236 627
rect 2308 624 2310 646
rect 2432 632 2434 653
rect 2430 631 2436 632
rect 2430 627 2431 631
rect 2435 627 2436 631
rect 2430 626 2436 627
rect 2508 624 2510 658
rect 2631 653 2635 654
rect 2655 658 2659 659
rect 2655 653 2659 654
rect 2632 632 2634 653
rect 2732 652 2734 690
rect 2854 685 2860 686
rect 2854 681 2855 685
rect 2859 681 2860 685
rect 2854 680 2860 681
rect 2856 659 2858 680
rect 2932 668 2934 690
rect 3046 685 3052 686
rect 3046 681 3047 685
rect 3051 681 3052 685
rect 3046 680 3052 681
rect 2930 667 2936 668
rect 2930 663 2931 667
rect 2935 663 2936 667
rect 2930 662 2936 663
rect 3048 659 3050 680
rect 3124 668 3126 690
rect 3238 685 3244 686
rect 3238 681 3239 685
rect 3243 681 3244 685
rect 3238 680 3244 681
rect 3122 667 3128 668
rect 3122 663 3123 667
rect 3127 663 3128 667
rect 3122 662 3128 663
rect 3240 659 3242 680
rect 3316 668 3318 690
rect 3438 685 3444 686
rect 3438 681 3439 685
rect 3443 681 3444 685
rect 3438 680 3444 681
rect 3314 667 3320 668
rect 3314 663 3315 667
rect 3319 663 3320 667
rect 3314 662 3320 663
rect 3440 659 3442 680
rect 3448 676 3450 774
rect 3502 768 3508 769
rect 3502 764 3503 768
rect 3507 764 3508 768
rect 3502 763 3508 764
rect 3718 768 3724 769
rect 3718 764 3719 768
rect 3723 764 3724 768
rect 3718 763 3724 764
rect 3504 735 3506 763
rect 3720 735 3722 763
rect 3503 734 3507 735
rect 3503 729 3507 730
rect 3639 734 3643 735
rect 3639 729 3643 730
rect 3719 734 3723 735
rect 3719 729 3723 730
rect 3640 705 3642 729
rect 3638 704 3644 705
rect 3638 700 3639 704
rect 3643 700 3644 704
rect 3638 699 3644 700
rect 3514 695 3520 696
rect 3514 691 3515 695
rect 3519 691 3520 695
rect 3514 690 3520 691
rect 3558 695 3564 696
rect 3558 691 3559 695
rect 3563 691 3564 695
rect 3558 690 3564 691
rect 3446 675 3452 676
rect 3446 671 3447 675
rect 3451 671 3452 675
rect 3446 670 3452 671
rect 3516 668 3518 690
rect 3514 667 3520 668
rect 3514 663 3515 667
rect 3519 663 3520 667
rect 3514 662 3520 663
rect 3560 660 3562 690
rect 3638 685 3644 686
rect 3638 681 3639 685
rect 3643 681 3644 685
rect 3638 680 3644 681
rect 3558 659 3564 660
rect 3640 659 3642 680
rect 2831 658 2835 659
rect 2831 653 2835 654
rect 2855 658 2859 659
rect 2855 653 2859 654
rect 3023 658 3027 659
rect 3023 653 3027 654
rect 3047 658 3051 659
rect 3047 653 3051 654
rect 3207 658 3211 659
rect 3207 653 3211 654
rect 3239 658 3243 659
rect 3239 653 3243 654
rect 3375 658 3379 659
rect 3375 653 3379 654
rect 3439 658 3443 659
rect 3439 653 3443 654
rect 3535 658 3539 659
rect 3558 655 3559 659
rect 3563 655 3564 659
rect 3558 654 3564 655
rect 3639 658 3643 659
rect 3535 653 3539 654
rect 3639 653 3643 654
rect 3695 658 3699 659
rect 3695 653 3699 654
rect 2722 651 2728 652
rect 2722 647 2723 651
rect 2727 647 2728 651
rect 2722 646 2728 647
rect 2730 651 2736 652
rect 2730 647 2731 651
rect 2735 647 2736 651
rect 2730 646 2736 647
rect 2630 631 2636 632
rect 2630 627 2631 631
rect 2635 627 2636 631
rect 2630 626 2636 627
rect 2724 624 2726 646
rect 2832 632 2834 653
rect 3024 632 3026 653
rect 3098 651 3104 652
rect 3098 647 3099 651
rect 3103 647 3104 651
rect 3098 646 3104 647
rect 2830 631 2836 632
rect 2830 627 2831 631
rect 2835 627 2836 631
rect 2830 626 2836 627
rect 3022 631 3028 632
rect 3022 627 3023 631
rect 3027 627 3028 631
rect 3022 626 3028 627
rect 3100 624 3102 646
rect 3208 632 3210 653
rect 3282 651 3288 652
rect 3282 647 3283 651
rect 3287 647 3288 651
rect 3282 646 3288 647
rect 3206 631 3212 632
rect 3206 627 3207 631
rect 3211 627 3212 631
rect 3206 626 3212 627
rect 3284 624 3286 646
rect 3376 632 3378 653
rect 3450 651 3456 652
rect 3450 647 3451 651
rect 3455 647 3456 651
rect 3450 646 3456 647
rect 3374 631 3380 632
rect 3374 627 3375 631
rect 3379 627 3380 631
rect 3374 626 3380 627
rect 3452 624 3454 646
rect 3536 632 3538 653
rect 3696 632 3698 653
rect 3534 631 3540 632
rect 3534 627 3535 631
rect 3539 627 3540 631
rect 3534 626 3540 627
rect 3694 631 3700 632
rect 3694 627 3695 631
rect 3699 627 3700 631
rect 3694 626 3700 627
rect 3772 624 3774 802
rect 3839 734 3843 735
rect 3839 729 3843 730
rect 3840 705 3842 729
rect 3838 704 3844 705
rect 3838 700 3839 704
rect 3843 700 3844 704
rect 3838 699 3844 700
rect 3838 685 3844 686
rect 3838 681 3839 685
rect 3843 681 3844 685
rect 3838 680 3844 681
rect 3840 659 3842 680
rect 3892 668 3894 846
rect 3916 824 3918 922
rect 3942 919 3943 923
rect 3947 919 3948 923
rect 3942 918 3948 919
rect 3944 891 3946 918
rect 3943 890 3947 891
rect 3943 885 3947 886
rect 3944 858 3946 885
rect 3942 857 3948 858
rect 3942 853 3943 857
rect 3947 853 3948 857
rect 3942 852 3948 853
rect 3942 840 3948 841
rect 3942 836 3943 840
rect 3947 836 3948 840
rect 3942 835 3948 836
rect 3914 823 3920 824
rect 3914 819 3915 823
rect 3919 819 3920 823
rect 3914 818 3920 819
rect 3944 815 3946 835
rect 3943 814 3947 815
rect 3943 809 3947 810
rect 3944 789 3946 809
rect 3942 788 3948 789
rect 3942 784 3943 788
rect 3947 784 3948 788
rect 3942 783 3948 784
rect 3942 771 3948 772
rect 3942 767 3943 771
rect 3947 767 3948 771
rect 3942 766 3948 767
rect 3944 735 3946 766
rect 3943 734 3947 735
rect 3943 729 3947 730
rect 3944 702 3946 729
rect 3942 701 3948 702
rect 3942 697 3943 701
rect 3947 697 3948 701
rect 3942 696 3948 697
rect 3906 695 3912 696
rect 3906 691 3907 695
rect 3911 691 3912 695
rect 3906 690 3912 691
rect 3890 667 3896 668
rect 3890 663 3891 667
rect 3895 663 3896 667
rect 3890 662 3896 663
rect 3839 658 3843 659
rect 3839 653 3843 654
rect 3778 651 3784 652
rect 3778 647 3779 651
rect 3783 647 3784 651
rect 3778 646 3784 647
rect 2146 623 2152 624
rect 2146 619 2147 623
rect 2151 619 2152 623
rect 2146 618 2152 619
rect 2306 623 2312 624
rect 2306 619 2307 623
rect 2311 619 2312 623
rect 2306 618 2312 619
rect 2506 623 2512 624
rect 2506 619 2507 623
rect 2511 619 2512 623
rect 2506 618 2512 619
rect 2598 623 2604 624
rect 2598 619 2599 623
rect 2603 619 2604 623
rect 2598 618 2604 619
rect 2722 623 2728 624
rect 2722 619 2723 623
rect 2727 619 2728 623
rect 2722 618 2728 619
rect 3098 623 3104 624
rect 3098 619 3099 623
rect 3103 619 3104 623
rect 3098 618 3104 619
rect 3282 623 3288 624
rect 3282 619 3283 623
rect 3287 619 3288 623
rect 3282 618 3288 619
rect 3450 623 3456 624
rect 3450 619 3451 623
rect 3455 619 3456 623
rect 3770 623 3776 624
rect 3450 618 3456 619
rect 3610 619 3616 620
rect 2230 612 2236 613
rect 2230 608 2231 612
rect 2235 608 2236 612
rect 2230 607 2236 608
rect 2430 612 2436 613
rect 2430 608 2431 612
rect 2435 608 2436 612
rect 2430 607 2436 608
rect 2232 579 2234 607
rect 2432 579 2434 607
rect 2215 578 2219 579
rect 2215 573 2219 574
rect 2231 578 2235 579
rect 2231 573 2235 574
rect 2399 578 2403 579
rect 2399 573 2403 574
rect 2431 578 2435 579
rect 2431 573 2435 574
rect 2583 578 2587 579
rect 2583 573 2587 574
rect 2110 555 2116 556
rect 2110 551 2111 555
rect 2115 551 2116 555
rect 2110 550 2116 551
rect 2216 549 2218 573
rect 2400 549 2402 573
rect 2584 549 2586 573
rect 2070 548 2076 549
rect 2006 545 2012 546
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2214 548 2220 549
rect 2214 544 2215 548
rect 2219 544 2220 548
rect 2214 543 2220 544
rect 2398 548 2404 549
rect 2398 544 2399 548
rect 2403 544 2404 548
rect 2398 543 2404 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2046 540 2052 541
rect 2138 539 2144 540
rect 2138 535 2139 539
rect 2143 535 2144 539
rect 2138 534 2144 535
rect 2530 539 2536 540
rect 2530 535 2531 539
rect 2535 535 2536 539
rect 2530 534 2536 535
rect 2070 529 2076 530
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2046 523 2052 524
rect 1850 511 1856 512
rect 1850 507 1851 511
rect 1855 507 1856 511
rect 1850 506 1856 507
rect 2008 503 2010 523
rect 1591 502 1595 503
rect 1591 497 1595 498
rect 1783 502 1787 503
rect 1783 497 1787 498
rect 2007 502 2011 503
rect 2048 499 2050 523
rect 2072 499 2074 524
rect 2007 497 2011 498
rect 2047 498 2051 499
rect 1466 495 1472 496
rect 1466 491 1467 495
rect 1471 491 1472 495
rect 1466 490 1472 491
rect 2008 477 2010 497
rect 2047 493 2051 494
rect 2071 498 2075 499
rect 2071 493 2075 494
rect 2006 476 2012 477
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2048 473 2050 493
rect 2006 471 2012 472
rect 2046 472 2052 473
rect 2072 472 2074 493
rect 2140 492 2142 534
rect 2214 529 2220 530
rect 2214 525 2215 529
rect 2219 525 2220 529
rect 2214 524 2220 525
rect 2398 529 2404 530
rect 2398 525 2399 529
rect 2403 525 2404 529
rect 2398 524 2404 525
rect 2216 499 2218 524
rect 2400 499 2402 524
rect 2532 512 2534 534
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2530 511 2536 512
rect 2530 507 2531 511
rect 2535 507 2536 511
rect 2530 506 2536 507
rect 2584 499 2586 524
rect 2600 520 2602 618
rect 3610 615 3611 619
rect 3615 615 3616 619
rect 3770 619 3771 623
rect 3775 619 3776 623
rect 3770 618 3776 619
rect 3610 614 3616 615
rect 2630 612 2636 613
rect 2630 608 2631 612
rect 2635 608 2636 612
rect 2630 607 2636 608
rect 2830 612 2836 613
rect 2830 608 2831 612
rect 2835 608 2836 612
rect 2830 607 2836 608
rect 3022 612 3028 613
rect 3022 608 3023 612
rect 3027 608 3028 612
rect 3022 607 3028 608
rect 3206 612 3212 613
rect 3206 608 3207 612
rect 3211 608 3212 612
rect 3206 607 3212 608
rect 3374 612 3380 613
rect 3374 608 3375 612
rect 3379 608 3380 612
rect 3374 607 3380 608
rect 3534 612 3540 613
rect 3534 608 3535 612
rect 3539 608 3540 612
rect 3534 607 3540 608
rect 2632 579 2634 607
rect 2832 579 2834 607
rect 3024 579 3026 607
rect 3208 579 3210 607
rect 3376 579 3378 607
rect 3536 579 3538 607
rect 2631 578 2635 579
rect 2631 573 2635 574
rect 2775 578 2779 579
rect 2775 573 2779 574
rect 2831 578 2835 579
rect 2831 573 2835 574
rect 2959 578 2963 579
rect 2959 573 2963 574
rect 3023 578 3027 579
rect 3023 573 3027 574
rect 3143 578 3147 579
rect 3143 573 3147 574
rect 3207 578 3211 579
rect 3207 573 3211 574
rect 3319 578 3323 579
rect 3319 573 3323 574
rect 3375 578 3379 579
rect 3375 573 3379 574
rect 3495 578 3499 579
rect 3495 573 3499 574
rect 3535 578 3539 579
rect 3535 573 3539 574
rect 2776 549 2778 573
rect 2960 549 2962 573
rect 3144 549 3146 573
rect 3320 549 3322 573
rect 3496 549 3498 573
rect 2774 548 2780 549
rect 2774 544 2775 548
rect 2779 544 2780 548
rect 2774 543 2780 544
rect 2958 548 2964 549
rect 2958 544 2959 548
rect 2963 544 2964 548
rect 2958 543 2964 544
rect 3142 548 3148 549
rect 3142 544 3143 548
rect 3147 544 3148 548
rect 3142 543 3148 544
rect 3318 548 3324 549
rect 3318 544 3319 548
rect 3323 544 3324 548
rect 3318 543 3324 544
rect 3494 548 3500 549
rect 3494 544 3495 548
rect 3499 544 3500 548
rect 3494 543 3500 544
rect 3034 539 3040 540
rect 3034 535 3035 539
rect 3039 535 3040 539
rect 3034 534 3040 535
rect 3230 539 3236 540
rect 3230 535 3231 539
rect 3235 535 3236 539
rect 3230 534 3236 535
rect 3238 539 3244 540
rect 3238 535 3239 539
rect 3243 535 3244 539
rect 3238 534 3244 535
rect 2774 529 2780 530
rect 2774 525 2775 529
rect 2779 525 2780 529
rect 2774 524 2780 525
rect 2958 529 2964 530
rect 2958 525 2959 529
rect 2963 525 2964 529
rect 2958 524 2964 525
rect 2598 519 2604 520
rect 2598 515 2599 519
rect 2603 515 2604 519
rect 2598 514 2604 515
rect 2776 499 2778 524
rect 2802 507 2808 508
rect 2802 503 2803 507
rect 2807 503 2808 507
rect 2802 502 2808 503
rect 2215 498 2219 499
rect 2215 493 2219 494
rect 2223 498 2227 499
rect 2223 493 2227 494
rect 2391 498 2395 499
rect 2391 493 2395 494
rect 2399 498 2403 499
rect 2399 493 2403 494
rect 2559 498 2563 499
rect 2559 493 2563 494
rect 2583 498 2587 499
rect 2583 493 2587 494
rect 2727 498 2731 499
rect 2727 493 2731 494
rect 2775 498 2779 499
rect 2775 493 2779 494
rect 2138 491 2144 492
rect 2138 487 2139 491
rect 2143 487 2144 491
rect 2138 486 2144 487
rect 2224 472 2226 493
rect 2262 491 2268 492
rect 2262 487 2263 491
rect 2267 487 2268 491
rect 2262 486 2268 487
rect 2298 491 2304 492
rect 2298 487 2299 491
rect 2303 487 2304 491
rect 2298 486 2304 487
rect 1414 470 1420 471
rect 2046 468 2047 472
rect 2051 468 2052 472
rect 978 467 984 468
rect 978 463 979 467
rect 983 463 984 467
rect 978 462 984 463
rect 1106 467 1112 468
rect 1106 463 1107 467
rect 1111 463 1112 467
rect 1106 462 1112 463
rect 1234 467 1240 468
rect 1234 463 1235 467
rect 1239 463 1240 467
rect 1406 467 1412 468
rect 2046 467 2052 468
rect 2070 471 2076 472
rect 2070 467 2071 471
rect 2075 467 2076 471
rect 1234 462 1240 463
rect 1398 463 1404 464
rect 1398 459 1399 463
rect 1403 459 1404 463
rect 1406 463 1407 467
rect 1411 463 1412 467
rect 2070 466 2076 467
rect 2222 471 2228 472
rect 2222 467 2223 471
rect 2227 467 2228 471
rect 2222 466 2228 467
rect 1406 462 1412 463
rect 2034 463 2040 464
rect 1398 458 1404 459
rect 2006 459 2012 460
rect 1030 456 1036 457
rect 1030 452 1031 456
rect 1035 452 1036 456
rect 1030 451 1036 452
rect 1158 456 1164 457
rect 1158 452 1159 456
rect 1163 452 1164 456
rect 1158 451 1164 452
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1286 451 1292 452
rect 1032 427 1034 451
rect 1160 427 1162 451
rect 1288 427 1290 451
rect 1031 426 1035 427
rect 1031 421 1035 422
rect 1079 426 1083 427
rect 1079 421 1083 422
rect 1159 426 1163 427
rect 1159 421 1163 422
rect 1271 426 1275 427
rect 1271 421 1275 422
rect 1287 426 1291 427
rect 1287 421 1291 422
rect 1080 397 1082 421
rect 1272 397 1274 421
rect 1078 396 1084 397
rect 1078 392 1079 396
rect 1083 392 1084 396
rect 1078 391 1084 392
rect 1270 396 1276 397
rect 1270 392 1271 396
rect 1275 392 1276 396
rect 1270 391 1276 392
rect 970 387 976 388
rect 970 383 971 387
rect 975 383 976 387
rect 970 382 976 383
rect 1210 387 1216 388
rect 1210 383 1211 387
rect 1215 383 1216 387
rect 1210 382 1216 383
rect 902 377 908 378
rect 902 373 903 377
rect 907 373 908 377
rect 902 372 908 373
rect 1078 377 1084 378
rect 1078 373 1079 377
rect 1083 373 1084 377
rect 1078 372 1084 373
rect 842 359 848 360
rect 842 355 843 359
rect 847 355 848 359
rect 842 354 848 355
rect 904 347 906 372
rect 1080 347 1082 372
rect 1212 360 1214 382
rect 1270 377 1276 378
rect 1270 373 1271 377
rect 1275 373 1276 377
rect 1270 372 1276 373
rect 1210 359 1216 360
rect 1210 355 1211 359
rect 1215 355 1216 359
rect 1210 354 1216 355
rect 1234 355 1240 356
rect 1234 351 1235 355
rect 1239 351 1240 355
rect 1234 350 1240 351
rect 551 346 555 347
rect 551 341 555 342
rect 599 346 603 347
rect 599 341 603 342
rect 751 346 755 347
rect 751 341 755 342
rect 759 346 763 347
rect 759 341 763 342
rect 903 346 907 347
rect 903 341 907 342
rect 959 346 963 347
rect 959 341 963 342
rect 1079 346 1083 347
rect 1079 341 1083 342
rect 1159 346 1163 347
rect 1159 341 1163 342
rect 522 339 528 340
rect 522 335 523 339
rect 527 335 528 339
rect 522 334 528 335
rect 552 320 554 341
rect 626 339 632 340
rect 626 335 627 339
rect 631 335 632 339
rect 626 334 632 335
rect 350 319 356 320
rect 350 315 351 319
rect 355 315 356 319
rect 350 314 356 315
rect 550 319 556 320
rect 550 315 551 319
rect 555 315 556 319
rect 550 314 556 315
rect 628 312 630 334
rect 760 320 762 341
rect 834 339 840 340
rect 834 335 835 339
rect 839 335 840 339
rect 834 334 840 335
rect 758 319 764 320
rect 758 315 759 319
rect 763 315 764 319
rect 758 314 764 315
rect 836 312 838 334
rect 960 320 962 341
rect 1160 320 1162 341
rect 958 319 964 320
rect 958 315 959 319
rect 963 315 964 319
rect 958 314 964 315
rect 1158 319 1164 320
rect 1158 315 1159 319
rect 1163 315 1164 319
rect 1158 314 1164 315
rect 1236 312 1238 350
rect 1272 347 1274 372
rect 1400 360 1402 458
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2034 459 2035 463
rect 2039 459 2040 463
rect 2034 458 2040 459
rect 2006 454 2012 455
rect 1414 451 1420 452
rect 1416 427 1418 451
rect 2008 427 2010 454
rect 1415 426 1419 427
rect 1415 421 1419 422
rect 1479 426 1483 427
rect 1479 421 1483 422
rect 1703 426 1707 427
rect 1703 421 1707 422
rect 1903 426 1907 427
rect 1903 421 1907 422
rect 2007 426 2011 427
rect 2007 421 2011 422
rect 1480 397 1482 421
rect 1704 397 1706 421
rect 1904 397 1906 421
rect 1478 396 1484 397
rect 1478 392 1479 396
rect 1483 392 1484 396
rect 1478 391 1484 392
rect 1702 396 1708 397
rect 1702 392 1703 396
rect 1707 392 1708 396
rect 1702 391 1708 392
rect 1902 396 1908 397
rect 1902 392 1903 396
rect 1907 392 1908 396
rect 2008 394 2010 421
rect 1902 391 1908 392
rect 2006 393 2012 394
rect 2006 389 2007 393
rect 2011 389 2012 393
rect 2006 388 2012 389
rect 1554 387 1560 388
rect 1554 383 1555 387
rect 1559 383 1560 387
rect 1554 382 1560 383
rect 1638 387 1644 388
rect 1638 383 1639 387
rect 1643 383 1644 387
rect 1638 382 1644 383
rect 1970 387 1976 388
rect 1970 383 1971 387
rect 1975 383 1976 387
rect 1970 382 1976 383
rect 1478 377 1484 378
rect 1478 373 1479 377
rect 1483 373 1484 377
rect 1478 372 1484 373
rect 1398 359 1404 360
rect 1398 355 1399 359
rect 1403 355 1404 359
rect 1398 354 1404 355
rect 1480 347 1482 372
rect 1556 360 1558 382
rect 1554 359 1560 360
rect 1554 355 1555 359
rect 1559 355 1560 359
rect 1554 354 1560 355
rect 1640 348 1642 382
rect 1702 377 1708 378
rect 1702 373 1703 377
rect 1707 373 1708 377
rect 1702 372 1708 373
rect 1902 377 1908 378
rect 1902 373 1903 377
rect 1907 373 1908 377
rect 1902 372 1908 373
rect 1638 347 1644 348
rect 1704 347 1706 372
rect 1904 347 1906 372
rect 1271 346 1275 347
rect 1271 341 1275 342
rect 1343 346 1347 347
rect 1343 341 1347 342
rect 1479 346 1483 347
rect 1479 341 1483 342
rect 1527 346 1531 347
rect 1638 343 1639 347
rect 1643 343 1644 347
rect 1638 342 1644 343
rect 1703 346 1707 347
rect 1527 341 1531 342
rect 1703 341 1707 342
rect 1711 346 1715 347
rect 1711 341 1715 342
rect 1895 346 1899 347
rect 1895 341 1899 342
rect 1903 346 1907 347
rect 1903 341 1907 342
rect 1344 320 1346 341
rect 1418 339 1424 340
rect 1418 335 1419 339
rect 1423 335 1424 339
rect 1418 334 1424 335
rect 1342 319 1348 320
rect 1342 315 1343 319
rect 1347 315 1348 319
rect 1342 314 1348 315
rect 1420 312 1422 334
rect 1528 320 1530 341
rect 1602 339 1608 340
rect 1602 335 1603 339
rect 1607 335 1608 339
rect 1602 334 1608 335
rect 1526 319 1532 320
rect 1526 315 1527 319
rect 1531 315 1532 319
rect 1526 314 1532 315
rect 1604 312 1606 334
rect 1712 320 1714 341
rect 1818 331 1824 332
rect 1818 327 1819 331
rect 1823 327 1824 331
rect 1818 326 1824 327
rect 1710 319 1716 320
rect 1710 315 1711 319
rect 1715 315 1716 319
rect 1710 314 1716 315
rect 1820 312 1822 326
rect 1896 320 1898 341
rect 1972 340 1974 382
rect 2006 376 2012 377
rect 2006 372 2007 376
rect 2011 372 2012 376
rect 2006 371 2012 372
rect 2008 347 2010 371
rect 2036 360 2038 458
rect 2046 455 2052 456
rect 2046 451 2047 455
rect 2051 451 2052 455
rect 2046 450 2052 451
rect 2070 452 2076 453
rect 2048 423 2050 450
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 2222 452 2228 453
rect 2222 448 2223 452
rect 2227 448 2228 452
rect 2222 447 2228 448
rect 2072 423 2074 447
rect 2224 423 2226 447
rect 2047 422 2051 423
rect 2047 417 2051 418
rect 2071 422 2075 423
rect 2071 417 2075 418
rect 2223 422 2227 423
rect 2223 417 2227 418
rect 2048 390 2050 417
rect 2046 389 2052 390
rect 2046 385 2047 389
rect 2051 385 2052 389
rect 2046 384 2052 385
rect 2264 384 2266 486
rect 2300 464 2302 486
rect 2392 472 2394 493
rect 2466 491 2472 492
rect 2466 487 2467 491
rect 2471 487 2472 491
rect 2466 486 2472 487
rect 2390 471 2396 472
rect 2390 467 2391 471
rect 2395 467 2396 471
rect 2390 466 2396 467
rect 2468 464 2470 486
rect 2560 472 2562 493
rect 2634 491 2640 492
rect 2634 487 2635 491
rect 2639 487 2640 491
rect 2634 486 2640 487
rect 2558 471 2564 472
rect 2558 467 2559 471
rect 2563 467 2564 471
rect 2558 466 2564 467
rect 2636 464 2638 486
rect 2728 472 2730 493
rect 2726 471 2732 472
rect 2726 467 2727 471
rect 2731 467 2732 471
rect 2726 466 2732 467
rect 2804 464 2806 502
rect 2960 499 2962 524
rect 3036 512 3038 534
rect 3142 529 3148 530
rect 3142 525 3143 529
rect 3147 525 3148 529
rect 3142 524 3148 525
rect 3034 511 3040 512
rect 3034 507 3035 511
rect 3039 507 3040 511
rect 3034 506 3040 507
rect 3144 499 3146 524
rect 2895 498 2899 499
rect 2895 493 2899 494
rect 2959 498 2963 499
rect 2959 493 2963 494
rect 3063 498 3067 499
rect 3063 493 3067 494
rect 3143 498 3147 499
rect 3143 493 3147 494
rect 3223 498 3227 499
rect 3223 493 3227 494
rect 2896 472 2898 493
rect 2978 491 2984 492
rect 2978 487 2979 491
rect 2983 487 2984 491
rect 2978 486 2984 487
rect 2894 471 2900 472
rect 2894 467 2895 471
rect 2899 467 2900 471
rect 2894 466 2900 467
rect 2980 464 2982 486
rect 3064 472 3066 493
rect 3118 491 3124 492
rect 3118 487 3119 491
rect 3123 487 3124 491
rect 3118 486 3124 487
rect 3120 477 3122 486
rect 3119 476 3123 477
rect 3224 472 3226 493
rect 3232 492 3234 534
rect 3240 520 3242 534
rect 3318 529 3324 530
rect 3318 525 3319 529
rect 3323 525 3324 529
rect 3318 524 3324 525
rect 3494 529 3500 530
rect 3494 525 3495 529
rect 3499 525 3500 529
rect 3494 524 3500 525
rect 3238 519 3244 520
rect 3238 515 3239 519
rect 3243 515 3244 519
rect 3238 514 3244 515
rect 3320 499 3322 524
rect 3496 499 3498 524
rect 3612 512 3614 614
rect 3694 612 3700 613
rect 3694 608 3695 612
rect 3699 608 3700 612
rect 3694 607 3700 608
rect 3696 579 3698 607
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3695 578 3699 579
rect 3695 573 3699 574
rect 3680 549 3682 573
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3678 543 3684 544
rect 3678 529 3684 530
rect 3678 525 3679 529
rect 3683 525 3684 529
rect 3678 524 3684 525
rect 3610 511 3616 512
rect 3610 507 3611 511
rect 3615 507 3616 511
rect 3610 506 3616 507
rect 3680 499 3682 524
rect 3319 498 3323 499
rect 3319 493 3323 494
rect 3383 498 3387 499
rect 3383 493 3387 494
rect 3495 498 3499 499
rect 3495 493 3499 494
rect 3543 498 3547 499
rect 3543 493 3547 494
rect 3679 498 3683 499
rect 3679 493 3683 494
rect 3703 498 3707 499
rect 3703 493 3707 494
rect 3230 491 3236 492
rect 3230 487 3231 491
rect 3235 487 3236 491
rect 3230 486 3236 487
rect 3298 491 3304 492
rect 3298 487 3299 491
rect 3303 487 3304 491
rect 3298 486 3304 487
rect 3062 471 3068 472
rect 3119 471 3123 472
rect 3222 471 3228 472
rect 3062 467 3063 471
rect 3067 467 3068 471
rect 3062 466 3068 467
rect 3222 467 3223 471
rect 3227 467 3228 471
rect 3222 466 3228 467
rect 3300 464 3302 486
rect 3319 476 3323 477
rect 3384 472 3386 493
rect 3544 472 3546 493
rect 3618 491 3624 492
rect 3618 487 3619 491
rect 3623 487 3624 491
rect 3618 486 3624 487
rect 3319 471 3323 472
rect 3382 471 3388 472
rect 3320 464 3322 471
rect 3382 467 3383 471
rect 3387 467 3388 471
rect 3382 466 3388 467
rect 3542 471 3548 472
rect 3542 467 3543 471
rect 3547 467 3548 471
rect 3542 466 3548 467
rect 3620 464 3622 486
rect 3704 472 3706 493
rect 3702 471 3708 472
rect 3702 467 3703 471
rect 3707 467 3708 471
rect 3702 466 3708 467
rect 3780 464 3782 646
rect 3840 632 3842 653
rect 3908 652 3910 690
rect 3942 684 3948 685
rect 3942 680 3943 684
rect 3947 680 3948 684
rect 3942 679 3948 680
rect 3944 659 3946 679
rect 3943 658 3947 659
rect 3943 653 3947 654
rect 3906 651 3912 652
rect 3906 647 3907 651
rect 3911 647 3912 651
rect 3906 646 3912 647
rect 3944 633 3946 653
rect 3942 632 3948 633
rect 3838 631 3844 632
rect 3838 627 3839 631
rect 3843 627 3844 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3838 626 3844 627
rect 3914 619 3920 620
rect 3914 615 3915 619
rect 3919 615 3920 619
rect 3914 614 3920 615
rect 3942 615 3948 616
rect 3838 612 3844 613
rect 3838 608 3839 612
rect 3843 608 3844 612
rect 3838 607 3844 608
rect 3840 579 3842 607
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3840 549 3842 573
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3906 539 3912 540
rect 3906 535 3907 539
rect 3911 535 3912 539
rect 3906 534 3912 535
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3840 499 3842 524
rect 3839 498 3843 499
rect 3839 493 3843 494
rect 3798 483 3804 484
rect 3798 479 3799 483
rect 3803 479 3804 483
rect 3798 478 3804 479
rect 3800 464 3802 478
rect 3840 472 3842 493
rect 3908 492 3910 534
rect 3916 512 3918 614
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3944 579 3946 610
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 3944 546 3946 573
rect 3942 545 3948 546
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 3942 523 3948 524
rect 3914 511 3920 512
rect 3914 507 3915 511
rect 3919 507 3920 511
rect 3914 506 3920 507
rect 3944 499 3946 523
rect 3943 498 3947 499
rect 3943 493 3947 494
rect 3906 491 3912 492
rect 3906 487 3907 491
rect 3911 487 3912 491
rect 3906 486 3912 487
rect 3944 473 3946 493
rect 3942 472 3948 473
rect 3838 471 3844 472
rect 3838 467 3839 471
rect 3843 467 3844 471
rect 3942 468 3943 472
rect 3947 468 3948 472
rect 3942 467 3948 468
rect 3838 466 3844 467
rect 2298 463 2304 464
rect 2298 459 2299 463
rect 2303 459 2304 463
rect 2298 458 2304 459
rect 2466 463 2472 464
rect 2466 459 2467 463
rect 2471 459 2472 463
rect 2466 458 2472 459
rect 2634 463 2640 464
rect 2634 459 2635 463
rect 2639 459 2640 463
rect 2634 458 2640 459
rect 2802 463 2808 464
rect 2802 459 2803 463
rect 2807 459 2808 463
rect 2802 458 2808 459
rect 2886 463 2892 464
rect 2886 459 2887 463
rect 2891 459 2892 463
rect 2886 458 2892 459
rect 2978 463 2984 464
rect 2978 459 2979 463
rect 2983 459 2984 463
rect 2978 458 2984 459
rect 3298 463 3304 464
rect 3298 459 3299 463
rect 3303 459 3304 463
rect 3298 458 3304 459
rect 3318 463 3324 464
rect 3318 459 3319 463
rect 3323 459 3324 463
rect 3318 458 3324 459
rect 3618 463 3624 464
rect 3618 459 3619 463
rect 3623 459 3624 463
rect 3618 458 3624 459
rect 3778 463 3784 464
rect 3778 459 3779 463
rect 3783 459 3784 463
rect 3778 458 3784 459
rect 3798 463 3804 464
rect 3798 459 3799 463
rect 3803 459 3804 463
rect 3798 458 3804 459
rect 2390 452 2396 453
rect 2390 448 2391 452
rect 2395 448 2396 452
rect 2390 447 2396 448
rect 2558 452 2564 453
rect 2558 448 2559 452
rect 2563 448 2564 452
rect 2558 447 2564 448
rect 2726 452 2732 453
rect 2726 448 2727 452
rect 2731 448 2732 452
rect 2726 447 2732 448
rect 2392 423 2394 447
rect 2560 423 2562 447
rect 2728 423 2730 447
rect 2391 422 2395 423
rect 2391 417 2395 418
rect 2463 422 2467 423
rect 2463 417 2467 418
rect 2559 422 2563 423
rect 2559 417 2563 418
rect 2655 422 2659 423
rect 2655 417 2659 418
rect 2727 422 2731 423
rect 2727 417 2731 418
rect 2751 422 2755 423
rect 2751 417 2755 418
rect 2847 422 2851 423
rect 2847 417 2851 418
rect 2464 393 2466 417
rect 2560 393 2562 417
rect 2656 393 2658 417
rect 2752 393 2754 417
rect 2848 393 2850 417
rect 2462 392 2468 393
rect 2462 388 2463 392
rect 2467 388 2468 392
rect 2462 387 2468 388
rect 2558 392 2564 393
rect 2558 388 2559 392
rect 2563 388 2564 392
rect 2558 387 2564 388
rect 2654 392 2660 393
rect 2654 388 2655 392
rect 2659 388 2660 392
rect 2654 387 2660 388
rect 2750 392 2756 393
rect 2750 388 2751 392
rect 2755 388 2756 392
rect 2750 387 2756 388
rect 2846 392 2852 393
rect 2846 388 2847 392
rect 2851 388 2852 392
rect 2846 387 2852 388
rect 2262 383 2268 384
rect 2262 379 2263 383
rect 2267 379 2268 383
rect 2262 378 2268 379
rect 2550 383 2556 384
rect 2550 379 2551 383
rect 2555 379 2556 383
rect 2550 378 2556 379
rect 2646 383 2652 384
rect 2646 379 2647 383
rect 2651 379 2652 383
rect 2646 378 2652 379
rect 2742 383 2748 384
rect 2742 379 2743 383
rect 2747 379 2748 383
rect 2742 378 2748 379
rect 2462 373 2468 374
rect 2046 372 2052 373
rect 2046 368 2047 372
rect 2051 368 2052 372
rect 2462 369 2463 373
rect 2467 369 2468 373
rect 2462 368 2468 369
rect 2046 367 2052 368
rect 2034 359 2040 360
rect 2034 355 2035 359
rect 2039 355 2040 359
rect 2034 354 2040 355
rect 2048 347 2050 367
rect 2464 347 2466 368
rect 2552 356 2554 378
rect 2558 373 2564 374
rect 2558 369 2559 373
rect 2563 369 2564 373
rect 2558 368 2564 369
rect 2550 355 2556 356
rect 2550 351 2551 355
rect 2555 351 2556 355
rect 2550 350 2556 351
rect 2560 347 2562 368
rect 2648 356 2650 378
rect 2654 373 2660 374
rect 2654 369 2655 373
rect 2659 369 2660 373
rect 2654 368 2660 369
rect 2646 355 2652 356
rect 2646 351 2647 355
rect 2651 351 2652 355
rect 2646 350 2652 351
rect 2656 347 2658 368
rect 2744 356 2746 378
rect 2750 373 2756 374
rect 2750 369 2751 373
rect 2755 369 2756 373
rect 2750 368 2756 369
rect 2846 373 2852 374
rect 2846 369 2847 373
rect 2851 369 2852 373
rect 2846 368 2852 369
rect 2742 355 2748 356
rect 2742 351 2743 355
rect 2747 351 2748 355
rect 2742 350 2748 351
rect 2752 347 2754 368
rect 2848 347 2850 368
rect 2888 356 2890 458
rect 3942 455 3948 456
rect 2894 452 2900 453
rect 2894 448 2895 452
rect 2899 448 2900 452
rect 2894 447 2900 448
rect 3062 452 3068 453
rect 3062 448 3063 452
rect 3067 448 3068 452
rect 3062 447 3068 448
rect 3222 452 3228 453
rect 3222 448 3223 452
rect 3227 448 3228 452
rect 3222 447 3228 448
rect 3382 452 3388 453
rect 3382 448 3383 452
rect 3387 448 3388 452
rect 3382 447 3388 448
rect 3542 452 3548 453
rect 3542 448 3543 452
rect 3547 448 3548 452
rect 3542 447 3548 448
rect 3702 452 3708 453
rect 3702 448 3703 452
rect 3707 448 3708 452
rect 3702 447 3708 448
rect 3838 452 3844 453
rect 3838 448 3839 452
rect 3843 448 3844 452
rect 3942 451 3943 455
rect 3947 451 3948 455
rect 3942 450 3948 451
rect 3838 447 3844 448
rect 2896 423 2898 447
rect 3064 423 3066 447
rect 3224 423 3226 447
rect 3384 423 3386 447
rect 3544 423 3546 447
rect 3704 423 3706 447
rect 3840 423 3842 447
rect 3944 423 3946 450
rect 2895 422 2899 423
rect 2895 417 2899 418
rect 2943 422 2947 423
rect 2943 417 2947 418
rect 3039 422 3043 423
rect 3039 417 3043 418
rect 3063 422 3067 423
rect 3063 417 3067 418
rect 3135 422 3139 423
rect 3135 417 3139 418
rect 3223 422 3227 423
rect 3223 417 3227 418
rect 3231 422 3235 423
rect 3231 417 3235 418
rect 3383 422 3387 423
rect 3383 417 3387 418
rect 3543 422 3547 423
rect 3543 417 3547 418
rect 3703 422 3707 423
rect 3703 417 3707 418
rect 3839 422 3843 423
rect 3839 417 3843 418
rect 3943 422 3947 423
rect 3943 417 3947 418
rect 2944 393 2946 417
rect 3040 393 3042 417
rect 3136 393 3138 417
rect 3232 393 3234 417
rect 2942 392 2948 393
rect 2942 388 2943 392
rect 2947 388 2948 392
rect 2942 387 2948 388
rect 3038 392 3044 393
rect 3038 388 3039 392
rect 3043 388 3044 392
rect 3038 387 3044 388
rect 3134 392 3140 393
rect 3134 388 3135 392
rect 3139 388 3140 392
rect 3134 387 3140 388
rect 3230 392 3236 393
rect 3230 388 3231 392
rect 3235 388 3236 392
rect 3944 390 3946 417
rect 3230 387 3236 388
rect 3942 389 3948 390
rect 3942 385 3943 389
rect 3947 385 3948 389
rect 3942 384 3948 385
rect 2922 383 2928 384
rect 2922 379 2923 383
rect 2927 379 2928 383
rect 2922 378 2928 379
rect 3018 383 3024 384
rect 3018 379 3019 383
rect 3023 379 3024 383
rect 3018 378 3024 379
rect 3114 383 3120 384
rect 3114 379 3115 383
rect 3119 379 3120 383
rect 3114 378 3120 379
rect 3210 383 3216 384
rect 3210 379 3211 383
rect 3215 379 3216 383
rect 3210 378 3216 379
rect 3298 383 3304 384
rect 3298 379 3299 383
rect 3303 379 3304 383
rect 3298 378 3304 379
rect 2924 356 2926 378
rect 2942 373 2948 374
rect 2942 369 2943 373
rect 2947 369 2948 373
rect 2942 368 2948 369
rect 2886 355 2892 356
rect 2858 351 2864 352
rect 2858 347 2859 351
rect 2863 347 2864 351
rect 2886 351 2887 355
rect 2891 351 2892 355
rect 2886 350 2892 351
rect 2922 355 2928 356
rect 2922 351 2923 355
rect 2927 351 2928 355
rect 2922 350 2928 351
rect 2944 347 2946 368
rect 3020 356 3022 378
rect 3038 373 3044 374
rect 3038 369 3039 373
rect 3043 369 3044 373
rect 3038 368 3044 369
rect 3018 355 3024 356
rect 3018 351 3019 355
rect 3023 351 3024 355
rect 3018 350 3024 351
rect 3040 347 3042 368
rect 3116 356 3118 378
rect 3134 373 3140 374
rect 3134 369 3135 373
rect 3139 369 3140 373
rect 3134 368 3140 369
rect 3114 355 3120 356
rect 3114 351 3115 355
rect 3119 351 3120 355
rect 3114 350 3120 351
rect 3136 347 3138 368
rect 3212 356 3214 378
rect 3230 373 3236 374
rect 3230 369 3231 373
rect 3235 369 3236 373
rect 3230 368 3236 369
rect 3210 355 3216 356
rect 3210 351 3211 355
rect 3215 351 3216 355
rect 3210 350 3216 351
rect 3232 347 3234 368
rect 2007 346 2011 347
rect 2007 341 2011 342
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2399 346 2403 347
rect 2399 341 2403 342
rect 2463 346 2467 347
rect 2463 341 2467 342
rect 2503 346 2507 347
rect 2503 341 2507 342
rect 2559 346 2563 347
rect 2559 341 2563 342
rect 2623 346 2627 347
rect 2623 341 2627 342
rect 2655 346 2659 347
rect 2655 341 2659 342
rect 2751 346 2755 347
rect 2751 341 2755 342
rect 2759 346 2763 347
rect 2759 341 2763 342
rect 2847 346 2851 347
rect 2858 346 2864 347
rect 2911 346 2915 347
rect 2847 341 2851 342
rect 1970 339 1976 340
rect 1970 335 1971 339
rect 1975 335 1976 339
rect 1970 334 1976 335
rect 2008 321 2010 341
rect 2048 321 2050 341
rect 2006 320 2012 321
rect 1894 319 1900 320
rect 1894 315 1895 319
rect 1899 315 1900 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 2400 320 2402 341
rect 2438 339 2444 340
rect 2438 335 2439 339
rect 2443 335 2444 339
rect 2438 334 2444 335
rect 2474 339 2480 340
rect 2474 335 2475 339
rect 2479 335 2480 339
rect 2474 334 2480 335
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2398 319 2404 320
rect 2398 315 2399 319
rect 2403 315 2404 319
rect 1894 314 1900 315
rect 2398 314 2404 315
rect 242 311 248 312
rect 242 307 243 311
rect 247 307 248 311
rect 242 306 248 307
rect 626 311 632 312
rect 626 307 627 311
rect 631 307 632 311
rect 626 306 632 307
rect 834 311 840 312
rect 834 307 835 311
rect 839 307 840 311
rect 834 306 840 307
rect 902 311 908 312
rect 902 307 903 311
rect 907 307 908 311
rect 902 306 908 307
rect 1234 311 1240 312
rect 1234 307 1235 311
rect 1239 307 1240 311
rect 1234 306 1240 307
rect 1418 311 1424 312
rect 1418 307 1419 311
rect 1423 307 1424 311
rect 1418 306 1424 307
rect 1602 311 1608 312
rect 1602 307 1603 311
rect 1607 307 1608 311
rect 1818 311 1824 312
rect 1602 306 1608 307
rect 1786 307 1792 308
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 110 298 116 299
rect 158 300 164 301
rect 112 263 114 298
rect 158 296 159 300
rect 163 296 164 300
rect 158 295 164 296
rect 350 300 356 301
rect 350 296 351 300
rect 355 296 356 300
rect 350 295 356 296
rect 550 300 556 301
rect 550 296 551 300
rect 555 296 556 300
rect 550 295 556 296
rect 758 300 764 301
rect 758 296 759 300
rect 763 296 764 300
rect 758 295 764 296
rect 160 263 162 295
rect 352 263 354 295
rect 552 263 554 295
rect 760 263 762 295
rect 111 262 115 263
rect 111 257 115 258
rect 159 262 163 263
rect 159 257 163 258
rect 223 262 227 263
rect 223 257 227 258
rect 351 262 355 263
rect 351 257 355 258
rect 383 262 387 263
rect 383 257 387 258
rect 543 262 547 263
rect 543 257 547 258
rect 551 262 555 263
rect 551 257 555 258
rect 703 262 707 263
rect 703 257 707 258
rect 759 262 763 263
rect 759 257 763 258
rect 863 262 867 263
rect 863 257 867 258
rect 112 230 114 257
rect 224 233 226 257
rect 384 233 386 257
rect 544 233 546 257
rect 704 233 706 257
rect 864 233 866 257
rect 222 232 228 233
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 222 228 223 232
rect 227 228 228 232
rect 222 227 228 228
rect 382 232 388 233
rect 382 228 383 232
rect 387 228 388 232
rect 382 227 388 228
rect 542 232 548 233
rect 542 228 543 232
rect 547 228 548 232
rect 542 227 548 228
rect 702 232 708 233
rect 702 228 703 232
rect 707 228 708 232
rect 702 227 708 228
rect 862 232 868 233
rect 862 228 863 232
rect 867 228 868 232
rect 862 227 868 228
rect 110 224 116 225
rect 298 223 304 224
rect 298 219 299 223
rect 303 219 304 223
rect 298 218 304 219
rect 618 223 624 224
rect 618 219 619 223
rect 623 219 624 223
rect 618 218 624 219
rect 798 223 804 224
rect 798 219 799 223
rect 803 219 804 223
rect 798 218 804 219
rect 222 213 228 214
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 222 209 223 213
rect 227 209 228 213
rect 222 208 228 209
rect 110 207 116 208
rect 112 167 114 207
rect 224 167 226 208
rect 300 196 302 218
rect 382 213 388 214
rect 382 209 383 213
rect 387 209 388 213
rect 382 208 388 209
rect 542 213 548 214
rect 542 209 543 213
rect 547 209 548 213
rect 542 208 548 209
rect 298 195 304 196
rect 298 191 299 195
rect 303 191 304 195
rect 298 190 304 191
rect 306 187 312 188
rect 306 183 307 187
rect 311 183 312 187
rect 306 182 312 183
rect 111 166 115 167
rect 111 161 115 162
rect 135 166 139 167
rect 135 161 139 162
rect 223 166 227 167
rect 223 161 227 162
rect 231 166 235 167
rect 231 161 235 162
rect 112 141 114 161
rect 110 140 116 141
rect 136 140 138 161
rect 210 159 216 160
rect 210 155 211 159
rect 215 155 216 159
rect 210 154 216 155
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 212 132 214 154
rect 232 140 234 161
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 308 132 310 182
rect 384 167 386 208
rect 544 167 546 208
rect 327 166 331 167
rect 327 161 331 162
rect 383 166 387 167
rect 383 161 387 162
rect 423 166 427 167
rect 423 161 427 162
rect 527 166 531 167
rect 527 161 531 162
rect 543 166 547 167
rect 543 161 547 162
rect 314 151 320 152
rect 314 147 315 151
rect 319 147 320 151
rect 314 146 320 147
rect 316 132 318 146
rect 328 140 330 161
rect 410 159 416 160
rect 410 155 411 159
rect 415 155 416 159
rect 410 154 416 155
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 412 132 414 154
rect 424 140 426 161
rect 506 159 512 160
rect 506 155 507 159
rect 511 155 512 159
rect 506 154 512 155
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 508 132 510 154
rect 528 140 530 161
rect 620 160 622 218
rect 702 213 708 214
rect 702 209 703 213
rect 707 209 708 213
rect 702 208 708 209
rect 704 167 706 208
rect 800 196 802 218
rect 862 213 868 214
rect 862 209 863 213
rect 867 209 868 213
rect 862 208 868 209
rect 798 195 804 196
rect 798 191 799 195
rect 803 191 804 195
rect 798 190 804 191
rect 864 167 866 208
rect 904 196 906 306
rect 1786 303 1787 307
rect 1791 303 1792 307
rect 1818 307 1819 311
rect 1823 307 1824 311
rect 1818 306 1824 307
rect 1786 302 1792 303
rect 2006 303 2012 304
rect 958 300 964 301
rect 958 296 959 300
rect 963 296 964 300
rect 958 295 964 296
rect 1158 300 1164 301
rect 1158 296 1159 300
rect 1163 296 1164 300
rect 1158 295 1164 296
rect 1342 300 1348 301
rect 1342 296 1343 300
rect 1347 296 1348 300
rect 1342 295 1348 296
rect 1526 300 1532 301
rect 1526 296 1527 300
rect 1531 296 1532 300
rect 1526 295 1532 296
rect 1710 300 1716 301
rect 1710 296 1711 300
rect 1715 296 1716 300
rect 1710 295 1716 296
rect 960 263 962 295
rect 1160 263 1162 295
rect 1344 263 1346 295
rect 1528 263 1530 295
rect 1712 263 1714 295
rect 959 262 963 263
rect 959 257 963 258
rect 1031 262 1035 263
rect 1031 257 1035 258
rect 1159 262 1163 263
rect 1159 257 1163 258
rect 1199 262 1203 263
rect 1199 257 1203 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1367 262 1371 263
rect 1367 257 1371 258
rect 1527 262 1531 263
rect 1527 257 1531 258
rect 1543 262 1547 263
rect 1543 257 1547 258
rect 1711 262 1715 263
rect 1711 257 1715 258
rect 1727 262 1731 263
rect 1727 257 1731 258
rect 1032 233 1034 257
rect 1200 233 1202 257
rect 1368 233 1370 257
rect 1544 233 1546 257
rect 1728 233 1730 257
rect 1030 232 1036 233
rect 1030 228 1031 232
rect 1035 228 1036 232
rect 1030 227 1036 228
rect 1198 232 1204 233
rect 1198 228 1199 232
rect 1203 228 1204 232
rect 1198 227 1204 228
rect 1366 232 1372 233
rect 1366 228 1367 232
rect 1371 228 1372 232
rect 1366 227 1372 228
rect 1542 232 1548 233
rect 1542 228 1543 232
rect 1547 228 1548 232
rect 1542 227 1548 228
rect 1726 232 1732 233
rect 1726 228 1727 232
rect 1731 228 1732 232
rect 1726 227 1732 228
rect 1098 223 1104 224
rect 1098 219 1099 223
rect 1103 219 1104 223
rect 1098 218 1104 219
rect 1114 223 1120 224
rect 1114 219 1115 223
rect 1119 219 1120 223
rect 1114 218 1120 219
rect 1626 223 1632 224
rect 1626 219 1627 223
rect 1631 219 1632 223
rect 1626 218 1632 219
rect 1030 213 1036 214
rect 1030 209 1031 213
rect 1035 209 1036 213
rect 1030 208 1036 209
rect 902 195 908 196
rect 902 191 903 195
rect 907 191 908 195
rect 902 190 908 191
rect 1032 167 1034 208
rect 647 166 651 167
rect 647 161 651 162
rect 703 166 707 167
rect 703 161 707 162
rect 775 166 779 167
rect 775 161 779 162
rect 863 166 867 167
rect 863 161 867 162
rect 903 166 907 167
rect 903 161 907 162
rect 1031 166 1035 167
rect 1031 161 1035 162
rect 618 159 624 160
rect 618 155 619 159
rect 623 155 624 159
rect 618 154 624 155
rect 648 140 650 161
rect 722 159 728 160
rect 722 155 723 159
rect 727 155 728 159
rect 722 154 728 155
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 724 132 726 154
rect 776 140 778 161
rect 850 159 856 160
rect 850 155 851 159
rect 855 155 856 159
rect 850 154 856 155
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 852 132 854 154
rect 858 151 864 152
rect 858 147 859 151
rect 863 147 864 151
rect 858 146 864 147
rect 860 132 862 146
rect 904 140 906 161
rect 1032 140 1034 161
rect 1100 160 1102 218
rect 1116 196 1118 218
rect 1198 213 1204 214
rect 1198 209 1199 213
rect 1203 209 1204 213
rect 1198 208 1204 209
rect 1366 213 1372 214
rect 1366 209 1367 213
rect 1371 209 1372 213
rect 1366 208 1372 209
rect 1542 213 1548 214
rect 1542 209 1543 213
rect 1547 209 1548 213
rect 1542 208 1548 209
rect 1114 195 1120 196
rect 1114 191 1115 195
rect 1119 191 1120 195
rect 1114 190 1120 191
rect 1200 167 1202 208
rect 1368 167 1370 208
rect 1544 167 1546 208
rect 1628 196 1630 218
rect 1726 213 1732 214
rect 1726 209 1727 213
rect 1731 209 1732 213
rect 1726 208 1732 209
rect 1626 195 1632 196
rect 1626 191 1627 195
rect 1631 191 1632 195
rect 1626 190 1632 191
rect 1728 167 1730 208
rect 1788 196 1790 302
rect 1894 300 1900 301
rect 1894 296 1895 300
rect 1899 296 1900 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 2046 298 2052 299
rect 2398 300 2404 301
rect 1894 295 1900 296
rect 1896 263 1898 295
rect 2008 263 2010 298
rect 2048 271 2050 298
rect 2398 296 2399 300
rect 2403 296 2404 300
rect 2398 295 2404 296
rect 2400 271 2402 295
rect 2047 270 2051 271
rect 2047 265 2051 266
rect 2191 270 2195 271
rect 2191 265 2195 266
rect 2351 270 2355 271
rect 2351 265 2355 266
rect 2399 270 2403 271
rect 2399 265 2403 266
rect 1895 262 1899 263
rect 1895 257 1899 258
rect 1903 262 1907 263
rect 1903 257 1907 258
rect 2007 262 2011 263
rect 2007 257 2011 258
rect 1904 233 1906 257
rect 1902 232 1908 233
rect 1902 228 1903 232
rect 1907 228 1908 232
rect 2008 230 2010 257
rect 2048 238 2050 265
rect 2192 241 2194 265
rect 2352 241 2354 265
rect 2440 248 2442 334
rect 2476 312 2478 334
rect 2504 320 2506 341
rect 2578 339 2584 340
rect 2578 335 2579 339
rect 2583 335 2584 339
rect 2578 334 2584 335
rect 2502 319 2508 320
rect 2502 315 2503 319
rect 2507 315 2508 319
rect 2502 314 2508 315
rect 2580 312 2582 334
rect 2624 320 2626 341
rect 2698 339 2704 340
rect 2698 335 2699 339
rect 2703 335 2704 339
rect 2698 334 2704 335
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2700 312 2702 334
rect 2760 320 2762 341
rect 2834 339 2840 340
rect 2834 335 2835 339
rect 2839 335 2840 339
rect 2834 334 2840 335
rect 2758 319 2764 320
rect 2758 315 2759 319
rect 2763 315 2764 319
rect 2758 314 2764 315
rect 2836 312 2838 334
rect 2860 312 2862 346
rect 2911 341 2915 342
rect 2943 346 2947 347
rect 2943 341 2947 342
rect 3039 346 3043 347
rect 3039 341 3043 342
rect 3071 346 3075 347
rect 3071 341 3075 342
rect 3135 346 3139 347
rect 3135 341 3139 342
rect 3231 346 3235 347
rect 3231 341 3235 342
rect 3247 346 3251 347
rect 3247 341 3251 342
rect 2912 320 2914 341
rect 3072 320 3074 341
rect 3154 339 3160 340
rect 3154 335 3155 339
rect 3159 335 3160 339
rect 3154 334 3160 335
rect 2910 319 2916 320
rect 2910 315 2911 319
rect 2915 315 2916 319
rect 2910 314 2916 315
rect 3070 319 3076 320
rect 3070 315 3071 319
rect 3075 315 3076 319
rect 3070 314 3076 315
rect 3156 312 3158 334
rect 3248 320 3250 341
rect 3300 340 3302 378
rect 3942 372 3948 373
rect 3942 368 3943 372
rect 3947 368 3948 372
rect 3942 367 3948 368
rect 3944 347 3946 367
rect 3423 346 3427 347
rect 3423 341 3427 342
rect 3607 346 3611 347
rect 3607 341 3611 342
rect 3791 346 3795 347
rect 3791 341 3795 342
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 3298 339 3304 340
rect 3298 335 3299 339
rect 3303 335 3304 339
rect 3298 334 3304 335
rect 3424 320 3426 341
rect 3558 339 3564 340
rect 3558 335 3559 339
rect 3563 335 3564 339
rect 3558 334 3564 335
rect 3498 331 3504 332
rect 3498 327 3499 331
rect 3503 327 3504 331
rect 3498 326 3504 327
rect 3246 319 3252 320
rect 3246 315 3247 319
rect 3251 315 3252 319
rect 3246 314 3252 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3500 312 3502 326
rect 2474 311 2480 312
rect 2474 307 2475 311
rect 2479 307 2480 311
rect 2474 306 2480 307
rect 2578 311 2584 312
rect 2578 307 2579 311
rect 2583 307 2584 311
rect 2578 306 2584 307
rect 2698 311 2704 312
rect 2698 307 2699 311
rect 2703 307 2704 311
rect 2698 306 2704 307
rect 2834 311 2840 312
rect 2834 307 2835 311
rect 2839 307 2840 311
rect 2834 306 2840 307
rect 2858 311 2864 312
rect 2858 307 2859 311
rect 2863 307 2864 311
rect 2858 306 2864 307
rect 3002 311 3008 312
rect 3002 307 3003 311
rect 3007 307 3008 311
rect 3002 306 3008 307
rect 3154 311 3160 312
rect 3154 307 3155 311
rect 3159 307 3160 311
rect 3154 306 3160 307
rect 3498 311 3504 312
rect 3498 307 3499 311
rect 3503 307 3504 311
rect 3498 306 3504 307
rect 2502 300 2508 301
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2758 300 2764 301
rect 2758 296 2759 300
rect 2763 296 2764 300
rect 2758 295 2764 296
rect 2910 300 2916 301
rect 2910 296 2911 300
rect 2915 296 2916 300
rect 2910 295 2916 296
rect 2504 271 2506 295
rect 2624 271 2626 295
rect 2760 271 2762 295
rect 2912 271 2914 295
rect 2503 270 2507 271
rect 2503 265 2507 266
rect 2519 270 2523 271
rect 2519 265 2523 266
rect 2623 270 2627 271
rect 2623 265 2627 266
rect 2687 270 2691 271
rect 2687 265 2691 266
rect 2759 270 2763 271
rect 2759 265 2763 266
rect 2855 270 2859 271
rect 2855 265 2859 266
rect 2911 270 2915 271
rect 2911 265 2915 266
rect 2438 247 2444 248
rect 2438 243 2439 247
rect 2443 243 2444 247
rect 2438 242 2444 243
rect 2520 241 2522 265
rect 2688 241 2690 265
rect 2856 241 2858 265
rect 2190 240 2196 241
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2190 236 2191 240
rect 2195 236 2196 240
rect 2190 235 2196 236
rect 2350 240 2356 241
rect 2350 236 2351 240
rect 2355 236 2356 240
rect 2350 235 2356 236
rect 2518 240 2524 241
rect 2518 236 2519 240
rect 2523 236 2524 240
rect 2518 235 2524 236
rect 2686 240 2692 241
rect 2686 236 2687 240
rect 2691 236 2692 240
rect 2686 235 2692 236
rect 2854 240 2860 241
rect 2854 236 2855 240
rect 2859 236 2860 240
rect 2854 235 2860 236
rect 2046 232 2052 233
rect 2266 231 2272 232
rect 1902 227 1908 228
rect 2006 229 2012 230
rect 2006 225 2007 229
rect 2011 225 2012 229
rect 2266 227 2267 231
rect 2271 227 2272 231
rect 2266 226 2272 227
rect 2426 231 2432 232
rect 2426 227 2427 231
rect 2431 227 2432 231
rect 2426 226 2432 227
rect 2594 231 2600 232
rect 2594 227 2595 231
rect 2599 227 2600 231
rect 2594 226 2600 227
rect 2930 231 2936 232
rect 2930 227 2931 231
rect 2935 227 2936 231
rect 2930 226 2936 227
rect 2006 224 2012 225
rect 1970 223 1976 224
rect 1970 219 1971 223
rect 1975 219 1976 223
rect 2190 221 2196 222
rect 1970 218 1976 219
rect 2046 220 2052 221
rect 1902 213 1908 214
rect 1902 209 1903 213
rect 1907 209 1908 213
rect 1902 208 1908 209
rect 1786 195 1792 196
rect 1786 191 1787 195
rect 1791 191 1792 195
rect 1786 190 1792 191
rect 1882 191 1888 192
rect 1882 187 1883 191
rect 1887 187 1888 191
rect 1882 186 1888 187
rect 1151 166 1155 167
rect 1151 161 1155 162
rect 1199 166 1203 167
rect 1199 161 1203 162
rect 1271 166 1275 167
rect 1271 161 1275 162
rect 1367 166 1371 167
rect 1367 161 1371 162
rect 1383 166 1387 167
rect 1383 161 1387 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1543 166 1547 167
rect 1543 161 1547 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1703 166 1707 167
rect 1703 161 1707 162
rect 1727 166 1731 167
rect 1727 161 1731 162
rect 1807 166 1811 167
rect 1807 161 1811 162
rect 1098 159 1104 160
rect 1098 155 1099 159
rect 1103 155 1104 159
rect 1098 154 1104 155
rect 1106 159 1112 160
rect 1106 155 1107 159
rect 1111 155 1112 159
rect 1106 154 1112 155
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1108 132 1110 154
rect 1152 140 1154 161
rect 1226 159 1232 160
rect 1226 155 1227 159
rect 1231 155 1232 159
rect 1226 154 1232 155
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1228 132 1230 154
rect 1272 140 1274 161
rect 1346 159 1352 160
rect 1346 155 1347 159
rect 1351 155 1352 159
rect 1346 154 1352 155
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1348 132 1350 154
rect 1384 140 1386 161
rect 1458 159 1464 160
rect 1458 155 1459 159
rect 1463 155 1464 159
rect 1458 154 1464 155
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1460 132 1462 154
rect 1488 140 1490 161
rect 1562 159 1568 160
rect 1562 155 1563 159
rect 1567 155 1568 159
rect 1562 154 1568 155
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1564 132 1566 154
rect 1592 140 1594 161
rect 1666 159 1672 160
rect 1666 155 1667 159
rect 1671 155 1672 159
rect 1666 154 1672 155
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1668 132 1670 154
rect 1704 140 1706 161
rect 1778 159 1784 160
rect 1778 155 1779 159
rect 1783 155 1784 159
rect 1778 154 1784 155
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1780 132 1782 154
rect 1808 140 1810 161
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1884 132 1886 186
rect 1904 167 1906 208
rect 1903 166 1907 167
rect 1903 161 1907 162
rect 1904 140 1906 161
rect 1972 160 1974 218
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2190 217 2191 221
rect 2195 217 2196 221
rect 2190 216 2196 217
rect 2046 215 2052 216
rect 2006 212 2012 213
rect 2006 208 2007 212
rect 2011 208 2012 212
rect 2006 207 2012 208
rect 2008 167 2010 207
rect 2007 166 2011 167
rect 2048 163 2050 215
rect 2192 163 2194 216
rect 2268 204 2270 226
rect 2350 221 2356 222
rect 2350 217 2351 221
rect 2355 217 2356 221
rect 2350 216 2356 217
rect 2266 203 2272 204
rect 2266 199 2267 203
rect 2271 199 2272 203
rect 2266 198 2272 199
rect 2352 163 2354 216
rect 2428 204 2430 226
rect 2518 221 2524 222
rect 2518 217 2519 221
rect 2523 217 2524 221
rect 2518 216 2524 217
rect 2426 203 2432 204
rect 2426 199 2427 203
rect 2431 199 2432 203
rect 2426 198 2432 199
rect 2520 163 2522 216
rect 2596 204 2598 226
rect 2686 221 2692 222
rect 2686 217 2687 221
rect 2691 217 2692 221
rect 2686 216 2692 217
rect 2854 221 2860 222
rect 2854 217 2855 221
rect 2859 217 2860 221
rect 2854 216 2860 217
rect 2594 203 2600 204
rect 2594 199 2595 203
rect 2599 199 2600 203
rect 2594 198 2600 199
rect 2688 163 2690 216
rect 2726 191 2732 192
rect 2726 187 2727 191
rect 2731 187 2732 191
rect 2726 186 2732 187
rect 2007 161 2011 162
rect 2047 162 2051 163
rect 1970 159 1976 160
rect 1970 155 1971 159
rect 1975 155 1976 159
rect 1970 154 1976 155
rect 1978 155 1984 156
rect 1978 151 1979 155
rect 1983 151 1984 155
rect 1978 150 1984 151
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 1902 134 1908 135
rect 1980 132 1982 150
rect 2008 141 2010 161
rect 2047 157 2051 158
rect 2071 162 2075 163
rect 2071 157 2075 158
rect 2167 162 2171 163
rect 2167 157 2171 158
rect 2191 162 2195 163
rect 2191 157 2195 158
rect 2263 162 2267 163
rect 2263 157 2267 158
rect 2351 162 2355 163
rect 2351 157 2355 158
rect 2367 162 2371 163
rect 2367 157 2371 158
rect 2487 162 2491 163
rect 2487 157 2491 158
rect 2519 162 2523 163
rect 2519 157 2523 158
rect 2615 162 2619 163
rect 2615 157 2619 158
rect 2687 162 2691 163
rect 2687 157 2691 158
rect 2006 140 2012 141
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2048 137 2050 157
rect 2006 135 2012 136
rect 2046 136 2052 137
rect 2072 136 2074 157
rect 2146 155 2152 156
rect 2146 151 2147 155
rect 2151 151 2152 155
rect 2146 150 2152 151
rect 2046 132 2047 136
rect 2051 132 2052 136
rect 210 131 216 132
rect 210 127 211 131
rect 215 127 216 131
rect 210 126 216 127
rect 306 131 312 132
rect 306 127 307 131
rect 311 127 312 131
rect 306 126 312 127
rect 314 131 320 132
rect 314 127 315 131
rect 319 127 320 131
rect 314 126 320 127
rect 410 131 416 132
rect 410 127 411 131
rect 415 127 416 131
rect 410 126 416 127
rect 506 131 512 132
rect 506 127 507 131
rect 511 127 512 131
rect 506 126 512 127
rect 722 131 728 132
rect 722 127 723 131
rect 727 127 728 131
rect 722 126 728 127
rect 850 131 856 132
rect 850 127 851 131
rect 855 127 856 131
rect 850 126 856 127
rect 858 131 864 132
rect 858 127 859 131
rect 863 127 864 131
rect 858 126 864 127
rect 1106 131 1112 132
rect 1106 127 1107 131
rect 1111 127 1112 131
rect 1106 126 1112 127
rect 1226 131 1232 132
rect 1226 127 1227 131
rect 1231 127 1232 131
rect 1226 126 1232 127
rect 1346 131 1352 132
rect 1346 127 1347 131
rect 1351 127 1352 131
rect 1346 126 1352 127
rect 1458 131 1464 132
rect 1458 127 1459 131
rect 1463 127 1464 131
rect 1458 126 1464 127
rect 1562 131 1568 132
rect 1562 127 1563 131
rect 1567 127 1568 131
rect 1562 126 1568 127
rect 1666 131 1672 132
rect 1666 127 1667 131
rect 1671 127 1672 131
rect 1666 126 1672 127
rect 1778 131 1784 132
rect 1778 127 1779 131
rect 1783 127 1784 131
rect 1778 126 1784 127
rect 1882 131 1888 132
rect 1882 127 1883 131
rect 1887 127 1888 131
rect 1882 126 1888 127
rect 1978 131 1984 132
rect 2046 131 2052 132
rect 2070 135 2076 136
rect 2070 131 2071 135
rect 2075 131 2076 135
rect 1978 127 1979 131
rect 1983 127 1984 131
rect 2070 130 2076 131
rect 2148 128 2150 150
rect 2168 136 2170 157
rect 2242 155 2248 156
rect 2242 151 2243 155
rect 2247 151 2248 155
rect 2242 150 2248 151
rect 2166 135 2172 136
rect 2166 131 2167 135
rect 2171 131 2172 135
rect 2166 130 2172 131
rect 2244 128 2246 150
rect 2264 136 2266 157
rect 2338 155 2344 156
rect 2338 151 2339 155
rect 2343 151 2344 155
rect 2338 150 2344 151
rect 2262 135 2268 136
rect 2262 131 2263 135
rect 2267 131 2268 135
rect 2262 130 2268 131
rect 2340 128 2342 150
rect 2368 136 2370 157
rect 2442 155 2448 156
rect 2442 151 2443 155
rect 2447 151 2448 155
rect 2442 150 2448 151
rect 2366 135 2372 136
rect 2366 131 2367 135
rect 2371 131 2372 135
rect 2366 130 2372 131
rect 2444 128 2446 150
rect 2488 136 2490 157
rect 2562 155 2568 156
rect 2562 151 2563 155
rect 2567 151 2568 155
rect 2562 150 2568 151
rect 2486 135 2492 136
rect 2486 131 2487 135
rect 2491 131 2492 135
rect 2486 130 2492 131
rect 2564 128 2566 150
rect 2616 136 2618 157
rect 2718 155 2724 156
rect 2718 151 2719 155
rect 2723 151 2724 155
rect 2718 150 2724 151
rect 2614 135 2620 136
rect 2614 131 2615 135
rect 2619 131 2620 135
rect 2614 130 2620 131
rect 2720 128 2722 150
rect 2728 128 2730 186
rect 2856 163 2858 216
rect 2932 204 2934 226
rect 3004 212 3006 306
rect 3070 300 3076 301
rect 3070 296 3071 300
rect 3075 296 3076 300
rect 3070 295 3076 296
rect 3246 300 3252 301
rect 3246 296 3247 300
rect 3251 296 3252 300
rect 3246 295 3252 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3072 271 3074 295
rect 3248 271 3250 295
rect 3424 271 3426 295
rect 3031 270 3035 271
rect 3031 265 3035 266
rect 3071 270 3075 271
rect 3071 265 3075 266
rect 3215 270 3219 271
rect 3215 265 3219 266
rect 3247 270 3251 271
rect 3247 265 3251 266
rect 3407 270 3411 271
rect 3407 265 3411 266
rect 3423 270 3427 271
rect 3423 265 3427 266
rect 3032 241 3034 265
rect 3216 241 3218 265
rect 3408 241 3410 265
rect 3030 240 3036 241
rect 3030 236 3031 240
rect 3035 236 3036 240
rect 3030 235 3036 236
rect 3214 240 3220 241
rect 3214 236 3215 240
rect 3219 236 3220 240
rect 3214 235 3220 236
rect 3406 240 3412 241
rect 3406 236 3407 240
rect 3411 236 3412 240
rect 3406 235 3412 236
rect 3560 232 3562 334
rect 3608 320 3610 341
rect 3682 339 3688 340
rect 3682 335 3683 339
rect 3687 335 3688 339
rect 3682 334 3688 335
rect 3606 319 3612 320
rect 3606 315 3607 319
rect 3611 315 3612 319
rect 3606 314 3612 315
rect 3684 312 3686 334
rect 3792 320 3794 341
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 3790 319 3796 320
rect 3790 315 3791 319
rect 3795 315 3796 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3790 314 3796 315
rect 3682 311 3688 312
rect 3682 307 3683 311
rect 3687 307 3688 311
rect 3682 306 3688 307
rect 3866 307 3872 308
rect 3866 303 3867 307
rect 3871 303 3872 307
rect 3866 302 3872 303
rect 3942 303 3948 304
rect 3606 300 3612 301
rect 3606 296 3607 300
rect 3611 296 3612 300
rect 3606 295 3612 296
rect 3790 300 3796 301
rect 3790 296 3791 300
rect 3795 296 3796 300
rect 3790 295 3796 296
rect 3608 271 3610 295
rect 3792 271 3794 295
rect 3607 270 3611 271
rect 3607 265 3611 266
rect 3791 270 3795 271
rect 3791 265 3795 266
rect 3807 270 3811 271
rect 3807 265 3811 266
rect 3608 241 3610 265
rect 3808 241 3810 265
rect 3606 240 3612 241
rect 3606 236 3607 240
rect 3611 236 3612 240
rect 3606 235 3612 236
rect 3806 240 3812 241
rect 3806 236 3807 240
rect 3811 236 3812 240
rect 3806 235 3812 236
rect 3106 231 3112 232
rect 3106 227 3107 231
rect 3111 227 3112 231
rect 3106 226 3112 227
rect 3290 231 3296 232
rect 3290 227 3291 231
rect 3295 227 3296 231
rect 3290 226 3296 227
rect 3378 231 3384 232
rect 3378 227 3379 231
rect 3383 227 3384 231
rect 3378 226 3384 227
rect 3558 231 3564 232
rect 3558 227 3559 231
rect 3563 227 3564 231
rect 3558 226 3564 227
rect 3782 231 3788 232
rect 3782 227 3783 231
rect 3787 227 3788 231
rect 3782 226 3788 227
rect 3030 221 3036 222
rect 3030 217 3031 221
rect 3035 217 3036 221
rect 3030 216 3036 217
rect 3002 211 3008 212
rect 3002 207 3003 211
rect 3007 207 3008 211
rect 3002 206 3008 207
rect 2930 203 2936 204
rect 2930 199 2931 203
rect 2935 199 2936 203
rect 2930 198 2936 199
rect 3032 163 3034 216
rect 3108 204 3110 226
rect 3214 221 3220 222
rect 3214 217 3215 221
rect 3219 217 3220 221
rect 3214 216 3220 217
rect 3106 203 3112 204
rect 3106 199 3107 203
rect 3111 199 3112 203
rect 3106 198 3112 199
rect 3216 163 3218 216
rect 3292 204 3294 226
rect 3290 203 3296 204
rect 3290 199 3291 203
rect 3295 199 3296 203
rect 3290 198 3296 199
rect 3380 164 3382 226
rect 3406 221 3412 222
rect 3406 217 3407 221
rect 3411 217 3412 221
rect 3406 216 3412 217
rect 3606 221 3612 222
rect 3606 217 3607 221
rect 3611 217 3612 221
rect 3606 216 3612 217
rect 3378 163 3384 164
rect 3408 163 3410 216
rect 3608 163 3610 216
rect 2743 162 2747 163
rect 2743 157 2747 158
rect 2855 162 2859 163
rect 2855 157 2859 158
rect 2871 162 2875 163
rect 2871 157 2875 158
rect 2991 162 2995 163
rect 2991 157 2995 158
rect 3031 162 3035 163
rect 3031 157 3035 158
rect 3111 162 3115 163
rect 3111 157 3115 158
rect 3215 162 3219 163
rect 3215 157 3219 158
rect 3223 162 3227 163
rect 3223 157 3227 158
rect 3327 162 3331 163
rect 3378 159 3379 163
rect 3383 159 3384 163
rect 3378 158 3384 159
rect 3407 162 3411 163
rect 3327 157 3331 158
rect 3407 157 3411 158
rect 3431 162 3435 163
rect 3431 157 3435 158
rect 3535 162 3539 163
rect 3535 157 3539 158
rect 3607 162 3611 163
rect 3607 157 3611 158
rect 3639 162 3643 163
rect 3639 157 3643 158
rect 3743 162 3747 163
rect 3743 157 3747 158
rect 2744 136 2746 157
rect 2872 136 2874 157
rect 2946 155 2952 156
rect 2946 151 2947 155
rect 2951 151 2952 155
rect 2946 150 2952 151
rect 2742 135 2748 136
rect 2742 131 2743 135
rect 2747 131 2748 135
rect 2742 130 2748 131
rect 2870 135 2876 136
rect 2870 131 2871 135
rect 2875 131 2876 135
rect 2870 130 2876 131
rect 2948 128 2950 150
rect 2992 136 2994 157
rect 3066 155 3072 156
rect 3066 151 3067 155
rect 3071 151 3072 155
rect 3066 150 3072 151
rect 2990 135 2996 136
rect 2990 131 2991 135
rect 2995 131 2996 135
rect 2990 130 2996 131
rect 3068 128 3070 150
rect 3112 136 3114 157
rect 3186 155 3192 156
rect 3186 151 3187 155
rect 3191 151 3192 155
rect 3186 150 3192 151
rect 3110 135 3116 136
rect 3110 131 3111 135
rect 3115 131 3116 135
rect 3110 130 3116 131
rect 3188 128 3190 150
rect 3224 136 3226 157
rect 3298 155 3304 156
rect 3298 151 3299 155
rect 3303 151 3304 155
rect 3298 150 3304 151
rect 3222 135 3228 136
rect 3222 131 3223 135
rect 3227 131 3228 135
rect 3222 130 3228 131
rect 3300 128 3302 150
rect 3328 136 3330 157
rect 3432 136 3434 157
rect 3506 155 3512 156
rect 3506 151 3507 155
rect 3511 151 3512 155
rect 3506 150 3512 151
rect 3326 135 3332 136
rect 3326 131 3327 135
rect 3331 131 3332 135
rect 3326 130 3332 131
rect 3430 135 3436 136
rect 3430 131 3431 135
rect 3435 131 3436 135
rect 3430 130 3436 131
rect 3508 128 3510 150
rect 3536 136 3538 157
rect 3640 136 3642 157
rect 3744 136 3746 157
rect 3784 156 3786 226
rect 3806 221 3812 222
rect 3806 217 3807 221
rect 3811 217 3812 221
rect 3806 216 3812 217
rect 3808 163 3810 216
rect 3868 204 3870 302
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3944 271 3946 298
rect 3943 270 3947 271
rect 3943 265 3947 266
rect 3944 238 3946 265
rect 3942 237 3948 238
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 3942 215 3948 216
rect 3866 203 3872 204
rect 3866 199 3867 203
rect 3871 199 3872 203
rect 3866 198 3872 199
rect 3944 163 3946 215
rect 3807 162 3811 163
rect 3807 157 3811 158
rect 3839 162 3843 163
rect 3839 157 3843 158
rect 3943 162 3947 163
rect 3943 157 3947 158
rect 3782 155 3788 156
rect 3782 151 3783 155
rect 3787 151 3788 155
rect 3782 150 3788 151
rect 3818 155 3824 156
rect 3818 151 3819 155
rect 3823 151 3824 155
rect 3818 150 3824 151
rect 3534 135 3540 136
rect 3534 131 3535 135
rect 3539 131 3540 135
rect 3534 130 3540 131
rect 3638 135 3644 136
rect 3638 131 3639 135
rect 3643 131 3644 135
rect 3638 130 3644 131
rect 3742 135 3748 136
rect 3742 131 3743 135
rect 3747 131 3748 135
rect 3742 130 3748 131
rect 3820 128 3822 150
rect 3840 136 3842 157
rect 3944 137 3946 157
rect 3942 136 3948 137
rect 3838 135 3844 136
rect 3838 131 3839 135
rect 3843 131 3844 135
rect 3942 132 3943 136
rect 3947 132 3948 136
rect 3942 131 3948 132
rect 3838 130 3844 131
rect 1978 126 1984 127
rect 2146 127 2152 128
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 112 91 114 118
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2146 123 2147 127
rect 2151 123 2152 127
rect 2146 122 2152 123
rect 2242 127 2248 128
rect 2242 123 2243 127
rect 2247 123 2248 127
rect 2242 122 2248 123
rect 2338 127 2344 128
rect 2338 123 2339 127
rect 2343 123 2344 127
rect 2338 122 2344 123
rect 2442 127 2448 128
rect 2442 123 2443 127
rect 2447 123 2448 127
rect 2442 122 2448 123
rect 2562 127 2568 128
rect 2562 123 2563 127
rect 2567 123 2568 127
rect 2562 122 2568 123
rect 2718 127 2724 128
rect 2718 123 2719 127
rect 2723 123 2724 127
rect 2718 122 2724 123
rect 2726 127 2732 128
rect 2726 123 2727 127
rect 2731 123 2732 127
rect 2726 122 2732 123
rect 2946 127 2952 128
rect 2946 123 2947 127
rect 2951 123 2952 127
rect 2946 122 2952 123
rect 3066 127 3072 128
rect 3066 123 3067 127
rect 3071 123 3072 127
rect 3066 122 3072 123
rect 3186 127 3192 128
rect 3186 123 3187 127
rect 3191 123 3192 127
rect 3186 122 3192 123
rect 3298 127 3304 128
rect 3298 123 3299 127
rect 3303 123 3304 127
rect 3298 122 3304 123
rect 3506 127 3512 128
rect 3506 123 3507 127
rect 3511 123 3512 127
rect 3506 122 3512 123
rect 3818 127 3824 128
rect 3818 123 3819 127
rect 3823 123 3824 127
rect 3818 122 3824 123
rect 2006 118 2012 119
rect 2046 119 2052 120
rect 1902 115 1908 116
rect 136 91 138 115
rect 232 91 234 115
rect 328 91 330 115
rect 424 91 426 115
rect 528 91 530 115
rect 648 91 650 115
rect 776 91 778 115
rect 904 91 906 115
rect 1032 91 1034 115
rect 1152 91 1154 115
rect 1272 91 1274 115
rect 1384 91 1386 115
rect 1488 91 1490 115
rect 1592 91 1594 115
rect 1704 91 1706 115
rect 1808 91 1810 115
rect 1904 91 1906 115
rect 2008 91 2010 118
rect 2046 115 2047 119
rect 2051 115 2052 119
rect 3942 119 3948 120
rect 2046 114 2052 115
rect 2070 116 2076 117
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 231 90 235 91
rect 231 85 235 86
rect 327 90 331 91
rect 327 85 331 86
rect 423 90 427 91
rect 423 85 427 86
rect 527 90 531 91
rect 527 85 531 86
rect 647 90 651 91
rect 647 85 651 86
rect 775 90 779 91
rect 775 85 779 86
rect 903 90 907 91
rect 903 85 907 86
rect 1031 90 1035 91
rect 1031 85 1035 86
rect 1151 90 1155 91
rect 1151 85 1155 86
rect 1271 90 1275 91
rect 1271 85 1275 86
rect 1383 90 1387 91
rect 1383 85 1387 86
rect 1487 90 1491 91
rect 1487 85 1491 86
rect 1591 90 1595 91
rect 1591 85 1595 86
rect 1703 90 1707 91
rect 1703 85 1707 86
rect 1807 90 1811 91
rect 1807 85 1811 86
rect 1903 90 1907 91
rect 1903 85 1907 86
rect 2007 90 2011 91
rect 2048 87 2050 114
rect 2070 112 2071 116
rect 2075 112 2076 116
rect 2070 111 2076 112
rect 2166 116 2172 117
rect 2166 112 2167 116
rect 2171 112 2172 116
rect 2166 111 2172 112
rect 2262 116 2268 117
rect 2262 112 2263 116
rect 2267 112 2268 116
rect 2262 111 2268 112
rect 2366 116 2372 117
rect 2366 112 2367 116
rect 2371 112 2372 116
rect 2366 111 2372 112
rect 2486 116 2492 117
rect 2486 112 2487 116
rect 2491 112 2492 116
rect 2486 111 2492 112
rect 2614 116 2620 117
rect 2614 112 2615 116
rect 2619 112 2620 116
rect 2614 111 2620 112
rect 2742 116 2748 117
rect 2742 112 2743 116
rect 2747 112 2748 116
rect 2742 111 2748 112
rect 2870 116 2876 117
rect 2870 112 2871 116
rect 2875 112 2876 116
rect 2870 111 2876 112
rect 2990 116 2996 117
rect 2990 112 2991 116
rect 2995 112 2996 116
rect 2990 111 2996 112
rect 3110 116 3116 117
rect 3110 112 3111 116
rect 3115 112 3116 116
rect 3110 111 3116 112
rect 3222 116 3228 117
rect 3222 112 3223 116
rect 3227 112 3228 116
rect 3222 111 3228 112
rect 3326 116 3332 117
rect 3326 112 3327 116
rect 3331 112 3332 116
rect 3326 111 3332 112
rect 3430 116 3436 117
rect 3430 112 3431 116
rect 3435 112 3436 116
rect 3430 111 3436 112
rect 3534 116 3540 117
rect 3534 112 3535 116
rect 3539 112 3540 116
rect 3534 111 3540 112
rect 3638 116 3644 117
rect 3638 112 3639 116
rect 3643 112 3644 116
rect 3638 111 3644 112
rect 3742 116 3748 117
rect 3742 112 3743 116
rect 3747 112 3748 116
rect 3742 111 3748 112
rect 3838 116 3844 117
rect 3838 112 3839 116
rect 3843 112 3844 116
rect 3942 115 3943 119
rect 3947 115 3948 119
rect 3942 114 3948 115
rect 3838 111 3844 112
rect 2072 87 2074 111
rect 2168 87 2170 111
rect 2264 87 2266 111
rect 2368 87 2370 111
rect 2488 87 2490 111
rect 2616 87 2618 111
rect 2744 87 2746 111
rect 2872 87 2874 111
rect 2992 87 2994 111
rect 3112 87 3114 111
rect 3224 87 3226 111
rect 3328 87 3330 111
rect 3432 87 3434 111
rect 3536 87 3538 111
rect 3640 87 3642 111
rect 3744 87 3746 111
rect 3840 87 3842 111
rect 3944 87 3946 114
rect 2007 85 2011 86
rect 2047 86 2051 87
rect 2047 81 2051 82
rect 2071 86 2075 87
rect 2071 81 2075 82
rect 2167 86 2171 87
rect 2167 81 2171 82
rect 2263 86 2267 87
rect 2263 81 2267 82
rect 2367 86 2371 87
rect 2367 81 2371 82
rect 2487 86 2491 87
rect 2487 81 2491 82
rect 2615 86 2619 87
rect 2615 81 2619 82
rect 2743 86 2747 87
rect 2743 81 2747 82
rect 2871 86 2875 87
rect 2871 81 2875 82
rect 2991 86 2995 87
rect 2991 81 2995 82
rect 3111 86 3115 87
rect 3111 81 3115 82
rect 3223 86 3227 87
rect 3223 81 3227 82
rect 3327 86 3331 87
rect 3327 81 3331 82
rect 3431 86 3435 87
rect 3431 81 3435 82
rect 3535 86 3539 87
rect 3535 81 3539 82
rect 3639 86 3643 87
rect 3639 81 3643 82
rect 3743 86 3747 87
rect 3743 81 3747 82
rect 3839 86 3843 87
rect 3839 81 3843 82
rect 3943 86 3947 87
rect 3943 81 3947 82
<< m4c >>
rect 2047 4026 2051 4030
rect 2071 4026 2075 4030
rect 3943 4026 3947 4030
rect 111 4006 115 4010
rect 151 4006 155 4010
rect 279 4006 283 4010
rect 431 4006 435 4010
rect 607 4006 611 4010
rect 791 4006 795 4010
rect 975 4006 979 4010
rect 1151 4006 1155 4010
rect 1311 4006 1315 4010
rect 1471 4006 1475 4010
rect 1623 4006 1627 4010
rect 1775 4006 1779 4010
rect 1903 4006 1907 4010
rect 111 3930 115 3934
rect 151 3930 155 3934
rect 279 3930 283 3934
rect 303 3930 307 3934
rect 423 3930 427 3934
rect 431 3930 435 3934
rect 551 3930 555 3934
rect 607 3930 611 3934
rect 687 3930 691 3934
rect 791 3930 795 3934
rect 815 3930 819 3934
rect 943 3930 947 3934
rect 975 3930 979 3934
rect 1071 3930 1075 3934
rect 1151 3930 1155 3934
rect 1199 3930 1203 3934
rect 1311 3930 1315 3934
rect 1327 3930 1331 3934
rect 2007 4006 2011 4010
rect 2047 3950 2051 3954
rect 2071 3950 2075 3954
rect 2079 3950 2083 3954
rect 1463 3930 1467 3934
rect 1471 3930 1475 3934
rect 1623 3930 1627 3934
rect 1775 3930 1779 3934
rect 1903 3930 1907 3934
rect 2007 3930 2011 3934
rect 111 3850 115 3854
rect 303 3850 307 3854
rect 415 3850 419 3854
rect 423 3850 427 3854
rect 551 3850 555 3854
rect 567 3850 571 3854
rect 687 3850 691 3854
rect 727 3850 731 3854
rect 815 3850 819 3854
rect 887 3850 891 3854
rect 943 3850 947 3854
rect 2215 3950 2219 3954
rect 2359 3950 2363 3954
rect 2503 3950 2507 3954
rect 2647 3950 2651 3954
rect 2791 3950 2795 3954
rect 2927 3950 2931 3954
rect 3055 3950 3059 3954
rect 3175 3950 3179 3954
rect 3295 3950 3299 3954
rect 3415 3950 3419 3954
rect 3535 3950 3539 3954
rect 3943 3950 3947 3954
rect 2047 3874 2051 3878
rect 2079 3874 2083 3878
rect 2215 3874 2219 3878
rect 2255 3874 2259 3878
rect 2359 3874 2363 3878
rect 2383 3874 2387 3878
rect 2503 3874 2507 3878
rect 2519 3874 2523 3878
rect 2647 3874 2651 3878
rect 2671 3874 2675 3878
rect 1039 3850 1043 3854
rect 1071 3850 1075 3854
rect 1191 3850 1195 3854
rect 1199 3850 1203 3854
rect 1327 3850 1331 3854
rect 1343 3850 1347 3854
rect 1463 3850 1467 3854
rect 1495 3850 1499 3854
rect 1647 3850 1651 3854
rect 2007 3850 2011 3854
rect 111 3770 115 3774
rect 399 3770 403 3774
rect 415 3770 419 3774
rect 567 3770 571 3774
rect 727 3770 731 3774
rect 751 3770 755 3774
rect 887 3770 891 3774
rect 935 3770 939 3774
rect 1039 3770 1043 3774
rect 1127 3770 1131 3774
rect 1191 3770 1195 3774
rect 1311 3770 1315 3774
rect 1343 3770 1347 3774
rect 1495 3770 1499 3774
rect 1503 3770 1507 3774
rect 2791 3874 2795 3878
rect 2831 3874 2835 3878
rect 2927 3874 2931 3878
rect 2991 3874 2995 3878
rect 3055 3874 3059 3878
rect 3159 3874 3163 3878
rect 2047 3798 2051 3802
rect 2071 3798 2075 3802
rect 2199 3798 2203 3802
rect 2255 3798 2259 3802
rect 2375 3798 2379 3802
rect 2383 3798 2387 3802
rect 2519 3798 2523 3802
rect 2559 3798 2563 3802
rect 1647 3770 1651 3774
rect 1695 3770 1699 3774
rect 1887 3770 1891 3774
rect 2007 3770 2011 3774
rect 111 3682 115 3686
rect 367 3682 371 3686
rect 399 3682 403 3686
rect 519 3682 523 3686
rect 567 3682 571 3686
rect 679 3682 683 3686
rect 751 3682 755 3686
rect 847 3682 851 3686
rect 935 3682 939 3686
rect 1015 3682 1019 3686
rect 1127 3682 1131 3686
rect 1175 3682 1179 3686
rect 1311 3682 1315 3686
rect 1327 3682 1331 3686
rect 1479 3682 1483 3686
rect 111 3598 115 3602
rect 271 3598 275 3602
rect 367 3598 371 3602
rect 415 3598 419 3602
rect 519 3598 523 3602
rect 575 3598 579 3602
rect 111 3514 115 3518
rect 159 3514 163 3518
rect 271 3514 275 3518
rect 287 3514 291 3518
rect 415 3514 419 3518
rect 423 3514 427 3518
rect 679 3598 683 3602
rect 735 3598 739 3602
rect 847 3598 851 3602
rect 895 3598 899 3602
rect 1015 3598 1019 3602
rect 1055 3598 1059 3602
rect 1175 3598 1179 3602
rect 1215 3598 1219 3602
rect 1327 3598 1331 3602
rect 1375 3598 1379 3602
rect 1503 3682 1507 3686
rect 1631 3682 1635 3686
rect 1695 3682 1699 3686
rect 1791 3682 1795 3686
rect 2047 3710 2051 3714
rect 2071 3710 2075 3714
rect 2671 3798 2675 3802
rect 2751 3798 2755 3802
rect 2831 3798 2835 3802
rect 2951 3798 2955 3802
rect 2991 3798 2995 3802
rect 3175 3874 3179 3878
rect 3295 3874 3299 3878
rect 3327 3874 3331 3878
rect 3415 3874 3419 3878
rect 3495 3874 3499 3878
rect 3535 3874 3539 3878
rect 3663 3874 3667 3878
rect 3943 3874 3947 3878
rect 3143 3798 3147 3802
rect 3159 3798 3163 3802
rect 3327 3798 3331 3802
rect 3335 3798 3339 3802
rect 2199 3710 2203 3714
rect 2263 3710 2267 3714
rect 2375 3710 2379 3714
rect 2479 3710 2483 3714
rect 2559 3710 2563 3714
rect 2695 3710 2699 3714
rect 2751 3710 2755 3714
rect 2911 3710 2915 3714
rect 2951 3710 2955 3714
rect 3119 3710 3123 3714
rect 3143 3710 3147 3714
rect 1887 3682 1891 3686
rect 2007 3682 2011 3686
rect 2047 3630 2051 3634
rect 2071 3630 2075 3634
rect 2111 3630 2115 3634
rect 2263 3630 2267 3634
rect 2271 3630 2275 3634
rect 2455 3630 2459 3634
rect 2479 3630 2483 3634
rect 2655 3630 2659 3634
rect 1479 3598 1483 3602
rect 1543 3598 1547 3602
rect 1631 3598 1635 3602
rect 1791 3598 1795 3602
rect 2007 3598 2011 3602
rect 559 3514 563 3518
rect 575 3514 579 3518
rect 695 3514 699 3518
rect 735 3514 739 3518
rect 831 3514 835 3518
rect 895 3514 899 3518
rect 967 3514 971 3518
rect 1055 3514 1059 3518
rect 1095 3514 1099 3518
rect 1215 3514 1219 3518
rect 1231 3514 1235 3518
rect 111 3430 115 3434
rect 135 3430 139 3434
rect 159 3430 163 3434
rect 247 3430 251 3434
rect 287 3430 291 3434
rect 111 3346 115 3350
rect 135 3346 139 3350
rect 383 3430 387 3434
rect 423 3430 427 3434
rect 527 3430 531 3434
rect 559 3430 563 3434
rect 671 3430 675 3434
rect 695 3430 699 3434
rect 815 3430 819 3434
rect 831 3430 835 3434
rect 2695 3630 2699 3634
rect 2871 3630 2875 3634
rect 2911 3630 2915 3634
rect 3495 3798 3499 3802
rect 3535 3798 3539 3802
rect 3663 3798 3667 3802
rect 3735 3798 3739 3802
rect 3943 3798 3947 3802
rect 3319 3710 3323 3714
rect 3335 3710 3339 3714
rect 3519 3710 3523 3714
rect 3535 3710 3539 3714
rect 3727 3710 3731 3714
rect 3735 3710 3739 3714
rect 3943 3710 3947 3714
rect 3095 3630 3099 3634
rect 3119 3630 3123 3634
rect 3319 3630 3323 3634
rect 3327 3630 3331 3634
rect 3519 3630 3523 3634
rect 3567 3630 3571 3634
rect 2047 3538 2051 3542
rect 2111 3538 2115 3542
rect 2271 3538 2275 3542
rect 2287 3538 2291 3542
rect 2383 3538 2387 3542
rect 2455 3538 2459 3542
rect 2479 3538 2483 3542
rect 2575 3538 2579 3542
rect 2655 3538 2659 3542
rect 2671 3538 2675 3542
rect 2767 3538 2771 3542
rect 1367 3514 1371 3518
rect 1375 3514 1379 3518
rect 1543 3514 1547 3518
rect 2007 3514 2011 3518
rect 2355 3496 2359 3500
rect 2871 3538 2875 3542
rect 2983 3538 2987 3542
rect 3095 3538 3099 3542
rect 3103 3538 3107 3542
rect 3223 3538 3227 3542
rect 3327 3538 3331 3542
rect 3351 3538 3355 3542
rect 2047 3462 2051 3466
rect 2287 3462 2291 3466
rect 2383 3462 2387 3466
rect 2479 3462 2483 3466
rect 2487 3462 2491 3466
rect 967 3430 971 3434
rect 1095 3430 1099 3434
rect 1119 3430 1123 3434
rect 1231 3430 1235 3434
rect 1271 3430 1275 3434
rect 1367 3430 1371 3434
rect 2007 3430 2011 3434
rect 2575 3462 2579 3466
rect 2583 3462 2587 3466
rect 2671 3462 2675 3466
rect 2679 3462 2683 3466
rect 2863 3496 2867 3500
rect 2767 3462 2771 3466
rect 2783 3462 2787 3466
rect 2871 3462 2875 3466
rect 2895 3462 2899 3466
rect 2983 3462 2987 3466
rect 3015 3462 3019 3466
rect 3103 3462 3107 3466
rect 3143 3462 3147 3466
rect 3223 3462 3227 3466
rect 3727 3630 3731 3634
rect 3943 3630 3947 3634
rect 3487 3538 3491 3542
rect 3567 3538 3571 3542
rect 3943 3538 3947 3542
rect 3271 3462 3275 3466
rect 3351 3462 3355 3466
rect 3407 3462 3411 3466
rect 247 3346 251 3350
rect 263 3346 267 3350
rect 383 3346 387 3350
rect 431 3346 435 3350
rect 527 3346 531 3350
rect 599 3346 603 3350
rect 671 3346 675 3350
rect 767 3346 771 3350
rect 815 3346 819 3350
rect 927 3346 931 3350
rect 967 3346 971 3350
rect 1087 3346 1091 3350
rect 1119 3346 1123 3350
rect 2047 3378 2051 3382
rect 2351 3378 2355 3382
rect 2479 3378 2483 3382
rect 2487 3378 2491 3382
rect 2583 3378 2587 3382
rect 2615 3378 2619 3382
rect 2679 3378 2683 3382
rect 2751 3378 2755 3382
rect 2783 3378 2787 3382
rect 2887 3378 2891 3382
rect 2895 3378 2899 3382
rect 3015 3378 3019 3382
rect 3023 3378 3027 3382
rect 1239 3346 1243 3350
rect 1271 3346 1275 3350
rect 1391 3346 1395 3350
rect 1551 3346 1555 3350
rect 2007 3346 2011 3350
rect 111 3262 115 3266
rect 135 3262 139 3266
rect 143 3262 147 3266
rect 263 3262 267 3266
rect 295 3262 299 3266
rect 431 3262 435 3266
rect 455 3262 459 3266
rect 599 3262 603 3266
rect 623 3262 627 3266
rect 183 3200 187 3204
rect 767 3262 771 3266
rect 791 3262 795 3266
rect 927 3262 931 3266
rect 959 3262 963 3266
rect 1087 3262 1091 3266
rect 1127 3262 1131 3266
rect 1239 3262 1243 3266
rect 1303 3262 1307 3266
rect 1391 3262 1395 3266
rect 1479 3262 1483 3266
rect 1551 3262 1555 3266
rect 2047 3298 2051 3302
rect 2127 3298 2131 3302
rect 2295 3298 2299 3302
rect 2351 3298 2355 3302
rect 2455 3298 2459 3302
rect 2479 3298 2483 3302
rect 2615 3298 2619 3302
rect 2007 3262 2011 3266
rect 2047 3222 2051 3226
rect 739 3200 743 3204
rect 2071 3222 2075 3226
rect 2127 3222 2131 3226
rect 2207 3222 2211 3226
rect 2751 3298 2755 3302
rect 2775 3298 2779 3302
rect 3143 3378 3147 3382
rect 3159 3378 3163 3382
rect 3271 3378 3275 3382
rect 3303 3378 3307 3382
rect 3487 3462 3491 3466
rect 3943 3462 3947 3466
rect 3407 3378 3411 3382
rect 3943 3378 3947 3382
rect 2887 3298 2891 3302
rect 2935 3298 2939 3302
rect 3023 3298 3027 3302
rect 3095 3298 3099 3302
rect 3159 3298 3163 3302
rect 2295 3222 2299 3226
rect 2375 3222 2379 3226
rect 2455 3222 2459 3226
rect 2543 3222 2547 3226
rect 2615 3222 2619 3226
rect 2703 3222 2707 3226
rect 2775 3222 2779 3226
rect 2863 3222 2867 3226
rect 2935 3222 2939 3226
rect 3015 3222 3019 3226
rect 111 3186 115 3190
rect 143 3186 147 3190
rect 295 3186 299 3190
rect 431 3186 435 3190
rect 455 3186 459 3190
rect 567 3186 571 3190
rect 623 3186 627 3190
rect 703 3186 707 3190
rect 791 3186 795 3190
rect 855 3186 859 3190
rect 959 3186 963 3190
rect 1031 3186 1035 3190
rect 1127 3186 1131 3190
rect 1231 3186 1235 3190
rect 1303 3186 1307 3190
rect 1455 3186 1459 3190
rect 1479 3186 1483 3190
rect 1687 3186 1691 3190
rect 111 3110 115 3114
rect 295 3110 299 3114
rect 311 3110 315 3114
rect 407 3110 411 3114
rect 431 3110 435 3114
rect 503 3110 507 3114
rect 567 3110 571 3114
rect 599 3110 603 3114
rect 695 3110 699 3114
rect 703 3110 707 3114
rect 807 3110 811 3114
rect 855 3110 859 3114
rect 1903 3186 1907 3190
rect 2007 3186 2011 3190
rect 943 3110 947 3114
rect 1031 3110 1035 3114
rect 1087 3110 1091 3114
rect 1231 3110 1235 3114
rect 1247 3110 1251 3114
rect 1407 3110 1411 3114
rect 1455 3110 1459 3114
rect 1575 3110 1579 3114
rect 1687 3110 1691 3114
rect 1751 3110 1755 3114
rect 1903 3110 1907 3114
rect 2047 3142 2051 3146
rect 463 3048 467 3052
rect 111 3034 115 3038
rect 311 3034 315 3038
rect 407 3034 411 3038
rect 423 3034 427 3038
rect 779 3048 783 3052
rect 503 3034 507 3038
rect 519 3034 523 3038
rect 599 3034 603 3038
rect 615 3034 619 3038
rect 695 3034 699 3038
rect 711 3034 715 3038
rect 807 3034 811 3038
rect 815 3034 819 3038
rect 935 3034 939 3038
rect 943 3034 947 3038
rect 1055 3034 1059 3038
rect 1087 3034 1091 3038
rect 1183 3034 1187 3038
rect 1247 3034 1251 3038
rect 1311 3034 1315 3038
rect 1407 3034 1411 3038
rect 1431 3034 1435 3038
rect 1551 3034 1555 3038
rect 1575 3034 1579 3038
rect 1671 3034 1675 3038
rect 1751 3034 1755 3038
rect 1799 3034 1803 3038
rect 2071 3142 2075 3146
rect 2007 3110 2011 3114
rect 2207 3142 2211 3146
rect 2343 3142 2347 3146
rect 2375 3142 2379 3146
rect 2543 3142 2547 3146
rect 2631 3142 2635 3146
rect 2703 3142 2707 3146
rect 3263 3298 3267 3302
rect 3303 3298 3307 3302
rect 3943 3298 3947 3302
rect 3095 3222 3099 3226
rect 3167 3222 3171 3226
rect 3263 3222 3267 3226
rect 3327 3222 3331 3226
rect 3943 3222 3947 3226
rect 2863 3142 2867 3146
rect 2903 3142 2907 3146
rect 3015 3142 3019 3146
rect 3167 3142 3171 3146
rect 3175 3142 3179 3146
rect 3327 3142 3331 3146
rect 2047 3062 2051 3066
rect 2071 3062 2075 3066
rect 2343 3062 2347 3066
rect 2487 3062 2491 3066
rect 2615 3062 2619 3066
rect 2631 3062 2635 3066
rect 2743 3062 2747 3066
rect 1903 3034 1907 3038
rect 2007 3034 2011 3038
rect 111 2934 115 2938
rect 423 2934 427 2938
rect 519 2934 523 2938
rect 615 2934 619 2938
rect 711 2934 715 2938
rect 815 2934 819 2938
rect 935 2934 939 2938
rect 1055 2934 1059 2938
rect 1183 2934 1187 2938
rect 1311 2934 1315 2938
rect 1431 2934 1435 2938
rect 1479 2934 1483 2938
rect 2047 2982 2051 2986
rect 2407 2982 2411 2986
rect 2487 2982 2491 2986
rect 2863 3062 2867 3066
rect 2903 3062 2907 3066
rect 2983 3062 2987 3066
rect 3447 3142 3451 3146
rect 3943 3142 3947 3146
rect 3103 3062 3107 3066
rect 3175 3062 3179 3066
rect 3215 3062 3219 3066
rect 3327 3062 3331 3066
rect 3431 3062 3435 3066
rect 3447 3062 3451 3066
rect 3535 3062 3539 3066
rect 3639 3062 3643 3066
rect 3743 3062 3747 3066
rect 3839 3062 3843 3066
rect 3943 3062 3947 3066
rect 2575 2982 2579 2986
rect 2615 2982 2619 2986
rect 2743 2982 2747 2986
rect 2767 2982 2771 2986
rect 2863 2982 2867 2986
rect 2967 2982 2971 2986
rect 2983 2982 2987 2986
rect 3103 2982 3107 2986
rect 3183 2982 3187 2986
rect 3215 2982 3219 2986
rect 3327 2982 3331 2986
rect 3399 2982 3403 2986
rect 3431 2982 3435 2986
rect 3535 2982 3539 2986
rect 3623 2982 3627 2986
rect 3639 2982 3643 2986
rect 3743 2982 3747 2986
rect 3839 2982 3843 2986
rect 1551 2934 1555 2938
rect 1575 2934 1579 2938
rect 1671 2934 1675 2938
rect 1767 2934 1771 2938
rect 1799 2934 1803 2938
rect 1863 2934 1867 2938
rect 1903 2934 1907 2938
rect 2007 2934 2011 2938
rect 111 2850 115 2854
rect 279 2850 283 2854
rect 447 2850 451 2854
rect 631 2850 635 2854
rect 815 2850 819 2854
rect 999 2850 1003 2854
rect 1183 2850 1187 2854
rect 1359 2850 1363 2854
rect 1479 2850 1483 2854
rect 1527 2850 1531 2854
rect 1575 2850 1579 2854
rect 1671 2850 1675 2854
rect 1695 2850 1699 2854
rect 1767 2850 1771 2854
rect 1863 2850 1867 2854
rect 111 2774 115 2778
rect 239 2774 243 2778
rect 279 2774 283 2778
rect 351 2774 355 2778
rect 2047 2890 2051 2894
rect 2407 2890 2411 2894
rect 2551 2890 2555 2894
rect 2575 2890 2579 2894
rect 2671 2890 2675 2894
rect 2767 2890 2771 2894
rect 2799 2890 2803 2894
rect 2927 2890 2931 2894
rect 2967 2890 2971 2894
rect 3055 2890 3059 2894
rect 2007 2850 2011 2854
rect 447 2774 451 2778
rect 471 2774 475 2778
rect 607 2774 611 2778
rect 631 2774 635 2778
rect 743 2774 747 2778
rect 815 2774 819 2778
rect 879 2774 883 2778
rect 111 2698 115 2702
rect 223 2698 227 2702
rect 239 2698 243 2702
rect 351 2698 355 2702
rect 367 2698 371 2702
rect 471 2698 475 2702
rect 503 2698 507 2702
rect 111 2622 115 2626
rect 175 2622 179 2626
rect 223 2622 227 2626
rect 367 2622 371 2626
rect 2047 2814 2051 2818
rect 2439 2814 2443 2818
rect 2551 2814 2555 2818
rect 2567 2814 2571 2818
rect 2671 2814 2675 2818
rect 2695 2814 2699 2818
rect 2799 2814 2803 2818
rect 2831 2814 2835 2818
rect 999 2774 1003 2778
rect 1015 2774 1019 2778
rect 1151 2774 1155 2778
rect 1183 2774 1187 2778
rect 1287 2774 1291 2778
rect 1359 2774 1363 2778
rect 1423 2774 1427 2778
rect 607 2698 611 2702
rect 639 2698 643 2702
rect 743 2698 747 2702
rect 767 2698 771 2702
rect 879 2698 883 2702
rect 887 2698 891 2702
rect 999 2698 1003 2702
rect 1015 2698 1019 2702
rect 1111 2698 1115 2702
rect 1151 2698 1155 2702
rect 1231 2698 1235 2702
rect 3943 2982 3947 2986
rect 3183 2890 3187 2894
rect 3311 2890 3315 2894
rect 3399 2890 3403 2894
rect 3439 2890 3443 2894
rect 3575 2890 3579 2894
rect 3623 2890 3627 2894
rect 3839 2890 3843 2894
rect 2927 2814 2931 2818
rect 2967 2814 2971 2818
rect 3055 2814 3059 2818
rect 3103 2814 3107 2818
rect 1527 2774 1531 2778
rect 1567 2774 1571 2778
rect 1695 2774 1699 2778
rect 1863 2774 1867 2778
rect 2007 2774 2011 2778
rect 3183 2814 3187 2818
rect 3247 2814 3251 2818
rect 3311 2814 3315 2818
rect 3391 2814 3395 2818
rect 3439 2814 3443 2818
rect 3543 2814 3547 2818
rect 3575 2814 3579 2818
rect 3703 2814 3707 2818
rect 3839 2814 3843 2818
rect 2047 2730 2051 2734
rect 2335 2730 2339 2734
rect 2439 2730 2443 2734
rect 2495 2730 2499 2734
rect 2567 2730 2571 2734
rect 2663 2730 2667 2734
rect 2695 2730 2699 2734
rect 2831 2730 2835 2734
rect 2967 2730 2971 2734
rect 2999 2730 3003 2734
rect 3103 2730 3107 2734
rect 3167 2730 3171 2734
rect 3247 2730 3251 2734
rect 1287 2698 1291 2702
rect 1351 2698 1355 2702
rect 1423 2698 1427 2702
rect 1567 2698 1571 2702
rect 2007 2698 2011 2702
rect 503 2622 507 2626
rect 543 2622 547 2626
rect 639 2622 643 2626
rect 711 2622 715 2626
rect 111 2542 115 2546
rect 135 2542 139 2546
rect 175 2542 179 2546
rect 271 2542 275 2546
rect 367 2542 371 2546
rect 439 2542 443 2546
rect 543 2542 547 2546
rect 607 2542 611 2546
rect 111 2462 115 2466
rect 135 2462 139 2466
rect 271 2462 275 2466
rect 311 2462 315 2466
rect 439 2462 443 2466
rect 767 2622 771 2626
rect 863 2622 867 2626
rect 2047 2650 2051 2654
rect 2127 2650 2131 2654
rect 2279 2650 2283 2654
rect 2335 2650 2339 2654
rect 887 2622 891 2626
rect 999 2622 1003 2626
rect 1007 2622 1011 2626
rect 1111 2622 1115 2626
rect 1143 2622 1147 2626
rect 1231 2622 1235 2626
rect 1279 2622 1283 2626
rect 1351 2622 1355 2626
rect 1423 2622 1427 2626
rect 2007 2622 2011 2626
rect 3335 2730 3339 2734
rect 3391 2730 3395 2734
rect 3511 2730 3515 2734
rect 3543 2730 3547 2734
rect 3687 2730 3691 2734
rect 3703 2730 3707 2734
rect 3839 2730 3843 2734
rect 3943 2890 3947 2894
rect 3943 2814 3947 2818
rect 3943 2730 3947 2734
rect 2447 2650 2451 2654
rect 2495 2650 2499 2654
rect 2623 2650 2627 2654
rect 2663 2650 2667 2654
rect 2807 2650 2811 2654
rect 2831 2650 2835 2654
rect 2991 2650 2995 2654
rect 2999 2650 3003 2654
rect 3167 2650 3171 2654
rect 3175 2650 3179 2654
rect 2167 2579 2171 2580
rect 2167 2576 2171 2579
rect 2599 2576 2603 2580
rect 2047 2566 2051 2570
rect 2071 2566 2075 2570
rect 2127 2566 2131 2570
rect 2183 2566 2187 2570
rect 2279 2566 2283 2570
rect 2319 2566 2323 2570
rect 2447 2566 2451 2570
rect 2471 2566 2475 2570
rect 711 2542 715 2546
rect 775 2542 779 2546
rect 863 2542 867 2546
rect 927 2542 931 2546
rect 1007 2542 1011 2546
rect 1079 2542 1083 2546
rect 1143 2542 1147 2546
rect 1223 2542 1227 2546
rect 1279 2542 1283 2546
rect 1359 2542 1363 2546
rect 1423 2542 1427 2546
rect 1495 2542 1499 2546
rect 1639 2542 1643 2546
rect 2007 2542 2011 2546
rect 511 2462 515 2466
rect 607 2462 611 2466
rect 711 2462 715 2466
rect 775 2462 779 2466
rect 903 2462 907 2466
rect 927 2462 931 2466
rect 111 2386 115 2390
rect 135 2386 139 2390
rect 311 2386 315 2390
rect 327 2386 331 2390
rect 511 2386 515 2390
rect 551 2386 555 2390
rect 111 2302 115 2306
rect 135 2302 139 2306
rect 271 2302 275 2306
rect 327 2302 331 2306
rect 1079 2462 1083 2466
rect 1223 2462 1227 2466
rect 1239 2462 1243 2466
rect 1359 2462 1363 2466
rect 1391 2462 1395 2466
rect 1495 2462 1499 2466
rect 1527 2462 1531 2466
rect 2047 2486 2051 2490
rect 2071 2486 2075 2490
rect 2183 2486 2187 2490
rect 2215 2486 2219 2490
rect 1639 2462 1643 2466
rect 1663 2462 1667 2466
rect 1791 2462 1795 2466
rect 1903 2462 1907 2466
rect 2007 2462 2011 2466
rect 2623 2566 2627 2570
rect 2639 2566 2643 2570
rect 2807 2566 2811 2570
rect 2823 2566 2827 2570
rect 3335 2650 3339 2654
rect 3351 2650 3355 2654
rect 3511 2650 3515 2654
rect 3519 2650 3523 2654
rect 3687 2650 3691 2654
rect 3839 2650 3843 2654
rect 2991 2566 2995 2570
rect 3031 2566 3035 2570
rect 3175 2566 3179 2570
rect 3263 2566 3267 2570
rect 3351 2566 3355 2570
rect 3503 2566 3507 2570
rect 3519 2566 3523 2570
rect 3687 2566 3691 2570
rect 2319 2486 2323 2490
rect 2383 2486 2387 2490
rect 2471 2486 2475 2490
rect 2559 2486 2563 2490
rect 2639 2486 2643 2490
rect 2751 2486 2755 2490
rect 2823 2486 2827 2490
rect 2951 2486 2955 2490
rect 3031 2486 3035 2490
rect 3167 2486 3171 2490
rect 3263 2486 3267 2490
rect 3391 2486 3395 2490
rect 2047 2394 2051 2398
rect 2071 2394 2075 2398
rect 2215 2394 2219 2398
rect 2247 2394 2251 2398
rect 2383 2394 2387 2398
rect 2431 2394 2435 2398
rect 711 2386 715 2390
rect 767 2386 771 2390
rect 903 2386 907 2390
rect 975 2386 979 2390
rect 1079 2386 1083 2390
rect 1175 2386 1179 2390
rect 1239 2386 1243 2390
rect 1367 2386 1371 2390
rect 1391 2386 1395 2390
rect 1527 2386 1531 2390
rect 1551 2386 1555 2390
rect 1663 2386 1667 2390
rect 1735 2386 1739 2390
rect 1791 2386 1795 2390
rect 1903 2386 1907 2390
rect 2007 2386 2011 2390
rect 431 2302 435 2306
rect 551 2302 555 2306
rect 591 2302 595 2306
rect 751 2302 755 2306
rect 767 2302 771 2306
rect 919 2302 923 2306
rect 111 2226 115 2230
rect 135 2226 139 2230
rect 159 2226 163 2230
rect 271 2226 275 2230
rect 327 2226 331 2230
rect 431 2226 435 2230
rect 495 2226 499 2230
rect 591 2226 595 2230
rect 975 2302 979 2306
rect 1087 2302 1091 2306
rect 1175 2302 1179 2306
rect 1263 2302 1267 2306
rect 1367 2302 1371 2306
rect 1447 2302 1451 2306
rect 1551 2302 1555 2306
rect 1631 2302 1635 2306
rect 679 2226 683 2230
rect 751 2226 755 2230
rect 879 2226 883 2230
rect 919 2226 923 2230
rect 111 2150 115 2154
rect 159 2150 163 2154
rect 223 2150 227 2154
rect 327 2150 331 2154
rect 359 2150 363 2154
rect 495 2150 499 2154
rect 1087 2226 1091 2230
rect 1095 2226 1099 2230
rect 1263 2226 1267 2230
rect 1327 2226 1331 2230
rect 1447 2226 1451 2230
rect 639 2150 643 2154
rect 679 2150 683 2154
rect 783 2150 787 2154
rect 111 2066 115 2070
rect 223 2066 227 2070
rect 359 2066 363 2070
rect 375 2066 379 2070
rect 495 2066 499 2070
rect 615 2066 619 2070
rect 639 2066 643 2070
rect 111 1982 115 1986
rect 375 1982 379 1986
rect 879 2150 883 2154
rect 935 2150 939 2154
rect 1095 2150 1099 2154
rect 2047 2318 2051 2322
rect 2071 2318 2075 2322
rect 2175 2318 2179 2322
rect 2247 2318 2251 2322
rect 1735 2302 1739 2306
rect 1815 2302 1819 2306
rect 1903 2302 1907 2306
rect 2007 2302 2011 2306
rect 3503 2486 3507 2490
rect 3623 2486 3627 2490
rect 3943 2650 3947 2654
rect 3743 2566 3747 2570
rect 3839 2566 3843 2570
rect 3743 2486 3747 2490
rect 3839 2486 3843 2490
rect 2559 2394 2563 2398
rect 2607 2394 2611 2398
rect 2751 2394 2755 2398
rect 2775 2394 2779 2398
rect 2935 2394 2939 2398
rect 2951 2394 2955 2398
rect 3103 2394 3107 2398
rect 3167 2394 3171 2398
rect 3391 2394 3395 2398
rect 3623 2394 3627 2398
rect 2311 2318 2315 2322
rect 2431 2318 2435 2322
rect 2447 2318 2451 2322
rect 2591 2318 2595 2322
rect 2607 2318 2611 2322
rect 2751 2318 2755 2322
rect 2775 2318 2779 2322
rect 2935 2318 2939 2322
rect 1567 2226 1571 2230
rect 1631 2226 1635 2230
rect 1815 2226 1819 2230
rect 2047 2234 2051 2238
rect 2071 2234 2075 2238
rect 2111 2234 2115 2238
rect 2175 2234 2179 2238
rect 2255 2234 2259 2238
rect 2311 2234 2315 2238
rect 2407 2234 2411 2238
rect 2447 2234 2451 2238
rect 2007 2226 2011 2230
rect 3103 2318 3107 2322
rect 3143 2318 3147 2322
rect 3375 2318 3379 2322
rect 3615 2318 3619 2322
rect 2559 2234 2563 2238
rect 2591 2234 2595 2238
rect 2719 2234 2723 2238
rect 2751 2234 2755 2238
rect 2879 2234 2883 2238
rect 2935 2234 2939 2238
rect 3047 2234 3051 2238
rect 3143 2234 3147 2238
rect 3223 2234 3227 2238
rect 3375 2234 3379 2238
rect 3407 2234 3411 2238
rect 3591 2234 3595 2238
rect 3615 2234 3619 2238
rect 1263 2150 1267 2154
rect 751 2066 755 2070
rect 783 2066 787 2070
rect 895 2066 899 2070
rect 935 2066 939 2070
rect 1327 2150 1331 2154
rect 1447 2150 1451 2154
rect 1567 2150 1571 2154
rect 1631 2150 1635 2154
rect 1815 2150 1819 2154
rect 1823 2150 1827 2154
rect 1047 2066 1051 2070
rect 1095 2066 1099 2070
rect 1215 2066 1219 2070
rect 1263 2066 1267 2070
rect 1399 2066 1403 2070
rect 1447 2066 1451 2070
rect 1583 2066 1587 2070
rect 495 1982 499 1986
rect 511 1982 515 1986
rect 615 1982 619 1986
rect 623 1982 627 1986
rect 743 1982 747 1986
rect 751 1982 755 1986
rect 871 1982 875 1986
rect 895 1982 899 1986
rect 1007 1982 1011 1986
rect 1047 1982 1051 1986
rect 1143 1982 1147 1986
rect 1215 1982 1219 1986
rect 1631 2066 1635 2070
rect 1775 2066 1779 2070
rect 2007 2150 2011 2154
rect 2047 2146 2051 2150
rect 2111 2146 2115 2150
rect 2255 2146 2259 2150
rect 2287 2146 2291 2150
rect 2407 2146 2411 2150
rect 2431 2146 2435 2150
rect 2559 2146 2563 2150
rect 2583 2146 2587 2150
rect 3839 2394 3843 2398
rect 3839 2318 3843 2322
rect 3943 2566 3947 2570
rect 3943 2486 3947 2490
rect 3943 2394 3947 2398
rect 3943 2318 3947 2322
rect 3783 2234 3787 2238
rect 3839 2234 3843 2238
rect 2719 2146 2723 2150
rect 2735 2146 2739 2150
rect 2879 2146 2883 2150
rect 2887 2146 2891 2150
rect 3047 2146 3051 2150
rect 3207 2146 3211 2150
rect 3223 2146 3227 2150
rect 3367 2146 3371 2150
rect 3407 2146 3411 2150
rect 3527 2146 3531 2150
rect 1823 2066 1827 2070
rect 2007 2066 2011 2070
rect 2047 2062 2051 2066
rect 2287 2062 2291 2066
rect 2431 2062 2435 2066
rect 2503 2062 2507 2066
rect 2583 2062 2587 2066
rect 2671 2062 2675 2066
rect 2735 2062 2739 2066
rect 2839 2062 2843 2066
rect 2887 2062 2891 2066
rect 1279 1982 1283 1986
rect 1399 1982 1403 1986
rect 1415 1982 1419 1986
rect 111 1898 115 1902
rect 511 1898 515 1902
rect 551 1898 555 1902
rect 623 1898 627 1902
rect 663 1898 667 1902
rect 743 1898 747 1902
rect 783 1898 787 1902
rect 871 1898 875 1902
rect 911 1898 915 1902
rect 1007 1898 1011 1902
rect 1047 1898 1051 1902
rect 111 1822 115 1826
rect 503 1822 507 1826
rect 551 1822 555 1826
rect 1143 1898 1147 1902
rect 1175 1898 1179 1902
rect 1279 1898 1283 1902
rect 1311 1898 1315 1902
rect 615 1822 619 1826
rect 663 1822 667 1826
rect 735 1822 739 1826
rect 783 1822 787 1826
rect 863 1822 867 1826
rect 911 1822 915 1826
rect 999 1822 1003 1826
rect 1047 1822 1051 1826
rect 1151 1822 1155 1826
rect 1175 1822 1179 1826
rect 1559 1982 1563 1986
rect 1583 1982 1587 1986
rect 1703 1982 1707 1986
rect 1775 1982 1779 1986
rect 2007 1982 2011 1986
rect 2047 1982 2051 1986
rect 2495 1982 2499 1986
rect 2503 1982 2507 1986
rect 3591 2146 3595 2150
rect 3695 2146 3699 2150
rect 3783 2146 3787 2150
rect 3839 2146 3843 2150
rect 3007 2062 3011 2066
rect 3047 2062 3051 2066
rect 3167 2062 3171 2066
rect 3207 2062 3211 2066
rect 3311 2062 3315 2066
rect 3367 2062 3371 2066
rect 3455 2062 3459 2066
rect 3527 2062 3531 2066
rect 3591 2062 3595 2066
rect 3695 2062 3699 2066
rect 3727 2062 3731 2066
rect 3839 2062 3843 2066
rect 2591 1982 2595 1986
rect 2671 1982 2675 1986
rect 2695 1982 2699 1986
rect 2807 1982 2811 1986
rect 2839 1982 2843 1986
rect 2927 1982 2931 1986
rect 3007 1982 3011 1986
rect 3047 1982 3051 1986
rect 3167 1982 3171 1986
rect 3175 1982 3179 1986
rect 3295 1982 3299 1986
rect 3311 1982 3315 1986
rect 3415 1982 3419 1986
rect 3455 1982 3459 1986
rect 3543 1982 3547 1986
rect 3591 1982 3595 1986
rect 3671 1982 3675 1986
rect 1415 1898 1419 1902
rect 1447 1898 1451 1902
rect 1559 1898 1563 1902
rect 1583 1898 1587 1902
rect 1703 1898 1707 1902
rect 1719 1898 1723 1902
rect 2007 1898 2011 1902
rect 2047 1902 2051 1906
rect 2071 1902 2075 1906
rect 2247 1902 2251 1906
rect 2439 1902 2443 1906
rect 2495 1902 2499 1906
rect 2591 1902 2595 1906
rect 2623 1902 2627 1906
rect 2695 1902 2699 1906
rect 2791 1902 2795 1906
rect 2807 1902 2811 1906
rect 1311 1822 1315 1826
rect 1319 1822 1323 1826
rect 1447 1822 1451 1826
rect 1487 1822 1491 1826
rect 1583 1822 1587 1826
rect 1663 1822 1667 1826
rect 111 1746 115 1750
rect 343 1746 347 1750
rect 463 1746 467 1750
rect 503 1746 507 1750
rect 591 1746 595 1750
rect 615 1746 619 1750
rect 719 1746 723 1750
rect 735 1746 739 1750
rect 111 1666 115 1670
rect 159 1666 163 1670
rect 295 1666 299 1670
rect 343 1666 347 1670
rect 455 1666 459 1670
rect 463 1666 467 1670
rect 591 1666 595 1670
rect 623 1666 627 1670
rect 719 1666 723 1670
rect 847 1746 851 1750
rect 863 1746 867 1750
rect 983 1746 987 1750
rect 999 1746 1003 1750
rect 1127 1746 1131 1750
rect 1151 1746 1155 1750
rect 1279 1746 1283 1750
rect 1319 1746 1323 1750
rect 799 1666 803 1670
rect 847 1666 851 1670
rect 983 1666 987 1670
rect 111 1590 115 1594
rect 135 1590 139 1594
rect 159 1590 163 1594
rect 255 1590 259 1594
rect 295 1590 299 1594
rect 423 1590 427 1594
rect 455 1590 459 1594
rect 607 1590 611 1594
rect 623 1590 627 1594
rect 799 1590 803 1594
rect 111 1510 115 1514
rect 135 1510 139 1514
rect 983 1590 987 1594
rect 991 1590 995 1594
rect 1127 1666 1131 1670
rect 1439 1746 1443 1750
rect 1487 1746 1491 1750
rect 1719 1822 1723 1826
rect 1847 1822 1851 1826
rect 2007 1822 2011 1826
rect 2047 1826 2051 1830
rect 2071 1826 2075 1830
rect 2095 1826 2099 1830
rect 2231 1826 2235 1830
rect 2247 1826 2251 1830
rect 2367 1826 2371 1830
rect 2439 1826 2443 1830
rect 3727 1982 3731 1986
rect 3799 1982 3803 1986
rect 3839 1982 3843 1986
rect 3943 2234 3947 2238
rect 3943 2146 3947 2150
rect 3943 2062 3947 2066
rect 2927 1902 2931 1906
rect 2959 1902 2963 1906
rect 3047 1902 3051 1906
rect 3127 1902 3131 1906
rect 3175 1902 3179 1906
rect 3295 1902 3299 1906
rect 3303 1902 3307 1906
rect 3415 1902 3419 1906
rect 3487 1902 3491 1906
rect 3543 1902 3547 1906
rect 3671 1902 3675 1906
rect 3799 1902 3803 1906
rect 3839 1902 3843 1906
rect 2511 1826 2515 1830
rect 2623 1826 2627 1830
rect 2671 1826 2675 1830
rect 2791 1826 2795 1830
rect 2855 1826 2859 1830
rect 2959 1826 2963 1830
rect 3071 1826 3075 1830
rect 3127 1826 3131 1830
rect 3303 1826 3307 1830
rect 3487 1826 3491 1830
rect 3543 1826 3547 1830
rect 1599 1746 1603 1750
rect 1663 1746 1667 1750
rect 1847 1746 1851 1750
rect 2007 1746 2011 1750
rect 2047 1750 2051 1754
rect 2095 1750 2099 1754
rect 2183 1750 2187 1754
rect 2231 1750 2235 1754
rect 2287 1750 2291 1754
rect 2367 1750 2371 1754
rect 2391 1750 2395 1754
rect 2495 1750 2499 1754
rect 2511 1750 2515 1754
rect 2599 1750 2603 1754
rect 2671 1750 2675 1754
rect 1167 1666 1171 1670
rect 1279 1666 1283 1670
rect 1351 1666 1355 1670
rect 1439 1666 1443 1670
rect 1543 1666 1547 1670
rect 2047 1674 2051 1678
rect 2183 1674 2187 1678
rect 2231 1674 2235 1678
rect 1599 1666 1603 1670
rect 1735 1666 1739 1670
rect 2007 1666 2011 1670
rect 1167 1590 1171 1594
rect 1183 1590 1187 1594
rect 1351 1590 1355 1594
rect 1367 1590 1371 1594
rect 247 1510 251 1514
rect 255 1510 259 1514
rect 399 1510 403 1514
rect 423 1510 427 1514
rect 559 1510 563 1514
rect 607 1510 611 1514
rect 719 1510 723 1514
rect 799 1510 803 1514
rect 879 1510 883 1514
rect 991 1510 995 1514
rect 1039 1510 1043 1514
rect 111 1434 115 1438
rect 135 1434 139 1438
rect 247 1434 251 1438
rect 263 1434 267 1438
rect 399 1434 403 1438
rect 431 1434 435 1438
rect 559 1434 563 1438
rect 607 1434 611 1438
rect 719 1434 723 1438
rect 791 1434 795 1438
rect 879 1434 883 1438
rect 111 1354 115 1358
rect 135 1354 139 1358
rect 159 1354 163 1358
rect 263 1354 267 1358
rect 311 1354 315 1358
rect 431 1354 435 1358
rect 479 1354 483 1358
rect 1183 1510 1187 1514
rect 1543 1590 1547 1594
rect 1551 1590 1555 1594
rect 1735 1590 1739 1594
rect 2287 1674 2291 1678
rect 2367 1674 2371 1678
rect 2391 1674 2395 1678
rect 2495 1674 2499 1678
rect 2519 1674 2523 1678
rect 2599 1674 2603 1678
rect 2703 1750 2707 1754
rect 3671 1826 3675 1830
rect 3791 1826 3795 1830
rect 3839 1826 3843 1830
rect 3943 1982 3947 1986
rect 3943 1902 3947 1906
rect 2807 1750 2811 1754
rect 2855 1750 2859 1754
rect 2911 1750 2915 1754
rect 3015 1750 3019 1754
rect 3071 1750 3075 1754
rect 3127 1750 3131 1754
rect 3303 1750 3307 1754
rect 3543 1750 3547 1754
rect 3791 1750 3795 1754
rect 2679 1674 2683 1678
rect 2703 1674 2707 1678
rect 2807 1674 2811 1678
rect 2847 1674 2851 1678
rect 2911 1674 2915 1678
rect 3015 1674 3019 1678
rect 3023 1674 3027 1678
rect 3127 1674 3131 1678
rect 3191 1674 3195 1678
rect 1903 1590 1907 1594
rect 2007 1590 2011 1594
rect 2047 1590 2051 1594
rect 2071 1590 2075 1594
rect 2231 1590 2235 1594
rect 2271 1590 2275 1594
rect 2367 1590 2371 1594
rect 2495 1590 2499 1594
rect 2519 1590 2523 1594
rect 1319 1510 1323 1514
rect 1367 1510 1371 1514
rect 1447 1510 1451 1514
rect 1551 1510 1555 1514
rect 1567 1510 1571 1514
rect 1687 1510 1691 1514
rect 1735 1510 1739 1514
rect 2679 1590 2683 1594
rect 2711 1590 2715 1594
rect 2847 1590 2851 1594
rect 2911 1590 2915 1594
rect 3023 1590 3027 1594
rect 3095 1590 3099 1594
rect 3359 1674 3363 1678
rect 3527 1674 3531 1678
rect 3695 1674 3699 1678
rect 3191 1590 3195 1594
rect 3263 1590 3267 1594
rect 3359 1590 3363 1594
rect 1807 1510 1811 1514
rect 1903 1510 1907 1514
rect 2007 1510 2011 1514
rect 2047 1514 2051 1518
rect 2071 1514 2075 1518
rect 2271 1514 2275 1518
rect 975 1434 979 1438
rect 1039 1434 1043 1438
rect 1159 1434 1163 1438
rect 1183 1434 1187 1438
rect 1319 1434 1323 1438
rect 1351 1434 1355 1438
rect 1447 1434 1451 1438
rect 1543 1434 1547 1438
rect 1567 1434 1571 1438
rect 1687 1434 1691 1438
rect 1735 1434 1739 1438
rect 1807 1434 1811 1438
rect 1903 1434 1907 1438
rect 2007 1434 2011 1438
rect 2431 1514 2435 1518
rect 2495 1514 2499 1518
rect 2711 1514 2715 1518
rect 2791 1514 2795 1518
rect 2911 1514 2915 1518
rect 3095 1514 3099 1518
rect 3127 1514 3131 1518
rect 3423 1590 3427 1594
rect 3527 1590 3531 1594
rect 3567 1590 3571 1594
rect 3695 1590 3699 1594
rect 3711 1590 3715 1594
rect 3839 1674 3843 1678
rect 3839 1590 3843 1594
rect 3943 1826 3947 1830
rect 3943 1750 3947 1754
rect 3943 1674 3947 1678
rect 3943 1590 3947 1594
rect 3263 1514 3267 1518
rect 3423 1514 3427 1518
rect 3463 1514 3467 1518
rect 3567 1514 3571 1518
rect 3711 1514 3715 1518
rect 3799 1514 3803 1518
rect 3839 1514 3843 1518
rect 3943 1514 3947 1518
rect 607 1354 611 1358
rect 663 1354 667 1358
rect 791 1354 795 1358
rect 855 1354 859 1358
rect 975 1354 979 1358
rect 1047 1354 1051 1358
rect 111 1274 115 1278
rect 159 1274 163 1278
rect 311 1274 315 1278
rect 407 1274 411 1278
rect 479 1274 483 1278
rect 543 1274 547 1278
rect 447 1267 451 1268
rect 447 1264 451 1267
rect 1159 1354 1163 1358
rect 1247 1354 1251 1358
rect 1351 1354 1355 1358
rect 1447 1354 1451 1358
rect 1543 1354 1547 1358
rect 1655 1354 1659 1358
rect 1735 1354 1739 1358
rect 2047 1430 2051 1434
rect 2071 1430 2075 1434
rect 2271 1430 2275 1434
rect 2431 1430 2435 1434
rect 2495 1430 2499 1434
rect 2711 1430 2715 1434
rect 2791 1430 2795 1434
rect 2911 1430 2915 1434
rect 3095 1430 3099 1434
rect 3127 1430 3131 1434
rect 3271 1430 3275 1434
rect 3439 1430 3443 1434
rect 3463 1430 3467 1434
rect 3607 1430 3611 1434
rect 3783 1430 3787 1434
rect 3799 1430 3803 1434
rect 1863 1354 1867 1358
rect 1903 1354 1907 1358
rect 2007 1354 2011 1358
rect 2047 1354 2051 1358
rect 2071 1354 2075 1358
rect 2207 1354 2211 1358
rect 2271 1354 2275 1358
rect 2383 1354 2387 1358
rect 2495 1354 2499 1358
rect 2567 1354 2571 1358
rect 663 1274 667 1278
rect 695 1274 699 1278
rect 855 1274 859 1278
rect 1023 1274 1027 1278
rect 1047 1274 1051 1278
rect 1191 1274 1195 1278
rect 1247 1274 1251 1278
rect 1367 1274 1371 1278
rect 1447 1274 1451 1278
rect 111 1198 115 1202
rect 407 1198 411 1202
rect 423 1198 427 1202
rect 543 1198 547 1202
rect 591 1198 595 1202
rect 979 1264 983 1268
rect 2711 1354 2715 1358
rect 2751 1354 2755 1358
rect 2911 1354 2915 1358
rect 2935 1354 2939 1358
rect 3095 1354 3099 1358
rect 3111 1354 3115 1358
rect 3271 1354 3275 1358
rect 3279 1354 3283 1358
rect 3439 1354 3443 1358
rect 3447 1354 3451 1358
rect 3943 1430 3947 1434
rect 3607 1354 3611 1358
rect 3623 1354 3627 1358
rect 3783 1354 3787 1358
rect 1543 1274 1547 1278
rect 1655 1274 1659 1278
rect 1719 1274 1723 1278
rect 1863 1274 1867 1278
rect 1895 1274 1899 1278
rect 2007 1274 2011 1278
rect 2047 1278 2051 1282
rect 2071 1278 2075 1282
rect 2151 1278 2155 1282
rect 2207 1278 2211 1282
rect 2287 1278 2291 1282
rect 2383 1278 2387 1282
rect 2431 1278 2435 1282
rect 2567 1278 2571 1282
rect 2583 1278 2587 1282
rect 2743 1278 2747 1282
rect 2751 1278 2755 1282
rect 2903 1278 2907 1282
rect 2935 1278 2939 1282
rect 695 1198 699 1202
rect 759 1198 763 1202
rect 855 1198 859 1202
rect 927 1198 931 1202
rect 1023 1198 1027 1202
rect 1095 1198 1099 1202
rect 1191 1198 1195 1202
rect 1247 1198 1251 1202
rect 111 1118 115 1122
rect 375 1118 379 1122
rect 423 1118 427 1122
rect 111 1042 115 1046
rect 303 1042 307 1046
rect 375 1042 379 1046
rect 487 1118 491 1122
rect 591 1118 595 1122
rect 599 1118 603 1122
rect 711 1118 715 1122
rect 759 1118 763 1122
rect 831 1118 835 1122
rect 927 1118 931 1122
rect 967 1118 971 1122
rect 1095 1118 1099 1122
rect 1119 1118 1123 1122
rect 1367 1198 1371 1202
rect 1399 1198 1403 1202
rect 1543 1198 1547 1202
rect 1687 1198 1691 1202
rect 1719 1198 1723 1202
rect 3071 1278 3075 1282
rect 3111 1278 3115 1282
rect 3247 1278 3251 1282
rect 3279 1278 3283 1282
rect 3431 1278 3435 1282
rect 3447 1278 3451 1282
rect 3615 1278 3619 1282
rect 3623 1278 3627 1282
rect 3807 1278 3811 1282
rect 1839 1198 1843 1202
rect 1895 1198 1899 1202
rect 2007 1198 2011 1202
rect 2047 1202 2051 1206
rect 2151 1202 2155 1206
rect 2287 1202 2291 1206
rect 2311 1202 2315 1206
rect 1247 1118 1251 1122
rect 1279 1118 1283 1122
rect 1399 1118 1403 1122
rect 1447 1118 1451 1122
rect 1543 1118 1547 1122
rect 447 1042 451 1046
rect 487 1042 491 1046
rect 591 1042 595 1046
rect 599 1042 603 1046
rect 711 1042 715 1046
rect 727 1042 731 1046
rect 111 966 115 970
rect 255 966 259 970
rect 303 966 307 970
rect 447 966 451 970
rect 111 886 115 890
rect 255 886 259 890
rect 591 966 595 970
rect 631 966 635 970
rect 831 1042 835 1046
rect 855 1042 859 1046
rect 967 1042 971 1046
rect 975 1042 979 1046
rect 1087 1042 1091 1046
rect 1119 1042 1123 1046
rect 1199 1042 1203 1046
rect 1279 1042 1283 1046
rect 1311 1042 1315 1046
rect 1431 1042 1435 1046
rect 1447 1042 1451 1046
rect 2415 1202 2419 1206
rect 2431 1202 2435 1206
rect 2527 1202 2531 1206
rect 2583 1202 2587 1206
rect 2639 1202 2643 1206
rect 2743 1202 2747 1206
rect 2767 1202 2771 1206
rect 2903 1202 2907 1206
rect 2911 1202 2915 1206
rect 3071 1202 3075 1206
rect 3247 1202 3251 1206
rect 3431 1202 3435 1206
rect 3439 1202 3443 1206
rect 3615 1202 3619 1206
rect 3631 1202 3635 1206
rect 3943 1354 3947 1358
rect 3943 1278 3947 1282
rect 3807 1202 3811 1206
rect 3831 1202 3835 1206
rect 2475 1136 2479 1140
rect 1623 1118 1627 1122
rect 1687 1118 1691 1122
rect 1839 1118 1843 1122
rect 2007 1118 2011 1122
rect 2047 1122 2051 1126
rect 2311 1122 2315 1126
rect 2407 1122 2411 1126
rect 2415 1122 2419 1126
rect 2723 1136 2727 1140
rect 2503 1122 2507 1126
rect 2527 1122 2531 1126
rect 2599 1122 2603 1126
rect 2639 1122 2643 1126
rect 2695 1122 2699 1126
rect 2767 1122 2771 1126
rect 2807 1122 2811 1126
rect 2911 1122 2915 1126
rect 2943 1122 2947 1126
rect 3071 1122 3075 1126
rect 3095 1122 3099 1126
rect 3247 1122 3251 1126
rect 3263 1122 3267 1126
rect 3439 1122 3443 1126
rect 3447 1122 3451 1126
rect 3631 1122 3635 1126
rect 3639 1122 3643 1126
rect 1623 1042 1627 1046
rect 2007 1042 2011 1046
rect 2047 1042 2051 1046
rect 2407 1042 2411 1046
rect 2455 1042 2459 1046
rect 2503 1042 2507 1046
rect 2551 1042 2555 1046
rect 2599 1042 2603 1046
rect 2647 1042 2651 1046
rect 727 966 731 970
rect 807 966 811 970
rect 855 966 859 970
rect 975 966 979 970
rect 1087 966 1091 970
rect 1127 966 1131 970
rect 1199 966 1203 970
rect 1271 966 1275 970
rect 1311 966 1315 970
rect 1415 966 1419 970
rect 1431 966 1435 970
rect 1551 966 1555 970
rect 1695 966 1699 970
rect 2007 966 2011 970
rect 2695 1042 2699 1046
rect 2759 1042 2763 1046
rect 2807 1042 2811 1046
rect 2887 1042 2891 1046
rect 447 886 451 890
rect 631 886 635 890
rect 639 886 643 890
rect 807 886 811 890
rect 823 886 827 890
rect 975 886 979 890
rect 999 886 1003 890
rect 111 806 115 810
rect 159 806 163 810
rect 255 806 259 810
rect 311 806 315 810
rect 447 806 451 810
rect 471 806 475 810
rect 111 730 115 734
rect 135 730 139 734
rect 159 730 163 734
rect 263 730 267 734
rect 311 730 315 734
rect 1127 886 1131 890
rect 1167 886 1171 890
rect 1271 886 1275 890
rect 1327 886 1331 890
rect 1415 886 1419 890
rect 1479 886 1483 890
rect 1551 886 1555 890
rect 1631 886 1635 890
rect 1695 886 1699 890
rect 2047 962 2051 966
rect 2423 962 2427 966
rect 2455 962 2459 966
rect 2519 962 2523 966
rect 2551 962 2555 966
rect 2615 962 2619 966
rect 2647 962 2651 966
rect 2711 962 2715 966
rect 2759 962 2763 966
rect 2823 962 2827 966
rect 2943 1042 2947 1046
rect 3031 1042 3035 1046
rect 3095 1042 3099 1046
rect 3183 1042 3187 1046
rect 3263 1042 3267 1046
rect 3343 1042 3347 1046
rect 2887 962 2891 966
rect 2951 962 2955 966
rect 3447 1042 3451 1046
rect 3503 1042 3507 1046
rect 3943 1202 3947 1206
rect 3831 1122 3835 1126
rect 3839 1122 3843 1126
rect 3943 1122 3947 1126
rect 3639 1042 3643 1046
rect 3671 1042 3675 1046
rect 3839 1042 3843 1046
rect 3031 962 3035 966
rect 3103 962 3107 966
rect 3183 962 3187 966
rect 3271 962 3275 966
rect 3343 962 3347 966
rect 3455 962 3459 966
rect 3503 962 3507 966
rect 3647 962 3651 966
rect 3671 962 3675 966
rect 1783 886 1787 890
rect 2007 886 2011 890
rect 2047 886 2051 890
rect 2343 886 2347 890
rect 2423 886 2427 890
rect 2439 886 2443 890
rect 2519 886 2523 890
rect 2535 886 2539 890
rect 2615 886 2619 890
rect 2631 886 2635 890
rect 2711 886 2715 890
rect 2735 886 2739 890
rect 2823 886 2827 890
rect 2863 886 2867 890
rect 2951 886 2955 890
rect 3015 886 3019 890
rect 3103 886 3107 890
rect 3191 886 3195 890
rect 3271 886 3275 890
rect 3391 886 3395 890
rect 3455 886 3459 890
rect 3607 886 3611 890
rect 3647 886 3651 890
rect 623 806 627 810
rect 639 806 643 810
rect 775 806 779 810
rect 823 806 827 810
rect 935 806 939 810
rect 999 806 1003 810
rect 1095 806 1099 810
rect 1167 806 1171 810
rect 1255 806 1259 810
rect 1327 806 1331 810
rect 1415 806 1419 810
rect 1479 806 1483 810
rect 431 730 435 734
rect 471 730 475 734
rect 623 730 627 734
rect 775 730 779 734
rect 823 730 827 734
rect 111 654 115 658
rect 135 654 139 658
rect 247 654 251 658
rect 263 654 267 658
rect 383 654 387 658
rect 111 574 115 578
rect 135 574 139 578
rect 247 574 251 578
rect 935 730 939 734
rect 1583 806 1587 810
rect 1631 806 1635 810
rect 1751 806 1755 810
rect 1783 806 1787 810
rect 1903 806 1907 810
rect 2007 806 2011 810
rect 2047 810 2051 814
rect 2311 810 2315 814
rect 2343 810 2347 814
rect 2439 810 2443 814
rect 2495 810 2499 814
rect 2535 810 2539 814
rect 2631 810 2635 814
rect 2687 810 2691 814
rect 2735 810 2739 814
rect 2863 810 2867 814
rect 2879 810 2883 814
rect 3015 810 3019 814
rect 3079 810 3083 814
rect 3191 810 3195 814
rect 3287 810 3291 814
rect 3391 810 3395 814
rect 3503 810 3507 814
rect 3607 810 3611 814
rect 1015 730 1019 734
rect 1095 730 1099 734
rect 1207 730 1211 734
rect 1255 730 1259 734
rect 1391 730 1395 734
rect 1415 730 1419 734
rect 1567 730 1571 734
rect 1583 730 1587 734
rect 1743 730 1747 734
rect 1751 730 1755 734
rect 431 654 435 658
rect 527 654 531 658
rect 623 654 627 658
rect 687 654 691 658
rect 823 654 827 658
rect 871 654 875 658
rect 1015 654 1019 658
rect 1079 654 1083 658
rect 1207 654 1211 658
rect 1303 654 1307 658
rect 1391 654 1395 658
rect 1543 654 1547 658
rect 1567 654 1571 658
rect 295 574 299 578
rect 383 574 387 578
rect 479 574 483 578
rect 527 574 531 578
rect 663 574 667 578
rect 687 574 691 578
rect 847 574 851 578
rect 871 574 875 578
rect 1903 730 1907 734
rect 3839 962 3843 966
rect 3943 1042 3947 1046
rect 3943 962 3947 966
rect 3823 886 3827 890
rect 3839 886 3843 890
rect 3719 810 3723 814
rect 3823 810 3827 814
rect 2007 730 2011 734
rect 2047 730 2051 734
rect 2071 730 2075 734
rect 2255 730 2259 734
rect 2311 730 2315 734
rect 2455 730 2459 734
rect 2495 730 2499 734
rect 2655 730 2659 734
rect 2687 730 2691 734
rect 2855 730 2859 734
rect 2879 730 2883 734
rect 3047 730 3051 734
rect 3079 730 3083 734
rect 3239 730 3243 734
rect 3287 730 3291 734
rect 3439 730 3443 734
rect 1743 654 1747 658
rect 1783 654 1787 658
rect 1903 654 1907 658
rect 2007 654 2011 658
rect 2047 654 2051 658
rect 2071 654 2075 658
rect 2231 654 2235 658
rect 2255 654 2259 658
rect 2431 654 2435 658
rect 2455 654 2459 658
rect 1031 574 1035 578
rect 1079 574 1083 578
rect 1215 574 1219 578
rect 1303 574 1307 578
rect 1399 574 1403 578
rect 1543 574 1547 578
rect 1591 574 1595 578
rect 1783 574 1787 578
rect 111 498 115 502
rect 135 498 139 502
rect 287 498 291 502
rect 295 498 299 502
rect 455 498 459 502
rect 479 498 483 502
rect 615 498 619 502
rect 663 498 667 502
rect 767 498 771 502
rect 847 498 851 502
rect 903 498 907 502
rect 111 422 115 426
rect 135 422 139 426
rect 287 422 291 426
rect 447 422 451 426
rect 455 422 459 426
rect 599 422 603 426
rect 615 422 619 426
rect 751 422 755 426
rect 767 422 771 426
rect 111 342 115 346
rect 135 342 139 346
rect 159 342 163 346
rect 287 342 291 346
rect 351 342 355 346
rect 447 342 451 346
rect 903 422 907 426
rect 1031 498 1035 502
rect 1159 498 1163 502
rect 1215 498 1219 502
rect 1287 498 1291 502
rect 1399 498 1403 502
rect 1415 498 1419 502
rect 2007 574 2011 578
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2631 654 2635 658
rect 2655 654 2659 658
rect 3503 730 3507 734
rect 3639 730 3643 734
rect 3719 730 3723 734
rect 2831 654 2835 658
rect 2855 654 2859 658
rect 3023 654 3027 658
rect 3047 654 3051 658
rect 3207 654 3211 658
rect 3239 654 3243 658
rect 3375 654 3379 658
rect 3439 654 3443 658
rect 3535 654 3539 658
rect 3639 654 3643 658
rect 3695 654 3699 658
rect 3839 730 3843 734
rect 3943 886 3947 890
rect 3943 810 3947 814
rect 3943 730 3947 734
rect 3839 654 3843 658
rect 2215 574 2219 578
rect 2231 574 2235 578
rect 2399 574 2403 578
rect 2431 574 2435 578
rect 2583 574 2587 578
rect 1591 498 1595 502
rect 1783 498 1787 502
rect 2007 498 2011 502
rect 2047 494 2051 498
rect 2071 494 2075 498
rect 2631 574 2635 578
rect 2775 574 2779 578
rect 2831 574 2835 578
rect 2959 574 2963 578
rect 3023 574 3027 578
rect 3143 574 3147 578
rect 3207 574 3211 578
rect 3319 574 3323 578
rect 3375 574 3379 578
rect 3495 574 3499 578
rect 3535 574 3539 578
rect 2215 494 2219 498
rect 2223 494 2227 498
rect 2391 494 2395 498
rect 2399 494 2403 498
rect 2559 494 2563 498
rect 2583 494 2587 498
rect 2727 494 2731 498
rect 2775 494 2779 498
rect 1031 422 1035 426
rect 1079 422 1083 426
rect 1159 422 1163 426
rect 1271 422 1275 426
rect 1287 422 1291 426
rect 551 342 555 346
rect 599 342 603 346
rect 751 342 755 346
rect 759 342 763 346
rect 903 342 907 346
rect 959 342 963 346
rect 1079 342 1083 346
rect 1159 342 1163 346
rect 1415 422 1419 426
rect 1479 422 1483 426
rect 1703 422 1707 426
rect 1903 422 1907 426
rect 2007 422 2011 426
rect 1271 342 1275 346
rect 1343 342 1347 346
rect 1479 342 1483 346
rect 1527 342 1531 346
rect 1703 342 1707 346
rect 1711 342 1715 346
rect 1895 342 1899 346
rect 1903 342 1907 346
rect 2047 418 2051 422
rect 2071 418 2075 422
rect 2223 418 2227 422
rect 2895 494 2899 498
rect 2959 494 2963 498
rect 3063 494 3067 498
rect 3143 494 3147 498
rect 3223 494 3227 498
rect 3119 472 3123 476
rect 3679 574 3683 578
rect 3695 574 3699 578
rect 3319 494 3323 498
rect 3383 494 3387 498
rect 3495 494 3499 498
rect 3543 494 3547 498
rect 3679 494 3683 498
rect 3703 494 3707 498
rect 3319 472 3323 476
rect 3943 654 3947 658
rect 3839 574 3843 578
rect 3839 494 3843 498
rect 3943 574 3947 578
rect 3943 494 3947 498
rect 2391 418 2395 422
rect 2463 418 2467 422
rect 2559 418 2563 422
rect 2655 418 2659 422
rect 2727 418 2731 422
rect 2751 418 2755 422
rect 2847 418 2851 422
rect 2895 418 2899 422
rect 2943 418 2947 422
rect 3039 418 3043 422
rect 3063 418 3067 422
rect 3135 418 3139 422
rect 3223 418 3227 422
rect 3231 418 3235 422
rect 3383 418 3387 422
rect 3543 418 3547 422
rect 3703 418 3707 422
rect 3839 418 3843 422
rect 3943 418 3947 422
rect 2007 342 2011 346
rect 2047 342 2051 346
rect 2399 342 2403 346
rect 2463 342 2467 346
rect 2503 342 2507 346
rect 2559 342 2563 346
rect 2623 342 2627 346
rect 2655 342 2659 346
rect 2751 342 2755 346
rect 2759 342 2763 346
rect 2847 342 2851 346
rect 111 258 115 262
rect 159 258 163 262
rect 223 258 227 262
rect 351 258 355 262
rect 383 258 387 262
rect 543 258 547 262
rect 551 258 555 262
rect 703 258 707 262
rect 759 258 763 262
rect 863 258 867 262
rect 111 162 115 166
rect 135 162 139 166
rect 223 162 227 166
rect 231 162 235 166
rect 327 162 331 166
rect 383 162 387 166
rect 423 162 427 166
rect 527 162 531 166
rect 543 162 547 166
rect 959 258 963 262
rect 1031 258 1035 262
rect 1159 258 1163 262
rect 1199 258 1203 262
rect 1343 258 1347 262
rect 1367 258 1371 262
rect 1527 258 1531 262
rect 1543 258 1547 262
rect 1711 258 1715 262
rect 1727 258 1731 262
rect 647 162 651 166
rect 703 162 707 166
rect 775 162 779 166
rect 863 162 867 166
rect 903 162 907 166
rect 1031 162 1035 166
rect 2047 266 2051 270
rect 2191 266 2195 270
rect 2351 266 2355 270
rect 2399 266 2403 270
rect 1895 258 1899 262
rect 1903 258 1907 262
rect 2007 258 2011 262
rect 2911 342 2915 346
rect 2943 342 2947 346
rect 3039 342 3043 346
rect 3071 342 3075 346
rect 3135 342 3139 346
rect 3231 342 3235 346
rect 3247 342 3251 346
rect 3423 342 3427 346
rect 3607 342 3611 346
rect 3791 342 3795 346
rect 3943 342 3947 346
rect 2503 266 2507 270
rect 2519 266 2523 270
rect 2623 266 2627 270
rect 2687 266 2691 270
rect 2759 266 2763 270
rect 2855 266 2859 270
rect 2911 266 2915 270
rect 1151 162 1155 166
rect 1199 162 1203 166
rect 1271 162 1275 166
rect 1367 162 1371 166
rect 1383 162 1387 166
rect 1487 162 1491 166
rect 1543 162 1547 166
rect 1591 162 1595 166
rect 1703 162 1707 166
rect 1727 162 1731 166
rect 1807 162 1811 166
rect 1903 162 1907 166
rect 2007 162 2011 166
rect 2047 158 2051 162
rect 2071 158 2075 162
rect 2167 158 2171 162
rect 2191 158 2195 162
rect 2263 158 2267 162
rect 2351 158 2355 162
rect 2367 158 2371 162
rect 2487 158 2491 162
rect 2519 158 2523 162
rect 2615 158 2619 162
rect 2687 158 2691 162
rect 3031 266 3035 270
rect 3071 266 3075 270
rect 3215 266 3219 270
rect 3247 266 3251 270
rect 3407 266 3411 270
rect 3423 266 3427 270
rect 3607 266 3611 270
rect 3791 266 3795 270
rect 3807 266 3811 270
rect 2743 158 2747 162
rect 2855 158 2859 162
rect 2871 158 2875 162
rect 2991 158 2995 162
rect 3031 158 3035 162
rect 3111 158 3115 162
rect 3215 158 3219 162
rect 3223 158 3227 162
rect 3327 158 3331 162
rect 3407 158 3411 162
rect 3431 158 3435 162
rect 3535 158 3539 162
rect 3607 158 3611 162
rect 3639 158 3643 162
rect 3743 158 3747 162
rect 3943 266 3947 270
rect 3807 158 3811 162
rect 3839 158 3843 162
rect 3943 158 3947 162
rect 111 86 115 90
rect 135 86 139 90
rect 231 86 235 90
rect 327 86 331 90
rect 423 86 427 90
rect 527 86 531 90
rect 647 86 651 90
rect 775 86 779 90
rect 903 86 907 90
rect 1031 86 1035 90
rect 1151 86 1155 90
rect 1271 86 1275 90
rect 1383 86 1387 90
rect 1487 86 1491 90
rect 1591 86 1595 90
rect 1703 86 1707 90
rect 1807 86 1811 90
rect 1903 86 1907 90
rect 2007 86 2011 90
rect 2047 82 2051 86
rect 2071 82 2075 86
rect 2167 82 2171 86
rect 2263 82 2267 86
rect 2367 82 2371 86
rect 2487 82 2491 86
rect 2615 82 2619 86
rect 2743 82 2747 86
rect 2871 82 2875 86
rect 2991 82 2995 86
rect 3111 82 3115 86
rect 3223 82 3227 86
rect 3327 82 3331 86
rect 3431 82 3435 86
rect 3535 82 3539 86
rect 3639 82 3643 86
rect 3743 82 3747 86
rect 3839 82 3843 86
rect 3943 82 3947 86
<< m4 >>
rect 2030 4025 2031 4031
rect 2037 4030 3979 4031
rect 2037 4026 2047 4030
rect 2051 4026 2071 4030
rect 2075 4026 3943 4030
rect 3947 4026 3979 4030
rect 2037 4025 3979 4026
rect 3985 4025 3986 4031
rect 96 4005 97 4011
rect 103 4010 2031 4011
rect 103 4006 111 4010
rect 115 4006 151 4010
rect 155 4006 279 4010
rect 283 4006 431 4010
rect 435 4006 607 4010
rect 611 4006 791 4010
rect 795 4006 975 4010
rect 979 4006 1151 4010
rect 1155 4006 1311 4010
rect 1315 4006 1471 4010
rect 1475 4006 1623 4010
rect 1627 4006 1775 4010
rect 1779 4006 1903 4010
rect 1907 4006 2007 4010
rect 2011 4006 2031 4010
rect 103 4005 2031 4006
rect 2037 4005 2038 4011
rect 2018 3949 2019 3955
rect 2025 3954 3967 3955
rect 2025 3950 2047 3954
rect 2051 3950 2071 3954
rect 2075 3950 2079 3954
rect 2083 3950 2215 3954
rect 2219 3950 2359 3954
rect 2363 3950 2503 3954
rect 2507 3950 2647 3954
rect 2651 3950 2791 3954
rect 2795 3950 2927 3954
rect 2931 3950 3055 3954
rect 3059 3950 3175 3954
rect 3179 3950 3295 3954
rect 3299 3950 3415 3954
rect 3419 3950 3535 3954
rect 3539 3950 3943 3954
rect 3947 3950 3967 3954
rect 2025 3949 3967 3950
rect 3973 3949 3974 3955
rect 84 3929 85 3935
rect 91 3934 2019 3935
rect 91 3930 111 3934
rect 115 3930 151 3934
rect 155 3930 279 3934
rect 283 3930 303 3934
rect 307 3930 423 3934
rect 427 3930 431 3934
rect 435 3930 551 3934
rect 555 3930 607 3934
rect 611 3930 687 3934
rect 691 3930 791 3934
rect 795 3930 815 3934
rect 819 3930 943 3934
rect 947 3930 975 3934
rect 979 3930 1071 3934
rect 1075 3930 1151 3934
rect 1155 3930 1199 3934
rect 1203 3930 1311 3934
rect 1315 3930 1327 3934
rect 1331 3930 1463 3934
rect 1467 3930 1471 3934
rect 1475 3930 1623 3934
rect 1627 3930 1775 3934
rect 1779 3930 1903 3934
rect 1907 3930 2007 3934
rect 2011 3930 2019 3934
rect 91 3929 2019 3930
rect 2025 3929 2026 3935
rect 2030 3873 2031 3879
rect 2037 3878 3979 3879
rect 2037 3874 2047 3878
rect 2051 3874 2079 3878
rect 2083 3874 2215 3878
rect 2219 3874 2255 3878
rect 2259 3874 2359 3878
rect 2363 3874 2383 3878
rect 2387 3874 2503 3878
rect 2507 3874 2519 3878
rect 2523 3874 2647 3878
rect 2651 3874 2671 3878
rect 2675 3874 2791 3878
rect 2795 3874 2831 3878
rect 2835 3874 2927 3878
rect 2931 3874 2991 3878
rect 2995 3874 3055 3878
rect 3059 3874 3159 3878
rect 3163 3874 3175 3878
rect 3179 3874 3295 3878
rect 3299 3874 3327 3878
rect 3331 3874 3415 3878
rect 3419 3874 3495 3878
rect 3499 3874 3535 3878
rect 3539 3874 3663 3878
rect 3667 3874 3943 3878
rect 3947 3874 3979 3878
rect 2037 3873 3979 3874
rect 3985 3873 3986 3879
rect 96 3849 97 3855
rect 103 3854 2031 3855
rect 103 3850 111 3854
rect 115 3850 303 3854
rect 307 3850 415 3854
rect 419 3850 423 3854
rect 427 3850 551 3854
rect 555 3850 567 3854
rect 571 3850 687 3854
rect 691 3850 727 3854
rect 731 3850 815 3854
rect 819 3850 887 3854
rect 891 3850 943 3854
rect 947 3850 1039 3854
rect 1043 3850 1071 3854
rect 1075 3850 1191 3854
rect 1195 3850 1199 3854
rect 1203 3850 1327 3854
rect 1331 3850 1343 3854
rect 1347 3850 1463 3854
rect 1467 3850 1495 3854
rect 1499 3850 1647 3854
rect 1651 3850 2007 3854
rect 2011 3850 2031 3854
rect 103 3849 2031 3850
rect 2037 3849 2038 3855
rect 2018 3797 2019 3803
rect 2025 3802 3967 3803
rect 2025 3798 2047 3802
rect 2051 3798 2071 3802
rect 2075 3798 2199 3802
rect 2203 3798 2255 3802
rect 2259 3798 2375 3802
rect 2379 3798 2383 3802
rect 2387 3798 2519 3802
rect 2523 3798 2559 3802
rect 2563 3798 2671 3802
rect 2675 3798 2751 3802
rect 2755 3798 2831 3802
rect 2835 3798 2951 3802
rect 2955 3798 2991 3802
rect 2995 3798 3143 3802
rect 3147 3798 3159 3802
rect 3163 3798 3327 3802
rect 3331 3798 3335 3802
rect 3339 3798 3495 3802
rect 3499 3798 3535 3802
rect 3539 3798 3663 3802
rect 3667 3798 3735 3802
rect 3739 3798 3943 3802
rect 3947 3798 3967 3802
rect 2025 3797 3967 3798
rect 3973 3797 3974 3803
rect 84 3769 85 3775
rect 91 3774 2019 3775
rect 91 3770 111 3774
rect 115 3770 399 3774
rect 403 3770 415 3774
rect 419 3770 567 3774
rect 571 3770 727 3774
rect 731 3770 751 3774
rect 755 3770 887 3774
rect 891 3770 935 3774
rect 939 3770 1039 3774
rect 1043 3770 1127 3774
rect 1131 3770 1191 3774
rect 1195 3770 1311 3774
rect 1315 3770 1343 3774
rect 1347 3770 1495 3774
rect 1499 3770 1503 3774
rect 1507 3770 1647 3774
rect 1651 3770 1695 3774
rect 1699 3770 1887 3774
rect 1891 3770 2007 3774
rect 2011 3770 2019 3774
rect 91 3769 2019 3770
rect 2025 3769 2026 3775
rect 2030 3709 2031 3715
rect 2037 3714 3979 3715
rect 2037 3710 2047 3714
rect 2051 3710 2071 3714
rect 2075 3710 2199 3714
rect 2203 3710 2263 3714
rect 2267 3710 2375 3714
rect 2379 3710 2479 3714
rect 2483 3710 2559 3714
rect 2563 3710 2695 3714
rect 2699 3710 2751 3714
rect 2755 3710 2911 3714
rect 2915 3710 2951 3714
rect 2955 3710 3119 3714
rect 3123 3710 3143 3714
rect 3147 3710 3319 3714
rect 3323 3710 3335 3714
rect 3339 3710 3519 3714
rect 3523 3710 3535 3714
rect 3539 3710 3727 3714
rect 3731 3710 3735 3714
rect 3739 3710 3943 3714
rect 3947 3710 3979 3714
rect 2037 3709 3979 3710
rect 3985 3709 3986 3715
rect 96 3681 97 3687
rect 103 3686 2031 3687
rect 103 3682 111 3686
rect 115 3682 367 3686
rect 371 3682 399 3686
rect 403 3682 519 3686
rect 523 3682 567 3686
rect 571 3682 679 3686
rect 683 3682 751 3686
rect 755 3682 847 3686
rect 851 3682 935 3686
rect 939 3682 1015 3686
rect 1019 3682 1127 3686
rect 1131 3682 1175 3686
rect 1179 3682 1311 3686
rect 1315 3682 1327 3686
rect 1331 3682 1479 3686
rect 1483 3682 1503 3686
rect 1507 3682 1631 3686
rect 1635 3682 1695 3686
rect 1699 3682 1791 3686
rect 1795 3682 1887 3686
rect 1891 3682 2007 3686
rect 2011 3682 2031 3686
rect 103 3681 2031 3682
rect 2037 3681 2038 3687
rect 2018 3629 2019 3635
rect 2025 3634 3967 3635
rect 2025 3630 2047 3634
rect 2051 3630 2071 3634
rect 2075 3630 2111 3634
rect 2115 3630 2263 3634
rect 2267 3630 2271 3634
rect 2275 3630 2455 3634
rect 2459 3630 2479 3634
rect 2483 3630 2655 3634
rect 2659 3630 2695 3634
rect 2699 3630 2871 3634
rect 2875 3630 2911 3634
rect 2915 3630 3095 3634
rect 3099 3630 3119 3634
rect 3123 3630 3319 3634
rect 3323 3630 3327 3634
rect 3331 3630 3519 3634
rect 3523 3630 3567 3634
rect 3571 3630 3727 3634
rect 3731 3630 3943 3634
rect 3947 3630 3967 3634
rect 2025 3629 3967 3630
rect 3973 3629 3974 3635
rect 84 3597 85 3603
rect 91 3602 2019 3603
rect 91 3598 111 3602
rect 115 3598 271 3602
rect 275 3598 367 3602
rect 371 3598 415 3602
rect 419 3598 519 3602
rect 523 3598 575 3602
rect 579 3598 679 3602
rect 683 3598 735 3602
rect 739 3598 847 3602
rect 851 3598 895 3602
rect 899 3598 1015 3602
rect 1019 3598 1055 3602
rect 1059 3598 1175 3602
rect 1179 3598 1215 3602
rect 1219 3598 1327 3602
rect 1331 3598 1375 3602
rect 1379 3598 1479 3602
rect 1483 3598 1543 3602
rect 1547 3598 1631 3602
rect 1635 3598 1791 3602
rect 1795 3598 2007 3602
rect 2011 3598 2019 3602
rect 91 3597 2019 3598
rect 2025 3597 2026 3603
rect 2030 3537 2031 3543
rect 2037 3542 3979 3543
rect 2037 3538 2047 3542
rect 2051 3538 2111 3542
rect 2115 3538 2271 3542
rect 2275 3538 2287 3542
rect 2291 3538 2383 3542
rect 2387 3538 2455 3542
rect 2459 3538 2479 3542
rect 2483 3538 2575 3542
rect 2579 3538 2655 3542
rect 2659 3538 2671 3542
rect 2675 3538 2767 3542
rect 2771 3538 2871 3542
rect 2875 3538 2983 3542
rect 2987 3538 3095 3542
rect 3099 3538 3103 3542
rect 3107 3538 3223 3542
rect 3227 3538 3327 3542
rect 3331 3538 3351 3542
rect 3355 3538 3487 3542
rect 3491 3538 3567 3542
rect 3571 3538 3943 3542
rect 3947 3538 3979 3542
rect 2037 3537 3979 3538
rect 3985 3537 3986 3543
rect 96 3513 97 3519
rect 103 3518 2031 3519
rect 103 3514 111 3518
rect 115 3514 159 3518
rect 163 3514 271 3518
rect 275 3514 287 3518
rect 291 3514 415 3518
rect 419 3514 423 3518
rect 427 3514 559 3518
rect 563 3514 575 3518
rect 579 3514 695 3518
rect 699 3514 735 3518
rect 739 3514 831 3518
rect 835 3514 895 3518
rect 899 3514 967 3518
rect 971 3514 1055 3518
rect 1059 3514 1095 3518
rect 1099 3514 1215 3518
rect 1219 3514 1231 3518
rect 1235 3514 1367 3518
rect 1371 3514 1375 3518
rect 1379 3514 1543 3518
rect 1547 3514 2007 3518
rect 2011 3514 2031 3518
rect 103 3513 2031 3514
rect 2037 3513 2038 3519
rect 2354 3500 2360 3501
rect 2862 3500 2868 3501
rect 2354 3496 2355 3500
rect 2359 3496 2863 3500
rect 2867 3496 2868 3500
rect 2354 3495 2360 3496
rect 2862 3495 2868 3496
rect 2018 3461 2019 3467
rect 2025 3466 3967 3467
rect 2025 3462 2047 3466
rect 2051 3462 2287 3466
rect 2291 3462 2383 3466
rect 2387 3462 2479 3466
rect 2483 3462 2487 3466
rect 2491 3462 2575 3466
rect 2579 3462 2583 3466
rect 2587 3462 2671 3466
rect 2675 3462 2679 3466
rect 2683 3462 2767 3466
rect 2771 3462 2783 3466
rect 2787 3462 2871 3466
rect 2875 3462 2895 3466
rect 2899 3462 2983 3466
rect 2987 3462 3015 3466
rect 3019 3462 3103 3466
rect 3107 3462 3143 3466
rect 3147 3462 3223 3466
rect 3227 3462 3271 3466
rect 3275 3462 3351 3466
rect 3355 3462 3407 3466
rect 3411 3462 3487 3466
rect 3491 3462 3943 3466
rect 3947 3462 3967 3466
rect 2025 3461 3967 3462
rect 3973 3461 3974 3467
rect 84 3429 85 3435
rect 91 3434 2019 3435
rect 91 3430 111 3434
rect 115 3430 135 3434
rect 139 3430 159 3434
rect 163 3430 247 3434
rect 251 3430 287 3434
rect 291 3430 383 3434
rect 387 3430 423 3434
rect 427 3430 527 3434
rect 531 3430 559 3434
rect 563 3430 671 3434
rect 675 3430 695 3434
rect 699 3430 815 3434
rect 819 3430 831 3434
rect 835 3430 967 3434
rect 971 3430 1095 3434
rect 1099 3430 1119 3434
rect 1123 3430 1231 3434
rect 1235 3430 1271 3434
rect 1275 3430 1367 3434
rect 1371 3430 2007 3434
rect 2011 3430 2019 3434
rect 91 3429 2019 3430
rect 2025 3429 2026 3435
rect 2030 3377 2031 3383
rect 2037 3382 3979 3383
rect 2037 3378 2047 3382
rect 2051 3378 2351 3382
rect 2355 3378 2479 3382
rect 2483 3378 2487 3382
rect 2491 3378 2583 3382
rect 2587 3378 2615 3382
rect 2619 3378 2679 3382
rect 2683 3378 2751 3382
rect 2755 3378 2783 3382
rect 2787 3378 2887 3382
rect 2891 3378 2895 3382
rect 2899 3378 3015 3382
rect 3019 3378 3023 3382
rect 3027 3378 3143 3382
rect 3147 3378 3159 3382
rect 3163 3378 3271 3382
rect 3275 3378 3303 3382
rect 3307 3378 3407 3382
rect 3411 3378 3943 3382
rect 3947 3378 3979 3382
rect 2037 3377 3979 3378
rect 3985 3377 3986 3383
rect 96 3345 97 3351
rect 103 3350 2031 3351
rect 103 3346 111 3350
rect 115 3346 135 3350
rect 139 3346 247 3350
rect 251 3346 263 3350
rect 267 3346 383 3350
rect 387 3346 431 3350
rect 435 3346 527 3350
rect 531 3346 599 3350
rect 603 3346 671 3350
rect 675 3346 767 3350
rect 771 3346 815 3350
rect 819 3346 927 3350
rect 931 3346 967 3350
rect 971 3346 1087 3350
rect 1091 3346 1119 3350
rect 1123 3346 1239 3350
rect 1243 3346 1271 3350
rect 1275 3346 1391 3350
rect 1395 3346 1551 3350
rect 1555 3346 2007 3350
rect 2011 3346 2031 3350
rect 103 3345 2031 3346
rect 2037 3345 2038 3351
rect 2018 3297 2019 3303
rect 2025 3302 3967 3303
rect 2025 3298 2047 3302
rect 2051 3298 2127 3302
rect 2131 3298 2295 3302
rect 2299 3298 2351 3302
rect 2355 3298 2455 3302
rect 2459 3298 2479 3302
rect 2483 3298 2615 3302
rect 2619 3298 2751 3302
rect 2755 3298 2775 3302
rect 2779 3298 2887 3302
rect 2891 3298 2935 3302
rect 2939 3298 3023 3302
rect 3027 3298 3095 3302
rect 3099 3298 3159 3302
rect 3163 3298 3263 3302
rect 3267 3298 3303 3302
rect 3307 3298 3943 3302
rect 3947 3298 3967 3302
rect 2025 3297 3967 3298
rect 3973 3297 3974 3303
rect 84 3261 85 3267
rect 91 3266 2019 3267
rect 91 3262 111 3266
rect 115 3262 135 3266
rect 139 3262 143 3266
rect 147 3262 263 3266
rect 267 3262 295 3266
rect 299 3262 431 3266
rect 435 3262 455 3266
rect 459 3262 599 3266
rect 603 3262 623 3266
rect 627 3262 767 3266
rect 771 3262 791 3266
rect 795 3262 927 3266
rect 931 3262 959 3266
rect 963 3262 1087 3266
rect 1091 3262 1127 3266
rect 1131 3262 1239 3266
rect 1243 3262 1303 3266
rect 1307 3262 1391 3266
rect 1395 3262 1479 3266
rect 1483 3262 1551 3266
rect 1555 3262 2007 3266
rect 2011 3262 2019 3266
rect 91 3261 2019 3262
rect 2025 3261 2026 3267
rect 2030 3221 2031 3227
rect 2037 3226 3979 3227
rect 2037 3222 2047 3226
rect 2051 3222 2071 3226
rect 2075 3222 2127 3226
rect 2131 3222 2207 3226
rect 2211 3222 2295 3226
rect 2299 3222 2375 3226
rect 2379 3222 2455 3226
rect 2459 3222 2543 3226
rect 2547 3222 2615 3226
rect 2619 3222 2703 3226
rect 2707 3222 2775 3226
rect 2779 3222 2863 3226
rect 2867 3222 2935 3226
rect 2939 3222 3015 3226
rect 3019 3222 3095 3226
rect 3099 3222 3167 3226
rect 3171 3222 3263 3226
rect 3267 3222 3327 3226
rect 3331 3222 3943 3226
rect 3947 3222 3979 3226
rect 2037 3221 3979 3222
rect 3985 3221 3986 3227
rect 182 3204 188 3205
rect 738 3204 744 3205
rect 182 3200 183 3204
rect 187 3200 739 3204
rect 743 3200 744 3204
rect 182 3199 188 3200
rect 738 3199 744 3200
rect 96 3185 97 3191
rect 103 3190 2031 3191
rect 103 3186 111 3190
rect 115 3186 143 3190
rect 147 3186 295 3190
rect 299 3186 431 3190
rect 435 3186 455 3190
rect 459 3186 567 3190
rect 571 3186 623 3190
rect 627 3186 703 3190
rect 707 3186 791 3190
rect 795 3186 855 3190
rect 859 3186 959 3190
rect 963 3186 1031 3190
rect 1035 3186 1127 3190
rect 1131 3186 1231 3190
rect 1235 3186 1303 3190
rect 1307 3186 1455 3190
rect 1459 3186 1479 3190
rect 1483 3186 1687 3190
rect 1691 3186 1903 3190
rect 1907 3186 2007 3190
rect 2011 3186 2031 3190
rect 103 3185 2031 3186
rect 2037 3185 2038 3191
rect 2018 3141 2019 3147
rect 2025 3146 3967 3147
rect 2025 3142 2047 3146
rect 2051 3142 2071 3146
rect 2075 3142 2207 3146
rect 2211 3142 2343 3146
rect 2347 3142 2375 3146
rect 2379 3142 2543 3146
rect 2547 3142 2631 3146
rect 2635 3142 2703 3146
rect 2707 3142 2863 3146
rect 2867 3142 2903 3146
rect 2907 3142 3015 3146
rect 3019 3142 3167 3146
rect 3171 3142 3175 3146
rect 3179 3142 3327 3146
rect 3331 3142 3447 3146
rect 3451 3142 3943 3146
rect 3947 3142 3967 3146
rect 2025 3141 3967 3142
rect 3973 3141 3974 3147
rect 84 3109 85 3115
rect 91 3114 2019 3115
rect 91 3110 111 3114
rect 115 3110 295 3114
rect 299 3110 311 3114
rect 315 3110 407 3114
rect 411 3110 431 3114
rect 435 3110 503 3114
rect 507 3110 567 3114
rect 571 3110 599 3114
rect 603 3110 695 3114
rect 699 3110 703 3114
rect 707 3110 807 3114
rect 811 3110 855 3114
rect 859 3110 943 3114
rect 947 3110 1031 3114
rect 1035 3110 1087 3114
rect 1091 3110 1231 3114
rect 1235 3110 1247 3114
rect 1251 3110 1407 3114
rect 1411 3110 1455 3114
rect 1459 3110 1575 3114
rect 1579 3110 1687 3114
rect 1691 3110 1751 3114
rect 1755 3110 1903 3114
rect 1907 3110 2007 3114
rect 2011 3110 2019 3114
rect 91 3109 2019 3110
rect 2025 3109 2026 3115
rect 2030 3061 2031 3067
rect 2037 3066 3979 3067
rect 2037 3062 2047 3066
rect 2051 3062 2071 3066
rect 2075 3062 2343 3066
rect 2347 3062 2487 3066
rect 2491 3062 2615 3066
rect 2619 3062 2631 3066
rect 2635 3062 2743 3066
rect 2747 3062 2863 3066
rect 2867 3062 2903 3066
rect 2907 3062 2983 3066
rect 2987 3062 3103 3066
rect 3107 3062 3175 3066
rect 3179 3062 3215 3066
rect 3219 3062 3327 3066
rect 3331 3062 3431 3066
rect 3435 3062 3447 3066
rect 3451 3062 3535 3066
rect 3539 3062 3639 3066
rect 3643 3062 3743 3066
rect 3747 3062 3839 3066
rect 3843 3062 3943 3066
rect 3947 3062 3979 3066
rect 2037 3061 3979 3062
rect 3985 3061 3986 3067
rect 462 3052 468 3053
rect 778 3052 784 3053
rect 462 3048 463 3052
rect 467 3048 779 3052
rect 783 3048 784 3052
rect 462 3047 468 3048
rect 778 3047 784 3048
rect 96 3033 97 3039
rect 103 3038 2031 3039
rect 103 3034 111 3038
rect 115 3034 311 3038
rect 315 3034 407 3038
rect 411 3034 423 3038
rect 427 3034 503 3038
rect 507 3034 519 3038
rect 523 3034 599 3038
rect 603 3034 615 3038
rect 619 3034 695 3038
rect 699 3034 711 3038
rect 715 3034 807 3038
rect 811 3034 815 3038
rect 819 3034 935 3038
rect 939 3034 943 3038
rect 947 3034 1055 3038
rect 1059 3034 1087 3038
rect 1091 3034 1183 3038
rect 1187 3034 1247 3038
rect 1251 3034 1311 3038
rect 1315 3034 1407 3038
rect 1411 3034 1431 3038
rect 1435 3034 1551 3038
rect 1555 3034 1575 3038
rect 1579 3034 1671 3038
rect 1675 3034 1751 3038
rect 1755 3034 1799 3038
rect 1803 3034 1903 3038
rect 1907 3034 2007 3038
rect 2011 3034 2031 3038
rect 103 3033 2031 3034
rect 2037 3033 2038 3039
rect 2018 2981 2019 2987
rect 2025 2986 3967 2987
rect 2025 2982 2047 2986
rect 2051 2982 2407 2986
rect 2411 2982 2487 2986
rect 2491 2982 2575 2986
rect 2579 2982 2615 2986
rect 2619 2982 2743 2986
rect 2747 2982 2767 2986
rect 2771 2982 2863 2986
rect 2867 2982 2967 2986
rect 2971 2982 2983 2986
rect 2987 2982 3103 2986
rect 3107 2982 3183 2986
rect 3187 2982 3215 2986
rect 3219 2982 3327 2986
rect 3331 2982 3399 2986
rect 3403 2982 3431 2986
rect 3435 2982 3535 2986
rect 3539 2982 3623 2986
rect 3627 2982 3639 2986
rect 3643 2982 3743 2986
rect 3747 2982 3839 2986
rect 3843 2982 3943 2986
rect 3947 2982 3967 2986
rect 2025 2981 3967 2982
rect 3973 2981 3974 2987
rect 84 2933 85 2939
rect 91 2938 2019 2939
rect 91 2934 111 2938
rect 115 2934 423 2938
rect 427 2934 519 2938
rect 523 2934 615 2938
rect 619 2934 711 2938
rect 715 2934 815 2938
rect 819 2934 935 2938
rect 939 2934 1055 2938
rect 1059 2934 1183 2938
rect 1187 2934 1311 2938
rect 1315 2934 1431 2938
rect 1435 2934 1479 2938
rect 1483 2934 1551 2938
rect 1555 2934 1575 2938
rect 1579 2934 1671 2938
rect 1675 2934 1767 2938
rect 1771 2934 1799 2938
rect 1803 2934 1863 2938
rect 1867 2934 1903 2938
rect 1907 2934 2007 2938
rect 2011 2934 2019 2938
rect 91 2933 2019 2934
rect 2025 2933 2026 2939
rect 2030 2889 2031 2895
rect 2037 2894 3979 2895
rect 2037 2890 2047 2894
rect 2051 2890 2407 2894
rect 2411 2890 2551 2894
rect 2555 2890 2575 2894
rect 2579 2890 2671 2894
rect 2675 2890 2767 2894
rect 2771 2890 2799 2894
rect 2803 2890 2927 2894
rect 2931 2890 2967 2894
rect 2971 2890 3055 2894
rect 3059 2890 3183 2894
rect 3187 2890 3311 2894
rect 3315 2890 3399 2894
rect 3403 2890 3439 2894
rect 3443 2890 3575 2894
rect 3579 2890 3623 2894
rect 3627 2890 3839 2894
rect 3843 2890 3943 2894
rect 3947 2890 3979 2894
rect 2037 2889 3979 2890
rect 3985 2889 3986 2895
rect 96 2849 97 2855
rect 103 2854 2031 2855
rect 103 2850 111 2854
rect 115 2850 279 2854
rect 283 2850 447 2854
rect 451 2850 631 2854
rect 635 2850 815 2854
rect 819 2850 999 2854
rect 1003 2850 1183 2854
rect 1187 2850 1359 2854
rect 1363 2850 1479 2854
rect 1483 2850 1527 2854
rect 1531 2850 1575 2854
rect 1579 2850 1671 2854
rect 1675 2850 1695 2854
rect 1699 2850 1767 2854
rect 1771 2850 1863 2854
rect 1867 2850 2007 2854
rect 2011 2850 2031 2854
rect 103 2849 2031 2850
rect 2037 2849 2038 2855
rect 2018 2813 2019 2819
rect 2025 2818 3967 2819
rect 2025 2814 2047 2818
rect 2051 2814 2439 2818
rect 2443 2814 2551 2818
rect 2555 2814 2567 2818
rect 2571 2814 2671 2818
rect 2675 2814 2695 2818
rect 2699 2814 2799 2818
rect 2803 2814 2831 2818
rect 2835 2814 2927 2818
rect 2931 2814 2967 2818
rect 2971 2814 3055 2818
rect 3059 2814 3103 2818
rect 3107 2814 3183 2818
rect 3187 2814 3247 2818
rect 3251 2814 3311 2818
rect 3315 2814 3391 2818
rect 3395 2814 3439 2818
rect 3443 2814 3543 2818
rect 3547 2814 3575 2818
rect 3579 2814 3703 2818
rect 3707 2814 3839 2818
rect 3843 2814 3943 2818
rect 3947 2814 3967 2818
rect 2025 2813 3967 2814
rect 3973 2813 3974 2819
rect 84 2773 85 2779
rect 91 2778 2019 2779
rect 91 2774 111 2778
rect 115 2774 239 2778
rect 243 2774 279 2778
rect 283 2774 351 2778
rect 355 2774 447 2778
rect 451 2774 471 2778
rect 475 2774 607 2778
rect 611 2774 631 2778
rect 635 2774 743 2778
rect 747 2774 815 2778
rect 819 2774 879 2778
rect 883 2774 999 2778
rect 1003 2774 1015 2778
rect 1019 2774 1151 2778
rect 1155 2774 1183 2778
rect 1187 2774 1287 2778
rect 1291 2774 1359 2778
rect 1363 2774 1423 2778
rect 1427 2774 1527 2778
rect 1531 2774 1567 2778
rect 1571 2774 1695 2778
rect 1699 2774 1863 2778
rect 1867 2774 2007 2778
rect 2011 2774 2019 2778
rect 91 2773 2019 2774
rect 2025 2773 2026 2779
rect 2030 2729 2031 2735
rect 2037 2734 3979 2735
rect 2037 2730 2047 2734
rect 2051 2730 2335 2734
rect 2339 2730 2439 2734
rect 2443 2730 2495 2734
rect 2499 2730 2567 2734
rect 2571 2730 2663 2734
rect 2667 2730 2695 2734
rect 2699 2730 2831 2734
rect 2835 2730 2967 2734
rect 2971 2730 2999 2734
rect 3003 2730 3103 2734
rect 3107 2730 3167 2734
rect 3171 2730 3247 2734
rect 3251 2730 3335 2734
rect 3339 2730 3391 2734
rect 3395 2730 3511 2734
rect 3515 2730 3543 2734
rect 3547 2730 3687 2734
rect 3691 2730 3703 2734
rect 3707 2730 3839 2734
rect 3843 2730 3943 2734
rect 3947 2730 3979 2734
rect 2037 2729 3979 2730
rect 3985 2729 3986 2735
rect 96 2697 97 2703
rect 103 2702 2031 2703
rect 103 2698 111 2702
rect 115 2698 223 2702
rect 227 2698 239 2702
rect 243 2698 351 2702
rect 355 2698 367 2702
rect 371 2698 471 2702
rect 475 2698 503 2702
rect 507 2698 607 2702
rect 611 2698 639 2702
rect 643 2698 743 2702
rect 747 2698 767 2702
rect 771 2698 879 2702
rect 883 2698 887 2702
rect 891 2698 999 2702
rect 1003 2698 1015 2702
rect 1019 2698 1111 2702
rect 1115 2698 1151 2702
rect 1155 2698 1231 2702
rect 1235 2698 1287 2702
rect 1291 2698 1351 2702
rect 1355 2698 1423 2702
rect 1427 2698 1567 2702
rect 1571 2698 2007 2702
rect 2011 2698 2031 2702
rect 103 2697 2031 2698
rect 2037 2697 2038 2703
rect 2018 2649 2019 2655
rect 2025 2654 3967 2655
rect 2025 2650 2047 2654
rect 2051 2650 2127 2654
rect 2131 2650 2279 2654
rect 2283 2650 2335 2654
rect 2339 2650 2447 2654
rect 2451 2650 2495 2654
rect 2499 2650 2623 2654
rect 2627 2650 2663 2654
rect 2667 2650 2807 2654
rect 2811 2650 2831 2654
rect 2835 2650 2991 2654
rect 2995 2650 2999 2654
rect 3003 2650 3167 2654
rect 3171 2650 3175 2654
rect 3179 2650 3335 2654
rect 3339 2650 3351 2654
rect 3355 2650 3511 2654
rect 3515 2650 3519 2654
rect 3523 2650 3687 2654
rect 3691 2650 3839 2654
rect 3843 2650 3943 2654
rect 3947 2650 3967 2654
rect 2025 2649 3967 2650
rect 3973 2649 3974 2655
rect 84 2621 85 2627
rect 91 2626 2019 2627
rect 91 2622 111 2626
rect 115 2622 175 2626
rect 179 2622 223 2626
rect 227 2622 367 2626
rect 371 2622 503 2626
rect 507 2622 543 2626
rect 547 2622 639 2626
rect 643 2622 711 2626
rect 715 2622 767 2626
rect 771 2622 863 2626
rect 867 2622 887 2626
rect 891 2622 999 2626
rect 1003 2622 1007 2626
rect 1011 2622 1111 2626
rect 1115 2622 1143 2626
rect 1147 2622 1231 2626
rect 1235 2622 1279 2626
rect 1283 2622 1351 2626
rect 1355 2622 1423 2626
rect 1427 2622 2007 2626
rect 2011 2622 2019 2626
rect 91 2621 2019 2622
rect 2025 2621 2026 2627
rect 2166 2580 2172 2581
rect 2598 2580 2604 2581
rect 2166 2576 2167 2580
rect 2171 2576 2599 2580
rect 2603 2576 2604 2580
rect 2166 2575 2172 2576
rect 2598 2575 2604 2576
rect 2030 2565 2031 2571
rect 2037 2570 3979 2571
rect 2037 2566 2047 2570
rect 2051 2566 2071 2570
rect 2075 2566 2127 2570
rect 2131 2566 2183 2570
rect 2187 2566 2279 2570
rect 2283 2566 2319 2570
rect 2323 2566 2447 2570
rect 2451 2566 2471 2570
rect 2475 2566 2623 2570
rect 2627 2566 2639 2570
rect 2643 2566 2807 2570
rect 2811 2566 2823 2570
rect 2827 2566 2991 2570
rect 2995 2566 3031 2570
rect 3035 2566 3175 2570
rect 3179 2566 3263 2570
rect 3267 2566 3351 2570
rect 3355 2566 3503 2570
rect 3507 2566 3519 2570
rect 3523 2566 3687 2570
rect 3691 2566 3743 2570
rect 3747 2566 3839 2570
rect 3843 2566 3943 2570
rect 3947 2566 3979 2570
rect 2037 2565 3979 2566
rect 3985 2565 3986 2571
rect 96 2541 97 2547
rect 103 2546 2031 2547
rect 103 2542 111 2546
rect 115 2542 135 2546
rect 139 2542 175 2546
rect 179 2542 271 2546
rect 275 2542 367 2546
rect 371 2542 439 2546
rect 443 2542 543 2546
rect 547 2542 607 2546
rect 611 2542 711 2546
rect 715 2542 775 2546
rect 779 2542 863 2546
rect 867 2542 927 2546
rect 931 2542 1007 2546
rect 1011 2542 1079 2546
rect 1083 2542 1143 2546
rect 1147 2542 1223 2546
rect 1227 2542 1279 2546
rect 1283 2542 1359 2546
rect 1363 2542 1423 2546
rect 1427 2542 1495 2546
rect 1499 2542 1639 2546
rect 1643 2542 2007 2546
rect 2011 2542 2031 2546
rect 103 2541 2031 2542
rect 2037 2541 2038 2547
rect 2018 2485 2019 2491
rect 2025 2490 3967 2491
rect 2025 2486 2047 2490
rect 2051 2486 2071 2490
rect 2075 2486 2183 2490
rect 2187 2486 2215 2490
rect 2219 2486 2319 2490
rect 2323 2486 2383 2490
rect 2387 2486 2471 2490
rect 2475 2486 2559 2490
rect 2563 2486 2639 2490
rect 2643 2486 2751 2490
rect 2755 2486 2823 2490
rect 2827 2486 2951 2490
rect 2955 2486 3031 2490
rect 3035 2486 3167 2490
rect 3171 2486 3263 2490
rect 3267 2486 3391 2490
rect 3395 2486 3503 2490
rect 3507 2486 3623 2490
rect 3627 2486 3743 2490
rect 3747 2486 3839 2490
rect 3843 2486 3943 2490
rect 3947 2486 3967 2490
rect 2025 2485 3967 2486
rect 3973 2485 3974 2491
rect 84 2461 85 2467
rect 91 2466 2019 2467
rect 91 2462 111 2466
rect 115 2462 135 2466
rect 139 2462 271 2466
rect 275 2462 311 2466
rect 315 2462 439 2466
rect 443 2462 511 2466
rect 515 2462 607 2466
rect 611 2462 711 2466
rect 715 2462 775 2466
rect 779 2462 903 2466
rect 907 2462 927 2466
rect 931 2462 1079 2466
rect 1083 2462 1223 2466
rect 1227 2462 1239 2466
rect 1243 2462 1359 2466
rect 1363 2462 1391 2466
rect 1395 2462 1495 2466
rect 1499 2462 1527 2466
rect 1531 2462 1639 2466
rect 1643 2462 1663 2466
rect 1667 2462 1791 2466
rect 1795 2462 1903 2466
rect 1907 2462 2007 2466
rect 2011 2462 2019 2466
rect 91 2461 2019 2462
rect 2025 2461 2026 2467
rect 2030 2393 2031 2399
rect 2037 2398 3979 2399
rect 2037 2394 2047 2398
rect 2051 2394 2071 2398
rect 2075 2394 2215 2398
rect 2219 2394 2247 2398
rect 2251 2394 2383 2398
rect 2387 2394 2431 2398
rect 2435 2394 2559 2398
rect 2563 2394 2607 2398
rect 2611 2394 2751 2398
rect 2755 2394 2775 2398
rect 2779 2394 2935 2398
rect 2939 2394 2951 2398
rect 2955 2394 3103 2398
rect 3107 2394 3167 2398
rect 3171 2394 3391 2398
rect 3395 2394 3623 2398
rect 3627 2394 3839 2398
rect 3843 2394 3943 2398
rect 3947 2394 3979 2398
rect 2037 2393 3979 2394
rect 3985 2393 3986 2399
rect 2030 2391 2038 2393
rect 96 2385 97 2391
rect 103 2390 2031 2391
rect 103 2386 111 2390
rect 115 2386 135 2390
rect 139 2386 311 2390
rect 315 2386 327 2390
rect 331 2386 511 2390
rect 515 2386 551 2390
rect 555 2386 711 2390
rect 715 2386 767 2390
rect 771 2386 903 2390
rect 907 2386 975 2390
rect 979 2386 1079 2390
rect 1083 2386 1175 2390
rect 1179 2386 1239 2390
rect 1243 2386 1367 2390
rect 1371 2386 1391 2390
rect 1395 2386 1527 2390
rect 1531 2386 1551 2390
rect 1555 2386 1663 2390
rect 1667 2386 1735 2390
rect 1739 2386 1791 2390
rect 1795 2386 1903 2390
rect 1907 2386 2007 2390
rect 2011 2386 2031 2390
rect 103 2385 2031 2386
rect 2037 2385 2038 2391
rect 2018 2317 2019 2323
rect 2025 2322 3967 2323
rect 2025 2318 2047 2322
rect 2051 2318 2071 2322
rect 2075 2318 2175 2322
rect 2179 2318 2247 2322
rect 2251 2318 2311 2322
rect 2315 2318 2431 2322
rect 2435 2318 2447 2322
rect 2451 2318 2591 2322
rect 2595 2318 2607 2322
rect 2611 2318 2751 2322
rect 2755 2318 2775 2322
rect 2779 2318 2935 2322
rect 2939 2318 3103 2322
rect 3107 2318 3143 2322
rect 3147 2318 3375 2322
rect 3379 2318 3615 2322
rect 3619 2318 3839 2322
rect 3843 2318 3943 2322
rect 3947 2318 3967 2322
rect 2025 2317 3967 2318
rect 3973 2317 3974 2323
rect 84 2301 85 2307
rect 91 2306 2019 2307
rect 91 2302 111 2306
rect 115 2302 135 2306
rect 139 2302 271 2306
rect 275 2302 327 2306
rect 331 2302 431 2306
rect 435 2302 551 2306
rect 555 2302 591 2306
rect 595 2302 751 2306
rect 755 2302 767 2306
rect 771 2302 919 2306
rect 923 2302 975 2306
rect 979 2302 1087 2306
rect 1091 2302 1175 2306
rect 1179 2302 1263 2306
rect 1267 2302 1367 2306
rect 1371 2302 1447 2306
rect 1451 2302 1551 2306
rect 1555 2302 1631 2306
rect 1635 2302 1735 2306
rect 1739 2302 1815 2306
rect 1819 2302 1903 2306
rect 1907 2302 2007 2306
rect 2011 2302 2019 2306
rect 91 2301 2019 2302
rect 2025 2301 2026 2307
rect 2030 2233 2031 2239
rect 2037 2238 3979 2239
rect 2037 2234 2047 2238
rect 2051 2234 2071 2238
rect 2075 2234 2111 2238
rect 2115 2234 2175 2238
rect 2179 2234 2255 2238
rect 2259 2234 2311 2238
rect 2315 2234 2407 2238
rect 2411 2234 2447 2238
rect 2451 2234 2559 2238
rect 2563 2234 2591 2238
rect 2595 2234 2719 2238
rect 2723 2234 2751 2238
rect 2755 2234 2879 2238
rect 2883 2234 2935 2238
rect 2939 2234 3047 2238
rect 3051 2234 3143 2238
rect 3147 2234 3223 2238
rect 3227 2234 3375 2238
rect 3379 2234 3407 2238
rect 3411 2234 3591 2238
rect 3595 2234 3615 2238
rect 3619 2234 3783 2238
rect 3787 2234 3839 2238
rect 3843 2234 3943 2238
rect 3947 2234 3979 2238
rect 2037 2233 3979 2234
rect 3985 2233 3986 2239
rect 2030 2231 2038 2233
rect 96 2225 97 2231
rect 103 2230 2031 2231
rect 103 2226 111 2230
rect 115 2226 135 2230
rect 139 2226 159 2230
rect 163 2226 271 2230
rect 275 2226 327 2230
rect 331 2226 431 2230
rect 435 2226 495 2230
rect 499 2226 591 2230
rect 595 2226 679 2230
rect 683 2226 751 2230
rect 755 2226 879 2230
rect 883 2226 919 2230
rect 923 2226 1087 2230
rect 1091 2226 1095 2230
rect 1099 2226 1263 2230
rect 1267 2226 1327 2230
rect 1331 2226 1447 2230
rect 1451 2226 1567 2230
rect 1571 2226 1631 2230
rect 1635 2226 1815 2230
rect 1819 2226 2007 2230
rect 2011 2226 2031 2230
rect 103 2225 2031 2226
rect 2037 2225 2038 2231
rect 84 2149 85 2155
rect 91 2154 2019 2155
rect 91 2150 111 2154
rect 115 2150 159 2154
rect 163 2150 223 2154
rect 227 2150 327 2154
rect 331 2150 359 2154
rect 363 2150 495 2154
rect 499 2150 639 2154
rect 643 2150 679 2154
rect 683 2150 783 2154
rect 787 2150 879 2154
rect 883 2150 935 2154
rect 939 2150 1095 2154
rect 1099 2150 1263 2154
rect 1267 2150 1327 2154
rect 1331 2150 1447 2154
rect 1451 2150 1567 2154
rect 1571 2150 1631 2154
rect 1635 2150 1815 2154
rect 1819 2150 1823 2154
rect 1827 2150 2007 2154
rect 2011 2150 2019 2154
rect 91 2149 2019 2150
rect 2025 2151 2026 2155
rect 2025 2150 3974 2151
rect 2025 2149 2047 2150
rect 2018 2146 2047 2149
rect 2051 2146 2111 2150
rect 2115 2146 2255 2150
rect 2259 2146 2287 2150
rect 2291 2146 2407 2150
rect 2411 2146 2431 2150
rect 2435 2146 2559 2150
rect 2563 2146 2583 2150
rect 2587 2146 2719 2150
rect 2723 2146 2735 2150
rect 2739 2146 2879 2150
rect 2883 2146 2887 2150
rect 2891 2146 3047 2150
rect 3051 2146 3207 2150
rect 3211 2146 3223 2150
rect 3227 2146 3367 2150
rect 3371 2146 3407 2150
rect 3411 2146 3527 2150
rect 3531 2146 3591 2150
rect 3595 2146 3695 2150
rect 3699 2146 3783 2150
rect 3787 2146 3839 2150
rect 3843 2146 3943 2150
rect 3947 2146 3974 2150
rect 2018 2145 3974 2146
rect 96 2065 97 2071
rect 103 2070 2031 2071
rect 103 2066 111 2070
rect 115 2066 223 2070
rect 227 2066 359 2070
rect 363 2066 375 2070
rect 379 2066 495 2070
rect 499 2066 615 2070
rect 619 2066 639 2070
rect 643 2066 751 2070
rect 755 2066 783 2070
rect 787 2066 895 2070
rect 899 2066 935 2070
rect 939 2066 1047 2070
rect 1051 2066 1095 2070
rect 1099 2066 1215 2070
rect 1219 2066 1263 2070
rect 1267 2066 1399 2070
rect 1403 2066 1447 2070
rect 1451 2066 1583 2070
rect 1587 2066 1631 2070
rect 1635 2066 1775 2070
rect 1779 2066 1823 2070
rect 1827 2066 2007 2070
rect 2011 2066 2031 2070
rect 103 2065 2031 2066
rect 2037 2067 2038 2071
rect 2037 2066 3986 2067
rect 2037 2065 2047 2066
rect 2030 2062 2047 2065
rect 2051 2062 2287 2066
rect 2291 2062 2431 2066
rect 2435 2062 2503 2066
rect 2507 2062 2583 2066
rect 2587 2062 2671 2066
rect 2675 2062 2735 2066
rect 2739 2062 2839 2066
rect 2843 2062 2887 2066
rect 2891 2062 3007 2066
rect 3011 2062 3047 2066
rect 3051 2062 3167 2066
rect 3171 2062 3207 2066
rect 3211 2062 3311 2066
rect 3315 2062 3367 2066
rect 3371 2062 3455 2066
rect 3459 2062 3527 2066
rect 3531 2062 3591 2066
rect 3595 2062 3695 2066
rect 3699 2062 3727 2066
rect 3731 2062 3839 2066
rect 3843 2062 3943 2066
rect 3947 2062 3986 2066
rect 2030 2061 3986 2062
rect 84 1981 85 1987
rect 91 1986 2019 1987
rect 91 1982 111 1986
rect 115 1982 375 1986
rect 379 1982 495 1986
rect 499 1982 511 1986
rect 515 1982 615 1986
rect 619 1982 623 1986
rect 627 1982 743 1986
rect 747 1982 751 1986
rect 755 1982 871 1986
rect 875 1982 895 1986
rect 899 1982 1007 1986
rect 1011 1982 1047 1986
rect 1051 1982 1143 1986
rect 1147 1982 1215 1986
rect 1219 1982 1279 1986
rect 1283 1982 1399 1986
rect 1403 1982 1415 1986
rect 1419 1982 1559 1986
rect 1563 1982 1583 1986
rect 1587 1982 1703 1986
rect 1707 1982 1775 1986
rect 1779 1982 2007 1986
rect 2011 1982 2019 1986
rect 91 1981 2019 1982
rect 2025 1986 3974 1987
rect 2025 1982 2047 1986
rect 2051 1982 2495 1986
rect 2499 1982 2503 1986
rect 2507 1982 2591 1986
rect 2595 1982 2671 1986
rect 2675 1982 2695 1986
rect 2699 1982 2807 1986
rect 2811 1982 2839 1986
rect 2843 1982 2927 1986
rect 2931 1982 3007 1986
rect 3011 1982 3047 1986
rect 3051 1982 3167 1986
rect 3171 1982 3175 1986
rect 3179 1982 3295 1986
rect 3299 1982 3311 1986
rect 3315 1982 3415 1986
rect 3419 1982 3455 1986
rect 3459 1982 3543 1986
rect 3547 1982 3591 1986
rect 3595 1982 3671 1986
rect 3675 1982 3727 1986
rect 3731 1982 3799 1986
rect 3803 1982 3839 1986
rect 3843 1982 3943 1986
rect 3947 1982 3974 1986
rect 2025 1981 3974 1982
rect 2030 1906 3986 1907
rect 2030 1903 2047 1906
rect 96 1897 97 1903
rect 103 1902 2031 1903
rect 103 1898 111 1902
rect 115 1898 511 1902
rect 515 1898 551 1902
rect 555 1898 623 1902
rect 627 1898 663 1902
rect 667 1898 743 1902
rect 747 1898 783 1902
rect 787 1898 871 1902
rect 875 1898 911 1902
rect 915 1898 1007 1902
rect 1011 1898 1047 1902
rect 1051 1898 1143 1902
rect 1147 1898 1175 1902
rect 1179 1898 1279 1902
rect 1283 1898 1311 1902
rect 1315 1898 1415 1902
rect 1419 1898 1447 1902
rect 1451 1898 1559 1902
rect 1563 1898 1583 1902
rect 1587 1898 1703 1902
rect 1707 1898 1719 1902
rect 1723 1898 2007 1902
rect 2011 1898 2031 1902
rect 103 1897 2031 1898
rect 2037 1902 2047 1903
rect 2051 1902 2071 1906
rect 2075 1902 2247 1906
rect 2251 1902 2439 1906
rect 2443 1902 2495 1906
rect 2499 1902 2591 1906
rect 2595 1902 2623 1906
rect 2627 1902 2695 1906
rect 2699 1902 2791 1906
rect 2795 1902 2807 1906
rect 2811 1902 2927 1906
rect 2931 1902 2959 1906
rect 2963 1902 3047 1906
rect 3051 1902 3127 1906
rect 3131 1902 3175 1906
rect 3179 1902 3295 1906
rect 3299 1902 3303 1906
rect 3307 1902 3415 1906
rect 3419 1902 3487 1906
rect 3491 1902 3543 1906
rect 3547 1902 3671 1906
rect 3675 1902 3799 1906
rect 3803 1902 3839 1906
rect 3843 1902 3943 1906
rect 3947 1902 3986 1906
rect 2037 1901 3986 1902
rect 2037 1897 2038 1901
rect 2018 1830 3974 1831
rect 2018 1827 2047 1830
rect 84 1821 85 1827
rect 91 1826 2019 1827
rect 91 1822 111 1826
rect 115 1822 503 1826
rect 507 1822 551 1826
rect 555 1822 615 1826
rect 619 1822 663 1826
rect 667 1822 735 1826
rect 739 1822 783 1826
rect 787 1822 863 1826
rect 867 1822 911 1826
rect 915 1822 999 1826
rect 1003 1822 1047 1826
rect 1051 1822 1151 1826
rect 1155 1822 1175 1826
rect 1179 1822 1311 1826
rect 1315 1822 1319 1826
rect 1323 1822 1447 1826
rect 1451 1822 1487 1826
rect 1491 1822 1583 1826
rect 1587 1822 1663 1826
rect 1667 1822 1719 1826
rect 1723 1822 1847 1826
rect 1851 1822 2007 1826
rect 2011 1822 2019 1826
rect 91 1821 2019 1822
rect 2025 1826 2047 1827
rect 2051 1826 2071 1830
rect 2075 1826 2095 1830
rect 2099 1826 2231 1830
rect 2235 1826 2247 1830
rect 2251 1826 2367 1830
rect 2371 1826 2439 1830
rect 2443 1826 2511 1830
rect 2515 1826 2623 1830
rect 2627 1826 2671 1830
rect 2675 1826 2791 1830
rect 2795 1826 2855 1830
rect 2859 1826 2959 1830
rect 2963 1826 3071 1830
rect 3075 1826 3127 1830
rect 3131 1826 3303 1830
rect 3307 1826 3487 1830
rect 3491 1826 3543 1830
rect 3547 1826 3671 1830
rect 3675 1826 3791 1830
rect 3795 1826 3839 1830
rect 3843 1826 3943 1830
rect 3947 1826 3974 1830
rect 2025 1825 3974 1826
rect 2025 1821 2026 1825
rect 2030 1754 3986 1755
rect 2030 1751 2047 1754
rect 96 1745 97 1751
rect 103 1750 2031 1751
rect 103 1746 111 1750
rect 115 1746 343 1750
rect 347 1746 463 1750
rect 467 1746 503 1750
rect 507 1746 591 1750
rect 595 1746 615 1750
rect 619 1746 719 1750
rect 723 1746 735 1750
rect 739 1746 847 1750
rect 851 1746 863 1750
rect 867 1746 983 1750
rect 987 1746 999 1750
rect 1003 1746 1127 1750
rect 1131 1746 1151 1750
rect 1155 1746 1279 1750
rect 1283 1746 1319 1750
rect 1323 1746 1439 1750
rect 1443 1746 1487 1750
rect 1491 1746 1599 1750
rect 1603 1746 1663 1750
rect 1667 1746 1847 1750
rect 1851 1746 2007 1750
rect 2011 1746 2031 1750
rect 103 1745 2031 1746
rect 2037 1750 2047 1751
rect 2051 1750 2095 1754
rect 2099 1750 2183 1754
rect 2187 1750 2231 1754
rect 2235 1750 2287 1754
rect 2291 1750 2367 1754
rect 2371 1750 2391 1754
rect 2395 1750 2495 1754
rect 2499 1750 2511 1754
rect 2515 1750 2599 1754
rect 2603 1750 2671 1754
rect 2675 1750 2703 1754
rect 2707 1750 2807 1754
rect 2811 1750 2855 1754
rect 2859 1750 2911 1754
rect 2915 1750 3015 1754
rect 3019 1750 3071 1754
rect 3075 1750 3127 1754
rect 3131 1750 3303 1754
rect 3307 1750 3543 1754
rect 3547 1750 3791 1754
rect 3795 1750 3943 1754
rect 3947 1750 3986 1754
rect 2037 1749 3986 1750
rect 2037 1745 2038 1749
rect 2018 1673 2019 1679
rect 2025 1678 3967 1679
rect 2025 1674 2047 1678
rect 2051 1674 2183 1678
rect 2187 1674 2231 1678
rect 2235 1674 2287 1678
rect 2291 1674 2367 1678
rect 2371 1674 2391 1678
rect 2395 1674 2495 1678
rect 2499 1674 2519 1678
rect 2523 1674 2599 1678
rect 2603 1674 2679 1678
rect 2683 1674 2703 1678
rect 2707 1674 2807 1678
rect 2811 1674 2847 1678
rect 2851 1674 2911 1678
rect 2915 1674 3015 1678
rect 3019 1674 3023 1678
rect 3027 1674 3127 1678
rect 3131 1674 3191 1678
rect 3195 1674 3359 1678
rect 3363 1674 3527 1678
rect 3531 1674 3695 1678
rect 3699 1674 3839 1678
rect 3843 1674 3943 1678
rect 3947 1674 3967 1678
rect 2025 1673 3967 1674
rect 3973 1673 3974 1679
rect 2018 1671 2026 1673
rect 84 1665 85 1671
rect 91 1670 2019 1671
rect 91 1666 111 1670
rect 115 1666 159 1670
rect 163 1666 295 1670
rect 299 1666 343 1670
rect 347 1666 455 1670
rect 459 1666 463 1670
rect 467 1666 591 1670
rect 595 1666 623 1670
rect 627 1666 719 1670
rect 723 1666 799 1670
rect 803 1666 847 1670
rect 851 1666 983 1670
rect 987 1666 1127 1670
rect 1131 1666 1167 1670
rect 1171 1666 1279 1670
rect 1283 1666 1351 1670
rect 1355 1666 1439 1670
rect 1443 1666 1543 1670
rect 1547 1666 1599 1670
rect 1603 1666 1735 1670
rect 1739 1666 2007 1670
rect 2011 1666 2019 1670
rect 91 1665 2019 1666
rect 2025 1665 2026 1671
rect 96 1589 97 1595
rect 103 1594 2031 1595
rect 103 1590 111 1594
rect 115 1590 135 1594
rect 139 1590 159 1594
rect 163 1590 255 1594
rect 259 1590 295 1594
rect 299 1590 423 1594
rect 427 1590 455 1594
rect 459 1590 607 1594
rect 611 1590 623 1594
rect 627 1590 799 1594
rect 803 1590 983 1594
rect 987 1590 991 1594
rect 995 1590 1167 1594
rect 1171 1590 1183 1594
rect 1187 1590 1351 1594
rect 1355 1590 1367 1594
rect 1371 1590 1543 1594
rect 1547 1590 1551 1594
rect 1555 1590 1735 1594
rect 1739 1590 1903 1594
rect 1907 1590 2007 1594
rect 2011 1590 2031 1594
rect 103 1589 2031 1590
rect 2037 1594 3986 1595
rect 2037 1590 2047 1594
rect 2051 1590 2071 1594
rect 2075 1590 2231 1594
rect 2235 1590 2271 1594
rect 2275 1590 2367 1594
rect 2371 1590 2495 1594
rect 2499 1590 2519 1594
rect 2523 1590 2679 1594
rect 2683 1590 2711 1594
rect 2715 1590 2847 1594
rect 2851 1590 2911 1594
rect 2915 1590 3023 1594
rect 3027 1590 3095 1594
rect 3099 1590 3191 1594
rect 3195 1590 3263 1594
rect 3267 1590 3359 1594
rect 3363 1590 3423 1594
rect 3427 1590 3527 1594
rect 3531 1590 3567 1594
rect 3571 1590 3695 1594
rect 3699 1590 3711 1594
rect 3715 1590 3839 1594
rect 3843 1590 3943 1594
rect 3947 1590 3986 1594
rect 2037 1589 3986 1590
rect 2018 1518 3974 1519
rect 2018 1515 2047 1518
rect 84 1509 85 1515
rect 91 1514 2019 1515
rect 91 1510 111 1514
rect 115 1510 135 1514
rect 139 1510 247 1514
rect 251 1510 255 1514
rect 259 1510 399 1514
rect 403 1510 423 1514
rect 427 1510 559 1514
rect 563 1510 607 1514
rect 611 1510 719 1514
rect 723 1510 799 1514
rect 803 1510 879 1514
rect 883 1510 991 1514
rect 995 1510 1039 1514
rect 1043 1510 1183 1514
rect 1187 1510 1319 1514
rect 1323 1510 1367 1514
rect 1371 1510 1447 1514
rect 1451 1510 1551 1514
rect 1555 1510 1567 1514
rect 1571 1510 1687 1514
rect 1691 1510 1735 1514
rect 1739 1510 1807 1514
rect 1811 1510 1903 1514
rect 1907 1510 2007 1514
rect 2011 1510 2019 1514
rect 91 1509 2019 1510
rect 2025 1514 2047 1515
rect 2051 1514 2071 1518
rect 2075 1514 2271 1518
rect 2275 1514 2431 1518
rect 2435 1514 2495 1518
rect 2499 1514 2711 1518
rect 2715 1514 2791 1518
rect 2795 1514 2911 1518
rect 2915 1514 3095 1518
rect 3099 1514 3127 1518
rect 3131 1514 3263 1518
rect 3267 1514 3423 1518
rect 3427 1514 3463 1518
rect 3467 1514 3567 1518
rect 3571 1514 3711 1518
rect 3715 1514 3799 1518
rect 3803 1514 3839 1518
rect 3843 1514 3943 1518
rect 3947 1514 3974 1518
rect 2025 1513 3974 1514
rect 2025 1509 2026 1513
rect 96 1433 97 1439
rect 103 1438 2031 1439
rect 103 1434 111 1438
rect 115 1434 135 1438
rect 139 1434 247 1438
rect 251 1434 263 1438
rect 267 1434 399 1438
rect 403 1434 431 1438
rect 435 1434 559 1438
rect 563 1434 607 1438
rect 611 1434 719 1438
rect 723 1434 791 1438
rect 795 1434 879 1438
rect 883 1434 975 1438
rect 979 1434 1039 1438
rect 1043 1434 1159 1438
rect 1163 1434 1183 1438
rect 1187 1434 1319 1438
rect 1323 1434 1351 1438
rect 1355 1434 1447 1438
rect 1451 1434 1543 1438
rect 1547 1434 1567 1438
rect 1571 1434 1687 1438
rect 1691 1434 1735 1438
rect 1739 1434 1807 1438
rect 1811 1434 1903 1438
rect 1907 1434 2007 1438
rect 2011 1434 2031 1438
rect 103 1433 2031 1434
rect 2037 1435 2038 1439
rect 2037 1434 3986 1435
rect 2037 1433 2047 1434
rect 2030 1430 2047 1433
rect 2051 1430 2071 1434
rect 2075 1430 2271 1434
rect 2275 1430 2431 1434
rect 2435 1430 2495 1434
rect 2499 1430 2711 1434
rect 2715 1430 2791 1434
rect 2795 1430 2911 1434
rect 2915 1430 3095 1434
rect 3099 1430 3127 1434
rect 3131 1430 3271 1434
rect 3275 1430 3439 1434
rect 3443 1430 3463 1434
rect 3467 1430 3607 1434
rect 3611 1430 3783 1434
rect 3787 1430 3799 1434
rect 3803 1430 3943 1434
rect 3947 1430 3986 1434
rect 2030 1429 3986 1430
rect 84 1353 85 1359
rect 91 1358 2019 1359
rect 91 1354 111 1358
rect 115 1354 135 1358
rect 139 1354 159 1358
rect 163 1354 263 1358
rect 267 1354 311 1358
rect 315 1354 431 1358
rect 435 1354 479 1358
rect 483 1354 607 1358
rect 611 1354 663 1358
rect 667 1354 791 1358
rect 795 1354 855 1358
rect 859 1354 975 1358
rect 979 1354 1047 1358
rect 1051 1354 1159 1358
rect 1163 1354 1247 1358
rect 1251 1354 1351 1358
rect 1355 1354 1447 1358
rect 1451 1354 1543 1358
rect 1547 1354 1655 1358
rect 1659 1354 1735 1358
rect 1739 1354 1863 1358
rect 1867 1354 1903 1358
rect 1907 1354 2007 1358
rect 2011 1354 2019 1358
rect 91 1353 2019 1354
rect 2025 1358 3974 1359
rect 2025 1354 2047 1358
rect 2051 1354 2071 1358
rect 2075 1354 2207 1358
rect 2211 1354 2271 1358
rect 2275 1354 2383 1358
rect 2387 1354 2495 1358
rect 2499 1354 2567 1358
rect 2571 1354 2711 1358
rect 2715 1354 2751 1358
rect 2755 1354 2911 1358
rect 2915 1354 2935 1358
rect 2939 1354 3095 1358
rect 3099 1354 3111 1358
rect 3115 1354 3271 1358
rect 3275 1354 3279 1358
rect 3283 1354 3439 1358
rect 3443 1354 3447 1358
rect 3451 1354 3607 1358
rect 3611 1354 3623 1358
rect 3627 1354 3783 1358
rect 3787 1354 3943 1358
rect 3947 1354 3974 1358
rect 2025 1353 3974 1354
rect 2030 1282 3986 1283
rect 2030 1279 2047 1282
rect 96 1273 97 1279
rect 103 1278 2031 1279
rect 103 1274 111 1278
rect 115 1274 159 1278
rect 163 1274 311 1278
rect 315 1274 407 1278
rect 411 1274 479 1278
rect 483 1274 543 1278
rect 547 1274 663 1278
rect 667 1274 695 1278
rect 699 1274 855 1278
rect 859 1274 1023 1278
rect 1027 1274 1047 1278
rect 1051 1274 1191 1278
rect 1195 1274 1247 1278
rect 1251 1274 1367 1278
rect 1371 1274 1447 1278
rect 1451 1274 1543 1278
rect 1547 1274 1655 1278
rect 1659 1274 1719 1278
rect 1723 1274 1863 1278
rect 1867 1274 1895 1278
rect 1899 1274 2007 1278
rect 2011 1274 2031 1278
rect 103 1273 2031 1274
rect 2037 1278 2047 1279
rect 2051 1278 2071 1282
rect 2075 1278 2151 1282
rect 2155 1278 2207 1282
rect 2211 1278 2287 1282
rect 2291 1278 2383 1282
rect 2387 1278 2431 1282
rect 2435 1278 2567 1282
rect 2571 1278 2583 1282
rect 2587 1278 2743 1282
rect 2747 1278 2751 1282
rect 2755 1278 2903 1282
rect 2907 1278 2935 1282
rect 2939 1278 3071 1282
rect 3075 1278 3111 1282
rect 3115 1278 3247 1282
rect 3251 1278 3279 1282
rect 3283 1278 3431 1282
rect 3435 1278 3447 1282
rect 3451 1278 3615 1282
rect 3619 1278 3623 1282
rect 3627 1278 3807 1282
rect 3811 1278 3943 1282
rect 3947 1278 3986 1282
rect 2037 1277 3986 1278
rect 2037 1273 2038 1277
rect 446 1268 452 1269
rect 978 1268 984 1269
rect 446 1264 447 1268
rect 451 1264 979 1268
rect 983 1264 984 1268
rect 446 1263 452 1264
rect 978 1263 984 1264
rect 2018 1206 3974 1207
rect 2018 1203 2047 1206
rect 84 1197 85 1203
rect 91 1202 2019 1203
rect 91 1198 111 1202
rect 115 1198 407 1202
rect 411 1198 423 1202
rect 427 1198 543 1202
rect 547 1198 591 1202
rect 595 1198 695 1202
rect 699 1198 759 1202
rect 763 1198 855 1202
rect 859 1198 927 1202
rect 931 1198 1023 1202
rect 1027 1198 1095 1202
rect 1099 1198 1191 1202
rect 1195 1198 1247 1202
rect 1251 1198 1367 1202
rect 1371 1198 1399 1202
rect 1403 1198 1543 1202
rect 1547 1198 1687 1202
rect 1691 1198 1719 1202
rect 1723 1198 1839 1202
rect 1843 1198 1895 1202
rect 1899 1198 2007 1202
rect 2011 1198 2019 1202
rect 91 1197 2019 1198
rect 2025 1202 2047 1203
rect 2051 1202 2151 1206
rect 2155 1202 2287 1206
rect 2291 1202 2311 1206
rect 2315 1202 2415 1206
rect 2419 1202 2431 1206
rect 2435 1202 2527 1206
rect 2531 1202 2583 1206
rect 2587 1202 2639 1206
rect 2643 1202 2743 1206
rect 2747 1202 2767 1206
rect 2771 1202 2903 1206
rect 2907 1202 2911 1206
rect 2915 1202 3071 1206
rect 3075 1202 3247 1206
rect 3251 1202 3431 1206
rect 3435 1202 3439 1206
rect 3443 1202 3615 1206
rect 3619 1202 3631 1206
rect 3635 1202 3807 1206
rect 3811 1202 3831 1206
rect 3835 1202 3943 1206
rect 3947 1202 3974 1206
rect 2025 1201 3974 1202
rect 2025 1197 2026 1201
rect 2474 1140 2480 1141
rect 2722 1140 2728 1141
rect 2474 1136 2475 1140
rect 2479 1136 2723 1140
rect 2727 1136 2728 1140
rect 2474 1135 2480 1136
rect 2722 1135 2728 1136
rect 2030 1126 3986 1127
rect 2030 1123 2047 1126
rect 96 1117 97 1123
rect 103 1122 2031 1123
rect 103 1118 111 1122
rect 115 1118 375 1122
rect 379 1118 423 1122
rect 427 1118 487 1122
rect 491 1118 591 1122
rect 595 1118 599 1122
rect 603 1118 711 1122
rect 715 1118 759 1122
rect 763 1118 831 1122
rect 835 1118 927 1122
rect 931 1118 967 1122
rect 971 1118 1095 1122
rect 1099 1118 1119 1122
rect 1123 1118 1247 1122
rect 1251 1118 1279 1122
rect 1283 1118 1399 1122
rect 1403 1118 1447 1122
rect 1451 1118 1543 1122
rect 1547 1118 1623 1122
rect 1627 1118 1687 1122
rect 1691 1118 1839 1122
rect 1843 1118 2007 1122
rect 2011 1118 2031 1122
rect 103 1117 2031 1118
rect 2037 1122 2047 1123
rect 2051 1122 2311 1126
rect 2315 1122 2407 1126
rect 2411 1122 2415 1126
rect 2419 1122 2503 1126
rect 2507 1122 2527 1126
rect 2531 1122 2599 1126
rect 2603 1122 2639 1126
rect 2643 1122 2695 1126
rect 2699 1122 2767 1126
rect 2771 1122 2807 1126
rect 2811 1122 2911 1126
rect 2915 1122 2943 1126
rect 2947 1122 3071 1126
rect 3075 1122 3095 1126
rect 3099 1122 3247 1126
rect 3251 1122 3263 1126
rect 3267 1122 3439 1126
rect 3443 1122 3447 1126
rect 3451 1122 3631 1126
rect 3635 1122 3639 1126
rect 3643 1122 3831 1126
rect 3835 1122 3839 1126
rect 3843 1122 3943 1126
rect 3947 1122 3986 1126
rect 2037 1121 3986 1122
rect 2037 1117 2038 1121
rect 84 1041 85 1047
rect 91 1046 2019 1047
rect 91 1042 111 1046
rect 115 1042 303 1046
rect 307 1042 375 1046
rect 379 1042 447 1046
rect 451 1042 487 1046
rect 491 1042 591 1046
rect 595 1042 599 1046
rect 603 1042 711 1046
rect 715 1042 727 1046
rect 731 1042 831 1046
rect 835 1042 855 1046
rect 859 1042 967 1046
rect 971 1042 975 1046
rect 979 1042 1087 1046
rect 1091 1042 1119 1046
rect 1123 1042 1199 1046
rect 1203 1042 1279 1046
rect 1283 1042 1311 1046
rect 1315 1042 1431 1046
rect 1435 1042 1447 1046
rect 1451 1042 1623 1046
rect 1627 1042 2007 1046
rect 2011 1042 2019 1046
rect 91 1041 2019 1042
rect 2025 1046 3974 1047
rect 2025 1042 2047 1046
rect 2051 1042 2407 1046
rect 2411 1042 2455 1046
rect 2459 1042 2503 1046
rect 2507 1042 2551 1046
rect 2555 1042 2599 1046
rect 2603 1042 2647 1046
rect 2651 1042 2695 1046
rect 2699 1042 2759 1046
rect 2763 1042 2807 1046
rect 2811 1042 2887 1046
rect 2891 1042 2943 1046
rect 2947 1042 3031 1046
rect 3035 1042 3095 1046
rect 3099 1042 3183 1046
rect 3187 1042 3263 1046
rect 3267 1042 3343 1046
rect 3347 1042 3447 1046
rect 3451 1042 3503 1046
rect 3507 1042 3639 1046
rect 3643 1042 3671 1046
rect 3675 1042 3839 1046
rect 3843 1042 3943 1046
rect 3947 1042 3974 1046
rect 2025 1041 3974 1042
rect 96 965 97 971
rect 103 970 2031 971
rect 103 966 111 970
rect 115 966 255 970
rect 259 966 303 970
rect 307 966 447 970
rect 451 966 591 970
rect 595 966 631 970
rect 635 966 727 970
rect 731 966 807 970
rect 811 966 855 970
rect 859 966 975 970
rect 979 966 1087 970
rect 1091 966 1127 970
rect 1131 966 1199 970
rect 1203 966 1271 970
rect 1275 966 1311 970
rect 1315 966 1415 970
rect 1419 966 1431 970
rect 1435 966 1551 970
rect 1555 966 1695 970
rect 1699 966 2007 970
rect 2011 966 2031 970
rect 103 965 2031 966
rect 2037 967 2038 971
rect 2037 966 3986 967
rect 2037 965 2047 966
rect 2030 962 2047 965
rect 2051 962 2423 966
rect 2427 962 2455 966
rect 2459 962 2519 966
rect 2523 962 2551 966
rect 2555 962 2615 966
rect 2619 962 2647 966
rect 2651 962 2711 966
rect 2715 962 2759 966
rect 2763 962 2823 966
rect 2827 962 2887 966
rect 2891 962 2951 966
rect 2955 962 3031 966
rect 3035 962 3103 966
rect 3107 962 3183 966
rect 3187 962 3271 966
rect 3275 962 3343 966
rect 3347 962 3455 966
rect 3459 962 3503 966
rect 3507 962 3647 966
rect 3651 962 3671 966
rect 3675 962 3839 966
rect 3843 962 3943 966
rect 3947 962 3986 966
rect 2030 961 3986 962
rect 84 885 85 891
rect 91 890 2019 891
rect 91 886 111 890
rect 115 886 255 890
rect 259 886 447 890
rect 451 886 631 890
rect 635 886 639 890
rect 643 886 807 890
rect 811 886 823 890
rect 827 886 975 890
rect 979 886 999 890
rect 1003 886 1127 890
rect 1131 886 1167 890
rect 1171 886 1271 890
rect 1275 886 1327 890
rect 1331 886 1415 890
rect 1419 886 1479 890
rect 1483 886 1551 890
rect 1555 886 1631 890
rect 1635 886 1695 890
rect 1699 886 1783 890
rect 1787 886 2007 890
rect 2011 886 2019 890
rect 91 885 2019 886
rect 2025 890 3974 891
rect 2025 886 2047 890
rect 2051 886 2343 890
rect 2347 886 2423 890
rect 2427 886 2439 890
rect 2443 886 2519 890
rect 2523 886 2535 890
rect 2539 886 2615 890
rect 2619 886 2631 890
rect 2635 886 2711 890
rect 2715 886 2735 890
rect 2739 886 2823 890
rect 2827 886 2863 890
rect 2867 886 2951 890
rect 2955 886 3015 890
rect 3019 886 3103 890
rect 3107 886 3191 890
rect 3195 886 3271 890
rect 3275 886 3391 890
rect 3395 886 3455 890
rect 3459 886 3607 890
rect 3611 886 3647 890
rect 3651 886 3823 890
rect 3827 886 3839 890
rect 3843 886 3943 890
rect 3947 886 3974 890
rect 2025 885 3974 886
rect 2030 814 3986 815
rect 2030 811 2047 814
rect 96 805 97 811
rect 103 810 2031 811
rect 103 806 111 810
rect 115 806 159 810
rect 163 806 255 810
rect 259 806 311 810
rect 315 806 447 810
rect 451 806 471 810
rect 475 806 623 810
rect 627 806 639 810
rect 643 806 775 810
rect 779 806 823 810
rect 827 806 935 810
rect 939 806 999 810
rect 1003 806 1095 810
rect 1099 806 1167 810
rect 1171 806 1255 810
rect 1259 806 1327 810
rect 1331 806 1415 810
rect 1419 806 1479 810
rect 1483 806 1583 810
rect 1587 806 1631 810
rect 1635 806 1751 810
rect 1755 806 1783 810
rect 1787 806 1903 810
rect 1907 806 2007 810
rect 2011 806 2031 810
rect 103 805 2031 806
rect 2037 810 2047 811
rect 2051 810 2311 814
rect 2315 810 2343 814
rect 2347 810 2439 814
rect 2443 810 2495 814
rect 2499 810 2535 814
rect 2539 810 2631 814
rect 2635 810 2687 814
rect 2691 810 2735 814
rect 2739 810 2863 814
rect 2867 810 2879 814
rect 2883 810 3015 814
rect 3019 810 3079 814
rect 3083 810 3191 814
rect 3195 810 3287 814
rect 3291 810 3391 814
rect 3395 810 3503 814
rect 3507 810 3607 814
rect 3611 810 3719 814
rect 3723 810 3823 814
rect 3827 810 3943 814
rect 3947 810 3986 814
rect 2037 809 3986 810
rect 2037 805 2038 809
rect 84 729 85 735
rect 91 734 2019 735
rect 91 730 111 734
rect 115 730 135 734
rect 139 730 159 734
rect 163 730 263 734
rect 267 730 311 734
rect 315 730 431 734
rect 435 730 471 734
rect 475 730 623 734
rect 627 730 775 734
rect 779 730 823 734
rect 827 730 935 734
rect 939 730 1015 734
rect 1019 730 1095 734
rect 1099 730 1207 734
rect 1211 730 1255 734
rect 1259 730 1391 734
rect 1395 730 1415 734
rect 1419 730 1567 734
rect 1571 730 1583 734
rect 1587 730 1743 734
rect 1747 730 1751 734
rect 1755 730 1903 734
rect 1907 730 2007 734
rect 2011 730 2019 734
rect 91 729 2019 730
rect 2025 734 3974 735
rect 2025 730 2047 734
rect 2051 730 2071 734
rect 2075 730 2255 734
rect 2259 730 2311 734
rect 2315 730 2455 734
rect 2459 730 2495 734
rect 2499 730 2655 734
rect 2659 730 2687 734
rect 2691 730 2855 734
rect 2859 730 2879 734
rect 2883 730 3047 734
rect 3051 730 3079 734
rect 3083 730 3239 734
rect 3243 730 3287 734
rect 3291 730 3439 734
rect 3443 730 3503 734
rect 3507 730 3639 734
rect 3643 730 3719 734
rect 3723 730 3839 734
rect 3843 730 3943 734
rect 3947 730 3974 734
rect 2025 729 3974 730
rect 96 653 97 659
rect 103 658 2031 659
rect 103 654 111 658
rect 115 654 135 658
rect 139 654 247 658
rect 251 654 263 658
rect 267 654 383 658
rect 387 654 431 658
rect 435 654 527 658
rect 531 654 623 658
rect 627 654 687 658
rect 691 654 823 658
rect 827 654 871 658
rect 875 654 1015 658
rect 1019 654 1079 658
rect 1083 654 1207 658
rect 1211 654 1303 658
rect 1307 654 1391 658
rect 1395 654 1543 658
rect 1547 654 1567 658
rect 1571 654 1743 658
rect 1747 654 1783 658
rect 1787 654 1903 658
rect 1907 654 2007 658
rect 2011 654 2031 658
rect 103 653 2031 654
rect 2037 658 3986 659
rect 2037 654 2047 658
rect 2051 654 2071 658
rect 2075 654 2231 658
rect 2235 654 2255 658
rect 2259 654 2431 658
rect 2435 654 2455 658
rect 2459 654 2631 658
rect 2635 654 2655 658
rect 2659 654 2831 658
rect 2835 654 2855 658
rect 2859 654 3023 658
rect 3027 654 3047 658
rect 3051 654 3207 658
rect 3211 654 3239 658
rect 3243 654 3375 658
rect 3379 654 3439 658
rect 3443 654 3535 658
rect 3539 654 3639 658
rect 3643 654 3695 658
rect 3699 654 3839 658
rect 3843 654 3943 658
rect 3947 654 3986 658
rect 2037 653 3986 654
rect 84 573 85 579
rect 91 578 2019 579
rect 91 574 111 578
rect 115 574 135 578
rect 139 574 247 578
rect 251 574 295 578
rect 299 574 383 578
rect 387 574 479 578
rect 483 574 527 578
rect 531 574 663 578
rect 667 574 687 578
rect 691 574 847 578
rect 851 574 871 578
rect 875 574 1031 578
rect 1035 574 1079 578
rect 1083 574 1215 578
rect 1219 574 1303 578
rect 1307 574 1399 578
rect 1403 574 1543 578
rect 1547 574 1591 578
rect 1595 574 1783 578
rect 1787 574 2007 578
rect 2011 574 2019 578
rect 91 573 2019 574
rect 2025 578 3974 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2215 578
rect 2219 574 2231 578
rect 2235 574 2399 578
rect 2403 574 2431 578
rect 2435 574 2583 578
rect 2587 574 2631 578
rect 2635 574 2775 578
rect 2779 574 2831 578
rect 2835 574 2959 578
rect 2963 574 3023 578
rect 3027 574 3143 578
rect 3147 574 3207 578
rect 3211 574 3319 578
rect 3323 574 3375 578
rect 3379 574 3495 578
rect 3499 574 3535 578
rect 3539 574 3679 578
rect 3683 574 3695 578
rect 3699 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3974 578
rect 2025 573 3974 574
rect 96 497 97 503
rect 103 502 2031 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 287 502
rect 291 498 295 502
rect 299 498 455 502
rect 459 498 479 502
rect 483 498 615 502
rect 619 498 663 502
rect 667 498 767 502
rect 771 498 847 502
rect 851 498 903 502
rect 907 498 1031 502
rect 1035 498 1159 502
rect 1163 498 1215 502
rect 1219 498 1287 502
rect 1291 498 1399 502
rect 1403 498 1415 502
rect 1419 498 1591 502
rect 1595 498 1783 502
rect 1787 498 2007 502
rect 2011 498 2031 502
rect 103 497 2031 498
rect 2037 499 2038 503
rect 2037 498 3986 499
rect 2037 497 2047 498
rect 2030 494 2047 497
rect 2051 494 2071 498
rect 2075 494 2215 498
rect 2219 494 2223 498
rect 2227 494 2391 498
rect 2395 494 2399 498
rect 2403 494 2559 498
rect 2563 494 2583 498
rect 2587 494 2727 498
rect 2731 494 2775 498
rect 2779 494 2895 498
rect 2899 494 2959 498
rect 2963 494 3063 498
rect 3067 494 3143 498
rect 3147 494 3223 498
rect 3227 494 3319 498
rect 3323 494 3383 498
rect 3387 494 3495 498
rect 3499 494 3543 498
rect 3547 494 3679 498
rect 3683 494 3703 498
rect 3707 494 3839 498
rect 3843 494 3943 498
rect 3947 494 3986 498
rect 2030 493 3986 494
rect 3118 476 3124 477
rect 3318 476 3324 477
rect 3118 472 3119 476
rect 3123 472 3319 476
rect 3323 472 3324 476
rect 3118 471 3124 472
rect 3318 471 3324 472
rect 84 421 85 427
rect 91 426 2019 427
rect 91 422 111 426
rect 115 422 135 426
rect 139 422 287 426
rect 291 422 447 426
rect 451 422 455 426
rect 459 422 599 426
rect 603 422 615 426
rect 619 422 751 426
rect 755 422 767 426
rect 771 422 903 426
rect 907 422 1031 426
rect 1035 422 1079 426
rect 1083 422 1159 426
rect 1163 422 1271 426
rect 1275 422 1287 426
rect 1291 422 1415 426
rect 1419 422 1479 426
rect 1483 422 1703 426
rect 1707 422 1903 426
rect 1907 422 2007 426
rect 2011 422 2019 426
rect 91 421 2019 422
rect 2025 423 2026 427
rect 2025 422 3974 423
rect 2025 421 2047 422
rect 2018 418 2047 421
rect 2051 418 2071 422
rect 2075 418 2223 422
rect 2227 418 2391 422
rect 2395 418 2463 422
rect 2467 418 2559 422
rect 2563 418 2655 422
rect 2659 418 2727 422
rect 2731 418 2751 422
rect 2755 418 2847 422
rect 2851 418 2895 422
rect 2899 418 2943 422
rect 2947 418 3039 422
rect 3043 418 3063 422
rect 3067 418 3135 422
rect 3139 418 3223 422
rect 3227 418 3231 422
rect 3235 418 3383 422
rect 3387 418 3543 422
rect 3547 418 3703 422
rect 3707 418 3839 422
rect 3843 418 3943 422
rect 3947 418 3974 422
rect 2018 417 3974 418
rect 96 341 97 347
rect 103 346 2031 347
rect 103 342 111 346
rect 115 342 135 346
rect 139 342 159 346
rect 163 342 287 346
rect 291 342 351 346
rect 355 342 447 346
rect 451 342 551 346
rect 555 342 599 346
rect 603 342 751 346
rect 755 342 759 346
rect 763 342 903 346
rect 907 342 959 346
rect 963 342 1079 346
rect 1083 342 1159 346
rect 1163 342 1271 346
rect 1275 342 1343 346
rect 1347 342 1479 346
rect 1483 342 1527 346
rect 1531 342 1703 346
rect 1707 342 1711 346
rect 1715 342 1895 346
rect 1899 342 1903 346
rect 1907 342 2007 346
rect 2011 342 2031 346
rect 103 341 2031 342
rect 2037 346 3986 347
rect 2037 342 2047 346
rect 2051 342 2399 346
rect 2403 342 2463 346
rect 2467 342 2503 346
rect 2507 342 2559 346
rect 2563 342 2623 346
rect 2627 342 2655 346
rect 2659 342 2751 346
rect 2755 342 2759 346
rect 2763 342 2847 346
rect 2851 342 2911 346
rect 2915 342 2943 346
rect 2947 342 3039 346
rect 3043 342 3071 346
rect 3075 342 3135 346
rect 3139 342 3231 346
rect 3235 342 3247 346
rect 3251 342 3423 346
rect 3427 342 3607 346
rect 3611 342 3791 346
rect 3795 342 3943 346
rect 3947 342 3986 346
rect 2037 341 3986 342
rect 2018 265 2019 271
rect 2025 270 3967 271
rect 2025 266 2047 270
rect 2051 266 2191 270
rect 2195 266 2351 270
rect 2355 266 2399 270
rect 2403 266 2503 270
rect 2507 266 2519 270
rect 2523 266 2623 270
rect 2627 266 2687 270
rect 2691 266 2759 270
rect 2763 266 2855 270
rect 2859 266 2911 270
rect 2915 266 3031 270
rect 3035 266 3071 270
rect 3075 266 3215 270
rect 3219 266 3247 270
rect 3251 266 3407 270
rect 3411 266 3423 270
rect 3427 266 3607 270
rect 3611 266 3791 270
rect 3795 266 3807 270
rect 3811 266 3943 270
rect 3947 266 3967 270
rect 2025 265 3967 266
rect 3973 265 3974 271
rect 2018 263 2026 265
rect 84 257 85 263
rect 91 262 2019 263
rect 91 258 111 262
rect 115 258 159 262
rect 163 258 223 262
rect 227 258 351 262
rect 355 258 383 262
rect 387 258 543 262
rect 547 258 551 262
rect 555 258 703 262
rect 707 258 759 262
rect 763 258 863 262
rect 867 258 959 262
rect 963 258 1031 262
rect 1035 258 1159 262
rect 1163 258 1199 262
rect 1203 258 1343 262
rect 1347 258 1367 262
rect 1371 258 1527 262
rect 1531 258 1543 262
rect 1547 258 1711 262
rect 1715 258 1727 262
rect 1731 258 1895 262
rect 1899 258 1903 262
rect 1907 258 2007 262
rect 2011 258 2019 262
rect 91 257 2019 258
rect 2025 257 2026 263
rect 96 161 97 167
rect 103 166 2031 167
rect 103 162 111 166
rect 115 162 135 166
rect 139 162 223 166
rect 227 162 231 166
rect 235 162 327 166
rect 331 162 383 166
rect 387 162 423 166
rect 427 162 527 166
rect 531 162 543 166
rect 547 162 647 166
rect 651 162 703 166
rect 707 162 775 166
rect 779 162 863 166
rect 867 162 903 166
rect 907 162 1031 166
rect 1035 162 1151 166
rect 1155 162 1199 166
rect 1203 162 1271 166
rect 1275 162 1367 166
rect 1371 162 1383 166
rect 1387 162 1487 166
rect 1491 162 1543 166
rect 1547 162 1591 166
rect 1595 162 1703 166
rect 1707 162 1727 166
rect 1731 162 1807 166
rect 1811 162 1903 166
rect 1907 162 2007 166
rect 2011 162 2031 166
rect 103 161 2031 162
rect 2037 163 2038 167
rect 2037 162 3986 163
rect 2037 161 2047 162
rect 2030 158 2047 161
rect 2051 158 2071 162
rect 2075 158 2167 162
rect 2171 158 2191 162
rect 2195 158 2263 162
rect 2267 158 2351 162
rect 2355 158 2367 162
rect 2371 158 2487 162
rect 2491 158 2519 162
rect 2523 158 2615 162
rect 2619 158 2687 162
rect 2691 158 2743 162
rect 2747 158 2855 162
rect 2859 158 2871 162
rect 2875 158 2991 162
rect 2995 158 3031 162
rect 3035 158 3111 162
rect 3115 158 3215 162
rect 3219 158 3223 162
rect 3227 158 3327 162
rect 3331 158 3407 162
rect 3411 158 3431 162
rect 3435 158 3535 162
rect 3539 158 3607 162
rect 3611 158 3639 162
rect 3643 158 3743 162
rect 3747 158 3807 162
rect 3811 158 3839 162
rect 3843 158 3943 162
rect 3947 158 3986 162
rect 2030 157 3986 158
rect 84 85 85 91
rect 91 90 2019 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 231 90
rect 235 86 327 90
rect 331 86 423 90
rect 427 86 527 90
rect 531 86 647 90
rect 651 86 775 90
rect 779 86 903 90
rect 907 86 1031 90
rect 1035 86 1151 90
rect 1155 86 1271 90
rect 1275 86 1383 90
rect 1387 86 1487 90
rect 1491 86 1591 90
rect 1595 86 1703 90
rect 1707 86 1807 90
rect 1811 86 1903 90
rect 1907 86 2007 90
rect 2011 86 2019 90
rect 91 85 2019 86
rect 2025 87 2026 91
rect 2025 86 3974 87
rect 2025 85 2047 86
rect 2018 82 2047 85
rect 2051 82 2071 86
rect 2075 82 2167 86
rect 2171 82 2263 86
rect 2267 82 2367 86
rect 2371 82 2487 86
rect 2491 82 2615 86
rect 2619 82 2743 86
rect 2747 82 2871 86
rect 2875 82 2991 86
rect 2995 82 3111 86
rect 3115 82 3223 86
rect 3227 82 3327 86
rect 3331 82 3431 86
rect 3435 82 3535 86
rect 3539 82 3639 86
rect 3643 82 3743 86
rect 3747 82 3839 86
rect 3843 82 3943 86
rect 3947 82 3974 86
rect 2018 81 3974 82
<< m5c >>
rect 2031 4025 2037 4031
rect 3979 4025 3985 4031
rect 97 4005 103 4011
rect 2031 4005 2037 4011
rect 2019 3949 2025 3955
rect 3967 3949 3973 3955
rect 85 3929 91 3935
rect 2019 3929 2025 3935
rect 2031 3873 2037 3879
rect 3979 3873 3985 3879
rect 97 3849 103 3855
rect 2031 3849 2037 3855
rect 2019 3797 2025 3803
rect 3967 3797 3973 3803
rect 85 3769 91 3775
rect 2019 3769 2025 3775
rect 2031 3709 2037 3715
rect 3979 3709 3985 3715
rect 97 3681 103 3687
rect 2031 3681 2037 3687
rect 2019 3629 2025 3635
rect 3967 3629 3973 3635
rect 85 3597 91 3603
rect 2019 3597 2025 3603
rect 2031 3537 2037 3543
rect 3979 3537 3985 3543
rect 97 3513 103 3519
rect 2031 3513 2037 3519
rect 2019 3461 2025 3467
rect 3967 3461 3973 3467
rect 85 3429 91 3435
rect 2019 3429 2025 3435
rect 2031 3377 2037 3383
rect 3979 3377 3985 3383
rect 97 3345 103 3351
rect 2031 3345 2037 3351
rect 2019 3297 2025 3303
rect 3967 3297 3973 3303
rect 85 3261 91 3267
rect 2019 3261 2025 3267
rect 2031 3221 2037 3227
rect 3979 3221 3985 3227
rect 97 3185 103 3191
rect 2031 3185 2037 3191
rect 2019 3141 2025 3147
rect 3967 3141 3973 3147
rect 85 3109 91 3115
rect 2019 3109 2025 3115
rect 2031 3061 2037 3067
rect 3979 3061 3985 3067
rect 97 3033 103 3039
rect 2031 3033 2037 3039
rect 2019 2981 2025 2987
rect 3967 2981 3973 2987
rect 85 2933 91 2939
rect 2019 2933 2025 2939
rect 2031 2889 2037 2895
rect 3979 2889 3985 2895
rect 97 2849 103 2855
rect 2031 2849 2037 2855
rect 2019 2813 2025 2819
rect 3967 2813 3973 2819
rect 85 2773 91 2779
rect 2019 2773 2025 2779
rect 2031 2729 2037 2735
rect 3979 2729 3985 2735
rect 97 2697 103 2703
rect 2031 2697 2037 2703
rect 2019 2649 2025 2655
rect 3967 2649 3973 2655
rect 85 2621 91 2627
rect 2019 2621 2025 2627
rect 2031 2565 2037 2571
rect 3979 2565 3985 2571
rect 97 2541 103 2547
rect 2031 2541 2037 2547
rect 2019 2485 2025 2491
rect 3967 2485 3973 2491
rect 85 2461 91 2467
rect 2019 2461 2025 2467
rect 2031 2393 2037 2399
rect 3979 2393 3985 2399
rect 97 2385 103 2391
rect 2031 2385 2037 2391
rect 2019 2317 2025 2323
rect 3967 2317 3973 2323
rect 85 2301 91 2307
rect 2019 2301 2025 2307
rect 2031 2233 2037 2239
rect 3979 2233 3985 2239
rect 97 2225 103 2231
rect 2031 2225 2037 2231
rect 85 2149 91 2155
rect 2019 2149 2025 2155
rect 97 2065 103 2071
rect 2031 2065 2037 2071
rect 85 1981 91 1987
rect 2019 1981 2025 1987
rect 97 1897 103 1903
rect 2031 1897 2037 1903
rect 85 1821 91 1827
rect 2019 1821 2025 1827
rect 97 1745 103 1751
rect 2031 1745 2037 1751
rect 2019 1673 2025 1679
rect 3967 1673 3973 1679
rect 85 1665 91 1671
rect 2019 1665 2025 1671
rect 97 1589 103 1595
rect 2031 1589 2037 1595
rect 85 1509 91 1515
rect 2019 1509 2025 1515
rect 97 1433 103 1439
rect 2031 1433 2037 1439
rect 85 1353 91 1359
rect 2019 1353 2025 1359
rect 97 1273 103 1279
rect 2031 1273 2037 1279
rect 85 1197 91 1203
rect 2019 1197 2025 1203
rect 97 1117 103 1123
rect 2031 1117 2037 1123
rect 85 1041 91 1047
rect 2019 1041 2025 1047
rect 97 965 103 971
rect 2031 965 2037 971
rect 85 885 91 891
rect 2019 885 2025 891
rect 97 805 103 811
rect 2031 805 2037 811
rect 85 729 91 735
rect 2019 729 2025 735
rect 97 653 103 659
rect 2031 653 2037 659
rect 85 573 91 579
rect 2019 573 2025 579
rect 97 497 103 503
rect 2031 497 2037 503
rect 85 421 91 427
rect 2019 421 2025 427
rect 97 341 103 347
rect 2031 341 2037 347
rect 2019 265 2025 271
rect 3967 265 3973 271
rect 85 257 91 263
rect 2019 257 2025 263
rect 97 161 103 167
rect 2031 161 2037 167
rect 85 85 91 91
rect 2019 85 2025 91
<< m5 >>
rect 84 3935 92 4032
rect 84 3929 85 3935
rect 91 3929 92 3935
rect 84 3775 92 3929
rect 84 3769 85 3775
rect 91 3769 92 3775
rect 84 3603 92 3769
rect 84 3597 85 3603
rect 91 3597 92 3603
rect 84 3435 92 3597
rect 84 3429 85 3435
rect 91 3429 92 3435
rect 84 3267 92 3429
rect 84 3261 85 3267
rect 91 3261 92 3267
rect 84 3115 92 3261
rect 84 3109 85 3115
rect 91 3109 92 3115
rect 84 2939 92 3109
rect 84 2933 85 2939
rect 91 2933 92 2939
rect 84 2779 92 2933
rect 84 2773 85 2779
rect 91 2773 92 2779
rect 84 2627 92 2773
rect 84 2621 85 2627
rect 91 2621 92 2627
rect 84 2467 92 2621
rect 84 2461 85 2467
rect 91 2461 92 2467
rect 84 2307 92 2461
rect 84 2301 85 2307
rect 91 2301 92 2307
rect 84 2155 92 2301
rect 84 2149 85 2155
rect 91 2149 92 2155
rect 84 1987 92 2149
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1827 92 1981
rect 84 1821 85 1827
rect 91 1821 92 1827
rect 84 1671 92 1821
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1515 92 1665
rect 84 1509 85 1515
rect 91 1509 92 1515
rect 84 1359 92 1509
rect 84 1353 85 1359
rect 91 1353 92 1359
rect 84 1203 92 1353
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1047 92 1197
rect 84 1041 85 1047
rect 91 1041 92 1047
rect 84 891 92 1041
rect 84 885 85 891
rect 91 885 92 891
rect 84 735 92 885
rect 84 729 85 735
rect 91 729 92 735
rect 84 579 92 729
rect 84 573 85 579
rect 91 573 92 579
rect 84 427 92 573
rect 84 421 85 427
rect 91 421 92 427
rect 84 263 92 421
rect 84 257 85 263
rect 91 257 92 263
rect 84 91 92 257
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 4011 104 4032
rect 96 4005 97 4011
rect 103 4005 104 4011
rect 96 3855 104 4005
rect 96 3849 97 3855
rect 103 3849 104 3855
rect 96 3687 104 3849
rect 96 3681 97 3687
rect 103 3681 104 3687
rect 96 3519 104 3681
rect 96 3513 97 3519
rect 103 3513 104 3519
rect 96 3351 104 3513
rect 96 3345 97 3351
rect 103 3345 104 3351
rect 96 3191 104 3345
rect 96 3185 97 3191
rect 103 3185 104 3191
rect 96 3039 104 3185
rect 96 3033 97 3039
rect 103 3033 104 3039
rect 96 2855 104 3033
rect 96 2849 97 2855
rect 103 2849 104 2855
rect 96 2703 104 2849
rect 96 2697 97 2703
rect 103 2697 104 2703
rect 96 2547 104 2697
rect 96 2541 97 2547
rect 103 2541 104 2547
rect 96 2391 104 2541
rect 96 2385 97 2391
rect 103 2385 104 2391
rect 96 2231 104 2385
rect 96 2225 97 2231
rect 103 2225 104 2231
rect 96 2071 104 2225
rect 96 2065 97 2071
rect 103 2065 104 2071
rect 96 1903 104 2065
rect 96 1897 97 1903
rect 103 1897 104 1903
rect 96 1751 104 1897
rect 96 1745 97 1751
rect 103 1745 104 1751
rect 96 1595 104 1745
rect 96 1589 97 1595
rect 103 1589 104 1595
rect 96 1439 104 1589
rect 96 1433 97 1439
rect 103 1433 104 1439
rect 96 1279 104 1433
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1123 104 1273
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 971 104 1117
rect 96 965 97 971
rect 103 965 104 971
rect 96 811 104 965
rect 96 805 97 811
rect 103 805 104 811
rect 96 659 104 805
rect 96 653 97 659
rect 103 653 104 659
rect 96 503 104 653
rect 96 497 97 503
rect 103 497 104 503
rect 96 347 104 497
rect 96 341 97 347
rect 103 341 104 347
rect 96 167 104 341
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 2018 3955 2026 4032
rect 2018 3949 2019 3955
rect 2025 3949 2026 3955
rect 2018 3935 2026 3949
rect 2018 3929 2019 3935
rect 2025 3929 2026 3935
rect 2018 3803 2026 3929
rect 2018 3797 2019 3803
rect 2025 3797 2026 3803
rect 2018 3775 2026 3797
rect 2018 3769 2019 3775
rect 2025 3769 2026 3775
rect 2018 3635 2026 3769
rect 2018 3629 2019 3635
rect 2025 3629 2026 3635
rect 2018 3603 2026 3629
rect 2018 3597 2019 3603
rect 2025 3597 2026 3603
rect 2018 3467 2026 3597
rect 2018 3461 2019 3467
rect 2025 3461 2026 3467
rect 2018 3435 2026 3461
rect 2018 3429 2019 3435
rect 2025 3429 2026 3435
rect 2018 3303 2026 3429
rect 2018 3297 2019 3303
rect 2025 3297 2026 3303
rect 2018 3267 2026 3297
rect 2018 3261 2019 3267
rect 2025 3261 2026 3267
rect 2018 3147 2026 3261
rect 2018 3141 2019 3147
rect 2025 3141 2026 3147
rect 2018 3115 2026 3141
rect 2018 3109 2019 3115
rect 2025 3109 2026 3115
rect 2018 2987 2026 3109
rect 2018 2981 2019 2987
rect 2025 2981 2026 2987
rect 2018 2939 2026 2981
rect 2018 2933 2019 2939
rect 2025 2933 2026 2939
rect 2018 2819 2026 2933
rect 2018 2813 2019 2819
rect 2025 2813 2026 2819
rect 2018 2779 2026 2813
rect 2018 2773 2019 2779
rect 2025 2773 2026 2779
rect 2018 2655 2026 2773
rect 2018 2649 2019 2655
rect 2025 2649 2026 2655
rect 2018 2627 2026 2649
rect 2018 2621 2019 2627
rect 2025 2621 2026 2627
rect 2018 2491 2026 2621
rect 2018 2485 2019 2491
rect 2025 2485 2026 2491
rect 2018 2467 2026 2485
rect 2018 2461 2019 2467
rect 2025 2461 2026 2467
rect 2018 2323 2026 2461
rect 2018 2317 2019 2323
rect 2025 2317 2026 2323
rect 2018 2307 2026 2317
rect 2018 2301 2019 2307
rect 2025 2301 2026 2307
rect 2018 2155 2026 2301
rect 2018 2149 2019 2155
rect 2025 2149 2026 2155
rect 2018 1987 2026 2149
rect 2018 1981 2019 1987
rect 2025 1981 2026 1987
rect 2018 1827 2026 1981
rect 2018 1821 2019 1827
rect 2025 1821 2026 1827
rect 2018 1679 2026 1821
rect 2018 1673 2019 1679
rect 2025 1673 2026 1679
rect 2018 1671 2026 1673
rect 2018 1665 2019 1671
rect 2025 1665 2026 1671
rect 2018 1515 2026 1665
rect 2018 1509 2019 1515
rect 2025 1509 2026 1515
rect 2018 1359 2026 1509
rect 2018 1353 2019 1359
rect 2025 1353 2026 1359
rect 2018 1203 2026 1353
rect 2018 1197 2019 1203
rect 2025 1197 2026 1203
rect 2018 1047 2026 1197
rect 2018 1041 2019 1047
rect 2025 1041 2026 1047
rect 2018 891 2026 1041
rect 2018 885 2019 891
rect 2025 885 2026 891
rect 2018 735 2026 885
rect 2018 729 2019 735
rect 2025 729 2026 735
rect 2018 579 2026 729
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 427 2026 573
rect 2018 421 2019 427
rect 2025 421 2026 427
rect 2018 271 2026 421
rect 2018 265 2019 271
rect 2025 265 2026 271
rect 2018 263 2026 265
rect 2018 257 2019 263
rect 2025 257 2026 263
rect 2018 91 2026 257
rect 2018 85 2019 91
rect 2025 85 2026 91
rect 2018 72 2026 85
rect 2030 4031 2038 4032
rect 2030 4025 2031 4031
rect 2037 4025 2038 4031
rect 2030 4011 2038 4025
rect 2030 4005 2031 4011
rect 2037 4005 2038 4011
rect 2030 3879 2038 4005
rect 2030 3873 2031 3879
rect 2037 3873 2038 3879
rect 2030 3855 2038 3873
rect 2030 3849 2031 3855
rect 2037 3849 2038 3855
rect 2030 3715 2038 3849
rect 2030 3709 2031 3715
rect 2037 3709 2038 3715
rect 2030 3687 2038 3709
rect 2030 3681 2031 3687
rect 2037 3681 2038 3687
rect 2030 3543 2038 3681
rect 2030 3537 2031 3543
rect 2037 3537 2038 3543
rect 2030 3519 2038 3537
rect 2030 3513 2031 3519
rect 2037 3513 2038 3519
rect 2030 3383 2038 3513
rect 2030 3377 2031 3383
rect 2037 3377 2038 3383
rect 2030 3351 2038 3377
rect 2030 3345 2031 3351
rect 2037 3345 2038 3351
rect 2030 3227 2038 3345
rect 2030 3221 2031 3227
rect 2037 3221 2038 3227
rect 2030 3191 2038 3221
rect 2030 3185 2031 3191
rect 2037 3185 2038 3191
rect 2030 3067 2038 3185
rect 2030 3061 2031 3067
rect 2037 3061 2038 3067
rect 2030 3039 2038 3061
rect 2030 3033 2031 3039
rect 2037 3033 2038 3039
rect 2030 2895 2038 3033
rect 2030 2889 2031 2895
rect 2037 2889 2038 2895
rect 2030 2855 2038 2889
rect 2030 2849 2031 2855
rect 2037 2849 2038 2855
rect 2030 2735 2038 2849
rect 2030 2729 2031 2735
rect 2037 2729 2038 2735
rect 2030 2703 2038 2729
rect 2030 2697 2031 2703
rect 2037 2697 2038 2703
rect 2030 2571 2038 2697
rect 2030 2565 2031 2571
rect 2037 2565 2038 2571
rect 2030 2547 2038 2565
rect 2030 2541 2031 2547
rect 2037 2541 2038 2547
rect 2030 2399 2038 2541
rect 2030 2393 2031 2399
rect 2037 2393 2038 2399
rect 2030 2391 2038 2393
rect 2030 2385 2031 2391
rect 2037 2385 2038 2391
rect 2030 2239 2038 2385
rect 2030 2233 2031 2239
rect 2037 2233 2038 2239
rect 2030 2231 2038 2233
rect 2030 2225 2031 2231
rect 2037 2225 2038 2231
rect 2030 2071 2038 2225
rect 2030 2065 2031 2071
rect 2037 2065 2038 2071
rect 2030 1903 2038 2065
rect 2030 1897 2031 1903
rect 2037 1897 2038 1903
rect 2030 1751 2038 1897
rect 2030 1745 2031 1751
rect 2037 1745 2038 1751
rect 2030 1595 2038 1745
rect 2030 1589 2031 1595
rect 2037 1589 2038 1595
rect 2030 1439 2038 1589
rect 2030 1433 2031 1439
rect 2037 1433 2038 1439
rect 2030 1279 2038 1433
rect 2030 1273 2031 1279
rect 2037 1273 2038 1279
rect 2030 1123 2038 1273
rect 2030 1117 2031 1123
rect 2037 1117 2038 1123
rect 2030 971 2038 1117
rect 2030 965 2031 971
rect 2037 965 2038 971
rect 2030 811 2038 965
rect 2030 805 2031 811
rect 2037 805 2038 811
rect 2030 659 2038 805
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 503 2038 653
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 347 2038 497
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 167 2038 341
rect 2030 161 2031 167
rect 2037 161 2038 167
rect 2030 72 2038 161
rect 3966 3955 3974 4032
rect 3966 3949 3967 3955
rect 3973 3949 3974 3955
rect 3966 3803 3974 3949
rect 3966 3797 3967 3803
rect 3973 3797 3974 3803
rect 3966 3635 3974 3797
rect 3966 3629 3967 3635
rect 3973 3629 3974 3635
rect 3966 3467 3974 3629
rect 3966 3461 3967 3467
rect 3973 3461 3974 3467
rect 3966 3303 3974 3461
rect 3966 3297 3967 3303
rect 3973 3297 3974 3303
rect 3966 3147 3974 3297
rect 3966 3141 3967 3147
rect 3973 3141 3974 3147
rect 3966 2987 3974 3141
rect 3966 2981 3967 2987
rect 3973 2981 3974 2987
rect 3966 2819 3974 2981
rect 3966 2813 3967 2819
rect 3973 2813 3974 2819
rect 3966 2655 3974 2813
rect 3966 2649 3967 2655
rect 3973 2649 3974 2655
rect 3966 2491 3974 2649
rect 3966 2485 3967 2491
rect 3973 2485 3974 2491
rect 3966 2323 3974 2485
rect 3966 2317 3967 2323
rect 3973 2317 3974 2323
rect 3966 1679 3974 2317
rect 3966 1673 3967 1679
rect 3973 1673 3974 1679
rect 3966 271 3974 1673
rect 3966 265 3967 271
rect 3973 265 3974 271
rect 3966 72 3974 265
rect 3978 4031 3986 4032
rect 3978 4025 3979 4031
rect 3985 4025 3986 4031
rect 3978 3879 3986 4025
rect 3978 3873 3979 3879
rect 3985 3873 3986 3879
rect 3978 3715 3986 3873
rect 3978 3709 3979 3715
rect 3985 3709 3986 3715
rect 3978 3543 3986 3709
rect 3978 3537 3979 3543
rect 3985 3537 3986 3543
rect 3978 3383 3986 3537
rect 3978 3377 3979 3383
rect 3985 3377 3986 3383
rect 3978 3227 3986 3377
rect 3978 3221 3979 3227
rect 3985 3221 3986 3227
rect 3978 3067 3986 3221
rect 3978 3061 3979 3067
rect 3985 3061 3986 3067
rect 3978 2895 3986 3061
rect 3978 2889 3979 2895
rect 3985 2889 3986 2895
rect 3978 2735 3986 2889
rect 3978 2729 3979 2735
rect 3985 2729 3986 2735
rect 3978 2571 3986 2729
rect 3978 2565 3979 2571
rect 3985 2565 3986 2571
rect 3978 2399 3986 2565
rect 3978 2393 3979 2399
rect 3985 2393 3986 2399
rect 3978 2239 3986 2393
rect 3978 2233 3979 2239
rect 3985 2233 3986 2239
rect 3978 72 3986 2233
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220370
transform 1 0 3936 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220370
transform 1 0 2040 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220370
transform 1 0 3936 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220370
transform 1 0 2040 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220370
transform 1 0 3936 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220370
transform 1 0 2040 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220370
transform 1 0 3936 0 -1 3772
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220370
transform 1 0 2040 0 -1 3772
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220370
transform 1 0 3936 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220370
transform 1 0 2040 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220370
transform 1 0 3936 0 -1 3604
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220370
transform 1 0 2040 0 -1 3604
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220370
transform 1 0 3936 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220370
transform 1 0 2040 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220370
transform 1 0 3936 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220370
transform 1 0 2040 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220370
transform 1 0 3936 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220370
transform 1 0 2040 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220370
transform 1 0 3936 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220370
transform 1 0 2040 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220370
transform 1 0 3936 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220370
transform 1 0 2040 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220370
transform 1 0 3936 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220370
transform 1 0 2040 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220370
transform 1 0 3936 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220370
transform 1 0 2040 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220370
transform 1 0 3936 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220370
transform 1 0 2040 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220370
transform 1 0 3936 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220370
transform 1 0 2040 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220370
transform 1 0 3936 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220370
transform 1 0 2040 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220370
transform 1 0 3936 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220370
transform 1 0 2040 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220370
transform 1 0 3936 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220370
transform 1 0 2040 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220370
transform 1 0 3936 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220370
transform 1 0 2040 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220370
transform 1 0 3936 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220370
transform 1 0 2040 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220370
transform 1 0 3936 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220370
transform 1 0 2040 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220370
transform 1 0 3936 0 -1 2292
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220370
transform 1 0 2040 0 -1 2292
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220370
transform 1 0 3936 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220370
transform 1 0 2040 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220370
transform 1 0 3936 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220370
transform 1 0 2040 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220370
transform 1 0 3936 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220370
transform 1 0 2040 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220370
transform 1 0 3936 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220370
transform 1 0 2040 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220370
transform 1 0 3936 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220370
transform 1 0 2040 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220370
transform 1 0 3936 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220370
transform 1 0 2040 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220370
transform 1 0 3936 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220370
transform 1 0 2040 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220370
transform 1 0 3936 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220370
transform 1 0 2040 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220370
transform 1 0 3936 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220370
transform 1 0 2040 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220370
transform 1 0 3936 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220370
transform 1 0 2040 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220370
transform 1 0 3936 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220370
transform 1 0 2040 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220370
transform 1 0 3936 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220370
transform 1 0 2040 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220370
transform 1 0 3936 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220370
transform 1 0 2040 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220370
transform 1 0 3936 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220370
transform 1 0 2040 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220370
transform 1 0 3936 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220370
transform 1 0 2040 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220370
transform 1 0 3936 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220370
transform 1 0 2040 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220370
transform 1 0 3936 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220370
transform 1 0 2040 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220370
transform 1 0 3936 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220370
transform 1 0 2040 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220370
transform 1 0 3936 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220370
transform 1 0 2040 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220370
transform 1 0 3936 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220370
transform 1 0 2040 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220370
transform 1 0 3936 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220370
transform 1 0 2040 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220370
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220370
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220370
transform 1 0 3936 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220370
transform 1 0 2040 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220370
transform 1 0 3936 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220370
transform 1 0 2040 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220370
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220370
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220370
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220370
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220370
transform 1 0 3936 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220370
transform 1 0 2040 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220370
transform 1 0 2000 0 1 3960
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220370
transform 1 0 104 0 1 3960
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220370
transform 1 0 2000 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220370
transform 1 0 104 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220370
transform 1 0 2000 0 1 3804
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220370
transform 1 0 104 0 1 3804
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220370
transform 1 0 2000 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220370
transform 1 0 104 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220370
transform 1 0 2000 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220370
transform 1 0 104 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220370
transform 1 0 2000 0 -1 3572
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220370
transform 1 0 104 0 -1 3572
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220370
transform 1 0 2000 0 1 3468
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220370
transform 1 0 104 0 1 3468
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220370
transform 1 0 2000 0 -1 3404
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220370
transform 1 0 104 0 -1 3404
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220370
transform 1 0 2000 0 1 3300
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220370
transform 1 0 104 0 1 3300
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220370
transform 1 0 2000 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220370
transform 1 0 104 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220370
transform 1 0 2000 0 1 3140
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220370
transform 1 0 104 0 1 3140
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220370
transform 1 0 2000 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220370
transform 1 0 104 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220370
transform 1 0 2000 0 1 2988
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220370
transform 1 0 104 0 1 2988
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220370
transform 1 0 2000 0 -1 2908
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220370
transform 1 0 104 0 -1 2908
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220370
transform 1 0 2000 0 1 2804
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220370
transform 1 0 104 0 1 2804
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220370
transform 1 0 2000 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220370
transform 1 0 104 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220370
transform 1 0 2000 0 1 2652
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220370
transform 1 0 104 0 1 2652
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220370
transform 1 0 2000 0 -1 2596
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220370
transform 1 0 104 0 -1 2596
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220370
transform 1 0 2000 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220370
transform 1 0 104 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220370
transform 1 0 2000 0 -1 2436
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220370
transform 1 0 104 0 -1 2436
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220370
transform 1 0 2000 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220370
transform 1 0 104 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220370
transform 1 0 2000 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220370
transform 1 0 104 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220370
transform 1 0 2000 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220370
transform 1 0 104 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220370
transform 1 0 2000 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220370
transform 1 0 104 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220370
transform 1 0 2000 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220370
transform 1 0 104 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220370
transform 1 0 2000 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220370
transform 1 0 104 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220370
transform 1 0 2000 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220370
transform 1 0 104 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220370
transform 1 0 2000 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220370
transform 1 0 104 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220370
transform 1 0 2000 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220370
transform 1 0 104 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220370
transform 1 0 2000 0 -1 1640
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220370
transform 1 0 104 0 -1 1640
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220370
transform 1 0 2000 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220370
transform 1 0 104 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220370
transform 1 0 2000 0 -1 1484
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220370
transform 1 0 104 0 -1 1484
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220370
transform 1 0 2000 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220370
transform 1 0 104 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220370
transform 1 0 2000 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220370
transform 1 0 104 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220370
transform 1 0 2000 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220370
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220370
transform 1 0 2000 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220370
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220370
transform 1 0 2000 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220370
transform 1 0 104 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220370
transform 1 0 2000 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220370
transform 1 0 104 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220370
transform 1 0 2000 0 1 920
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220370
transform 1 0 104 0 1 920
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220370
transform 1 0 2000 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220370
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220370
transform 1 0 2000 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220370
transform 1 0 104 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220370
transform 1 0 2000 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220370
transform 1 0 104 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220370
transform 1 0 2000 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220370
transform 1 0 104 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220370
transform 1 0 2000 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220370
transform 1 0 104 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220370
transform 1 0 2000 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220370
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220370
transform 1 0 2000 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220370
transform 1 0 104 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220370
transform 1 0 2000 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220370
transform 1 0 104 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220370
transform 1 0 2000 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220370
transform 1 0 104 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220370
transform 1 0 2000 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220370
transform 1 0 104 0 1 116
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220370
transform 1 0 3832 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220370
transform 1 0 3736 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220370
transform 1 0 3800 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220370
transform 1 0 3784 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220370
transform 1 0 3600 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220370
transform 1 0 3416 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220370
transform 1 0 3600 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220370
transform 1 0 3632 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220370
transform 1 0 3528 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220370
transform 1 0 3424 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220370
transform 1 0 3320 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220370
transform 1 0 3216 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220370
transform 1 0 3104 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220370
transform 1 0 2984 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220370
transform 1 0 2864 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220370
transform 1 0 3400 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220370
transform 1 0 3208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220370
transform 1 0 3024 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220370
transform 1 0 2848 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220370
transform 1 0 3064 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220370
transform 1 0 3240 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220370
transform 1 0 3224 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220370
transform 1 0 3128 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220370
transform 1 0 3032 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220370
transform 1 0 2936 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220370
transform 1 0 2840 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220370
transform 1 0 2888 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220370
transform 1 0 3056 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220370
transform 1 0 3376 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220370
transform 1 0 3216 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220370
transform 1 0 3136 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220370
transform 1 0 2952 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220370
transform 1 0 3312 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220370
transform 1 0 3488 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220370
transform 1 0 3672 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220370
transform 1 0 3528 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220370
transform 1 0 3368 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220370
transform 1 0 3200 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220370
transform 1 0 3016 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220370
transform 1 0 3632 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220370
transform 1 0 3432 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220370
transform 1 0 3232 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220370
transform 1 0 3040 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220370
transform 1 0 2848 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220370
transform 1 0 3496 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220370
transform 1 0 3280 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220370
transform 1 0 3072 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220370
transform 1 0 2872 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220370
transform 1 0 3600 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220370
transform 1 0 3384 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220370
transform 1 0 3184 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220370
transform 1 0 3008 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220370
transform 1 0 2856 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220370
transform 1 0 3448 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220370
transform 1 0 3264 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220370
transform 1 0 3096 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220370
transform 1 0 2944 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220370
transform 1 0 3024 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220370
transform 1 0 2816 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220370
transform 1 0 2752 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220370
transform 1 0 2704 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220370
transform 1 0 2640 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220370
transform 1 0 2880 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220370
transform 1 0 2800 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220370
transform 1 0 2936 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220370
transform 1 0 3176 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220370
transform 1 0 3336 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220370
transform 1 0 3440 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220370
transform 1 0 3256 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220370
transform 1 0 3088 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220370
transform 1 0 3064 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220370
transform 1 0 2904 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220370
transform 1 0 3432 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220370
transform 1 0 3240 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220370
transform 1 0 3064 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220370
transform 1 0 2896 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220370
transform 1 0 3240 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220370
transform 1 0 3424 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220370
transform 1 0 3272 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220370
transform 1 0 3104 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220370
transform 1 0 2928 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220370
transform 1 0 3264 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220370
transform 1 0 3432 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220370
transform 1 0 3600 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220370
transform 1 0 3440 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220370
transform 1 0 3616 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220370
transform 1 0 3608 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220370
transform 1 0 3624 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220370
transform 1 0 3632 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220370
transform 1 0 3496 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220370
transform 1 0 3664 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220370
transform 1 0 3640 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220370
transform 1 0 3712 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220370
transform 1 0 3688 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220370
transform 1 0 3696 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220370
transform 1 0 3536 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220370
transform 1 0 3832 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220370
transform 1 0 3832 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220370
transform 1 0 3832 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220370
transform 1 0 3832 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220370
transform 1 0 3816 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220370
transform 1 0 3832 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220370
transform 1 0 3832 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220370
transform 1 0 3832 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220370
transform 1 0 3824 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220370
transform 1 0 3800 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220370
transform 1 0 3776 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220370
transform 1 0 3792 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220370
transform 1 0 3456 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220370
transform 1 0 3560 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220370
transform 1 0 3688 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220370
transform 1 0 3520 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220370
transform 1 0 3352 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220370
transform 1 0 3416 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220370
transform 1 0 3256 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220370
transform 1 0 3120 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220370
transform 1 0 3088 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220370
transform 1 0 2904 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220370
transform 1 0 2784 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220370
transform 1 0 2424 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220370
transform 1 0 2904 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220370
transform 1 0 3088 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220370
transform 1 0 3016 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220370
transform 1 0 3184 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220370
transform 1 0 3120 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220370
transform 1 0 3008 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220370
transform 1 0 2904 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220370
transform 1 0 2800 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220370
transform 1 0 2696 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220370
transform 1 0 2848 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220370
transform 1 0 3064 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220370
transform 1 0 3296 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220370
transform 1 0 3536 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220370
transform 1 0 3664 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220370
transform 1 0 3480 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220370
transform 1 0 3296 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220370
transform 1 0 3120 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220370
transform 1 0 2952 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220370
transform 1 0 3288 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220370
transform 1 0 3408 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220370
transform 1 0 3536 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220370
transform 1 0 3664 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220370
transform 1 0 3720 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220370
transform 1 0 3584 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220370
transform 1 0 3448 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220370
transform 1 0 3304 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220370
transform 1 0 3160 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220370
transform 1 0 3688 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220370
transform 1 0 3520 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220370
transform 1 0 3360 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220370
transform 1 0 3200 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220370
transform 1 0 3040 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220370
transform 1 0 3584 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220370
transform 1 0 3400 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220370
transform 1 0 3216 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220370
transform 1 0 3040 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220370
transform 1 0 2872 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220370
transform 1 0 3608 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220370
transform 1 0 3368 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220370
transform 1 0 3136 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220370
transform 1 0 2928 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220370
transform 1 0 2744 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220370
transform 1 0 3096 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220370
transform 1 0 2928 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220370
transform 1 0 2768 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220370
transform 1 0 2600 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220370
transform 1 0 2424 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220370
transform 1 0 2552 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220370
transform 1 0 2744 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220370
transform 1 0 2944 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220370
transform 1 0 3160 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220370
transform 1 0 3384 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220370
transform 1 0 3496 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220370
transform 1 0 3256 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220370
transform 1 0 3024 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220370
transform 1 0 2816 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220370
transform 1 0 2984 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220370
transform 1 0 3168 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220370
transform 1 0 3160 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220370
transform 1 0 2992 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220370
transform 1 0 3328 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220370
transform 1 0 3240 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220370
transform 1 0 3096 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220370
transform 1 0 3176 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220370
transform 1 0 3304 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220370
transform 1 0 3568 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220370
transform 1 0 3432 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220370
transform 1 0 3384 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220370
transform 1 0 3536 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220370
transform 1 0 3696 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220370
transform 1 0 3680 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220370
transform 1 0 3504 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220370
transform 1 0 3512 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220370
transform 1 0 3344 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220370
transform 1 0 3680 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220370
transform 1 0 3736 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220370
transform 1 0 3616 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220370
transform 1 0 3776 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220370
transform 1 0 3792 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220370
transform 1 0 3784 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220370
transform 1 0 3704 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220370
transform 1 0 3832 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220370
transform 1 0 3832 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220370
transform 1 0 3832 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220370
transform 1 0 3832 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220370
transform 1 0 3832 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220370
transform 1 0 3832 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220370
transform 1 0 3832 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220370
transform 1 0 3832 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220370
transform 1 0 3832 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220370
transform 1 0 3832 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220370
transform 1 0 3832 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220370
transform 1 0 3832 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220370
transform 1 0 3736 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220370
transform 1 0 3632 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220370
transform 1 0 3528 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220370
transform 1 0 3616 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220370
transform 1 0 3392 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220370
transform 1 0 3424 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220370
transform 1 0 3320 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220370
transform 1 0 3208 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220370
transform 1 0 3096 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220370
transform 1 0 2976 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220370
transform 1 0 2896 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220370
transform 1 0 3168 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220370
transform 1 0 3440 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220370
transform 1 0 3320 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220370
transform 1 0 3160 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220370
transform 1 0 3008 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220370
transform 1 0 2928 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220370
transform 1 0 3088 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220370
transform 1 0 3256 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220370
transform 1 0 3152 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220370
transform 1 0 3296 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220370
transform 1 0 3264 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220370
transform 1 0 3400 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220370
transform 1 0 3480 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220370
transform 1 0 3344 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220370
transform 1 0 3320 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220370
transform 1 0 3560 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220370
transform 1 0 3512 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220370
transform 1 0 3312 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220370
transform 1 0 3720 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220370
transform 1 0 3728 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220370
transform 1 0 3528 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220370
transform 1 0 3328 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220370
transform 1 0 3320 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220370
transform 1 0 3488 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220370
transform 1 0 3656 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220370
transform 1 0 3528 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220370
transform 1 0 3408 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220370
transform 1 0 3288 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220370
transform 1 0 3168 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220370
transform 1 0 3048 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220370
transform 1 0 2920 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220370
transform 1 0 2784 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220370
transform 1 0 3152 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220370
transform 1 0 2984 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220370
transform 1 0 2944 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220370
transform 1 0 3136 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220370
transform 1 0 3112 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220370
transform 1 0 2904 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220370
transform 1 0 3088 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220370
transform 1 0 3216 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220370
transform 1 0 3136 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220370
transform 1 0 3016 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220370
transform 1 0 2880 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220370
transform 1 0 2768 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220370
transform 1 0 2856 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220370
transform 1 0 2696 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220370
transform 1 0 2624 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220370
transform 1 0 2336 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220370
transform 1 0 2856 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220370
transform 1 0 2736 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220370
transform 1 0 2608 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220370
transform 1 0 2480 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220370
transform 1 0 2400 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220370
transform 1 0 2568 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220370
transform 1 0 2760 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220370
transform 1 0 2960 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220370
transform 1 0 3176 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220370
transform 1 0 3048 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220370
transform 1 0 2920 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220370
transform 1 0 2792 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220370
transform 1 0 2664 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220370
transform 1 0 2544 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220370
transform 1 0 2960 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220370
transform 1 0 2824 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220370
transform 1 0 2688 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220370
transform 1 0 2560 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220370
transform 1 0 2432 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220370
transform 1 0 2824 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220370
transform 1 0 2656 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220370
transform 1 0 2488 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220370
transform 1 0 2328 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220370
transform 1 0 2800 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220370
transform 1 0 2616 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220370
transform 1 0 2440 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220370
transform 1 0 2272 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220370
transform 1 0 2120 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220370
transform 1 0 2632 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220370
transform 1 0 2464 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220370
transform 1 0 2312 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220370
transform 1 0 2176 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220370
transform 1 0 2064 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220370
transform 1 0 2376 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220370
transform 1 0 2208 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220370
transform 1 0 2064 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220370
transform 1 0 1896 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220370
transform 1 0 1784 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220370
transform 1 0 1656 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220370
transform 1 0 1896 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220370
transform 1 0 2064 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220370
transform 1 0 2240 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220370
transform 1 0 2168 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220370
transform 1 0 2064 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220370
transform 1 0 2304 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220370
transform 1 0 2584 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220370
transform 1 0 2440 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220370
transform 1 0 2400 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220370
transform 1 0 2248 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220370
transform 1 0 2104 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220370
transform 1 0 2552 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220370
transform 1 0 2712 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220370
transform 1 0 2576 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220370
transform 1 0 2424 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220370
transform 1 0 2280 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220370
transform 1 0 2728 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220370
transform 1 0 2880 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220370
transform 1 0 3000 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220370
transform 1 0 2832 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220370
transform 1 0 2664 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220370
transform 1 0 2496 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220370
transform 1 0 2488 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220370
transform 1 0 2584 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220370
transform 1 0 2688 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220370
transform 1 0 2800 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220370
transform 1 0 3168 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220370
transform 1 0 3040 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220370
transform 1 0 2920 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220370
transform 1 0 2784 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220370
transform 1 0 2616 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220370
transform 1 0 2432 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220370
transform 1 0 2240 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220370
transform 1 0 2504 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220370
transform 1 0 2664 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220370
transform 1 0 2592 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220370
transform 1 0 2488 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220370
transform 1 0 2672 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220370
transform 1 0 2840 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220370
transform 1 0 2704 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220370
transform 1 0 2512 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220370
transform 1 0 2360 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220370
transform 1 0 2224 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220370
transform 1 0 2176 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220370
transform 1 0 2280 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220370
transform 1 0 2384 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220370
transform 1 0 2360 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220370
transform 1 0 2224 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220370
transform 1 0 2088 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220370
transform 1 0 2064 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220370
transform 1 0 1840 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220370
transform 1 0 1576 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220370
transform 1 0 1440 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220370
transform 1 0 1304 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220370
transform 1 0 1272 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220370
transform 1 0 1552 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220370
transform 1 0 1408 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220370
transform 1 0 1392 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220370
transform 1 0 1576 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220370
transform 1 0 1624 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220370
transform 1 0 1440 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220370
transform 1 0 1256 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220370
transform 1 0 1320 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220370
transform 1 0 1560 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220370
transform 1 0 1440 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220370
transform 1 0 1256 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220370
transform 1 0 1080 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220370
transform 1 0 912 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220370
transform 1 0 1088 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220370
transform 1 0 1088 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220370
transform 1 0 928 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220370
transform 1 0 1040 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220370
transform 1 0 1208 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220370
transform 1 0 1136 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220370
transform 1 0 1168 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220370
transform 1 0 1144 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220370
transform 1 0 1312 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220370
transform 1 0 1432 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220370
transform 1 0 1272 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220370
transform 1 0 1120 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220370
transform 1 0 1160 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220370
transform 1 0 1344 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220370
transform 1 0 1360 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220370
transform 1 0 1176 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220370
transform 1 0 1176 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220370
transform 1 0 1344 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220370
transform 1 0 1536 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220370
transform 1 0 1728 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220370
transform 1 0 1648 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220370
transform 1 0 1856 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220370
transform 1 0 1888 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220370
transform 1 0 1712 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220370
transform 1 0 1832 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220370
transform 1 0 1680 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220370
transform 1 0 1536 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220370
transform 1 0 1616 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220370
transform 1 0 1392 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220370
transform 1 0 1240 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220370
transform 1 0 1184 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220370
transform 1 0 1360 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220370
transform 1 0 1536 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220370
transform 1 0 1440 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220370
transform 1 0 1240 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220370
transform 1 0 1040 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220370
transform 1 0 1152 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220370
transform 1 0 968 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220370
transform 1 0 872 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220370
transform 1 0 1032 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220370
transform 1 0 984 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220370
transform 1 0 976 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220370
transform 1 0 976 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220370
transform 1 0 840 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220370
transform 1 0 856 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220370
transform 1 0 992 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220370
transform 1 0 1040 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220370
transform 1 0 1000 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220370
transform 1 0 864 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220370
transform 1 0 888 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220370
transform 1 0 744 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220370
transform 1 0 776 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220370
transform 1 0 872 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220370
transform 1 0 672 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220370
transform 1 0 584 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220370
transform 1 0 744 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220370
transform 1 0 968 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220370
transform 1 0 760 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220370
transform 1 0 544 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220370
transform 1 0 704 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220370
transform 1 0 896 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220370
transform 1 0 920 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220370
transform 1 0 768 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220370
transform 1 0 600 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220370
transform 1 0 536 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220370
transform 1 0 704 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220370
transform 1 0 760 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220370
transform 1 0 632 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220370
transform 1 0 496 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220370
transform 1 0 600 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220370
transform 1 0 736 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220370
transform 1 0 872 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220370
transform 1 0 992 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220370
transform 1 0 808 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220370
transform 1 0 624 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220370
transform 1 0 440 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220370
transform 1 0 272 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220370
transform 1 0 464 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220370
transform 1 0 344 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220370
transform 1 0 232 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220370
transform 1 0 216 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220370
transform 1 0 360 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220370
transform 1 0 360 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220370
transform 1 0 168 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220370
transform 1 0 128 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220370
transform 1 0 264 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220370
transform 1 0 432 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220370
transform 1 0 504 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220370
transform 1 0 304 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220370
transform 1 0 128 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220370
transform 1 0 128 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220370
transform 1 0 320 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220370
transform 1 0 264 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220370
transform 1 0 128 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220370
transform 1 0 424 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220370
transform 1 0 320 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220370
transform 1 0 152 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220370
transform 1 0 488 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220370
transform 1 0 488 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220370
transform 1 0 352 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220370
transform 1 0 216 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220370
transform 1 0 632 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220370
transform 1 0 608 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220370
transform 1 0 488 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220370
transform 1 0 368 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220370
transform 1 0 504 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220370
transform 1 0 616 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220370
transform 1 0 736 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220370
transform 1 0 904 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220370
transform 1 0 776 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220370
transform 1 0 656 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220370
transform 1 0 544 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220370
transform 1 0 496 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220370
transform 1 0 608 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220370
transform 1 0 728 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220370
transform 1 0 712 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220370
transform 1 0 584 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220370
transform 1 0 456 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220370
transform 1 0 336 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220370
transform 1 0 792 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220370
transform 1 0 616 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220370
transform 1 0 448 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220370
transform 1 0 288 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220370
transform 1 0 152 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220370
transform 1 0 792 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220370
transform 1 0 600 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220370
transform 1 0 416 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220370
transform 1 0 248 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220370
transform 1 0 128 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220370
transform 1 0 712 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220370
transform 1 0 552 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220370
transform 1 0 392 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220370
transform 1 0 240 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220370
transform 1 0 128 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220370
transform 1 0 128 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220370
transform 1 0 256 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220370
transform 1 0 424 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220370
transform 1 0 784 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220370
transform 1 0 600 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220370
transform 1 0 472 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220370
transform 1 0 304 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220370
transform 1 0 152 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220370
transform 1 0 848 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220370
transform 1 0 656 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220370
transform 1 0 536 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220370
transform 1 0 400 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220370
transform 1 0 1016 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220370
transform 1 0 848 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220370
transform 1 0 688 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220370
transform 1 0 584 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220370
transform 1 0 416 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220370
transform 1 0 368 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220370
transform 1 0 296 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220370
transform 1 0 440 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220370
transform 1 0 440 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220370
transform 1 0 248 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220370
transform 1 0 248 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220370
transform 1 0 152 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220370
transform 1 0 304 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220370
transform 1 0 256 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220370
transform 1 0 128 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220370
transform 1 0 128 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220370
transform 1 0 240 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220370
transform 1 0 288 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220370
transform 1 0 128 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220370
transform 1 0 128 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220370
transform 1 0 280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220370
transform 1 0 280 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220370
transform 1 0 128 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220370
transform 1 0 152 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220370
transform 1 0 344 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220370
transform 1 0 376 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220370
transform 1 0 216 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220370
transform 1 0 224 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220370
transform 1 0 128 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220370
transform 1 0 320 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220370
transform 1 0 416 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220370
transform 1 0 520 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220370
transform 1 0 896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220370
transform 1 0 768 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220370
transform 1 0 640 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220370
transform 1 0 536 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220370
transform 1 0 696 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220370
transform 1 0 856 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220370
transform 1 0 952 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220370
transform 1 0 752 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220370
transform 1 0 544 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220370
transform 1 0 440 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220370
transform 1 0 592 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220370
transform 1 0 744 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220370
transform 1 0 760 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220370
transform 1 0 608 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220370
transform 1 0 448 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220370
transform 1 0 472 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220370
transform 1 0 656 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220370
transform 1 0 680 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220370
transform 1 0 520 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220370
transform 1 0 376 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220370
transform 1 0 424 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220370
transform 1 0 616 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220370
transform 1 0 816 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220370
transform 1 0 768 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220370
transform 1 0 616 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220370
transform 1 0 464 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220370
transform 1 0 440 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220370
transform 1 0 632 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220370
transform 1 0 816 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220370
transform 1 0 992 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220370
transform 1 0 968 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220370
transform 1 0 800 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220370
transform 1 0 624 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220370
transform 1 0 584 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220370
transform 1 0 848 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220370
transform 1 0 720 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220370
transform 1 0 704 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220370
transform 1 0 592 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220370
transform 1 0 480 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220370
transform 1 0 752 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220370
transform 1 0 920 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220370
transform 1 0 1088 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220370
transform 1 0 1112 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220370
transform 1 0 960 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220370
transform 1 0 824 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220370
transform 1 0 1272 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220370
transform 1 0 1440 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220370
transform 1 0 1424 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220370
transform 1 0 1304 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220370
transform 1 0 1192 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220370
transform 1 0 1080 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220370
transform 1 0 968 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220370
transform 1 0 1120 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220370
transform 1 0 1264 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220370
transform 1 0 1408 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220370
transform 1 0 1544 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220370
transform 1 0 1688 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220370
transform 1 0 1776 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220370
transform 1 0 1624 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220370
transform 1 0 1472 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220370
transform 1 0 1320 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220370
transform 1 0 1160 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220370
transform 1 0 1576 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220370
transform 1 0 1408 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220370
transform 1 0 1248 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220370
transform 1 0 1088 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220370
transform 1 0 928 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220370
transform 1 0 1008 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220370
transform 1 0 1200 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220370
transform 1 0 1536 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220370
transform 1 0 1296 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220370
transform 1 0 1072 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220370
transform 1 0 864 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220370
transform 1 0 840 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220370
transform 1 0 1208 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220370
transform 1 0 1024 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220370
transform 1 0 896 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220370
transform 1 0 896 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220370
transform 1 0 1072 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220370
transform 1 0 1264 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220370
transform 1 0 1152 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220370
transform 1 0 1696 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220370
transform 1 0 1472 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220370
transform 1 0 1280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220370
transform 1 0 1152 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220370
transform 1 0 1024 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220370
transform 1 0 1408 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220370
transform 1 0 1392 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220370
transform 1 0 1584 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220370
transform 1 0 1776 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220370
transform 1 0 1776 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220370
transform 1 0 1560 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220370
transform 1 0 1384 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220370
transform 1 0 1736 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220370
transform 1 0 1896 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220370
transform 1 0 1744 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220370
transform 1 0 1896 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220370
transform 1 0 2064 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220370
transform 1 0 2248 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220370
transform 1 0 2448 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220370
transform 1 0 2424 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220370
transform 1 0 2224 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220370
transform 1 0 2064 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220370
transform 1 0 2392 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220370
transform 1 0 2576 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220370
transform 1 0 2768 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220370
transform 1 0 2720 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220370
transform 1 0 2552 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220370
transform 1 0 2384 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220370
transform 1 0 2216 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220370
transform 1 0 2456 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220370
transform 1 0 2552 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220370
transform 1 0 2648 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220370
transform 1 0 2744 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220370
transform 1 0 2904 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220370
transform 1 0 2752 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220370
transform 1 0 2616 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220370
transform 1 0 2496 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220370
transform 1 0 2392 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220370
transform 1 0 2680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220370
transform 1 0 2512 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220370
transform 1 0 2344 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220370
transform 1 0 2184 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220370
transform 1 0 2736 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220370
transform 1 0 2608 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220370
transform 1 0 2480 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220370
transform 1 0 2360 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220370
transform 1 0 2256 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220370
transform 1 0 2160 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220370
transform 1 0 2064 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220370
transform 1 0 1896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220370
transform 1 0 1896 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220370
transform 1 0 1800 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220370
transform 1 0 1696 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220370
transform 1 0 1584 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220370
transform 1 0 1480 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220370
transform 1 0 1376 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220370
transform 1 0 1264 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220370
transform 1 0 1144 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220370
transform 1 0 1024 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220370
transform 1 0 1024 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220370
transform 1 0 1192 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220370
transform 1 0 1360 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220370
transform 1 0 1536 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220370
transform 1 0 1720 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220370
transform 1 0 1704 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220370
transform 1 0 1520 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220370
transform 1 0 1336 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220370
transform 1 0 1888 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220370
transform 1 0 1896 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220370
transform 1 0 2064 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220370
transform 1 0 2064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220370
transform 1 0 2208 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220370
transform 1 0 2624 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220370
transform 1 0 2824 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220370
transform 1 0 2648 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220370
transform 1 0 2680 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220370
transform 1 0 2488 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220370
transform 1 0 2304 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220370
transform 1 0 2336 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220370
transform 1 0 2432 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220370
transform 1 0 2528 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220370
transform 1 0 2728 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220370
transform 1 0 2624 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220370
transform 1 0 2608 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220370
transform 1 0 2512 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220370
transform 1 0 2416 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220370
transform 1 0 2448 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220370
transform 1 0 2544 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220370
transform 1 0 2688 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220370
transform 1 0 2592 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220370
transform 1 0 2496 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220370
transform 1 0 2400 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220370
transform 1 0 2760 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220370
transform 1 0 2632 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220370
transform 1 0 2520 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220370
transform 1 0 2408 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220370
transform 1 0 2304 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220370
transform 1 0 2736 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220370
transform 1 0 2576 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220370
transform 1 0 2424 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220370
transform 1 0 2280 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220370
transform 1 0 2144 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220370
transform 1 0 2744 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220370
transform 1 0 2560 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220370
transform 1 0 2376 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220370
transform 1 0 2200 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220370
transform 1 0 2064 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220370
transform 1 0 2704 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220370
transform 1 0 2488 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220370
transform 1 0 2264 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220370
transform 1 0 2064 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220370
transform 1 0 1896 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220370
transform 1 0 1800 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220370
transform 1 0 1896 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220370
transform 1 0 2064 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220370
transform 1 0 2488 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220370
transform 1 0 2264 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220370
transform 1 0 2064 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220370
transform 1 0 1896 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220370
transform 1 0 1680 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220370
transform 1 0 1560 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220370
transform 1 0 1440 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220370
transform 1 0 1312 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220370
transform 1 0 1544 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220370
transform 1 0 1728 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220370
transform 1 0 1728 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220370
transform 1 0 1536 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220370
transform 1 0 1592 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220370
transform 1 0 1480 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220370
transform 1 0 1656 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220370
transform 1 0 1712 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220370
transform 1 0 1696 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220370
transform 1 0 1768 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220370
transform 1 0 1816 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220370
transform 1 0 1808 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220370
transform 1 0 1808 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220370
transform 1 0 1624 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220370
transform 1 0 1728 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220370
transform 1 0 1544 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220370
transform 1 0 1360 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220370
transform 1 0 1168 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220370
transform 1 0 1520 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220370
transform 1 0 1384 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220370
transform 1 0 1232 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220370
transform 1 0 1072 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220370
transform 1 0 1632 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220370
transform 1 0 1488 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220370
transform 1 0 1352 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220370
transform 1 0 1216 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220370
transform 1 0 1072 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220370
transform 1 0 1416 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220370
transform 1 0 1272 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220370
transform 1 0 1136 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220370
transform 1 0 1000 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220370
transform 1 0 856 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220370
transform 1 0 880 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220370
transform 1 0 992 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220370
transform 1 0 1104 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220370
transform 1 0 1344 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220370
transform 1 0 1224 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220370
transform 1 0 1144 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220370
transform 1 0 1008 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220370
transform 1 0 1280 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220370
transform 1 0 1560 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220370
transform 1 0 1416 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220370
transform 1 0 1352 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220370
transform 1 0 1176 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220370
transform 1 0 1520 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220370
transform 1 0 1688 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220370
transform 1 0 1856 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220370
transform 1 0 1856 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220370
transform 1 0 1760 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220370
transform 1 0 1664 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220370
transform 1 0 1568 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220370
transform 1 0 1472 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220370
transform 1 0 1424 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220370
transform 1 0 1544 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220370
transform 1 0 1664 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220370
transform 1 0 1896 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220370
transform 1 0 1792 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220370
transform 1 0 1744 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220370
transform 1 0 1568 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220370
transform 1 0 1896 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220370
transform 1 0 1896 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220370
transform 1 0 2064 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220370
transform 1 0 2064 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220370
transform 1 0 2536 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220370
transform 1 0 2368 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220370
transform 1 0 2200 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220370
transform 1 0 2120 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220370
transform 1 0 2288 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220370
transform 1 0 2448 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220370
transform 1 0 2608 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220370
transform 1 0 2608 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220370
transform 1 0 2472 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220370
transform 1 0 2344 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220370
transform 1 0 2744 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220370
transform 1 0 2776 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220370
transform 1 0 2888 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220370
transform 1 0 3008 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220370
transform 1 0 3096 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220370
transform 1 0 2976 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220370
transform 1 0 2864 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220370
transform 1 0 2760 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220370
transform 1 0 2664 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220370
transform 1 0 2672 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220370
transform 1 0 2576 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220370
transform 1 0 2480 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220370
transform 1 0 2568 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220370
transform 1 0 2472 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220370
transform 1 0 2376 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220370
transform 1 0 2280 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220370
transform 1 0 2864 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220370
transform 1 0 2648 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220370
transform 1 0 2448 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220370
transform 1 0 2264 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220370
transform 1 0 2104 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220370
transform 1 0 2688 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220370
transform 1 0 2472 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220370
transform 1 0 2256 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220370
transform 1 0 2064 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220370
transform 1 0 2064 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220370
transform 1 0 2192 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220370
transform 1 0 2368 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220370
transform 1 0 2744 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220370
transform 1 0 2552 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220370
transform 1 0 2512 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220370
transform 1 0 2376 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220370
transform 1 0 2248 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220370
transform 1 0 2824 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220370
transform 1 0 2664 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220370
transform 1 0 2640 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220370
transform 1 0 2496 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220370
transform 1 0 2352 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220370
transform 1 0 2208 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220370
transform 1 0 2072 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220370
transform 1 0 2064 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220370
transform 1 0 1896 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220370
transform 1 0 1768 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220370
transform 1 0 1616 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220370
transform 1 0 1464 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220370
transform 1 0 1304 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220370
transform 1 0 1144 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220370
transform 1 0 1456 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220370
transform 1 0 1320 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220370
transform 1 0 1192 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220370
transform 1 0 1064 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220370
transform 1 0 936 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220370
transform 1 0 1032 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220370
transform 1 0 1184 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220370
transform 1 0 1336 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220370
transform 1 0 1488 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220370
transform 1 0 1640 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220370
transform 1 0 1496 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220370
transform 1 0 1304 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220370
transform 1 0 1688 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220370
transform 1 0 1880 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220370
transform 1 0 1784 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220370
transform 1 0 1624 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220370
transform 1 0 1472 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220370
transform 1 0 1320 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220370
transform 1 0 1168 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220370
transform 1 0 1536 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220370
transform 1 0 1368 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220370
transform 1 0 1208 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220370
transform 1 0 1048 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220370
transform 1 0 1360 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220370
transform 1 0 1224 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220370
transform 1 0 1088 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220370
transform 1 0 960 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220370
transform 1 0 824 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220370
transform 1 0 808 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220370
transform 1 0 960 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220370
transform 1 0 1264 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220370
transform 1 0 1112 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220370
transform 1 0 1080 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220370
transform 1 0 920 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220370
transform 1 0 1232 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220370
transform 1 0 1384 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220370
transform 1 0 1544 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220370
transform 1 0 1472 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220370
transform 1 0 1296 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220370
transform 1 0 1120 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220370
transform 1 0 952 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220370
transform 1 0 1680 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220370
transform 1 0 1448 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220370
transform 1 0 1224 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220370
transform 1 0 1024 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220370
transform 1 0 848 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220370
transform 1 0 1400 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220370
transform 1 0 1240 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220370
transform 1 0 1080 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220370
transform 1 0 936 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220370
transform 1 0 1304 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220370
transform 1 0 1176 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220370
transform 1 0 1048 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220370
transform 1 0 928 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220370
transform 1 0 808 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220370
transform 1 0 704 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220370
transform 1 0 608 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220370
transform 1 0 512 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220370
transform 1 0 416 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220370
transform 1 0 800 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220370
transform 1 0 688 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220370
transform 1 0 592 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220370
transform 1 0 496 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220370
transform 1 0 400 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220370
transform 1 0 304 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220370
transform 1 0 696 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220370
transform 1 0 560 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220370
transform 1 0 424 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220370
transform 1 0 288 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220370
transform 1 0 784 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220370
transform 1 0 616 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220370
transform 1 0 448 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220370
transform 1 0 288 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220370
transform 1 0 136 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220370
transform 1 0 760 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220370
transform 1 0 592 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220370
transform 1 0 424 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220370
transform 1 0 256 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220370
transform 1 0 128 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220370
transform 1 0 128 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220370
transform 1 0 240 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220370
transform 1 0 664 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220370
transform 1 0 520 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220370
transform 1 0 376 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220370
transform 1 0 280 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220370
transform 1 0 152 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220370
transform 1 0 688 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220370
transform 1 0 552 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220370
transform 1 0 416 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220370
transform 1 0 408 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220370
transform 1 0 264 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220370
transform 1 0 888 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220370
transform 1 0 728 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220370
transform 1 0 568 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220370
transform 1 0 512 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220370
transform 1 0 360 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220370
transform 1 0 672 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220370
transform 1 0 840 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220370
transform 1 0 1008 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220370
transform 1 0 1120 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220370
transform 1 0 928 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220370
transform 1 0 744 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220370
transform 1 0 560 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220370
transform 1 0 392 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220370
transform 1 0 880 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220370
transform 1 0 720 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220370
transform 1 0 560 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220370
transform 1 0 408 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220370
transform 1 0 808 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220370
transform 1 0 680 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220370
transform 1 0 544 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220370
transform 1 0 416 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220370
transform 1 0 296 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220370
transform 1 0 968 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220370
transform 1 0 784 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220370
transform 1 0 600 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220370
transform 1 0 424 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220370
transform 1 0 272 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220370
transform 1 0 144 0 1 3932
box 8 5 92 72
<< end >>
