magic
tech sky130l
timestamp 1731220636
<< m2 >>
rect 1534 2508 1540 2509
rect 1534 2504 1535 2508
rect 1539 2504 1540 2508
rect 1534 2503 1540 2504
rect 1574 2508 1580 2509
rect 1574 2504 1575 2508
rect 1579 2504 1580 2508
rect 1574 2503 1580 2504
rect 1614 2508 1620 2509
rect 1614 2504 1615 2508
rect 1619 2504 1620 2508
rect 1614 2503 1620 2504
rect 1654 2508 1660 2509
rect 1654 2504 1655 2508
rect 1659 2504 1660 2508
rect 1654 2503 1660 2504
rect 1694 2508 1700 2509
rect 1694 2504 1695 2508
rect 1699 2504 1700 2508
rect 1694 2503 1700 2504
rect 1734 2508 1740 2509
rect 1734 2504 1735 2508
rect 1739 2504 1740 2508
rect 1734 2503 1740 2504
rect 1774 2508 1780 2509
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1814 2503 1820 2504
rect 1854 2508 1860 2509
rect 1854 2504 1855 2508
rect 1859 2504 1860 2508
rect 1854 2503 1860 2504
rect 1894 2508 1900 2509
rect 1894 2504 1895 2508
rect 1899 2504 1900 2508
rect 1894 2503 1900 2504
rect 1934 2508 1940 2509
rect 1934 2504 1935 2508
rect 1939 2504 1940 2508
rect 1934 2503 1940 2504
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 1974 2503 1980 2504
rect 1278 2501 1284 2502
rect 1278 2497 1279 2501
rect 1283 2497 1284 2501
rect 1278 2496 1284 2497
rect 2406 2501 2412 2502
rect 2406 2497 2407 2501
rect 2411 2497 2412 2501
rect 2406 2496 2412 2497
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 174 2487 180 2488
rect 174 2483 175 2487
rect 179 2483 180 2487
rect 174 2482 180 2483
rect 214 2487 220 2488
rect 214 2483 215 2487
rect 219 2483 220 2487
rect 214 2482 220 2483
rect 254 2487 260 2488
rect 254 2483 255 2487
rect 259 2483 260 2487
rect 254 2482 260 2483
rect 310 2487 316 2488
rect 310 2483 311 2487
rect 315 2483 316 2487
rect 310 2482 316 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 478 2487 484 2488
rect 478 2483 479 2487
rect 483 2483 484 2487
rect 478 2482 484 2483
rect 566 2487 572 2488
rect 566 2483 567 2487
rect 571 2483 572 2487
rect 566 2482 572 2483
rect 654 2487 660 2488
rect 654 2483 655 2487
rect 659 2483 660 2487
rect 654 2482 660 2483
rect 742 2487 748 2488
rect 742 2483 743 2487
rect 747 2483 748 2487
rect 742 2482 748 2483
rect 830 2487 836 2488
rect 830 2483 831 2487
rect 835 2483 836 2487
rect 830 2482 836 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 1278 2484 1284 2485
rect 1278 2480 1279 2484
rect 1283 2480 1284 2484
rect 1278 2479 1284 2480
rect 2406 2484 2412 2485
rect 2406 2480 2407 2484
rect 2411 2480 2412 2484
rect 2406 2479 2412 2480
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 110 2459 116 2460
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 1534 2461 1540 2462
rect 1534 2457 1535 2461
rect 1539 2457 1540 2461
rect 1534 2456 1540 2457
rect 1574 2461 1580 2462
rect 1574 2457 1575 2461
rect 1579 2457 1580 2461
rect 1574 2456 1580 2457
rect 1614 2461 1620 2462
rect 1614 2457 1615 2461
rect 1619 2457 1620 2461
rect 1614 2456 1620 2457
rect 1654 2461 1660 2462
rect 1654 2457 1655 2461
rect 1659 2457 1660 2461
rect 1654 2456 1660 2457
rect 1694 2461 1700 2462
rect 1694 2457 1695 2461
rect 1699 2457 1700 2461
rect 1694 2456 1700 2457
rect 1734 2461 1740 2462
rect 1734 2457 1735 2461
rect 1739 2457 1740 2461
rect 1734 2456 1740 2457
rect 1774 2461 1780 2462
rect 1774 2457 1775 2461
rect 1779 2457 1780 2461
rect 1774 2456 1780 2457
rect 1814 2461 1820 2462
rect 1814 2457 1815 2461
rect 1819 2457 1820 2461
rect 1814 2456 1820 2457
rect 1854 2461 1860 2462
rect 1854 2457 1855 2461
rect 1859 2457 1860 2461
rect 1854 2456 1860 2457
rect 1894 2461 1900 2462
rect 1894 2457 1895 2461
rect 1899 2457 1900 2461
rect 1894 2456 1900 2457
rect 1934 2461 1940 2462
rect 1934 2457 1935 2461
rect 1939 2457 1940 2461
rect 1934 2456 1940 2457
rect 1974 2461 1980 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 110 2447 116 2448
rect 110 2443 111 2447
rect 115 2443 116 2447
rect 110 2442 116 2443
rect 1238 2447 1244 2448
rect 1238 2443 1239 2447
rect 1243 2443 1244 2447
rect 1238 2442 1244 2443
rect 134 2440 140 2441
rect 134 2436 135 2440
rect 139 2436 140 2440
rect 134 2435 140 2436
rect 174 2440 180 2441
rect 174 2436 175 2440
rect 179 2436 180 2440
rect 174 2435 180 2436
rect 214 2440 220 2441
rect 214 2436 215 2440
rect 219 2436 220 2440
rect 214 2435 220 2436
rect 254 2440 260 2441
rect 254 2436 255 2440
rect 259 2436 260 2440
rect 254 2435 260 2436
rect 310 2440 316 2441
rect 310 2436 311 2440
rect 315 2436 316 2440
rect 310 2435 316 2436
rect 390 2440 396 2441
rect 390 2436 391 2440
rect 395 2436 396 2440
rect 390 2435 396 2436
rect 478 2440 484 2441
rect 478 2436 479 2440
rect 483 2436 484 2440
rect 478 2435 484 2436
rect 566 2440 572 2441
rect 566 2436 567 2440
rect 571 2436 572 2440
rect 566 2435 572 2436
rect 654 2440 660 2441
rect 654 2436 655 2440
rect 659 2436 660 2440
rect 654 2435 660 2436
rect 742 2440 748 2441
rect 742 2436 743 2440
rect 747 2436 748 2440
rect 742 2435 748 2436
rect 830 2440 836 2441
rect 830 2436 831 2440
rect 835 2436 836 2440
rect 830 2435 836 2436
rect 926 2440 932 2441
rect 926 2436 927 2440
rect 931 2436 932 2440
rect 926 2435 932 2436
rect 1358 2431 1364 2432
rect 134 2428 140 2429
rect 134 2424 135 2428
rect 139 2424 140 2428
rect 134 2423 140 2424
rect 182 2428 188 2429
rect 182 2424 183 2428
rect 187 2424 188 2428
rect 182 2423 188 2424
rect 246 2428 252 2429
rect 246 2424 247 2428
rect 251 2424 252 2428
rect 246 2423 252 2424
rect 318 2428 324 2429
rect 318 2424 319 2428
rect 323 2424 324 2428
rect 318 2423 324 2424
rect 390 2428 396 2429
rect 390 2424 391 2428
rect 395 2424 396 2428
rect 390 2423 396 2424
rect 470 2428 476 2429
rect 470 2424 471 2428
rect 475 2424 476 2428
rect 470 2423 476 2424
rect 542 2428 548 2429
rect 542 2424 543 2428
rect 547 2424 548 2428
rect 542 2423 548 2424
rect 614 2428 620 2429
rect 614 2424 615 2428
rect 619 2424 620 2428
rect 614 2423 620 2424
rect 678 2428 684 2429
rect 678 2424 679 2428
rect 683 2424 684 2428
rect 678 2423 684 2424
rect 734 2428 740 2429
rect 734 2424 735 2428
rect 739 2424 740 2428
rect 734 2423 740 2424
rect 790 2428 796 2429
rect 790 2424 791 2428
rect 795 2424 796 2428
rect 790 2423 796 2424
rect 838 2428 844 2429
rect 838 2424 839 2428
rect 843 2424 844 2428
rect 838 2423 844 2424
rect 886 2428 892 2429
rect 886 2424 887 2428
rect 891 2424 892 2428
rect 886 2423 892 2424
rect 934 2428 940 2429
rect 934 2424 935 2428
rect 939 2424 940 2428
rect 934 2423 940 2424
rect 990 2428 996 2429
rect 990 2424 991 2428
rect 995 2424 996 2428
rect 990 2423 996 2424
rect 1046 2428 1052 2429
rect 1046 2424 1047 2428
rect 1051 2424 1052 2428
rect 1358 2427 1359 2431
rect 1363 2427 1364 2431
rect 1358 2426 1364 2427
rect 1398 2431 1404 2432
rect 1398 2427 1399 2431
rect 1403 2427 1404 2431
rect 1398 2426 1404 2427
rect 1454 2431 1460 2432
rect 1454 2427 1455 2431
rect 1459 2427 1460 2431
rect 1454 2426 1460 2427
rect 1518 2431 1524 2432
rect 1518 2427 1519 2431
rect 1523 2427 1524 2431
rect 1518 2426 1524 2427
rect 1598 2431 1604 2432
rect 1598 2427 1599 2431
rect 1603 2427 1604 2431
rect 1598 2426 1604 2427
rect 1678 2431 1684 2432
rect 1678 2427 1679 2431
rect 1683 2427 1684 2431
rect 1678 2426 1684 2427
rect 1758 2431 1764 2432
rect 1758 2427 1759 2431
rect 1763 2427 1764 2431
rect 1758 2426 1764 2427
rect 1838 2431 1844 2432
rect 1838 2427 1839 2431
rect 1843 2427 1844 2431
rect 1838 2426 1844 2427
rect 1918 2431 1924 2432
rect 1918 2427 1919 2431
rect 1923 2427 1924 2431
rect 1918 2426 1924 2427
rect 1998 2431 2004 2432
rect 1998 2427 1999 2431
rect 2003 2427 2004 2431
rect 1998 2426 2004 2427
rect 2078 2431 2084 2432
rect 2078 2427 2079 2431
rect 2083 2427 2084 2431
rect 2078 2426 2084 2427
rect 2158 2431 2164 2432
rect 2158 2427 2159 2431
rect 2163 2427 2164 2431
rect 2158 2426 2164 2427
rect 2246 2431 2252 2432
rect 2246 2427 2247 2431
rect 2251 2427 2252 2431
rect 2246 2426 2252 2427
rect 2334 2431 2340 2432
rect 2334 2427 2335 2431
rect 2339 2427 2340 2431
rect 2334 2426 2340 2427
rect 1046 2423 1052 2424
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 110 2416 116 2417
rect 1238 2421 1244 2422
rect 1238 2417 1239 2421
rect 1243 2417 1244 2421
rect 1238 2416 1244 2417
rect 1278 2408 1284 2409
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 110 2399 116 2400
rect 1238 2404 1244 2405
rect 1238 2400 1239 2404
rect 1243 2400 1244 2404
rect 1278 2404 1279 2408
rect 1283 2404 1284 2408
rect 1278 2403 1284 2404
rect 2406 2408 2412 2409
rect 2406 2404 2407 2408
rect 2411 2404 2412 2408
rect 2406 2403 2412 2404
rect 1238 2399 1244 2400
rect 1278 2391 1284 2392
rect 1278 2387 1279 2391
rect 1283 2387 1284 2391
rect 1278 2386 1284 2387
rect 2406 2391 2412 2392
rect 2406 2387 2407 2391
rect 2411 2387 2412 2391
rect 2406 2386 2412 2387
rect 1358 2384 1364 2385
rect 134 2381 140 2382
rect 134 2377 135 2381
rect 139 2377 140 2381
rect 134 2376 140 2377
rect 182 2381 188 2382
rect 182 2377 183 2381
rect 187 2377 188 2381
rect 182 2376 188 2377
rect 246 2381 252 2382
rect 246 2377 247 2381
rect 251 2377 252 2381
rect 246 2376 252 2377
rect 318 2381 324 2382
rect 318 2377 319 2381
rect 323 2377 324 2381
rect 318 2376 324 2377
rect 390 2381 396 2382
rect 390 2377 391 2381
rect 395 2377 396 2381
rect 390 2376 396 2377
rect 470 2381 476 2382
rect 470 2377 471 2381
rect 475 2377 476 2381
rect 470 2376 476 2377
rect 542 2381 548 2382
rect 542 2377 543 2381
rect 547 2377 548 2381
rect 542 2376 548 2377
rect 614 2381 620 2382
rect 614 2377 615 2381
rect 619 2377 620 2381
rect 614 2376 620 2377
rect 678 2381 684 2382
rect 678 2377 679 2381
rect 683 2377 684 2381
rect 678 2376 684 2377
rect 734 2381 740 2382
rect 734 2377 735 2381
rect 739 2377 740 2381
rect 734 2376 740 2377
rect 790 2381 796 2382
rect 790 2377 791 2381
rect 795 2377 796 2381
rect 790 2376 796 2377
rect 838 2381 844 2382
rect 838 2377 839 2381
rect 843 2377 844 2381
rect 838 2376 844 2377
rect 886 2381 892 2382
rect 886 2377 887 2381
rect 891 2377 892 2381
rect 886 2376 892 2377
rect 934 2381 940 2382
rect 934 2377 935 2381
rect 939 2377 940 2381
rect 934 2376 940 2377
rect 990 2381 996 2382
rect 990 2377 991 2381
rect 995 2377 996 2381
rect 990 2376 996 2377
rect 1046 2381 1052 2382
rect 1046 2377 1047 2381
rect 1051 2377 1052 2381
rect 1358 2380 1359 2384
rect 1363 2380 1364 2384
rect 1358 2379 1364 2380
rect 1398 2384 1404 2385
rect 1398 2380 1399 2384
rect 1403 2380 1404 2384
rect 1398 2379 1404 2380
rect 1454 2384 1460 2385
rect 1454 2380 1455 2384
rect 1459 2380 1460 2384
rect 1454 2379 1460 2380
rect 1518 2384 1524 2385
rect 1518 2380 1519 2384
rect 1523 2380 1524 2384
rect 1518 2379 1524 2380
rect 1598 2384 1604 2385
rect 1598 2380 1599 2384
rect 1603 2380 1604 2384
rect 1598 2379 1604 2380
rect 1678 2384 1684 2385
rect 1678 2380 1679 2384
rect 1683 2380 1684 2384
rect 1678 2379 1684 2380
rect 1758 2384 1764 2385
rect 1758 2380 1759 2384
rect 1763 2380 1764 2384
rect 1758 2379 1764 2380
rect 1838 2384 1844 2385
rect 1838 2380 1839 2384
rect 1843 2380 1844 2384
rect 1838 2379 1844 2380
rect 1918 2384 1924 2385
rect 1918 2380 1919 2384
rect 1923 2380 1924 2384
rect 1918 2379 1924 2380
rect 1998 2384 2004 2385
rect 1998 2380 1999 2384
rect 2003 2380 2004 2384
rect 1998 2379 2004 2380
rect 2078 2384 2084 2385
rect 2078 2380 2079 2384
rect 2083 2380 2084 2384
rect 2078 2379 2084 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2246 2384 2252 2385
rect 2246 2380 2247 2384
rect 2251 2380 2252 2384
rect 2246 2379 2252 2380
rect 2334 2384 2340 2385
rect 2334 2380 2335 2384
rect 2339 2380 2340 2384
rect 2334 2379 2340 2380
rect 1046 2376 1052 2377
rect 1358 2372 1364 2373
rect 1358 2368 1359 2372
rect 1363 2368 1364 2372
rect 1358 2367 1364 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1470 2372 1476 2373
rect 1470 2368 1471 2372
rect 1475 2368 1476 2372
rect 1470 2367 1476 2368
rect 1542 2372 1548 2373
rect 1542 2368 1543 2372
rect 1547 2368 1548 2372
rect 1542 2367 1548 2368
rect 1614 2372 1620 2373
rect 1614 2368 1615 2372
rect 1619 2368 1620 2372
rect 1614 2367 1620 2368
rect 1694 2372 1700 2373
rect 1694 2368 1695 2372
rect 1699 2368 1700 2372
rect 1694 2367 1700 2368
rect 1774 2372 1780 2373
rect 1774 2368 1775 2372
rect 1779 2368 1780 2372
rect 1774 2367 1780 2368
rect 1854 2372 1860 2373
rect 1854 2368 1855 2372
rect 1859 2368 1860 2372
rect 1854 2367 1860 2368
rect 1926 2372 1932 2373
rect 1926 2368 1927 2372
rect 1931 2368 1932 2372
rect 1926 2367 1932 2368
rect 1998 2372 2004 2373
rect 1998 2368 1999 2372
rect 2003 2368 2004 2372
rect 1998 2367 2004 2368
rect 2070 2372 2076 2373
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 2142 2372 2148 2373
rect 2142 2368 2143 2372
rect 2147 2368 2148 2372
rect 2142 2367 2148 2368
rect 2222 2372 2228 2373
rect 2222 2368 2223 2372
rect 2227 2368 2228 2372
rect 2222 2367 2228 2368
rect 2302 2372 2308 2373
rect 2302 2368 2303 2372
rect 2307 2368 2308 2372
rect 2302 2367 2308 2368
rect 2358 2372 2364 2373
rect 2358 2368 2359 2372
rect 2363 2368 2364 2372
rect 2358 2367 2364 2368
rect 1278 2365 1284 2366
rect 1278 2361 1279 2365
rect 1283 2361 1284 2365
rect 1278 2360 1284 2361
rect 2406 2365 2412 2366
rect 2406 2361 2407 2365
rect 2411 2361 2412 2365
rect 2406 2360 2412 2361
rect 1278 2348 1284 2349
rect 1278 2344 1279 2348
rect 1283 2344 1284 2348
rect 134 2343 140 2344
rect 134 2339 135 2343
rect 139 2339 140 2343
rect 134 2338 140 2339
rect 174 2343 180 2344
rect 174 2339 175 2343
rect 179 2339 180 2343
rect 174 2338 180 2339
rect 214 2343 220 2344
rect 214 2339 215 2343
rect 219 2339 220 2343
rect 214 2338 220 2339
rect 270 2343 276 2344
rect 270 2339 271 2343
rect 275 2339 276 2343
rect 270 2338 276 2339
rect 350 2343 356 2344
rect 350 2339 351 2343
rect 355 2339 356 2343
rect 350 2338 356 2339
rect 430 2343 436 2344
rect 430 2339 431 2343
rect 435 2339 436 2343
rect 430 2338 436 2339
rect 518 2343 524 2344
rect 518 2339 519 2343
rect 523 2339 524 2343
rect 518 2338 524 2339
rect 598 2343 604 2344
rect 598 2339 599 2343
rect 603 2339 604 2343
rect 598 2338 604 2339
rect 678 2343 684 2344
rect 678 2339 679 2343
rect 683 2339 684 2343
rect 678 2338 684 2339
rect 750 2343 756 2344
rect 750 2339 751 2343
rect 755 2339 756 2343
rect 750 2338 756 2339
rect 822 2343 828 2344
rect 822 2339 823 2343
rect 827 2339 828 2343
rect 822 2338 828 2339
rect 886 2343 892 2344
rect 886 2339 887 2343
rect 891 2339 892 2343
rect 886 2338 892 2339
rect 958 2343 964 2344
rect 958 2339 959 2343
rect 963 2339 964 2343
rect 958 2338 964 2339
rect 1030 2343 1036 2344
rect 1278 2343 1284 2344
rect 2406 2348 2412 2349
rect 2406 2344 2407 2348
rect 2411 2344 2412 2348
rect 2406 2343 2412 2344
rect 1030 2339 1031 2343
rect 1035 2339 1036 2343
rect 1030 2338 1036 2339
rect 1358 2325 1364 2326
rect 1358 2321 1359 2325
rect 1363 2321 1364 2325
rect 110 2320 116 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 1238 2320 1244 2321
rect 1358 2320 1364 2321
rect 1406 2325 1412 2326
rect 1406 2321 1407 2325
rect 1411 2321 1412 2325
rect 1406 2320 1412 2321
rect 1470 2325 1476 2326
rect 1470 2321 1471 2325
rect 1475 2321 1476 2325
rect 1470 2320 1476 2321
rect 1542 2325 1548 2326
rect 1542 2321 1543 2325
rect 1547 2321 1548 2325
rect 1542 2320 1548 2321
rect 1614 2325 1620 2326
rect 1614 2321 1615 2325
rect 1619 2321 1620 2325
rect 1614 2320 1620 2321
rect 1694 2325 1700 2326
rect 1694 2321 1695 2325
rect 1699 2321 1700 2325
rect 1694 2320 1700 2321
rect 1774 2325 1780 2326
rect 1774 2321 1775 2325
rect 1779 2321 1780 2325
rect 1774 2320 1780 2321
rect 1854 2325 1860 2326
rect 1854 2321 1855 2325
rect 1859 2321 1860 2325
rect 1854 2320 1860 2321
rect 1926 2325 1932 2326
rect 1926 2321 1927 2325
rect 1931 2321 1932 2325
rect 1926 2320 1932 2321
rect 1998 2325 2004 2326
rect 1998 2321 1999 2325
rect 2003 2321 2004 2325
rect 1998 2320 2004 2321
rect 2070 2325 2076 2326
rect 2070 2321 2071 2325
rect 2075 2321 2076 2325
rect 2070 2320 2076 2321
rect 2142 2325 2148 2326
rect 2142 2321 2143 2325
rect 2147 2321 2148 2325
rect 2142 2320 2148 2321
rect 2222 2325 2228 2326
rect 2222 2321 2223 2325
rect 2227 2321 2228 2325
rect 2222 2320 2228 2321
rect 2302 2325 2308 2326
rect 2302 2321 2303 2325
rect 2307 2321 2308 2325
rect 2302 2320 2308 2321
rect 2358 2325 2364 2326
rect 2358 2321 2359 2325
rect 2363 2321 2364 2325
rect 2358 2320 2364 2321
rect 1238 2316 1239 2320
rect 1243 2316 1244 2320
rect 1238 2315 1244 2316
rect 110 2303 116 2304
rect 110 2299 111 2303
rect 115 2299 116 2303
rect 110 2298 116 2299
rect 1238 2303 1244 2304
rect 1238 2299 1239 2303
rect 1243 2299 1244 2303
rect 1238 2298 1244 2299
rect 134 2296 140 2297
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 174 2296 180 2297
rect 174 2292 175 2296
rect 179 2292 180 2296
rect 174 2291 180 2292
rect 214 2296 220 2297
rect 214 2292 215 2296
rect 219 2292 220 2296
rect 214 2291 220 2292
rect 270 2296 276 2297
rect 270 2292 271 2296
rect 275 2292 276 2296
rect 270 2291 276 2292
rect 350 2296 356 2297
rect 350 2292 351 2296
rect 355 2292 356 2296
rect 350 2291 356 2292
rect 430 2296 436 2297
rect 430 2292 431 2296
rect 435 2292 436 2296
rect 430 2291 436 2292
rect 518 2296 524 2297
rect 518 2292 519 2296
rect 523 2292 524 2296
rect 518 2291 524 2292
rect 598 2296 604 2297
rect 598 2292 599 2296
rect 603 2292 604 2296
rect 598 2291 604 2292
rect 678 2296 684 2297
rect 678 2292 679 2296
rect 683 2292 684 2296
rect 678 2291 684 2292
rect 750 2296 756 2297
rect 750 2292 751 2296
rect 755 2292 756 2296
rect 750 2291 756 2292
rect 822 2296 828 2297
rect 822 2292 823 2296
rect 827 2292 828 2296
rect 822 2291 828 2292
rect 886 2296 892 2297
rect 886 2292 887 2296
rect 891 2292 892 2296
rect 886 2291 892 2292
rect 958 2296 964 2297
rect 958 2292 959 2296
rect 963 2292 964 2296
rect 958 2291 964 2292
rect 1030 2296 1036 2297
rect 1030 2292 1031 2296
rect 1035 2292 1036 2296
rect 1030 2291 1036 2292
rect 1502 2291 1508 2292
rect 1502 2287 1503 2291
rect 1507 2287 1508 2291
rect 1502 2286 1508 2287
rect 1542 2291 1548 2292
rect 1542 2287 1543 2291
rect 1547 2287 1548 2291
rect 1542 2286 1548 2287
rect 1582 2291 1588 2292
rect 1582 2287 1583 2291
rect 1587 2287 1588 2291
rect 1582 2286 1588 2287
rect 1622 2291 1628 2292
rect 1622 2287 1623 2291
rect 1627 2287 1628 2291
rect 1622 2286 1628 2287
rect 1662 2291 1668 2292
rect 1662 2287 1663 2291
rect 1667 2287 1668 2291
rect 1662 2286 1668 2287
rect 1702 2291 1708 2292
rect 1702 2287 1703 2291
rect 1707 2287 1708 2291
rect 1702 2286 1708 2287
rect 1758 2291 1764 2292
rect 1758 2287 1759 2291
rect 1763 2287 1764 2291
rect 1758 2286 1764 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1894 2291 1900 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1894 2286 1900 2287
rect 1966 2291 1972 2292
rect 1966 2287 1967 2291
rect 1971 2287 1972 2291
rect 1966 2286 1972 2287
rect 2046 2291 2052 2292
rect 2046 2287 2047 2291
rect 2051 2287 2052 2291
rect 2046 2286 2052 2287
rect 2126 2291 2132 2292
rect 2126 2287 2127 2291
rect 2131 2287 2132 2291
rect 2126 2286 2132 2287
rect 2206 2291 2212 2292
rect 2206 2287 2207 2291
rect 2211 2287 2212 2291
rect 2206 2286 2212 2287
rect 2294 2291 2300 2292
rect 2294 2287 2295 2291
rect 2299 2287 2300 2291
rect 2294 2286 2300 2287
rect 2358 2291 2364 2292
rect 2358 2287 2359 2291
rect 2363 2287 2364 2291
rect 2358 2286 2364 2287
rect 134 2280 140 2281
rect 134 2276 135 2280
rect 139 2276 140 2280
rect 134 2275 140 2276
rect 174 2280 180 2281
rect 174 2276 175 2280
rect 179 2276 180 2280
rect 174 2275 180 2276
rect 230 2280 236 2281
rect 230 2276 231 2280
rect 235 2276 236 2280
rect 230 2275 236 2276
rect 302 2280 308 2281
rect 302 2276 303 2280
rect 307 2276 308 2280
rect 302 2275 308 2276
rect 374 2280 380 2281
rect 374 2276 375 2280
rect 379 2276 380 2280
rect 374 2275 380 2276
rect 454 2280 460 2281
rect 454 2276 455 2280
rect 459 2276 460 2280
rect 454 2275 460 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 614 2280 620 2281
rect 614 2276 615 2280
rect 619 2276 620 2280
rect 614 2275 620 2276
rect 686 2280 692 2281
rect 686 2276 687 2280
rect 691 2276 692 2280
rect 686 2275 692 2276
rect 758 2280 764 2281
rect 758 2276 759 2280
rect 763 2276 764 2280
rect 758 2275 764 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 110 2268 116 2269
rect 1238 2273 1244 2274
rect 1238 2269 1239 2273
rect 1243 2269 1244 2273
rect 1238 2268 1244 2269
rect 1278 2268 1284 2269
rect 1278 2264 1279 2268
rect 1283 2264 1284 2268
rect 1278 2263 1284 2264
rect 2406 2268 2412 2269
rect 2406 2264 2407 2268
rect 2411 2264 2412 2268
rect 2406 2263 2412 2264
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 110 2251 116 2252
rect 1238 2256 1244 2257
rect 1238 2252 1239 2256
rect 1243 2252 1244 2256
rect 1238 2251 1244 2252
rect 1278 2251 1284 2252
rect 1278 2247 1279 2251
rect 1283 2247 1284 2251
rect 1278 2246 1284 2247
rect 2406 2251 2412 2252
rect 2406 2247 2407 2251
rect 2411 2247 2412 2251
rect 2406 2246 2412 2247
rect 1502 2244 1508 2245
rect 1502 2240 1503 2244
rect 1507 2240 1508 2244
rect 1502 2239 1508 2240
rect 1542 2244 1548 2245
rect 1542 2240 1543 2244
rect 1547 2240 1548 2244
rect 1542 2239 1548 2240
rect 1582 2244 1588 2245
rect 1582 2240 1583 2244
rect 1587 2240 1588 2244
rect 1582 2239 1588 2240
rect 1622 2244 1628 2245
rect 1622 2240 1623 2244
rect 1627 2240 1628 2244
rect 1622 2239 1628 2240
rect 1662 2244 1668 2245
rect 1662 2240 1663 2244
rect 1667 2240 1668 2244
rect 1662 2239 1668 2240
rect 1702 2244 1708 2245
rect 1702 2240 1703 2244
rect 1707 2240 1708 2244
rect 1702 2239 1708 2240
rect 1758 2244 1764 2245
rect 1758 2240 1759 2244
rect 1763 2240 1764 2244
rect 1758 2239 1764 2240
rect 1822 2244 1828 2245
rect 1822 2240 1823 2244
rect 1827 2240 1828 2244
rect 1822 2239 1828 2240
rect 1894 2244 1900 2245
rect 1894 2240 1895 2244
rect 1899 2240 1900 2244
rect 1894 2239 1900 2240
rect 1966 2244 1972 2245
rect 1966 2240 1967 2244
rect 1971 2240 1972 2244
rect 1966 2239 1972 2240
rect 2046 2244 2052 2245
rect 2046 2240 2047 2244
rect 2051 2240 2052 2244
rect 2046 2239 2052 2240
rect 2126 2244 2132 2245
rect 2126 2240 2127 2244
rect 2131 2240 2132 2244
rect 2126 2239 2132 2240
rect 2206 2244 2212 2245
rect 2206 2240 2207 2244
rect 2211 2240 2212 2244
rect 2206 2239 2212 2240
rect 2294 2244 2300 2245
rect 2294 2240 2295 2244
rect 2299 2240 2300 2244
rect 2294 2239 2300 2240
rect 2358 2244 2364 2245
rect 2358 2240 2359 2244
rect 2363 2240 2364 2244
rect 2358 2239 2364 2240
rect 134 2233 140 2234
rect 134 2229 135 2233
rect 139 2229 140 2233
rect 134 2228 140 2229
rect 174 2233 180 2234
rect 174 2229 175 2233
rect 179 2229 180 2233
rect 174 2228 180 2229
rect 230 2233 236 2234
rect 230 2229 231 2233
rect 235 2229 236 2233
rect 230 2228 236 2229
rect 302 2233 308 2234
rect 302 2229 303 2233
rect 307 2229 308 2233
rect 302 2228 308 2229
rect 374 2233 380 2234
rect 374 2229 375 2233
rect 379 2229 380 2233
rect 374 2228 380 2229
rect 454 2233 460 2234
rect 454 2229 455 2233
rect 459 2229 460 2233
rect 454 2228 460 2229
rect 534 2233 540 2234
rect 534 2229 535 2233
rect 539 2229 540 2233
rect 534 2228 540 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 686 2233 692 2234
rect 686 2229 687 2233
rect 691 2229 692 2233
rect 686 2228 692 2229
rect 758 2233 764 2234
rect 758 2229 759 2233
rect 763 2229 764 2233
rect 758 2228 764 2229
rect 830 2233 836 2234
rect 830 2229 831 2233
rect 835 2229 836 2233
rect 830 2228 836 2229
rect 910 2233 916 2234
rect 910 2229 911 2233
rect 915 2229 916 2233
rect 910 2228 916 2229
rect 990 2233 996 2234
rect 990 2229 991 2233
rect 995 2229 996 2233
rect 990 2228 996 2229
rect 1302 2224 1308 2225
rect 1302 2220 1303 2224
rect 1307 2220 1308 2224
rect 1302 2219 1308 2220
rect 1342 2224 1348 2225
rect 1342 2220 1343 2224
rect 1347 2220 1348 2224
rect 1342 2219 1348 2220
rect 1382 2224 1388 2225
rect 1382 2220 1383 2224
rect 1387 2220 1388 2224
rect 1382 2219 1388 2220
rect 1430 2224 1436 2225
rect 1430 2220 1431 2224
rect 1435 2220 1436 2224
rect 1430 2219 1436 2220
rect 1494 2224 1500 2225
rect 1494 2220 1495 2224
rect 1499 2220 1500 2224
rect 1494 2219 1500 2220
rect 1566 2224 1572 2225
rect 1566 2220 1567 2224
rect 1571 2220 1572 2224
rect 1566 2219 1572 2220
rect 1638 2224 1644 2225
rect 1638 2220 1639 2224
rect 1643 2220 1644 2224
rect 1638 2219 1644 2220
rect 1710 2224 1716 2225
rect 1710 2220 1711 2224
rect 1715 2220 1716 2224
rect 1710 2219 1716 2220
rect 1782 2224 1788 2225
rect 1782 2220 1783 2224
rect 1787 2220 1788 2224
rect 1782 2219 1788 2220
rect 1854 2224 1860 2225
rect 1854 2220 1855 2224
rect 1859 2220 1860 2224
rect 1854 2219 1860 2220
rect 1934 2224 1940 2225
rect 1934 2220 1935 2224
rect 1939 2220 1940 2224
rect 1934 2219 1940 2220
rect 2014 2224 2020 2225
rect 2014 2220 2015 2224
rect 2019 2220 2020 2224
rect 2014 2219 2020 2220
rect 2094 2224 2100 2225
rect 2094 2220 2095 2224
rect 2099 2220 2100 2224
rect 2094 2219 2100 2220
rect 2182 2224 2188 2225
rect 2182 2220 2183 2224
rect 2187 2220 2188 2224
rect 2182 2219 2188 2220
rect 2278 2224 2284 2225
rect 2278 2220 2279 2224
rect 2283 2220 2284 2224
rect 2278 2219 2284 2220
rect 2358 2224 2364 2225
rect 2358 2220 2359 2224
rect 2363 2220 2364 2224
rect 2358 2219 2364 2220
rect 1278 2217 1284 2218
rect 1278 2213 1279 2217
rect 1283 2213 1284 2217
rect 1278 2212 1284 2213
rect 2406 2217 2412 2218
rect 2406 2213 2407 2217
rect 2411 2213 2412 2217
rect 2406 2212 2412 2213
rect 246 2203 252 2204
rect 246 2199 247 2203
rect 251 2199 252 2203
rect 246 2198 252 2199
rect 286 2203 292 2204
rect 286 2199 287 2203
rect 291 2199 292 2203
rect 286 2198 292 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 374 2203 380 2204
rect 374 2199 375 2203
rect 379 2199 380 2203
rect 374 2198 380 2199
rect 430 2203 436 2204
rect 430 2199 431 2203
rect 435 2199 436 2203
rect 430 2198 436 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 550 2203 556 2204
rect 550 2199 551 2203
rect 555 2199 556 2203
rect 550 2198 556 2199
rect 606 2203 612 2204
rect 606 2199 607 2203
rect 611 2199 612 2203
rect 606 2198 612 2199
rect 662 2203 668 2204
rect 662 2199 663 2203
rect 667 2199 668 2203
rect 662 2198 668 2199
rect 718 2203 724 2204
rect 718 2199 719 2203
rect 723 2199 724 2203
rect 718 2198 724 2199
rect 782 2203 788 2204
rect 782 2199 783 2203
rect 787 2199 788 2203
rect 782 2198 788 2199
rect 846 2203 852 2204
rect 846 2199 847 2203
rect 851 2199 852 2203
rect 846 2198 852 2199
rect 910 2203 916 2204
rect 910 2199 911 2203
rect 915 2199 916 2203
rect 910 2198 916 2199
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 2406 2200 2412 2201
rect 2406 2196 2407 2200
rect 2411 2196 2412 2200
rect 2406 2195 2412 2196
rect 110 2180 116 2181
rect 110 2176 111 2180
rect 115 2176 116 2180
rect 110 2175 116 2176
rect 1238 2180 1244 2181
rect 1238 2176 1239 2180
rect 1243 2176 1244 2180
rect 1238 2175 1244 2176
rect 1302 2177 1308 2178
rect 1302 2173 1303 2177
rect 1307 2173 1308 2177
rect 1302 2172 1308 2173
rect 1342 2177 1348 2178
rect 1342 2173 1343 2177
rect 1347 2173 1348 2177
rect 1342 2172 1348 2173
rect 1382 2177 1388 2178
rect 1382 2173 1383 2177
rect 1387 2173 1388 2177
rect 1382 2172 1388 2173
rect 1430 2177 1436 2178
rect 1430 2173 1431 2177
rect 1435 2173 1436 2177
rect 1430 2172 1436 2173
rect 1494 2177 1500 2178
rect 1494 2173 1495 2177
rect 1499 2173 1500 2177
rect 1494 2172 1500 2173
rect 1566 2177 1572 2178
rect 1566 2173 1567 2177
rect 1571 2173 1572 2177
rect 1566 2172 1572 2173
rect 1638 2177 1644 2178
rect 1638 2173 1639 2177
rect 1643 2173 1644 2177
rect 1638 2172 1644 2173
rect 1710 2177 1716 2178
rect 1710 2173 1711 2177
rect 1715 2173 1716 2177
rect 1710 2172 1716 2173
rect 1782 2177 1788 2178
rect 1782 2173 1783 2177
rect 1787 2173 1788 2177
rect 1782 2172 1788 2173
rect 1854 2177 1860 2178
rect 1854 2173 1855 2177
rect 1859 2173 1860 2177
rect 1854 2172 1860 2173
rect 1934 2177 1940 2178
rect 1934 2173 1935 2177
rect 1939 2173 1940 2177
rect 1934 2172 1940 2173
rect 2014 2177 2020 2178
rect 2014 2173 2015 2177
rect 2019 2173 2020 2177
rect 2014 2172 2020 2173
rect 2094 2177 2100 2178
rect 2094 2173 2095 2177
rect 2099 2173 2100 2177
rect 2094 2172 2100 2173
rect 2182 2177 2188 2178
rect 2182 2173 2183 2177
rect 2187 2173 2188 2177
rect 2182 2172 2188 2173
rect 2278 2177 2284 2178
rect 2278 2173 2279 2177
rect 2283 2173 2284 2177
rect 2278 2172 2284 2173
rect 2358 2177 2364 2178
rect 2358 2173 2359 2177
rect 2363 2173 2364 2177
rect 2358 2172 2364 2173
rect 110 2163 116 2164
rect 110 2159 111 2163
rect 115 2159 116 2163
rect 110 2158 116 2159
rect 1238 2163 1244 2164
rect 1238 2159 1239 2163
rect 1243 2159 1244 2163
rect 1238 2158 1244 2159
rect 246 2156 252 2157
rect 246 2152 247 2156
rect 251 2152 252 2156
rect 246 2151 252 2152
rect 286 2156 292 2157
rect 286 2152 287 2156
rect 291 2152 292 2156
rect 286 2151 292 2152
rect 326 2156 332 2157
rect 326 2152 327 2156
rect 331 2152 332 2156
rect 326 2151 332 2152
rect 374 2156 380 2157
rect 374 2152 375 2156
rect 379 2152 380 2156
rect 374 2151 380 2152
rect 430 2156 436 2157
rect 430 2152 431 2156
rect 435 2152 436 2156
rect 430 2151 436 2152
rect 494 2156 500 2157
rect 494 2152 495 2156
rect 499 2152 500 2156
rect 494 2151 500 2152
rect 550 2156 556 2157
rect 550 2152 551 2156
rect 555 2152 556 2156
rect 550 2151 556 2152
rect 606 2156 612 2157
rect 606 2152 607 2156
rect 611 2152 612 2156
rect 606 2151 612 2152
rect 662 2156 668 2157
rect 662 2152 663 2156
rect 667 2152 668 2156
rect 662 2151 668 2152
rect 718 2156 724 2157
rect 718 2152 719 2156
rect 723 2152 724 2156
rect 718 2151 724 2152
rect 782 2156 788 2157
rect 782 2152 783 2156
rect 787 2152 788 2156
rect 782 2151 788 2152
rect 846 2156 852 2157
rect 846 2152 847 2156
rect 851 2152 852 2156
rect 846 2151 852 2152
rect 910 2156 916 2157
rect 910 2152 911 2156
rect 915 2152 916 2156
rect 910 2151 916 2152
rect 1302 2147 1308 2148
rect 1302 2143 1303 2147
rect 1307 2143 1308 2147
rect 1302 2142 1308 2143
rect 1350 2147 1356 2148
rect 1350 2143 1351 2147
rect 1355 2143 1356 2147
rect 1350 2142 1356 2143
rect 1438 2147 1444 2148
rect 1438 2143 1439 2147
rect 1443 2143 1444 2147
rect 1438 2142 1444 2143
rect 1534 2147 1540 2148
rect 1534 2143 1535 2147
rect 1539 2143 1540 2147
rect 1534 2142 1540 2143
rect 1630 2147 1636 2148
rect 1630 2143 1631 2147
rect 1635 2143 1636 2147
rect 1630 2142 1636 2143
rect 1726 2147 1732 2148
rect 1726 2143 1727 2147
rect 1731 2143 1732 2147
rect 1726 2142 1732 2143
rect 1814 2147 1820 2148
rect 1814 2143 1815 2147
rect 1819 2143 1820 2147
rect 1814 2142 1820 2143
rect 1894 2147 1900 2148
rect 1894 2143 1895 2147
rect 1899 2143 1900 2147
rect 1894 2142 1900 2143
rect 1974 2147 1980 2148
rect 1974 2143 1975 2147
rect 1979 2143 1980 2147
rect 1974 2142 1980 2143
rect 2046 2147 2052 2148
rect 2046 2143 2047 2147
rect 2051 2143 2052 2147
rect 2046 2142 2052 2143
rect 2110 2147 2116 2148
rect 2110 2143 2111 2147
rect 2115 2143 2116 2147
rect 2110 2142 2116 2143
rect 2174 2147 2180 2148
rect 2174 2143 2175 2147
rect 2179 2143 2180 2147
rect 2174 2142 2180 2143
rect 2238 2147 2244 2148
rect 2238 2143 2239 2147
rect 2243 2143 2244 2147
rect 2238 2142 2244 2143
rect 2310 2147 2316 2148
rect 2310 2143 2311 2147
rect 2315 2143 2316 2147
rect 2310 2142 2316 2143
rect 2358 2147 2364 2148
rect 2358 2143 2359 2147
rect 2363 2143 2364 2147
rect 2358 2142 2364 2143
rect 382 2136 388 2137
rect 382 2132 383 2136
rect 387 2132 388 2136
rect 382 2131 388 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 462 2136 468 2137
rect 462 2132 463 2136
rect 467 2132 468 2136
rect 462 2131 468 2132
rect 502 2136 508 2137
rect 502 2132 503 2136
rect 507 2132 508 2136
rect 502 2131 508 2132
rect 550 2136 556 2137
rect 550 2132 551 2136
rect 555 2132 556 2136
rect 550 2131 556 2132
rect 606 2136 612 2137
rect 606 2132 607 2136
rect 611 2132 612 2136
rect 606 2131 612 2132
rect 662 2136 668 2137
rect 662 2132 663 2136
rect 667 2132 668 2136
rect 662 2131 668 2132
rect 726 2136 732 2137
rect 726 2132 727 2136
rect 731 2132 732 2136
rect 726 2131 732 2132
rect 790 2136 796 2137
rect 790 2132 791 2136
rect 795 2132 796 2136
rect 790 2131 796 2132
rect 854 2136 860 2137
rect 854 2132 855 2136
rect 859 2132 860 2136
rect 854 2131 860 2132
rect 910 2136 916 2137
rect 910 2132 911 2136
rect 915 2132 916 2136
rect 910 2131 916 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1022 2136 1028 2137
rect 1022 2132 1023 2136
rect 1027 2132 1028 2136
rect 1022 2131 1028 2132
rect 1078 2136 1084 2137
rect 1078 2132 1079 2136
rect 1083 2132 1084 2136
rect 1078 2131 1084 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 110 2129 116 2130
rect 110 2125 111 2129
rect 115 2125 116 2129
rect 110 2124 116 2125
rect 1238 2129 1244 2130
rect 1238 2125 1239 2129
rect 1243 2125 1244 2129
rect 1238 2124 1244 2125
rect 1278 2124 1284 2125
rect 1278 2120 1279 2124
rect 1283 2120 1284 2124
rect 1278 2119 1284 2120
rect 2406 2124 2412 2125
rect 2406 2120 2407 2124
rect 2411 2120 2412 2124
rect 2406 2119 2412 2120
rect 110 2112 116 2113
rect 110 2108 111 2112
rect 115 2108 116 2112
rect 110 2107 116 2108
rect 1238 2112 1244 2113
rect 1238 2108 1239 2112
rect 1243 2108 1244 2112
rect 1238 2107 1244 2108
rect 1278 2107 1284 2108
rect 1278 2103 1279 2107
rect 1283 2103 1284 2107
rect 1278 2102 1284 2103
rect 2406 2107 2412 2108
rect 2406 2103 2407 2107
rect 2411 2103 2412 2107
rect 2406 2102 2412 2103
rect 1302 2100 1308 2101
rect 1302 2096 1303 2100
rect 1307 2096 1308 2100
rect 1302 2095 1308 2096
rect 1350 2100 1356 2101
rect 1350 2096 1351 2100
rect 1355 2096 1356 2100
rect 1350 2095 1356 2096
rect 1438 2100 1444 2101
rect 1438 2096 1439 2100
rect 1443 2096 1444 2100
rect 1438 2095 1444 2096
rect 1534 2100 1540 2101
rect 1534 2096 1535 2100
rect 1539 2096 1540 2100
rect 1534 2095 1540 2096
rect 1630 2100 1636 2101
rect 1630 2096 1631 2100
rect 1635 2096 1636 2100
rect 1630 2095 1636 2096
rect 1726 2100 1732 2101
rect 1726 2096 1727 2100
rect 1731 2096 1732 2100
rect 1726 2095 1732 2096
rect 1814 2100 1820 2101
rect 1814 2096 1815 2100
rect 1819 2096 1820 2100
rect 1814 2095 1820 2096
rect 1894 2100 1900 2101
rect 1894 2096 1895 2100
rect 1899 2096 1900 2100
rect 1894 2095 1900 2096
rect 1974 2100 1980 2101
rect 1974 2096 1975 2100
rect 1979 2096 1980 2100
rect 1974 2095 1980 2096
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2046 2095 2052 2096
rect 2110 2100 2116 2101
rect 2110 2096 2111 2100
rect 2115 2096 2116 2100
rect 2110 2095 2116 2096
rect 2174 2100 2180 2101
rect 2174 2096 2175 2100
rect 2179 2096 2180 2100
rect 2174 2095 2180 2096
rect 2238 2100 2244 2101
rect 2238 2096 2239 2100
rect 2243 2096 2244 2100
rect 2238 2095 2244 2096
rect 2310 2100 2316 2101
rect 2310 2096 2311 2100
rect 2315 2096 2316 2100
rect 2310 2095 2316 2096
rect 2358 2100 2364 2101
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 382 2089 388 2090
rect 382 2085 383 2089
rect 387 2085 388 2089
rect 382 2084 388 2085
rect 422 2089 428 2090
rect 422 2085 423 2089
rect 427 2085 428 2089
rect 422 2084 428 2085
rect 462 2089 468 2090
rect 462 2085 463 2089
rect 467 2085 468 2089
rect 462 2084 468 2085
rect 502 2089 508 2090
rect 502 2085 503 2089
rect 507 2085 508 2089
rect 502 2084 508 2085
rect 550 2089 556 2090
rect 550 2085 551 2089
rect 555 2085 556 2089
rect 550 2084 556 2085
rect 606 2089 612 2090
rect 606 2085 607 2089
rect 611 2085 612 2089
rect 606 2084 612 2085
rect 662 2089 668 2090
rect 662 2085 663 2089
rect 667 2085 668 2089
rect 662 2084 668 2085
rect 726 2089 732 2090
rect 726 2085 727 2089
rect 731 2085 732 2089
rect 726 2084 732 2085
rect 790 2089 796 2090
rect 790 2085 791 2089
rect 795 2085 796 2089
rect 790 2084 796 2085
rect 854 2089 860 2090
rect 854 2085 855 2089
rect 859 2085 860 2089
rect 854 2084 860 2085
rect 910 2089 916 2090
rect 910 2085 911 2089
rect 915 2085 916 2089
rect 910 2084 916 2085
rect 966 2089 972 2090
rect 966 2085 967 2089
rect 971 2085 972 2089
rect 966 2084 972 2085
rect 1022 2089 1028 2090
rect 1022 2085 1023 2089
rect 1027 2085 1028 2089
rect 1022 2084 1028 2085
rect 1078 2089 1084 2090
rect 1078 2085 1079 2089
rect 1083 2085 1084 2089
rect 1078 2084 1084 2085
rect 1142 2089 1148 2090
rect 1142 2085 1143 2089
rect 1147 2085 1148 2089
rect 1142 2084 1148 2085
rect 1302 2084 1308 2085
rect 1302 2080 1303 2084
rect 1307 2080 1308 2084
rect 1302 2079 1308 2080
rect 1342 2084 1348 2085
rect 1342 2080 1343 2084
rect 1347 2080 1348 2084
rect 1342 2079 1348 2080
rect 1398 2084 1404 2085
rect 1398 2080 1399 2084
rect 1403 2080 1404 2084
rect 1398 2079 1404 2080
rect 1478 2084 1484 2085
rect 1478 2080 1479 2084
rect 1483 2080 1484 2084
rect 1478 2079 1484 2080
rect 1566 2084 1572 2085
rect 1566 2080 1567 2084
rect 1571 2080 1572 2084
rect 1566 2079 1572 2080
rect 1662 2084 1668 2085
rect 1662 2080 1663 2084
rect 1667 2080 1668 2084
rect 1662 2079 1668 2080
rect 1758 2084 1764 2085
rect 1758 2080 1759 2084
rect 1763 2080 1764 2084
rect 1758 2079 1764 2080
rect 1846 2084 1852 2085
rect 1846 2080 1847 2084
rect 1851 2080 1852 2084
rect 1846 2079 1852 2080
rect 1934 2084 1940 2085
rect 1934 2080 1935 2084
rect 1939 2080 1940 2084
rect 1934 2079 1940 2080
rect 2014 2084 2020 2085
rect 2014 2080 2015 2084
rect 2019 2080 2020 2084
rect 2014 2079 2020 2080
rect 2094 2084 2100 2085
rect 2094 2080 2095 2084
rect 2099 2080 2100 2084
rect 2094 2079 2100 2080
rect 2166 2084 2172 2085
rect 2166 2080 2167 2084
rect 2171 2080 2172 2084
rect 2166 2079 2172 2080
rect 2238 2084 2244 2085
rect 2238 2080 2239 2084
rect 2243 2080 2244 2084
rect 2238 2079 2244 2080
rect 2310 2084 2316 2085
rect 2310 2080 2311 2084
rect 2315 2080 2316 2084
rect 2310 2079 2316 2080
rect 2358 2084 2364 2085
rect 2358 2080 2359 2084
rect 2363 2080 2364 2084
rect 2358 2079 2364 2080
rect 1278 2077 1284 2078
rect 1278 2073 1279 2077
rect 1283 2073 1284 2077
rect 1278 2072 1284 2073
rect 2406 2077 2412 2078
rect 2406 2073 2407 2077
rect 2411 2073 2412 2077
rect 2406 2072 2412 2073
rect 1278 2060 1284 2061
rect 382 2059 388 2060
rect 382 2055 383 2059
rect 387 2055 388 2059
rect 382 2054 388 2055
rect 422 2059 428 2060
rect 422 2055 423 2059
rect 427 2055 428 2059
rect 422 2054 428 2055
rect 462 2059 468 2060
rect 462 2055 463 2059
rect 467 2055 468 2059
rect 462 2054 468 2055
rect 502 2059 508 2060
rect 502 2055 503 2059
rect 507 2055 508 2059
rect 502 2054 508 2055
rect 542 2059 548 2060
rect 542 2055 543 2059
rect 547 2055 548 2059
rect 542 2054 548 2055
rect 582 2059 588 2060
rect 582 2055 583 2059
rect 587 2055 588 2059
rect 582 2054 588 2055
rect 630 2059 636 2060
rect 630 2055 631 2059
rect 635 2055 636 2059
rect 630 2054 636 2055
rect 686 2059 692 2060
rect 686 2055 687 2059
rect 691 2055 692 2059
rect 686 2054 692 2055
rect 742 2059 748 2060
rect 742 2055 743 2059
rect 747 2055 748 2059
rect 742 2054 748 2055
rect 798 2059 804 2060
rect 798 2055 799 2059
rect 803 2055 804 2059
rect 798 2054 804 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 902 2059 908 2060
rect 902 2055 903 2059
rect 907 2055 908 2059
rect 902 2054 908 2055
rect 958 2059 964 2060
rect 958 2055 959 2059
rect 963 2055 964 2059
rect 958 2054 964 2055
rect 1014 2059 1020 2060
rect 1014 2055 1015 2059
rect 1019 2055 1020 2059
rect 1014 2054 1020 2055
rect 1070 2059 1076 2060
rect 1070 2055 1071 2059
rect 1075 2055 1076 2059
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 1070 2054 1076 2055
rect 1302 2037 1308 2038
rect 110 2036 116 2037
rect 110 2032 111 2036
rect 115 2032 116 2036
rect 110 2031 116 2032
rect 1238 2036 1244 2037
rect 1238 2032 1239 2036
rect 1243 2032 1244 2036
rect 1302 2033 1303 2037
rect 1307 2033 1308 2037
rect 1302 2032 1308 2033
rect 1342 2037 1348 2038
rect 1342 2033 1343 2037
rect 1347 2033 1348 2037
rect 1342 2032 1348 2033
rect 1398 2037 1404 2038
rect 1398 2033 1399 2037
rect 1403 2033 1404 2037
rect 1398 2032 1404 2033
rect 1478 2037 1484 2038
rect 1478 2033 1479 2037
rect 1483 2033 1484 2037
rect 1478 2032 1484 2033
rect 1566 2037 1572 2038
rect 1566 2033 1567 2037
rect 1571 2033 1572 2037
rect 1566 2032 1572 2033
rect 1662 2037 1668 2038
rect 1662 2033 1663 2037
rect 1667 2033 1668 2037
rect 1662 2032 1668 2033
rect 1758 2037 1764 2038
rect 1758 2033 1759 2037
rect 1763 2033 1764 2037
rect 1758 2032 1764 2033
rect 1846 2037 1852 2038
rect 1846 2033 1847 2037
rect 1851 2033 1852 2037
rect 1846 2032 1852 2033
rect 1934 2037 1940 2038
rect 1934 2033 1935 2037
rect 1939 2033 1940 2037
rect 1934 2032 1940 2033
rect 2014 2037 2020 2038
rect 2014 2033 2015 2037
rect 2019 2033 2020 2037
rect 2014 2032 2020 2033
rect 2094 2037 2100 2038
rect 2094 2033 2095 2037
rect 2099 2033 2100 2037
rect 2094 2032 2100 2033
rect 2166 2037 2172 2038
rect 2166 2033 2167 2037
rect 2171 2033 2172 2037
rect 2166 2032 2172 2033
rect 2238 2037 2244 2038
rect 2238 2033 2239 2037
rect 2243 2033 2244 2037
rect 2238 2032 2244 2033
rect 2310 2037 2316 2038
rect 2310 2033 2311 2037
rect 2315 2033 2316 2037
rect 2310 2032 2316 2033
rect 2358 2037 2364 2038
rect 2358 2033 2359 2037
rect 2363 2033 2364 2037
rect 2358 2032 2364 2033
rect 1238 2031 1244 2032
rect 110 2019 116 2020
rect 110 2015 111 2019
rect 115 2015 116 2019
rect 110 2014 116 2015
rect 1238 2019 1244 2020
rect 1238 2015 1239 2019
rect 1243 2015 1244 2019
rect 1238 2014 1244 2015
rect 382 2012 388 2013
rect 382 2008 383 2012
rect 387 2008 388 2012
rect 382 2007 388 2008
rect 422 2012 428 2013
rect 422 2008 423 2012
rect 427 2008 428 2012
rect 422 2007 428 2008
rect 462 2012 468 2013
rect 462 2008 463 2012
rect 467 2008 468 2012
rect 462 2007 468 2008
rect 502 2012 508 2013
rect 502 2008 503 2012
rect 507 2008 508 2012
rect 502 2007 508 2008
rect 542 2012 548 2013
rect 542 2008 543 2012
rect 547 2008 548 2012
rect 542 2007 548 2008
rect 582 2012 588 2013
rect 582 2008 583 2012
rect 587 2008 588 2012
rect 582 2007 588 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 686 2012 692 2013
rect 686 2008 687 2012
rect 691 2008 692 2012
rect 686 2007 692 2008
rect 742 2012 748 2013
rect 742 2008 743 2012
rect 747 2008 748 2012
rect 742 2007 748 2008
rect 798 2012 804 2013
rect 798 2008 799 2012
rect 803 2008 804 2012
rect 798 2007 804 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 902 2012 908 2013
rect 902 2008 903 2012
rect 907 2008 908 2012
rect 902 2007 908 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1014 2012 1020 2013
rect 1014 2008 1015 2012
rect 1019 2008 1020 2012
rect 1014 2007 1020 2008
rect 1070 2012 1076 2013
rect 1070 2008 1071 2012
rect 1075 2008 1076 2012
rect 1070 2007 1076 2008
rect 1302 1999 1308 2000
rect 1302 1995 1303 1999
rect 1307 1995 1308 1999
rect 1302 1994 1308 1995
rect 1350 1999 1356 2000
rect 1350 1995 1351 1999
rect 1355 1995 1356 1999
rect 1350 1994 1356 1995
rect 1422 1999 1428 2000
rect 1422 1995 1423 1999
rect 1427 1995 1428 1999
rect 1422 1994 1428 1995
rect 1494 1999 1500 2000
rect 1494 1995 1495 1999
rect 1499 1995 1500 1999
rect 1494 1994 1500 1995
rect 1574 1999 1580 2000
rect 1574 1995 1575 1999
rect 1579 1995 1580 1999
rect 1574 1994 1580 1995
rect 1662 1999 1668 2000
rect 1662 1995 1663 1999
rect 1667 1995 1668 1999
rect 1662 1994 1668 1995
rect 1750 1999 1756 2000
rect 1750 1995 1751 1999
rect 1755 1995 1756 1999
rect 1750 1994 1756 1995
rect 1838 1999 1844 2000
rect 1838 1995 1839 1999
rect 1843 1995 1844 1999
rect 1838 1994 1844 1995
rect 1918 1999 1924 2000
rect 1918 1995 1919 1999
rect 1923 1995 1924 1999
rect 1918 1994 1924 1995
rect 1998 1999 2004 2000
rect 1998 1995 1999 1999
rect 2003 1995 2004 1999
rect 1998 1994 2004 1995
rect 2070 1999 2076 2000
rect 2070 1995 2071 1999
rect 2075 1995 2076 1999
rect 2070 1994 2076 1995
rect 2134 1999 2140 2000
rect 2134 1995 2135 1999
rect 2139 1995 2140 1999
rect 2134 1994 2140 1995
rect 2190 1999 2196 2000
rect 2190 1995 2191 1999
rect 2195 1995 2196 1999
rect 2190 1994 2196 1995
rect 2254 1999 2260 2000
rect 2254 1995 2255 1999
rect 2259 1995 2260 1999
rect 2254 1994 2260 1995
rect 2318 1999 2324 2000
rect 2318 1995 2319 1999
rect 2323 1995 2324 1999
rect 2318 1994 2324 1995
rect 2358 1999 2364 2000
rect 2358 1995 2359 1999
rect 2363 1995 2364 1999
rect 2358 1994 2364 1995
rect 366 1992 372 1993
rect 366 1988 367 1992
rect 371 1988 372 1992
rect 366 1987 372 1988
rect 406 1992 412 1993
rect 406 1988 407 1992
rect 411 1988 412 1992
rect 406 1987 412 1988
rect 454 1992 460 1993
rect 454 1988 455 1992
rect 459 1988 460 1992
rect 454 1987 460 1988
rect 510 1992 516 1993
rect 510 1988 511 1992
rect 515 1988 516 1992
rect 510 1987 516 1988
rect 566 1992 572 1993
rect 566 1988 567 1992
rect 571 1988 572 1992
rect 566 1987 572 1988
rect 630 1992 636 1993
rect 630 1988 631 1992
rect 635 1988 636 1992
rect 630 1987 636 1988
rect 694 1992 700 1993
rect 694 1988 695 1992
rect 699 1988 700 1992
rect 694 1987 700 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 870 1992 876 1993
rect 870 1988 871 1992
rect 875 1988 876 1992
rect 870 1987 876 1988
rect 934 1992 940 1993
rect 934 1988 935 1992
rect 939 1988 940 1992
rect 934 1987 940 1988
rect 998 1992 1004 1993
rect 998 1988 999 1992
rect 1003 1988 1004 1992
rect 998 1987 1004 1988
rect 1062 1992 1068 1993
rect 1062 1988 1063 1992
rect 1067 1988 1068 1992
rect 1062 1987 1068 1988
rect 110 1985 116 1986
rect 110 1981 111 1985
rect 115 1981 116 1985
rect 110 1980 116 1981
rect 1238 1985 1244 1986
rect 1238 1981 1239 1985
rect 1243 1981 1244 1985
rect 1238 1980 1244 1981
rect 1278 1976 1284 1977
rect 1278 1972 1279 1976
rect 1283 1972 1284 1976
rect 1278 1971 1284 1972
rect 2406 1976 2412 1977
rect 2406 1972 2407 1976
rect 2411 1972 2412 1976
rect 2406 1971 2412 1972
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 1238 1968 1244 1969
rect 1238 1964 1239 1968
rect 1243 1964 1244 1968
rect 1238 1963 1244 1964
rect 1278 1959 1284 1960
rect 1278 1955 1279 1959
rect 1283 1955 1284 1959
rect 1278 1954 1284 1955
rect 2406 1959 2412 1960
rect 2406 1955 2407 1959
rect 2411 1955 2412 1959
rect 2406 1954 2412 1955
rect 1302 1952 1308 1953
rect 1302 1948 1303 1952
rect 1307 1948 1308 1952
rect 1302 1947 1308 1948
rect 1350 1952 1356 1953
rect 1350 1948 1351 1952
rect 1355 1948 1356 1952
rect 1350 1947 1356 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1494 1952 1500 1953
rect 1494 1948 1495 1952
rect 1499 1948 1500 1952
rect 1494 1947 1500 1948
rect 1574 1952 1580 1953
rect 1574 1948 1575 1952
rect 1579 1948 1580 1952
rect 1574 1947 1580 1948
rect 1662 1952 1668 1953
rect 1662 1948 1663 1952
rect 1667 1948 1668 1952
rect 1662 1947 1668 1948
rect 1750 1952 1756 1953
rect 1750 1948 1751 1952
rect 1755 1948 1756 1952
rect 1750 1947 1756 1948
rect 1838 1952 1844 1953
rect 1838 1948 1839 1952
rect 1843 1948 1844 1952
rect 1838 1947 1844 1948
rect 1918 1952 1924 1953
rect 1918 1948 1919 1952
rect 1923 1948 1924 1952
rect 1918 1947 1924 1948
rect 1998 1952 2004 1953
rect 1998 1948 1999 1952
rect 2003 1948 2004 1952
rect 1998 1947 2004 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2134 1952 2140 1953
rect 2134 1948 2135 1952
rect 2139 1948 2140 1952
rect 2134 1947 2140 1948
rect 2190 1952 2196 1953
rect 2190 1948 2191 1952
rect 2195 1948 2196 1952
rect 2190 1947 2196 1948
rect 2254 1952 2260 1953
rect 2254 1948 2255 1952
rect 2259 1948 2260 1952
rect 2254 1947 2260 1948
rect 2318 1952 2324 1953
rect 2318 1948 2319 1952
rect 2323 1948 2324 1952
rect 2318 1947 2324 1948
rect 2358 1952 2364 1953
rect 2358 1948 2359 1952
rect 2363 1948 2364 1952
rect 2358 1947 2364 1948
rect 366 1945 372 1946
rect 366 1941 367 1945
rect 371 1941 372 1945
rect 366 1940 372 1941
rect 406 1945 412 1946
rect 406 1941 407 1945
rect 411 1941 412 1945
rect 406 1940 412 1941
rect 454 1945 460 1946
rect 454 1941 455 1945
rect 459 1941 460 1945
rect 454 1940 460 1941
rect 510 1945 516 1946
rect 510 1941 511 1945
rect 515 1941 516 1945
rect 510 1940 516 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 630 1945 636 1946
rect 630 1941 631 1945
rect 635 1941 636 1945
rect 630 1940 636 1941
rect 694 1945 700 1946
rect 694 1941 695 1945
rect 699 1941 700 1945
rect 694 1940 700 1941
rect 758 1945 764 1946
rect 758 1941 759 1945
rect 763 1941 764 1945
rect 758 1940 764 1941
rect 814 1945 820 1946
rect 814 1941 815 1945
rect 819 1941 820 1945
rect 814 1940 820 1941
rect 870 1945 876 1946
rect 870 1941 871 1945
rect 875 1941 876 1945
rect 870 1940 876 1941
rect 934 1945 940 1946
rect 934 1941 935 1945
rect 939 1941 940 1945
rect 934 1940 940 1941
rect 998 1945 1004 1946
rect 998 1941 999 1945
rect 1003 1941 1004 1945
rect 998 1940 1004 1941
rect 1062 1945 1068 1946
rect 1062 1941 1063 1945
rect 1067 1941 1068 1945
rect 1062 1940 1068 1941
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1358 1940 1364 1941
rect 1358 1936 1359 1940
rect 1363 1936 1364 1940
rect 1358 1935 1364 1936
rect 1446 1940 1452 1941
rect 1446 1936 1447 1940
rect 1451 1936 1452 1940
rect 1446 1935 1452 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1622 1940 1628 1941
rect 1622 1936 1623 1940
rect 1627 1936 1628 1940
rect 1622 1935 1628 1936
rect 1710 1940 1716 1941
rect 1710 1936 1711 1940
rect 1715 1936 1716 1940
rect 1710 1935 1716 1936
rect 1790 1940 1796 1941
rect 1790 1936 1791 1940
rect 1795 1936 1796 1940
rect 1790 1935 1796 1936
rect 1862 1940 1868 1941
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 1934 1940 1940 1941
rect 1934 1936 1935 1940
rect 1939 1936 1940 1940
rect 1934 1935 1940 1936
rect 2006 1940 2012 1941
rect 2006 1936 2007 1940
rect 2011 1936 2012 1940
rect 2006 1935 2012 1936
rect 2078 1940 2084 1941
rect 2078 1936 2079 1940
rect 2083 1936 2084 1940
rect 2078 1935 2084 1936
rect 2150 1940 2156 1941
rect 2150 1936 2151 1940
rect 2155 1936 2156 1940
rect 2150 1935 2156 1936
rect 2222 1940 2228 1941
rect 2222 1936 2223 1940
rect 2227 1936 2228 1940
rect 2222 1935 2228 1936
rect 2302 1940 2308 1941
rect 2302 1936 2303 1940
rect 2307 1936 2308 1940
rect 2302 1935 2308 1936
rect 2358 1940 2364 1941
rect 2358 1936 2359 1940
rect 2363 1936 2364 1940
rect 2358 1935 2364 1936
rect 1278 1933 1284 1934
rect 1278 1929 1279 1933
rect 1283 1929 1284 1933
rect 1278 1928 1284 1929
rect 2406 1933 2412 1934
rect 2406 1929 2407 1933
rect 2411 1929 2412 1933
rect 2406 1928 2412 1929
rect 1278 1916 1284 1917
rect 1278 1912 1279 1916
rect 1283 1912 1284 1916
rect 174 1911 180 1912
rect 174 1907 175 1911
rect 179 1907 180 1911
rect 174 1906 180 1907
rect 214 1911 220 1912
rect 214 1907 215 1911
rect 219 1907 220 1911
rect 214 1906 220 1907
rect 262 1911 268 1912
rect 262 1907 263 1911
rect 267 1907 268 1911
rect 262 1906 268 1907
rect 318 1911 324 1912
rect 318 1907 319 1911
rect 323 1907 324 1911
rect 318 1906 324 1907
rect 390 1911 396 1912
rect 390 1907 391 1911
rect 395 1907 396 1911
rect 390 1906 396 1907
rect 470 1911 476 1912
rect 470 1907 471 1911
rect 475 1907 476 1911
rect 470 1906 476 1907
rect 550 1911 556 1912
rect 550 1907 551 1911
rect 555 1907 556 1911
rect 550 1906 556 1907
rect 638 1911 644 1912
rect 638 1907 639 1911
rect 643 1907 644 1911
rect 638 1906 644 1907
rect 718 1911 724 1912
rect 718 1907 719 1911
rect 723 1907 724 1911
rect 718 1906 724 1907
rect 798 1911 804 1912
rect 798 1907 799 1911
rect 803 1907 804 1911
rect 798 1906 804 1907
rect 878 1911 884 1912
rect 878 1907 879 1911
rect 883 1907 884 1911
rect 878 1906 884 1907
rect 958 1911 964 1912
rect 958 1907 959 1911
rect 963 1907 964 1911
rect 958 1906 964 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1118 1911 1124 1912
rect 1278 1911 1284 1912
rect 2406 1916 2412 1917
rect 2406 1912 2407 1916
rect 2411 1912 2412 1916
rect 2406 1911 2412 1912
rect 1118 1907 1119 1911
rect 1123 1907 1124 1911
rect 1118 1906 1124 1907
rect 1302 1893 1308 1894
rect 1302 1889 1303 1893
rect 1307 1889 1308 1893
rect 110 1888 116 1889
rect 110 1884 111 1888
rect 115 1884 116 1888
rect 110 1883 116 1884
rect 1238 1888 1244 1889
rect 1302 1888 1308 1889
rect 1358 1893 1364 1894
rect 1358 1889 1359 1893
rect 1363 1889 1364 1893
rect 1358 1888 1364 1889
rect 1446 1893 1452 1894
rect 1446 1889 1447 1893
rect 1451 1889 1452 1893
rect 1446 1888 1452 1889
rect 1534 1893 1540 1894
rect 1534 1889 1535 1893
rect 1539 1889 1540 1893
rect 1534 1888 1540 1889
rect 1622 1893 1628 1894
rect 1622 1889 1623 1893
rect 1627 1889 1628 1893
rect 1622 1888 1628 1889
rect 1710 1893 1716 1894
rect 1710 1889 1711 1893
rect 1715 1889 1716 1893
rect 1710 1888 1716 1889
rect 1790 1893 1796 1894
rect 1790 1889 1791 1893
rect 1795 1889 1796 1893
rect 1790 1888 1796 1889
rect 1862 1893 1868 1894
rect 1862 1889 1863 1893
rect 1867 1889 1868 1893
rect 1862 1888 1868 1889
rect 1934 1893 1940 1894
rect 1934 1889 1935 1893
rect 1939 1889 1940 1893
rect 1934 1888 1940 1889
rect 2006 1893 2012 1894
rect 2006 1889 2007 1893
rect 2011 1889 2012 1893
rect 2006 1888 2012 1889
rect 2078 1893 2084 1894
rect 2078 1889 2079 1893
rect 2083 1889 2084 1893
rect 2078 1888 2084 1889
rect 2150 1893 2156 1894
rect 2150 1889 2151 1893
rect 2155 1889 2156 1893
rect 2150 1888 2156 1889
rect 2222 1893 2228 1894
rect 2222 1889 2223 1893
rect 2227 1889 2228 1893
rect 2222 1888 2228 1889
rect 2302 1893 2308 1894
rect 2302 1889 2303 1893
rect 2307 1889 2308 1893
rect 2302 1888 2308 1889
rect 2358 1893 2364 1894
rect 2358 1889 2359 1893
rect 2363 1889 2364 1893
rect 2358 1888 2364 1889
rect 1238 1884 1239 1888
rect 1243 1884 1244 1888
rect 1238 1883 1244 1884
rect 110 1871 116 1872
rect 110 1867 111 1871
rect 115 1867 116 1871
rect 110 1866 116 1867
rect 1238 1871 1244 1872
rect 1238 1867 1239 1871
rect 1243 1867 1244 1871
rect 1238 1866 1244 1867
rect 174 1864 180 1865
rect 174 1860 175 1864
rect 179 1860 180 1864
rect 174 1859 180 1860
rect 214 1864 220 1865
rect 214 1860 215 1864
rect 219 1860 220 1864
rect 214 1859 220 1860
rect 262 1864 268 1865
rect 262 1860 263 1864
rect 267 1860 268 1864
rect 262 1859 268 1860
rect 318 1864 324 1865
rect 318 1860 319 1864
rect 323 1860 324 1864
rect 318 1859 324 1860
rect 390 1864 396 1865
rect 390 1860 391 1864
rect 395 1860 396 1864
rect 390 1859 396 1860
rect 470 1864 476 1865
rect 470 1860 471 1864
rect 475 1860 476 1864
rect 470 1859 476 1860
rect 550 1864 556 1865
rect 550 1860 551 1864
rect 555 1860 556 1864
rect 550 1859 556 1860
rect 638 1864 644 1865
rect 638 1860 639 1864
rect 643 1860 644 1864
rect 638 1859 644 1860
rect 718 1864 724 1865
rect 718 1860 719 1864
rect 723 1860 724 1864
rect 718 1859 724 1860
rect 798 1864 804 1865
rect 798 1860 799 1864
rect 803 1860 804 1864
rect 798 1859 804 1860
rect 878 1864 884 1865
rect 878 1860 879 1864
rect 883 1860 884 1864
rect 878 1859 884 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1038 1864 1044 1865
rect 1038 1860 1039 1864
rect 1043 1860 1044 1864
rect 1038 1859 1044 1860
rect 1118 1864 1124 1865
rect 1118 1860 1119 1864
rect 1123 1860 1124 1864
rect 1118 1859 1124 1860
rect 1310 1863 1316 1864
rect 1310 1859 1311 1863
rect 1315 1859 1316 1863
rect 1310 1858 1316 1859
rect 1358 1863 1364 1864
rect 1358 1859 1359 1863
rect 1363 1859 1364 1863
rect 1358 1858 1364 1859
rect 1414 1863 1420 1864
rect 1414 1859 1415 1863
rect 1419 1859 1420 1863
rect 1414 1858 1420 1859
rect 1478 1863 1484 1864
rect 1478 1859 1479 1863
rect 1483 1859 1484 1863
rect 1478 1858 1484 1859
rect 1542 1863 1548 1864
rect 1542 1859 1543 1863
rect 1547 1859 1548 1863
rect 1542 1858 1548 1859
rect 1614 1863 1620 1864
rect 1614 1859 1615 1863
rect 1619 1859 1620 1863
rect 1614 1858 1620 1859
rect 1686 1863 1692 1864
rect 1686 1859 1687 1863
rect 1691 1859 1692 1863
rect 1686 1858 1692 1859
rect 1766 1863 1772 1864
rect 1766 1859 1767 1863
rect 1771 1859 1772 1863
rect 1766 1858 1772 1859
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 1974 1863 1980 1864
rect 1974 1859 1975 1863
rect 1979 1859 1980 1863
rect 1974 1858 1980 1859
rect 2094 1863 2100 1864
rect 2094 1859 2095 1863
rect 2099 1859 2100 1863
rect 2094 1858 2100 1859
rect 2222 1863 2228 1864
rect 2222 1859 2223 1863
rect 2227 1859 2228 1863
rect 2222 1858 2228 1859
rect 2358 1863 2364 1864
rect 2358 1859 2359 1863
rect 2363 1859 2364 1863
rect 2358 1858 2364 1859
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 214 1844 220 1845
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 270 1844 276 1845
rect 270 1840 271 1844
rect 275 1840 276 1844
rect 270 1839 276 1840
rect 350 1844 356 1845
rect 350 1840 351 1844
rect 355 1840 356 1844
rect 350 1839 356 1840
rect 438 1844 444 1845
rect 438 1840 439 1844
rect 443 1840 444 1844
rect 438 1839 444 1840
rect 534 1844 540 1845
rect 534 1840 535 1844
rect 539 1840 540 1844
rect 534 1839 540 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 726 1844 732 1845
rect 726 1840 727 1844
rect 731 1840 732 1844
rect 726 1839 732 1840
rect 822 1844 828 1845
rect 822 1840 823 1844
rect 827 1840 828 1844
rect 822 1839 828 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 990 1844 996 1845
rect 990 1840 991 1844
rect 995 1840 996 1844
rect 990 1839 996 1840
rect 1062 1844 1068 1845
rect 1062 1840 1063 1844
rect 1067 1840 1068 1844
rect 1062 1839 1068 1840
rect 1134 1844 1140 1845
rect 1134 1840 1135 1844
rect 1139 1840 1140 1844
rect 1134 1839 1140 1840
rect 1190 1844 1196 1845
rect 1190 1840 1191 1844
rect 1195 1840 1196 1844
rect 1190 1839 1196 1840
rect 1278 1840 1284 1841
rect 110 1837 116 1838
rect 110 1833 111 1837
rect 115 1833 116 1837
rect 110 1832 116 1833
rect 1238 1837 1244 1838
rect 1238 1833 1239 1837
rect 1243 1833 1244 1837
rect 1278 1836 1279 1840
rect 1283 1836 1284 1840
rect 1278 1835 1284 1836
rect 2406 1840 2412 1841
rect 2406 1836 2407 1840
rect 2411 1836 2412 1840
rect 2406 1835 2412 1836
rect 1238 1832 1244 1833
rect 1278 1823 1284 1824
rect 110 1820 116 1821
rect 110 1816 111 1820
rect 115 1816 116 1820
rect 110 1815 116 1816
rect 1238 1820 1244 1821
rect 1238 1816 1239 1820
rect 1243 1816 1244 1820
rect 1278 1819 1279 1823
rect 1283 1819 1284 1823
rect 1278 1818 1284 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 1238 1815 1244 1816
rect 1310 1816 1316 1817
rect 1310 1812 1311 1816
rect 1315 1812 1316 1816
rect 1310 1811 1316 1812
rect 1358 1816 1364 1817
rect 1358 1812 1359 1816
rect 1363 1812 1364 1816
rect 1358 1811 1364 1812
rect 1414 1816 1420 1817
rect 1414 1812 1415 1816
rect 1419 1812 1420 1816
rect 1414 1811 1420 1812
rect 1478 1816 1484 1817
rect 1478 1812 1479 1816
rect 1483 1812 1484 1816
rect 1478 1811 1484 1812
rect 1542 1816 1548 1817
rect 1542 1812 1543 1816
rect 1547 1812 1548 1816
rect 1542 1811 1548 1812
rect 1614 1816 1620 1817
rect 1614 1812 1615 1816
rect 1619 1812 1620 1816
rect 1614 1811 1620 1812
rect 1686 1816 1692 1817
rect 1686 1812 1687 1816
rect 1691 1812 1692 1816
rect 1686 1811 1692 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1862 1816 1868 1817
rect 1862 1812 1863 1816
rect 1867 1812 1868 1816
rect 1862 1811 1868 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2094 1816 2100 1817
rect 2094 1812 2095 1816
rect 2099 1812 2100 1816
rect 2094 1811 2100 1812
rect 2222 1816 2228 1817
rect 2222 1812 2223 1816
rect 2227 1812 2228 1816
rect 2222 1811 2228 1812
rect 2358 1816 2364 1817
rect 2358 1812 2359 1816
rect 2363 1812 2364 1816
rect 2358 1811 2364 1812
rect 1406 1800 1412 1801
rect 134 1797 140 1798
rect 134 1793 135 1797
rect 139 1793 140 1797
rect 134 1792 140 1793
rect 174 1797 180 1798
rect 174 1793 175 1797
rect 179 1793 180 1797
rect 174 1792 180 1793
rect 214 1797 220 1798
rect 214 1793 215 1797
rect 219 1793 220 1797
rect 214 1792 220 1793
rect 270 1797 276 1798
rect 270 1793 271 1797
rect 275 1793 276 1797
rect 270 1792 276 1793
rect 350 1797 356 1798
rect 350 1793 351 1797
rect 355 1793 356 1797
rect 350 1792 356 1793
rect 438 1797 444 1798
rect 438 1793 439 1797
rect 443 1793 444 1797
rect 438 1792 444 1793
rect 534 1797 540 1798
rect 534 1793 535 1797
rect 539 1793 540 1797
rect 534 1792 540 1793
rect 630 1797 636 1798
rect 630 1793 631 1797
rect 635 1793 636 1797
rect 630 1792 636 1793
rect 726 1797 732 1798
rect 726 1793 727 1797
rect 731 1793 732 1797
rect 726 1792 732 1793
rect 822 1797 828 1798
rect 822 1793 823 1797
rect 827 1793 828 1797
rect 822 1792 828 1793
rect 910 1797 916 1798
rect 910 1793 911 1797
rect 915 1793 916 1797
rect 910 1792 916 1793
rect 990 1797 996 1798
rect 990 1793 991 1797
rect 995 1793 996 1797
rect 990 1792 996 1793
rect 1062 1797 1068 1798
rect 1062 1793 1063 1797
rect 1067 1793 1068 1797
rect 1062 1792 1068 1793
rect 1134 1797 1140 1798
rect 1134 1793 1135 1797
rect 1139 1793 1140 1797
rect 1134 1792 1140 1793
rect 1190 1797 1196 1798
rect 1190 1793 1191 1797
rect 1195 1793 1196 1797
rect 1406 1796 1407 1800
rect 1411 1796 1412 1800
rect 1406 1795 1412 1796
rect 1470 1800 1476 1801
rect 1470 1796 1471 1800
rect 1475 1796 1476 1800
rect 1470 1795 1476 1796
rect 1534 1800 1540 1801
rect 1534 1796 1535 1800
rect 1539 1796 1540 1800
rect 1534 1795 1540 1796
rect 1598 1800 1604 1801
rect 1598 1796 1599 1800
rect 1603 1796 1604 1800
rect 1598 1795 1604 1796
rect 1662 1800 1668 1801
rect 1662 1796 1663 1800
rect 1667 1796 1668 1800
rect 1662 1795 1668 1796
rect 1726 1800 1732 1801
rect 1726 1796 1727 1800
rect 1731 1796 1732 1800
rect 1726 1795 1732 1796
rect 1782 1800 1788 1801
rect 1782 1796 1783 1800
rect 1787 1796 1788 1800
rect 1782 1795 1788 1796
rect 1838 1800 1844 1801
rect 1838 1796 1839 1800
rect 1843 1796 1844 1800
rect 1838 1795 1844 1796
rect 1894 1800 1900 1801
rect 1894 1796 1895 1800
rect 1899 1796 1900 1800
rect 1894 1795 1900 1796
rect 1958 1800 1964 1801
rect 1958 1796 1959 1800
rect 1963 1796 1964 1800
rect 1958 1795 1964 1796
rect 1190 1792 1196 1793
rect 1278 1793 1284 1794
rect 1278 1789 1279 1793
rect 1283 1789 1284 1793
rect 1278 1788 1284 1789
rect 2406 1793 2412 1794
rect 2406 1789 2407 1793
rect 2411 1789 2412 1793
rect 2406 1788 2412 1789
rect 1278 1776 1284 1777
rect 1278 1772 1279 1776
rect 1283 1772 1284 1776
rect 1278 1771 1284 1772
rect 2406 1776 2412 1777
rect 2406 1772 2407 1776
rect 2411 1772 2412 1776
rect 2406 1771 2412 1772
rect 134 1767 140 1768
rect 134 1763 135 1767
rect 139 1763 140 1767
rect 134 1762 140 1763
rect 174 1767 180 1768
rect 174 1763 175 1767
rect 179 1763 180 1767
rect 174 1762 180 1763
rect 214 1767 220 1768
rect 214 1763 215 1767
rect 219 1763 220 1767
rect 214 1762 220 1763
rect 286 1767 292 1768
rect 286 1763 287 1767
rect 291 1763 292 1767
rect 286 1762 292 1763
rect 374 1767 380 1768
rect 374 1763 375 1767
rect 379 1763 380 1767
rect 374 1762 380 1763
rect 470 1767 476 1768
rect 470 1763 471 1767
rect 475 1763 476 1767
rect 470 1762 476 1763
rect 566 1767 572 1768
rect 566 1763 567 1767
rect 571 1763 572 1767
rect 566 1762 572 1763
rect 662 1767 668 1768
rect 662 1763 663 1767
rect 667 1763 668 1767
rect 662 1762 668 1763
rect 750 1767 756 1768
rect 750 1763 751 1767
rect 755 1763 756 1767
rect 750 1762 756 1763
rect 830 1767 836 1768
rect 830 1763 831 1767
rect 835 1763 836 1767
rect 830 1762 836 1763
rect 902 1767 908 1768
rect 902 1763 903 1767
rect 907 1763 908 1767
rect 902 1762 908 1763
rect 966 1767 972 1768
rect 966 1763 967 1767
rect 971 1763 972 1767
rect 966 1762 972 1763
rect 1030 1767 1036 1768
rect 1030 1763 1031 1767
rect 1035 1763 1036 1767
rect 1030 1762 1036 1763
rect 1086 1767 1092 1768
rect 1086 1763 1087 1767
rect 1091 1763 1092 1767
rect 1086 1762 1092 1763
rect 1150 1767 1156 1768
rect 1150 1763 1151 1767
rect 1155 1763 1156 1767
rect 1150 1762 1156 1763
rect 1190 1767 1196 1768
rect 1190 1763 1191 1767
rect 1195 1763 1196 1767
rect 1190 1762 1196 1763
rect 1406 1753 1412 1754
rect 1406 1749 1407 1753
rect 1411 1749 1412 1753
rect 1406 1748 1412 1749
rect 1470 1753 1476 1754
rect 1470 1749 1471 1753
rect 1475 1749 1476 1753
rect 1470 1748 1476 1749
rect 1534 1753 1540 1754
rect 1534 1749 1535 1753
rect 1539 1749 1540 1753
rect 1534 1748 1540 1749
rect 1598 1753 1604 1754
rect 1598 1749 1599 1753
rect 1603 1749 1604 1753
rect 1598 1748 1604 1749
rect 1662 1753 1668 1754
rect 1662 1749 1663 1753
rect 1667 1749 1668 1753
rect 1662 1748 1668 1749
rect 1726 1753 1732 1754
rect 1726 1749 1727 1753
rect 1731 1749 1732 1753
rect 1726 1748 1732 1749
rect 1782 1753 1788 1754
rect 1782 1749 1783 1753
rect 1787 1749 1788 1753
rect 1782 1748 1788 1749
rect 1838 1753 1844 1754
rect 1838 1749 1839 1753
rect 1843 1749 1844 1753
rect 1838 1748 1844 1749
rect 1894 1753 1900 1754
rect 1894 1749 1895 1753
rect 1899 1749 1900 1753
rect 1894 1748 1900 1749
rect 1958 1753 1964 1754
rect 1958 1749 1959 1753
rect 1963 1749 1964 1753
rect 1958 1748 1964 1749
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 1238 1744 1244 1745
rect 1238 1740 1239 1744
rect 1243 1740 1244 1744
rect 1238 1739 1244 1740
rect 110 1727 116 1728
rect 110 1723 111 1727
rect 115 1723 116 1727
rect 110 1722 116 1723
rect 1238 1727 1244 1728
rect 1238 1723 1239 1727
rect 1243 1723 1244 1727
rect 1238 1722 1244 1723
rect 1302 1723 1308 1724
rect 134 1720 140 1721
rect 134 1716 135 1720
rect 139 1716 140 1720
rect 134 1715 140 1716
rect 174 1720 180 1721
rect 174 1716 175 1720
rect 179 1716 180 1720
rect 174 1715 180 1716
rect 214 1720 220 1721
rect 214 1716 215 1720
rect 219 1716 220 1720
rect 214 1715 220 1716
rect 286 1720 292 1721
rect 286 1716 287 1720
rect 291 1716 292 1720
rect 286 1715 292 1716
rect 374 1720 380 1721
rect 374 1716 375 1720
rect 379 1716 380 1720
rect 374 1715 380 1716
rect 470 1720 476 1721
rect 470 1716 471 1720
rect 475 1716 476 1720
rect 470 1715 476 1716
rect 566 1720 572 1721
rect 566 1716 567 1720
rect 571 1716 572 1720
rect 566 1715 572 1716
rect 662 1720 668 1721
rect 662 1716 663 1720
rect 667 1716 668 1720
rect 662 1715 668 1716
rect 750 1720 756 1721
rect 750 1716 751 1720
rect 755 1716 756 1720
rect 750 1715 756 1716
rect 830 1720 836 1721
rect 830 1716 831 1720
rect 835 1716 836 1720
rect 830 1715 836 1716
rect 902 1720 908 1721
rect 902 1716 903 1720
rect 907 1716 908 1720
rect 902 1715 908 1716
rect 966 1720 972 1721
rect 966 1716 967 1720
rect 971 1716 972 1720
rect 966 1715 972 1716
rect 1030 1720 1036 1721
rect 1030 1716 1031 1720
rect 1035 1716 1036 1720
rect 1030 1715 1036 1716
rect 1086 1720 1092 1721
rect 1086 1716 1087 1720
rect 1091 1716 1092 1720
rect 1086 1715 1092 1716
rect 1150 1720 1156 1721
rect 1150 1716 1151 1720
rect 1155 1716 1156 1720
rect 1150 1715 1156 1716
rect 1190 1720 1196 1721
rect 1190 1716 1191 1720
rect 1195 1716 1196 1720
rect 1302 1719 1303 1723
rect 1307 1719 1308 1723
rect 1302 1718 1308 1719
rect 1350 1723 1356 1724
rect 1350 1719 1351 1723
rect 1355 1719 1356 1723
rect 1350 1718 1356 1719
rect 1422 1723 1428 1724
rect 1422 1719 1423 1723
rect 1427 1719 1428 1723
rect 1422 1718 1428 1719
rect 1502 1723 1508 1724
rect 1502 1719 1503 1723
rect 1507 1719 1508 1723
rect 1502 1718 1508 1719
rect 1582 1723 1588 1724
rect 1582 1719 1583 1723
rect 1587 1719 1588 1723
rect 1582 1718 1588 1719
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1719 1668 1723
rect 1662 1718 1668 1719
rect 1734 1723 1740 1724
rect 1734 1719 1735 1723
rect 1739 1719 1740 1723
rect 1734 1718 1740 1719
rect 1806 1723 1812 1724
rect 1806 1719 1807 1723
rect 1811 1719 1812 1723
rect 1806 1718 1812 1719
rect 1870 1723 1876 1724
rect 1870 1719 1871 1723
rect 1875 1719 1876 1723
rect 1870 1718 1876 1719
rect 1934 1723 1940 1724
rect 1934 1719 1935 1723
rect 1939 1719 1940 1723
rect 1934 1718 1940 1719
rect 1998 1723 2004 1724
rect 1998 1719 1999 1723
rect 2003 1719 2004 1723
rect 1998 1718 2004 1719
rect 2062 1723 2068 1724
rect 2062 1719 2063 1723
rect 2067 1719 2068 1723
rect 2062 1718 2068 1719
rect 1190 1715 1196 1716
rect 134 1704 140 1705
rect 134 1700 135 1704
rect 139 1700 140 1704
rect 134 1699 140 1700
rect 174 1704 180 1705
rect 174 1700 175 1704
rect 179 1700 180 1704
rect 174 1699 180 1700
rect 238 1704 244 1705
rect 238 1700 239 1704
rect 243 1700 244 1704
rect 238 1699 244 1700
rect 318 1704 324 1705
rect 318 1700 319 1704
rect 323 1700 324 1704
rect 318 1699 324 1700
rect 414 1704 420 1705
rect 414 1700 415 1704
rect 419 1700 420 1704
rect 414 1699 420 1700
rect 510 1704 516 1705
rect 510 1700 511 1704
rect 515 1700 516 1704
rect 510 1699 516 1700
rect 614 1704 620 1705
rect 614 1700 615 1704
rect 619 1700 620 1704
rect 614 1699 620 1700
rect 710 1704 716 1705
rect 710 1700 711 1704
rect 715 1700 716 1704
rect 710 1699 716 1700
rect 798 1704 804 1705
rect 798 1700 799 1704
rect 803 1700 804 1704
rect 798 1699 804 1700
rect 878 1704 884 1705
rect 878 1700 879 1704
rect 883 1700 884 1704
rect 878 1699 884 1700
rect 950 1704 956 1705
rect 950 1700 951 1704
rect 955 1700 956 1704
rect 950 1699 956 1700
rect 1014 1704 1020 1705
rect 1014 1700 1015 1704
rect 1019 1700 1020 1704
rect 1014 1699 1020 1700
rect 1086 1704 1092 1705
rect 1086 1700 1087 1704
rect 1091 1700 1092 1704
rect 1086 1699 1092 1700
rect 1158 1704 1164 1705
rect 1158 1700 1159 1704
rect 1163 1700 1164 1704
rect 1158 1699 1164 1700
rect 1278 1700 1284 1701
rect 110 1697 116 1698
rect 110 1693 111 1697
rect 115 1693 116 1697
rect 110 1692 116 1693
rect 1238 1697 1244 1698
rect 1238 1693 1239 1697
rect 1243 1693 1244 1697
rect 1278 1696 1279 1700
rect 1283 1696 1284 1700
rect 1278 1695 1284 1696
rect 2406 1700 2412 1701
rect 2406 1696 2407 1700
rect 2411 1696 2412 1700
rect 2406 1695 2412 1696
rect 1238 1692 1244 1693
rect 1278 1683 1284 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1238 1680 1244 1681
rect 1238 1676 1239 1680
rect 1243 1676 1244 1680
rect 1278 1679 1279 1683
rect 1283 1679 1284 1683
rect 1278 1678 1284 1679
rect 2406 1683 2412 1684
rect 2406 1679 2407 1683
rect 2411 1679 2412 1683
rect 2406 1678 2412 1679
rect 1238 1675 1244 1676
rect 1302 1676 1308 1677
rect 1302 1672 1303 1676
rect 1307 1672 1308 1676
rect 1302 1671 1308 1672
rect 1350 1676 1356 1677
rect 1350 1672 1351 1676
rect 1355 1672 1356 1676
rect 1350 1671 1356 1672
rect 1422 1676 1428 1677
rect 1422 1672 1423 1676
rect 1427 1672 1428 1676
rect 1422 1671 1428 1672
rect 1502 1676 1508 1677
rect 1502 1672 1503 1676
rect 1507 1672 1508 1676
rect 1502 1671 1508 1672
rect 1582 1676 1588 1677
rect 1582 1672 1583 1676
rect 1587 1672 1588 1676
rect 1582 1671 1588 1672
rect 1662 1676 1668 1677
rect 1662 1672 1663 1676
rect 1667 1672 1668 1676
rect 1662 1671 1668 1672
rect 1734 1676 1740 1677
rect 1734 1672 1735 1676
rect 1739 1672 1740 1676
rect 1734 1671 1740 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1870 1676 1876 1677
rect 1870 1672 1871 1676
rect 1875 1672 1876 1676
rect 1870 1671 1876 1672
rect 1934 1676 1940 1677
rect 1934 1672 1935 1676
rect 1939 1672 1940 1676
rect 1934 1671 1940 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2062 1676 2068 1677
rect 2062 1672 2063 1676
rect 2067 1672 2068 1676
rect 2062 1671 2068 1672
rect 1302 1664 1308 1665
rect 1302 1660 1303 1664
rect 1307 1660 1308 1664
rect 1302 1659 1308 1660
rect 1358 1664 1364 1665
rect 1358 1660 1359 1664
rect 1363 1660 1364 1664
rect 1358 1659 1364 1660
rect 1446 1664 1452 1665
rect 1446 1660 1447 1664
rect 1451 1660 1452 1664
rect 1446 1659 1452 1660
rect 1542 1664 1548 1665
rect 1542 1660 1543 1664
rect 1547 1660 1548 1664
rect 1542 1659 1548 1660
rect 1638 1664 1644 1665
rect 1638 1660 1639 1664
rect 1643 1660 1644 1664
rect 1638 1659 1644 1660
rect 1726 1664 1732 1665
rect 1726 1660 1727 1664
rect 1731 1660 1732 1664
rect 1726 1659 1732 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1894 1664 1900 1665
rect 1894 1660 1895 1664
rect 1899 1660 1900 1664
rect 1894 1659 1900 1660
rect 1966 1664 1972 1665
rect 1966 1660 1967 1664
rect 1971 1660 1972 1664
rect 1966 1659 1972 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2094 1664 2100 1665
rect 2094 1660 2095 1664
rect 2099 1660 2100 1664
rect 2094 1659 2100 1660
rect 2158 1664 2164 1665
rect 2158 1660 2159 1664
rect 2163 1660 2164 1664
rect 2158 1659 2164 1660
rect 2222 1664 2228 1665
rect 2222 1660 2223 1664
rect 2227 1660 2228 1664
rect 2222 1659 2228 1660
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 174 1657 180 1658
rect 174 1653 175 1657
rect 179 1653 180 1657
rect 174 1652 180 1653
rect 238 1657 244 1658
rect 238 1653 239 1657
rect 243 1653 244 1657
rect 238 1652 244 1653
rect 318 1657 324 1658
rect 318 1653 319 1657
rect 323 1653 324 1657
rect 318 1652 324 1653
rect 414 1657 420 1658
rect 414 1653 415 1657
rect 419 1653 420 1657
rect 414 1652 420 1653
rect 510 1657 516 1658
rect 510 1653 511 1657
rect 515 1653 516 1657
rect 510 1652 516 1653
rect 614 1657 620 1658
rect 614 1653 615 1657
rect 619 1653 620 1657
rect 614 1652 620 1653
rect 710 1657 716 1658
rect 710 1653 711 1657
rect 715 1653 716 1657
rect 710 1652 716 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 878 1657 884 1658
rect 878 1653 879 1657
rect 883 1653 884 1657
rect 878 1652 884 1653
rect 950 1657 956 1658
rect 950 1653 951 1657
rect 955 1653 956 1657
rect 950 1652 956 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1086 1657 1092 1658
rect 1086 1653 1087 1657
rect 1091 1653 1092 1657
rect 1086 1652 1092 1653
rect 1158 1657 1164 1658
rect 1158 1653 1159 1657
rect 1163 1653 1164 1657
rect 1158 1652 1164 1653
rect 1278 1657 1284 1658
rect 1278 1653 1279 1657
rect 1283 1653 1284 1657
rect 1278 1652 1284 1653
rect 2406 1657 2412 1658
rect 2406 1653 2407 1657
rect 2411 1653 2412 1657
rect 2406 1652 2412 1653
rect 1278 1640 1284 1641
rect 1278 1636 1279 1640
rect 1283 1636 1284 1640
rect 1278 1635 1284 1636
rect 2406 1640 2412 1641
rect 2406 1636 2407 1640
rect 2411 1636 2412 1640
rect 2406 1635 2412 1636
rect 270 1623 276 1624
rect 270 1619 271 1623
rect 275 1619 276 1623
rect 270 1618 276 1619
rect 310 1623 316 1624
rect 310 1619 311 1623
rect 315 1619 316 1623
rect 310 1618 316 1619
rect 358 1623 364 1624
rect 358 1619 359 1623
rect 363 1619 364 1623
rect 358 1618 364 1619
rect 414 1623 420 1624
rect 414 1619 415 1623
rect 419 1619 420 1623
rect 414 1618 420 1619
rect 470 1623 476 1624
rect 470 1619 471 1623
rect 475 1619 476 1623
rect 470 1618 476 1619
rect 534 1623 540 1624
rect 534 1619 535 1623
rect 539 1619 540 1623
rect 534 1618 540 1619
rect 598 1623 604 1624
rect 598 1619 599 1623
rect 603 1619 604 1623
rect 598 1618 604 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 718 1623 724 1624
rect 718 1619 719 1623
rect 723 1619 724 1623
rect 718 1618 724 1619
rect 774 1623 780 1624
rect 774 1619 775 1623
rect 779 1619 780 1623
rect 774 1618 780 1619
rect 830 1623 836 1624
rect 830 1619 831 1623
rect 835 1619 836 1623
rect 830 1618 836 1619
rect 886 1623 892 1624
rect 886 1619 887 1623
rect 891 1619 892 1623
rect 886 1618 892 1619
rect 942 1623 948 1624
rect 942 1619 943 1623
rect 947 1619 948 1623
rect 942 1618 948 1619
rect 998 1623 1004 1624
rect 998 1619 999 1623
rect 1003 1619 1004 1623
rect 998 1618 1004 1619
rect 1302 1617 1308 1618
rect 1302 1613 1303 1617
rect 1307 1613 1308 1617
rect 1302 1612 1308 1613
rect 1358 1617 1364 1618
rect 1358 1613 1359 1617
rect 1363 1613 1364 1617
rect 1358 1612 1364 1613
rect 1446 1617 1452 1618
rect 1446 1613 1447 1617
rect 1451 1613 1452 1617
rect 1446 1612 1452 1613
rect 1542 1617 1548 1618
rect 1542 1613 1543 1617
rect 1547 1613 1548 1617
rect 1542 1612 1548 1613
rect 1638 1617 1644 1618
rect 1638 1613 1639 1617
rect 1643 1613 1644 1617
rect 1638 1612 1644 1613
rect 1726 1617 1732 1618
rect 1726 1613 1727 1617
rect 1731 1613 1732 1617
rect 1726 1612 1732 1613
rect 1814 1617 1820 1618
rect 1814 1613 1815 1617
rect 1819 1613 1820 1617
rect 1814 1612 1820 1613
rect 1894 1617 1900 1618
rect 1894 1613 1895 1617
rect 1899 1613 1900 1617
rect 1894 1612 1900 1613
rect 1966 1617 1972 1618
rect 1966 1613 1967 1617
rect 1971 1613 1972 1617
rect 1966 1612 1972 1613
rect 2030 1617 2036 1618
rect 2030 1613 2031 1617
rect 2035 1613 2036 1617
rect 2030 1612 2036 1613
rect 2094 1617 2100 1618
rect 2094 1613 2095 1617
rect 2099 1613 2100 1617
rect 2094 1612 2100 1613
rect 2158 1617 2164 1618
rect 2158 1613 2159 1617
rect 2163 1613 2164 1617
rect 2158 1612 2164 1613
rect 2222 1617 2228 1618
rect 2222 1613 2223 1617
rect 2227 1613 2228 1617
rect 2222 1612 2228 1613
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 110 1595 116 1596
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 1238 1595 1244 1596
rect 1326 1587 1332 1588
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 110 1578 116 1579
rect 1238 1583 1244 1584
rect 1238 1579 1239 1583
rect 1243 1579 1244 1583
rect 1326 1583 1327 1587
rect 1331 1583 1332 1587
rect 1326 1582 1332 1583
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1583 1404 1587
rect 1398 1582 1404 1583
rect 1478 1587 1484 1588
rect 1478 1583 1479 1587
rect 1483 1583 1484 1587
rect 1478 1582 1484 1583
rect 1566 1587 1572 1588
rect 1566 1583 1567 1587
rect 1571 1583 1572 1587
rect 1566 1582 1572 1583
rect 1654 1587 1660 1588
rect 1654 1583 1655 1587
rect 1659 1583 1660 1587
rect 1654 1582 1660 1583
rect 1742 1587 1748 1588
rect 1742 1583 1743 1587
rect 1747 1583 1748 1587
rect 1742 1582 1748 1583
rect 1830 1587 1836 1588
rect 1830 1583 1831 1587
rect 1835 1583 1836 1587
rect 1830 1582 1836 1583
rect 1910 1587 1916 1588
rect 1910 1583 1911 1587
rect 1915 1583 1916 1587
rect 1910 1582 1916 1583
rect 1982 1587 1988 1588
rect 1982 1583 1983 1587
rect 1987 1583 1988 1587
rect 1982 1582 1988 1583
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 2046 1582 2052 1583
rect 2110 1587 2116 1588
rect 2110 1583 2111 1587
rect 2115 1583 2116 1587
rect 2110 1582 2116 1583
rect 2166 1587 2172 1588
rect 2166 1583 2167 1587
rect 2171 1583 2172 1587
rect 2166 1582 2172 1583
rect 2214 1587 2220 1588
rect 2214 1583 2215 1587
rect 2219 1583 2220 1587
rect 2214 1582 2220 1583
rect 2270 1587 2276 1588
rect 2270 1583 2271 1587
rect 2275 1583 2276 1587
rect 2270 1582 2276 1583
rect 2318 1587 2324 1588
rect 2318 1583 2319 1587
rect 2323 1583 2324 1587
rect 2318 1582 2324 1583
rect 2358 1587 2364 1588
rect 2358 1583 2359 1587
rect 2363 1583 2364 1587
rect 2358 1582 2364 1583
rect 1238 1578 1244 1579
rect 270 1576 276 1577
rect 270 1572 271 1576
rect 275 1572 276 1576
rect 270 1571 276 1572
rect 310 1576 316 1577
rect 310 1572 311 1576
rect 315 1572 316 1576
rect 310 1571 316 1572
rect 358 1576 364 1577
rect 358 1572 359 1576
rect 363 1572 364 1576
rect 358 1571 364 1572
rect 414 1576 420 1577
rect 414 1572 415 1576
rect 419 1572 420 1576
rect 414 1571 420 1572
rect 470 1576 476 1577
rect 470 1572 471 1576
rect 475 1572 476 1576
rect 470 1571 476 1572
rect 534 1576 540 1577
rect 534 1572 535 1576
rect 539 1572 540 1576
rect 534 1571 540 1572
rect 598 1576 604 1577
rect 598 1572 599 1576
rect 603 1572 604 1576
rect 598 1571 604 1572
rect 662 1576 668 1577
rect 662 1572 663 1576
rect 667 1572 668 1576
rect 662 1571 668 1572
rect 718 1576 724 1577
rect 718 1572 719 1576
rect 723 1572 724 1576
rect 718 1571 724 1572
rect 774 1576 780 1577
rect 774 1572 775 1576
rect 779 1572 780 1576
rect 774 1571 780 1572
rect 830 1576 836 1577
rect 830 1572 831 1576
rect 835 1572 836 1576
rect 830 1571 836 1572
rect 886 1576 892 1577
rect 886 1572 887 1576
rect 891 1572 892 1576
rect 886 1571 892 1572
rect 942 1576 948 1577
rect 942 1572 943 1576
rect 947 1572 948 1576
rect 942 1571 948 1572
rect 998 1576 1004 1577
rect 998 1572 999 1576
rect 1003 1572 1004 1576
rect 998 1571 1004 1572
rect 1278 1564 1284 1565
rect 1278 1560 1279 1564
rect 1283 1560 1284 1564
rect 1278 1559 1284 1560
rect 2406 1564 2412 1565
rect 2406 1560 2407 1564
rect 2411 1560 2412 1564
rect 2406 1559 2412 1560
rect 326 1556 332 1557
rect 326 1552 327 1556
rect 331 1552 332 1556
rect 326 1551 332 1552
rect 366 1556 372 1557
rect 366 1552 367 1556
rect 371 1552 372 1556
rect 366 1551 372 1552
rect 406 1556 412 1557
rect 406 1552 407 1556
rect 411 1552 412 1556
rect 406 1551 412 1552
rect 446 1556 452 1557
rect 446 1552 447 1556
rect 451 1552 452 1556
rect 446 1551 452 1552
rect 486 1556 492 1557
rect 486 1552 487 1556
rect 491 1552 492 1556
rect 486 1551 492 1552
rect 526 1556 532 1557
rect 526 1552 527 1556
rect 531 1552 532 1556
rect 526 1551 532 1552
rect 566 1556 572 1557
rect 566 1552 567 1556
rect 571 1552 572 1556
rect 566 1551 572 1552
rect 606 1556 612 1557
rect 606 1552 607 1556
rect 611 1552 612 1556
rect 606 1551 612 1552
rect 646 1556 652 1557
rect 646 1552 647 1556
rect 651 1552 652 1556
rect 646 1551 652 1552
rect 686 1556 692 1557
rect 686 1552 687 1556
rect 691 1552 692 1556
rect 686 1551 692 1552
rect 726 1556 732 1557
rect 726 1552 727 1556
rect 731 1552 732 1556
rect 726 1551 732 1552
rect 766 1556 772 1557
rect 766 1552 767 1556
rect 771 1552 772 1556
rect 766 1551 772 1552
rect 806 1556 812 1557
rect 806 1552 807 1556
rect 811 1552 812 1556
rect 806 1551 812 1552
rect 846 1556 852 1557
rect 846 1552 847 1556
rect 851 1552 852 1556
rect 846 1551 852 1552
rect 886 1556 892 1557
rect 886 1552 887 1556
rect 891 1552 892 1556
rect 886 1551 892 1552
rect 926 1556 932 1557
rect 926 1552 927 1556
rect 931 1552 932 1556
rect 926 1551 932 1552
rect 110 1549 116 1550
rect 110 1545 111 1549
rect 115 1545 116 1549
rect 110 1544 116 1545
rect 1238 1549 1244 1550
rect 1238 1545 1239 1549
rect 1243 1545 1244 1549
rect 1238 1544 1244 1545
rect 1278 1547 1284 1548
rect 1278 1543 1279 1547
rect 1283 1543 1284 1547
rect 1278 1542 1284 1543
rect 2406 1547 2412 1548
rect 2406 1543 2407 1547
rect 2411 1543 2412 1547
rect 2406 1542 2412 1543
rect 1326 1540 1332 1541
rect 1326 1536 1327 1540
rect 1331 1536 1332 1540
rect 1326 1535 1332 1536
rect 1398 1540 1404 1541
rect 1398 1536 1399 1540
rect 1403 1536 1404 1540
rect 1398 1535 1404 1536
rect 1478 1540 1484 1541
rect 1478 1536 1479 1540
rect 1483 1536 1484 1540
rect 1478 1535 1484 1536
rect 1566 1540 1572 1541
rect 1566 1536 1567 1540
rect 1571 1536 1572 1540
rect 1566 1535 1572 1536
rect 1654 1540 1660 1541
rect 1654 1536 1655 1540
rect 1659 1536 1660 1540
rect 1654 1535 1660 1536
rect 1742 1540 1748 1541
rect 1742 1536 1743 1540
rect 1747 1536 1748 1540
rect 1742 1535 1748 1536
rect 1830 1540 1836 1541
rect 1830 1536 1831 1540
rect 1835 1536 1836 1540
rect 1830 1535 1836 1536
rect 1910 1540 1916 1541
rect 1910 1536 1911 1540
rect 1915 1536 1916 1540
rect 1910 1535 1916 1536
rect 1982 1540 1988 1541
rect 1982 1536 1983 1540
rect 1987 1536 1988 1540
rect 1982 1535 1988 1536
rect 2046 1540 2052 1541
rect 2046 1536 2047 1540
rect 2051 1536 2052 1540
rect 2046 1535 2052 1536
rect 2110 1540 2116 1541
rect 2110 1536 2111 1540
rect 2115 1536 2116 1540
rect 2110 1535 2116 1536
rect 2166 1540 2172 1541
rect 2166 1536 2167 1540
rect 2171 1536 2172 1540
rect 2166 1535 2172 1536
rect 2214 1540 2220 1541
rect 2214 1536 2215 1540
rect 2219 1536 2220 1540
rect 2214 1535 2220 1536
rect 2270 1540 2276 1541
rect 2270 1536 2271 1540
rect 2275 1536 2276 1540
rect 2270 1535 2276 1536
rect 2318 1540 2324 1541
rect 2318 1536 2319 1540
rect 2323 1536 2324 1540
rect 2318 1535 2324 1536
rect 2358 1540 2364 1541
rect 2358 1536 2359 1540
rect 2363 1536 2364 1540
rect 2358 1535 2364 1536
rect 110 1532 116 1533
rect 110 1528 111 1532
rect 115 1528 116 1532
rect 110 1527 116 1528
rect 1238 1532 1244 1533
rect 1238 1528 1239 1532
rect 1243 1528 1244 1532
rect 1238 1527 1244 1528
rect 1334 1524 1340 1525
rect 1334 1520 1335 1524
rect 1339 1520 1340 1524
rect 1334 1519 1340 1520
rect 1414 1524 1420 1525
rect 1414 1520 1415 1524
rect 1419 1520 1420 1524
rect 1414 1519 1420 1520
rect 1502 1524 1508 1525
rect 1502 1520 1503 1524
rect 1507 1520 1508 1524
rect 1502 1519 1508 1520
rect 1614 1524 1620 1525
rect 1614 1520 1615 1524
rect 1619 1520 1620 1524
rect 1614 1519 1620 1520
rect 1742 1524 1748 1525
rect 1742 1520 1743 1524
rect 1747 1520 1748 1524
rect 1742 1519 1748 1520
rect 1886 1524 1892 1525
rect 1886 1520 1887 1524
rect 1891 1520 1892 1524
rect 1886 1519 1892 1520
rect 2046 1524 2052 1525
rect 2046 1520 2047 1524
rect 2051 1520 2052 1524
rect 2046 1519 2052 1520
rect 2214 1524 2220 1525
rect 2214 1520 2215 1524
rect 2219 1520 2220 1524
rect 2214 1519 2220 1520
rect 2358 1524 2364 1525
rect 2358 1520 2359 1524
rect 2363 1520 2364 1524
rect 2358 1519 2364 1520
rect 1278 1517 1284 1518
rect 1278 1513 1279 1517
rect 1283 1513 1284 1517
rect 1278 1512 1284 1513
rect 2406 1517 2412 1518
rect 2406 1513 2407 1517
rect 2411 1513 2412 1517
rect 2406 1512 2412 1513
rect 326 1509 332 1510
rect 326 1505 327 1509
rect 331 1505 332 1509
rect 326 1504 332 1505
rect 366 1509 372 1510
rect 366 1505 367 1509
rect 371 1505 372 1509
rect 366 1504 372 1505
rect 406 1509 412 1510
rect 406 1505 407 1509
rect 411 1505 412 1509
rect 406 1504 412 1505
rect 446 1509 452 1510
rect 446 1505 447 1509
rect 451 1505 452 1509
rect 446 1504 452 1505
rect 486 1509 492 1510
rect 486 1505 487 1509
rect 491 1505 492 1509
rect 486 1504 492 1505
rect 526 1509 532 1510
rect 526 1505 527 1509
rect 531 1505 532 1509
rect 526 1504 532 1505
rect 566 1509 572 1510
rect 566 1505 567 1509
rect 571 1505 572 1509
rect 566 1504 572 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 646 1509 652 1510
rect 646 1505 647 1509
rect 651 1505 652 1509
rect 646 1504 652 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 726 1509 732 1510
rect 726 1505 727 1509
rect 731 1505 732 1509
rect 726 1504 732 1505
rect 766 1509 772 1510
rect 766 1505 767 1509
rect 771 1505 772 1509
rect 766 1504 772 1505
rect 806 1509 812 1510
rect 806 1505 807 1509
rect 811 1505 812 1509
rect 806 1504 812 1505
rect 846 1509 852 1510
rect 846 1505 847 1509
rect 851 1505 852 1509
rect 846 1504 852 1505
rect 886 1509 892 1510
rect 886 1505 887 1509
rect 891 1505 892 1509
rect 886 1504 892 1505
rect 926 1509 932 1510
rect 926 1505 927 1509
rect 931 1505 932 1509
rect 926 1504 932 1505
rect 1278 1500 1284 1501
rect 1278 1496 1279 1500
rect 1283 1496 1284 1500
rect 1278 1495 1284 1496
rect 2406 1500 2412 1501
rect 2406 1496 2407 1500
rect 2411 1496 2412 1500
rect 2406 1495 2412 1496
rect 1334 1477 1340 1478
rect 1334 1473 1335 1477
rect 1339 1473 1340 1477
rect 1334 1472 1340 1473
rect 1414 1477 1420 1478
rect 1414 1473 1415 1477
rect 1419 1473 1420 1477
rect 1414 1472 1420 1473
rect 1502 1477 1508 1478
rect 1502 1473 1503 1477
rect 1507 1473 1508 1477
rect 1502 1472 1508 1473
rect 1614 1477 1620 1478
rect 1614 1473 1615 1477
rect 1619 1473 1620 1477
rect 1614 1472 1620 1473
rect 1742 1477 1748 1478
rect 1742 1473 1743 1477
rect 1747 1473 1748 1477
rect 1742 1472 1748 1473
rect 1886 1477 1892 1478
rect 1886 1473 1887 1477
rect 1891 1473 1892 1477
rect 1886 1472 1892 1473
rect 2046 1477 2052 1478
rect 2046 1473 2047 1477
rect 2051 1473 2052 1477
rect 2046 1472 2052 1473
rect 2214 1477 2220 1478
rect 2214 1473 2215 1477
rect 2219 1473 2220 1477
rect 2214 1472 2220 1473
rect 2358 1477 2364 1478
rect 2358 1473 2359 1477
rect 2363 1473 2364 1477
rect 2358 1472 2364 1473
rect 1374 1447 1380 1448
rect 1374 1443 1375 1447
rect 1379 1443 1380 1447
rect 1374 1442 1380 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1550 1447 1556 1448
rect 1550 1443 1551 1447
rect 1555 1443 1556 1447
rect 1550 1442 1556 1443
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1726 1447 1732 1448
rect 1726 1443 1727 1447
rect 1731 1443 1732 1447
rect 1726 1442 1732 1443
rect 1806 1447 1812 1448
rect 1806 1443 1807 1447
rect 1811 1443 1812 1447
rect 1806 1442 1812 1443
rect 1878 1447 1884 1448
rect 1878 1443 1879 1447
rect 1883 1443 1884 1447
rect 1878 1442 1884 1443
rect 1942 1447 1948 1448
rect 1942 1443 1943 1447
rect 1947 1443 1948 1447
rect 1942 1442 1948 1443
rect 1998 1447 2004 1448
rect 1998 1443 1999 1447
rect 2003 1443 2004 1447
rect 1998 1442 2004 1443
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2046 1442 2052 1443
rect 2094 1447 2100 1448
rect 2094 1443 2095 1447
rect 2099 1443 2100 1447
rect 2094 1442 2100 1443
rect 2142 1447 2148 1448
rect 2142 1443 2143 1447
rect 2147 1443 2148 1447
rect 2142 1442 2148 1443
rect 2190 1447 2196 1448
rect 2190 1443 2191 1447
rect 2195 1443 2196 1447
rect 2190 1442 2196 1443
rect 2238 1447 2244 1448
rect 2238 1443 2239 1447
rect 2243 1443 2244 1447
rect 2238 1442 2244 1443
rect 2278 1447 2284 1448
rect 2278 1443 2279 1447
rect 2283 1443 2284 1447
rect 2278 1442 2284 1443
rect 2318 1447 2324 1448
rect 2318 1443 2319 1447
rect 2323 1443 2324 1447
rect 2318 1442 2324 1443
rect 2358 1447 2364 1448
rect 2358 1443 2359 1447
rect 2363 1443 2364 1447
rect 2358 1442 2364 1443
rect 142 1439 148 1440
rect 142 1435 143 1439
rect 147 1435 148 1439
rect 142 1434 148 1435
rect 182 1439 188 1440
rect 182 1435 183 1439
rect 187 1435 188 1439
rect 182 1434 188 1435
rect 222 1439 228 1440
rect 222 1435 223 1439
rect 227 1435 228 1439
rect 222 1434 228 1435
rect 262 1439 268 1440
rect 262 1435 263 1439
rect 267 1435 268 1439
rect 262 1434 268 1435
rect 318 1439 324 1440
rect 318 1435 319 1439
rect 323 1435 324 1439
rect 318 1434 324 1435
rect 390 1439 396 1440
rect 390 1435 391 1439
rect 395 1435 396 1439
rect 390 1434 396 1435
rect 470 1439 476 1440
rect 470 1435 471 1439
rect 475 1435 476 1439
rect 470 1434 476 1435
rect 558 1439 564 1440
rect 558 1435 559 1439
rect 563 1435 564 1439
rect 558 1434 564 1435
rect 646 1439 652 1440
rect 646 1435 647 1439
rect 651 1435 652 1439
rect 646 1434 652 1435
rect 726 1439 732 1440
rect 726 1435 727 1439
rect 731 1435 732 1439
rect 726 1434 732 1435
rect 806 1439 812 1440
rect 806 1435 807 1439
rect 811 1435 812 1439
rect 806 1434 812 1435
rect 878 1439 884 1440
rect 878 1435 879 1439
rect 883 1435 884 1439
rect 878 1434 884 1435
rect 942 1439 948 1440
rect 942 1435 943 1439
rect 947 1435 948 1439
rect 942 1434 948 1435
rect 998 1439 1004 1440
rect 998 1435 999 1439
rect 1003 1435 1004 1439
rect 998 1434 1004 1435
rect 1046 1439 1052 1440
rect 1046 1435 1047 1439
rect 1051 1435 1052 1439
rect 1046 1434 1052 1435
rect 1102 1439 1108 1440
rect 1102 1435 1103 1439
rect 1107 1435 1108 1439
rect 1102 1434 1108 1435
rect 1150 1439 1156 1440
rect 1150 1435 1151 1439
rect 1155 1435 1156 1439
rect 1150 1434 1156 1435
rect 1190 1439 1196 1440
rect 1190 1435 1191 1439
rect 1195 1435 1196 1439
rect 1190 1434 1196 1435
rect 1278 1424 1284 1425
rect 1278 1420 1279 1424
rect 1283 1420 1284 1424
rect 1278 1419 1284 1420
rect 2406 1424 2412 1425
rect 2406 1420 2407 1424
rect 2411 1420 2412 1424
rect 2406 1419 2412 1420
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1238 1416 1244 1417
rect 1238 1412 1239 1416
rect 1243 1412 1244 1416
rect 1238 1411 1244 1412
rect 1278 1407 1284 1408
rect 1278 1403 1279 1407
rect 1283 1403 1284 1407
rect 1278 1402 1284 1403
rect 2406 1407 2412 1408
rect 2406 1403 2407 1407
rect 2411 1403 2412 1407
rect 2406 1402 2412 1403
rect 1374 1400 1380 1401
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 1238 1399 1244 1400
rect 1238 1395 1239 1399
rect 1243 1395 1244 1399
rect 1374 1396 1375 1400
rect 1379 1396 1380 1400
rect 1374 1395 1380 1396
rect 1462 1400 1468 1401
rect 1462 1396 1463 1400
rect 1467 1396 1468 1400
rect 1462 1395 1468 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1806 1400 1812 1401
rect 1806 1396 1807 1400
rect 1811 1396 1812 1400
rect 1806 1395 1812 1396
rect 1878 1400 1884 1401
rect 1878 1396 1879 1400
rect 1883 1396 1884 1400
rect 1878 1395 1884 1396
rect 1942 1400 1948 1401
rect 1942 1396 1943 1400
rect 1947 1396 1948 1400
rect 1942 1395 1948 1396
rect 1998 1400 2004 1401
rect 1998 1396 1999 1400
rect 2003 1396 2004 1400
rect 1998 1395 2004 1396
rect 2046 1400 2052 1401
rect 2046 1396 2047 1400
rect 2051 1396 2052 1400
rect 2046 1395 2052 1396
rect 2094 1400 2100 1401
rect 2094 1396 2095 1400
rect 2099 1396 2100 1400
rect 2094 1395 2100 1396
rect 2142 1400 2148 1401
rect 2142 1396 2143 1400
rect 2147 1396 2148 1400
rect 2142 1395 2148 1396
rect 2190 1400 2196 1401
rect 2190 1396 2191 1400
rect 2195 1396 2196 1400
rect 2190 1395 2196 1396
rect 2238 1400 2244 1401
rect 2238 1396 2239 1400
rect 2243 1396 2244 1400
rect 2238 1395 2244 1396
rect 2278 1400 2284 1401
rect 2278 1396 2279 1400
rect 2283 1396 2284 1400
rect 2278 1395 2284 1396
rect 2318 1400 2324 1401
rect 2318 1396 2319 1400
rect 2323 1396 2324 1400
rect 2318 1395 2324 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 1238 1394 1244 1395
rect 142 1392 148 1393
rect 142 1388 143 1392
rect 147 1388 148 1392
rect 142 1387 148 1388
rect 182 1392 188 1393
rect 182 1388 183 1392
rect 187 1388 188 1392
rect 182 1387 188 1388
rect 222 1392 228 1393
rect 222 1388 223 1392
rect 227 1388 228 1392
rect 222 1387 228 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 318 1392 324 1393
rect 318 1388 319 1392
rect 323 1388 324 1392
rect 318 1387 324 1388
rect 390 1392 396 1393
rect 390 1388 391 1392
rect 395 1388 396 1392
rect 390 1387 396 1388
rect 470 1392 476 1393
rect 470 1388 471 1392
rect 475 1388 476 1392
rect 470 1387 476 1388
rect 558 1392 564 1393
rect 558 1388 559 1392
rect 563 1388 564 1392
rect 558 1387 564 1388
rect 646 1392 652 1393
rect 646 1388 647 1392
rect 651 1388 652 1392
rect 646 1387 652 1388
rect 726 1392 732 1393
rect 726 1388 727 1392
rect 731 1388 732 1392
rect 726 1387 732 1388
rect 806 1392 812 1393
rect 806 1388 807 1392
rect 811 1388 812 1392
rect 806 1387 812 1388
rect 878 1392 884 1393
rect 878 1388 879 1392
rect 883 1388 884 1392
rect 878 1387 884 1388
rect 942 1392 948 1393
rect 942 1388 943 1392
rect 947 1388 948 1392
rect 942 1387 948 1388
rect 998 1392 1004 1393
rect 998 1388 999 1392
rect 1003 1388 1004 1392
rect 998 1387 1004 1388
rect 1046 1392 1052 1393
rect 1046 1388 1047 1392
rect 1051 1388 1052 1392
rect 1046 1387 1052 1388
rect 1102 1392 1108 1393
rect 1102 1388 1103 1392
rect 1107 1388 1108 1392
rect 1102 1387 1108 1388
rect 1150 1392 1156 1393
rect 1150 1388 1151 1392
rect 1155 1388 1156 1392
rect 1150 1387 1156 1388
rect 1190 1392 1196 1393
rect 1190 1388 1191 1392
rect 1195 1388 1196 1392
rect 1190 1387 1196 1388
rect 166 1380 172 1381
rect 166 1376 167 1380
rect 171 1376 172 1380
rect 166 1375 172 1376
rect 206 1380 212 1381
rect 206 1376 207 1380
rect 211 1376 212 1380
rect 206 1375 212 1376
rect 246 1380 252 1381
rect 246 1376 247 1380
rect 251 1376 252 1380
rect 246 1375 252 1376
rect 302 1380 308 1381
rect 302 1376 303 1380
rect 307 1376 308 1380
rect 302 1375 308 1376
rect 366 1380 372 1381
rect 366 1376 367 1380
rect 371 1376 372 1380
rect 366 1375 372 1376
rect 438 1380 444 1381
rect 438 1376 439 1380
rect 443 1376 444 1380
rect 438 1375 444 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 598 1380 604 1381
rect 598 1376 599 1380
rect 603 1376 604 1380
rect 598 1375 604 1376
rect 678 1380 684 1381
rect 678 1376 679 1380
rect 683 1376 684 1380
rect 678 1375 684 1376
rect 750 1380 756 1381
rect 750 1376 751 1380
rect 755 1376 756 1380
rect 750 1375 756 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 886 1380 892 1381
rect 886 1376 887 1380
rect 891 1376 892 1380
rect 886 1375 892 1376
rect 950 1380 956 1381
rect 950 1376 951 1380
rect 955 1376 956 1380
rect 950 1375 956 1376
rect 1014 1380 1020 1381
rect 1014 1376 1015 1380
rect 1019 1376 1020 1380
rect 1014 1375 1020 1376
rect 1078 1380 1084 1381
rect 1078 1376 1079 1380
rect 1083 1376 1084 1380
rect 1078 1375 1084 1376
rect 1142 1380 1148 1381
rect 1142 1376 1143 1380
rect 1147 1376 1148 1380
rect 1142 1375 1148 1376
rect 1190 1380 1196 1381
rect 1190 1376 1191 1380
rect 1195 1376 1196 1380
rect 1190 1375 1196 1376
rect 1302 1380 1308 1381
rect 1302 1376 1303 1380
rect 1307 1376 1308 1380
rect 1302 1375 1308 1376
rect 1342 1380 1348 1381
rect 1342 1376 1343 1380
rect 1347 1376 1348 1380
rect 1342 1375 1348 1376
rect 1398 1380 1404 1381
rect 1398 1376 1399 1380
rect 1403 1376 1404 1380
rect 1398 1375 1404 1376
rect 1462 1380 1468 1381
rect 1462 1376 1463 1380
rect 1467 1376 1468 1380
rect 1462 1375 1468 1376
rect 1534 1380 1540 1381
rect 1534 1376 1535 1380
rect 1539 1376 1540 1380
rect 1534 1375 1540 1376
rect 1606 1380 1612 1381
rect 1606 1376 1607 1380
rect 1611 1376 1612 1380
rect 1606 1375 1612 1376
rect 1686 1380 1692 1381
rect 1686 1376 1687 1380
rect 1691 1376 1692 1380
rect 1686 1375 1692 1376
rect 1766 1380 1772 1381
rect 1766 1376 1767 1380
rect 1771 1376 1772 1380
rect 1766 1375 1772 1376
rect 1846 1380 1852 1381
rect 1846 1376 1847 1380
rect 1851 1376 1852 1380
rect 1846 1375 1852 1376
rect 1934 1380 1940 1381
rect 1934 1376 1935 1380
rect 1939 1376 1940 1380
rect 1934 1375 1940 1376
rect 2022 1380 2028 1381
rect 2022 1376 2023 1380
rect 2027 1376 2028 1380
rect 2022 1375 2028 1376
rect 2110 1380 2116 1381
rect 2110 1376 2111 1380
rect 2115 1376 2116 1380
rect 2110 1375 2116 1376
rect 2198 1380 2204 1381
rect 2198 1376 2199 1380
rect 2203 1376 2204 1380
rect 2198 1375 2204 1376
rect 2286 1380 2292 1381
rect 2286 1376 2287 1380
rect 2291 1376 2292 1380
rect 2286 1375 2292 1376
rect 2358 1380 2364 1381
rect 2358 1376 2359 1380
rect 2363 1376 2364 1380
rect 2358 1375 2364 1376
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1278 1373 1284 1374
rect 1278 1369 1279 1373
rect 1283 1369 1284 1373
rect 1278 1368 1284 1369
rect 2406 1373 2412 1374
rect 2406 1369 2407 1373
rect 2411 1369 2412 1373
rect 2406 1368 2412 1369
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 110 1351 116 1352
rect 1238 1356 1244 1357
rect 1238 1352 1239 1356
rect 1243 1352 1244 1356
rect 1238 1351 1244 1352
rect 1278 1356 1284 1357
rect 1278 1352 1279 1356
rect 1283 1352 1284 1356
rect 1278 1351 1284 1352
rect 2406 1356 2412 1357
rect 2406 1352 2407 1356
rect 2411 1352 2412 1356
rect 2406 1351 2412 1352
rect 166 1333 172 1334
rect 166 1329 167 1333
rect 171 1329 172 1333
rect 166 1328 172 1329
rect 206 1333 212 1334
rect 206 1329 207 1333
rect 211 1329 212 1333
rect 206 1328 212 1329
rect 246 1333 252 1334
rect 246 1329 247 1333
rect 251 1329 252 1333
rect 246 1328 252 1329
rect 302 1333 308 1334
rect 302 1329 303 1333
rect 307 1329 308 1333
rect 302 1328 308 1329
rect 366 1333 372 1334
rect 366 1329 367 1333
rect 371 1329 372 1333
rect 366 1328 372 1329
rect 438 1333 444 1334
rect 438 1329 439 1333
rect 443 1329 444 1333
rect 438 1328 444 1329
rect 518 1333 524 1334
rect 518 1329 519 1333
rect 523 1329 524 1333
rect 518 1328 524 1329
rect 598 1333 604 1334
rect 598 1329 599 1333
rect 603 1329 604 1333
rect 598 1328 604 1329
rect 678 1333 684 1334
rect 678 1329 679 1333
rect 683 1329 684 1333
rect 678 1328 684 1329
rect 750 1333 756 1334
rect 750 1329 751 1333
rect 755 1329 756 1333
rect 750 1328 756 1329
rect 822 1333 828 1334
rect 822 1329 823 1333
rect 827 1329 828 1333
rect 822 1328 828 1329
rect 886 1333 892 1334
rect 886 1329 887 1333
rect 891 1329 892 1333
rect 886 1328 892 1329
rect 950 1333 956 1334
rect 950 1329 951 1333
rect 955 1329 956 1333
rect 950 1328 956 1329
rect 1014 1333 1020 1334
rect 1014 1329 1015 1333
rect 1019 1329 1020 1333
rect 1014 1328 1020 1329
rect 1078 1333 1084 1334
rect 1078 1329 1079 1333
rect 1083 1329 1084 1333
rect 1078 1328 1084 1329
rect 1142 1333 1148 1334
rect 1142 1329 1143 1333
rect 1147 1329 1148 1333
rect 1142 1328 1148 1329
rect 1190 1333 1196 1334
rect 1190 1329 1191 1333
rect 1195 1329 1196 1333
rect 1190 1328 1196 1329
rect 1302 1333 1308 1334
rect 1302 1329 1303 1333
rect 1307 1329 1308 1333
rect 1302 1328 1308 1329
rect 1342 1333 1348 1334
rect 1342 1329 1343 1333
rect 1347 1329 1348 1333
rect 1342 1328 1348 1329
rect 1398 1333 1404 1334
rect 1398 1329 1399 1333
rect 1403 1329 1404 1333
rect 1398 1328 1404 1329
rect 1462 1333 1468 1334
rect 1462 1329 1463 1333
rect 1467 1329 1468 1333
rect 1462 1328 1468 1329
rect 1534 1333 1540 1334
rect 1534 1329 1535 1333
rect 1539 1329 1540 1333
rect 1534 1328 1540 1329
rect 1606 1333 1612 1334
rect 1606 1329 1607 1333
rect 1611 1329 1612 1333
rect 1606 1328 1612 1329
rect 1686 1333 1692 1334
rect 1686 1329 1687 1333
rect 1691 1329 1692 1333
rect 1686 1328 1692 1329
rect 1766 1333 1772 1334
rect 1766 1329 1767 1333
rect 1771 1329 1772 1333
rect 1766 1328 1772 1329
rect 1846 1333 1852 1334
rect 1846 1329 1847 1333
rect 1851 1329 1852 1333
rect 1846 1328 1852 1329
rect 1934 1333 1940 1334
rect 1934 1329 1935 1333
rect 1939 1329 1940 1333
rect 1934 1328 1940 1329
rect 2022 1333 2028 1334
rect 2022 1329 2023 1333
rect 2027 1329 2028 1333
rect 2022 1328 2028 1329
rect 2110 1333 2116 1334
rect 2110 1329 2111 1333
rect 2115 1329 2116 1333
rect 2110 1328 2116 1329
rect 2198 1333 2204 1334
rect 2198 1329 2199 1333
rect 2203 1329 2204 1333
rect 2198 1328 2204 1329
rect 2286 1333 2292 1334
rect 2286 1329 2287 1333
rect 2291 1329 2292 1333
rect 2286 1328 2292 1329
rect 2358 1333 2364 1334
rect 2358 1329 2359 1333
rect 2363 1329 2364 1333
rect 2358 1328 2364 1329
rect 1302 1303 1308 1304
rect 182 1299 188 1300
rect 182 1295 183 1299
rect 187 1295 188 1299
rect 182 1294 188 1295
rect 230 1299 236 1300
rect 230 1295 231 1299
rect 235 1295 236 1299
rect 230 1294 236 1295
rect 286 1299 292 1300
rect 286 1295 287 1299
rect 291 1295 292 1299
rect 286 1294 292 1295
rect 350 1299 356 1300
rect 350 1295 351 1299
rect 355 1295 356 1299
rect 350 1294 356 1295
rect 422 1299 428 1300
rect 422 1295 423 1299
rect 427 1295 428 1299
rect 422 1294 428 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 566 1299 572 1300
rect 566 1295 567 1299
rect 571 1295 572 1299
rect 566 1294 572 1295
rect 638 1299 644 1300
rect 638 1295 639 1299
rect 643 1295 644 1299
rect 638 1294 644 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 766 1299 772 1300
rect 766 1295 767 1299
rect 771 1295 772 1299
rect 766 1294 772 1295
rect 822 1299 828 1300
rect 822 1295 823 1299
rect 827 1295 828 1299
rect 822 1294 828 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 934 1299 940 1300
rect 934 1295 935 1299
rect 939 1295 940 1299
rect 934 1294 940 1295
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1295 1004 1299
rect 1302 1299 1303 1303
rect 1307 1299 1308 1303
rect 1302 1298 1308 1299
rect 1342 1303 1348 1304
rect 1342 1299 1343 1303
rect 1347 1299 1348 1303
rect 1342 1298 1348 1299
rect 1382 1303 1388 1304
rect 1382 1299 1383 1303
rect 1387 1299 1388 1303
rect 1382 1298 1388 1299
rect 1422 1303 1428 1304
rect 1422 1299 1423 1303
rect 1427 1299 1428 1303
rect 1422 1298 1428 1299
rect 1462 1303 1468 1304
rect 1462 1299 1463 1303
rect 1467 1299 1468 1303
rect 1462 1298 1468 1299
rect 1502 1303 1508 1304
rect 1502 1299 1503 1303
rect 1507 1299 1508 1303
rect 1502 1298 1508 1299
rect 1542 1303 1548 1304
rect 1542 1299 1543 1303
rect 1547 1299 1548 1303
rect 1542 1298 1548 1299
rect 1582 1303 1588 1304
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1622 1303 1628 1304
rect 1622 1299 1623 1303
rect 1627 1299 1628 1303
rect 1622 1298 1628 1299
rect 1678 1303 1684 1304
rect 1678 1299 1679 1303
rect 1683 1299 1684 1303
rect 1678 1298 1684 1299
rect 1734 1303 1740 1304
rect 1734 1299 1735 1303
rect 1739 1299 1740 1303
rect 1734 1298 1740 1299
rect 1790 1303 1796 1304
rect 1790 1299 1791 1303
rect 1795 1299 1796 1303
rect 1790 1298 1796 1299
rect 1846 1303 1852 1304
rect 1846 1299 1847 1303
rect 1851 1299 1852 1303
rect 1846 1298 1852 1299
rect 1902 1303 1908 1304
rect 1902 1299 1903 1303
rect 1907 1299 1908 1303
rect 1902 1298 1908 1299
rect 1966 1303 1972 1304
rect 1966 1299 1967 1303
rect 1971 1299 1972 1303
rect 1966 1298 1972 1299
rect 2038 1303 2044 1304
rect 2038 1299 2039 1303
rect 2043 1299 2044 1303
rect 2038 1298 2044 1299
rect 2118 1303 2124 1304
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2198 1303 2204 1304
rect 2198 1299 2199 1303
rect 2203 1299 2204 1303
rect 2198 1298 2204 1299
rect 2286 1303 2292 1304
rect 2286 1299 2287 1303
rect 2291 1299 2292 1303
rect 2286 1298 2292 1299
rect 2358 1303 2364 1304
rect 2358 1299 2359 1303
rect 2363 1299 2364 1303
rect 2358 1298 2364 1299
rect 998 1294 1004 1295
rect 1278 1280 1284 1281
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 110 1271 116 1272
rect 1238 1276 1244 1277
rect 1238 1272 1239 1276
rect 1243 1272 1244 1276
rect 1278 1276 1279 1280
rect 1283 1276 1284 1280
rect 1278 1275 1284 1276
rect 2406 1280 2412 1281
rect 2406 1276 2407 1280
rect 2411 1276 2412 1280
rect 2406 1275 2412 1276
rect 1238 1271 1244 1272
rect 1278 1263 1284 1264
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 1238 1259 1244 1260
rect 1238 1255 1239 1259
rect 1243 1255 1244 1259
rect 1278 1259 1279 1263
rect 1283 1259 1284 1263
rect 1278 1258 1284 1259
rect 2406 1263 2412 1264
rect 2406 1259 2407 1263
rect 2411 1259 2412 1263
rect 2406 1258 2412 1259
rect 1238 1254 1244 1255
rect 1302 1256 1308 1257
rect 182 1252 188 1253
rect 182 1248 183 1252
rect 187 1248 188 1252
rect 182 1247 188 1248
rect 230 1252 236 1253
rect 230 1248 231 1252
rect 235 1248 236 1252
rect 230 1247 236 1248
rect 286 1252 292 1253
rect 286 1248 287 1252
rect 291 1248 292 1252
rect 286 1247 292 1248
rect 350 1252 356 1253
rect 350 1248 351 1252
rect 355 1248 356 1252
rect 350 1247 356 1248
rect 422 1252 428 1253
rect 422 1248 423 1252
rect 427 1248 428 1252
rect 422 1247 428 1248
rect 494 1252 500 1253
rect 494 1248 495 1252
rect 499 1248 500 1252
rect 494 1247 500 1248
rect 566 1252 572 1253
rect 566 1248 567 1252
rect 571 1248 572 1252
rect 566 1247 572 1248
rect 638 1252 644 1253
rect 638 1248 639 1252
rect 643 1248 644 1252
rect 638 1247 644 1248
rect 702 1252 708 1253
rect 702 1248 703 1252
rect 707 1248 708 1252
rect 702 1247 708 1248
rect 766 1252 772 1253
rect 766 1248 767 1252
rect 771 1248 772 1252
rect 766 1247 772 1248
rect 822 1252 828 1253
rect 822 1248 823 1252
rect 827 1248 828 1252
rect 822 1247 828 1248
rect 878 1252 884 1253
rect 878 1248 879 1252
rect 883 1248 884 1252
rect 878 1247 884 1248
rect 934 1252 940 1253
rect 934 1248 935 1252
rect 939 1248 940 1252
rect 934 1247 940 1248
rect 998 1252 1004 1253
rect 998 1248 999 1252
rect 1003 1248 1004 1252
rect 1302 1252 1303 1256
rect 1307 1252 1308 1256
rect 1302 1251 1308 1252
rect 1342 1256 1348 1257
rect 1342 1252 1343 1256
rect 1347 1252 1348 1256
rect 1342 1251 1348 1252
rect 1382 1256 1388 1257
rect 1382 1252 1383 1256
rect 1387 1252 1388 1256
rect 1382 1251 1388 1252
rect 1422 1256 1428 1257
rect 1422 1252 1423 1256
rect 1427 1252 1428 1256
rect 1422 1251 1428 1252
rect 1462 1256 1468 1257
rect 1462 1252 1463 1256
rect 1467 1252 1468 1256
rect 1462 1251 1468 1252
rect 1502 1256 1508 1257
rect 1502 1252 1503 1256
rect 1507 1252 1508 1256
rect 1502 1251 1508 1252
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1582 1256 1588 1257
rect 1582 1252 1583 1256
rect 1587 1252 1588 1256
rect 1582 1251 1588 1252
rect 1622 1256 1628 1257
rect 1622 1252 1623 1256
rect 1627 1252 1628 1256
rect 1622 1251 1628 1252
rect 1678 1256 1684 1257
rect 1678 1252 1679 1256
rect 1683 1252 1684 1256
rect 1678 1251 1684 1252
rect 1734 1256 1740 1257
rect 1734 1252 1735 1256
rect 1739 1252 1740 1256
rect 1734 1251 1740 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1846 1256 1852 1257
rect 1846 1252 1847 1256
rect 1851 1252 1852 1256
rect 1846 1251 1852 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2198 1256 2204 1257
rect 2198 1252 2199 1256
rect 2203 1252 2204 1256
rect 2198 1251 2204 1252
rect 2286 1256 2292 1257
rect 2286 1252 2287 1256
rect 2291 1252 2292 1256
rect 2286 1251 2292 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 998 1247 1004 1248
rect 134 1236 140 1237
rect 134 1232 135 1236
rect 139 1232 140 1236
rect 134 1231 140 1232
rect 174 1236 180 1237
rect 174 1232 175 1236
rect 179 1232 180 1236
rect 174 1231 180 1232
rect 230 1236 236 1237
rect 230 1232 231 1236
rect 235 1232 236 1236
rect 230 1231 236 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 398 1236 404 1237
rect 398 1232 399 1236
rect 403 1232 404 1236
rect 398 1231 404 1232
rect 486 1236 492 1237
rect 486 1232 487 1236
rect 491 1232 492 1236
rect 486 1231 492 1232
rect 574 1236 580 1237
rect 574 1232 575 1236
rect 579 1232 580 1236
rect 574 1231 580 1232
rect 662 1236 668 1237
rect 662 1232 663 1236
rect 667 1232 668 1236
rect 662 1231 668 1232
rect 742 1236 748 1237
rect 742 1232 743 1236
rect 747 1232 748 1236
rect 742 1231 748 1232
rect 814 1236 820 1237
rect 814 1232 815 1236
rect 819 1232 820 1236
rect 814 1231 820 1232
rect 878 1236 884 1237
rect 878 1232 879 1236
rect 883 1232 884 1236
rect 878 1231 884 1232
rect 942 1236 948 1237
rect 942 1232 943 1236
rect 947 1232 948 1236
rect 942 1231 948 1232
rect 1006 1236 1012 1237
rect 1006 1232 1007 1236
rect 1011 1232 1012 1236
rect 1006 1231 1012 1232
rect 1070 1236 1076 1237
rect 1070 1232 1071 1236
rect 1075 1232 1076 1236
rect 1070 1231 1076 1232
rect 1302 1236 1308 1237
rect 1302 1232 1303 1236
rect 1307 1232 1308 1236
rect 1302 1231 1308 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1478 1236 1484 1237
rect 1478 1232 1479 1236
rect 1483 1232 1484 1236
rect 1478 1231 1484 1232
rect 1582 1236 1588 1237
rect 1582 1232 1583 1236
rect 1587 1232 1588 1236
rect 1582 1231 1588 1232
rect 1686 1236 1692 1237
rect 1686 1232 1687 1236
rect 1691 1232 1692 1236
rect 1686 1231 1692 1232
rect 1790 1236 1796 1237
rect 1790 1232 1791 1236
rect 1795 1232 1796 1236
rect 1790 1231 1796 1232
rect 1886 1236 1892 1237
rect 1886 1232 1887 1236
rect 1891 1232 1892 1236
rect 1886 1231 1892 1232
rect 1982 1236 1988 1237
rect 1982 1232 1983 1236
rect 1987 1232 1988 1236
rect 1982 1231 1988 1232
rect 2070 1236 2076 1237
rect 2070 1232 2071 1236
rect 2075 1232 2076 1236
rect 2070 1231 2076 1232
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2222 1236 2228 1237
rect 2222 1232 2223 1236
rect 2227 1232 2228 1236
rect 2222 1231 2228 1232
rect 2302 1236 2308 1237
rect 2302 1232 2303 1236
rect 2307 1232 2308 1236
rect 2302 1231 2308 1232
rect 2358 1236 2364 1237
rect 2358 1232 2359 1236
rect 2363 1232 2364 1236
rect 2358 1231 2364 1232
rect 110 1229 116 1230
rect 110 1225 111 1229
rect 115 1225 116 1229
rect 110 1224 116 1225
rect 1238 1229 1244 1230
rect 1238 1225 1239 1229
rect 1243 1225 1244 1229
rect 1238 1224 1244 1225
rect 1278 1229 1284 1230
rect 1278 1225 1279 1229
rect 1283 1225 1284 1229
rect 1278 1224 1284 1225
rect 2406 1229 2412 1230
rect 2406 1225 2407 1229
rect 2411 1225 2412 1229
rect 2406 1224 2412 1225
rect 110 1212 116 1213
rect 110 1208 111 1212
rect 115 1208 116 1212
rect 110 1207 116 1208
rect 1238 1212 1244 1213
rect 1238 1208 1239 1212
rect 1243 1208 1244 1212
rect 1238 1207 1244 1208
rect 1278 1212 1284 1213
rect 1278 1208 1279 1212
rect 1283 1208 1284 1212
rect 1278 1207 1284 1208
rect 2406 1212 2412 1213
rect 2406 1208 2407 1212
rect 2411 1208 2412 1212
rect 2406 1207 2412 1208
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 174 1189 180 1190
rect 174 1185 175 1189
rect 179 1185 180 1189
rect 174 1184 180 1185
rect 230 1189 236 1190
rect 230 1185 231 1189
rect 235 1185 236 1189
rect 230 1184 236 1185
rect 310 1189 316 1190
rect 310 1185 311 1189
rect 315 1185 316 1189
rect 310 1184 316 1185
rect 398 1189 404 1190
rect 398 1185 399 1189
rect 403 1185 404 1189
rect 398 1184 404 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 574 1189 580 1190
rect 574 1185 575 1189
rect 579 1185 580 1189
rect 574 1184 580 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 742 1189 748 1190
rect 742 1185 743 1189
rect 747 1185 748 1189
rect 742 1184 748 1185
rect 814 1189 820 1190
rect 814 1185 815 1189
rect 819 1185 820 1189
rect 814 1184 820 1185
rect 878 1189 884 1190
rect 878 1185 879 1189
rect 883 1185 884 1189
rect 878 1184 884 1185
rect 942 1189 948 1190
rect 942 1185 943 1189
rect 947 1185 948 1189
rect 942 1184 948 1185
rect 1006 1189 1012 1190
rect 1006 1185 1007 1189
rect 1011 1185 1012 1189
rect 1006 1184 1012 1185
rect 1070 1189 1076 1190
rect 1070 1185 1071 1189
rect 1075 1185 1076 1189
rect 1070 1184 1076 1185
rect 1302 1189 1308 1190
rect 1302 1185 1303 1189
rect 1307 1185 1308 1189
rect 1302 1184 1308 1185
rect 1374 1189 1380 1190
rect 1374 1185 1375 1189
rect 1379 1185 1380 1189
rect 1374 1184 1380 1185
rect 1478 1189 1484 1190
rect 1478 1185 1479 1189
rect 1483 1185 1484 1189
rect 1478 1184 1484 1185
rect 1582 1189 1588 1190
rect 1582 1185 1583 1189
rect 1587 1185 1588 1189
rect 1582 1184 1588 1185
rect 1686 1189 1692 1190
rect 1686 1185 1687 1189
rect 1691 1185 1692 1189
rect 1686 1184 1692 1185
rect 1790 1189 1796 1190
rect 1790 1185 1791 1189
rect 1795 1185 1796 1189
rect 1790 1184 1796 1185
rect 1886 1189 1892 1190
rect 1886 1185 1887 1189
rect 1891 1185 1892 1189
rect 1886 1184 1892 1185
rect 1982 1189 1988 1190
rect 1982 1185 1983 1189
rect 1987 1185 1988 1189
rect 1982 1184 1988 1185
rect 2070 1189 2076 1190
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 2150 1189 2156 1190
rect 2150 1185 2151 1189
rect 2155 1185 2156 1189
rect 2150 1184 2156 1185
rect 2222 1189 2228 1190
rect 2222 1185 2223 1189
rect 2227 1185 2228 1189
rect 2222 1184 2228 1185
rect 2302 1189 2308 1190
rect 2302 1185 2303 1189
rect 2307 1185 2308 1189
rect 2302 1184 2308 1185
rect 2358 1189 2364 1190
rect 2358 1185 2359 1189
rect 2363 1185 2364 1189
rect 2358 1184 2364 1185
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1155 140 1159
rect 134 1154 140 1155
rect 174 1159 180 1160
rect 174 1155 175 1159
rect 179 1155 180 1159
rect 174 1154 180 1155
rect 238 1159 244 1160
rect 238 1155 239 1159
rect 243 1155 244 1159
rect 238 1154 244 1155
rect 326 1159 332 1160
rect 326 1155 327 1159
rect 331 1155 332 1159
rect 326 1154 332 1155
rect 430 1159 436 1160
rect 430 1155 431 1159
rect 435 1155 436 1159
rect 430 1154 436 1155
rect 534 1159 540 1160
rect 534 1155 535 1159
rect 539 1155 540 1159
rect 534 1154 540 1155
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1155 644 1159
rect 638 1154 644 1155
rect 742 1159 748 1160
rect 742 1155 743 1159
rect 747 1155 748 1159
rect 742 1154 748 1155
rect 838 1159 844 1160
rect 838 1155 839 1159
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 918 1159 924 1160
rect 918 1155 919 1159
rect 923 1155 924 1159
rect 918 1154 924 1155
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1070 1159 1076 1160
rect 1070 1155 1071 1159
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 1142 1159 1148 1160
rect 1142 1155 1143 1159
rect 1147 1155 1148 1159
rect 1142 1154 1148 1155
rect 1190 1159 1196 1160
rect 1190 1155 1191 1159
rect 1195 1155 1196 1159
rect 1190 1154 1196 1155
rect 1302 1159 1308 1160
rect 1302 1155 1303 1159
rect 1307 1155 1308 1159
rect 1302 1154 1308 1155
rect 1342 1159 1348 1160
rect 1342 1155 1343 1159
rect 1347 1155 1348 1159
rect 1342 1154 1348 1155
rect 1406 1159 1412 1160
rect 1406 1155 1407 1159
rect 1411 1155 1412 1159
rect 1406 1154 1412 1155
rect 1486 1159 1492 1160
rect 1486 1155 1487 1159
rect 1491 1155 1492 1159
rect 1486 1154 1492 1155
rect 1582 1159 1588 1160
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1686 1159 1692 1160
rect 1686 1155 1687 1159
rect 1691 1155 1692 1159
rect 1686 1154 1692 1155
rect 1798 1159 1804 1160
rect 1798 1155 1799 1159
rect 1803 1155 1804 1159
rect 1798 1154 1804 1155
rect 1902 1159 1908 1160
rect 1902 1155 1903 1159
rect 1907 1155 1908 1159
rect 1902 1154 1908 1155
rect 1998 1159 2004 1160
rect 1998 1155 1999 1159
rect 2003 1155 2004 1159
rect 1998 1154 2004 1155
rect 2078 1159 2084 1160
rect 2078 1155 2079 1159
rect 2083 1155 2084 1159
rect 2078 1154 2084 1155
rect 2158 1159 2164 1160
rect 2158 1155 2159 1159
rect 2163 1155 2164 1159
rect 2158 1154 2164 1155
rect 2230 1159 2236 1160
rect 2230 1155 2231 1159
rect 2235 1155 2236 1159
rect 2230 1154 2236 1155
rect 2302 1159 2308 1160
rect 2302 1155 2303 1159
rect 2307 1155 2308 1159
rect 2302 1154 2308 1155
rect 2358 1159 2364 1160
rect 2358 1155 2359 1159
rect 2363 1155 2364 1159
rect 2358 1154 2364 1155
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 110 1131 116 1132
rect 1238 1136 1244 1137
rect 1238 1132 1239 1136
rect 1243 1132 1244 1136
rect 1238 1131 1244 1132
rect 1278 1136 1284 1137
rect 1278 1132 1279 1136
rect 1283 1132 1284 1136
rect 1278 1131 1284 1132
rect 2406 1136 2412 1137
rect 2406 1132 2407 1136
rect 2411 1132 2412 1136
rect 2406 1131 2412 1132
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 110 1114 116 1115
rect 1238 1119 1244 1120
rect 1238 1115 1239 1119
rect 1243 1115 1244 1119
rect 1238 1114 1244 1115
rect 1278 1119 1284 1120
rect 1278 1115 1279 1119
rect 1283 1115 1284 1119
rect 1278 1114 1284 1115
rect 2406 1119 2412 1120
rect 2406 1115 2407 1119
rect 2411 1115 2412 1119
rect 2406 1114 2412 1115
rect 134 1112 140 1113
rect 134 1108 135 1112
rect 139 1108 140 1112
rect 134 1107 140 1108
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 238 1112 244 1113
rect 238 1108 239 1112
rect 243 1108 244 1112
rect 238 1107 244 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 430 1112 436 1113
rect 430 1108 431 1112
rect 435 1108 436 1112
rect 430 1107 436 1108
rect 534 1112 540 1113
rect 534 1108 535 1112
rect 539 1108 540 1112
rect 534 1107 540 1108
rect 638 1112 644 1113
rect 638 1108 639 1112
rect 643 1108 644 1112
rect 638 1107 644 1108
rect 742 1112 748 1113
rect 742 1108 743 1112
rect 747 1108 748 1112
rect 742 1107 748 1108
rect 838 1112 844 1113
rect 838 1108 839 1112
rect 843 1108 844 1112
rect 838 1107 844 1108
rect 918 1112 924 1113
rect 918 1108 919 1112
rect 923 1108 924 1112
rect 918 1107 924 1108
rect 998 1112 1004 1113
rect 998 1108 999 1112
rect 1003 1108 1004 1112
rect 998 1107 1004 1108
rect 1070 1112 1076 1113
rect 1070 1108 1071 1112
rect 1075 1108 1076 1112
rect 1070 1107 1076 1108
rect 1142 1112 1148 1113
rect 1142 1108 1143 1112
rect 1147 1108 1148 1112
rect 1142 1107 1148 1108
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 1302 1112 1308 1113
rect 1302 1108 1303 1112
rect 1307 1108 1308 1112
rect 1302 1107 1308 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1406 1112 1412 1113
rect 1406 1108 1407 1112
rect 1411 1108 1412 1112
rect 1406 1107 1412 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1582 1112 1588 1113
rect 1582 1108 1583 1112
rect 1587 1108 1588 1112
rect 1582 1107 1588 1108
rect 1686 1112 1692 1113
rect 1686 1108 1687 1112
rect 1691 1108 1692 1112
rect 1686 1107 1692 1108
rect 1798 1112 1804 1113
rect 1798 1108 1799 1112
rect 1803 1108 1804 1112
rect 1798 1107 1804 1108
rect 1902 1112 1908 1113
rect 1902 1108 1903 1112
rect 1907 1108 1908 1112
rect 1902 1107 1908 1108
rect 1998 1112 2004 1113
rect 1998 1108 1999 1112
rect 2003 1108 2004 1112
rect 1998 1107 2004 1108
rect 2078 1112 2084 1113
rect 2078 1108 2079 1112
rect 2083 1108 2084 1112
rect 2078 1107 2084 1108
rect 2158 1112 2164 1113
rect 2158 1108 2159 1112
rect 2163 1108 2164 1112
rect 2158 1107 2164 1108
rect 2230 1112 2236 1113
rect 2230 1108 2231 1112
rect 2235 1108 2236 1112
rect 2230 1107 2236 1108
rect 2302 1112 2308 1113
rect 2302 1108 2303 1112
rect 2307 1108 2308 1112
rect 2302 1107 2308 1108
rect 2358 1112 2364 1113
rect 2358 1108 2359 1112
rect 2363 1108 2364 1112
rect 2358 1107 2364 1108
rect 1430 1100 1436 1101
rect 134 1096 140 1097
rect 134 1092 135 1096
rect 139 1092 140 1096
rect 134 1091 140 1092
rect 174 1096 180 1097
rect 174 1092 175 1096
rect 179 1092 180 1096
rect 174 1091 180 1092
rect 246 1096 252 1097
rect 246 1092 247 1096
rect 251 1092 252 1096
rect 246 1091 252 1092
rect 326 1096 332 1097
rect 326 1092 327 1096
rect 331 1092 332 1096
rect 326 1091 332 1092
rect 414 1096 420 1097
rect 414 1092 415 1096
rect 419 1092 420 1096
rect 414 1091 420 1092
rect 502 1096 508 1097
rect 502 1092 503 1096
rect 507 1092 508 1096
rect 502 1091 508 1092
rect 582 1096 588 1097
rect 582 1092 583 1096
rect 587 1092 588 1096
rect 582 1091 588 1092
rect 662 1096 668 1097
rect 662 1092 663 1096
rect 667 1092 668 1096
rect 662 1091 668 1092
rect 734 1096 740 1097
rect 734 1092 735 1096
rect 739 1092 740 1096
rect 734 1091 740 1092
rect 798 1096 804 1097
rect 798 1092 799 1096
rect 803 1092 804 1096
rect 798 1091 804 1092
rect 862 1096 868 1097
rect 862 1092 863 1096
rect 867 1092 868 1096
rect 862 1091 868 1092
rect 918 1096 924 1097
rect 918 1092 919 1096
rect 923 1092 924 1096
rect 918 1091 924 1092
rect 982 1096 988 1097
rect 982 1092 983 1096
rect 987 1092 988 1096
rect 982 1091 988 1092
rect 1046 1096 1052 1097
rect 1046 1092 1047 1096
rect 1051 1092 1052 1096
rect 1430 1096 1431 1100
rect 1435 1096 1436 1100
rect 1430 1095 1436 1096
rect 1470 1100 1476 1101
rect 1470 1096 1471 1100
rect 1475 1096 1476 1100
rect 1470 1095 1476 1096
rect 1510 1100 1516 1101
rect 1510 1096 1511 1100
rect 1515 1096 1516 1100
rect 1510 1095 1516 1096
rect 1558 1100 1564 1101
rect 1558 1096 1559 1100
rect 1563 1096 1564 1100
rect 1558 1095 1564 1096
rect 1614 1100 1620 1101
rect 1614 1096 1615 1100
rect 1619 1096 1620 1100
rect 1614 1095 1620 1096
rect 1670 1100 1676 1101
rect 1670 1096 1671 1100
rect 1675 1096 1676 1100
rect 1670 1095 1676 1096
rect 1726 1100 1732 1101
rect 1726 1096 1727 1100
rect 1731 1096 1732 1100
rect 1726 1095 1732 1096
rect 1774 1100 1780 1101
rect 1774 1096 1775 1100
rect 1779 1096 1780 1100
rect 1774 1095 1780 1096
rect 1822 1100 1828 1101
rect 1822 1096 1823 1100
rect 1827 1096 1828 1100
rect 1822 1095 1828 1096
rect 1870 1100 1876 1101
rect 1870 1096 1871 1100
rect 1875 1096 1876 1100
rect 1870 1095 1876 1096
rect 1918 1100 1924 1101
rect 1918 1096 1919 1100
rect 1923 1096 1924 1100
rect 1918 1095 1924 1096
rect 1966 1100 1972 1101
rect 1966 1096 1967 1100
rect 1971 1096 1972 1100
rect 1966 1095 1972 1096
rect 2014 1100 2020 1101
rect 2014 1096 2015 1100
rect 2019 1096 2020 1100
rect 2014 1095 2020 1096
rect 2062 1100 2068 1101
rect 2062 1096 2063 1100
rect 2067 1096 2068 1100
rect 2062 1095 2068 1096
rect 2118 1100 2124 1101
rect 2118 1096 2119 1100
rect 2123 1096 2124 1100
rect 2118 1095 2124 1096
rect 2174 1100 2180 1101
rect 2174 1096 2175 1100
rect 2179 1096 2180 1100
rect 2174 1095 2180 1096
rect 2230 1100 2236 1101
rect 2230 1096 2231 1100
rect 2235 1096 2236 1100
rect 2230 1095 2236 1096
rect 1046 1091 1052 1092
rect 1278 1093 1284 1094
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 110 1084 116 1085
rect 1238 1089 1244 1090
rect 1238 1085 1239 1089
rect 1243 1085 1244 1089
rect 1278 1089 1279 1093
rect 1283 1089 1284 1093
rect 1278 1088 1284 1089
rect 2406 1093 2412 1094
rect 2406 1089 2407 1093
rect 2411 1089 2412 1093
rect 2406 1088 2412 1089
rect 1238 1084 1244 1085
rect 1278 1076 1284 1077
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 110 1067 116 1068
rect 1238 1072 1244 1073
rect 1238 1068 1239 1072
rect 1243 1068 1244 1072
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 2406 1076 2412 1077
rect 2406 1072 2407 1076
rect 2411 1072 2412 1076
rect 2406 1071 2412 1072
rect 1238 1067 1244 1068
rect 1430 1053 1436 1054
rect 134 1049 140 1050
rect 134 1045 135 1049
rect 139 1045 140 1049
rect 134 1044 140 1045
rect 174 1049 180 1050
rect 174 1045 175 1049
rect 179 1045 180 1049
rect 174 1044 180 1045
rect 246 1049 252 1050
rect 246 1045 247 1049
rect 251 1045 252 1049
rect 246 1044 252 1045
rect 326 1049 332 1050
rect 326 1045 327 1049
rect 331 1045 332 1049
rect 326 1044 332 1045
rect 414 1049 420 1050
rect 414 1045 415 1049
rect 419 1045 420 1049
rect 414 1044 420 1045
rect 502 1049 508 1050
rect 502 1045 503 1049
rect 507 1045 508 1049
rect 502 1044 508 1045
rect 582 1049 588 1050
rect 582 1045 583 1049
rect 587 1045 588 1049
rect 582 1044 588 1045
rect 662 1049 668 1050
rect 662 1045 663 1049
rect 667 1045 668 1049
rect 662 1044 668 1045
rect 734 1049 740 1050
rect 734 1045 735 1049
rect 739 1045 740 1049
rect 734 1044 740 1045
rect 798 1049 804 1050
rect 798 1045 799 1049
rect 803 1045 804 1049
rect 798 1044 804 1045
rect 862 1049 868 1050
rect 862 1045 863 1049
rect 867 1045 868 1049
rect 862 1044 868 1045
rect 918 1049 924 1050
rect 918 1045 919 1049
rect 923 1045 924 1049
rect 918 1044 924 1045
rect 982 1049 988 1050
rect 982 1045 983 1049
rect 987 1045 988 1049
rect 982 1044 988 1045
rect 1046 1049 1052 1050
rect 1046 1045 1047 1049
rect 1051 1045 1052 1049
rect 1430 1049 1431 1053
rect 1435 1049 1436 1053
rect 1430 1048 1436 1049
rect 1470 1053 1476 1054
rect 1470 1049 1471 1053
rect 1475 1049 1476 1053
rect 1470 1048 1476 1049
rect 1510 1053 1516 1054
rect 1510 1049 1511 1053
rect 1515 1049 1516 1053
rect 1510 1048 1516 1049
rect 1558 1053 1564 1054
rect 1558 1049 1559 1053
rect 1563 1049 1564 1053
rect 1558 1048 1564 1049
rect 1614 1053 1620 1054
rect 1614 1049 1615 1053
rect 1619 1049 1620 1053
rect 1614 1048 1620 1049
rect 1670 1053 1676 1054
rect 1670 1049 1671 1053
rect 1675 1049 1676 1053
rect 1670 1048 1676 1049
rect 1726 1053 1732 1054
rect 1726 1049 1727 1053
rect 1731 1049 1732 1053
rect 1726 1048 1732 1049
rect 1774 1053 1780 1054
rect 1774 1049 1775 1053
rect 1779 1049 1780 1053
rect 1774 1048 1780 1049
rect 1822 1053 1828 1054
rect 1822 1049 1823 1053
rect 1827 1049 1828 1053
rect 1822 1048 1828 1049
rect 1870 1053 1876 1054
rect 1870 1049 1871 1053
rect 1875 1049 1876 1053
rect 1870 1048 1876 1049
rect 1918 1053 1924 1054
rect 1918 1049 1919 1053
rect 1923 1049 1924 1053
rect 1918 1048 1924 1049
rect 1966 1053 1972 1054
rect 1966 1049 1967 1053
rect 1971 1049 1972 1053
rect 1966 1048 1972 1049
rect 2014 1053 2020 1054
rect 2014 1049 2015 1053
rect 2019 1049 2020 1053
rect 2014 1048 2020 1049
rect 2062 1053 2068 1054
rect 2062 1049 2063 1053
rect 2067 1049 2068 1053
rect 2062 1048 2068 1049
rect 2118 1053 2124 1054
rect 2118 1049 2119 1053
rect 2123 1049 2124 1053
rect 2118 1048 2124 1049
rect 2174 1053 2180 1054
rect 2174 1049 2175 1053
rect 2179 1049 2180 1053
rect 2174 1048 2180 1049
rect 2230 1053 2236 1054
rect 2230 1049 2231 1053
rect 2235 1049 2236 1053
rect 2230 1048 2236 1049
rect 1046 1044 1052 1045
rect 1574 1023 1580 1024
rect 174 1019 180 1020
rect 174 1015 175 1019
rect 179 1015 180 1019
rect 174 1014 180 1015
rect 254 1019 260 1020
rect 254 1015 255 1019
rect 259 1015 260 1019
rect 254 1014 260 1015
rect 326 1019 332 1020
rect 326 1015 327 1019
rect 331 1015 332 1019
rect 326 1014 332 1015
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 462 1019 468 1020
rect 462 1015 463 1019
rect 467 1015 468 1019
rect 462 1014 468 1015
rect 518 1019 524 1020
rect 518 1015 519 1019
rect 523 1015 524 1019
rect 518 1014 524 1015
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 574 1014 580 1015
rect 622 1019 628 1020
rect 622 1015 623 1019
rect 627 1015 628 1019
rect 622 1014 628 1015
rect 670 1019 676 1020
rect 670 1015 671 1019
rect 675 1015 676 1019
rect 670 1014 676 1015
rect 734 1019 740 1020
rect 734 1015 735 1019
rect 739 1015 740 1019
rect 734 1014 740 1015
rect 806 1019 812 1020
rect 806 1015 807 1019
rect 811 1015 812 1019
rect 806 1014 812 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 998 1019 1004 1020
rect 998 1015 999 1019
rect 1003 1015 1004 1019
rect 998 1014 1004 1015
rect 1102 1019 1108 1020
rect 1102 1015 1103 1019
rect 1107 1015 1108 1019
rect 1102 1014 1108 1015
rect 1190 1019 1196 1020
rect 1190 1015 1191 1019
rect 1195 1015 1196 1019
rect 1574 1019 1575 1023
rect 1579 1019 1580 1023
rect 1574 1018 1580 1019
rect 1614 1023 1620 1024
rect 1614 1019 1615 1023
rect 1619 1019 1620 1023
rect 1614 1018 1620 1019
rect 1654 1023 1660 1024
rect 1654 1019 1655 1023
rect 1659 1019 1660 1023
rect 1654 1018 1660 1019
rect 1694 1023 1700 1024
rect 1694 1019 1695 1023
rect 1699 1019 1700 1023
rect 1694 1018 1700 1019
rect 1734 1023 1740 1024
rect 1734 1019 1735 1023
rect 1739 1019 1740 1023
rect 1734 1018 1740 1019
rect 1774 1023 1780 1024
rect 1774 1019 1775 1023
rect 1779 1019 1780 1023
rect 1774 1018 1780 1019
rect 1822 1023 1828 1024
rect 1822 1019 1823 1023
rect 1827 1019 1828 1023
rect 1822 1018 1828 1019
rect 1878 1023 1884 1024
rect 1878 1019 1879 1023
rect 1883 1019 1884 1023
rect 1878 1018 1884 1019
rect 1942 1023 1948 1024
rect 1942 1019 1943 1023
rect 1947 1019 1948 1023
rect 1942 1018 1948 1019
rect 2014 1023 2020 1024
rect 2014 1019 2015 1023
rect 2019 1019 2020 1023
rect 2014 1018 2020 1019
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2174 1023 2180 1024
rect 2174 1019 2175 1023
rect 2179 1019 2180 1023
rect 2174 1018 2180 1019
rect 2254 1023 2260 1024
rect 2254 1019 2255 1023
rect 2259 1019 2260 1023
rect 2254 1018 2260 1019
rect 1190 1014 1196 1015
rect 1278 1000 1284 1001
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1238 996 1244 997
rect 1238 992 1239 996
rect 1243 992 1244 996
rect 1278 996 1279 1000
rect 1283 996 1284 1000
rect 1278 995 1284 996
rect 2406 1000 2412 1001
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 2406 995 2412 996
rect 1238 991 1244 992
rect 1278 983 1284 984
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 1238 979 1244 980
rect 1238 975 1239 979
rect 1243 975 1244 979
rect 1278 979 1279 983
rect 1283 979 1284 983
rect 1278 978 1284 979
rect 2406 983 2412 984
rect 2406 979 2407 983
rect 2411 979 2412 983
rect 2406 978 2412 979
rect 1238 974 1244 975
rect 1574 976 1580 977
rect 174 972 180 973
rect 174 968 175 972
rect 179 968 180 972
rect 174 967 180 968
rect 254 972 260 973
rect 254 968 255 972
rect 259 968 260 972
rect 254 967 260 968
rect 326 972 332 973
rect 326 968 327 972
rect 331 968 332 972
rect 326 967 332 968
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 462 972 468 973
rect 462 968 463 972
rect 467 968 468 972
rect 462 967 468 968
rect 518 972 524 973
rect 518 968 519 972
rect 523 968 524 972
rect 518 967 524 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 622 972 628 973
rect 622 968 623 972
rect 627 968 628 972
rect 622 967 628 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 806 972 812 973
rect 806 968 807 972
rect 811 968 812 972
rect 806 967 812 968
rect 894 972 900 973
rect 894 968 895 972
rect 899 968 900 972
rect 894 967 900 968
rect 998 972 1004 973
rect 998 968 999 972
rect 1003 968 1004 972
rect 998 967 1004 968
rect 1102 972 1108 973
rect 1102 968 1103 972
rect 1107 968 1108 972
rect 1102 967 1108 968
rect 1190 972 1196 973
rect 1190 968 1191 972
rect 1195 968 1196 972
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1614 976 1620 977
rect 1614 972 1615 976
rect 1619 972 1620 976
rect 1614 971 1620 972
rect 1654 976 1660 977
rect 1654 972 1655 976
rect 1659 972 1660 976
rect 1654 971 1660 972
rect 1694 976 1700 977
rect 1694 972 1695 976
rect 1699 972 1700 976
rect 1694 971 1700 972
rect 1734 976 1740 977
rect 1734 972 1735 976
rect 1739 972 1740 976
rect 1734 971 1740 972
rect 1774 976 1780 977
rect 1774 972 1775 976
rect 1779 972 1780 976
rect 1774 971 1780 972
rect 1822 976 1828 977
rect 1822 972 1823 976
rect 1827 972 1828 976
rect 1822 971 1828 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1942 976 1948 977
rect 1942 972 1943 976
rect 1947 972 1948 976
rect 1942 971 1948 972
rect 2014 976 2020 977
rect 2014 972 2015 976
rect 2019 972 2020 976
rect 2014 971 2020 972
rect 2094 976 2100 977
rect 2094 972 2095 976
rect 2099 972 2100 976
rect 2094 971 2100 972
rect 2174 976 2180 977
rect 2174 972 2175 976
rect 2179 972 2180 976
rect 2174 971 2180 972
rect 2254 976 2260 977
rect 2254 972 2255 976
rect 2259 972 2260 976
rect 2254 971 2260 972
rect 1190 967 1196 968
rect 214 960 220 961
rect 214 956 215 960
rect 219 956 220 960
rect 214 955 220 956
rect 254 960 260 961
rect 254 956 255 960
rect 259 956 260 960
rect 254 955 260 956
rect 302 960 308 961
rect 302 956 303 960
rect 307 956 308 960
rect 302 955 308 956
rect 358 960 364 961
rect 358 956 359 960
rect 363 956 364 960
rect 358 955 364 956
rect 414 960 420 961
rect 414 956 415 960
rect 419 956 420 960
rect 414 955 420 956
rect 462 960 468 961
rect 462 956 463 960
rect 467 956 468 960
rect 462 955 468 956
rect 518 960 524 961
rect 518 956 519 960
rect 523 956 524 960
rect 518 955 524 956
rect 574 960 580 961
rect 574 956 575 960
rect 579 956 580 960
rect 574 955 580 956
rect 638 960 644 961
rect 638 956 639 960
rect 643 956 644 960
rect 638 955 644 956
rect 710 960 716 961
rect 710 956 711 960
rect 715 956 716 960
rect 710 955 716 956
rect 782 960 788 961
rect 782 956 783 960
rect 787 956 788 960
rect 782 955 788 956
rect 854 960 860 961
rect 854 956 855 960
rect 859 956 860 960
rect 854 955 860 956
rect 926 960 932 961
rect 926 956 927 960
rect 931 956 932 960
rect 926 955 932 956
rect 998 960 1004 961
rect 998 956 999 960
rect 1003 956 1004 960
rect 998 955 1004 956
rect 1070 960 1076 961
rect 1070 956 1071 960
rect 1075 956 1076 960
rect 1070 955 1076 956
rect 1142 960 1148 961
rect 1142 956 1143 960
rect 1147 956 1148 960
rect 1142 955 1148 956
rect 1190 960 1196 961
rect 1190 956 1191 960
rect 1195 956 1196 960
rect 1190 955 1196 956
rect 1302 956 1308 957
rect 110 953 116 954
rect 110 949 111 953
rect 115 949 116 953
rect 110 948 116 949
rect 1238 953 1244 954
rect 1238 949 1239 953
rect 1243 949 1244 953
rect 1302 952 1303 956
rect 1307 952 1308 956
rect 1302 951 1308 952
rect 1350 956 1356 957
rect 1350 952 1351 956
rect 1355 952 1356 956
rect 1350 951 1356 952
rect 1430 956 1436 957
rect 1430 952 1431 956
rect 1435 952 1436 956
rect 1430 951 1436 952
rect 1510 956 1516 957
rect 1510 952 1511 956
rect 1515 952 1516 956
rect 1510 951 1516 952
rect 1590 956 1596 957
rect 1590 952 1591 956
rect 1595 952 1596 956
rect 1590 951 1596 952
rect 1678 956 1684 957
rect 1678 952 1679 956
rect 1683 952 1684 956
rect 1678 951 1684 952
rect 1766 956 1772 957
rect 1766 952 1767 956
rect 1771 952 1772 956
rect 1766 951 1772 952
rect 1854 956 1860 957
rect 1854 952 1855 956
rect 1859 952 1860 956
rect 1854 951 1860 952
rect 1942 956 1948 957
rect 1942 952 1943 956
rect 1947 952 1948 956
rect 1942 951 1948 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2102 956 2108 957
rect 2102 952 2103 956
rect 2107 952 2108 956
rect 2102 951 2108 952
rect 2182 956 2188 957
rect 2182 952 2183 956
rect 2187 952 2188 956
rect 2182 951 2188 952
rect 2270 956 2276 957
rect 2270 952 2271 956
rect 2275 952 2276 956
rect 2270 951 2276 952
rect 1238 948 1244 949
rect 1278 949 1284 950
rect 1278 945 1279 949
rect 1283 945 1284 949
rect 1278 944 1284 945
rect 2406 949 2412 950
rect 2406 945 2407 949
rect 2411 945 2412 949
rect 2406 944 2412 945
rect 110 936 116 937
rect 110 932 111 936
rect 115 932 116 936
rect 110 931 116 932
rect 1238 936 1244 937
rect 1238 932 1239 936
rect 1243 932 1244 936
rect 1238 931 1244 932
rect 1278 932 1284 933
rect 1278 928 1279 932
rect 1283 928 1284 932
rect 1278 927 1284 928
rect 2406 932 2412 933
rect 2406 928 2407 932
rect 2411 928 2412 932
rect 2406 927 2412 928
rect 214 913 220 914
rect 214 909 215 913
rect 219 909 220 913
rect 214 908 220 909
rect 254 913 260 914
rect 254 909 255 913
rect 259 909 260 913
rect 254 908 260 909
rect 302 913 308 914
rect 302 909 303 913
rect 307 909 308 913
rect 302 908 308 909
rect 358 913 364 914
rect 358 909 359 913
rect 363 909 364 913
rect 358 908 364 909
rect 414 913 420 914
rect 414 909 415 913
rect 419 909 420 913
rect 414 908 420 909
rect 462 913 468 914
rect 462 909 463 913
rect 467 909 468 913
rect 462 908 468 909
rect 518 913 524 914
rect 518 909 519 913
rect 523 909 524 913
rect 518 908 524 909
rect 574 913 580 914
rect 574 909 575 913
rect 579 909 580 913
rect 574 908 580 909
rect 638 913 644 914
rect 638 909 639 913
rect 643 909 644 913
rect 638 908 644 909
rect 710 913 716 914
rect 710 909 711 913
rect 715 909 716 913
rect 710 908 716 909
rect 782 913 788 914
rect 782 909 783 913
rect 787 909 788 913
rect 782 908 788 909
rect 854 913 860 914
rect 854 909 855 913
rect 859 909 860 913
rect 854 908 860 909
rect 926 913 932 914
rect 926 909 927 913
rect 931 909 932 913
rect 926 908 932 909
rect 998 913 1004 914
rect 998 909 999 913
rect 1003 909 1004 913
rect 998 908 1004 909
rect 1070 913 1076 914
rect 1070 909 1071 913
rect 1075 909 1076 913
rect 1070 908 1076 909
rect 1142 913 1148 914
rect 1142 909 1143 913
rect 1147 909 1148 913
rect 1142 908 1148 909
rect 1190 913 1196 914
rect 1190 909 1191 913
rect 1195 909 1196 913
rect 1190 908 1196 909
rect 1302 909 1308 910
rect 1302 905 1303 909
rect 1307 905 1308 909
rect 1302 904 1308 905
rect 1350 909 1356 910
rect 1350 905 1351 909
rect 1355 905 1356 909
rect 1350 904 1356 905
rect 1430 909 1436 910
rect 1430 905 1431 909
rect 1435 905 1436 909
rect 1430 904 1436 905
rect 1510 909 1516 910
rect 1510 905 1511 909
rect 1515 905 1516 909
rect 1510 904 1516 905
rect 1590 909 1596 910
rect 1590 905 1591 909
rect 1595 905 1596 909
rect 1590 904 1596 905
rect 1678 909 1684 910
rect 1678 905 1679 909
rect 1683 905 1684 909
rect 1678 904 1684 905
rect 1766 909 1772 910
rect 1766 905 1767 909
rect 1771 905 1772 909
rect 1766 904 1772 905
rect 1854 909 1860 910
rect 1854 905 1855 909
rect 1859 905 1860 909
rect 1854 904 1860 905
rect 1942 909 1948 910
rect 1942 905 1943 909
rect 1947 905 1948 909
rect 1942 904 1948 905
rect 2022 909 2028 910
rect 2022 905 2023 909
rect 2027 905 2028 909
rect 2022 904 2028 905
rect 2102 909 2108 910
rect 2102 905 2103 909
rect 2107 905 2108 909
rect 2102 904 2108 905
rect 2182 909 2188 910
rect 2182 905 2183 909
rect 2187 905 2188 909
rect 2182 904 2188 905
rect 2270 909 2276 910
rect 2270 905 2271 909
rect 2275 905 2276 909
rect 2270 904 2276 905
rect 1438 879 1444 880
rect 190 875 196 876
rect 190 871 191 875
rect 195 871 196 875
rect 190 870 196 871
rect 230 875 236 876
rect 230 871 231 875
rect 235 871 236 875
rect 230 870 236 871
rect 286 875 292 876
rect 286 871 287 875
rect 291 871 292 875
rect 286 870 292 871
rect 358 875 364 876
rect 358 871 359 875
rect 363 871 364 875
rect 358 870 364 871
rect 446 875 452 876
rect 446 871 447 875
rect 451 871 452 875
rect 446 870 452 871
rect 542 875 548 876
rect 542 871 543 875
rect 547 871 548 875
rect 542 870 548 871
rect 638 875 644 876
rect 638 871 639 875
rect 643 871 644 875
rect 638 870 644 871
rect 726 875 732 876
rect 726 871 727 875
rect 731 871 732 875
rect 726 870 732 871
rect 806 875 812 876
rect 806 871 807 875
rect 811 871 812 875
rect 806 870 812 871
rect 886 875 892 876
rect 886 871 887 875
rect 891 871 892 875
rect 886 870 892 871
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 958 870 964 871
rect 1022 875 1028 876
rect 1022 871 1023 875
rect 1027 871 1028 875
rect 1022 870 1028 871
rect 1086 875 1092 876
rect 1086 871 1087 875
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 1158 875 1164 876
rect 1158 871 1159 875
rect 1163 871 1164 875
rect 1438 875 1439 879
rect 1443 875 1444 879
rect 1438 874 1444 875
rect 1478 879 1484 880
rect 1478 875 1479 879
rect 1483 875 1484 879
rect 1478 874 1484 875
rect 1518 879 1524 880
rect 1518 875 1519 879
rect 1523 875 1524 879
rect 1518 874 1524 875
rect 1558 879 1564 880
rect 1558 875 1559 879
rect 1563 875 1564 879
rect 1558 874 1564 875
rect 1606 879 1612 880
rect 1606 875 1607 879
rect 1611 875 1612 879
rect 1606 874 1612 875
rect 1654 879 1660 880
rect 1654 875 1655 879
rect 1659 875 1660 879
rect 1654 874 1660 875
rect 1710 879 1716 880
rect 1710 875 1711 879
rect 1715 875 1716 879
rect 1710 874 1716 875
rect 1774 879 1780 880
rect 1774 875 1775 879
rect 1779 875 1780 879
rect 1774 874 1780 875
rect 1846 879 1852 880
rect 1846 875 1847 879
rect 1851 875 1852 879
rect 1846 874 1852 875
rect 1918 879 1924 880
rect 1918 875 1919 879
rect 1923 875 1924 879
rect 1918 874 1924 875
rect 1990 879 1996 880
rect 1990 875 1991 879
rect 1995 875 1996 879
rect 1990 874 1996 875
rect 2062 879 2068 880
rect 2062 875 2063 879
rect 2067 875 2068 879
rect 2062 874 2068 875
rect 2134 879 2140 880
rect 2134 875 2135 879
rect 2139 875 2140 879
rect 2134 874 2140 875
rect 2214 879 2220 880
rect 2214 875 2215 879
rect 2219 875 2220 879
rect 2214 874 2220 875
rect 2294 879 2300 880
rect 2294 875 2295 879
rect 2299 875 2300 879
rect 2294 874 2300 875
rect 1158 870 1164 871
rect 1278 856 1284 857
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 110 847 116 848
rect 1238 852 1244 853
rect 1238 848 1239 852
rect 1243 848 1244 852
rect 1278 852 1279 856
rect 1283 852 1284 856
rect 1278 851 1284 852
rect 2406 856 2412 857
rect 2406 852 2407 856
rect 2411 852 2412 856
rect 2406 851 2412 852
rect 1238 847 1244 848
rect 1278 839 1284 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 1238 835 1244 836
rect 1238 831 1239 835
rect 1243 831 1244 835
rect 1278 835 1279 839
rect 1283 835 1284 839
rect 1278 834 1284 835
rect 2406 839 2412 840
rect 2406 835 2407 839
rect 2411 835 2412 839
rect 2406 834 2412 835
rect 1238 830 1244 831
rect 1438 832 1444 833
rect 190 828 196 829
rect 190 824 191 828
rect 195 824 196 828
rect 190 823 196 824
rect 230 828 236 829
rect 230 824 231 828
rect 235 824 236 828
rect 230 823 236 824
rect 286 828 292 829
rect 286 824 287 828
rect 291 824 292 828
rect 286 823 292 824
rect 358 828 364 829
rect 358 824 359 828
rect 363 824 364 828
rect 358 823 364 824
rect 446 828 452 829
rect 446 824 447 828
rect 451 824 452 828
rect 446 823 452 824
rect 542 828 548 829
rect 542 824 543 828
rect 547 824 548 828
rect 542 823 548 824
rect 638 828 644 829
rect 638 824 639 828
rect 643 824 644 828
rect 638 823 644 824
rect 726 828 732 829
rect 726 824 727 828
rect 731 824 732 828
rect 726 823 732 824
rect 806 828 812 829
rect 806 824 807 828
rect 811 824 812 828
rect 806 823 812 824
rect 886 828 892 829
rect 886 824 887 828
rect 891 824 892 828
rect 886 823 892 824
rect 958 828 964 829
rect 958 824 959 828
rect 963 824 964 828
rect 958 823 964 824
rect 1022 828 1028 829
rect 1022 824 1023 828
rect 1027 824 1028 828
rect 1022 823 1028 824
rect 1086 828 1092 829
rect 1086 824 1087 828
rect 1091 824 1092 828
rect 1086 823 1092 824
rect 1158 828 1164 829
rect 1158 824 1159 828
rect 1163 824 1164 828
rect 1438 828 1439 832
rect 1443 828 1444 832
rect 1438 827 1444 828
rect 1478 832 1484 833
rect 1478 828 1479 832
rect 1483 828 1484 832
rect 1478 827 1484 828
rect 1518 832 1524 833
rect 1518 828 1519 832
rect 1523 828 1524 832
rect 1518 827 1524 828
rect 1558 832 1564 833
rect 1558 828 1559 832
rect 1563 828 1564 832
rect 1558 827 1564 828
rect 1606 832 1612 833
rect 1606 828 1607 832
rect 1611 828 1612 832
rect 1606 827 1612 828
rect 1654 832 1660 833
rect 1654 828 1655 832
rect 1659 828 1660 832
rect 1654 827 1660 828
rect 1710 832 1716 833
rect 1710 828 1711 832
rect 1715 828 1716 832
rect 1710 827 1716 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1846 832 1852 833
rect 1846 828 1847 832
rect 1851 828 1852 832
rect 1846 827 1852 828
rect 1918 832 1924 833
rect 1918 828 1919 832
rect 1923 828 1924 832
rect 1918 827 1924 828
rect 1990 832 1996 833
rect 1990 828 1991 832
rect 1995 828 1996 832
rect 1990 827 1996 828
rect 2062 832 2068 833
rect 2062 828 2063 832
rect 2067 828 2068 832
rect 2062 827 2068 828
rect 2134 832 2140 833
rect 2134 828 2135 832
rect 2139 828 2140 832
rect 2134 827 2140 828
rect 2214 832 2220 833
rect 2214 828 2215 832
rect 2219 828 2220 832
rect 2214 827 2220 828
rect 2294 832 2300 833
rect 2294 828 2295 832
rect 2299 828 2300 832
rect 2294 827 2300 828
rect 1158 823 1164 824
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 174 816 180 817
rect 174 812 175 816
rect 179 812 180 816
rect 174 811 180 812
rect 238 816 244 817
rect 238 812 239 816
rect 243 812 244 816
rect 238 811 244 812
rect 326 816 332 817
rect 326 812 327 816
rect 331 812 332 816
rect 326 811 332 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 590 816 596 817
rect 590 812 591 816
rect 595 812 596 816
rect 590 811 596 812
rect 670 816 676 817
rect 670 812 671 816
rect 675 812 676 816
rect 670 811 676 812
rect 742 816 748 817
rect 742 812 743 816
rect 747 812 748 816
rect 742 811 748 812
rect 814 816 820 817
rect 814 812 815 816
rect 819 812 820 816
rect 814 811 820 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 942 816 948 817
rect 942 812 943 816
rect 947 812 948 816
rect 942 811 948 812
rect 1014 816 1020 817
rect 1014 812 1015 816
rect 1019 812 1020 816
rect 1014 811 1020 812
rect 110 809 116 810
rect 110 805 111 809
rect 115 805 116 809
rect 110 804 116 805
rect 1238 809 1244 810
rect 1238 805 1239 809
rect 1243 805 1244 809
rect 1238 804 1244 805
rect 1358 808 1364 809
rect 1358 804 1359 808
rect 1363 804 1364 808
rect 1358 803 1364 804
rect 1414 808 1420 809
rect 1414 804 1415 808
rect 1419 804 1420 808
rect 1414 803 1420 804
rect 1470 808 1476 809
rect 1470 804 1471 808
rect 1475 804 1476 808
rect 1470 803 1476 804
rect 1534 808 1540 809
rect 1534 804 1535 808
rect 1539 804 1540 808
rect 1534 803 1540 804
rect 1590 808 1596 809
rect 1590 804 1591 808
rect 1595 804 1596 808
rect 1590 803 1596 804
rect 1646 808 1652 809
rect 1646 804 1647 808
rect 1651 804 1652 808
rect 1646 803 1652 804
rect 1702 808 1708 809
rect 1702 804 1703 808
rect 1707 804 1708 808
rect 1702 803 1708 804
rect 1758 808 1764 809
rect 1758 804 1759 808
rect 1763 804 1764 808
rect 1758 803 1764 804
rect 1814 808 1820 809
rect 1814 804 1815 808
rect 1819 804 1820 808
rect 1814 803 1820 804
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 1934 808 1940 809
rect 1934 804 1935 808
rect 1939 804 1940 808
rect 1934 803 1940 804
rect 1998 808 2004 809
rect 1998 804 1999 808
rect 2003 804 2004 808
rect 1998 803 2004 804
rect 2070 808 2076 809
rect 2070 804 2071 808
rect 2075 804 2076 808
rect 2070 803 2076 804
rect 2142 808 2148 809
rect 2142 804 2143 808
rect 2147 804 2148 808
rect 2142 803 2148 804
rect 2222 808 2228 809
rect 2222 804 2223 808
rect 2227 804 2228 808
rect 2222 803 2228 804
rect 2302 808 2308 809
rect 2302 804 2303 808
rect 2307 804 2308 808
rect 2302 803 2308 804
rect 2358 808 2364 809
rect 2358 804 2359 808
rect 2363 804 2364 808
rect 2358 803 2364 804
rect 1278 801 1284 802
rect 1278 797 1279 801
rect 1283 797 1284 801
rect 1278 796 1284 797
rect 2406 801 2412 802
rect 2406 797 2407 801
rect 2411 797 2412 801
rect 2406 796 2412 797
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 110 787 116 788
rect 1238 792 1244 793
rect 1238 788 1239 792
rect 1243 788 1244 792
rect 1238 787 1244 788
rect 1278 784 1284 785
rect 1278 780 1279 784
rect 1283 780 1284 784
rect 1278 779 1284 780
rect 2406 784 2412 785
rect 2406 780 2407 784
rect 2411 780 2412 784
rect 2406 779 2412 780
rect 134 769 140 770
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 174 769 180 770
rect 174 765 175 769
rect 179 765 180 769
rect 174 764 180 765
rect 238 769 244 770
rect 238 765 239 769
rect 243 765 244 769
rect 238 764 244 765
rect 326 769 332 770
rect 326 765 327 769
rect 331 765 332 769
rect 326 764 332 765
rect 414 769 420 770
rect 414 765 415 769
rect 419 765 420 769
rect 414 764 420 765
rect 502 769 508 770
rect 502 765 503 769
rect 507 765 508 769
rect 502 764 508 765
rect 590 769 596 770
rect 590 765 591 769
rect 595 765 596 769
rect 590 764 596 765
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 742 769 748 770
rect 742 765 743 769
rect 747 765 748 769
rect 742 764 748 765
rect 814 769 820 770
rect 814 765 815 769
rect 819 765 820 769
rect 814 764 820 765
rect 878 769 884 770
rect 878 765 879 769
rect 883 765 884 769
rect 878 764 884 765
rect 942 769 948 770
rect 942 765 943 769
rect 947 765 948 769
rect 942 764 948 765
rect 1014 769 1020 770
rect 1014 765 1015 769
rect 1019 765 1020 769
rect 1014 764 1020 765
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1534 761 1540 762
rect 1534 757 1535 761
rect 1539 757 1540 761
rect 1534 756 1540 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1590 756 1596 757
rect 1646 761 1652 762
rect 1646 757 1647 761
rect 1651 757 1652 761
rect 1646 756 1652 757
rect 1702 761 1708 762
rect 1702 757 1703 761
rect 1707 757 1708 761
rect 1702 756 1708 757
rect 1758 761 1764 762
rect 1758 757 1759 761
rect 1763 757 1764 761
rect 1758 756 1764 757
rect 1814 761 1820 762
rect 1814 757 1815 761
rect 1819 757 1820 761
rect 1814 756 1820 757
rect 1870 761 1876 762
rect 1870 757 1871 761
rect 1875 757 1876 761
rect 1870 756 1876 757
rect 1934 761 1940 762
rect 1934 757 1935 761
rect 1939 757 1940 761
rect 1934 756 1940 757
rect 1998 761 2004 762
rect 1998 757 1999 761
rect 2003 757 2004 761
rect 1998 756 2004 757
rect 2070 761 2076 762
rect 2070 757 2071 761
rect 2075 757 2076 761
rect 2070 756 2076 757
rect 2142 761 2148 762
rect 2142 757 2143 761
rect 2147 757 2148 761
rect 2142 756 2148 757
rect 2222 761 2228 762
rect 2222 757 2223 761
rect 2227 757 2228 761
rect 2222 756 2228 757
rect 2302 761 2308 762
rect 2302 757 2303 761
rect 2307 757 2308 761
rect 2302 756 2308 757
rect 2358 761 2364 762
rect 2358 757 2359 761
rect 2363 757 2364 761
rect 2358 756 2364 757
rect 134 735 140 736
rect 134 731 135 735
rect 139 731 140 735
rect 134 730 140 731
rect 190 735 196 736
rect 190 731 191 735
rect 195 731 196 735
rect 190 730 196 731
rect 262 735 268 736
rect 262 731 263 735
rect 267 731 268 735
rect 262 730 268 731
rect 334 735 340 736
rect 334 731 335 735
rect 339 731 340 735
rect 334 730 340 731
rect 398 735 404 736
rect 398 731 399 735
rect 403 731 404 735
rect 398 730 404 731
rect 454 735 460 736
rect 454 731 455 735
rect 459 731 460 735
rect 454 730 460 731
rect 502 735 508 736
rect 502 731 503 735
rect 507 731 508 735
rect 502 730 508 731
rect 542 735 548 736
rect 542 731 543 735
rect 547 731 548 735
rect 542 730 548 731
rect 582 735 588 736
rect 582 731 583 735
rect 587 731 588 735
rect 582 730 588 731
rect 622 735 628 736
rect 622 731 623 735
rect 627 731 628 735
rect 622 730 628 731
rect 670 735 676 736
rect 670 731 671 735
rect 675 731 676 735
rect 670 730 676 731
rect 718 735 724 736
rect 718 731 719 735
rect 723 731 724 735
rect 718 730 724 731
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 814 735 820 736
rect 814 731 815 735
rect 819 731 820 735
rect 814 730 820 731
rect 862 735 868 736
rect 862 731 863 735
rect 867 731 868 735
rect 862 730 868 731
rect 910 735 916 736
rect 910 731 911 735
rect 915 731 916 735
rect 910 730 916 731
rect 1302 731 1308 732
rect 1302 727 1303 731
rect 1307 727 1308 731
rect 1302 726 1308 727
rect 1342 731 1348 732
rect 1342 727 1343 731
rect 1347 727 1348 731
rect 1342 726 1348 727
rect 1406 731 1412 732
rect 1406 727 1407 731
rect 1411 727 1412 731
rect 1406 726 1412 727
rect 1486 731 1492 732
rect 1486 727 1487 731
rect 1491 727 1492 731
rect 1486 726 1492 727
rect 1574 731 1580 732
rect 1574 727 1575 731
rect 1579 727 1580 731
rect 1574 726 1580 727
rect 1662 731 1668 732
rect 1662 727 1663 731
rect 1667 727 1668 731
rect 1662 726 1668 727
rect 1750 731 1756 732
rect 1750 727 1751 731
rect 1755 727 1756 731
rect 1750 726 1756 727
rect 1830 731 1836 732
rect 1830 727 1831 731
rect 1835 727 1836 731
rect 1830 726 1836 727
rect 1910 731 1916 732
rect 1910 727 1911 731
rect 1915 727 1916 731
rect 1910 726 1916 727
rect 1990 731 1996 732
rect 1990 727 1991 731
rect 1995 727 1996 731
rect 1990 726 1996 727
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 727 2084 731
rect 2078 726 2084 727
rect 2174 731 2180 732
rect 2174 727 2175 731
rect 2179 727 2180 731
rect 2174 726 2180 727
rect 2278 731 2284 732
rect 2278 727 2279 731
rect 2283 727 2284 731
rect 2278 726 2284 727
rect 2358 731 2364 732
rect 2358 727 2359 731
rect 2363 727 2364 731
rect 2358 726 2364 727
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 1238 712 1244 713
rect 1238 708 1239 712
rect 1243 708 1244 712
rect 1238 707 1244 708
rect 1278 708 1284 709
rect 1278 704 1279 708
rect 1283 704 1284 708
rect 1278 703 1284 704
rect 2406 708 2412 709
rect 2406 704 2407 708
rect 2411 704 2412 708
rect 2406 703 2412 704
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 1238 695 1244 696
rect 1238 691 1239 695
rect 1243 691 1244 695
rect 1238 690 1244 691
rect 1278 691 1284 692
rect 134 688 140 689
rect 134 684 135 688
rect 139 684 140 688
rect 134 683 140 684
rect 190 688 196 689
rect 190 684 191 688
rect 195 684 196 688
rect 190 683 196 684
rect 262 688 268 689
rect 262 684 263 688
rect 267 684 268 688
rect 262 683 268 684
rect 334 688 340 689
rect 334 684 335 688
rect 339 684 340 688
rect 334 683 340 684
rect 398 688 404 689
rect 398 684 399 688
rect 403 684 404 688
rect 398 683 404 684
rect 454 688 460 689
rect 454 684 455 688
rect 459 684 460 688
rect 454 683 460 684
rect 502 688 508 689
rect 502 684 503 688
rect 507 684 508 688
rect 502 683 508 684
rect 542 688 548 689
rect 542 684 543 688
rect 547 684 548 688
rect 542 683 548 684
rect 582 688 588 689
rect 582 684 583 688
rect 587 684 588 688
rect 582 683 588 684
rect 622 688 628 689
rect 622 684 623 688
rect 627 684 628 688
rect 622 683 628 684
rect 670 688 676 689
rect 670 684 671 688
rect 675 684 676 688
rect 670 683 676 684
rect 718 688 724 689
rect 718 684 719 688
rect 723 684 724 688
rect 718 683 724 684
rect 766 688 772 689
rect 766 684 767 688
rect 771 684 772 688
rect 766 683 772 684
rect 814 688 820 689
rect 814 684 815 688
rect 819 684 820 688
rect 814 683 820 684
rect 862 688 868 689
rect 862 684 863 688
rect 867 684 868 688
rect 862 683 868 684
rect 910 688 916 689
rect 910 684 911 688
rect 915 684 916 688
rect 1278 687 1279 691
rect 1283 687 1284 691
rect 1278 686 1284 687
rect 2406 691 2412 692
rect 2406 687 2407 691
rect 2411 687 2412 691
rect 2406 686 2412 687
rect 910 683 916 684
rect 1302 684 1308 685
rect 1302 680 1303 684
rect 1307 680 1308 684
rect 1302 679 1308 680
rect 1342 684 1348 685
rect 1342 680 1343 684
rect 1347 680 1348 684
rect 1342 679 1348 680
rect 1406 684 1412 685
rect 1406 680 1407 684
rect 1411 680 1412 684
rect 1406 679 1412 680
rect 1486 684 1492 685
rect 1486 680 1487 684
rect 1491 680 1492 684
rect 1486 679 1492 680
rect 1574 684 1580 685
rect 1574 680 1575 684
rect 1579 680 1580 684
rect 1574 679 1580 680
rect 1662 684 1668 685
rect 1662 680 1663 684
rect 1667 680 1668 684
rect 1662 679 1668 680
rect 1750 684 1756 685
rect 1750 680 1751 684
rect 1755 680 1756 684
rect 1750 679 1756 680
rect 1830 684 1836 685
rect 1830 680 1831 684
rect 1835 680 1836 684
rect 1830 679 1836 680
rect 1910 684 1916 685
rect 1910 680 1911 684
rect 1915 680 1916 684
rect 1910 679 1916 680
rect 1990 684 1996 685
rect 1990 680 1991 684
rect 1995 680 1996 684
rect 1990 679 1996 680
rect 2078 684 2084 685
rect 2078 680 2079 684
rect 2083 680 2084 684
rect 2078 679 2084 680
rect 2174 684 2180 685
rect 2174 680 2175 684
rect 2179 680 2180 684
rect 2174 679 2180 680
rect 2278 684 2284 685
rect 2278 680 2279 684
rect 2283 680 2284 684
rect 2278 679 2284 680
rect 2358 684 2364 685
rect 2358 680 2359 684
rect 2363 680 2364 684
rect 2358 679 2364 680
rect 134 672 140 673
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 198 672 204 673
rect 198 668 199 672
rect 203 668 204 672
rect 198 667 204 668
rect 278 672 284 673
rect 278 668 279 672
rect 283 668 284 672
rect 278 667 284 668
rect 350 672 356 673
rect 350 668 351 672
rect 355 668 356 672
rect 350 667 356 668
rect 414 672 420 673
rect 414 668 415 672
rect 419 668 420 672
rect 414 667 420 668
rect 486 672 492 673
rect 486 668 487 672
rect 491 668 492 672
rect 486 667 492 668
rect 558 672 564 673
rect 558 668 559 672
rect 563 668 564 672
rect 558 667 564 668
rect 638 672 644 673
rect 638 668 639 672
rect 643 668 644 672
rect 638 667 644 668
rect 710 672 716 673
rect 710 668 711 672
rect 715 668 716 672
rect 710 667 716 668
rect 782 672 788 673
rect 782 668 783 672
rect 787 668 788 672
rect 782 667 788 668
rect 854 672 860 673
rect 854 668 855 672
rect 859 668 860 672
rect 854 667 860 668
rect 918 672 924 673
rect 918 668 919 672
rect 923 668 924 672
rect 918 667 924 668
rect 982 672 988 673
rect 982 668 983 672
rect 987 668 988 672
rect 982 667 988 668
rect 1038 672 1044 673
rect 1038 668 1039 672
rect 1043 668 1044 672
rect 1038 667 1044 668
rect 1094 672 1100 673
rect 1094 668 1095 672
rect 1099 668 1100 672
rect 1094 667 1100 668
rect 1150 672 1156 673
rect 1150 668 1151 672
rect 1155 668 1156 672
rect 1150 667 1156 668
rect 1190 672 1196 673
rect 1190 668 1191 672
rect 1195 668 1196 672
rect 1190 667 1196 668
rect 1302 668 1308 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 1238 665 1244 666
rect 1238 661 1239 665
rect 1243 661 1244 665
rect 1302 664 1303 668
rect 1307 664 1308 668
rect 1302 663 1308 664
rect 1398 668 1404 669
rect 1398 664 1399 668
rect 1403 664 1404 668
rect 1398 663 1404 664
rect 1510 668 1516 669
rect 1510 664 1511 668
rect 1515 664 1516 668
rect 1510 663 1516 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1726 668 1732 669
rect 1726 664 1727 668
rect 1731 664 1732 668
rect 1726 663 1732 664
rect 1814 668 1820 669
rect 1814 664 1815 668
rect 1819 664 1820 668
rect 1814 663 1820 664
rect 1894 668 1900 669
rect 1894 664 1895 668
rect 1899 664 1900 668
rect 1894 663 1900 664
rect 1974 668 1980 669
rect 1974 664 1975 668
rect 1979 664 1980 668
rect 1974 663 1980 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2110 668 2116 669
rect 2110 664 2111 668
rect 2115 664 2116 668
rect 2110 663 2116 664
rect 2174 668 2180 669
rect 2174 664 2175 668
rect 2179 664 2180 668
rect 2174 663 2180 664
rect 2238 668 2244 669
rect 2238 664 2239 668
rect 2243 664 2244 668
rect 2238 663 2244 664
rect 2310 668 2316 669
rect 2310 664 2311 668
rect 2315 664 2316 668
rect 2310 663 2316 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 1238 660 1244 661
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 110 648 116 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 1238 648 1244 649
rect 1238 644 1239 648
rect 1243 644 1244 648
rect 1238 643 1244 644
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1278 639 1284 640
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 134 625 140 626
rect 134 621 135 625
rect 139 621 140 625
rect 134 620 140 621
rect 198 625 204 626
rect 198 621 199 625
rect 203 621 204 625
rect 198 620 204 621
rect 278 625 284 626
rect 278 621 279 625
rect 283 621 284 625
rect 278 620 284 621
rect 350 625 356 626
rect 350 621 351 625
rect 355 621 356 625
rect 350 620 356 621
rect 414 625 420 626
rect 414 621 415 625
rect 419 621 420 625
rect 414 620 420 621
rect 486 625 492 626
rect 486 621 487 625
rect 491 621 492 625
rect 486 620 492 621
rect 558 625 564 626
rect 558 621 559 625
rect 563 621 564 625
rect 558 620 564 621
rect 638 625 644 626
rect 638 621 639 625
rect 643 621 644 625
rect 638 620 644 621
rect 710 625 716 626
rect 710 621 711 625
rect 715 621 716 625
rect 710 620 716 621
rect 782 625 788 626
rect 782 621 783 625
rect 787 621 788 625
rect 782 620 788 621
rect 854 625 860 626
rect 854 621 855 625
rect 859 621 860 625
rect 854 620 860 621
rect 918 625 924 626
rect 918 621 919 625
rect 923 621 924 625
rect 918 620 924 621
rect 982 625 988 626
rect 982 621 983 625
rect 987 621 988 625
rect 982 620 988 621
rect 1038 625 1044 626
rect 1038 621 1039 625
rect 1043 621 1044 625
rect 1038 620 1044 621
rect 1094 625 1100 626
rect 1094 621 1095 625
rect 1099 621 1100 625
rect 1094 620 1100 621
rect 1150 625 1156 626
rect 1150 621 1151 625
rect 1155 621 1156 625
rect 1150 620 1156 621
rect 1190 625 1196 626
rect 1190 621 1191 625
rect 1195 621 1196 625
rect 1190 620 1196 621
rect 1302 621 1308 622
rect 1302 617 1303 621
rect 1307 617 1308 621
rect 1302 616 1308 617
rect 1398 621 1404 622
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1622 621 1628 622
rect 1622 617 1623 621
rect 1627 617 1628 621
rect 1622 616 1628 617
rect 1726 621 1732 622
rect 1726 617 1727 621
rect 1731 617 1732 621
rect 1726 616 1732 617
rect 1814 621 1820 622
rect 1814 617 1815 621
rect 1819 617 1820 621
rect 1814 616 1820 617
rect 1894 621 1900 622
rect 1894 617 1895 621
rect 1899 617 1900 621
rect 1894 616 1900 617
rect 1974 621 1980 622
rect 1974 617 1975 621
rect 1979 617 1980 621
rect 1974 616 1980 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2110 621 2116 622
rect 2110 617 2111 621
rect 2115 617 2116 621
rect 2110 616 2116 617
rect 2174 621 2180 622
rect 2174 617 2175 621
rect 2179 617 2180 621
rect 2174 616 2180 617
rect 2238 621 2244 622
rect 2238 617 2239 621
rect 2243 617 2244 621
rect 2238 616 2244 617
rect 2310 621 2316 622
rect 2310 617 2311 621
rect 2315 617 2316 621
rect 2310 616 2316 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 134 587 140 588
rect 134 583 135 587
rect 139 583 140 587
rect 134 582 140 583
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 270 587 276 588
rect 270 583 271 587
rect 275 583 276 587
rect 270 582 276 583
rect 358 587 364 588
rect 358 583 359 587
rect 363 583 364 587
rect 358 582 364 583
rect 446 587 452 588
rect 446 583 447 587
rect 451 583 452 587
rect 446 582 452 583
rect 534 587 540 588
rect 534 583 535 587
rect 539 583 540 587
rect 534 582 540 583
rect 622 587 628 588
rect 622 583 623 587
rect 627 583 628 587
rect 622 582 628 583
rect 702 587 708 588
rect 702 583 703 587
rect 707 583 708 587
rect 702 582 708 583
rect 782 587 788 588
rect 782 583 783 587
rect 787 583 788 587
rect 782 582 788 583
rect 854 587 860 588
rect 854 583 855 587
rect 859 583 860 587
rect 854 582 860 583
rect 918 587 924 588
rect 918 583 919 587
rect 923 583 924 587
rect 918 582 924 583
rect 974 587 980 588
rect 974 583 975 587
rect 979 583 980 587
rect 974 582 980 583
rect 1022 587 1028 588
rect 1022 583 1023 587
rect 1027 583 1028 587
rect 1022 582 1028 583
rect 1078 587 1084 588
rect 1078 583 1079 587
rect 1083 583 1084 587
rect 1078 582 1084 583
rect 1134 587 1140 588
rect 1134 583 1135 587
rect 1139 583 1140 587
rect 1134 582 1140 583
rect 1190 587 1196 588
rect 1190 583 1191 587
rect 1195 583 1196 587
rect 1190 582 1196 583
rect 1414 587 1420 588
rect 1414 583 1415 587
rect 1419 583 1420 587
rect 1414 582 1420 583
rect 1454 587 1460 588
rect 1454 583 1455 587
rect 1459 583 1460 587
rect 1454 582 1460 583
rect 1494 587 1500 588
rect 1494 583 1495 587
rect 1499 583 1500 587
rect 1494 582 1500 583
rect 1542 587 1548 588
rect 1542 583 1543 587
rect 1547 583 1548 587
rect 1542 582 1548 583
rect 1598 587 1604 588
rect 1598 583 1599 587
rect 1603 583 1604 587
rect 1598 582 1604 583
rect 1662 587 1668 588
rect 1662 583 1663 587
rect 1667 583 1668 587
rect 1662 582 1668 583
rect 1726 587 1732 588
rect 1726 583 1727 587
rect 1731 583 1732 587
rect 1726 582 1732 583
rect 1790 587 1796 588
rect 1790 583 1791 587
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1846 587 1852 588
rect 1846 583 1847 587
rect 1851 583 1852 587
rect 1846 582 1852 583
rect 1910 587 1916 588
rect 1910 583 1911 587
rect 1915 583 1916 587
rect 1910 582 1916 583
rect 1974 587 1980 588
rect 1974 583 1975 587
rect 1979 583 1980 587
rect 1974 582 1980 583
rect 2046 587 2052 588
rect 2046 583 2047 587
rect 2051 583 2052 587
rect 2046 582 2052 583
rect 2118 587 2124 588
rect 2118 583 2119 587
rect 2123 583 2124 587
rect 2118 582 2124 583
rect 2198 587 2204 588
rect 2198 583 2199 587
rect 2203 583 2204 587
rect 2198 582 2204 583
rect 2286 587 2292 588
rect 2286 583 2287 587
rect 2291 583 2292 587
rect 2286 582 2292 583
rect 2358 587 2364 588
rect 2358 583 2359 587
rect 2363 583 2364 587
rect 2358 582 2364 583
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 110 559 116 560
rect 1238 564 1244 565
rect 1238 560 1239 564
rect 1243 560 1244 564
rect 1238 559 1244 560
rect 1278 564 1284 565
rect 1278 560 1279 564
rect 1283 560 1284 564
rect 1278 559 1284 560
rect 2406 564 2412 565
rect 2406 560 2407 564
rect 2411 560 2412 564
rect 2406 559 2412 560
rect 110 547 116 548
rect 110 543 111 547
rect 115 543 116 547
rect 110 542 116 543
rect 1238 547 1244 548
rect 1238 543 1239 547
rect 1243 543 1244 547
rect 1238 542 1244 543
rect 1278 547 1284 548
rect 1278 543 1279 547
rect 1283 543 1284 547
rect 1278 542 1284 543
rect 2406 547 2412 548
rect 2406 543 2407 547
rect 2411 543 2412 547
rect 2406 542 2412 543
rect 134 540 140 541
rect 134 536 135 540
rect 139 536 140 540
rect 134 535 140 536
rect 190 540 196 541
rect 190 536 191 540
rect 195 536 196 540
rect 190 535 196 536
rect 270 540 276 541
rect 270 536 271 540
rect 275 536 276 540
rect 270 535 276 536
rect 358 540 364 541
rect 358 536 359 540
rect 363 536 364 540
rect 358 535 364 536
rect 446 540 452 541
rect 446 536 447 540
rect 451 536 452 540
rect 446 535 452 536
rect 534 540 540 541
rect 534 536 535 540
rect 539 536 540 540
rect 534 535 540 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 782 540 788 541
rect 782 536 783 540
rect 787 536 788 540
rect 782 535 788 536
rect 854 540 860 541
rect 854 536 855 540
rect 859 536 860 540
rect 854 535 860 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 974 540 980 541
rect 974 536 975 540
rect 979 536 980 540
rect 974 535 980 536
rect 1022 540 1028 541
rect 1022 536 1023 540
rect 1027 536 1028 540
rect 1022 535 1028 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 1134 540 1140 541
rect 1134 536 1135 540
rect 1139 536 1140 540
rect 1134 535 1140 536
rect 1190 540 1196 541
rect 1190 536 1191 540
rect 1195 536 1196 540
rect 1190 535 1196 536
rect 1414 540 1420 541
rect 1414 536 1415 540
rect 1419 536 1420 540
rect 1414 535 1420 536
rect 1454 540 1460 541
rect 1454 536 1455 540
rect 1459 536 1460 540
rect 1454 535 1460 536
rect 1494 540 1500 541
rect 1494 536 1495 540
rect 1499 536 1500 540
rect 1494 535 1500 536
rect 1542 540 1548 541
rect 1542 536 1543 540
rect 1547 536 1548 540
rect 1542 535 1548 536
rect 1598 540 1604 541
rect 1598 536 1599 540
rect 1603 536 1604 540
rect 1598 535 1604 536
rect 1662 540 1668 541
rect 1662 536 1663 540
rect 1667 536 1668 540
rect 1662 535 1668 536
rect 1726 540 1732 541
rect 1726 536 1727 540
rect 1731 536 1732 540
rect 1726 535 1732 536
rect 1790 540 1796 541
rect 1790 536 1791 540
rect 1795 536 1796 540
rect 1790 535 1796 536
rect 1846 540 1852 541
rect 1846 536 1847 540
rect 1851 536 1852 540
rect 1846 535 1852 536
rect 1910 540 1916 541
rect 1910 536 1911 540
rect 1915 536 1916 540
rect 1910 535 1916 536
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 1974 535 1980 536
rect 2046 540 2052 541
rect 2046 536 2047 540
rect 2051 536 2052 540
rect 2046 535 2052 536
rect 2118 540 2124 541
rect 2118 536 2119 540
rect 2123 536 2124 540
rect 2118 535 2124 536
rect 2198 540 2204 541
rect 2198 536 2199 540
rect 2203 536 2204 540
rect 2198 535 2204 536
rect 2286 540 2292 541
rect 2286 536 2287 540
rect 2291 536 2292 540
rect 2286 535 2292 536
rect 2358 540 2364 541
rect 2358 536 2359 540
rect 2363 536 2364 540
rect 2358 535 2364 536
rect 1302 528 1308 529
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1374 528 1380 529
rect 1374 524 1375 528
rect 1379 524 1380 528
rect 1374 523 1380 524
rect 1478 528 1484 529
rect 1478 524 1479 528
rect 1483 524 1484 528
rect 1478 523 1484 524
rect 1582 528 1588 529
rect 1582 524 1583 528
rect 1587 524 1588 528
rect 1582 523 1588 524
rect 1694 528 1700 529
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1798 528 1804 529
rect 1798 524 1799 528
rect 1803 524 1804 528
rect 1798 523 1804 524
rect 1902 528 1908 529
rect 1902 524 1903 528
rect 1907 524 1908 528
rect 1902 523 1908 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2190 528 2196 529
rect 2190 524 2191 528
rect 2195 524 2196 528
rect 2190 523 2196 524
rect 2286 528 2292 529
rect 2286 524 2287 528
rect 2291 524 2292 528
rect 2286 523 2292 524
rect 2358 528 2364 529
rect 2358 524 2359 528
rect 2363 524 2364 528
rect 2358 523 2364 524
rect 1278 521 1284 522
rect 134 520 140 521
rect 134 516 135 520
rect 139 516 140 520
rect 134 515 140 516
rect 190 520 196 521
rect 190 516 191 520
rect 195 516 196 520
rect 190 515 196 516
rect 262 520 268 521
rect 262 516 263 520
rect 267 516 268 520
rect 262 515 268 516
rect 334 520 340 521
rect 334 516 335 520
rect 339 516 340 520
rect 334 515 340 516
rect 414 520 420 521
rect 414 516 415 520
rect 419 516 420 520
rect 414 515 420 516
rect 494 520 500 521
rect 494 516 495 520
rect 499 516 500 520
rect 494 515 500 516
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 646 520 652 521
rect 646 516 647 520
rect 651 516 652 520
rect 646 515 652 516
rect 718 520 724 521
rect 718 516 719 520
rect 723 516 724 520
rect 718 515 724 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 846 520 852 521
rect 846 516 847 520
rect 851 516 852 520
rect 846 515 852 516
rect 902 520 908 521
rect 902 516 903 520
rect 907 516 908 520
rect 902 515 908 516
rect 958 520 964 521
rect 958 516 959 520
rect 963 516 964 520
rect 958 515 964 516
rect 1022 520 1028 521
rect 1022 516 1023 520
rect 1027 516 1028 520
rect 1022 515 1028 516
rect 1086 520 1092 521
rect 1086 516 1087 520
rect 1091 516 1092 520
rect 1086 515 1092 516
rect 1150 520 1156 521
rect 1150 516 1151 520
rect 1155 516 1156 520
rect 1150 515 1156 516
rect 1190 520 1196 521
rect 1190 516 1191 520
rect 1195 516 1196 520
rect 1278 517 1279 521
rect 1283 517 1284 521
rect 1278 516 1284 517
rect 2406 521 2412 522
rect 2406 517 2407 521
rect 2411 517 2412 521
rect 2406 516 2412 517
rect 1190 515 1196 516
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 1238 513 1244 514
rect 1238 509 1239 513
rect 1243 509 1244 513
rect 1238 508 1244 509
rect 1278 504 1284 505
rect 1278 500 1279 504
rect 1283 500 1284 504
rect 1278 499 1284 500
rect 2406 504 2412 505
rect 2406 500 2407 504
rect 2411 500 2412 504
rect 2406 499 2412 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1238 496 1244 497
rect 1238 492 1239 496
rect 1243 492 1244 496
rect 1238 491 1244 492
rect 1302 481 1308 482
rect 1302 477 1303 481
rect 1307 477 1308 481
rect 1302 476 1308 477
rect 1374 481 1380 482
rect 1374 477 1375 481
rect 1379 477 1380 481
rect 1374 476 1380 477
rect 1478 481 1484 482
rect 1478 477 1479 481
rect 1483 477 1484 481
rect 1478 476 1484 477
rect 1582 481 1588 482
rect 1582 477 1583 481
rect 1587 477 1588 481
rect 1582 476 1588 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1798 481 1804 482
rect 1798 477 1799 481
rect 1803 477 1804 481
rect 1798 476 1804 477
rect 1902 481 1908 482
rect 1902 477 1903 481
rect 1907 477 1908 481
rect 1902 476 1908 477
rect 2006 481 2012 482
rect 2006 477 2007 481
rect 2011 477 2012 481
rect 2006 476 2012 477
rect 2102 481 2108 482
rect 2102 477 2103 481
rect 2107 477 2108 481
rect 2102 476 2108 477
rect 2190 481 2196 482
rect 2190 477 2191 481
rect 2195 477 2196 481
rect 2190 476 2196 477
rect 2286 481 2292 482
rect 2286 477 2287 481
rect 2291 477 2292 481
rect 2286 476 2292 477
rect 2358 481 2364 482
rect 2358 477 2359 481
rect 2363 477 2364 481
rect 2358 476 2364 477
rect 134 473 140 474
rect 134 469 135 473
rect 139 469 140 473
rect 134 468 140 469
rect 190 473 196 474
rect 190 469 191 473
rect 195 469 196 473
rect 190 468 196 469
rect 262 473 268 474
rect 262 469 263 473
rect 267 469 268 473
rect 262 468 268 469
rect 334 473 340 474
rect 334 469 335 473
rect 339 469 340 473
rect 334 468 340 469
rect 414 473 420 474
rect 414 469 415 473
rect 419 469 420 473
rect 414 468 420 469
rect 494 473 500 474
rect 494 469 495 473
rect 499 469 500 473
rect 494 468 500 469
rect 574 473 580 474
rect 574 469 575 473
rect 579 469 580 473
rect 574 468 580 469
rect 646 473 652 474
rect 646 469 647 473
rect 651 469 652 473
rect 646 468 652 469
rect 718 473 724 474
rect 718 469 719 473
rect 723 469 724 473
rect 718 468 724 469
rect 782 473 788 474
rect 782 469 783 473
rect 787 469 788 473
rect 782 468 788 469
rect 846 473 852 474
rect 846 469 847 473
rect 851 469 852 473
rect 846 468 852 469
rect 902 473 908 474
rect 902 469 903 473
rect 907 469 908 473
rect 902 468 908 469
rect 958 473 964 474
rect 958 469 959 473
rect 963 469 964 473
rect 958 468 964 469
rect 1022 473 1028 474
rect 1022 469 1023 473
rect 1027 469 1028 473
rect 1022 468 1028 469
rect 1086 473 1092 474
rect 1086 469 1087 473
rect 1091 469 1092 473
rect 1086 468 1092 469
rect 1150 473 1156 474
rect 1150 469 1151 473
rect 1155 469 1156 473
rect 1150 468 1156 469
rect 1190 473 1196 474
rect 1190 469 1191 473
rect 1195 469 1196 473
rect 1190 468 1196 469
rect 1302 447 1308 448
rect 182 443 188 444
rect 182 439 183 443
rect 187 439 188 443
rect 182 438 188 439
rect 222 443 228 444
rect 222 439 223 443
rect 227 439 228 443
rect 222 438 228 439
rect 262 443 268 444
rect 262 439 263 443
rect 267 439 268 443
rect 262 438 268 439
rect 310 443 316 444
rect 310 439 311 443
rect 315 439 316 443
rect 310 438 316 439
rect 366 443 372 444
rect 366 439 367 443
rect 371 439 372 443
rect 366 438 372 439
rect 430 443 436 444
rect 430 439 431 443
rect 435 439 436 443
rect 430 438 436 439
rect 494 443 500 444
rect 494 439 495 443
rect 499 439 500 443
rect 494 438 500 439
rect 558 443 564 444
rect 558 439 559 443
rect 563 439 564 443
rect 558 438 564 439
rect 614 443 620 444
rect 614 439 615 443
rect 619 439 620 443
rect 614 438 620 439
rect 670 443 676 444
rect 670 439 671 443
rect 675 439 676 443
rect 670 438 676 439
rect 718 443 724 444
rect 718 439 719 443
rect 723 439 724 443
rect 718 438 724 439
rect 774 443 780 444
rect 774 439 775 443
rect 779 439 780 443
rect 774 438 780 439
rect 830 443 836 444
rect 830 439 831 443
rect 835 439 836 443
rect 830 438 836 439
rect 886 443 892 444
rect 886 439 887 443
rect 891 439 892 443
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1398 447 1404 448
rect 1398 443 1399 447
rect 1403 443 1404 447
rect 1398 442 1404 443
rect 1462 447 1468 448
rect 1462 443 1463 447
rect 1467 443 1468 447
rect 1462 442 1468 443
rect 1526 447 1532 448
rect 1526 443 1527 447
rect 1531 443 1532 447
rect 1526 442 1532 443
rect 1590 447 1596 448
rect 1590 443 1591 447
rect 1595 443 1596 447
rect 1590 442 1596 443
rect 1662 447 1668 448
rect 1662 443 1663 447
rect 1667 443 1668 447
rect 1662 442 1668 443
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1814 447 1820 448
rect 1814 443 1815 447
rect 1819 443 1820 447
rect 1814 442 1820 443
rect 1894 447 1900 448
rect 1894 443 1895 447
rect 1899 443 1900 447
rect 1894 442 1900 443
rect 1974 447 1980 448
rect 1974 443 1975 447
rect 1979 443 1980 447
rect 1974 442 1980 443
rect 2054 447 2060 448
rect 2054 443 2055 447
rect 2059 443 2060 447
rect 2054 442 2060 443
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2214 447 2220 448
rect 2214 443 2215 447
rect 2219 443 2220 447
rect 2214 442 2220 443
rect 2294 447 2300 448
rect 2294 443 2295 447
rect 2299 443 2300 447
rect 2294 442 2300 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 886 438 892 439
rect 1278 424 1284 425
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 1238 420 1244 421
rect 1238 416 1239 420
rect 1243 416 1244 420
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1278 419 1284 420
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2406 419 2412 420
rect 1238 415 1244 416
rect 1278 407 1284 408
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 110 398 116 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1278 402 1284 403
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 1238 398 1244 399
rect 1302 400 1308 401
rect 182 396 188 397
rect 182 392 183 396
rect 187 392 188 396
rect 182 391 188 392
rect 222 396 228 397
rect 222 392 223 396
rect 227 392 228 396
rect 222 391 228 392
rect 262 396 268 397
rect 262 392 263 396
rect 267 392 268 396
rect 262 391 268 392
rect 310 396 316 397
rect 310 392 311 396
rect 315 392 316 396
rect 310 391 316 392
rect 366 396 372 397
rect 366 392 367 396
rect 371 392 372 396
rect 366 391 372 392
rect 430 396 436 397
rect 430 392 431 396
rect 435 392 436 396
rect 430 391 436 392
rect 494 396 500 397
rect 494 392 495 396
rect 499 392 500 396
rect 494 391 500 392
rect 558 396 564 397
rect 558 392 559 396
rect 563 392 564 396
rect 558 391 564 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 718 396 724 397
rect 718 392 719 396
rect 723 392 724 396
rect 718 391 724 392
rect 774 396 780 397
rect 774 392 775 396
rect 779 392 780 396
rect 774 391 780 392
rect 830 396 836 397
rect 830 392 831 396
rect 835 392 836 396
rect 830 391 836 392
rect 886 396 892 397
rect 886 392 887 396
rect 891 392 892 396
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1398 400 1404 401
rect 1398 396 1399 400
rect 1403 396 1404 400
rect 1398 395 1404 396
rect 1462 400 1468 401
rect 1462 396 1463 400
rect 1467 396 1468 400
rect 1462 395 1468 396
rect 1526 400 1532 401
rect 1526 396 1527 400
rect 1531 396 1532 400
rect 1526 395 1532 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1662 400 1668 401
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1814 400 1820 401
rect 1814 396 1815 400
rect 1819 396 1820 400
rect 1814 395 1820 396
rect 1894 400 1900 401
rect 1894 396 1895 400
rect 1899 396 1900 400
rect 1894 395 1900 396
rect 1974 400 1980 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 2054 400 2060 401
rect 2054 396 2055 400
rect 2059 396 2060 400
rect 2054 395 2060 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2214 400 2220 401
rect 2214 396 2215 400
rect 2219 396 2220 400
rect 2214 395 2220 396
rect 2294 400 2300 401
rect 2294 396 2295 400
rect 2299 396 2300 400
rect 2294 395 2300 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 886 391 892 392
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 174 384 180 385
rect 174 380 175 384
rect 179 380 180 384
rect 174 379 180 380
rect 230 384 236 385
rect 230 380 231 384
rect 235 380 236 384
rect 230 379 236 380
rect 286 384 292 385
rect 286 380 287 384
rect 291 380 292 384
rect 286 379 292 380
rect 342 384 348 385
rect 342 380 343 384
rect 347 380 348 384
rect 342 379 348 380
rect 390 384 396 385
rect 390 380 391 384
rect 395 380 396 384
rect 390 379 396 380
rect 438 384 444 385
rect 438 380 439 384
rect 443 380 444 384
rect 438 379 444 380
rect 486 384 492 385
rect 486 380 487 384
rect 491 380 492 384
rect 486 379 492 380
rect 534 384 540 385
rect 534 380 535 384
rect 539 380 540 384
rect 534 379 540 380
rect 582 384 588 385
rect 582 380 583 384
rect 587 380 588 384
rect 582 379 588 380
rect 630 384 636 385
rect 630 380 631 384
rect 635 380 636 384
rect 630 379 636 380
rect 678 384 684 385
rect 678 380 679 384
rect 683 380 684 384
rect 678 379 684 380
rect 726 384 732 385
rect 726 380 727 384
rect 731 380 732 384
rect 726 379 732 380
rect 774 384 780 385
rect 774 380 775 384
rect 779 380 780 384
rect 774 379 780 380
rect 1446 384 1452 385
rect 1446 380 1447 384
rect 1451 380 1452 384
rect 1446 379 1452 380
rect 1486 384 1492 385
rect 1486 380 1487 384
rect 1491 380 1492 384
rect 1486 379 1492 380
rect 1534 384 1540 385
rect 1534 380 1535 384
rect 1539 380 1540 384
rect 1534 379 1540 380
rect 1590 384 1596 385
rect 1590 380 1591 384
rect 1595 380 1596 384
rect 1590 379 1596 380
rect 1662 384 1668 385
rect 1662 380 1663 384
rect 1667 380 1668 384
rect 1662 379 1668 380
rect 1734 384 1740 385
rect 1734 380 1735 384
rect 1739 380 1740 384
rect 1734 379 1740 380
rect 1814 384 1820 385
rect 1814 380 1815 384
rect 1819 380 1820 384
rect 1814 379 1820 380
rect 1894 384 1900 385
rect 1894 380 1895 384
rect 1899 380 1900 384
rect 1894 379 1900 380
rect 1966 384 1972 385
rect 1966 380 1967 384
rect 1971 380 1972 384
rect 1966 379 1972 380
rect 2038 384 2044 385
rect 2038 380 2039 384
rect 2043 380 2044 384
rect 2038 379 2044 380
rect 2110 384 2116 385
rect 2110 380 2111 384
rect 2115 380 2116 384
rect 2110 379 2116 380
rect 2174 384 2180 385
rect 2174 380 2175 384
rect 2179 380 2180 384
rect 2174 379 2180 380
rect 2238 384 2244 385
rect 2238 380 2239 384
rect 2243 380 2244 384
rect 2238 379 2244 380
rect 2302 384 2308 385
rect 2302 380 2303 384
rect 2307 380 2308 384
rect 2302 379 2308 380
rect 2358 384 2364 385
rect 2358 380 2359 384
rect 2363 380 2364 384
rect 2358 379 2364 380
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 1238 377 1244 378
rect 1238 373 1239 377
rect 1243 373 1244 377
rect 1238 372 1244 373
rect 1278 377 1284 378
rect 1278 373 1279 377
rect 1283 373 1284 377
rect 1278 372 1284 373
rect 2406 377 2412 378
rect 2406 373 2407 377
rect 2411 373 2412 377
rect 2406 372 2412 373
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 110 355 116 356
rect 1238 360 1244 361
rect 1238 356 1239 360
rect 1243 356 1244 360
rect 1238 355 1244 356
rect 1278 360 1284 361
rect 1278 356 1279 360
rect 1283 356 1284 360
rect 1278 355 1284 356
rect 2406 360 2412 361
rect 2406 356 2407 360
rect 2411 356 2412 360
rect 2406 355 2412 356
rect 134 337 140 338
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 174 337 180 338
rect 174 333 175 337
rect 179 333 180 337
rect 174 332 180 333
rect 230 337 236 338
rect 230 333 231 337
rect 235 333 236 337
rect 230 332 236 333
rect 286 337 292 338
rect 286 333 287 337
rect 291 333 292 337
rect 286 332 292 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 390 337 396 338
rect 390 333 391 337
rect 395 333 396 337
rect 390 332 396 333
rect 438 337 444 338
rect 438 333 439 337
rect 443 333 444 337
rect 438 332 444 333
rect 486 337 492 338
rect 486 333 487 337
rect 491 333 492 337
rect 486 332 492 333
rect 534 337 540 338
rect 534 333 535 337
rect 539 333 540 337
rect 534 332 540 333
rect 582 337 588 338
rect 582 333 583 337
rect 587 333 588 337
rect 582 332 588 333
rect 630 337 636 338
rect 630 333 631 337
rect 635 333 636 337
rect 630 332 636 333
rect 678 337 684 338
rect 678 333 679 337
rect 683 333 684 337
rect 678 332 684 333
rect 726 337 732 338
rect 726 333 727 337
rect 731 333 732 337
rect 726 332 732 333
rect 774 337 780 338
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 1446 337 1452 338
rect 1446 333 1447 337
rect 1451 333 1452 337
rect 1446 332 1452 333
rect 1486 337 1492 338
rect 1486 333 1487 337
rect 1491 333 1492 337
rect 1486 332 1492 333
rect 1534 337 1540 338
rect 1534 333 1535 337
rect 1539 333 1540 337
rect 1534 332 1540 333
rect 1590 337 1596 338
rect 1590 333 1591 337
rect 1595 333 1596 337
rect 1590 332 1596 333
rect 1662 337 1668 338
rect 1662 333 1663 337
rect 1667 333 1668 337
rect 1662 332 1668 333
rect 1734 337 1740 338
rect 1734 333 1735 337
rect 1739 333 1740 337
rect 1734 332 1740 333
rect 1814 337 1820 338
rect 1814 333 1815 337
rect 1819 333 1820 337
rect 1814 332 1820 333
rect 1894 337 1900 338
rect 1894 333 1895 337
rect 1899 333 1900 337
rect 1894 332 1900 333
rect 1966 337 1972 338
rect 1966 333 1967 337
rect 1971 333 1972 337
rect 1966 332 1972 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2110 337 2116 338
rect 2110 333 2111 337
rect 2115 333 2116 337
rect 2110 332 2116 333
rect 2174 337 2180 338
rect 2174 333 2175 337
rect 2179 333 2180 337
rect 2174 332 2180 333
rect 2238 337 2244 338
rect 2238 333 2239 337
rect 2243 333 2244 337
rect 2238 332 2244 333
rect 2302 337 2308 338
rect 2302 333 2303 337
rect 2307 333 2308 337
rect 2302 332 2308 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 134 303 140 304
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 182 303 188 304
rect 182 299 183 303
rect 187 299 188 303
rect 182 298 188 299
rect 254 303 260 304
rect 254 299 255 303
rect 259 299 260 303
rect 254 298 260 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 446 303 452 304
rect 446 299 447 303
rect 451 299 452 303
rect 446 298 452 299
rect 502 303 508 304
rect 502 299 503 303
rect 507 299 508 303
rect 502 298 508 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 550 298 556 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 630 303 636 304
rect 630 299 631 303
rect 635 299 636 303
rect 630 298 636 299
rect 678 303 684 304
rect 678 299 679 303
rect 683 299 684 303
rect 678 298 684 299
rect 726 303 732 304
rect 726 299 727 303
rect 731 299 732 303
rect 726 298 732 299
rect 774 303 780 304
rect 774 299 775 303
rect 779 299 780 303
rect 774 298 780 299
rect 822 303 828 304
rect 822 299 823 303
rect 827 299 828 303
rect 822 298 828 299
rect 870 303 876 304
rect 870 299 871 303
rect 875 299 876 303
rect 870 298 876 299
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 918 298 924 299
rect 1494 303 1500 304
rect 1494 299 1495 303
rect 1499 299 1500 303
rect 1494 298 1500 299
rect 1534 303 1540 304
rect 1534 299 1535 303
rect 1539 299 1540 303
rect 1534 298 1540 299
rect 1574 303 1580 304
rect 1574 299 1575 303
rect 1579 299 1580 303
rect 1574 298 1580 299
rect 1614 303 1620 304
rect 1614 299 1615 303
rect 1619 299 1620 303
rect 1614 298 1620 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1694 303 1700 304
rect 1694 299 1695 303
rect 1699 299 1700 303
rect 1694 298 1700 299
rect 1742 303 1748 304
rect 1742 299 1743 303
rect 1747 299 1748 303
rect 1742 298 1748 299
rect 1798 303 1804 304
rect 1798 299 1799 303
rect 1803 299 1804 303
rect 1798 298 1804 299
rect 1862 303 1868 304
rect 1862 299 1863 303
rect 1867 299 1868 303
rect 1862 298 1868 299
rect 1934 303 1940 304
rect 1934 299 1935 303
rect 1939 299 1940 303
rect 1934 298 1940 299
rect 2006 303 2012 304
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2070 303 2076 304
rect 2070 299 2071 303
rect 2075 299 2076 303
rect 2070 298 2076 299
rect 2134 303 2140 304
rect 2134 299 2135 303
rect 2139 299 2140 303
rect 2134 298 2140 299
rect 2190 303 2196 304
rect 2190 299 2191 303
rect 2195 299 2196 303
rect 2190 298 2196 299
rect 2254 303 2260 304
rect 2254 299 2255 303
rect 2259 299 2260 303
rect 2254 298 2260 299
rect 2318 303 2324 304
rect 2318 299 2319 303
rect 2323 299 2324 303
rect 2318 298 2324 299
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 110 280 116 281
rect 110 276 111 280
rect 115 276 116 280
rect 110 275 116 276
rect 1238 280 1244 281
rect 1238 276 1239 280
rect 1243 276 1244 280
rect 1238 275 1244 276
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 1278 275 1284 276
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2406 275 2412 276
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 1238 263 1244 264
rect 1238 259 1239 263
rect 1243 259 1244 263
rect 1238 258 1244 259
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1278 258 1284 259
rect 2406 263 2412 264
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 134 256 140 257
rect 134 252 135 256
rect 139 252 140 256
rect 134 251 140 252
rect 182 256 188 257
rect 182 252 183 256
rect 187 252 188 256
rect 182 251 188 252
rect 254 256 260 257
rect 254 252 255 256
rect 259 252 260 256
rect 254 251 260 252
rect 326 256 332 257
rect 326 252 327 256
rect 331 252 332 256
rect 326 251 332 252
rect 390 256 396 257
rect 390 252 391 256
rect 395 252 396 256
rect 390 251 396 252
rect 446 256 452 257
rect 446 252 447 256
rect 451 252 452 256
rect 446 251 452 252
rect 502 256 508 257
rect 502 252 503 256
rect 507 252 508 256
rect 502 251 508 252
rect 550 256 556 257
rect 550 252 551 256
rect 555 252 556 256
rect 550 251 556 252
rect 590 256 596 257
rect 590 252 591 256
rect 595 252 596 256
rect 590 251 596 252
rect 630 256 636 257
rect 630 252 631 256
rect 635 252 636 256
rect 630 251 636 252
rect 678 256 684 257
rect 678 252 679 256
rect 683 252 684 256
rect 678 251 684 252
rect 726 256 732 257
rect 726 252 727 256
rect 731 252 732 256
rect 726 251 732 252
rect 774 256 780 257
rect 774 252 775 256
rect 779 252 780 256
rect 774 251 780 252
rect 822 256 828 257
rect 822 252 823 256
rect 827 252 828 256
rect 822 251 828 252
rect 870 256 876 257
rect 870 252 871 256
rect 875 252 876 256
rect 870 251 876 252
rect 918 256 924 257
rect 918 252 919 256
rect 923 252 924 256
rect 918 251 924 252
rect 1494 256 1500 257
rect 1494 252 1495 256
rect 1499 252 1500 256
rect 1494 251 1500 252
rect 1534 256 1540 257
rect 1534 252 1535 256
rect 1539 252 1540 256
rect 1534 251 1540 252
rect 1574 256 1580 257
rect 1574 252 1575 256
rect 1579 252 1580 256
rect 1574 251 1580 252
rect 1614 256 1620 257
rect 1614 252 1615 256
rect 1619 252 1620 256
rect 1614 251 1620 252
rect 1654 256 1660 257
rect 1654 252 1655 256
rect 1659 252 1660 256
rect 1654 251 1660 252
rect 1694 256 1700 257
rect 1694 252 1695 256
rect 1699 252 1700 256
rect 1694 251 1700 252
rect 1742 256 1748 257
rect 1742 252 1743 256
rect 1747 252 1748 256
rect 1742 251 1748 252
rect 1798 256 1804 257
rect 1798 252 1799 256
rect 1803 252 1804 256
rect 1798 251 1804 252
rect 1862 256 1868 257
rect 1862 252 1863 256
rect 1867 252 1868 256
rect 1862 251 1868 252
rect 1934 256 1940 257
rect 1934 252 1935 256
rect 1939 252 1940 256
rect 1934 251 1940 252
rect 2006 256 2012 257
rect 2006 252 2007 256
rect 2011 252 2012 256
rect 2006 251 2012 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2134 256 2140 257
rect 2134 252 2135 256
rect 2139 252 2140 256
rect 2134 251 2140 252
rect 2190 256 2196 257
rect 2190 252 2191 256
rect 2195 252 2196 256
rect 2190 251 2196 252
rect 2254 256 2260 257
rect 2254 252 2255 256
rect 2259 252 2260 256
rect 2254 251 2260 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 1366 240 1372 241
rect 134 236 140 237
rect 134 232 135 236
rect 139 232 140 236
rect 134 231 140 232
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 246 236 252 237
rect 246 232 247 236
rect 251 232 252 236
rect 246 231 252 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 414 236 420 237
rect 414 232 415 236
rect 419 232 420 236
rect 414 231 420 232
rect 494 236 500 237
rect 494 232 495 236
rect 499 232 500 236
rect 494 231 500 232
rect 574 236 580 237
rect 574 232 575 236
rect 579 232 580 236
rect 574 231 580 232
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 726 236 732 237
rect 726 232 727 236
rect 731 232 732 236
rect 726 231 732 232
rect 790 236 796 237
rect 790 232 791 236
rect 795 232 796 236
rect 790 231 796 232
rect 846 236 852 237
rect 846 232 847 236
rect 851 232 852 236
rect 846 231 852 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 958 236 964 237
rect 958 232 959 236
rect 963 232 964 236
rect 958 231 964 232
rect 1022 236 1028 237
rect 1022 232 1023 236
rect 1027 232 1028 236
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1446 240 1452 241
rect 1446 236 1447 240
rect 1451 236 1452 240
rect 1446 235 1452 236
rect 1494 240 1500 241
rect 1494 236 1495 240
rect 1499 236 1500 240
rect 1494 235 1500 236
rect 1550 240 1556 241
rect 1550 236 1551 240
rect 1555 236 1556 240
rect 1550 235 1556 236
rect 1606 240 1612 241
rect 1606 236 1607 240
rect 1611 236 1612 240
rect 1606 235 1612 236
rect 1670 240 1676 241
rect 1670 236 1671 240
rect 1675 236 1676 240
rect 1670 235 1676 236
rect 1734 240 1740 241
rect 1734 236 1735 240
rect 1739 236 1740 240
rect 1734 235 1740 236
rect 1806 240 1812 241
rect 1806 236 1807 240
rect 1811 236 1812 240
rect 1806 235 1812 236
rect 1886 240 1892 241
rect 1886 236 1887 240
rect 1891 236 1892 240
rect 1886 235 1892 236
rect 1974 240 1980 241
rect 1974 236 1975 240
rect 1979 236 1980 240
rect 1974 235 1980 236
rect 2070 240 2076 241
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2166 240 2172 241
rect 2166 236 2167 240
rect 2171 236 2172 240
rect 2166 235 2172 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 1022 231 1028 232
rect 1278 233 1284 234
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 1238 229 1244 230
rect 1238 225 1239 229
rect 1243 225 1244 229
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 1238 224 1244 225
rect 1278 216 1284 217
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 110 207 116 208
rect 1238 212 1244 213
rect 1238 208 1239 212
rect 1243 208 1244 212
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1278 211 1284 212
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 1238 207 1244 208
rect 1366 193 1372 194
rect 134 189 140 190
rect 134 185 135 189
rect 139 185 140 189
rect 134 184 140 185
rect 174 189 180 190
rect 174 185 175 189
rect 179 185 180 189
rect 174 184 180 185
rect 246 189 252 190
rect 246 185 247 189
rect 251 185 252 189
rect 246 184 252 185
rect 326 189 332 190
rect 326 185 327 189
rect 331 185 332 189
rect 326 184 332 185
rect 414 189 420 190
rect 414 185 415 189
rect 419 185 420 189
rect 414 184 420 185
rect 494 189 500 190
rect 494 185 495 189
rect 499 185 500 189
rect 494 184 500 185
rect 574 189 580 190
rect 574 185 575 189
rect 579 185 580 189
rect 574 184 580 185
rect 654 189 660 190
rect 654 185 655 189
rect 659 185 660 189
rect 654 184 660 185
rect 726 189 732 190
rect 726 185 727 189
rect 731 185 732 189
rect 726 184 732 185
rect 790 189 796 190
rect 790 185 791 189
rect 795 185 796 189
rect 790 184 796 185
rect 846 189 852 190
rect 846 185 847 189
rect 851 185 852 189
rect 846 184 852 185
rect 902 189 908 190
rect 902 185 903 189
rect 907 185 908 189
rect 902 184 908 185
rect 958 189 964 190
rect 958 185 959 189
rect 963 185 964 189
rect 958 184 964 185
rect 1022 189 1028 190
rect 1022 185 1023 189
rect 1027 185 1028 189
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1446 193 1452 194
rect 1446 189 1447 193
rect 1451 189 1452 193
rect 1446 188 1452 189
rect 1494 193 1500 194
rect 1494 189 1495 193
rect 1499 189 1500 193
rect 1494 188 1500 189
rect 1550 193 1556 194
rect 1550 189 1551 193
rect 1555 189 1556 193
rect 1550 188 1556 189
rect 1606 193 1612 194
rect 1606 189 1607 193
rect 1611 189 1612 193
rect 1606 188 1612 189
rect 1670 193 1676 194
rect 1670 189 1671 193
rect 1675 189 1676 193
rect 1670 188 1676 189
rect 1734 193 1740 194
rect 1734 189 1735 193
rect 1739 189 1740 193
rect 1734 188 1740 189
rect 1806 193 1812 194
rect 1806 189 1807 193
rect 1811 189 1812 193
rect 1806 188 1812 189
rect 1886 193 1892 194
rect 1886 189 1887 193
rect 1891 189 1892 193
rect 1886 188 1892 189
rect 1974 193 1980 194
rect 1974 189 1975 193
rect 1979 189 1980 193
rect 1974 188 1980 189
rect 2070 193 2076 194
rect 2070 189 2071 193
rect 2075 189 2076 193
rect 2070 188 2076 189
rect 2166 193 2172 194
rect 2166 189 2167 193
rect 2171 189 2172 193
rect 2166 188 2172 189
rect 2270 193 2276 194
rect 2270 189 2271 193
rect 2275 189 2276 193
rect 2270 188 2276 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1022 184 1028 185
rect 1302 147 1308 148
rect 1302 143 1303 147
rect 1307 143 1308 147
rect 1302 142 1308 143
rect 1342 147 1348 148
rect 1342 143 1343 147
rect 1347 143 1348 147
rect 1342 142 1348 143
rect 1382 147 1388 148
rect 1382 143 1383 147
rect 1387 143 1388 147
rect 1382 142 1388 143
rect 1422 147 1428 148
rect 1422 143 1423 147
rect 1427 143 1428 147
rect 1422 142 1428 143
rect 1462 147 1468 148
rect 1462 143 1463 147
rect 1467 143 1468 147
rect 1462 142 1468 143
rect 1518 147 1524 148
rect 1518 143 1519 147
rect 1523 143 1524 147
rect 1518 142 1524 143
rect 1582 147 1588 148
rect 1582 143 1583 147
rect 1587 143 1588 147
rect 1582 142 1588 143
rect 1646 147 1652 148
rect 1646 143 1647 147
rect 1651 143 1652 147
rect 1646 142 1652 143
rect 1710 147 1716 148
rect 1710 143 1711 147
rect 1715 143 1716 147
rect 1710 142 1716 143
rect 1766 147 1772 148
rect 1766 143 1767 147
rect 1771 143 1772 147
rect 1766 142 1772 143
rect 1822 147 1828 148
rect 1822 143 1823 147
rect 1827 143 1828 147
rect 1822 142 1828 143
rect 1870 147 1876 148
rect 1870 143 1871 147
rect 1875 143 1876 147
rect 1870 142 1876 143
rect 1918 147 1924 148
rect 1918 143 1919 147
rect 1923 143 1924 147
rect 1918 142 1924 143
rect 1966 147 1972 148
rect 1966 143 1967 147
rect 1971 143 1972 147
rect 1966 142 1972 143
rect 2014 147 2020 148
rect 2014 143 2015 147
rect 2019 143 2020 147
rect 2014 142 2020 143
rect 2062 147 2068 148
rect 2062 143 2063 147
rect 2067 143 2068 147
rect 2062 142 2068 143
rect 2110 147 2116 148
rect 2110 143 2111 147
rect 2115 143 2116 147
rect 2110 142 2116 143
rect 2158 147 2164 148
rect 2158 143 2159 147
rect 2163 143 2164 147
rect 2158 142 2164 143
rect 2214 147 2220 148
rect 2214 143 2215 147
rect 2219 143 2220 147
rect 2214 142 2220 143
rect 2270 147 2276 148
rect 2270 143 2271 147
rect 2275 143 2276 147
rect 2270 142 2276 143
rect 2318 147 2324 148
rect 2318 143 2319 147
rect 2323 143 2324 147
rect 2318 142 2324 143
rect 2358 147 2364 148
rect 2358 143 2359 147
rect 2363 143 2364 147
rect 2358 142 2364 143
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 174 139 180 140
rect 174 135 175 139
rect 179 135 180 139
rect 174 134 180 135
rect 214 139 220 140
rect 214 135 215 139
rect 219 135 220 139
rect 214 134 220 135
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 294 139 300 140
rect 294 135 295 139
rect 299 135 300 139
rect 294 134 300 135
rect 334 139 340 140
rect 334 135 335 139
rect 339 135 340 139
rect 334 134 340 135
rect 374 139 380 140
rect 374 135 375 139
rect 379 135 380 139
rect 374 134 380 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 582 139 588 140
rect 582 135 583 139
rect 587 135 588 139
rect 582 134 588 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 678 139 684 140
rect 678 135 679 139
rect 683 135 684 139
rect 678 134 684 135
rect 726 139 732 140
rect 726 135 727 139
rect 731 135 732 139
rect 726 134 732 135
rect 766 139 772 140
rect 766 135 767 139
rect 771 135 772 139
rect 766 134 772 135
rect 806 139 812 140
rect 806 135 807 139
rect 811 135 812 139
rect 806 134 812 135
rect 846 139 852 140
rect 846 135 847 139
rect 851 135 852 139
rect 846 134 852 135
rect 886 139 892 140
rect 886 135 887 139
rect 891 135 892 139
rect 886 134 892 135
rect 926 139 932 140
rect 926 135 927 139
rect 931 135 932 139
rect 926 134 932 135
rect 974 139 980 140
rect 974 135 975 139
rect 979 135 980 139
rect 974 134 980 135
rect 1022 139 1028 140
rect 1022 135 1023 139
rect 1027 135 1028 139
rect 1022 134 1028 135
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1278 124 1284 125
rect 1278 120 1279 124
rect 1283 120 1284 124
rect 1278 119 1284 120
rect 2406 124 2412 125
rect 2406 120 2407 124
rect 2411 120 2412 124
rect 2406 119 2412 120
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 110 111 116 112
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1238 111 1244 112
rect 1278 107 1284 108
rect 1278 103 1279 107
rect 1283 103 1284 107
rect 1278 102 1284 103
rect 2406 107 2412 108
rect 2406 103 2407 107
rect 2411 103 2412 107
rect 2406 102 2412 103
rect 1302 100 1308 101
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1302 96 1303 100
rect 1307 96 1308 100
rect 1302 95 1308 96
rect 1342 100 1348 101
rect 1342 96 1343 100
rect 1347 96 1348 100
rect 1342 95 1348 96
rect 1382 100 1388 101
rect 1382 96 1383 100
rect 1387 96 1388 100
rect 1382 95 1388 96
rect 1422 100 1428 101
rect 1422 96 1423 100
rect 1427 96 1428 100
rect 1422 95 1428 96
rect 1462 100 1468 101
rect 1462 96 1463 100
rect 1467 96 1468 100
rect 1462 95 1468 96
rect 1518 100 1524 101
rect 1518 96 1519 100
rect 1523 96 1524 100
rect 1518 95 1524 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1646 100 1652 101
rect 1646 96 1647 100
rect 1651 96 1652 100
rect 1646 95 1652 96
rect 1710 100 1716 101
rect 1710 96 1711 100
rect 1715 96 1716 100
rect 1710 95 1716 96
rect 1766 100 1772 101
rect 1766 96 1767 100
rect 1771 96 1772 100
rect 1766 95 1772 96
rect 1822 100 1828 101
rect 1822 96 1823 100
rect 1827 96 1828 100
rect 1822 95 1828 96
rect 1870 100 1876 101
rect 1870 96 1871 100
rect 1875 96 1876 100
rect 1870 95 1876 96
rect 1918 100 1924 101
rect 1918 96 1919 100
rect 1923 96 1924 100
rect 1918 95 1924 96
rect 1966 100 1972 101
rect 1966 96 1967 100
rect 1971 96 1972 100
rect 1966 95 1972 96
rect 2014 100 2020 101
rect 2014 96 2015 100
rect 2019 96 2020 100
rect 2014 95 2020 96
rect 2062 100 2068 101
rect 2062 96 2063 100
rect 2067 96 2068 100
rect 2062 95 2068 96
rect 2110 100 2116 101
rect 2110 96 2111 100
rect 2115 96 2116 100
rect 2110 95 2116 96
rect 2158 100 2164 101
rect 2158 96 2159 100
rect 2163 96 2164 100
rect 2158 95 2164 96
rect 2214 100 2220 101
rect 2214 96 2215 100
rect 2219 96 2220 100
rect 2214 95 2220 96
rect 2270 100 2276 101
rect 2270 96 2271 100
rect 2275 96 2276 100
rect 2270 95 2276 96
rect 2318 100 2324 101
rect 2318 96 2319 100
rect 2323 96 2324 100
rect 2318 95 2324 96
rect 2358 100 2364 101
rect 2358 96 2359 100
rect 2363 96 2364 100
rect 2358 95 2364 96
rect 1238 94 1244 95
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 526 92 532 93
rect 526 88 527 92
rect 531 88 532 92
rect 526 87 532 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 678 92 684 93
rect 678 88 679 92
rect 683 88 684 92
rect 678 87 684 88
rect 726 92 732 93
rect 726 88 727 92
rect 731 88 732 92
rect 726 87 732 88
rect 766 92 772 93
rect 766 88 767 92
rect 771 88 772 92
rect 766 87 772 88
rect 806 92 812 93
rect 806 88 807 92
rect 811 88 812 92
rect 806 87 812 88
rect 846 92 852 93
rect 846 88 847 92
rect 851 88 852 92
rect 846 87 852 88
rect 886 92 892 93
rect 886 88 887 92
rect 891 88 892 92
rect 886 87 892 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 974 92 980 93
rect 974 88 975 92
rect 979 88 980 92
rect 974 87 980 88
rect 1022 92 1028 93
rect 1022 88 1023 92
rect 1027 88 1028 92
rect 1022 87 1028 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
<< m3c >>
rect 1535 2504 1539 2508
rect 1575 2504 1579 2508
rect 1615 2504 1619 2508
rect 1655 2504 1659 2508
rect 1695 2504 1699 2508
rect 1735 2504 1739 2508
rect 1775 2504 1779 2508
rect 1815 2504 1819 2508
rect 1855 2504 1859 2508
rect 1895 2504 1899 2508
rect 1935 2504 1939 2508
rect 1975 2504 1979 2508
rect 1279 2497 1283 2501
rect 2407 2497 2411 2501
rect 135 2483 139 2487
rect 175 2483 179 2487
rect 215 2483 219 2487
rect 255 2483 259 2487
rect 311 2483 315 2487
rect 391 2483 395 2487
rect 479 2483 483 2487
rect 567 2483 571 2487
rect 655 2483 659 2487
rect 743 2483 747 2487
rect 831 2483 835 2487
rect 927 2483 931 2487
rect 1279 2480 1283 2484
rect 2407 2480 2411 2484
rect 111 2460 115 2464
rect 1239 2460 1243 2464
rect 1535 2457 1539 2461
rect 1575 2457 1579 2461
rect 1615 2457 1619 2461
rect 1655 2457 1659 2461
rect 1695 2457 1699 2461
rect 1735 2457 1739 2461
rect 1775 2457 1779 2461
rect 1815 2457 1819 2461
rect 1855 2457 1859 2461
rect 1895 2457 1899 2461
rect 1935 2457 1939 2461
rect 1975 2457 1979 2461
rect 111 2443 115 2447
rect 1239 2443 1243 2447
rect 135 2436 139 2440
rect 175 2436 179 2440
rect 215 2436 219 2440
rect 255 2436 259 2440
rect 311 2436 315 2440
rect 391 2436 395 2440
rect 479 2436 483 2440
rect 567 2436 571 2440
rect 655 2436 659 2440
rect 743 2436 747 2440
rect 831 2436 835 2440
rect 927 2436 931 2440
rect 135 2424 139 2428
rect 183 2424 187 2428
rect 247 2424 251 2428
rect 319 2424 323 2428
rect 391 2424 395 2428
rect 471 2424 475 2428
rect 543 2424 547 2428
rect 615 2424 619 2428
rect 679 2424 683 2428
rect 735 2424 739 2428
rect 791 2424 795 2428
rect 839 2424 843 2428
rect 887 2424 891 2428
rect 935 2424 939 2428
rect 991 2424 995 2428
rect 1047 2424 1051 2428
rect 1359 2427 1363 2431
rect 1399 2427 1403 2431
rect 1455 2427 1459 2431
rect 1519 2427 1523 2431
rect 1599 2427 1603 2431
rect 1679 2427 1683 2431
rect 1759 2427 1763 2431
rect 1839 2427 1843 2431
rect 1919 2427 1923 2431
rect 1999 2427 2003 2431
rect 2079 2427 2083 2431
rect 2159 2427 2163 2431
rect 2247 2427 2251 2431
rect 2335 2427 2339 2431
rect 111 2417 115 2421
rect 1239 2417 1243 2421
rect 111 2400 115 2404
rect 1239 2400 1243 2404
rect 1279 2404 1283 2408
rect 2407 2404 2411 2408
rect 1279 2387 1283 2391
rect 2407 2387 2411 2391
rect 135 2377 139 2381
rect 183 2377 187 2381
rect 247 2377 251 2381
rect 319 2377 323 2381
rect 391 2377 395 2381
rect 471 2377 475 2381
rect 543 2377 547 2381
rect 615 2377 619 2381
rect 679 2377 683 2381
rect 735 2377 739 2381
rect 791 2377 795 2381
rect 839 2377 843 2381
rect 887 2377 891 2381
rect 935 2377 939 2381
rect 991 2377 995 2381
rect 1047 2377 1051 2381
rect 1359 2380 1363 2384
rect 1399 2380 1403 2384
rect 1455 2380 1459 2384
rect 1519 2380 1523 2384
rect 1599 2380 1603 2384
rect 1679 2380 1683 2384
rect 1759 2380 1763 2384
rect 1839 2380 1843 2384
rect 1919 2380 1923 2384
rect 1999 2380 2003 2384
rect 2079 2380 2083 2384
rect 2159 2380 2163 2384
rect 2247 2380 2251 2384
rect 2335 2380 2339 2384
rect 1359 2368 1363 2372
rect 1407 2368 1411 2372
rect 1471 2368 1475 2372
rect 1543 2368 1547 2372
rect 1615 2368 1619 2372
rect 1695 2368 1699 2372
rect 1775 2368 1779 2372
rect 1855 2368 1859 2372
rect 1927 2368 1931 2372
rect 1999 2368 2003 2372
rect 2071 2368 2075 2372
rect 2143 2368 2147 2372
rect 2223 2368 2227 2372
rect 2303 2368 2307 2372
rect 2359 2368 2363 2372
rect 1279 2361 1283 2365
rect 2407 2361 2411 2365
rect 1279 2344 1283 2348
rect 135 2339 139 2343
rect 175 2339 179 2343
rect 215 2339 219 2343
rect 271 2339 275 2343
rect 351 2339 355 2343
rect 431 2339 435 2343
rect 519 2339 523 2343
rect 599 2339 603 2343
rect 679 2339 683 2343
rect 751 2339 755 2343
rect 823 2339 827 2343
rect 887 2339 891 2343
rect 959 2339 963 2343
rect 2407 2344 2411 2348
rect 1031 2339 1035 2343
rect 1359 2321 1363 2325
rect 111 2316 115 2320
rect 1407 2321 1411 2325
rect 1471 2321 1475 2325
rect 1543 2321 1547 2325
rect 1615 2321 1619 2325
rect 1695 2321 1699 2325
rect 1775 2321 1779 2325
rect 1855 2321 1859 2325
rect 1927 2321 1931 2325
rect 1999 2321 2003 2325
rect 2071 2321 2075 2325
rect 2143 2321 2147 2325
rect 2223 2321 2227 2325
rect 2303 2321 2307 2325
rect 2359 2321 2363 2325
rect 1239 2316 1243 2320
rect 111 2299 115 2303
rect 1239 2299 1243 2303
rect 135 2292 139 2296
rect 175 2292 179 2296
rect 215 2292 219 2296
rect 271 2292 275 2296
rect 351 2292 355 2296
rect 431 2292 435 2296
rect 519 2292 523 2296
rect 599 2292 603 2296
rect 679 2292 683 2296
rect 751 2292 755 2296
rect 823 2292 827 2296
rect 887 2292 891 2296
rect 959 2292 963 2296
rect 1031 2292 1035 2296
rect 1503 2287 1507 2291
rect 1543 2287 1547 2291
rect 1583 2287 1587 2291
rect 1623 2287 1627 2291
rect 1663 2287 1667 2291
rect 1703 2287 1707 2291
rect 1759 2287 1763 2291
rect 1823 2287 1827 2291
rect 1895 2287 1899 2291
rect 1967 2287 1971 2291
rect 2047 2287 2051 2291
rect 2127 2287 2131 2291
rect 2207 2287 2211 2291
rect 2295 2287 2299 2291
rect 2359 2287 2363 2291
rect 135 2276 139 2280
rect 175 2276 179 2280
rect 231 2276 235 2280
rect 303 2276 307 2280
rect 375 2276 379 2280
rect 455 2276 459 2280
rect 535 2276 539 2280
rect 615 2276 619 2280
rect 687 2276 691 2280
rect 759 2276 763 2280
rect 831 2276 835 2280
rect 911 2276 915 2280
rect 991 2276 995 2280
rect 111 2269 115 2273
rect 1239 2269 1243 2273
rect 1279 2264 1283 2268
rect 2407 2264 2411 2268
rect 111 2252 115 2256
rect 1239 2252 1243 2256
rect 1279 2247 1283 2251
rect 2407 2247 2411 2251
rect 1503 2240 1507 2244
rect 1543 2240 1547 2244
rect 1583 2240 1587 2244
rect 1623 2240 1627 2244
rect 1663 2240 1667 2244
rect 1703 2240 1707 2244
rect 1759 2240 1763 2244
rect 1823 2240 1827 2244
rect 1895 2240 1899 2244
rect 1967 2240 1971 2244
rect 2047 2240 2051 2244
rect 2127 2240 2131 2244
rect 2207 2240 2211 2244
rect 2295 2240 2299 2244
rect 2359 2240 2363 2244
rect 135 2229 139 2233
rect 175 2229 179 2233
rect 231 2229 235 2233
rect 303 2229 307 2233
rect 375 2229 379 2233
rect 455 2229 459 2233
rect 535 2229 539 2233
rect 615 2229 619 2233
rect 687 2229 691 2233
rect 759 2229 763 2233
rect 831 2229 835 2233
rect 911 2229 915 2233
rect 991 2229 995 2233
rect 1303 2220 1307 2224
rect 1343 2220 1347 2224
rect 1383 2220 1387 2224
rect 1431 2220 1435 2224
rect 1495 2220 1499 2224
rect 1567 2220 1571 2224
rect 1639 2220 1643 2224
rect 1711 2220 1715 2224
rect 1783 2220 1787 2224
rect 1855 2220 1859 2224
rect 1935 2220 1939 2224
rect 2015 2220 2019 2224
rect 2095 2220 2099 2224
rect 2183 2220 2187 2224
rect 2279 2220 2283 2224
rect 2359 2220 2363 2224
rect 1279 2213 1283 2217
rect 2407 2213 2411 2217
rect 247 2199 251 2203
rect 287 2199 291 2203
rect 327 2199 331 2203
rect 375 2199 379 2203
rect 431 2199 435 2203
rect 495 2199 499 2203
rect 551 2199 555 2203
rect 607 2199 611 2203
rect 663 2199 667 2203
rect 719 2199 723 2203
rect 783 2199 787 2203
rect 847 2199 851 2203
rect 911 2199 915 2203
rect 1279 2196 1283 2200
rect 2407 2196 2411 2200
rect 111 2176 115 2180
rect 1239 2176 1243 2180
rect 1303 2173 1307 2177
rect 1343 2173 1347 2177
rect 1383 2173 1387 2177
rect 1431 2173 1435 2177
rect 1495 2173 1499 2177
rect 1567 2173 1571 2177
rect 1639 2173 1643 2177
rect 1711 2173 1715 2177
rect 1783 2173 1787 2177
rect 1855 2173 1859 2177
rect 1935 2173 1939 2177
rect 2015 2173 2019 2177
rect 2095 2173 2099 2177
rect 2183 2173 2187 2177
rect 2279 2173 2283 2177
rect 2359 2173 2363 2177
rect 111 2159 115 2163
rect 1239 2159 1243 2163
rect 247 2152 251 2156
rect 287 2152 291 2156
rect 327 2152 331 2156
rect 375 2152 379 2156
rect 431 2152 435 2156
rect 495 2152 499 2156
rect 551 2152 555 2156
rect 607 2152 611 2156
rect 663 2152 667 2156
rect 719 2152 723 2156
rect 783 2152 787 2156
rect 847 2152 851 2156
rect 911 2152 915 2156
rect 1303 2143 1307 2147
rect 1351 2143 1355 2147
rect 1439 2143 1443 2147
rect 1535 2143 1539 2147
rect 1631 2143 1635 2147
rect 1727 2143 1731 2147
rect 1815 2143 1819 2147
rect 1895 2143 1899 2147
rect 1975 2143 1979 2147
rect 2047 2143 2051 2147
rect 2111 2143 2115 2147
rect 2175 2143 2179 2147
rect 2239 2143 2243 2147
rect 2311 2143 2315 2147
rect 2359 2143 2363 2147
rect 383 2132 387 2136
rect 423 2132 427 2136
rect 463 2132 467 2136
rect 503 2132 507 2136
rect 551 2132 555 2136
rect 607 2132 611 2136
rect 663 2132 667 2136
rect 727 2132 731 2136
rect 791 2132 795 2136
rect 855 2132 859 2136
rect 911 2132 915 2136
rect 967 2132 971 2136
rect 1023 2132 1027 2136
rect 1079 2132 1083 2136
rect 1143 2132 1147 2136
rect 111 2125 115 2129
rect 1239 2125 1243 2129
rect 1279 2120 1283 2124
rect 2407 2120 2411 2124
rect 111 2108 115 2112
rect 1239 2108 1243 2112
rect 1279 2103 1283 2107
rect 2407 2103 2411 2107
rect 1303 2096 1307 2100
rect 1351 2096 1355 2100
rect 1439 2096 1443 2100
rect 1535 2096 1539 2100
rect 1631 2096 1635 2100
rect 1727 2096 1731 2100
rect 1815 2096 1819 2100
rect 1895 2096 1899 2100
rect 1975 2096 1979 2100
rect 2047 2096 2051 2100
rect 2111 2096 2115 2100
rect 2175 2096 2179 2100
rect 2239 2096 2243 2100
rect 2311 2096 2315 2100
rect 2359 2096 2363 2100
rect 383 2085 387 2089
rect 423 2085 427 2089
rect 463 2085 467 2089
rect 503 2085 507 2089
rect 551 2085 555 2089
rect 607 2085 611 2089
rect 663 2085 667 2089
rect 727 2085 731 2089
rect 791 2085 795 2089
rect 855 2085 859 2089
rect 911 2085 915 2089
rect 967 2085 971 2089
rect 1023 2085 1027 2089
rect 1079 2085 1083 2089
rect 1143 2085 1147 2089
rect 1303 2080 1307 2084
rect 1343 2080 1347 2084
rect 1399 2080 1403 2084
rect 1479 2080 1483 2084
rect 1567 2080 1571 2084
rect 1663 2080 1667 2084
rect 1759 2080 1763 2084
rect 1847 2080 1851 2084
rect 1935 2080 1939 2084
rect 2015 2080 2019 2084
rect 2095 2080 2099 2084
rect 2167 2080 2171 2084
rect 2239 2080 2243 2084
rect 2311 2080 2315 2084
rect 2359 2080 2363 2084
rect 1279 2073 1283 2077
rect 2407 2073 2411 2077
rect 383 2055 387 2059
rect 423 2055 427 2059
rect 463 2055 467 2059
rect 503 2055 507 2059
rect 543 2055 547 2059
rect 583 2055 587 2059
rect 631 2055 635 2059
rect 687 2055 691 2059
rect 743 2055 747 2059
rect 799 2055 803 2059
rect 847 2055 851 2059
rect 903 2055 907 2059
rect 959 2055 963 2059
rect 1015 2055 1019 2059
rect 1071 2055 1075 2059
rect 1279 2056 1283 2060
rect 2407 2056 2411 2060
rect 111 2032 115 2036
rect 1239 2032 1243 2036
rect 1303 2033 1307 2037
rect 1343 2033 1347 2037
rect 1399 2033 1403 2037
rect 1479 2033 1483 2037
rect 1567 2033 1571 2037
rect 1663 2033 1667 2037
rect 1759 2033 1763 2037
rect 1847 2033 1851 2037
rect 1935 2033 1939 2037
rect 2015 2033 2019 2037
rect 2095 2033 2099 2037
rect 2167 2033 2171 2037
rect 2239 2033 2243 2037
rect 2311 2033 2315 2037
rect 2359 2033 2363 2037
rect 111 2015 115 2019
rect 1239 2015 1243 2019
rect 383 2008 387 2012
rect 423 2008 427 2012
rect 463 2008 467 2012
rect 503 2008 507 2012
rect 543 2008 547 2012
rect 583 2008 587 2012
rect 631 2008 635 2012
rect 687 2008 691 2012
rect 743 2008 747 2012
rect 799 2008 803 2012
rect 847 2008 851 2012
rect 903 2008 907 2012
rect 959 2008 963 2012
rect 1015 2008 1019 2012
rect 1071 2008 1075 2012
rect 1303 1995 1307 1999
rect 1351 1995 1355 1999
rect 1423 1995 1427 1999
rect 1495 1995 1499 1999
rect 1575 1995 1579 1999
rect 1663 1995 1667 1999
rect 1751 1995 1755 1999
rect 1839 1995 1843 1999
rect 1919 1995 1923 1999
rect 1999 1995 2003 1999
rect 2071 1995 2075 1999
rect 2135 1995 2139 1999
rect 2191 1995 2195 1999
rect 2255 1995 2259 1999
rect 2319 1995 2323 1999
rect 2359 1995 2363 1999
rect 367 1988 371 1992
rect 407 1988 411 1992
rect 455 1988 459 1992
rect 511 1988 515 1992
rect 567 1988 571 1992
rect 631 1988 635 1992
rect 695 1988 699 1992
rect 759 1988 763 1992
rect 815 1988 819 1992
rect 871 1988 875 1992
rect 935 1988 939 1992
rect 999 1988 1003 1992
rect 1063 1988 1067 1992
rect 111 1981 115 1985
rect 1239 1981 1243 1985
rect 1279 1972 1283 1976
rect 2407 1972 2411 1976
rect 111 1964 115 1968
rect 1239 1964 1243 1968
rect 1279 1955 1283 1959
rect 2407 1955 2411 1959
rect 1303 1948 1307 1952
rect 1351 1948 1355 1952
rect 1423 1948 1427 1952
rect 1495 1948 1499 1952
rect 1575 1948 1579 1952
rect 1663 1948 1667 1952
rect 1751 1948 1755 1952
rect 1839 1948 1843 1952
rect 1919 1948 1923 1952
rect 1999 1948 2003 1952
rect 2071 1948 2075 1952
rect 2135 1948 2139 1952
rect 2191 1948 2195 1952
rect 2255 1948 2259 1952
rect 2319 1948 2323 1952
rect 2359 1948 2363 1952
rect 367 1941 371 1945
rect 407 1941 411 1945
rect 455 1941 459 1945
rect 511 1941 515 1945
rect 567 1941 571 1945
rect 631 1941 635 1945
rect 695 1941 699 1945
rect 759 1941 763 1945
rect 815 1941 819 1945
rect 871 1941 875 1945
rect 935 1941 939 1945
rect 999 1941 1003 1945
rect 1063 1941 1067 1945
rect 1303 1936 1307 1940
rect 1359 1936 1363 1940
rect 1447 1936 1451 1940
rect 1535 1936 1539 1940
rect 1623 1936 1627 1940
rect 1711 1936 1715 1940
rect 1791 1936 1795 1940
rect 1863 1936 1867 1940
rect 1935 1936 1939 1940
rect 2007 1936 2011 1940
rect 2079 1936 2083 1940
rect 2151 1936 2155 1940
rect 2223 1936 2227 1940
rect 2303 1936 2307 1940
rect 2359 1936 2363 1940
rect 1279 1929 1283 1933
rect 2407 1929 2411 1933
rect 1279 1912 1283 1916
rect 175 1907 179 1911
rect 215 1907 219 1911
rect 263 1907 267 1911
rect 319 1907 323 1911
rect 391 1907 395 1911
rect 471 1907 475 1911
rect 551 1907 555 1911
rect 639 1907 643 1911
rect 719 1907 723 1911
rect 799 1907 803 1911
rect 879 1907 883 1911
rect 959 1907 963 1911
rect 1039 1907 1043 1911
rect 2407 1912 2411 1916
rect 1119 1907 1123 1911
rect 1303 1889 1307 1893
rect 111 1884 115 1888
rect 1359 1889 1363 1893
rect 1447 1889 1451 1893
rect 1535 1889 1539 1893
rect 1623 1889 1627 1893
rect 1711 1889 1715 1893
rect 1791 1889 1795 1893
rect 1863 1889 1867 1893
rect 1935 1889 1939 1893
rect 2007 1889 2011 1893
rect 2079 1889 2083 1893
rect 2151 1889 2155 1893
rect 2223 1889 2227 1893
rect 2303 1889 2307 1893
rect 2359 1889 2363 1893
rect 1239 1884 1243 1888
rect 111 1867 115 1871
rect 1239 1867 1243 1871
rect 175 1860 179 1864
rect 215 1860 219 1864
rect 263 1860 267 1864
rect 319 1860 323 1864
rect 391 1860 395 1864
rect 471 1860 475 1864
rect 551 1860 555 1864
rect 639 1860 643 1864
rect 719 1860 723 1864
rect 799 1860 803 1864
rect 879 1860 883 1864
rect 959 1860 963 1864
rect 1039 1860 1043 1864
rect 1119 1860 1123 1864
rect 1311 1859 1315 1863
rect 1359 1859 1363 1863
rect 1415 1859 1419 1863
rect 1479 1859 1483 1863
rect 1543 1859 1547 1863
rect 1615 1859 1619 1863
rect 1687 1859 1691 1863
rect 1767 1859 1771 1863
rect 1863 1859 1867 1863
rect 1975 1859 1979 1863
rect 2095 1859 2099 1863
rect 2223 1859 2227 1863
rect 2359 1859 2363 1863
rect 135 1840 139 1844
rect 175 1840 179 1844
rect 215 1840 219 1844
rect 271 1840 275 1844
rect 351 1840 355 1844
rect 439 1840 443 1844
rect 535 1840 539 1844
rect 631 1840 635 1844
rect 727 1840 731 1844
rect 823 1840 827 1844
rect 911 1840 915 1844
rect 991 1840 995 1844
rect 1063 1840 1067 1844
rect 1135 1840 1139 1844
rect 1191 1840 1195 1844
rect 111 1833 115 1837
rect 1239 1833 1243 1837
rect 1279 1836 1283 1840
rect 2407 1836 2411 1840
rect 111 1816 115 1820
rect 1239 1816 1243 1820
rect 1279 1819 1283 1823
rect 2407 1819 2411 1823
rect 1311 1812 1315 1816
rect 1359 1812 1363 1816
rect 1415 1812 1419 1816
rect 1479 1812 1483 1816
rect 1543 1812 1547 1816
rect 1615 1812 1619 1816
rect 1687 1812 1691 1816
rect 1767 1812 1771 1816
rect 1863 1812 1867 1816
rect 1975 1812 1979 1816
rect 2095 1812 2099 1816
rect 2223 1812 2227 1816
rect 2359 1812 2363 1816
rect 135 1793 139 1797
rect 175 1793 179 1797
rect 215 1793 219 1797
rect 271 1793 275 1797
rect 351 1793 355 1797
rect 439 1793 443 1797
rect 535 1793 539 1797
rect 631 1793 635 1797
rect 727 1793 731 1797
rect 823 1793 827 1797
rect 911 1793 915 1797
rect 991 1793 995 1797
rect 1063 1793 1067 1797
rect 1135 1793 1139 1797
rect 1191 1793 1195 1797
rect 1407 1796 1411 1800
rect 1471 1796 1475 1800
rect 1535 1796 1539 1800
rect 1599 1796 1603 1800
rect 1663 1796 1667 1800
rect 1727 1796 1731 1800
rect 1783 1796 1787 1800
rect 1839 1796 1843 1800
rect 1895 1796 1899 1800
rect 1959 1796 1963 1800
rect 1279 1789 1283 1793
rect 2407 1789 2411 1793
rect 1279 1772 1283 1776
rect 2407 1772 2411 1776
rect 135 1763 139 1767
rect 175 1763 179 1767
rect 215 1763 219 1767
rect 287 1763 291 1767
rect 375 1763 379 1767
rect 471 1763 475 1767
rect 567 1763 571 1767
rect 663 1763 667 1767
rect 751 1763 755 1767
rect 831 1763 835 1767
rect 903 1763 907 1767
rect 967 1763 971 1767
rect 1031 1763 1035 1767
rect 1087 1763 1091 1767
rect 1151 1763 1155 1767
rect 1191 1763 1195 1767
rect 1407 1749 1411 1753
rect 1471 1749 1475 1753
rect 1535 1749 1539 1753
rect 1599 1749 1603 1753
rect 1663 1749 1667 1753
rect 1727 1749 1731 1753
rect 1783 1749 1787 1753
rect 1839 1749 1843 1753
rect 1895 1749 1899 1753
rect 1959 1749 1963 1753
rect 111 1740 115 1744
rect 1239 1740 1243 1744
rect 111 1723 115 1727
rect 1239 1723 1243 1727
rect 135 1716 139 1720
rect 175 1716 179 1720
rect 215 1716 219 1720
rect 287 1716 291 1720
rect 375 1716 379 1720
rect 471 1716 475 1720
rect 567 1716 571 1720
rect 663 1716 667 1720
rect 751 1716 755 1720
rect 831 1716 835 1720
rect 903 1716 907 1720
rect 967 1716 971 1720
rect 1031 1716 1035 1720
rect 1087 1716 1091 1720
rect 1151 1716 1155 1720
rect 1191 1716 1195 1720
rect 1303 1719 1307 1723
rect 1351 1719 1355 1723
rect 1423 1719 1427 1723
rect 1503 1719 1507 1723
rect 1583 1719 1587 1723
rect 1663 1719 1667 1723
rect 1735 1719 1739 1723
rect 1807 1719 1811 1723
rect 1871 1719 1875 1723
rect 1935 1719 1939 1723
rect 1999 1719 2003 1723
rect 2063 1719 2067 1723
rect 135 1700 139 1704
rect 175 1700 179 1704
rect 239 1700 243 1704
rect 319 1700 323 1704
rect 415 1700 419 1704
rect 511 1700 515 1704
rect 615 1700 619 1704
rect 711 1700 715 1704
rect 799 1700 803 1704
rect 879 1700 883 1704
rect 951 1700 955 1704
rect 1015 1700 1019 1704
rect 1087 1700 1091 1704
rect 1159 1700 1163 1704
rect 111 1693 115 1697
rect 1239 1693 1243 1697
rect 1279 1696 1283 1700
rect 2407 1696 2411 1700
rect 111 1676 115 1680
rect 1239 1676 1243 1680
rect 1279 1679 1283 1683
rect 2407 1679 2411 1683
rect 1303 1672 1307 1676
rect 1351 1672 1355 1676
rect 1423 1672 1427 1676
rect 1503 1672 1507 1676
rect 1583 1672 1587 1676
rect 1663 1672 1667 1676
rect 1735 1672 1739 1676
rect 1807 1672 1811 1676
rect 1871 1672 1875 1676
rect 1935 1672 1939 1676
rect 1999 1672 2003 1676
rect 2063 1672 2067 1676
rect 1303 1660 1307 1664
rect 1359 1660 1363 1664
rect 1447 1660 1451 1664
rect 1543 1660 1547 1664
rect 1639 1660 1643 1664
rect 1727 1660 1731 1664
rect 1815 1660 1819 1664
rect 1895 1660 1899 1664
rect 1967 1660 1971 1664
rect 2031 1660 2035 1664
rect 2095 1660 2099 1664
rect 2159 1660 2163 1664
rect 2223 1660 2227 1664
rect 135 1653 139 1657
rect 175 1653 179 1657
rect 239 1653 243 1657
rect 319 1653 323 1657
rect 415 1653 419 1657
rect 511 1653 515 1657
rect 615 1653 619 1657
rect 711 1653 715 1657
rect 799 1653 803 1657
rect 879 1653 883 1657
rect 951 1653 955 1657
rect 1015 1653 1019 1657
rect 1087 1653 1091 1657
rect 1159 1653 1163 1657
rect 1279 1653 1283 1657
rect 2407 1653 2411 1657
rect 1279 1636 1283 1640
rect 2407 1636 2411 1640
rect 271 1619 275 1623
rect 311 1619 315 1623
rect 359 1619 363 1623
rect 415 1619 419 1623
rect 471 1619 475 1623
rect 535 1619 539 1623
rect 599 1619 603 1623
rect 663 1619 667 1623
rect 719 1619 723 1623
rect 775 1619 779 1623
rect 831 1619 835 1623
rect 887 1619 891 1623
rect 943 1619 947 1623
rect 999 1619 1003 1623
rect 1303 1613 1307 1617
rect 1359 1613 1363 1617
rect 1447 1613 1451 1617
rect 1543 1613 1547 1617
rect 1639 1613 1643 1617
rect 1727 1613 1731 1617
rect 1815 1613 1819 1617
rect 1895 1613 1899 1617
rect 1967 1613 1971 1617
rect 2031 1613 2035 1617
rect 2095 1613 2099 1617
rect 2159 1613 2163 1617
rect 2223 1613 2227 1617
rect 111 1596 115 1600
rect 1239 1596 1243 1600
rect 111 1579 115 1583
rect 1239 1579 1243 1583
rect 1327 1583 1331 1587
rect 1399 1583 1403 1587
rect 1479 1583 1483 1587
rect 1567 1583 1571 1587
rect 1655 1583 1659 1587
rect 1743 1583 1747 1587
rect 1831 1583 1835 1587
rect 1911 1583 1915 1587
rect 1983 1583 1987 1587
rect 2047 1583 2051 1587
rect 2111 1583 2115 1587
rect 2167 1583 2171 1587
rect 2215 1583 2219 1587
rect 2271 1583 2275 1587
rect 2319 1583 2323 1587
rect 2359 1583 2363 1587
rect 271 1572 275 1576
rect 311 1572 315 1576
rect 359 1572 363 1576
rect 415 1572 419 1576
rect 471 1572 475 1576
rect 535 1572 539 1576
rect 599 1572 603 1576
rect 663 1572 667 1576
rect 719 1572 723 1576
rect 775 1572 779 1576
rect 831 1572 835 1576
rect 887 1572 891 1576
rect 943 1572 947 1576
rect 999 1572 1003 1576
rect 1279 1560 1283 1564
rect 2407 1560 2411 1564
rect 327 1552 331 1556
rect 367 1552 371 1556
rect 407 1552 411 1556
rect 447 1552 451 1556
rect 487 1552 491 1556
rect 527 1552 531 1556
rect 567 1552 571 1556
rect 607 1552 611 1556
rect 647 1552 651 1556
rect 687 1552 691 1556
rect 727 1552 731 1556
rect 767 1552 771 1556
rect 807 1552 811 1556
rect 847 1552 851 1556
rect 887 1552 891 1556
rect 927 1552 931 1556
rect 111 1545 115 1549
rect 1239 1545 1243 1549
rect 1279 1543 1283 1547
rect 2407 1543 2411 1547
rect 1327 1536 1331 1540
rect 1399 1536 1403 1540
rect 1479 1536 1483 1540
rect 1567 1536 1571 1540
rect 1655 1536 1659 1540
rect 1743 1536 1747 1540
rect 1831 1536 1835 1540
rect 1911 1536 1915 1540
rect 1983 1536 1987 1540
rect 2047 1536 2051 1540
rect 2111 1536 2115 1540
rect 2167 1536 2171 1540
rect 2215 1536 2219 1540
rect 2271 1536 2275 1540
rect 2319 1536 2323 1540
rect 2359 1536 2363 1540
rect 111 1528 115 1532
rect 1239 1528 1243 1532
rect 1335 1520 1339 1524
rect 1415 1520 1419 1524
rect 1503 1520 1507 1524
rect 1615 1520 1619 1524
rect 1743 1520 1747 1524
rect 1887 1520 1891 1524
rect 2047 1520 2051 1524
rect 2215 1520 2219 1524
rect 2359 1520 2363 1524
rect 1279 1513 1283 1517
rect 2407 1513 2411 1517
rect 327 1505 331 1509
rect 367 1505 371 1509
rect 407 1505 411 1509
rect 447 1505 451 1509
rect 487 1505 491 1509
rect 527 1505 531 1509
rect 567 1505 571 1509
rect 607 1505 611 1509
rect 647 1505 651 1509
rect 687 1505 691 1509
rect 727 1505 731 1509
rect 767 1505 771 1509
rect 807 1505 811 1509
rect 847 1505 851 1509
rect 887 1505 891 1509
rect 927 1505 931 1509
rect 1279 1496 1283 1500
rect 2407 1496 2411 1500
rect 1335 1473 1339 1477
rect 1415 1473 1419 1477
rect 1503 1473 1507 1477
rect 1615 1473 1619 1477
rect 1743 1473 1747 1477
rect 1887 1473 1891 1477
rect 2047 1473 2051 1477
rect 2215 1473 2219 1477
rect 2359 1473 2363 1477
rect 1375 1443 1379 1447
rect 1463 1443 1467 1447
rect 1551 1443 1555 1447
rect 1639 1443 1643 1447
rect 1727 1443 1731 1447
rect 1807 1443 1811 1447
rect 1879 1443 1883 1447
rect 1943 1443 1947 1447
rect 1999 1443 2003 1447
rect 2047 1443 2051 1447
rect 2095 1443 2099 1447
rect 2143 1443 2147 1447
rect 2191 1443 2195 1447
rect 2239 1443 2243 1447
rect 2279 1443 2283 1447
rect 2319 1443 2323 1447
rect 2359 1443 2363 1447
rect 143 1435 147 1439
rect 183 1435 187 1439
rect 223 1435 227 1439
rect 263 1435 267 1439
rect 319 1435 323 1439
rect 391 1435 395 1439
rect 471 1435 475 1439
rect 559 1435 563 1439
rect 647 1435 651 1439
rect 727 1435 731 1439
rect 807 1435 811 1439
rect 879 1435 883 1439
rect 943 1435 947 1439
rect 999 1435 1003 1439
rect 1047 1435 1051 1439
rect 1103 1435 1107 1439
rect 1151 1435 1155 1439
rect 1191 1435 1195 1439
rect 1279 1420 1283 1424
rect 2407 1420 2411 1424
rect 111 1412 115 1416
rect 1239 1412 1243 1416
rect 1279 1403 1283 1407
rect 2407 1403 2411 1407
rect 111 1395 115 1399
rect 1239 1395 1243 1399
rect 1375 1396 1379 1400
rect 1463 1396 1467 1400
rect 1551 1396 1555 1400
rect 1639 1396 1643 1400
rect 1727 1396 1731 1400
rect 1807 1396 1811 1400
rect 1879 1396 1883 1400
rect 1943 1396 1947 1400
rect 1999 1396 2003 1400
rect 2047 1396 2051 1400
rect 2095 1396 2099 1400
rect 2143 1396 2147 1400
rect 2191 1396 2195 1400
rect 2239 1396 2243 1400
rect 2279 1396 2283 1400
rect 2319 1396 2323 1400
rect 2359 1396 2363 1400
rect 143 1388 147 1392
rect 183 1388 187 1392
rect 223 1388 227 1392
rect 263 1388 267 1392
rect 319 1388 323 1392
rect 391 1388 395 1392
rect 471 1388 475 1392
rect 559 1388 563 1392
rect 647 1388 651 1392
rect 727 1388 731 1392
rect 807 1388 811 1392
rect 879 1388 883 1392
rect 943 1388 947 1392
rect 999 1388 1003 1392
rect 1047 1388 1051 1392
rect 1103 1388 1107 1392
rect 1151 1388 1155 1392
rect 1191 1388 1195 1392
rect 167 1376 171 1380
rect 207 1376 211 1380
rect 247 1376 251 1380
rect 303 1376 307 1380
rect 367 1376 371 1380
rect 439 1376 443 1380
rect 519 1376 523 1380
rect 599 1376 603 1380
rect 679 1376 683 1380
rect 751 1376 755 1380
rect 823 1376 827 1380
rect 887 1376 891 1380
rect 951 1376 955 1380
rect 1015 1376 1019 1380
rect 1079 1376 1083 1380
rect 1143 1376 1147 1380
rect 1191 1376 1195 1380
rect 1303 1376 1307 1380
rect 1343 1376 1347 1380
rect 1399 1376 1403 1380
rect 1463 1376 1467 1380
rect 1535 1376 1539 1380
rect 1607 1376 1611 1380
rect 1687 1376 1691 1380
rect 1767 1376 1771 1380
rect 1847 1376 1851 1380
rect 1935 1376 1939 1380
rect 2023 1376 2027 1380
rect 2111 1376 2115 1380
rect 2199 1376 2203 1380
rect 2287 1376 2291 1380
rect 2359 1376 2363 1380
rect 111 1369 115 1373
rect 1239 1369 1243 1373
rect 1279 1369 1283 1373
rect 2407 1369 2411 1373
rect 111 1352 115 1356
rect 1239 1352 1243 1356
rect 1279 1352 1283 1356
rect 2407 1352 2411 1356
rect 167 1329 171 1333
rect 207 1329 211 1333
rect 247 1329 251 1333
rect 303 1329 307 1333
rect 367 1329 371 1333
rect 439 1329 443 1333
rect 519 1329 523 1333
rect 599 1329 603 1333
rect 679 1329 683 1333
rect 751 1329 755 1333
rect 823 1329 827 1333
rect 887 1329 891 1333
rect 951 1329 955 1333
rect 1015 1329 1019 1333
rect 1079 1329 1083 1333
rect 1143 1329 1147 1333
rect 1191 1329 1195 1333
rect 1303 1329 1307 1333
rect 1343 1329 1347 1333
rect 1399 1329 1403 1333
rect 1463 1329 1467 1333
rect 1535 1329 1539 1333
rect 1607 1329 1611 1333
rect 1687 1329 1691 1333
rect 1767 1329 1771 1333
rect 1847 1329 1851 1333
rect 1935 1329 1939 1333
rect 2023 1329 2027 1333
rect 2111 1329 2115 1333
rect 2199 1329 2203 1333
rect 2287 1329 2291 1333
rect 2359 1329 2363 1333
rect 183 1295 187 1299
rect 231 1295 235 1299
rect 287 1295 291 1299
rect 351 1295 355 1299
rect 423 1295 427 1299
rect 495 1295 499 1299
rect 567 1295 571 1299
rect 639 1295 643 1299
rect 703 1295 707 1299
rect 767 1295 771 1299
rect 823 1295 827 1299
rect 879 1295 883 1299
rect 935 1295 939 1299
rect 999 1295 1003 1299
rect 1303 1299 1307 1303
rect 1343 1299 1347 1303
rect 1383 1299 1387 1303
rect 1423 1299 1427 1303
rect 1463 1299 1467 1303
rect 1503 1299 1507 1303
rect 1543 1299 1547 1303
rect 1583 1299 1587 1303
rect 1623 1299 1627 1303
rect 1679 1299 1683 1303
rect 1735 1299 1739 1303
rect 1791 1299 1795 1303
rect 1847 1299 1851 1303
rect 1903 1299 1907 1303
rect 1967 1299 1971 1303
rect 2039 1299 2043 1303
rect 2119 1299 2123 1303
rect 2199 1299 2203 1303
rect 2287 1299 2291 1303
rect 2359 1299 2363 1303
rect 111 1272 115 1276
rect 1239 1272 1243 1276
rect 1279 1276 1283 1280
rect 2407 1276 2411 1280
rect 111 1255 115 1259
rect 1239 1255 1243 1259
rect 1279 1259 1283 1263
rect 2407 1259 2411 1263
rect 183 1248 187 1252
rect 231 1248 235 1252
rect 287 1248 291 1252
rect 351 1248 355 1252
rect 423 1248 427 1252
rect 495 1248 499 1252
rect 567 1248 571 1252
rect 639 1248 643 1252
rect 703 1248 707 1252
rect 767 1248 771 1252
rect 823 1248 827 1252
rect 879 1248 883 1252
rect 935 1248 939 1252
rect 999 1248 1003 1252
rect 1303 1252 1307 1256
rect 1343 1252 1347 1256
rect 1383 1252 1387 1256
rect 1423 1252 1427 1256
rect 1463 1252 1467 1256
rect 1503 1252 1507 1256
rect 1543 1252 1547 1256
rect 1583 1252 1587 1256
rect 1623 1252 1627 1256
rect 1679 1252 1683 1256
rect 1735 1252 1739 1256
rect 1791 1252 1795 1256
rect 1847 1252 1851 1256
rect 1903 1252 1907 1256
rect 1967 1252 1971 1256
rect 2039 1252 2043 1256
rect 2119 1252 2123 1256
rect 2199 1252 2203 1256
rect 2287 1252 2291 1256
rect 2359 1252 2363 1256
rect 135 1232 139 1236
rect 175 1232 179 1236
rect 231 1232 235 1236
rect 311 1232 315 1236
rect 399 1232 403 1236
rect 487 1232 491 1236
rect 575 1232 579 1236
rect 663 1232 667 1236
rect 743 1232 747 1236
rect 815 1232 819 1236
rect 879 1232 883 1236
rect 943 1232 947 1236
rect 1007 1232 1011 1236
rect 1071 1232 1075 1236
rect 1303 1232 1307 1236
rect 1375 1232 1379 1236
rect 1479 1232 1483 1236
rect 1583 1232 1587 1236
rect 1687 1232 1691 1236
rect 1791 1232 1795 1236
rect 1887 1232 1891 1236
rect 1983 1232 1987 1236
rect 2071 1232 2075 1236
rect 2151 1232 2155 1236
rect 2223 1232 2227 1236
rect 2303 1232 2307 1236
rect 2359 1232 2363 1236
rect 111 1225 115 1229
rect 1239 1225 1243 1229
rect 1279 1225 1283 1229
rect 2407 1225 2411 1229
rect 111 1208 115 1212
rect 1239 1208 1243 1212
rect 1279 1208 1283 1212
rect 2407 1208 2411 1212
rect 135 1185 139 1189
rect 175 1185 179 1189
rect 231 1185 235 1189
rect 311 1185 315 1189
rect 399 1185 403 1189
rect 487 1185 491 1189
rect 575 1185 579 1189
rect 663 1185 667 1189
rect 743 1185 747 1189
rect 815 1185 819 1189
rect 879 1185 883 1189
rect 943 1185 947 1189
rect 1007 1185 1011 1189
rect 1071 1185 1075 1189
rect 1303 1185 1307 1189
rect 1375 1185 1379 1189
rect 1479 1185 1483 1189
rect 1583 1185 1587 1189
rect 1687 1185 1691 1189
rect 1791 1185 1795 1189
rect 1887 1185 1891 1189
rect 1983 1185 1987 1189
rect 2071 1185 2075 1189
rect 2151 1185 2155 1189
rect 2223 1185 2227 1189
rect 2303 1185 2307 1189
rect 2359 1185 2363 1189
rect 135 1155 139 1159
rect 175 1155 179 1159
rect 239 1155 243 1159
rect 327 1155 331 1159
rect 431 1155 435 1159
rect 535 1155 539 1159
rect 639 1155 643 1159
rect 743 1155 747 1159
rect 839 1155 843 1159
rect 919 1155 923 1159
rect 999 1155 1003 1159
rect 1071 1155 1075 1159
rect 1143 1155 1147 1159
rect 1191 1155 1195 1159
rect 1303 1155 1307 1159
rect 1343 1155 1347 1159
rect 1407 1155 1411 1159
rect 1487 1155 1491 1159
rect 1583 1155 1587 1159
rect 1687 1155 1691 1159
rect 1799 1155 1803 1159
rect 1903 1155 1907 1159
rect 1999 1155 2003 1159
rect 2079 1155 2083 1159
rect 2159 1155 2163 1159
rect 2231 1155 2235 1159
rect 2303 1155 2307 1159
rect 2359 1155 2363 1159
rect 111 1132 115 1136
rect 1239 1132 1243 1136
rect 1279 1132 1283 1136
rect 2407 1132 2411 1136
rect 111 1115 115 1119
rect 1239 1115 1243 1119
rect 1279 1115 1283 1119
rect 2407 1115 2411 1119
rect 135 1108 139 1112
rect 175 1108 179 1112
rect 239 1108 243 1112
rect 327 1108 331 1112
rect 431 1108 435 1112
rect 535 1108 539 1112
rect 639 1108 643 1112
rect 743 1108 747 1112
rect 839 1108 843 1112
rect 919 1108 923 1112
rect 999 1108 1003 1112
rect 1071 1108 1075 1112
rect 1143 1108 1147 1112
rect 1191 1108 1195 1112
rect 1303 1108 1307 1112
rect 1343 1108 1347 1112
rect 1407 1108 1411 1112
rect 1487 1108 1491 1112
rect 1583 1108 1587 1112
rect 1687 1108 1691 1112
rect 1799 1108 1803 1112
rect 1903 1108 1907 1112
rect 1999 1108 2003 1112
rect 2079 1108 2083 1112
rect 2159 1108 2163 1112
rect 2231 1108 2235 1112
rect 2303 1108 2307 1112
rect 2359 1108 2363 1112
rect 135 1092 139 1096
rect 175 1092 179 1096
rect 247 1092 251 1096
rect 327 1092 331 1096
rect 415 1092 419 1096
rect 503 1092 507 1096
rect 583 1092 587 1096
rect 663 1092 667 1096
rect 735 1092 739 1096
rect 799 1092 803 1096
rect 863 1092 867 1096
rect 919 1092 923 1096
rect 983 1092 987 1096
rect 1047 1092 1051 1096
rect 1431 1096 1435 1100
rect 1471 1096 1475 1100
rect 1511 1096 1515 1100
rect 1559 1096 1563 1100
rect 1615 1096 1619 1100
rect 1671 1096 1675 1100
rect 1727 1096 1731 1100
rect 1775 1096 1779 1100
rect 1823 1096 1827 1100
rect 1871 1096 1875 1100
rect 1919 1096 1923 1100
rect 1967 1096 1971 1100
rect 2015 1096 2019 1100
rect 2063 1096 2067 1100
rect 2119 1096 2123 1100
rect 2175 1096 2179 1100
rect 2231 1096 2235 1100
rect 111 1085 115 1089
rect 1239 1085 1243 1089
rect 1279 1089 1283 1093
rect 2407 1089 2411 1093
rect 111 1068 115 1072
rect 1239 1068 1243 1072
rect 1279 1072 1283 1076
rect 2407 1072 2411 1076
rect 135 1045 139 1049
rect 175 1045 179 1049
rect 247 1045 251 1049
rect 327 1045 331 1049
rect 415 1045 419 1049
rect 503 1045 507 1049
rect 583 1045 587 1049
rect 663 1045 667 1049
rect 735 1045 739 1049
rect 799 1045 803 1049
rect 863 1045 867 1049
rect 919 1045 923 1049
rect 983 1045 987 1049
rect 1047 1045 1051 1049
rect 1431 1049 1435 1053
rect 1471 1049 1475 1053
rect 1511 1049 1515 1053
rect 1559 1049 1563 1053
rect 1615 1049 1619 1053
rect 1671 1049 1675 1053
rect 1727 1049 1731 1053
rect 1775 1049 1779 1053
rect 1823 1049 1827 1053
rect 1871 1049 1875 1053
rect 1919 1049 1923 1053
rect 1967 1049 1971 1053
rect 2015 1049 2019 1053
rect 2063 1049 2067 1053
rect 2119 1049 2123 1053
rect 2175 1049 2179 1053
rect 2231 1049 2235 1053
rect 175 1015 179 1019
rect 255 1015 259 1019
rect 327 1015 331 1019
rect 399 1015 403 1019
rect 463 1015 467 1019
rect 519 1015 523 1019
rect 575 1015 579 1019
rect 623 1015 627 1019
rect 671 1015 675 1019
rect 735 1015 739 1019
rect 807 1015 811 1019
rect 895 1015 899 1019
rect 999 1015 1003 1019
rect 1103 1015 1107 1019
rect 1191 1015 1195 1019
rect 1575 1019 1579 1023
rect 1615 1019 1619 1023
rect 1655 1019 1659 1023
rect 1695 1019 1699 1023
rect 1735 1019 1739 1023
rect 1775 1019 1779 1023
rect 1823 1019 1827 1023
rect 1879 1019 1883 1023
rect 1943 1019 1947 1023
rect 2015 1019 2019 1023
rect 2095 1019 2099 1023
rect 2175 1019 2179 1023
rect 2255 1019 2259 1023
rect 111 992 115 996
rect 1239 992 1243 996
rect 1279 996 1283 1000
rect 2407 996 2411 1000
rect 111 975 115 979
rect 1239 975 1243 979
rect 1279 979 1283 983
rect 2407 979 2411 983
rect 175 968 179 972
rect 255 968 259 972
rect 327 968 331 972
rect 399 968 403 972
rect 463 968 467 972
rect 519 968 523 972
rect 575 968 579 972
rect 623 968 627 972
rect 671 968 675 972
rect 735 968 739 972
rect 807 968 811 972
rect 895 968 899 972
rect 999 968 1003 972
rect 1103 968 1107 972
rect 1191 968 1195 972
rect 1575 972 1579 976
rect 1615 972 1619 976
rect 1655 972 1659 976
rect 1695 972 1699 976
rect 1735 972 1739 976
rect 1775 972 1779 976
rect 1823 972 1827 976
rect 1879 972 1883 976
rect 1943 972 1947 976
rect 2015 972 2019 976
rect 2095 972 2099 976
rect 2175 972 2179 976
rect 2255 972 2259 976
rect 215 956 219 960
rect 255 956 259 960
rect 303 956 307 960
rect 359 956 363 960
rect 415 956 419 960
rect 463 956 467 960
rect 519 956 523 960
rect 575 956 579 960
rect 639 956 643 960
rect 711 956 715 960
rect 783 956 787 960
rect 855 956 859 960
rect 927 956 931 960
rect 999 956 1003 960
rect 1071 956 1075 960
rect 1143 956 1147 960
rect 1191 956 1195 960
rect 111 949 115 953
rect 1239 949 1243 953
rect 1303 952 1307 956
rect 1351 952 1355 956
rect 1431 952 1435 956
rect 1511 952 1515 956
rect 1591 952 1595 956
rect 1679 952 1683 956
rect 1767 952 1771 956
rect 1855 952 1859 956
rect 1943 952 1947 956
rect 2023 952 2027 956
rect 2103 952 2107 956
rect 2183 952 2187 956
rect 2271 952 2275 956
rect 1279 945 1283 949
rect 2407 945 2411 949
rect 111 932 115 936
rect 1239 932 1243 936
rect 1279 928 1283 932
rect 2407 928 2411 932
rect 215 909 219 913
rect 255 909 259 913
rect 303 909 307 913
rect 359 909 363 913
rect 415 909 419 913
rect 463 909 467 913
rect 519 909 523 913
rect 575 909 579 913
rect 639 909 643 913
rect 711 909 715 913
rect 783 909 787 913
rect 855 909 859 913
rect 927 909 931 913
rect 999 909 1003 913
rect 1071 909 1075 913
rect 1143 909 1147 913
rect 1191 909 1195 913
rect 1303 905 1307 909
rect 1351 905 1355 909
rect 1431 905 1435 909
rect 1511 905 1515 909
rect 1591 905 1595 909
rect 1679 905 1683 909
rect 1767 905 1771 909
rect 1855 905 1859 909
rect 1943 905 1947 909
rect 2023 905 2027 909
rect 2103 905 2107 909
rect 2183 905 2187 909
rect 2271 905 2275 909
rect 191 871 195 875
rect 231 871 235 875
rect 287 871 291 875
rect 359 871 363 875
rect 447 871 451 875
rect 543 871 547 875
rect 639 871 643 875
rect 727 871 731 875
rect 807 871 811 875
rect 887 871 891 875
rect 959 871 963 875
rect 1023 871 1027 875
rect 1087 871 1091 875
rect 1159 871 1163 875
rect 1439 875 1443 879
rect 1479 875 1483 879
rect 1519 875 1523 879
rect 1559 875 1563 879
rect 1607 875 1611 879
rect 1655 875 1659 879
rect 1711 875 1715 879
rect 1775 875 1779 879
rect 1847 875 1851 879
rect 1919 875 1923 879
rect 1991 875 1995 879
rect 2063 875 2067 879
rect 2135 875 2139 879
rect 2215 875 2219 879
rect 2295 875 2299 879
rect 111 848 115 852
rect 1239 848 1243 852
rect 1279 852 1283 856
rect 2407 852 2411 856
rect 111 831 115 835
rect 1239 831 1243 835
rect 1279 835 1283 839
rect 2407 835 2411 839
rect 191 824 195 828
rect 231 824 235 828
rect 287 824 291 828
rect 359 824 363 828
rect 447 824 451 828
rect 543 824 547 828
rect 639 824 643 828
rect 727 824 731 828
rect 807 824 811 828
rect 887 824 891 828
rect 959 824 963 828
rect 1023 824 1027 828
rect 1087 824 1091 828
rect 1159 824 1163 828
rect 1439 828 1443 832
rect 1479 828 1483 832
rect 1519 828 1523 832
rect 1559 828 1563 832
rect 1607 828 1611 832
rect 1655 828 1659 832
rect 1711 828 1715 832
rect 1775 828 1779 832
rect 1847 828 1851 832
rect 1919 828 1923 832
rect 1991 828 1995 832
rect 2063 828 2067 832
rect 2135 828 2139 832
rect 2215 828 2219 832
rect 2295 828 2299 832
rect 135 812 139 816
rect 175 812 179 816
rect 239 812 243 816
rect 327 812 331 816
rect 415 812 419 816
rect 503 812 507 816
rect 591 812 595 816
rect 671 812 675 816
rect 743 812 747 816
rect 815 812 819 816
rect 879 812 883 816
rect 943 812 947 816
rect 1015 812 1019 816
rect 111 805 115 809
rect 1239 805 1243 809
rect 1359 804 1363 808
rect 1415 804 1419 808
rect 1471 804 1475 808
rect 1535 804 1539 808
rect 1591 804 1595 808
rect 1647 804 1651 808
rect 1703 804 1707 808
rect 1759 804 1763 808
rect 1815 804 1819 808
rect 1871 804 1875 808
rect 1935 804 1939 808
rect 1999 804 2003 808
rect 2071 804 2075 808
rect 2143 804 2147 808
rect 2223 804 2227 808
rect 2303 804 2307 808
rect 2359 804 2363 808
rect 1279 797 1283 801
rect 2407 797 2411 801
rect 111 788 115 792
rect 1239 788 1243 792
rect 1279 780 1283 784
rect 2407 780 2411 784
rect 135 765 139 769
rect 175 765 179 769
rect 239 765 243 769
rect 327 765 331 769
rect 415 765 419 769
rect 503 765 507 769
rect 591 765 595 769
rect 671 765 675 769
rect 743 765 747 769
rect 815 765 819 769
rect 879 765 883 769
rect 943 765 947 769
rect 1015 765 1019 769
rect 1359 757 1363 761
rect 1415 757 1419 761
rect 1471 757 1475 761
rect 1535 757 1539 761
rect 1591 757 1595 761
rect 1647 757 1651 761
rect 1703 757 1707 761
rect 1759 757 1763 761
rect 1815 757 1819 761
rect 1871 757 1875 761
rect 1935 757 1939 761
rect 1999 757 2003 761
rect 2071 757 2075 761
rect 2143 757 2147 761
rect 2223 757 2227 761
rect 2303 757 2307 761
rect 2359 757 2363 761
rect 135 731 139 735
rect 191 731 195 735
rect 263 731 267 735
rect 335 731 339 735
rect 399 731 403 735
rect 455 731 459 735
rect 503 731 507 735
rect 543 731 547 735
rect 583 731 587 735
rect 623 731 627 735
rect 671 731 675 735
rect 719 731 723 735
rect 767 731 771 735
rect 815 731 819 735
rect 863 731 867 735
rect 911 731 915 735
rect 1303 727 1307 731
rect 1343 727 1347 731
rect 1407 727 1411 731
rect 1487 727 1491 731
rect 1575 727 1579 731
rect 1663 727 1667 731
rect 1751 727 1755 731
rect 1831 727 1835 731
rect 1911 727 1915 731
rect 1991 727 1995 731
rect 2079 727 2083 731
rect 2175 727 2179 731
rect 2279 727 2283 731
rect 2359 727 2363 731
rect 111 708 115 712
rect 1239 708 1243 712
rect 1279 704 1283 708
rect 2407 704 2411 708
rect 111 691 115 695
rect 1239 691 1243 695
rect 135 684 139 688
rect 191 684 195 688
rect 263 684 267 688
rect 335 684 339 688
rect 399 684 403 688
rect 455 684 459 688
rect 503 684 507 688
rect 543 684 547 688
rect 583 684 587 688
rect 623 684 627 688
rect 671 684 675 688
rect 719 684 723 688
rect 767 684 771 688
rect 815 684 819 688
rect 863 684 867 688
rect 911 684 915 688
rect 1279 687 1283 691
rect 2407 687 2411 691
rect 1303 680 1307 684
rect 1343 680 1347 684
rect 1407 680 1411 684
rect 1487 680 1491 684
rect 1575 680 1579 684
rect 1663 680 1667 684
rect 1751 680 1755 684
rect 1831 680 1835 684
rect 1911 680 1915 684
rect 1991 680 1995 684
rect 2079 680 2083 684
rect 2175 680 2179 684
rect 2279 680 2283 684
rect 2359 680 2363 684
rect 135 668 139 672
rect 199 668 203 672
rect 279 668 283 672
rect 351 668 355 672
rect 415 668 419 672
rect 487 668 491 672
rect 559 668 563 672
rect 639 668 643 672
rect 711 668 715 672
rect 783 668 787 672
rect 855 668 859 672
rect 919 668 923 672
rect 983 668 987 672
rect 1039 668 1043 672
rect 1095 668 1099 672
rect 1151 668 1155 672
rect 1191 668 1195 672
rect 111 661 115 665
rect 1239 661 1243 665
rect 1303 664 1307 668
rect 1399 664 1403 668
rect 1511 664 1515 668
rect 1623 664 1627 668
rect 1727 664 1731 668
rect 1815 664 1819 668
rect 1895 664 1899 668
rect 1975 664 1979 668
rect 2047 664 2051 668
rect 2111 664 2115 668
rect 2175 664 2179 668
rect 2239 664 2243 668
rect 2311 664 2315 668
rect 2359 664 2363 668
rect 1279 657 1283 661
rect 2407 657 2411 661
rect 111 644 115 648
rect 1239 644 1243 648
rect 1279 640 1283 644
rect 2407 640 2411 644
rect 135 621 139 625
rect 199 621 203 625
rect 279 621 283 625
rect 351 621 355 625
rect 415 621 419 625
rect 487 621 491 625
rect 559 621 563 625
rect 639 621 643 625
rect 711 621 715 625
rect 783 621 787 625
rect 855 621 859 625
rect 919 621 923 625
rect 983 621 987 625
rect 1039 621 1043 625
rect 1095 621 1099 625
rect 1151 621 1155 625
rect 1191 621 1195 625
rect 1303 617 1307 621
rect 1399 617 1403 621
rect 1511 617 1515 621
rect 1623 617 1627 621
rect 1727 617 1731 621
rect 1815 617 1819 621
rect 1895 617 1899 621
rect 1975 617 1979 621
rect 2047 617 2051 621
rect 2111 617 2115 621
rect 2175 617 2179 621
rect 2239 617 2243 621
rect 2311 617 2315 621
rect 2359 617 2363 621
rect 135 583 139 587
rect 191 583 195 587
rect 271 583 275 587
rect 359 583 363 587
rect 447 583 451 587
rect 535 583 539 587
rect 623 583 627 587
rect 703 583 707 587
rect 783 583 787 587
rect 855 583 859 587
rect 919 583 923 587
rect 975 583 979 587
rect 1023 583 1027 587
rect 1079 583 1083 587
rect 1135 583 1139 587
rect 1191 583 1195 587
rect 1415 583 1419 587
rect 1455 583 1459 587
rect 1495 583 1499 587
rect 1543 583 1547 587
rect 1599 583 1603 587
rect 1663 583 1667 587
rect 1727 583 1731 587
rect 1791 583 1795 587
rect 1847 583 1851 587
rect 1911 583 1915 587
rect 1975 583 1979 587
rect 2047 583 2051 587
rect 2119 583 2123 587
rect 2199 583 2203 587
rect 2287 583 2291 587
rect 2359 583 2363 587
rect 111 560 115 564
rect 1239 560 1243 564
rect 1279 560 1283 564
rect 2407 560 2411 564
rect 111 543 115 547
rect 1239 543 1243 547
rect 1279 543 1283 547
rect 2407 543 2411 547
rect 135 536 139 540
rect 191 536 195 540
rect 271 536 275 540
rect 359 536 363 540
rect 447 536 451 540
rect 535 536 539 540
rect 623 536 627 540
rect 703 536 707 540
rect 783 536 787 540
rect 855 536 859 540
rect 919 536 923 540
rect 975 536 979 540
rect 1023 536 1027 540
rect 1079 536 1083 540
rect 1135 536 1139 540
rect 1191 536 1195 540
rect 1415 536 1419 540
rect 1455 536 1459 540
rect 1495 536 1499 540
rect 1543 536 1547 540
rect 1599 536 1603 540
rect 1663 536 1667 540
rect 1727 536 1731 540
rect 1791 536 1795 540
rect 1847 536 1851 540
rect 1911 536 1915 540
rect 1975 536 1979 540
rect 2047 536 2051 540
rect 2119 536 2123 540
rect 2199 536 2203 540
rect 2287 536 2291 540
rect 2359 536 2363 540
rect 1303 524 1307 528
rect 1375 524 1379 528
rect 1479 524 1483 528
rect 1583 524 1587 528
rect 1695 524 1699 528
rect 1799 524 1803 528
rect 1903 524 1907 528
rect 2007 524 2011 528
rect 2103 524 2107 528
rect 2191 524 2195 528
rect 2287 524 2291 528
rect 2359 524 2363 528
rect 135 516 139 520
rect 191 516 195 520
rect 263 516 267 520
rect 335 516 339 520
rect 415 516 419 520
rect 495 516 499 520
rect 575 516 579 520
rect 647 516 651 520
rect 719 516 723 520
rect 783 516 787 520
rect 847 516 851 520
rect 903 516 907 520
rect 959 516 963 520
rect 1023 516 1027 520
rect 1087 516 1091 520
rect 1151 516 1155 520
rect 1191 516 1195 520
rect 1279 517 1283 521
rect 2407 517 2411 521
rect 111 509 115 513
rect 1239 509 1243 513
rect 1279 500 1283 504
rect 2407 500 2411 504
rect 111 492 115 496
rect 1239 492 1243 496
rect 1303 477 1307 481
rect 1375 477 1379 481
rect 1479 477 1483 481
rect 1583 477 1587 481
rect 1695 477 1699 481
rect 1799 477 1803 481
rect 1903 477 1907 481
rect 2007 477 2011 481
rect 2103 477 2107 481
rect 2191 477 2195 481
rect 2287 477 2291 481
rect 2359 477 2363 481
rect 135 469 139 473
rect 191 469 195 473
rect 263 469 267 473
rect 335 469 339 473
rect 415 469 419 473
rect 495 469 499 473
rect 575 469 579 473
rect 647 469 651 473
rect 719 469 723 473
rect 783 469 787 473
rect 847 469 851 473
rect 903 469 907 473
rect 959 469 963 473
rect 1023 469 1027 473
rect 1087 469 1091 473
rect 1151 469 1155 473
rect 1191 469 1195 473
rect 183 439 187 443
rect 223 439 227 443
rect 263 439 267 443
rect 311 439 315 443
rect 367 439 371 443
rect 431 439 435 443
rect 495 439 499 443
rect 559 439 563 443
rect 615 439 619 443
rect 671 439 675 443
rect 719 439 723 443
rect 775 439 779 443
rect 831 439 835 443
rect 887 439 891 443
rect 1303 443 1307 447
rect 1343 443 1347 447
rect 1399 443 1403 447
rect 1463 443 1467 447
rect 1527 443 1531 447
rect 1591 443 1595 447
rect 1663 443 1667 447
rect 1735 443 1739 447
rect 1815 443 1819 447
rect 1895 443 1899 447
rect 1975 443 1979 447
rect 2055 443 2059 447
rect 2135 443 2139 447
rect 2215 443 2219 447
rect 2295 443 2299 447
rect 2359 443 2363 447
rect 111 416 115 420
rect 1239 416 1243 420
rect 1279 420 1283 424
rect 2407 420 2411 424
rect 111 399 115 403
rect 1239 399 1243 403
rect 1279 403 1283 407
rect 2407 403 2411 407
rect 183 392 187 396
rect 223 392 227 396
rect 263 392 267 396
rect 311 392 315 396
rect 367 392 371 396
rect 431 392 435 396
rect 495 392 499 396
rect 559 392 563 396
rect 615 392 619 396
rect 671 392 675 396
rect 719 392 723 396
rect 775 392 779 396
rect 831 392 835 396
rect 887 392 891 396
rect 1303 396 1307 400
rect 1343 396 1347 400
rect 1399 396 1403 400
rect 1463 396 1467 400
rect 1527 396 1531 400
rect 1591 396 1595 400
rect 1663 396 1667 400
rect 1735 396 1739 400
rect 1815 396 1819 400
rect 1895 396 1899 400
rect 1975 396 1979 400
rect 2055 396 2059 400
rect 2135 396 2139 400
rect 2215 396 2219 400
rect 2295 396 2299 400
rect 2359 396 2363 400
rect 135 380 139 384
rect 175 380 179 384
rect 231 380 235 384
rect 287 380 291 384
rect 343 380 347 384
rect 391 380 395 384
rect 439 380 443 384
rect 487 380 491 384
rect 535 380 539 384
rect 583 380 587 384
rect 631 380 635 384
rect 679 380 683 384
rect 727 380 731 384
rect 775 380 779 384
rect 1447 380 1451 384
rect 1487 380 1491 384
rect 1535 380 1539 384
rect 1591 380 1595 384
rect 1663 380 1667 384
rect 1735 380 1739 384
rect 1815 380 1819 384
rect 1895 380 1899 384
rect 1967 380 1971 384
rect 2039 380 2043 384
rect 2111 380 2115 384
rect 2175 380 2179 384
rect 2239 380 2243 384
rect 2303 380 2307 384
rect 2359 380 2363 384
rect 111 373 115 377
rect 1239 373 1243 377
rect 1279 373 1283 377
rect 2407 373 2411 377
rect 111 356 115 360
rect 1239 356 1243 360
rect 1279 356 1283 360
rect 2407 356 2411 360
rect 135 333 139 337
rect 175 333 179 337
rect 231 333 235 337
rect 287 333 291 337
rect 343 333 347 337
rect 391 333 395 337
rect 439 333 443 337
rect 487 333 491 337
rect 535 333 539 337
rect 583 333 587 337
rect 631 333 635 337
rect 679 333 683 337
rect 727 333 731 337
rect 775 333 779 337
rect 1447 333 1451 337
rect 1487 333 1491 337
rect 1535 333 1539 337
rect 1591 333 1595 337
rect 1663 333 1667 337
rect 1735 333 1739 337
rect 1815 333 1819 337
rect 1895 333 1899 337
rect 1967 333 1971 337
rect 2039 333 2043 337
rect 2111 333 2115 337
rect 2175 333 2179 337
rect 2239 333 2243 337
rect 2303 333 2307 337
rect 2359 333 2363 337
rect 135 299 139 303
rect 183 299 187 303
rect 255 299 259 303
rect 327 299 331 303
rect 391 299 395 303
rect 447 299 451 303
rect 503 299 507 303
rect 551 299 555 303
rect 591 299 595 303
rect 631 299 635 303
rect 679 299 683 303
rect 727 299 731 303
rect 775 299 779 303
rect 823 299 827 303
rect 871 299 875 303
rect 919 299 923 303
rect 1495 299 1499 303
rect 1535 299 1539 303
rect 1575 299 1579 303
rect 1615 299 1619 303
rect 1655 299 1659 303
rect 1695 299 1699 303
rect 1743 299 1747 303
rect 1799 299 1803 303
rect 1863 299 1867 303
rect 1935 299 1939 303
rect 2007 299 2011 303
rect 2071 299 2075 303
rect 2135 299 2139 303
rect 2191 299 2195 303
rect 2255 299 2259 303
rect 2319 299 2323 303
rect 2359 299 2363 303
rect 111 276 115 280
rect 1239 276 1243 280
rect 1279 276 1283 280
rect 2407 276 2411 280
rect 111 259 115 263
rect 1239 259 1243 263
rect 1279 259 1283 263
rect 2407 259 2411 263
rect 135 252 139 256
rect 183 252 187 256
rect 255 252 259 256
rect 327 252 331 256
rect 391 252 395 256
rect 447 252 451 256
rect 503 252 507 256
rect 551 252 555 256
rect 591 252 595 256
rect 631 252 635 256
rect 679 252 683 256
rect 727 252 731 256
rect 775 252 779 256
rect 823 252 827 256
rect 871 252 875 256
rect 919 252 923 256
rect 1495 252 1499 256
rect 1535 252 1539 256
rect 1575 252 1579 256
rect 1615 252 1619 256
rect 1655 252 1659 256
rect 1695 252 1699 256
rect 1743 252 1747 256
rect 1799 252 1803 256
rect 1863 252 1867 256
rect 1935 252 1939 256
rect 2007 252 2011 256
rect 2071 252 2075 256
rect 2135 252 2139 256
rect 2191 252 2195 256
rect 2255 252 2259 256
rect 2319 252 2323 256
rect 2359 252 2363 256
rect 135 232 139 236
rect 175 232 179 236
rect 247 232 251 236
rect 327 232 331 236
rect 415 232 419 236
rect 495 232 499 236
rect 575 232 579 236
rect 655 232 659 236
rect 727 232 731 236
rect 791 232 795 236
rect 847 232 851 236
rect 903 232 907 236
rect 959 232 963 236
rect 1023 232 1027 236
rect 1367 236 1371 240
rect 1407 236 1411 240
rect 1447 236 1451 240
rect 1495 236 1499 240
rect 1551 236 1555 240
rect 1607 236 1611 240
rect 1671 236 1675 240
rect 1735 236 1739 240
rect 1807 236 1811 240
rect 1887 236 1891 240
rect 1975 236 1979 240
rect 2071 236 2075 240
rect 2167 236 2171 240
rect 2271 236 2275 240
rect 2359 236 2363 240
rect 111 225 115 229
rect 1239 225 1243 229
rect 1279 229 1283 233
rect 2407 229 2411 233
rect 111 208 115 212
rect 1239 208 1243 212
rect 1279 212 1283 216
rect 2407 212 2411 216
rect 135 185 139 189
rect 175 185 179 189
rect 247 185 251 189
rect 327 185 331 189
rect 415 185 419 189
rect 495 185 499 189
rect 575 185 579 189
rect 655 185 659 189
rect 727 185 731 189
rect 791 185 795 189
rect 847 185 851 189
rect 903 185 907 189
rect 959 185 963 189
rect 1023 185 1027 189
rect 1367 189 1371 193
rect 1407 189 1411 193
rect 1447 189 1451 193
rect 1495 189 1499 193
rect 1551 189 1555 193
rect 1607 189 1611 193
rect 1671 189 1675 193
rect 1735 189 1739 193
rect 1807 189 1811 193
rect 1887 189 1891 193
rect 1975 189 1979 193
rect 2071 189 2075 193
rect 2167 189 2171 193
rect 2271 189 2275 193
rect 2359 189 2363 193
rect 1303 143 1307 147
rect 1343 143 1347 147
rect 1383 143 1387 147
rect 1423 143 1427 147
rect 1463 143 1467 147
rect 1519 143 1523 147
rect 1583 143 1587 147
rect 1647 143 1651 147
rect 1711 143 1715 147
rect 1767 143 1771 147
rect 1823 143 1827 147
rect 1871 143 1875 147
rect 1919 143 1923 147
rect 1967 143 1971 147
rect 2015 143 2019 147
rect 2063 143 2067 147
rect 2111 143 2115 147
rect 2159 143 2163 147
rect 2215 143 2219 147
rect 2271 143 2275 147
rect 2319 143 2323 147
rect 2359 143 2363 147
rect 135 135 139 139
rect 175 135 179 139
rect 215 135 219 139
rect 255 135 259 139
rect 295 135 299 139
rect 335 135 339 139
rect 375 135 379 139
rect 423 135 427 139
rect 471 135 475 139
rect 527 135 531 139
rect 583 135 587 139
rect 631 135 635 139
rect 679 135 683 139
rect 727 135 731 139
rect 767 135 771 139
rect 807 135 811 139
rect 847 135 851 139
rect 887 135 891 139
rect 927 135 931 139
rect 975 135 979 139
rect 1023 135 1027 139
rect 1071 135 1075 139
rect 1111 135 1115 139
rect 1151 135 1155 139
rect 1191 135 1195 139
rect 1279 120 1283 124
rect 2407 120 2411 124
rect 111 112 115 116
rect 1239 112 1243 116
rect 1279 103 1283 107
rect 2407 103 2411 107
rect 111 95 115 99
rect 1239 95 1243 99
rect 1303 96 1307 100
rect 1343 96 1347 100
rect 1383 96 1387 100
rect 1423 96 1427 100
rect 1463 96 1467 100
rect 1519 96 1523 100
rect 1583 96 1587 100
rect 1647 96 1651 100
rect 1711 96 1715 100
rect 1767 96 1771 100
rect 1823 96 1827 100
rect 1871 96 1875 100
rect 1919 96 1923 100
rect 1967 96 1971 100
rect 2015 96 2019 100
rect 2063 96 2067 100
rect 2111 96 2115 100
rect 2159 96 2163 100
rect 2215 96 2219 100
rect 2271 96 2275 100
rect 2319 96 2323 100
rect 2359 96 2363 100
rect 135 88 139 92
rect 175 88 179 92
rect 215 88 219 92
rect 255 88 259 92
rect 295 88 299 92
rect 335 88 339 92
rect 375 88 379 92
rect 423 88 427 92
rect 471 88 475 92
rect 527 88 531 92
rect 583 88 587 92
rect 631 88 635 92
rect 679 88 683 92
rect 727 88 731 92
rect 767 88 771 92
rect 807 88 811 92
rect 847 88 851 92
rect 887 88 891 92
rect 927 88 931 92
rect 975 88 979 92
rect 1023 88 1027 92
rect 1071 88 1075 92
rect 1111 88 1115 92
rect 1151 88 1155 92
rect 1191 88 1195 92
<< m3 >>
rect 1279 2514 1283 2515
rect 1279 2509 1283 2510
rect 1535 2514 1539 2515
rect 1535 2509 1539 2510
rect 1575 2514 1579 2515
rect 1575 2509 1579 2510
rect 1615 2514 1619 2515
rect 1615 2509 1619 2510
rect 1655 2514 1659 2515
rect 1655 2509 1659 2510
rect 1695 2514 1699 2515
rect 1695 2509 1699 2510
rect 1735 2514 1739 2515
rect 1735 2509 1739 2510
rect 1775 2514 1779 2515
rect 1775 2509 1779 2510
rect 1815 2514 1819 2515
rect 1815 2509 1819 2510
rect 1855 2514 1859 2515
rect 1855 2509 1859 2510
rect 1895 2514 1899 2515
rect 1895 2509 1899 2510
rect 1935 2514 1939 2515
rect 1935 2509 1939 2510
rect 1975 2514 1979 2515
rect 1975 2509 1979 2510
rect 2407 2514 2411 2515
rect 2407 2509 2411 2510
rect 111 2502 115 2503
rect 111 2497 115 2498
rect 135 2502 139 2503
rect 135 2497 139 2498
rect 175 2502 179 2503
rect 175 2497 179 2498
rect 215 2502 219 2503
rect 215 2497 219 2498
rect 255 2502 259 2503
rect 255 2497 259 2498
rect 311 2502 315 2503
rect 311 2497 315 2498
rect 391 2502 395 2503
rect 391 2497 395 2498
rect 479 2502 483 2503
rect 479 2497 483 2498
rect 567 2502 571 2503
rect 567 2497 571 2498
rect 655 2502 659 2503
rect 655 2497 659 2498
rect 743 2502 747 2503
rect 743 2497 747 2498
rect 831 2502 835 2503
rect 831 2497 835 2498
rect 927 2502 931 2503
rect 927 2497 931 2498
rect 1239 2502 1243 2503
rect 1280 2502 1282 2509
rect 1534 2508 1540 2509
rect 1534 2504 1535 2508
rect 1539 2504 1540 2508
rect 1534 2503 1540 2504
rect 1574 2508 1580 2509
rect 1574 2504 1575 2508
rect 1579 2504 1580 2508
rect 1574 2503 1580 2504
rect 1614 2508 1620 2509
rect 1614 2504 1615 2508
rect 1619 2504 1620 2508
rect 1614 2503 1620 2504
rect 1654 2508 1660 2509
rect 1654 2504 1655 2508
rect 1659 2504 1660 2508
rect 1654 2503 1660 2504
rect 1694 2508 1700 2509
rect 1694 2504 1695 2508
rect 1699 2504 1700 2508
rect 1694 2503 1700 2504
rect 1734 2508 1740 2509
rect 1734 2504 1735 2508
rect 1739 2504 1740 2508
rect 1734 2503 1740 2504
rect 1774 2508 1780 2509
rect 1774 2504 1775 2508
rect 1779 2504 1780 2508
rect 1774 2503 1780 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1814 2503 1820 2504
rect 1854 2508 1860 2509
rect 1854 2504 1855 2508
rect 1859 2504 1860 2508
rect 1854 2503 1860 2504
rect 1894 2508 1900 2509
rect 1894 2504 1895 2508
rect 1899 2504 1900 2508
rect 1894 2503 1900 2504
rect 1934 2508 1940 2509
rect 1934 2504 1935 2508
rect 1939 2504 1940 2508
rect 1934 2503 1940 2504
rect 1974 2508 1980 2509
rect 1974 2504 1975 2508
rect 1979 2504 1980 2508
rect 1974 2503 1980 2504
rect 2408 2502 2410 2509
rect 1239 2497 1243 2498
rect 1278 2501 1284 2502
rect 1278 2497 1279 2501
rect 1283 2497 1284 2501
rect 112 2465 114 2497
rect 136 2488 138 2497
rect 176 2488 178 2497
rect 216 2488 218 2497
rect 256 2488 258 2497
rect 312 2488 314 2497
rect 392 2488 394 2497
rect 480 2488 482 2497
rect 568 2488 570 2497
rect 656 2488 658 2497
rect 744 2488 746 2497
rect 832 2488 834 2497
rect 928 2488 930 2497
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 174 2487 180 2488
rect 174 2483 175 2487
rect 179 2483 180 2487
rect 174 2482 180 2483
rect 214 2487 220 2488
rect 214 2483 215 2487
rect 219 2483 220 2487
rect 214 2482 220 2483
rect 254 2487 260 2488
rect 254 2483 255 2487
rect 259 2483 260 2487
rect 254 2482 260 2483
rect 310 2487 316 2488
rect 310 2483 311 2487
rect 315 2483 316 2487
rect 310 2482 316 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 478 2487 484 2488
rect 478 2483 479 2487
rect 483 2483 484 2487
rect 478 2482 484 2483
rect 566 2487 572 2488
rect 566 2483 567 2487
rect 571 2483 572 2487
rect 566 2482 572 2483
rect 654 2487 660 2488
rect 654 2483 655 2487
rect 659 2483 660 2487
rect 654 2482 660 2483
rect 742 2487 748 2488
rect 742 2483 743 2487
rect 747 2483 748 2487
rect 742 2482 748 2483
rect 830 2487 836 2488
rect 830 2483 831 2487
rect 835 2483 836 2487
rect 830 2482 836 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 1240 2465 1242 2497
rect 1278 2496 1284 2497
rect 2406 2501 2412 2502
rect 2406 2497 2407 2501
rect 2411 2497 2412 2501
rect 2406 2496 2412 2497
rect 1278 2484 1284 2485
rect 1278 2480 1279 2484
rect 1283 2480 1284 2484
rect 1278 2479 1284 2480
rect 2406 2484 2412 2485
rect 2406 2480 2407 2484
rect 2411 2480 2412 2484
rect 2406 2479 2412 2480
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 110 2459 116 2460
rect 1238 2464 1244 2465
rect 1238 2460 1239 2464
rect 1243 2460 1244 2464
rect 1238 2459 1244 2460
rect 110 2447 116 2448
rect 110 2443 111 2447
rect 115 2443 116 2447
rect 110 2442 116 2443
rect 1238 2447 1244 2448
rect 1280 2447 1282 2479
rect 1534 2461 1540 2462
rect 1534 2457 1535 2461
rect 1539 2457 1540 2461
rect 1534 2456 1540 2457
rect 1574 2461 1580 2462
rect 1574 2457 1575 2461
rect 1579 2457 1580 2461
rect 1574 2456 1580 2457
rect 1614 2461 1620 2462
rect 1614 2457 1615 2461
rect 1619 2457 1620 2461
rect 1614 2456 1620 2457
rect 1654 2461 1660 2462
rect 1654 2457 1655 2461
rect 1659 2457 1660 2461
rect 1654 2456 1660 2457
rect 1694 2461 1700 2462
rect 1694 2457 1695 2461
rect 1699 2457 1700 2461
rect 1694 2456 1700 2457
rect 1734 2461 1740 2462
rect 1734 2457 1735 2461
rect 1739 2457 1740 2461
rect 1734 2456 1740 2457
rect 1774 2461 1780 2462
rect 1774 2457 1775 2461
rect 1779 2457 1780 2461
rect 1774 2456 1780 2457
rect 1814 2461 1820 2462
rect 1814 2457 1815 2461
rect 1819 2457 1820 2461
rect 1814 2456 1820 2457
rect 1854 2461 1860 2462
rect 1854 2457 1855 2461
rect 1859 2457 1860 2461
rect 1854 2456 1860 2457
rect 1894 2461 1900 2462
rect 1894 2457 1895 2461
rect 1899 2457 1900 2461
rect 1894 2456 1900 2457
rect 1934 2461 1940 2462
rect 1934 2457 1935 2461
rect 1939 2457 1940 2461
rect 1934 2456 1940 2457
rect 1974 2461 1980 2462
rect 1974 2457 1975 2461
rect 1979 2457 1980 2461
rect 1974 2456 1980 2457
rect 1536 2447 1538 2456
rect 1576 2447 1578 2456
rect 1616 2447 1618 2456
rect 1656 2447 1658 2456
rect 1696 2447 1698 2456
rect 1736 2447 1738 2456
rect 1776 2447 1778 2456
rect 1816 2447 1818 2456
rect 1856 2447 1858 2456
rect 1896 2447 1898 2456
rect 1936 2447 1938 2456
rect 1976 2447 1978 2456
rect 2408 2447 2410 2479
rect 1238 2443 1239 2447
rect 1243 2443 1244 2447
rect 1238 2442 1244 2443
rect 1279 2446 1283 2447
rect 112 2435 114 2442
rect 134 2440 140 2441
rect 134 2436 135 2440
rect 139 2436 140 2440
rect 134 2435 140 2436
rect 174 2440 180 2441
rect 174 2436 175 2440
rect 179 2436 180 2440
rect 174 2435 180 2436
rect 214 2440 220 2441
rect 214 2436 215 2440
rect 219 2436 220 2440
rect 214 2435 220 2436
rect 254 2440 260 2441
rect 254 2436 255 2440
rect 259 2436 260 2440
rect 254 2435 260 2436
rect 310 2440 316 2441
rect 310 2436 311 2440
rect 315 2436 316 2440
rect 310 2435 316 2436
rect 390 2440 396 2441
rect 390 2436 391 2440
rect 395 2436 396 2440
rect 390 2435 396 2436
rect 478 2440 484 2441
rect 478 2436 479 2440
rect 483 2436 484 2440
rect 478 2435 484 2436
rect 566 2440 572 2441
rect 566 2436 567 2440
rect 571 2436 572 2440
rect 566 2435 572 2436
rect 654 2440 660 2441
rect 654 2436 655 2440
rect 659 2436 660 2440
rect 654 2435 660 2436
rect 742 2440 748 2441
rect 742 2436 743 2440
rect 747 2436 748 2440
rect 742 2435 748 2436
rect 830 2440 836 2441
rect 830 2436 831 2440
rect 835 2436 836 2440
rect 830 2435 836 2436
rect 926 2440 932 2441
rect 926 2436 927 2440
rect 931 2436 932 2440
rect 926 2435 932 2436
rect 1240 2435 1242 2442
rect 1279 2441 1283 2442
rect 1359 2446 1363 2447
rect 1359 2441 1363 2442
rect 1399 2446 1403 2447
rect 1399 2441 1403 2442
rect 1455 2446 1459 2447
rect 1455 2441 1459 2442
rect 1519 2446 1523 2447
rect 1519 2441 1523 2442
rect 1535 2446 1539 2447
rect 1535 2441 1539 2442
rect 1575 2446 1579 2447
rect 1575 2441 1579 2442
rect 1599 2446 1603 2447
rect 1599 2441 1603 2442
rect 1615 2446 1619 2447
rect 1615 2441 1619 2442
rect 1655 2446 1659 2447
rect 1655 2441 1659 2442
rect 1679 2446 1683 2447
rect 1679 2441 1683 2442
rect 1695 2446 1699 2447
rect 1695 2441 1699 2442
rect 1735 2446 1739 2447
rect 1735 2441 1739 2442
rect 1759 2446 1763 2447
rect 1759 2441 1763 2442
rect 1775 2446 1779 2447
rect 1775 2441 1779 2442
rect 1815 2446 1819 2447
rect 1815 2441 1819 2442
rect 1839 2446 1843 2447
rect 1839 2441 1843 2442
rect 1855 2446 1859 2447
rect 1855 2441 1859 2442
rect 1895 2446 1899 2447
rect 1895 2441 1899 2442
rect 1919 2446 1923 2447
rect 1919 2441 1923 2442
rect 1935 2446 1939 2447
rect 1935 2441 1939 2442
rect 1975 2446 1979 2447
rect 1975 2441 1979 2442
rect 1999 2446 2003 2447
rect 1999 2441 2003 2442
rect 2079 2446 2083 2447
rect 2079 2441 2083 2442
rect 2159 2446 2163 2447
rect 2159 2441 2163 2442
rect 2247 2446 2251 2447
rect 2247 2441 2251 2442
rect 2335 2446 2339 2447
rect 2335 2441 2339 2442
rect 2407 2446 2411 2447
rect 2407 2441 2411 2442
rect 111 2434 115 2435
rect 111 2429 115 2430
rect 135 2434 139 2435
rect 135 2429 139 2430
rect 175 2434 179 2435
rect 175 2429 179 2430
rect 183 2434 187 2435
rect 183 2429 187 2430
rect 215 2434 219 2435
rect 215 2429 219 2430
rect 247 2434 251 2435
rect 247 2429 251 2430
rect 255 2434 259 2435
rect 255 2429 259 2430
rect 311 2434 315 2435
rect 311 2429 315 2430
rect 319 2434 323 2435
rect 319 2429 323 2430
rect 391 2434 395 2435
rect 391 2429 395 2430
rect 471 2434 475 2435
rect 471 2429 475 2430
rect 479 2434 483 2435
rect 479 2429 483 2430
rect 543 2434 547 2435
rect 543 2429 547 2430
rect 567 2434 571 2435
rect 567 2429 571 2430
rect 615 2434 619 2435
rect 615 2429 619 2430
rect 655 2434 659 2435
rect 655 2429 659 2430
rect 679 2434 683 2435
rect 679 2429 683 2430
rect 735 2434 739 2435
rect 735 2429 739 2430
rect 743 2434 747 2435
rect 743 2429 747 2430
rect 791 2434 795 2435
rect 791 2429 795 2430
rect 831 2434 835 2435
rect 831 2429 835 2430
rect 839 2434 843 2435
rect 839 2429 843 2430
rect 887 2434 891 2435
rect 887 2429 891 2430
rect 927 2434 931 2435
rect 927 2429 931 2430
rect 935 2434 939 2435
rect 935 2429 939 2430
rect 991 2434 995 2435
rect 991 2429 995 2430
rect 1047 2434 1051 2435
rect 1047 2429 1051 2430
rect 1239 2434 1243 2435
rect 1239 2429 1243 2430
rect 112 2422 114 2429
rect 134 2428 140 2429
rect 134 2424 135 2428
rect 139 2424 140 2428
rect 134 2423 140 2424
rect 182 2428 188 2429
rect 182 2424 183 2428
rect 187 2424 188 2428
rect 182 2423 188 2424
rect 246 2428 252 2429
rect 246 2424 247 2428
rect 251 2424 252 2428
rect 246 2423 252 2424
rect 318 2428 324 2429
rect 318 2424 319 2428
rect 323 2424 324 2428
rect 318 2423 324 2424
rect 390 2428 396 2429
rect 390 2424 391 2428
rect 395 2424 396 2428
rect 390 2423 396 2424
rect 470 2428 476 2429
rect 470 2424 471 2428
rect 475 2424 476 2428
rect 470 2423 476 2424
rect 542 2428 548 2429
rect 542 2424 543 2428
rect 547 2424 548 2428
rect 542 2423 548 2424
rect 614 2428 620 2429
rect 614 2424 615 2428
rect 619 2424 620 2428
rect 614 2423 620 2424
rect 678 2428 684 2429
rect 678 2424 679 2428
rect 683 2424 684 2428
rect 678 2423 684 2424
rect 734 2428 740 2429
rect 734 2424 735 2428
rect 739 2424 740 2428
rect 734 2423 740 2424
rect 790 2428 796 2429
rect 790 2424 791 2428
rect 795 2424 796 2428
rect 790 2423 796 2424
rect 838 2428 844 2429
rect 838 2424 839 2428
rect 843 2424 844 2428
rect 838 2423 844 2424
rect 886 2428 892 2429
rect 886 2424 887 2428
rect 891 2424 892 2428
rect 886 2423 892 2424
rect 934 2428 940 2429
rect 934 2424 935 2428
rect 939 2424 940 2428
rect 934 2423 940 2424
rect 990 2428 996 2429
rect 990 2424 991 2428
rect 995 2424 996 2428
rect 990 2423 996 2424
rect 1046 2428 1052 2429
rect 1046 2424 1047 2428
rect 1051 2424 1052 2428
rect 1046 2423 1052 2424
rect 1240 2422 1242 2429
rect 110 2421 116 2422
rect 110 2417 111 2421
rect 115 2417 116 2421
rect 110 2416 116 2417
rect 1238 2421 1244 2422
rect 1238 2417 1239 2421
rect 1243 2417 1244 2421
rect 1238 2416 1244 2417
rect 1280 2409 1282 2441
rect 1360 2432 1362 2441
rect 1400 2432 1402 2441
rect 1456 2432 1458 2441
rect 1520 2432 1522 2441
rect 1600 2432 1602 2441
rect 1680 2432 1682 2441
rect 1760 2432 1762 2441
rect 1840 2432 1842 2441
rect 1920 2432 1922 2441
rect 2000 2432 2002 2441
rect 2080 2432 2082 2441
rect 2160 2432 2162 2441
rect 2248 2432 2250 2441
rect 2336 2432 2338 2441
rect 1358 2431 1364 2432
rect 1358 2427 1359 2431
rect 1363 2427 1364 2431
rect 1358 2426 1364 2427
rect 1398 2431 1404 2432
rect 1398 2427 1399 2431
rect 1403 2427 1404 2431
rect 1398 2426 1404 2427
rect 1454 2431 1460 2432
rect 1454 2427 1455 2431
rect 1459 2427 1460 2431
rect 1454 2426 1460 2427
rect 1518 2431 1524 2432
rect 1518 2427 1519 2431
rect 1523 2427 1524 2431
rect 1518 2426 1524 2427
rect 1598 2431 1604 2432
rect 1598 2427 1599 2431
rect 1603 2427 1604 2431
rect 1598 2426 1604 2427
rect 1678 2431 1684 2432
rect 1678 2427 1679 2431
rect 1683 2427 1684 2431
rect 1678 2426 1684 2427
rect 1758 2431 1764 2432
rect 1758 2427 1759 2431
rect 1763 2427 1764 2431
rect 1758 2426 1764 2427
rect 1838 2431 1844 2432
rect 1838 2427 1839 2431
rect 1843 2427 1844 2431
rect 1838 2426 1844 2427
rect 1918 2431 1924 2432
rect 1918 2427 1919 2431
rect 1923 2427 1924 2431
rect 1918 2426 1924 2427
rect 1998 2431 2004 2432
rect 1998 2427 1999 2431
rect 2003 2427 2004 2431
rect 1998 2426 2004 2427
rect 2078 2431 2084 2432
rect 2078 2427 2079 2431
rect 2083 2427 2084 2431
rect 2078 2426 2084 2427
rect 2158 2431 2164 2432
rect 2158 2427 2159 2431
rect 2163 2427 2164 2431
rect 2158 2426 2164 2427
rect 2246 2431 2252 2432
rect 2246 2427 2247 2431
rect 2251 2427 2252 2431
rect 2246 2426 2252 2427
rect 2334 2431 2340 2432
rect 2334 2427 2335 2431
rect 2339 2427 2340 2431
rect 2334 2426 2340 2427
rect 2408 2409 2410 2441
rect 1278 2408 1284 2409
rect 110 2404 116 2405
rect 110 2400 111 2404
rect 115 2400 116 2404
rect 110 2399 116 2400
rect 1238 2404 1244 2405
rect 1238 2400 1239 2404
rect 1243 2400 1244 2404
rect 1278 2404 1279 2408
rect 1283 2404 1284 2408
rect 1278 2403 1284 2404
rect 2406 2408 2412 2409
rect 2406 2404 2407 2408
rect 2411 2404 2412 2408
rect 2406 2403 2412 2404
rect 1238 2399 1244 2400
rect 112 2359 114 2399
rect 134 2381 140 2382
rect 134 2377 135 2381
rect 139 2377 140 2381
rect 134 2376 140 2377
rect 182 2381 188 2382
rect 182 2377 183 2381
rect 187 2377 188 2381
rect 182 2376 188 2377
rect 246 2381 252 2382
rect 246 2377 247 2381
rect 251 2377 252 2381
rect 246 2376 252 2377
rect 318 2381 324 2382
rect 318 2377 319 2381
rect 323 2377 324 2381
rect 318 2376 324 2377
rect 390 2381 396 2382
rect 390 2377 391 2381
rect 395 2377 396 2381
rect 390 2376 396 2377
rect 470 2381 476 2382
rect 470 2377 471 2381
rect 475 2377 476 2381
rect 470 2376 476 2377
rect 542 2381 548 2382
rect 542 2377 543 2381
rect 547 2377 548 2381
rect 542 2376 548 2377
rect 614 2381 620 2382
rect 614 2377 615 2381
rect 619 2377 620 2381
rect 614 2376 620 2377
rect 678 2381 684 2382
rect 678 2377 679 2381
rect 683 2377 684 2381
rect 678 2376 684 2377
rect 734 2381 740 2382
rect 734 2377 735 2381
rect 739 2377 740 2381
rect 734 2376 740 2377
rect 790 2381 796 2382
rect 790 2377 791 2381
rect 795 2377 796 2381
rect 790 2376 796 2377
rect 838 2381 844 2382
rect 838 2377 839 2381
rect 843 2377 844 2381
rect 838 2376 844 2377
rect 886 2381 892 2382
rect 886 2377 887 2381
rect 891 2377 892 2381
rect 886 2376 892 2377
rect 934 2381 940 2382
rect 934 2377 935 2381
rect 939 2377 940 2381
rect 934 2376 940 2377
rect 990 2381 996 2382
rect 990 2377 991 2381
rect 995 2377 996 2381
rect 990 2376 996 2377
rect 1046 2381 1052 2382
rect 1046 2377 1047 2381
rect 1051 2377 1052 2381
rect 1046 2376 1052 2377
rect 136 2359 138 2376
rect 184 2359 186 2376
rect 248 2359 250 2376
rect 320 2359 322 2376
rect 392 2359 394 2376
rect 472 2359 474 2376
rect 544 2359 546 2376
rect 616 2359 618 2376
rect 680 2359 682 2376
rect 736 2359 738 2376
rect 792 2359 794 2376
rect 840 2359 842 2376
rect 888 2359 890 2376
rect 936 2359 938 2376
rect 992 2359 994 2376
rect 1048 2359 1050 2376
rect 1240 2359 1242 2399
rect 1278 2391 1284 2392
rect 1278 2387 1279 2391
rect 1283 2387 1284 2391
rect 1278 2386 1284 2387
rect 2406 2391 2412 2392
rect 2406 2387 2407 2391
rect 2411 2387 2412 2391
rect 2406 2386 2412 2387
rect 1280 2379 1282 2386
rect 1358 2384 1364 2385
rect 1358 2380 1359 2384
rect 1363 2380 1364 2384
rect 1358 2379 1364 2380
rect 1398 2384 1404 2385
rect 1398 2380 1399 2384
rect 1403 2380 1404 2384
rect 1398 2379 1404 2380
rect 1454 2384 1460 2385
rect 1454 2380 1455 2384
rect 1459 2380 1460 2384
rect 1454 2379 1460 2380
rect 1518 2384 1524 2385
rect 1518 2380 1519 2384
rect 1523 2380 1524 2384
rect 1518 2379 1524 2380
rect 1598 2384 1604 2385
rect 1598 2380 1599 2384
rect 1603 2380 1604 2384
rect 1598 2379 1604 2380
rect 1678 2384 1684 2385
rect 1678 2380 1679 2384
rect 1683 2380 1684 2384
rect 1678 2379 1684 2380
rect 1758 2384 1764 2385
rect 1758 2380 1759 2384
rect 1763 2380 1764 2384
rect 1758 2379 1764 2380
rect 1838 2384 1844 2385
rect 1838 2380 1839 2384
rect 1843 2380 1844 2384
rect 1838 2379 1844 2380
rect 1918 2384 1924 2385
rect 1918 2380 1919 2384
rect 1923 2380 1924 2384
rect 1918 2379 1924 2380
rect 1998 2384 2004 2385
rect 1998 2380 1999 2384
rect 2003 2380 2004 2384
rect 1998 2379 2004 2380
rect 2078 2384 2084 2385
rect 2078 2380 2079 2384
rect 2083 2380 2084 2384
rect 2078 2379 2084 2380
rect 2158 2384 2164 2385
rect 2158 2380 2159 2384
rect 2163 2380 2164 2384
rect 2158 2379 2164 2380
rect 2246 2384 2252 2385
rect 2246 2380 2247 2384
rect 2251 2380 2252 2384
rect 2246 2379 2252 2380
rect 2334 2384 2340 2385
rect 2334 2380 2335 2384
rect 2339 2380 2340 2384
rect 2334 2379 2340 2380
rect 2408 2379 2410 2386
rect 1279 2378 1283 2379
rect 1279 2373 1283 2374
rect 1359 2378 1363 2379
rect 1359 2373 1363 2374
rect 1399 2378 1403 2379
rect 1399 2373 1403 2374
rect 1407 2378 1411 2379
rect 1407 2373 1411 2374
rect 1455 2378 1459 2379
rect 1455 2373 1459 2374
rect 1471 2378 1475 2379
rect 1471 2373 1475 2374
rect 1519 2378 1523 2379
rect 1519 2373 1523 2374
rect 1543 2378 1547 2379
rect 1543 2373 1547 2374
rect 1599 2378 1603 2379
rect 1599 2373 1603 2374
rect 1615 2378 1619 2379
rect 1615 2373 1619 2374
rect 1679 2378 1683 2379
rect 1679 2373 1683 2374
rect 1695 2378 1699 2379
rect 1695 2373 1699 2374
rect 1759 2378 1763 2379
rect 1759 2373 1763 2374
rect 1775 2378 1779 2379
rect 1775 2373 1779 2374
rect 1839 2378 1843 2379
rect 1839 2373 1843 2374
rect 1855 2378 1859 2379
rect 1855 2373 1859 2374
rect 1919 2378 1923 2379
rect 1919 2373 1923 2374
rect 1927 2378 1931 2379
rect 1927 2373 1931 2374
rect 1999 2378 2003 2379
rect 1999 2373 2003 2374
rect 2071 2378 2075 2379
rect 2071 2373 2075 2374
rect 2079 2378 2083 2379
rect 2079 2373 2083 2374
rect 2143 2378 2147 2379
rect 2143 2373 2147 2374
rect 2159 2378 2163 2379
rect 2159 2373 2163 2374
rect 2223 2378 2227 2379
rect 2223 2373 2227 2374
rect 2247 2378 2251 2379
rect 2247 2373 2251 2374
rect 2303 2378 2307 2379
rect 2303 2373 2307 2374
rect 2335 2378 2339 2379
rect 2335 2373 2339 2374
rect 2359 2378 2363 2379
rect 2359 2373 2363 2374
rect 2407 2378 2411 2379
rect 2407 2373 2411 2374
rect 1280 2366 1282 2373
rect 1358 2372 1364 2373
rect 1358 2368 1359 2372
rect 1363 2368 1364 2372
rect 1358 2367 1364 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1470 2372 1476 2373
rect 1470 2368 1471 2372
rect 1475 2368 1476 2372
rect 1470 2367 1476 2368
rect 1542 2372 1548 2373
rect 1542 2368 1543 2372
rect 1547 2368 1548 2372
rect 1542 2367 1548 2368
rect 1614 2372 1620 2373
rect 1614 2368 1615 2372
rect 1619 2368 1620 2372
rect 1614 2367 1620 2368
rect 1694 2372 1700 2373
rect 1694 2368 1695 2372
rect 1699 2368 1700 2372
rect 1694 2367 1700 2368
rect 1774 2372 1780 2373
rect 1774 2368 1775 2372
rect 1779 2368 1780 2372
rect 1774 2367 1780 2368
rect 1854 2372 1860 2373
rect 1854 2368 1855 2372
rect 1859 2368 1860 2372
rect 1854 2367 1860 2368
rect 1926 2372 1932 2373
rect 1926 2368 1927 2372
rect 1931 2368 1932 2372
rect 1926 2367 1932 2368
rect 1998 2372 2004 2373
rect 1998 2368 1999 2372
rect 2003 2368 2004 2372
rect 1998 2367 2004 2368
rect 2070 2372 2076 2373
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 2142 2372 2148 2373
rect 2142 2368 2143 2372
rect 2147 2368 2148 2372
rect 2142 2367 2148 2368
rect 2222 2372 2228 2373
rect 2222 2368 2223 2372
rect 2227 2368 2228 2372
rect 2222 2367 2228 2368
rect 2302 2372 2308 2373
rect 2302 2368 2303 2372
rect 2307 2368 2308 2372
rect 2302 2367 2308 2368
rect 2358 2372 2364 2373
rect 2358 2368 2359 2372
rect 2363 2368 2364 2372
rect 2358 2367 2364 2368
rect 2408 2366 2410 2373
rect 1278 2365 1284 2366
rect 1278 2361 1279 2365
rect 1283 2361 1284 2365
rect 1278 2360 1284 2361
rect 2406 2365 2412 2366
rect 2406 2361 2407 2365
rect 2411 2361 2412 2365
rect 2406 2360 2412 2361
rect 111 2358 115 2359
rect 111 2353 115 2354
rect 135 2358 139 2359
rect 135 2353 139 2354
rect 175 2358 179 2359
rect 175 2353 179 2354
rect 183 2358 187 2359
rect 183 2353 187 2354
rect 215 2358 219 2359
rect 215 2353 219 2354
rect 247 2358 251 2359
rect 247 2353 251 2354
rect 271 2358 275 2359
rect 271 2353 275 2354
rect 319 2358 323 2359
rect 319 2353 323 2354
rect 351 2358 355 2359
rect 351 2353 355 2354
rect 391 2358 395 2359
rect 391 2353 395 2354
rect 431 2358 435 2359
rect 431 2353 435 2354
rect 471 2358 475 2359
rect 471 2353 475 2354
rect 519 2358 523 2359
rect 519 2353 523 2354
rect 543 2358 547 2359
rect 543 2353 547 2354
rect 599 2358 603 2359
rect 599 2353 603 2354
rect 615 2358 619 2359
rect 615 2353 619 2354
rect 679 2358 683 2359
rect 679 2353 683 2354
rect 735 2358 739 2359
rect 735 2353 739 2354
rect 751 2358 755 2359
rect 751 2353 755 2354
rect 791 2358 795 2359
rect 791 2353 795 2354
rect 823 2358 827 2359
rect 823 2353 827 2354
rect 839 2358 843 2359
rect 839 2353 843 2354
rect 887 2358 891 2359
rect 887 2353 891 2354
rect 935 2358 939 2359
rect 935 2353 939 2354
rect 959 2358 963 2359
rect 959 2353 963 2354
rect 991 2358 995 2359
rect 991 2353 995 2354
rect 1031 2358 1035 2359
rect 1031 2353 1035 2354
rect 1047 2358 1051 2359
rect 1047 2353 1051 2354
rect 1239 2358 1243 2359
rect 1239 2353 1243 2354
rect 112 2321 114 2353
rect 136 2344 138 2353
rect 176 2344 178 2353
rect 216 2344 218 2353
rect 272 2344 274 2353
rect 352 2344 354 2353
rect 432 2344 434 2353
rect 520 2344 522 2353
rect 600 2344 602 2353
rect 680 2344 682 2353
rect 752 2344 754 2353
rect 824 2344 826 2353
rect 888 2344 890 2353
rect 960 2344 962 2353
rect 1032 2344 1034 2353
rect 134 2343 140 2344
rect 134 2339 135 2343
rect 139 2339 140 2343
rect 134 2338 140 2339
rect 174 2343 180 2344
rect 174 2339 175 2343
rect 179 2339 180 2343
rect 174 2338 180 2339
rect 214 2343 220 2344
rect 214 2339 215 2343
rect 219 2339 220 2343
rect 214 2338 220 2339
rect 270 2343 276 2344
rect 270 2339 271 2343
rect 275 2339 276 2343
rect 270 2338 276 2339
rect 350 2343 356 2344
rect 350 2339 351 2343
rect 355 2339 356 2343
rect 350 2338 356 2339
rect 430 2343 436 2344
rect 430 2339 431 2343
rect 435 2339 436 2343
rect 430 2338 436 2339
rect 518 2343 524 2344
rect 518 2339 519 2343
rect 523 2339 524 2343
rect 518 2338 524 2339
rect 598 2343 604 2344
rect 598 2339 599 2343
rect 603 2339 604 2343
rect 598 2338 604 2339
rect 678 2343 684 2344
rect 678 2339 679 2343
rect 683 2339 684 2343
rect 678 2338 684 2339
rect 750 2343 756 2344
rect 750 2339 751 2343
rect 755 2339 756 2343
rect 750 2338 756 2339
rect 822 2343 828 2344
rect 822 2339 823 2343
rect 827 2339 828 2343
rect 822 2338 828 2339
rect 886 2343 892 2344
rect 886 2339 887 2343
rect 891 2339 892 2343
rect 886 2338 892 2339
rect 958 2343 964 2344
rect 958 2339 959 2343
rect 963 2339 964 2343
rect 958 2338 964 2339
rect 1030 2343 1036 2344
rect 1030 2339 1031 2343
rect 1035 2339 1036 2343
rect 1030 2338 1036 2339
rect 1240 2321 1242 2353
rect 1278 2348 1284 2349
rect 1278 2344 1279 2348
rect 1283 2344 1284 2348
rect 1278 2343 1284 2344
rect 2406 2348 2412 2349
rect 2406 2344 2407 2348
rect 2411 2344 2412 2348
rect 2406 2343 2412 2344
rect 110 2320 116 2321
rect 110 2316 111 2320
rect 115 2316 116 2320
rect 110 2315 116 2316
rect 1238 2320 1244 2321
rect 1238 2316 1239 2320
rect 1243 2316 1244 2320
rect 1238 2315 1244 2316
rect 1280 2307 1282 2343
rect 1358 2325 1364 2326
rect 1358 2321 1359 2325
rect 1363 2321 1364 2325
rect 1358 2320 1364 2321
rect 1406 2325 1412 2326
rect 1406 2321 1407 2325
rect 1411 2321 1412 2325
rect 1406 2320 1412 2321
rect 1470 2325 1476 2326
rect 1470 2321 1471 2325
rect 1475 2321 1476 2325
rect 1470 2320 1476 2321
rect 1542 2325 1548 2326
rect 1542 2321 1543 2325
rect 1547 2321 1548 2325
rect 1542 2320 1548 2321
rect 1614 2325 1620 2326
rect 1614 2321 1615 2325
rect 1619 2321 1620 2325
rect 1614 2320 1620 2321
rect 1694 2325 1700 2326
rect 1694 2321 1695 2325
rect 1699 2321 1700 2325
rect 1694 2320 1700 2321
rect 1774 2325 1780 2326
rect 1774 2321 1775 2325
rect 1779 2321 1780 2325
rect 1774 2320 1780 2321
rect 1854 2325 1860 2326
rect 1854 2321 1855 2325
rect 1859 2321 1860 2325
rect 1854 2320 1860 2321
rect 1926 2325 1932 2326
rect 1926 2321 1927 2325
rect 1931 2321 1932 2325
rect 1926 2320 1932 2321
rect 1998 2325 2004 2326
rect 1998 2321 1999 2325
rect 2003 2321 2004 2325
rect 1998 2320 2004 2321
rect 2070 2325 2076 2326
rect 2070 2321 2071 2325
rect 2075 2321 2076 2325
rect 2070 2320 2076 2321
rect 2142 2325 2148 2326
rect 2142 2321 2143 2325
rect 2147 2321 2148 2325
rect 2142 2320 2148 2321
rect 2222 2325 2228 2326
rect 2222 2321 2223 2325
rect 2227 2321 2228 2325
rect 2222 2320 2228 2321
rect 2302 2325 2308 2326
rect 2302 2321 2303 2325
rect 2307 2321 2308 2325
rect 2302 2320 2308 2321
rect 2358 2325 2364 2326
rect 2358 2321 2359 2325
rect 2363 2321 2364 2325
rect 2358 2320 2364 2321
rect 1360 2307 1362 2320
rect 1408 2307 1410 2320
rect 1472 2307 1474 2320
rect 1544 2307 1546 2320
rect 1616 2307 1618 2320
rect 1696 2307 1698 2320
rect 1776 2307 1778 2320
rect 1856 2307 1858 2320
rect 1928 2307 1930 2320
rect 2000 2307 2002 2320
rect 2072 2307 2074 2320
rect 2144 2307 2146 2320
rect 2224 2307 2226 2320
rect 2304 2307 2306 2320
rect 2360 2307 2362 2320
rect 2408 2307 2410 2343
rect 1279 2306 1283 2307
rect 110 2303 116 2304
rect 110 2299 111 2303
rect 115 2299 116 2303
rect 110 2298 116 2299
rect 1238 2303 1244 2304
rect 1238 2299 1239 2303
rect 1243 2299 1244 2303
rect 1279 2301 1283 2302
rect 1359 2306 1363 2307
rect 1359 2301 1363 2302
rect 1407 2306 1411 2307
rect 1407 2301 1411 2302
rect 1471 2306 1475 2307
rect 1471 2301 1475 2302
rect 1503 2306 1507 2307
rect 1503 2301 1507 2302
rect 1543 2306 1547 2307
rect 1543 2301 1547 2302
rect 1583 2306 1587 2307
rect 1583 2301 1587 2302
rect 1615 2306 1619 2307
rect 1615 2301 1619 2302
rect 1623 2306 1627 2307
rect 1623 2301 1627 2302
rect 1663 2306 1667 2307
rect 1663 2301 1667 2302
rect 1695 2306 1699 2307
rect 1695 2301 1699 2302
rect 1703 2306 1707 2307
rect 1703 2301 1707 2302
rect 1759 2306 1763 2307
rect 1759 2301 1763 2302
rect 1775 2306 1779 2307
rect 1775 2301 1779 2302
rect 1823 2306 1827 2307
rect 1823 2301 1827 2302
rect 1855 2306 1859 2307
rect 1855 2301 1859 2302
rect 1895 2306 1899 2307
rect 1895 2301 1899 2302
rect 1927 2306 1931 2307
rect 1927 2301 1931 2302
rect 1967 2306 1971 2307
rect 1967 2301 1971 2302
rect 1999 2306 2003 2307
rect 1999 2301 2003 2302
rect 2047 2306 2051 2307
rect 2047 2301 2051 2302
rect 2071 2306 2075 2307
rect 2071 2301 2075 2302
rect 2127 2306 2131 2307
rect 2127 2301 2131 2302
rect 2143 2306 2147 2307
rect 2143 2301 2147 2302
rect 2207 2306 2211 2307
rect 2207 2301 2211 2302
rect 2223 2306 2227 2307
rect 2223 2301 2227 2302
rect 2295 2306 2299 2307
rect 2295 2301 2299 2302
rect 2303 2306 2307 2307
rect 2303 2301 2307 2302
rect 2359 2306 2363 2307
rect 2359 2301 2363 2302
rect 2407 2306 2411 2307
rect 2407 2301 2411 2302
rect 1238 2298 1244 2299
rect 112 2287 114 2298
rect 134 2296 140 2297
rect 134 2292 135 2296
rect 139 2292 140 2296
rect 134 2291 140 2292
rect 174 2296 180 2297
rect 174 2292 175 2296
rect 179 2292 180 2296
rect 174 2291 180 2292
rect 214 2296 220 2297
rect 214 2292 215 2296
rect 219 2292 220 2296
rect 214 2291 220 2292
rect 270 2296 276 2297
rect 270 2292 271 2296
rect 275 2292 276 2296
rect 270 2291 276 2292
rect 350 2296 356 2297
rect 350 2292 351 2296
rect 355 2292 356 2296
rect 350 2291 356 2292
rect 430 2296 436 2297
rect 430 2292 431 2296
rect 435 2292 436 2296
rect 430 2291 436 2292
rect 518 2296 524 2297
rect 518 2292 519 2296
rect 523 2292 524 2296
rect 518 2291 524 2292
rect 598 2296 604 2297
rect 598 2292 599 2296
rect 603 2292 604 2296
rect 598 2291 604 2292
rect 678 2296 684 2297
rect 678 2292 679 2296
rect 683 2292 684 2296
rect 678 2291 684 2292
rect 750 2296 756 2297
rect 750 2292 751 2296
rect 755 2292 756 2296
rect 750 2291 756 2292
rect 822 2296 828 2297
rect 822 2292 823 2296
rect 827 2292 828 2296
rect 822 2291 828 2292
rect 886 2296 892 2297
rect 886 2292 887 2296
rect 891 2292 892 2296
rect 886 2291 892 2292
rect 958 2296 964 2297
rect 958 2292 959 2296
rect 963 2292 964 2296
rect 958 2291 964 2292
rect 1030 2296 1036 2297
rect 1030 2292 1031 2296
rect 1035 2292 1036 2296
rect 1030 2291 1036 2292
rect 136 2287 138 2291
rect 176 2287 178 2291
rect 216 2287 218 2291
rect 272 2287 274 2291
rect 352 2287 354 2291
rect 432 2287 434 2291
rect 520 2287 522 2291
rect 600 2287 602 2291
rect 680 2287 682 2291
rect 752 2287 754 2291
rect 824 2287 826 2291
rect 888 2287 890 2291
rect 960 2287 962 2291
rect 1032 2287 1034 2291
rect 1240 2287 1242 2298
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 135 2286 139 2287
rect 135 2281 139 2282
rect 175 2286 179 2287
rect 175 2281 179 2282
rect 215 2286 219 2287
rect 215 2281 219 2282
rect 231 2286 235 2287
rect 231 2281 235 2282
rect 271 2286 275 2287
rect 271 2281 275 2282
rect 303 2286 307 2287
rect 303 2281 307 2282
rect 351 2286 355 2287
rect 351 2281 355 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 431 2286 435 2287
rect 431 2281 435 2282
rect 455 2286 459 2287
rect 455 2281 459 2282
rect 519 2286 523 2287
rect 519 2281 523 2282
rect 535 2286 539 2287
rect 535 2281 539 2282
rect 599 2286 603 2287
rect 599 2281 603 2282
rect 615 2286 619 2287
rect 615 2281 619 2282
rect 679 2286 683 2287
rect 679 2281 683 2282
rect 687 2286 691 2287
rect 687 2281 691 2282
rect 751 2286 755 2287
rect 751 2281 755 2282
rect 759 2286 763 2287
rect 759 2281 763 2282
rect 823 2286 827 2287
rect 823 2281 827 2282
rect 831 2286 835 2287
rect 831 2281 835 2282
rect 887 2286 891 2287
rect 887 2281 891 2282
rect 911 2286 915 2287
rect 911 2281 915 2282
rect 959 2286 963 2287
rect 959 2281 963 2282
rect 991 2286 995 2287
rect 991 2281 995 2282
rect 1031 2286 1035 2287
rect 1031 2281 1035 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 112 2274 114 2281
rect 134 2280 140 2281
rect 134 2276 135 2280
rect 139 2276 140 2280
rect 134 2275 140 2276
rect 174 2280 180 2281
rect 174 2276 175 2280
rect 179 2276 180 2280
rect 174 2275 180 2276
rect 230 2280 236 2281
rect 230 2276 231 2280
rect 235 2276 236 2280
rect 230 2275 236 2276
rect 302 2280 308 2281
rect 302 2276 303 2280
rect 307 2276 308 2280
rect 302 2275 308 2276
rect 374 2280 380 2281
rect 374 2276 375 2280
rect 379 2276 380 2280
rect 374 2275 380 2276
rect 454 2280 460 2281
rect 454 2276 455 2280
rect 459 2276 460 2280
rect 454 2275 460 2276
rect 534 2280 540 2281
rect 534 2276 535 2280
rect 539 2276 540 2280
rect 534 2275 540 2276
rect 614 2280 620 2281
rect 614 2276 615 2280
rect 619 2276 620 2280
rect 614 2275 620 2276
rect 686 2280 692 2281
rect 686 2276 687 2280
rect 691 2276 692 2280
rect 686 2275 692 2276
rect 758 2280 764 2281
rect 758 2276 759 2280
rect 763 2276 764 2280
rect 758 2275 764 2276
rect 830 2280 836 2281
rect 830 2276 831 2280
rect 835 2276 836 2280
rect 830 2275 836 2276
rect 910 2280 916 2281
rect 910 2276 911 2280
rect 915 2276 916 2280
rect 910 2275 916 2276
rect 990 2280 996 2281
rect 990 2276 991 2280
rect 995 2276 996 2280
rect 990 2275 996 2276
rect 1240 2274 1242 2281
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 110 2268 116 2269
rect 1238 2273 1244 2274
rect 1238 2269 1239 2273
rect 1243 2269 1244 2273
rect 1280 2269 1282 2301
rect 1504 2292 1506 2301
rect 1544 2292 1546 2301
rect 1584 2292 1586 2301
rect 1624 2292 1626 2301
rect 1664 2292 1666 2301
rect 1704 2292 1706 2301
rect 1760 2292 1762 2301
rect 1824 2292 1826 2301
rect 1896 2292 1898 2301
rect 1968 2292 1970 2301
rect 2048 2292 2050 2301
rect 2128 2292 2130 2301
rect 2208 2292 2210 2301
rect 2296 2292 2298 2301
rect 2360 2292 2362 2301
rect 1502 2291 1508 2292
rect 1502 2287 1503 2291
rect 1507 2287 1508 2291
rect 1502 2286 1508 2287
rect 1542 2291 1548 2292
rect 1542 2287 1543 2291
rect 1547 2287 1548 2291
rect 1542 2286 1548 2287
rect 1582 2291 1588 2292
rect 1582 2287 1583 2291
rect 1587 2287 1588 2291
rect 1582 2286 1588 2287
rect 1622 2291 1628 2292
rect 1622 2287 1623 2291
rect 1627 2287 1628 2291
rect 1622 2286 1628 2287
rect 1662 2291 1668 2292
rect 1662 2287 1663 2291
rect 1667 2287 1668 2291
rect 1662 2286 1668 2287
rect 1702 2291 1708 2292
rect 1702 2287 1703 2291
rect 1707 2287 1708 2291
rect 1702 2286 1708 2287
rect 1758 2291 1764 2292
rect 1758 2287 1759 2291
rect 1763 2287 1764 2291
rect 1758 2286 1764 2287
rect 1822 2291 1828 2292
rect 1822 2287 1823 2291
rect 1827 2287 1828 2291
rect 1822 2286 1828 2287
rect 1894 2291 1900 2292
rect 1894 2287 1895 2291
rect 1899 2287 1900 2291
rect 1894 2286 1900 2287
rect 1966 2291 1972 2292
rect 1966 2287 1967 2291
rect 1971 2287 1972 2291
rect 1966 2286 1972 2287
rect 2046 2291 2052 2292
rect 2046 2287 2047 2291
rect 2051 2287 2052 2291
rect 2046 2286 2052 2287
rect 2126 2291 2132 2292
rect 2126 2287 2127 2291
rect 2131 2287 2132 2291
rect 2126 2286 2132 2287
rect 2206 2291 2212 2292
rect 2206 2287 2207 2291
rect 2211 2287 2212 2291
rect 2206 2286 2212 2287
rect 2294 2291 2300 2292
rect 2294 2287 2295 2291
rect 2299 2287 2300 2291
rect 2294 2286 2300 2287
rect 2358 2291 2364 2292
rect 2358 2287 2359 2291
rect 2363 2287 2364 2291
rect 2358 2286 2364 2287
rect 2408 2269 2410 2301
rect 1238 2268 1244 2269
rect 1278 2268 1284 2269
rect 1278 2264 1279 2268
rect 1283 2264 1284 2268
rect 1278 2263 1284 2264
rect 2406 2268 2412 2269
rect 2406 2264 2407 2268
rect 2411 2264 2412 2268
rect 2406 2263 2412 2264
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 110 2251 116 2252
rect 1238 2256 1244 2257
rect 1238 2252 1239 2256
rect 1243 2252 1244 2256
rect 1238 2251 1244 2252
rect 1278 2251 1284 2252
rect 112 2219 114 2251
rect 134 2233 140 2234
rect 134 2229 135 2233
rect 139 2229 140 2233
rect 134 2228 140 2229
rect 174 2233 180 2234
rect 174 2229 175 2233
rect 179 2229 180 2233
rect 174 2228 180 2229
rect 230 2233 236 2234
rect 230 2229 231 2233
rect 235 2229 236 2233
rect 230 2228 236 2229
rect 302 2233 308 2234
rect 302 2229 303 2233
rect 307 2229 308 2233
rect 302 2228 308 2229
rect 374 2233 380 2234
rect 374 2229 375 2233
rect 379 2229 380 2233
rect 374 2228 380 2229
rect 454 2233 460 2234
rect 454 2229 455 2233
rect 459 2229 460 2233
rect 454 2228 460 2229
rect 534 2233 540 2234
rect 534 2229 535 2233
rect 539 2229 540 2233
rect 534 2228 540 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 686 2233 692 2234
rect 686 2229 687 2233
rect 691 2229 692 2233
rect 686 2228 692 2229
rect 758 2233 764 2234
rect 758 2229 759 2233
rect 763 2229 764 2233
rect 758 2228 764 2229
rect 830 2233 836 2234
rect 830 2229 831 2233
rect 835 2229 836 2233
rect 830 2228 836 2229
rect 910 2233 916 2234
rect 910 2229 911 2233
rect 915 2229 916 2233
rect 910 2228 916 2229
rect 990 2233 996 2234
rect 990 2229 991 2233
rect 995 2229 996 2233
rect 990 2228 996 2229
rect 136 2219 138 2228
rect 176 2219 178 2228
rect 232 2219 234 2228
rect 304 2219 306 2228
rect 376 2219 378 2228
rect 456 2219 458 2228
rect 536 2219 538 2228
rect 616 2219 618 2228
rect 688 2219 690 2228
rect 760 2219 762 2228
rect 832 2219 834 2228
rect 912 2219 914 2228
rect 992 2219 994 2228
rect 1240 2219 1242 2251
rect 1278 2247 1279 2251
rect 1283 2247 1284 2251
rect 1278 2246 1284 2247
rect 2406 2251 2412 2252
rect 2406 2247 2407 2251
rect 2411 2247 2412 2251
rect 2406 2246 2412 2247
rect 1280 2231 1282 2246
rect 1502 2244 1508 2245
rect 1502 2240 1503 2244
rect 1507 2240 1508 2244
rect 1502 2239 1508 2240
rect 1542 2244 1548 2245
rect 1542 2240 1543 2244
rect 1547 2240 1548 2244
rect 1542 2239 1548 2240
rect 1582 2244 1588 2245
rect 1582 2240 1583 2244
rect 1587 2240 1588 2244
rect 1582 2239 1588 2240
rect 1622 2244 1628 2245
rect 1622 2240 1623 2244
rect 1627 2240 1628 2244
rect 1622 2239 1628 2240
rect 1662 2244 1668 2245
rect 1662 2240 1663 2244
rect 1667 2240 1668 2244
rect 1662 2239 1668 2240
rect 1702 2244 1708 2245
rect 1702 2240 1703 2244
rect 1707 2240 1708 2244
rect 1702 2239 1708 2240
rect 1758 2244 1764 2245
rect 1758 2240 1759 2244
rect 1763 2240 1764 2244
rect 1758 2239 1764 2240
rect 1822 2244 1828 2245
rect 1822 2240 1823 2244
rect 1827 2240 1828 2244
rect 1822 2239 1828 2240
rect 1894 2244 1900 2245
rect 1894 2240 1895 2244
rect 1899 2240 1900 2244
rect 1894 2239 1900 2240
rect 1966 2244 1972 2245
rect 1966 2240 1967 2244
rect 1971 2240 1972 2244
rect 1966 2239 1972 2240
rect 2046 2244 2052 2245
rect 2046 2240 2047 2244
rect 2051 2240 2052 2244
rect 2046 2239 2052 2240
rect 2126 2244 2132 2245
rect 2126 2240 2127 2244
rect 2131 2240 2132 2244
rect 2126 2239 2132 2240
rect 2206 2244 2212 2245
rect 2206 2240 2207 2244
rect 2211 2240 2212 2244
rect 2206 2239 2212 2240
rect 2294 2244 2300 2245
rect 2294 2240 2295 2244
rect 2299 2240 2300 2244
rect 2294 2239 2300 2240
rect 2358 2244 2364 2245
rect 2358 2240 2359 2244
rect 2363 2240 2364 2244
rect 2358 2239 2364 2240
rect 1504 2231 1506 2239
rect 1544 2231 1546 2239
rect 1584 2231 1586 2239
rect 1624 2231 1626 2239
rect 1664 2231 1666 2239
rect 1704 2231 1706 2239
rect 1760 2231 1762 2239
rect 1824 2231 1826 2239
rect 1896 2231 1898 2239
rect 1968 2231 1970 2239
rect 2048 2231 2050 2239
rect 2128 2231 2130 2239
rect 2208 2231 2210 2239
rect 2296 2231 2298 2239
rect 2360 2231 2362 2239
rect 2408 2231 2410 2246
rect 1279 2230 1283 2231
rect 1279 2225 1283 2226
rect 1303 2230 1307 2231
rect 1303 2225 1307 2226
rect 1343 2230 1347 2231
rect 1343 2225 1347 2226
rect 1383 2230 1387 2231
rect 1383 2225 1387 2226
rect 1431 2230 1435 2231
rect 1431 2225 1435 2226
rect 1495 2230 1499 2231
rect 1495 2225 1499 2226
rect 1503 2230 1507 2231
rect 1503 2225 1507 2226
rect 1543 2230 1547 2231
rect 1543 2225 1547 2226
rect 1567 2230 1571 2231
rect 1567 2225 1571 2226
rect 1583 2230 1587 2231
rect 1583 2225 1587 2226
rect 1623 2230 1627 2231
rect 1623 2225 1627 2226
rect 1639 2230 1643 2231
rect 1639 2225 1643 2226
rect 1663 2230 1667 2231
rect 1663 2225 1667 2226
rect 1703 2230 1707 2231
rect 1703 2225 1707 2226
rect 1711 2230 1715 2231
rect 1711 2225 1715 2226
rect 1759 2230 1763 2231
rect 1759 2225 1763 2226
rect 1783 2230 1787 2231
rect 1783 2225 1787 2226
rect 1823 2230 1827 2231
rect 1823 2225 1827 2226
rect 1855 2230 1859 2231
rect 1855 2225 1859 2226
rect 1895 2230 1899 2231
rect 1895 2225 1899 2226
rect 1935 2230 1939 2231
rect 1935 2225 1939 2226
rect 1967 2230 1971 2231
rect 1967 2225 1971 2226
rect 2015 2230 2019 2231
rect 2015 2225 2019 2226
rect 2047 2230 2051 2231
rect 2047 2225 2051 2226
rect 2095 2230 2099 2231
rect 2095 2225 2099 2226
rect 2127 2230 2131 2231
rect 2127 2225 2131 2226
rect 2183 2230 2187 2231
rect 2183 2225 2187 2226
rect 2207 2230 2211 2231
rect 2207 2225 2211 2226
rect 2279 2230 2283 2231
rect 2279 2225 2283 2226
rect 2295 2230 2299 2231
rect 2295 2225 2299 2226
rect 2359 2230 2363 2231
rect 2359 2225 2363 2226
rect 2407 2230 2411 2231
rect 2407 2225 2411 2226
rect 111 2218 115 2219
rect 111 2213 115 2214
rect 135 2218 139 2219
rect 135 2213 139 2214
rect 175 2218 179 2219
rect 175 2213 179 2214
rect 231 2218 235 2219
rect 231 2213 235 2214
rect 247 2218 251 2219
rect 247 2213 251 2214
rect 287 2218 291 2219
rect 287 2213 291 2214
rect 303 2218 307 2219
rect 303 2213 307 2214
rect 327 2218 331 2219
rect 327 2213 331 2214
rect 375 2218 379 2219
rect 375 2213 379 2214
rect 431 2218 435 2219
rect 431 2213 435 2214
rect 455 2218 459 2219
rect 455 2213 459 2214
rect 495 2218 499 2219
rect 495 2213 499 2214
rect 535 2218 539 2219
rect 535 2213 539 2214
rect 551 2218 555 2219
rect 551 2213 555 2214
rect 607 2218 611 2219
rect 607 2213 611 2214
rect 615 2218 619 2219
rect 615 2213 619 2214
rect 663 2218 667 2219
rect 663 2213 667 2214
rect 687 2218 691 2219
rect 687 2213 691 2214
rect 719 2218 723 2219
rect 719 2213 723 2214
rect 759 2218 763 2219
rect 759 2213 763 2214
rect 783 2218 787 2219
rect 783 2213 787 2214
rect 831 2218 835 2219
rect 831 2213 835 2214
rect 847 2218 851 2219
rect 847 2213 851 2214
rect 911 2218 915 2219
rect 911 2213 915 2214
rect 991 2218 995 2219
rect 991 2213 995 2214
rect 1239 2218 1243 2219
rect 1280 2218 1282 2225
rect 1302 2224 1308 2225
rect 1302 2220 1303 2224
rect 1307 2220 1308 2224
rect 1302 2219 1308 2220
rect 1342 2224 1348 2225
rect 1342 2220 1343 2224
rect 1347 2220 1348 2224
rect 1342 2219 1348 2220
rect 1382 2224 1388 2225
rect 1382 2220 1383 2224
rect 1387 2220 1388 2224
rect 1382 2219 1388 2220
rect 1430 2224 1436 2225
rect 1430 2220 1431 2224
rect 1435 2220 1436 2224
rect 1430 2219 1436 2220
rect 1494 2224 1500 2225
rect 1494 2220 1495 2224
rect 1499 2220 1500 2224
rect 1494 2219 1500 2220
rect 1566 2224 1572 2225
rect 1566 2220 1567 2224
rect 1571 2220 1572 2224
rect 1566 2219 1572 2220
rect 1638 2224 1644 2225
rect 1638 2220 1639 2224
rect 1643 2220 1644 2224
rect 1638 2219 1644 2220
rect 1710 2224 1716 2225
rect 1710 2220 1711 2224
rect 1715 2220 1716 2224
rect 1710 2219 1716 2220
rect 1782 2224 1788 2225
rect 1782 2220 1783 2224
rect 1787 2220 1788 2224
rect 1782 2219 1788 2220
rect 1854 2224 1860 2225
rect 1854 2220 1855 2224
rect 1859 2220 1860 2224
rect 1854 2219 1860 2220
rect 1934 2224 1940 2225
rect 1934 2220 1935 2224
rect 1939 2220 1940 2224
rect 1934 2219 1940 2220
rect 2014 2224 2020 2225
rect 2014 2220 2015 2224
rect 2019 2220 2020 2224
rect 2014 2219 2020 2220
rect 2094 2224 2100 2225
rect 2094 2220 2095 2224
rect 2099 2220 2100 2224
rect 2094 2219 2100 2220
rect 2182 2224 2188 2225
rect 2182 2220 2183 2224
rect 2187 2220 2188 2224
rect 2182 2219 2188 2220
rect 2278 2224 2284 2225
rect 2278 2220 2279 2224
rect 2283 2220 2284 2224
rect 2278 2219 2284 2220
rect 2358 2224 2364 2225
rect 2358 2220 2359 2224
rect 2363 2220 2364 2224
rect 2358 2219 2364 2220
rect 2408 2218 2410 2225
rect 1239 2213 1243 2214
rect 1278 2217 1284 2218
rect 1278 2213 1279 2217
rect 1283 2213 1284 2217
rect 112 2181 114 2213
rect 248 2204 250 2213
rect 288 2204 290 2213
rect 328 2204 330 2213
rect 376 2204 378 2213
rect 432 2204 434 2213
rect 496 2204 498 2213
rect 552 2204 554 2213
rect 608 2204 610 2213
rect 664 2204 666 2213
rect 720 2204 722 2213
rect 784 2204 786 2213
rect 848 2204 850 2213
rect 912 2204 914 2213
rect 246 2203 252 2204
rect 246 2199 247 2203
rect 251 2199 252 2203
rect 246 2198 252 2199
rect 286 2203 292 2204
rect 286 2199 287 2203
rect 291 2199 292 2203
rect 286 2198 292 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 374 2203 380 2204
rect 374 2199 375 2203
rect 379 2199 380 2203
rect 374 2198 380 2199
rect 430 2203 436 2204
rect 430 2199 431 2203
rect 435 2199 436 2203
rect 430 2198 436 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 550 2203 556 2204
rect 550 2199 551 2203
rect 555 2199 556 2203
rect 550 2198 556 2199
rect 606 2203 612 2204
rect 606 2199 607 2203
rect 611 2199 612 2203
rect 606 2198 612 2199
rect 662 2203 668 2204
rect 662 2199 663 2203
rect 667 2199 668 2203
rect 662 2198 668 2199
rect 718 2203 724 2204
rect 718 2199 719 2203
rect 723 2199 724 2203
rect 718 2198 724 2199
rect 782 2203 788 2204
rect 782 2199 783 2203
rect 787 2199 788 2203
rect 782 2198 788 2199
rect 846 2203 852 2204
rect 846 2199 847 2203
rect 851 2199 852 2203
rect 846 2198 852 2199
rect 910 2203 916 2204
rect 910 2199 911 2203
rect 915 2199 916 2203
rect 910 2198 916 2199
rect 1240 2181 1242 2213
rect 1278 2212 1284 2213
rect 2406 2217 2412 2218
rect 2406 2213 2407 2217
rect 2411 2213 2412 2217
rect 2406 2212 2412 2213
rect 1278 2200 1284 2201
rect 1278 2196 1279 2200
rect 1283 2196 1284 2200
rect 1278 2195 1284 2196
rect 2406 2200 2412 2201
rect 2406 2196 2407 2200
rect 2411 2196 2412 2200
rect 2406 2195 2412 2196
rect 110 2180 116 2181
rect 110 2176 111 2180
rect 115 2176 116 2180
rect 110 2175 116 2176
rect 1238 2180 1244 2181
rect 1238 2176 1239 2180
rect 1243 2176 1244 2180
rect 1238 2175 1244 2176
rect 110 2163 116 2164
rect 110 2159 111 2163
rect 115 2159 116 2163
rect 110 2158 116 2159
rect 1238 2163 1244 2164
rect 1280 2163 1282 2195
rect 1302 2177 1308 2178
rect 1302 2173 1303 2177
rect 1307 2173 1308 2177
rect 1302 2172 1308 2173
rect 1342 2177 1348 2178
rect 1342 2173 1343 2177
rect 1347 2173 1348 2177
rect 1342 2172 1348 2173
rect 1382 2177 1388 2178
rect 1382 2173 1383 2177
rect 1387 2173 1388 2177
rect 1382 2172 1388 2173
rect 1430 2177 1436 2178
rect 1430 2173 1431 2177
rect 1435 2173 1436 2177
rect 1430 2172 1436 2173
rect 1494 2177 1500 2178
rect 1494 2173 1495 2177
rect 1499 2173 1500 2177
rect 1494 2172 1500 2173
rect 1566 2177 1572 2178
rect 1566 2173 1567 2177
rect 1571 2173 1572 2177
rect 1566 2172 1572 2173
rect 1638 2177 1644 2178
rect 1638 2173 1639 2177
rect 1643 2173 1644 2177
rect 1638 2172 1644 2173
rect 1710 2177 1716 2178
rect 1710 2173 1711 2177
rect 1715 2173 1716 2177
rect 1710 2172 1716 2173
rect 1782 2177 1788 2178
rect 1782 2173 1783 2177
rect 1787 2173 1788 2177
rect 1782 2172 1788 2173
rect 1854 2177 1860 2178
rect 1854 2173 1855 2177
rect 1859 2173 1860 2177
rect 1854 2172 1860 2173
rect 1934 2177 1940 2178
rect 1934 2173 1935 2177
rect 1939 2173 1940 2177
rect 1934 2172 1940 2173
rect 2014 2177 2020 2178
rect 2014 2173 2015 2177
rect 2019 2173 2020 2177
rect 2014 2172 2020 2173
rect 2094 2177 2100 2178
rect 2094 2173 2095 2177
rect 2099 2173 2100 2177
rect 2094 2172 2100 2173
rect 2182 2177 2188 2178
rect 2182 2173 2183 2177
rect 2187 2173 2188 2177
rect 2182 2172 2188 2173
rect 2278 2177 2284 2178
rect 2278 2173 2279 2177
rect 2283 2173 2284 2177
rect 2278 2172 2284 2173
rect 2358 2177 2364 2178
rect 2358 2173 2359 2177
rect 2363 2173 2364 2177
rect 2358 2172 2364 2173
rect 1304 2163 1306 2172
rect 1344 2163 1346 2172
rect 1384 2163 1386 2172
rect 1432 2163 1434 2172
rect 1496 2163 1498 2172
rect 1568 2163 1570 2172
rect 1640 2163 1642 2172
rect 1712 2163 1714 2172
rect 1784 2163 1786 2172
rect 1856 2163 1858 2172
rect 1936 2163 1938 2172
rect 2016 2163 2018 2172
rect 2096 2163 2098 2172
rect 2184 2163 2186 2172
rect 2280 2163 2282 2172
rect 2360 2163 2362 2172
rect 2408 2163 2410 2195
rect 1238 2159 1239 2163
rect 1243 2159 1244 2163
rect 1238 2158 1244 2159
rect 1279 2162 1283 2163
rect 112 2143 114 2158
rect 246 2156 252 2157
rect 246 2152 247 2156
rect 251 2152 252 2156
rect 246 2151 252 2152
rect 286 2156 292 2157
rect 286 2152 287 2156
rect 291 2152 292 2156
rect 286 2151 292 2152
rect 326 2156 332 2157
rect 326 2152 327 2156
rect 331 2152 332 2156
rect 326 2151 332 2152
rect 374 2156 380 2157
rect 374 2152 375 2156
rect 379 2152 380 2156
rect 374 2151 380 2152
rect 430 2156 436 2157
rect 430 2152 431 2156
rect 435 2152 436 2156
rect 430 2151 436 2152
rect 494 2156 500 2157
rect 494 2152 495 2156
rect 499 2152 500 2156
rect 494 2151 500 2152
rect 550 2156 556 2157
rect 550 2152 551 2156
rect 555 2152 556 2156
rect 550 2151 556 2152
rect 606 2156 612 2157
rect 606 2152 607 2156
rect 611 2152 612 2156
rect 606 2151 612 2152
rect 662 2156 668 2157
rect 662 2152 663 2156
rect 667 2152 668 2156
rect 662 2151 668 2152
rect 718 2156 724 2157
rect 718 2152 719 2156
rect 723 2152 724 2156
rect 718 2151 724 2152
rect 782 2156 788 2157
rect 782 2152 783 2156
rect 787 2152 788 2156
rect 782 2151 788 2152
rect 846 2156 852 2157
rect 846 2152 847 2156
rect 851 2152 852 2156
rect 846 2151 852 2152
rect 910 2156 916 2157
rect 910 2152 911 2156
rect 915 2152 916 2156
rect 910 2151 916 2152
rect 248 2143 250 2151
rect 288 2143 290 2151
rect 328 2143 330 2151
rect 376 2143 378 2151
rect 432 2143 434 2151
rect 496 2143 498 2151
rect 552 2143 554 2151
rect 608 2143 610 2151
rect 664 2143 666 2151
rect 720 2143 722 2151
rect 784 2143 786 2151
rect 848 2143 850 2151
rect 912 2143 914 2151
rect 1240 2143 1242 2158
rect 1279 2157 1283 2158
rect 1303 2162 1307 2163
rect 1303 2157 1307 2158
rect 1343 2162 1347 2163
rect 1343 2157 1347 2158
rect 1351 2162 1355 2163
rect 1351 2157 1355 2158
rect 1383 2162 1387 2163
rect 1383 2157 1387 2158
rect 1431 2162 1435 2163
rect 1431 2157 1435 2158
rect 1439 2162 1443 2163
rect 1439 2157 1443 2158
rect 1495 2162 1499 2163
rect 1495 2157 1499 2158
rect 1535 2162 1539 2163
rect 1535 2157 1539 2158
rect 1567 2162 1571 2163
rect 1567 2157 1571 2158
rect 1631 2162 1635 2163
rect 1631 2157 1635 2158
rect 1639 2162 1643 2163
rect 1639 2157 1643 2158
rect 1711 2162 1715 2163
rect 1711 2157 1715 2158
rect 1727 2162 1731 2163
rect 1727 2157 1731 2158
rect 1783 2162 1787 2163
rect 1783 2157 1787 2158
rect 1815 2162 1819 2163
rect 1815 2157 1819 2158
rect 1855 2162 1859 2163
rect 1855 2157 1859 2158
rect 1895 2162 1899 2163
rect 1895 2157 1899 2158
rect 1935 2162 1939 2163
rect 1935 2157 1939 2158
rect 1975 2162 1979 2163
rect 1975 2157 1979 2158
rect 2015 2162 2019 2163
rect 2015 2157 2019 2158
rect 2047 2162 2051 2163
rect 2047 2157 2051 2158
rect 2095 2162 2099 2163
rect 2095 2157 2099 2158
rect 2111 2162 2115 2163
rect 2111 2157 2115 2158
rect 2175 2162 2179 2163
rect 2175 2157 2179 2158
rect 2183 2162 2187 2163
rect 2183 2157 2187 2158
rect 2239 2162 2243 2163
rect 2239 2157 2243 2158
rect 2279 2162 2283 2163
rect 2279 2157 2283 2158
rect 2311 2162 2315 2163
rect 2311 2157 2315 2158
rect 2359 2162 2363 2163
rect 2359 2157 2363 2158
rect 2407 2162 2411 2163
rect 2407 2157 2411 2158
rect 111 2142 115 2143
rect 111 2137 115 2138
rect 247 2142 251 2143
rect 247 2137 251 2138
rect 287 2142 291 2143
rect 287 2137 291 2138
rect 327 2142 331 2143
rect 327 2137 331 2138
rect 375 2142 379 2143
rect 375 2137 379 2138
rect 383 2142 387 2143
rect 383 2137 387 2138
rect 423 2142 427 2143
rect 423 2137 427 2138
rect 431 2142 435 2143
rect 431 2137 435 2138
rect 463 2142 467 2143
rect 463 2137 467 2138
rect 495 2142 499 2143
rect 495 2137 499 2138
rect 503 2142 507 2143
rect 503 2137 507 2138
rect 551 2142 555 2143
rect 551 2137 555 2138
rect 607 2142 611 2143
rect 607 2137 611 2138
rect 663 2142 667 2143
rect 663 2137 667 2138
rect 719 2142 723 2143
rect 719 2137 723 2138
rect 727 2142 731 2143
rect 727 2137 731 2138
rect 783 2142 787 2143
rect 783 2137 787 2138
rect 791 2142 795 2143
rect 791 2137 795 2138
rect 847 2142 851 2143
rect 847 2137 851 2138
rect 855 2142 859 2143
rect 855 2137 859 2138
rect 911 2142 915 2143
rect 911 2137 915 2138
rect 967 2142 971 2143
rect 967 2137 971 2138
rect 1023 2142 1027 2143
rect 1023 2137 1027 2138
rect 1079 2142 1083 2143
rect 1079 2137 1083 2138
rect 1143 2142 1147 2143
rect 1143 2137 1147 2138
rect 1239 2142 1243 2143
rect 1239 2137 1243 2138
rect 112 2130 114 2137
rect 382 2136 388 2137
rect 382 2132 383 2136
rect 387 2132 388 2136
rect 382 2131 388 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 462 2136 468 2137
rect 462 2132 463 2136
rect 467 2132 468 2136
rect 462 2131 468 2132
rect 502 2136 508 2137
rect 502 2132 503 2136
rect 507 2132 508 2136
rect 502 2131 508 2132
rect 550 2136 556 2137
rect 550 2132 551 2136
rect 555 2132 556 2136
rect 550 2131 556 2132
rect 606 2136 612 2137
rect 606 2132 607 2136
rect 611 2132 612 2136
rect 606 2131 612 2132
rect 662 2136 668 2137
rect 662 2132 663 2136
rect 667 2132 668 2136
rect 662 2131 668 2132
rect 726 2136 732 2137
rect 726 2132 727 2136
rect 731 2132 732 2136
rect 726 2131 732 2132
rect 790 2136 796 2137
rect 790 2132 791 2136
rect 795 2132 796 2136
rect 790 2131 796 2132
rect 854 2136 860 2137
rect 854 2132 855 2136
rect 859 2132 860 2136
rect 854 2131 860 2132
rect 910 2136 916 2137
rect 910 2132 911 2136
rect 915 2132 916 2136
rect 910 2131 916 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1022 2136 1028 2137
rect 1022 2132 1023 2136
rect 1027 2132 1028 2136
rect 1022 2131 1028 2132
rect 1078 2136 1084 2137
rect 1078 2132 1079 2136
rect 1083 2132 1084 2136
rect 1078 2131 1084 2132
rect 1142 2136 1148 2137
rect 1142 2132 1143 2136
rect 1147 2132 1148 2136
rect 1142 2131 1148 2132
rect 1240 2130 1242 2137
rect 110 2129 116 2130
rect 110 2125 111 2129
rect 115 2125 116 2129
rect 110 2124 116 2125
rect 1238 2129 1244 2130
rect 1238 2125 1239 2129
rect 1243 2125 1244 2129
rect 1280 2125 1282 2157
rect 1304 2148 1306 2157
rect 1352 2148 1354 2157
rect 1440 2148 1442 2157
rect 1536 2148 1538 2157
rect 1632 2148 1634 2157
rect 1728 2148 1730 2157
rect 1816 2148 1818 2157
rect 1896 2148 1898 2157
rect 1976 2148 1978 2157
rect 2048 2148 2050 2157
rect 2112 2148 2114 2157
rect 2176 2148 2178 2157
rect 2240 2148 2242 2157
rect 2312 2148 2314 2157
rect 2360 2148 2362 2157
rect 1302 2147 1308 2148
rect 1302 2143 1303 2147
rect 1307 2143 1308 2147
rect 1302 2142 1308 2143
rect 1350 2147 1356 2148
rect 1350 2143 1351 2147
rect 1355 2143 1356 2147
rect 1350 2142 1356 2143
rect 1438 2147 1444 2148
rect 1438 2143 1439 2147
rect 1443 2143 1444 2147
rect 1438 2142 1444 2143
rect 1534 2147 1540 2148
rect 1534 2143 1535 2147
rect 1539 2143 1540 2147
rect 1534 2142 1540 2143
rect 1630 2147 1636 2148
rect 1630 2143 1631 2147
rect 1635 2143 1636 2147
rect 1630 2142 1636 2143
rect 1726 2147 1732 2148
rect 1726 2143 1727 2147
rect 1731 2143 1732 2147
rect 1726 2142 1732 2143
rect 1814 2147 1820 2148
rect 1814 2143 1815 2147
rect 1819 2143 1820 2147
rect 1814 2142 1820 2143
rect 1894 2147 1900 2148
rect 1894 2143 1895 2147
rect 1899 2143 1900 2147
rect 1894 2142 1900 2143
rect 1974 2147 1980 2148
rect 1974 2143 1975 2147
rect 1979 2143 1980 2147
rect 1974 2142 1980 2143
rect 2046 2147 2052 2148
rect 2046 2143 2047 2147
rect 2051 2143 2052 2147
rect 2046 2142 2052 2143
rect 2110 2147 2116 2148
rect 2110 2143 2111 2147
rect 2115 2143 2116 2147
rect 2110 2142 2116 2143
rect 2174 2147 2180 2148
rect 2174 2143 2175 2147
rect 2179 2143 2180 2147
rect 2174 2142 2180 2143
rect 2238 2147 2244 2148
rect 2238 2143 2239 2147
rect 2243 2143 2244 2147
rect 2238 2142 2244 2143
rect 2310 2147 2316 2148
rect 2310 2143 2311 2147
rect 2315 2143 2316 2147
rect 2310 2142 2316 2143
rect 2358 2147 2364 2148
rect 2358 2143 2359 2147
rect 2363 2143 2364 2147
rect 2358 2142 2364 2143
rect 2408 2125 2410 2157
rect 1238 2124 1244 2125
rect 1278 2124 1284 2125
rect 1278 2120 1279 2124
rect 1283 2120 1284 2124
rect 1278 2119 1284 2120
rect 2406 2124 2412 2125
rect 2406 2120 2407 2124
rect 2411 2120 2412 2124
rect 2406 2119 2412 2120
rect 110 2112 116 2113
rect 110 2108 111 2112
rect 115 2108 116 2112
rect 110 2107 116 2108
rect 1238 2112 1244 2113
rect 1238 2108 1239 2112
rect 1243 2108 1244 2112
rect 1238 2107 1244 2108
rect 1278 2107 1284 2108
rect 112 2075 114 2107
rect 382 2089 388 2090
rect 382 2085 383 2089
rect 387 2085 388 2089
rect 382 2084 388 2085
rect 422 2089 428 2090
rect 422 2085 423 2089
rect 427 2085 428 2089
rect 422 2084 428 2085
rect 462 2089 468 2090
rect 462 2085 463 2089
rect 467 2085 468 2089
rect 462 2084 468 2085
rect 502 2089 508 2090
rect 502 2085 503 2089
rect 507 2085 508 2089
rect 502 2084 508 2085
rect 550 2089 556 2090
rect 550 2085 551 2089
rect 555 2085 556 2089
rect 550 2084 556 2085
rect 606 2089 612 2090
rect 606 2085 607 2089
rect 611 2085 612 2089
rect 606 2084 612 2085
rect 662 2089 668 2090
rect 662 2085 663 2089
rect 667 2085 668 2089
rect 662 2084 668 2085
rect 726 2089 732 2090
rect 726 2085 727 2089
rect 731 2085 732 2089
rect 726 2084 732 2085
rect 790 2089 796 2090
rect 790 2085 791 2089
rect 795 2085 796 2089
rect 790 2084 796 2085
rect 854 2089 860 2090
rect 854 2085 855 2089
rect 859 2085 860 2089
rect 854 2084 860 2085
rect 910 2089 916 2090
rect 910 2085 911 2089
rect 915 2085 916 2089
rect 910 2084 916 2085
rect 966 2089 972 2090
rect 966 2085 967 2089
rect 971 2085 972 2089
rect 966 2084 972 2085
rect 1022 2089 1028 2090
rect 1022 2085 1023 2089
rect 1027 2085 1028 2089
rect 1022 2084 1028 2085
rect 1078 2089 1084 2090
rect 1078 2085 1079 2089
rect 1083 2085 1084 2089
rect 1078 2084 1084 2085
rect 1142 2089 1148 2090
rect 1142 2085 1143 2089
rect 1147 2085 1148 2089
rect 1142 2084 1148 2085
rect 384 2075 386 2084
rect 424 2075 426 2084
rect 464 2075 466 2084
rect 504 2075 506 2084
rect 552 2075 554 2084
rect 608 2075 610 2084
rect 664 2075 666 2084
rect 728 2075 730 2084
rect 792 2075 794 2084
rect 856 2075 858 2084
rect 912 2075 914 2084
rect 968 2075 970 2084
rect 1024 2075 1026 2084
rect 1080 2075 1082 2084
rect 1144 2075 1146 2084
rect 1240 2075 1242 2107
rect 1278 2103 1279 2107
rect 1283 2103 1284 2107
rect 1278 2102 1284 2103
rect 2406 2107 2412 2108
rect 2406 2103 2407 2107
rect 2411 2103 2412 2107
rect 2406 2102 2412 2103
rect 1280 2091 1282 2102
rect 1302 2100 1308 2101
rect 1302 2096 1303 2100
rect 1307 2096 1308 2100
rect 1302 2095 1308 2096
rect 1350 2100 1356 2101
rect 1350 2096 1351 2100
rect 1355 2096 1356 2100
rect 1350 2095 1356 2096
rect 1438 2100 1444 2101
rect 1438 2096 1439 2100
rect 1443 2096 1444 2100
rect 1438 2095 1444 2096
rect 1534 2100 1540 2101
rect 1534 2096 1535 2100
rect 1539 2096 1540 2100
rect 1534 2095 1540 2096
rect 1630 2100 1636 2101
rect 1630 2096 1631 2100
rect 1635 2096 1636 2100
rect 1630 2095 1636 2096
rect 1726 2100 1732 2101
rect 1726 2096 1727 2100
rect 1731 2096 1732 2100
rect 1726 2095 1732 2096
rect 1814 2100 1820 2101
rect 1814 2096 1815 2100
rect 1819 2096 1820 2100
rect 1814 2095 1820 2096
rect 1894 2100 1900 2101
rect 1894 2096 1895 2100
rect 1899 2096 1900 2100
rect 1894 2095 1900 2096
rect 1974 2100 1980 2101
rect 1974 2096 1975 2100
rect 1979 2096 1980 2100
rect 1974 2095 1980 2096
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2046 2095 2052 2096
rect 2110 2100 2116 2101
rect 2110 2096 2111 2100
rect 2115 2096 2116 2100
rect 2110 2095 2116 2096
rect 2174 2100 2180 2101
rect 2174 2096 2175 2100
rect 2179 2096 2180 2100
rect 2174 2095 2180 2096
rect 2238 2100 2244 2101
rect 2238 2096 2239 2100
rect 2243 2096 2244 2100
rect 2238 2095 2244 2096
rect 2310 2100 2316 2101
rect 2310 2096 2311 2100
rect 2315 2096 2316 2100
rect 2310 2095 2316 2096
rect 2358 2100 2364 2101
rect 2358 2096 2359 2100
rect 2363 2096 2364 2100
rect 2358 2095 2364 2096
rect 1304 2091 1306 2095
rect 1352 2091 1354 2095
rect 1440 2091 1442 2095
rect 1536 2091 1538 2095
rect 1632 2091 1634 2095
rect 1728 2091 1730 2095
rect 1816 2091 1818 2095
rect 1896 2091 1898 2095
rect 1976 2091 1978 2095
rect 2048 2091 2050 2095
rect 2112 2091 2114 2095
rect 2176 2091 2178 2095
rect 2240 2091 2242 2095
rect 2312 2091 2314 2095
rect 2360 2091 2362 2095
rect 2408 2091 2410 2102
rect 1279 2090 1283 2091
rect 1279 2085 1283 2086
rect 1303 2090 1307 2091
rect 1303 2085 1307 2086
rect 1343 2090 1347 2091
rect 1343 2085 1347 2086
rect 1351 2090 1355 2091
rect 1351 2085 1355 2086
rect 1399 2090 1403 2091
rect 1399 2085 1403 2086
rect 1439 2090 1443 2091
rect 1439 2085 1443 2086
rect 1479 2090 1483 2091
rect 1479 2085 1483 2086
rect 1535 2090 1539 2091
rect 1535 2085 1539 2086
rect 1567 2090 1571 2091
rect 1567 2085 1571 2086
rect 1631 2090 1635 2091
rect 1631 2085 1635 2086
rect 1663 2090 1667 2091
rect 1663 2085 1667 2086
rect 1727 2090 1731 2091
rect 1727 2085 1731 2086
rect 1759 2090 1763 2091
rect 1759 2085 1763 2086
rect 1815 2090 1819 2091
rect 1815 2085 1819 2086
rect 1847 2090 1851 2091
rect 1847 2085 1851 2086
rect 1895 2090 1899 2091
rect 1895 2085 1899 2086
rect 1935 2090 1939 2091
rect 1935 2085 1939 2086
rect 1975 2090 1979 2091
rect 1975 2085 1979 2086
rect 2015 2090 2019 2091
rect 2015 2085 2019 2086
rect 2047 2090 2051 2091
rect 2047 2085 2051 2086
rect 2095 2090 2099 2091
rect 2095 2085 2099 2086
rect 2111 2090 2115 2091
rect 2111 2085 2115 2086
rect 2167 2090 2171 2091
rect 2167 2085 2171 2086
rect 2175 2090 2179 2091
rect 2175 2085 2179 2086
rect 2239 2090 2243 2091
rect 2239 2085 2243 2086
rect 2311 2090 2315 2091
rect 2311 2085 2315 2086
rect 2359 2090 2363 2091
rect 2359 2085 2363 2086
rect 2407 2090 2411 2091
rect 2407 2085 2411 2086
rect 1280 2078 1282 2085
rect 1302 2084 1308 2085
rect 1302 2080 1303 2084
rect 1307 2080 1308 2084
rect 1302 2079 1308 2080
rect 1342 2084 1348 2085
rect 1342 2080 1343 2084
rect 1347 2080 1348 2084
rect 1342 2079 1348 2080
rect 1398 2084 1404 2085
rect 1398 2080 1399 2084
rect 1403 2080 1404 2084
rect 1398 2079 1404 2080
rect 1478 2084 1484 2085
rect 1478 2080 1479 2084
rect 1483 2080 1484 2084
rect 1478 2079 1484 2080
rect 1566 2084 1572 2085
rect 1566 2080 1567 2084
rect 1571 2080 1572 2084
rect 1566 2079 1572 2080
rect 1662 2084 1668 2085
rect 1662 2080 1663 2084
rect 1667 2080 1668 2084
rect 1662 2079 1668 2080
rect 1758 2084 1764 2085
rect 1758 2080 1759 2084
rect 1763 2080 1764 2084
rect 1758 2079 1764 2080
rect 1846 2084 1852 2085
rect 1846 2080 1847 2084
rect 1851 2080 1852 2084
rect 1846 2079 1852 2080
rect 1934 2084 1940 2085
rect 1934 2080 1935 2084
rect 1939 2080 1940 2084
rect 1934 2079 1940 2080
rect 2014 2084 2020 2085
rect 2014 2080 2015 2084
rect 2019 2080 2020 2084
rect 2014 2079 2020 2080
rect 2094 2084 2100 2085
rect 2094 2080 2095 2084
rect 2099 2080 2100 2084
rect 2094 2079 2100 2080
rect 2166 2084 2172 2085
rect 2166 2080 2167 2084
rect 2171 2080 2172 2084
rect 2166 2079 2172 2080
rect 2238 2084 2244 2085
rect 2238 2080 2239 2084
rect 2243 2080 2244 2084
rect 2238 2079 2244 2080
rect 2310 2084 2316 2085
rect 2310 2080 2311 2084
rect 2315 2080 2316 2084
rect 2310 2079 2316 2080
rect 2358 2084 2364 2085
rect 2358 2080 2359 2084
rect 2363 2080 2364 2084
rect 2358 2079 2364 2080
rect 2408 2078 2410 2085
rect 1278 2077 1284 2078
rect 111 2074 115 2075
rect 111 2069 115 2070
rect 383 2074 387 2075
rect 383 2069 387 2070
rect 423 2074 427 2075
rect 423 2069 427 2070
rect 463 2074 467 2075
rect 463 2069 467 2070
rect 503 2074 507 2075
rect 503 2069 507 2070
rect 543 2074 547 2075
rect 543 2069 547 2070
rect 551 2074 555 2075
rect 551 2069 555 2070
rect 583 2074 587 2075
rect 583 2069 587 2070
rect 607 2074 611 2075
rect 607 2069 611 2070
rect 631 2074 635 2075
rect 631 2069 635 2070
rect 663 2074 667 2075
rect 663 2069 667 2070
rect 687 2074 691 2075
rect 687 2069 691 2070
rect 727 2074 731 2075
rect 727 2069 731 2070
rect 743 2074 747 2075
rect 743 2069 747 2070
rect 791 2074 795 2075
rect 791 2069 795 2070
rect 799 2074 803 2075
rect 799 2069 803 2070
rect 847 2074 851 2075
rect 847 2069 851 2070
rect 855 2074 859 2075
rect 855 2069 859 2070
rect 903 2074 907 2075
rect 903 2069 907 2070
rect 911 2074 915 2075
rect 911 2069 915 2070
rect 959 2074 963 2075
rect 959 2069 963 2070
rect 967 2074 971 2075
rect 967 2069 971 2070
rect 1015 2074 1019 2075
rect 1015 2069 1019 2070
rect 1023 2074 1027 2075
rect 1023 2069 1027 2070
rect 1071 2074 1075 2075
rect 1071 2069 1075 2070
rect 1079 2074 1083 2075
rect 1079 2069 1083 2070
rect 1143 2074 1147 2075
rect 1143 2069 1147 2070
rect 1239 2074 1243 2075
rect 1278 2073 1279 2077
rect 1283 2073 1284 2077
rect 1278 2072 1284 2073
rect 2406 2077 2412 2078
rect 2406 2073 2407 2077
rect 2411 2073 2412 2077
rect 2406 2072 2412 2073
rect 1239 2069 1243 2070
rect 112 2037 114 2069
rect 384 2060 386 2069
rect 424 2060 426 2069
rect 464 2060 466 2069
rect 504 2060 506 2069
rect 544 2060 546 2069
rect 584 2060 586 2069
rect 632 2060 634 2069
rect 688 2060 690 2069
rect 744 2060 746 2069
rect 800 2060 802 2069
rect 848 2060 850 2069
rect 904 2060 906 2069
rect 960 2060 962 2069
rect 1016 2060 1018 2069
rect 1072 2060 1074 2069
rect 382 2059 388 2060
rect 382 2055 383 2059
rect 387 2055 388 2059
rect 382 2054 388 2055
rect 422 2059 428 2060
rect 422 2055 423 2059
rect 427 2055 428 2059
rect 422 2054 428 2055
rect 462 2059 468 2060
rect 462 2055 463 2059
rect 467 2055 468 2059
rect 462 2054 468 2055
rect 502 2059 508 2060
rect 502 2055 503 2059
rect 507 2055 508 2059
rect 502 2054 508 2055
rect 542 2059 548 2060
rect 542 2055 543 2059
rect 547 2055 548 2059
rect 542 2054 548 2055
rect 582 2059 588 2060
rect 582 2055 583 2059
rect 587 2055 588 2059
rect 582 2054 588 2055
rect 630 2059 636 2060
rect 630 2055 631 2059
rect 635 2055 636 2059
rect 630 2054 636 2055
rect 686 2059 692 2060
rect 686 2055 687 2059
rect 691 2055 692 2059
rect 686 2054 692 2055
rect 742 2059 748 2060
rect 742 2055 743 2059
rect 747 2055 748 2059
rect 742 2054 748 2055
rect 798 2059 804 2060
rect 798 2055 799 2059
rect 803 2055 804 2059
rect 798 2054 804 2055
rect 846 2059 852 2060
rect 846 2055 847 2059
rect 851 2055 852 2059
rect 846 2054 852 2055
rect 902 2059 908 2060
rect 902 2055 903 2059
rect 907 2055 908 2059
rect 902 2054 908 2055
rect 958 2059 964 2060
rect 958 2055 959 2059
rect 963 2055 964 2059
rect 958 2054 964 2055
rect 1014 2059 1020 2060
rect 1014 2055 1015 2059
rect 1019 2055 1020 2059
rect 1014 2054 1020 2055
rect 1070 2059 1076 2060
rect 1070 2055 1071 2059
rect 1075 2055 1076 2059
rect 1070 2054 1076 2055
rect 1240 2037 1242 2069
rect 1278 2060 1284 2061
rect 1278 2056 1279 2060
rect 1283 2056 1284 2060
rect 1278 2055 1284 2056
rect 2406 2060 2412 2061
rect 2406 2056 2407 2060
rect 2411 2056 2412 2060
rect 2406 2055 2412 2056
rect 110 2036 116 2037
rect 110 2032 111 2036
rect 115 2032 116 2036
rect 110 2031 116 2032
rect 1238 2036 1244 2037
rect 1238 2032 1239 2036
rect 1243 2032 1244 2036
rect 1238 2031 1244 2032
rect 110 2019 116 2020
rect 110 2015 111 2019
rect 115 2015 116 2019
rect 110 2014 116 2015
rect 1238 2019 1244 2020
rect 1238 2015 1239 2019
rect 1243 2015 1244 2019
rect 1280 2015 1282 2055
rect 1302 2037 1308 2038
rect 1302 2033 1303 2037
rect 1307 2033 1308 2037
rect 1302 2032 1308 2033
rect 1342 2037 1348 2038
rect 1342 2033 1343 2037
rect 1347 2033 1348 2037
rect 1342 2032 1348 2033
rect 1398 2037 1404 2038
rect 1398 2033 1399 2037
rect 1403 2033 1404 2037
rect 1398 2032 1404 2033
rect 1478 2037 1484 2038
rect 1478 2033 1479 2037
rect 1483 2033 1484 2037
rect 1478 2032 1484 2033
rect 1566 2037 1572 2038
rect 1566 2033 1567 2037
rect 1571 2033 1572 2037
rect 1566 2032 1572 2033
rect 1662 2037 1668 2038
rect 1662 2033 1663 2037
rect 1667 2033 1668 2037
rect 1662 2032 1668 2033
rect 1758 2037 1764 2038
rect 1758 2033 1759 2037
rect 1763 2033 1764 2037
rect 1758 2032 1764 2033
rect 1846 2037 1852 2038
rect 1846 2033 1847 2037
rect 1851 2033 1852 2037
rect 1846 2032 1852 2033
rect 1934 2037 1940 2038
rect 1934 2033 1935 2037
rect 1939 2033 1940 2037
rect 1934 2032 1940 2033
rect 2014 2037 2020 2038
rect 2014 2033 2015 2037
rect 2019 2033 2020 2037
rect 2014 2032 2020 2033
rect 2094 2037 2100 2038
rect 2094 2033 2095 2037
rect 2099 2033 2100 2037
rect 2094 2032 2100 2033
rect 2166 2037 2172 2038
rect 2166 2033 2167 2037
rect 2171 2033 2172 2037
rect 2166 2032 2172 2033
rect 2238 2037 2244 2038
rect 2238 2033 2239 2037
rect 2243 2033 2244 2037
rect 2238 2032 2244 2033
rect 2310 2037 2316 2038
rect 2310 2033 2311 2037
rect 2315 2033 2316 2037
rect 2310 2032 2316 2033
rect 2358 2037 2364 2038
rect 2358 2033 2359 2037
rect 2363 2033 2364 2037
rect 2358 2032 2364 2033
rect 1304 2015 1306 2032
rect 1344 2015 1346 2032
rect 1400 2015 1402 2032
rect 1480 2015 1482 2032
rect 1568 2015 1570 2032
rect 1664 2015 1666 2032
rect 1760 2015 1762 2032
rect 1848 2015 1850 2032
rect 1936 2015 1938 2032
rect 2016 2015 2018 2032
rect 2096 2015 2098 2032
rect 2168 2015 2170 2032
rect 2240 2015 2242 2032
rect 2312 2015 2314 2032
rect 2360 2015 2362 2032
rect 2408 2015 2410 2055
rect 1238 2014 1244 2015
rect 1279 2014 1283 2015
rect 112 1999 114 2014
rect 382 2012 388 2013
rect 382 2008 383 2012
rect 387 2008 388 2012
rect 382 2007 388 2008
rect 422 2012 428 2013
rect 422 2008 423 2012
rect 427 2008 428 2012
rect 422 2007 428 2008
rect 462 2012 468 2013
rect 462 2008 463 2012
rect 467 2008 468 2012
rect 462 2007 468 2008
rect 502 2012 508 2013
rect 502 2008 503 2012
rect 507 2008 508 2012
rect 502 2007 508 2008
rect 542 2012 548 2013
rect 542 2008 543 2012
rect 547 2008 548 2012
rect 542 2007 548 2008
rect 582 2012 588 2013
rect 582 2008 583 2012
rect 587 2008 588 2012
rect 582 2007 588 2008
rect 630 2012 636 2013
rect 630 2008 631 2012
rect 635 2008 636 2012
rect 630 2007 636 2008
rect 686 2012 692 2013
rect 686 2008 687 2012
rect 691 2008 692 2012
rect 686 2007 692 2008
rect 742 2012 748 2013
rect 742 2008 743 2012
rect 747 2008 748 2012
rect 742 2007 748 2008
rect 798 2012 804 2013
rect 798 2008 799 2012
rect 803 2008 804 2012
rect 798 2007 804 2008
rect 846 2012 852 2013
rect 846 2008 847 2012
rect 851 2008 852 2012
rect 846 2007 852 2008
rect 902 2012 908 2013
rect 902 2008 903 2012
rect 907 2008 908 2012
rect 902 2007 908 2008
rect 958 2012 964 2013
rect 958 2008 959 2012
rect 963 2008 964 2012
rect 958 2007 964 2008
rect 1014 2012 1020 2013
rect 1014 2008 1015 2012
rect 1019 2008 1020 2012
rect 1014 2007 1020 2008
rect 1070 2012 1076 2013
rect 1070 2008 1071 2012
rect 1075 2008 1076 2012
rect 1070 2007 1076 2008
rect 384 1999 386 2007
rect 424 1999 426 2007
rect 464 1999 466 2007
rect 504 1999 506 2007
rect 544 1999 546 2007
rect 584 1999 586 2007
rect 632 1999 634 2007
rect 688 1999 690 2007
rect 744 1999 746 2007
rect 800 1999 802 2007
rect 848 1999 850 2007
rect 904 1999 906 2007
rect 960 1999 962 2007
rect 1016 1999 1018 2007
rect 1072 1999 1074 2007
rect 1240 1999 1242 2014
rect 1279 2009 1283 2010
rect 1303 2014 1307 2015
rect 1303 2009 1307 2010
rect 1343 2014 1347 2015
rect 1343 2009 1347 2010
rect 1351 2014 1355 2015
rect 1351 2009 1355 2010
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1423 2014 1427 2015
rect 1423 2009 1427 2010
rect 1479 2014 1483 2015
rect 1479 2009 1483 2010
rect 1495 2014 1499 2015
rect 1495 2009 1499 2010
rect 1567 2014 1571 2015
rect 1567 2009 1571 2010
rect 1575 2014 1579 2015
rect 1575 2009 1579 2010
rect 1663 2014 1667 2015
rect 1663 2009 1667 2010
rect 1751 2014 1755 2015
rect 1751 2009 1755 2010
rect 1759 2014 1763 2015
rect 1759 2009 1763 2010
rect 1839 2014 1843 2015
rect 1839 2009 1843 2010
rect 1847 2014 1851 2015
rect 1847 2009 1851 2010
rect 1919 2014 1923 2015
rect 1919 2009 1923 2010
rect 1935 2014 1939 2015
rect 1935 2009 1939 2010
rect 1999 2014 2003 2015
rect 1999 2009 2003 2010
rect 2015 2014 2019 2015
rect 2015 2009 2019 2010
rect 2071 2014 2075 2015
rect 2071 2009 2075 2010
rect 2095 2014 2099 2015
rect 2095 2009 2099 2010
rect 2135 2014 2139 2015
rect 2135 2009 2139 2010
rect 2167 2014 2171 2015
rect 2167 2009 2171 2010
rect 2191 2014 2195 2015
rect 2191 2009 2195 2010
rect 2239 2014 2243 2015
rect 2239 2009 2243 2010
rect 2255 2014 2259 2015
rect 2255 2009 2259 2010
rect 2311 2014 2315 2015
rect 2311 2009 2315 2010
rect 2319 2014 2323 2015
rect 2319 2009 2323 2010
rect 2359 2014 2363 2015
rect 2359 2009 2363 2010
rect 2407 2014 2411 2015
rect 2407 2009 2411 2010
rect 111 1998 115 1999
rect 111 1993 115 1994
rect 367 1998 371 1999
rect 367 1993 371 1994
rect 383 1998 387 1999
rect 383 1993 387 1994
rect 407 1998 411 1999
rect 407 1993 411 1994
rect 423 1998 427 1999
rect 423 1993 427 1994
rect 455 1998 459 1999
rect 455 1993 459 1994
rect 463 1998 467 1999
rect 463 1993 467 1994
rect 503 1998 507 1999
rect 503 1993 507 1994
rect 511 1998 515 1999
rect 511 1993 515 1994
rect 543 1998 547 1999
rect 543 1993 547 1994
rect 567 1998 571 1999
rect 567 1993 571 1994
rect 583 1998 587 1999
rect 583 1993 587 1994
rect 631 1998 635 1999
rect 631 1993 635 1994
rect 687 1998 691 1999
rect 687 1993 691 1994
rect 695 1998 699 1999
rect 695 1993 699 1994
rect 743 1998 747 1999
rect 743 1993 747 1994
rect 759 1998 763 1999
rect 759 1993 763 1994
rect 799 1998 803 1999
rect 799 1993 803 1994
rect 815 1998 819 1999
rect 815 1993 819 1994
rect 847 1998 851 1999
rect 847 1993 851 1994
rect 871 1998 875 1999
rect 871 1993 875 1994
rect 903 1998 907 1999
rect 903 1993 907 1994
rect 935 1998 939 1999
rect 935 1993 939 1994
rect 959 1998 963 1999
rect 959 1993 963 1994
rect 999 1998 1003 1999
rect 999 1993 1003 1994
rect 1015 1998 1019 1999
rect 1015 1993 1019 1994
rect 1063 1998 1067 1999
rect 1063 1993 1067 1994
rect 1071 1998 1075 1999
rect 1071 1993 1075 1994
rect 1239 1998 1243 1999
rect 1239 1993 1243 1994
rect 112 1986 114 1993
rect 366 1992 372 1993
rect 366 1988 367 1992
rect 371 1988 372 1992
rect 366 1987 372 1988
rect 406 1992 412 1993
rect 406 1988 407 1992
rect 411 1988 412 1992
rect 406 1987 412 1988
rect 454 1992 460 1993
rect 454 1988 455 1992
rect 459 1988 460 1992
rect 454 1987 460 1988
rect 510 1992 516 1993
rect 510 1988 511 1992
rect 515 1988 516 1992
rect 510 1987 516 1988
rect 566 1992 572 1993
rect 566 1988 567 1992
rect 571 1988 572 1992
rect 566 1987 572 1988
rect 630 1992 636 1993
rect 630 1988 631 1992
rect 635 1988 636 1992
rect 630 1987 636 1988
rect 694 1992 700 1993
rect 694 1988 695 1992
rect 699 1988 700 1992
rect 694 1987 700 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 870 1992 876 1993
rect 870 1988 871 1992
rect 875 1988 876 1992
rect 870 1987 876 1988
rect 934 1992 940 1993
rect 934 1988 935 1992
rect 939 1988 940 1992
rect 934 1987 940 1988
rect 998 1992 1004 1993
rect 998 1988 999 1992
rect 1003 1988 1004 1992
rect 998 1987 1004 1988
rect 1062 1992 1068 1993
rect 1062 1988 1063 1992
rect 1067 1988 1068 1992
rect 1062 1987 1068 1988
rect 1240 1986 1242 1993
rect 110 1985 116 1986
rect 110 1981 111 1985
rect 115 1981 116 1985
rect 110 1980 116 1981
rect 1238 1985 1244 1986
rect 1238 1981 1239 1985
rect 1243 1981 1244 1985
rect 1238 1980 1244 1981
rect 1280 1977 1282 2009
rect 1304 2000 1306 2009
rect 1352 2000 1354 2009
rect 1424 2000 1426 2009
rect 1496 2000 1498 2009
rect 1576 2000 1578 2009
rect 1664 2000 1666 2009
rect 1752 2000 1754 2009
rect 1840 2000 1842 2009
rect 1920 2000 1922 2009
rect 2000 2000 2002 2009
rect 2072 2000 2074 2009
rect 2136 2000 2138 2009
rect 2192 2000 2194 2009
rect 2256 2000 2258 2009
rect 2320 2000 2322 2009
rect 2360 2000 2362 2009
rect 1302 1999 1308 2000
rect 1302 1995 1303 1999
rect 1307 1995 1308 1999
rect 1302 1994 1308 1995
rect 1350 1999 1356 2000
rect 1350 1995 1351 1999
rect 1355 1995 1356 1999
rect 1350 1994 1356 1995
rect 1422 1999 1428 2000
rect 1422 1995 1423 1999
rect 1427 1995 1428 1999
rect 1422 1994 1428 1995
rect 1494 1999 1500 2000
rect 1494 1995 1495 1999
rect 1499 1995 1500 1999
rect 1494 1994 1500 1995
rect 1574 1999 1580 2000
rect 1574 1995 1575 1999
rect 1579 1995 1580 1999
rect 1574 1994 1580 1995
rect 1662 1999 1668 2000
rect 1662 1995 1663 1999
rect 1667 1995 1668 1999
rect 1662 1994 1668 1995
rect 1750 1999 1756 2000
rect 1750 1995 1751 1999
rect 1755 1995 1756 1999
rect 1750 1994 1756 1995
rect 1838 1999 1844 2000
rect 1838 1995 1839 1999
rect 1843 1995 1844 1999
rect 1838 1994 1844 1995
rect 1918 1999 1924 2000
rect 1918 1995 1919 1999
rect 1923 1995 1924 1999
rect 1918 1994 1924 1995
rect 1998 1999 2004 2000
rect 1998 1995 1999 1999
rect 2003 1995 2004 1999
rect 1998 1994 2004 1995
rect 2070 1999 2076 2000
rect 2070 1995 2071 1999
rect 2075 1995 2076 1999
rect 2070 1994 2076 1995
rect 2134 1999 2140 2000
rect 2134 1995 2135 1999
rect 2139 1995 2140 1999
rect 2134 1994 2140 1995
rect 2190 1999 2196 2000
rect 2190 1995 2191 1999
rect 2195 1995 2196 1999
rect 2190 1994 2196 1995
rect 2254 1999 2260 2000
rect 2254 1995 2255 1999
rect 2259 1995 2260 1999
rect 2254 1994 2260 1995
rect 2318 1999 2324 2000
rect 2318 1995 2319 1999
rect 2323 1995 2324 1999
rect 2318 1994 2324 1995
rect 2358 1999 2364 2000
rect 2358 1995 2359 1999
rect 2363 1995 2364 1999
rect 2358 1994 2364 1995
rect 2408 1977 2410 2009
rect 1278 1976 1284 1977
rect 1278 1972 1279 1976
rect 1283 1972 1284 1976
rect 1278 1971 1284 1972
rect 2406 1976 2412 1977
rect 2406 1972 2407 1976
rect 2411 1972 2412 1976
rect 2406 1971 2412 1972
rect 110 1968 116 1969
rect 110 1964 111 1968
rect 115 1964 116 1968
rect 110 1963 116 1964
rect 1238 1968 1244 1969
rect 1238 1964 1239 1968
rect 1243 1964 1244 1968
rect 1238 1963 1244 1964
rect 112 1927 114 1963
rect 366 1945 372 1946
rect 366 1941 367 1945
rect 371 1941 372 1945
rect 366 1940 372 1941
rect 406 1945 412 1946
rect 406 1941 407 1945
rect 411 1941 412 1945
rect 406 1940 412 1941
rect 454 1945 460 1946
rect 454 1941 455 1945
rect 459 1941 460 1945
rect 454 1940 460 1941
rect 510 1945 516 1946
rect 510 1941 511 1945
rect 515 1941 516 1945
rect 510 1940 516 1941
rect 566 1945 572 1946
rect 566 1941 567 1945
rect 571 1941 572 1945
rect 566 1940 572 1941
rect 630 1945 636 1946
rect 630 1941 631 1945
rect 635 1941 636 1945
rect 630 1940 636 1941
rect 694 1945 700 1946
rect 694 1941 695 1945
rect 699 1941 700 1945
rect 694 1940 700 1941
rect 758 1945 764 1946
rect 758 1941 759 1945
rect 763 1941 764 1945
rect 758 1940 764 1941
rect 814 1945 820 1946
rect 814 1941 815 1945
rect 819 1941 820 1945
rect 814 1940 820 1941
rect 870 1945 876 1946
rect 870 1941 871 1945
rect 875 1941 876 1945
rect 870 1940 876 1941
rect 934 1945 940 1946
rect 934 1941 935 1945
rect 939 1941 940 1945
rect 934 1940 940 1941
rect 998 1945 1004 1946
rect 998 1941 999 1945
rect 1003 1941 1004 1945
rect 998 1940 1004 1941
rect 1062 1945 1068 1946
rect 1062 1941 1063 1945
rect 1067 1941 1068 1945
rect 1062 1940 1068 1941
rect 368 1927 370 1940
rect 408 1927 410 1940
rect 456 1927 458 1940
rect 512 1927 514 1940
rect 568 1927 570 1940
rect 632 1927 634 1940
rect 696 1927 698 1940
rect 760 1927 762 1940
rect 816 1927 818 1940
rect 872 1927 874 1940
rect 936 1927 938 1940
rect 1000 1927 1002 1940
rect 1064 1927 1066 1940
rect 1240 1927 1242 1963
rect 1278 1959 1284 1960
rect 1278 1955 1279 1959
rect 1283 1955 1284 1959
rect 1278 1954 1284 1955
rect 2406 1959 2412 1960
rect 2406 1955 2407 1959
rect 2411 1955 2412 1959
rect 2406 1954 2412 1955
rect 1280 1947 1282 1954
rect 1302 1952 1308 1953
rect 1302 1948 1303 1952
rect 1307 1948 1308 1952
rect 1302 1947 1308 1948
rect 1350 1952 1356 1953
rect 1350 1948 1351 1952
rect 1355 1948 1356 1952
rect 1350 1947 1356 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1494 1952 1500 1953
rect 1494 1948 1495 1952
rect 1499 1948 1500 1952
rect 1494 1947 1500 1948
rect 1574 1952 1580 1953
rect 1574 1948 1575 1952
rect 1579 1948 1580 1952
rect 1574 1947 1580 1948
rect 1662 1952 1668 1953
rect 1662 1948 1663 1952
rect 1667 1948 1668 1952
rect 1662 1947 1668 1948
rect 1750 1952 1756 1953
rect 1750 1948 1751 1952
rect 1755 1948 1756 1952
rect 1750 1947 1756 1948
rect 1838 1952 1844 1953
rect 1838 1948 1839 1952
rect 1843 1948 1844 1952
rect 1838 1947 1844 1948
rect 1918 1952 1924 1953
rect 1918 1948 1919 1952
rect 1923 1948 1924 1952
rect 1918 1947 1924 1948
rect 1998 1952 2004 1953
rect 1998 1948 1999 1952
rect 2003 1948 2004 1952
rect 1998 1947 2004 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2134 1952 2140 1953
rect 2134 1948 2135 1952
rect 2139 1948 2140 1952
rect 2134 1947 2140 1948
rect 2190 1952 2196 1953
rect 2190 1948 2191 1952
rect 2195 1948 2196 1952
rect 2190 1947 2196 1948
rect 2254 1952 2260 1953
rect 2254 1948 2255 1952
rect 2259 1948 2260 1952
rect 2254 1947 2260 1948
rect 2318 1952 2324 1953
rect 2318 1948 2319 1952
rect 2323 1948 2324 1952
rect 2318 1947 2324 1948
rect 2358 1952 2364 1953
rect 2358 1948 2359 1952
rect 2363 1948 2364 1952
rect 2358 1947 2364 1948
rect 2408 1947 2410 1954
rect 1279 1946 1283 1947
rect 1279 1941 1283 1942
rect 1303 1946 1307 1947
rect 1303 1941 1307 1942
rect 1351 1946 1355 1947
rect 1351 1941 1355 1942
rect 1359 1946 1363 1947
rect 1359 1941 1363 1942
rect 1423 1946 1427 1947
rect 1423 1941 1427 1942
rect 1447 1946 1451 1947
rect 1447 1941 1451 1942
rect 1495 1946 1499 1947
rect 1495 1941 1499 1942
rect 1535 1946 1539 1947
rect 1535 1941 1539 1942
rect 1575 1946 1579 1947
rect 1575 1941 1579 1942
rect 1623 1946 1627 1947
rect 1623 1941 1627 1942
rect 1663 1946 1667 1947
rect 1663 1941 1667 1942
rect 1711 1946 1715 1947
rect 1711 1941 1715 1942
rect 1751 1946 1755 1947
rect 1751 1941 1755 1942
rect 1791 1946 1795 1947
rect 1791 1941 1795 1942
rect 1839 1946 1843 1947
rect 1839 1941 1843 1942
rect 1863 1946 1867 1947
rect 1863 1941 1867 1942
rect 1919 1946 1923 1947
rect 1919 1941 1923 1942
rect 1935 1946 1939 1947
rect 1935 1941 1939 1942
rect 1999 1946 2003 1947
rect 1999 1941 2003 1942
rect 2007 1946 2011 1947
rect 2007 1941 2011 1942
rect 2071 1946 2075 1947
rect 2071 1941 2075 1942
rect 2079 1946 2083 1947
rect 2079 1941 2083 1942
rect 2135 1946 2139 1947
rect 2135 1941 2139 1942
rect 2151 1946 2155 1947
rect 2151 1941 2155 1942
rect 2191 1946 2195 1947
rect 2191 1941 2195 1942
rect 2223 1946 2227 1947
rect 2223 1941 2227 1942
rect 2255 1946 2259 1947
rect 2255 1941 2259 1942
rect 2303 1946 2307 1947
rect 2303 1941 2307 1942
rect 2319 1946 2323 1947
rect 2319 1941 2323 1942
rect 2359 1946 2363 1947
rect 2359 1941 2363 1942
rect 2407 1946 2411 1947
rect 2407 1941 2411 1942
rect 1280 1934 1282 1941
rect 1302 1940 1308 1941
rect 1302 1936 1303 1940
rect 1307 1936 1308 1940
rect 1302 1935 1308 1936
rect 1358 1940 1364 1941
rect 1358 1936 1359 1940
rect 1363 1936 1364 1940
rect 1358 1935 1364 1936
rect 1446 1940 1452 1941
rect 1446 1936 1447 1940
rect 1451 1936 1452 1940
rect 1446 1935 1452 1936
rect 1534 1940 1540 1941
rect 1534 1936 1535 1940
rect 1539 1936 1540 1940
rect 1534 1935 1540 1936
rect 1622 1940 1628 1941
rect 1622 1936 1623 1940
rect 1627 1936 1628 1940
rect 1622 1935 1628 1936
rect 1710 1940 1716 1941
rect 1710 1936 1711 1940
rect 1715 1936 1716 1940
rect 1710 1935 1716 1936
rect 1790 1940 1796 1941
rect 1790 1936 1791 1940
rect 1795 1936 1796 1940
rect 1790 1935 1796 1936
rect 1862 1940 1868 1941
rect 1862 1936 1863 1940
rect 1867 1936 1868 1940
rect 1862 1935 1868 1936
rect 1934 1940 1940 1941
rect 1934 1936 1935 1940
rect 1939 1936 1940 1940
rect 1934 1935 1940 1936
rect 2006 1940 2012 1941
rect 2006 1936 2007 1940
rect 2011 1936 2012 1940
rect 2006 1935 2012 1936
rect 2078 1940 2084 1941
rect 2078 1936 2079 1940
rect 2083 1936 2084 1940
rect 2078 1935 2084 1936
rect 2150 1940 2156 1941
rect 2150 1936 2151 1940
rect 2155 1936 2156 1940
rect 2150 1935 2156 1936
rect 2222 1940 2228 1941
rect 2222 1936 2223 1940
rect 2227 1936 2228 1940
rect 2222 1935 2228 1936
rect 2302 1940 2308 1941
rect 2302 1936 2303 1940
rect 2307 1936 2308 1940
rect 2302 1935 2308 1936
rect 2358 1940 2364 1941
rect 2358 1936 2359 1940
rect 2363 1936 2364 1940
rect 2358 1935 2364 1936
rect 2408 1934 2410 1941
rect 1278 1933 1284 1934
rect 1278 1929 1279 1933
rect 1283 1929 1284 1933
rect 1278 1928 1284 1929
rect 2406 1933 2412 1934
rect 2406 1929 2407 1933
rect 2411 1929 2412 1933
rect 2406 1928 2412 1929
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 175 1926 179 1927
rect 175 1921 179 1922
rect 215 1926 219 1927
rect 215 1921 219 1922
rect 263 1926 267 1927
rect 263 1921 267 1922
rect 319 1926 323 1927
rect 319 1921 323 1922
rect 367 1926 371 1927
rect 367 1921 371 1922
rect 391 1926 395 1927
rect 391 1921 395 1922
rect 407 1926 411 1927
rect 407 1921 411 1922
rect 455 1926 459 1927
rect 455 1921 459 1922
rect 471 1926 475 1927
rect 471 1921 475 1922
rect 511 1926 515 1927
rect 511 1921 515 1922
rect 551 1926 555 1927
rect 551 1921 555 1922
rect 567 1926 571 1927
rect 567 1921 571 1922
rect 631 1926 635 1927
rect 631 1921 635 1922
rect 639 1926 643 1927
rect 639 1921 643 1922
rect 695 1926 699 1927
rect 695 1921 699 1922
rect 719 1926 723 1927
rect 719 1921 723 1922
rect 759 1926 763 1927
rect 759 1921 763 1922
rect 799 1926 803 1927
rect 799 1921 803 1922
rect 815 1926 819 1927
rect 815 1921 819 1922
rect 871 1926 875 1927
rect 871 1921 875 1922
rect 879 1926 883 1927
rect 879 1921 883 1922
rect 935 1926 939 1927
rect 935 1921 939 1922
rect 959 1926 963 1927
rect 959 1921 963 1922
rect 999 1926 1003 1927
rect 999 1921 1003 1922
rect 1039 1926 1043 1927
rect 1039 1921 1043 1922
rect 1063 1926 1067 1927
rect 1063 1921 1067 1922
rect 1119 1926 1123 1927
rect 1119 1921 1123 1922
rect 1239 1926 1243 1927
rect 1239 1921 1243 1922
rect 112 1889 114 1921
rect 176 1912 178 1921
rect 216 1912 218 1921
rect 264 1912 266 1921
rect 320 1912 322 1921
rect 392 1912 394 1921
rect 472 1912 474 1921
rect 552 1912 554 1921
rect 640 1912 642 1921
rect 720 1912 722 1921
rect 800 1912 802 1921
rect 880 1912 882 1921
rect 960 1912 962 1921
rect 1040 1912 1042 1921
rect 1120 1912 1122 1921
rect 174 1911 180 1912
rect 174 1907 175 1911
rect 179 1907 180 1911
rect 174 1906 180 1907
rect 214 1911 220 1912
rect 214 1907 215 1911
rect 219 1907 220 1911
rect 214 1906 220 1907
rect 262 1911 268 1912
rect 262 1907 263 1911
rect 267 1907 268 1911
rect 262 1906 268 1907
rect 318 1911 324 1912
rect 318 1907 319 1911
rect 323 1907 324 1911
rect 318 1906 324 1907
rect 390 1911 396 1912
rect 390 1907 391 1911
rect 395 1907 396 1911
rect 390 1906 396 1907
rect 470 1911 476 1912
rect 470 1907 471 1911
rect 475 1907 476 1911
rect 470 1906 476 1907
rect 550 1911 556 1912
rect 550 1907 551 1911
rect 555 1907 556 1911
rect 550 1906 556 1907
rect 638 1911 644 1912
rect 638 1907 639 1911
rect 643 1907 644 1911
rect 638 1906 644 1907
rect 718 1911 724 1912
rect 718 1907 719 1911
rect 723 1907 724 1911
rect 718 1906 724 1907
rect 798 1911 804 1912
rect 798 1907 799 1911
rect 803 1907 804 1911
rect 798 1906 804 1907
rect 878 1911 884 1912
rect 878 1907 879 1911
rect 883 1907 884 1911
rect 878 1906 884 1907
rect 958 1911 964 1912
rect 958 1907 959 1911
rect 963 1907 964 1911
rect 958 1906 964 1907
rect 1038 1911 1044 1912
rect 1038 1907 1039 1911
rect 1043 1907 1044 1911
rect 1038 1906 1044 1907
rect 1118 1911 1124 1912
rect 1118 1907 1119 1911
rect 1123 1907 1124 1911
rect 1118 1906 1124 1907
rect 1240 1889 1242 1921
rect 1278 1916 1284 1917
rect 1278 1912 1279 1916
rect 1283 1912 1284 1916
rect 1278 1911 1284 1912
rect 2406 1916 2412 1917
rect 2406 1912 2407 1916
rect 2411 1912 2412 1916
rect 2406 1911 2412 1912
rect 110 1888 116 1889
rect 110 1884 111 1888
rect 115 1884 116 1888
rect 110 1883 116 1884
rect 1238 1888 1244 1889
rect 1238 1884 1239 1888
rect 1243 1884 1244 1888
rect 1238 1883 1244 1884
rect 1280 1879 1282 1911
rect 1302 1893 1308 1894
rect 1302 1889 1303 1893
rect 1307 1889 1308 1893
rect 1302 1888 1308 1889
rect 1358 1893 1364 1894
rect 1358 1889 1359 1893
rect 1363 1889 1364 1893
rect 1358 1888 1364 1889
rect 1446 1893 1452 1894
rect 1446 1889 1447 1893
rect 1451 1889 1452 1893
rect 1446 1888 1452 1889
rect 1534 1893 1540 1894
rect 1534 1889 1535 1893
rect 1539 1889 1540 1893
rect 1534 1888 1540 1889
rect 1622 1893 1628 1894
rect 1622 1889 1623 1893
rect 1627 1889 1628 1893
rect 1622 1888 1628 1889
rect 1710 1893 1716 1894
rect 1710 1889 1711 1893
rect 1715 1889 1716 1893
rect 1710 1888 1716 1889
rect 1790 1893 1796 1894
rect 1790 1889 1791 1893
rect 1795 1889 1796 1893
rect 1790 1888 1796 1889
rect 1862 1893 1868 1894
rect 1862 1889 1863 1893
rect 1867 1889 1868 1893
rect 1862 1888 1868 1889
rect 1934 1893 1940 1894
rect 1934 1889 1935 1893
rect 1939 1889 1940 1893
rect 1934 1888 1940 1889
rect 2006 1893 2012 1894
rect 2006 1889 2007 1893
rect 2011 1889 2012 1893
rect 2006 1888 2012 1889
rect 2078 1893 2084 1894
rect 2078 1889 2079 1893
rect 2083 1889 2084 1893
rect 2078 1888 2084 1889
rect 2150 1893 2156 1894
rect 2150 1889 2151 1893
rect 2155 1889 2156 1893
rect 2150 1888 2156 1889
rect 2222 1893 2228 1894
rect 2222 1889 2223 1893
rect 2227 1889 2228 1893
rect 2222 1888 2228 1889
rect 2302 1893 2308 1894
rect 2302 1889 2303 1893
rect 2307 1889 2308 1893
rect 2302 1888 2308 1889
rect 2358 1893 2364 1894
rect 2358 1889 2359 1893
rect 2363 1889 2364 1893
rect 2358 1888 2364 1889
rect 1304 1879 1306 1888
rect 1360 1879 1362 1888
rect 1448 1879 1450 1888
rect 1536 1879 1538 1888
rect 1624 1879 1626 1888
rect 1712 1879 1714 1888
rect 1792 1879 1794 1888
rect 1864 1879 1866 1888
rect 1936 1879 1938 1888
rect 2008 1879 2010 1888
rect 2080 1879 2082 1888
rect 2152 1879 2154 1888
rect 2224 1879 2226 1888
rect 2304 1879 2306 1888
rect 2360 1879 2362 1888
rect 2408 1879 2410 1911
rect 1279 1878 1283 1879
rect 1279 1873 1283 1874
rect 1303 1878 1307 1879
rect 1303 1873 1307 1874
rect 1311 1878 1315 1879
rect 1311 1873 1315 1874
rect 1359 1878 1363 1879
rect 1359 1873 1363 1874
rect 1415 1878 1419 1879
rect 1415 1873 1419 1874
rect 1447 1878 1451 1879
rect 1447 1873 1451 1874
rect 1479 1878 1483 1879
rect 1479 1873 1483 1874
rect 1535 1878 1539 1879
rect 1535 1873 1539 1874
rect 1543 1878 1547 1879
rect 1543 1873 1547 1874
rect 1615 1878 1619 1879
rect 1615 1873 1619 1874
rect 1623 1878 1627 1879
rect 1623 1873 1627 1874
rect 1687 1878 1691 1879
rect 1687 1873 1691 1874
rect 1711 1878 1715 1879
rect 1711 1873 1715 1874
rect 1767 1878 1771 1879
rect 1767 1873 1771 1874
rect 1791 1878 1795 1879
rect 1791 1873 1795 1874
rect 1863 1878 1867 1879
rect 1863 1873 1867 1874
rect 1935 1878 1939 1879
rect 1935 1873 1939 1874
rect 1975 1878 1979 1879
rect 1975 1873 1979 1874
rect 2007 1878 2011 1879
rect 2007 1873 2011 1874
rect 2079 1878 2083 1879
rect 2079 1873 2083 1874
rect 2095 1878 2099 1879
rect 2095 1873 2099 1874
rect 2151 1878 2155 1879
rect 2151 1873 2155 1874
rect 2223 1878 2227 1879
rect 2223 1873 2227 1874
rect 2303 1878 2307 1879
rect 2303 1873 2307 1874
rect 2359 1878 2363 1879
rect 2359 1873 2363 1874
rect 2407 1878 2411 1879
rect 2407 1873 2411 1874
rect 110 1871 116 1872
rect 110 1867 111 1871
rect 115 1867 116 1871
rect 110 1866 116 1867
rect 1238 1871 1244 1872
rect 1238 1867 1239 1871
rect 1243 1867 1244 1871
rect 1238 1866 1244 1867
rect 112 1851 114 1866
rect 174 1864 180 1865
rect 174 1860 175 1864
rect 179 1860 180 1864
rect 174 1859 180 1860
rect 214 1864 220 1865
rect 214 1860 215 1864
rect 219 1860 220 1864
rect 214 1859 220 1860
rect 262 1864 268 1865
rect 262 1860 263 1864
rect 267 1860 268 1864
rect 262 1859 268 1860
rect 318 1864 324 1865
rect 318 1860 319 1864
rect 323 1860 324 1864
rect 318 1859 324 1860
rect 390 1864 396 1865
rect 390 1860 391 1864
rect 395 1860 396 1864
rect 390 1859 396 1860
rect 470 1864 476 1865
rect 470 1860 471 1864
rect 475 1860 476 1864
rect 470 1859 476 1860
rect 550 1864 556 1865
rect 550 1860 551 1864
rect 555 1860 556 1864
rect 550 1859 556 1860
rect 638 1864 644 1865
rect 638 1860 639 1864
rect 643 1860 644 1864
rect 638 1859 644 1860
rect 718 1864 724 1865
rect 718 1860 719 1864
rect 723 1860 724 1864
rect 718 1859 724 1860
rect 798 1864 804 1865
rect 798 1860 799 1864
rect 803 1860 804 1864
rect 798 1859 804 1860
rect 878 1864 884 1865
rect 878 1860 879 1864
rect 883 1860 884 1864
rect 878 1859 884 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1038 1864 1044 1865
rect 1038 1860 1039 1864
rect 1043 1860 1044 1864
rect 1038 1859 1044 1860
rect 1118 1864 1124 1865
rect 1118 1860 1119 1864
rect 1123 1860 1124 1864
rect 1118 1859 1124 1860
rect 176 1851 178 1859
rect 216 1851 218 1859
rect 264 1851 266 1859
rect 320 1851 322 1859
rect 392 1851 394 1859
rect 472 1851 474 1859
rect 552 1851 554 1859
rect 640 1851 642 1859
rect 720 1851 722 1859
rect 800 1851 802 1859
rect 880 1851 882 1859
rect 960 1851 962 1859
rect 1040 1851 1042 1859
rect 1120 1851 1122 1859
rect 1240 1851 1242 1866
rect 111 1850 115 1851
rect 111 1845 115 1846
rect 135 1850 139 1851
rect 135 1845 139 1846
rect 175 1850 179 1851
rect 175 1845 179 1846
rect 215 1850 219 1851
rect 215 1845 219 1846
rect 263 1850 267 1851
rect 263 1845 267 1846
rect 271 1850 275 1851
rect 271 1845 275 1846
rect 319 1850 323 1851
rect 319 1845 323 1846
rect 351 1850 355 1851
rect 351 1845 355 1846
rect 391 1850 395 1851
rect 391 1845 395 1846
rect 439 1850 443 1851
rect 439 1845 443 1846
rect 471 1850 475 1851
rect 471 1845 475 1846
rect 535 1850 539 1851
rect 535 1845 539 1846
rect 551 1850 555 1851
rect 551 1845 555 1846
rect 631 1850 635 1851
rect 631 1845 635 1846
rect 639 1850 643 1851
rect 639 1845 643 1846
rect 719 1850 723 1851
rect 719 1845 723 1846
rect 727 1850 731 1851
rect 727 1845 731 1846
rect 799 1850 803 1851
rect 799 1845 803 1846
rect 823 1850 827 1851
rect 823 1845 827 1846
rect 879 1850 883 1851
rect 879 1845 883 1846
rect 911 1850 915 1851
rect 911 1845 915 1846
rect 959 1850 963 1851
rect 959 1845 963 1846
rect 991 1850 995 1851
rect 991 1845 995 1846
rect 1039 1850 1043 1851
rect 1039 1845 1043 1846
rect 1063 1850 1067 1851
rect 1063 1845 1067 1846
rect 1119 1850 1123 1851
rect 1119 1845 1123 1846
rect 1135 1850 1139 1851
rect 1135 1845 1139 1846
rect 1191 1850 1195 1851
rect 1191 1845 1195 1846
rect 1239 1850 1243 1851
rect 1239 1845 1243 1846
rect 112 1838 114 1845
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 214 1844 220 1845
rect 214 1840 215 1844
rect 219 1840 220 1844
rect 214 1839 220 1840
rect 270 1844 276 1845
rect 270 1840 271 1844
rect 275 1840 276 1844
rect 270 1839 276 1840
rect 350 1844 356 1845
rect 350 1840 351 1844
rect 355 1840 356 1844
rect 350 1839 356 1840
rect 438 1844 444 1845
rect 438 1840 439 1844
rect 443 1840 444 1844
rect 438 1839 444 1840
rect 534 1844 540 1845
rect 534 1840 535 1844
rect 539 1840 540 1844
rect 534 1839 540 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 726 1844 732 1845
rect 726 1840 727 1844
rect 731 1840 732 1844
rect 726 1839 732 1840
rect 822 1844 828 1845
rect 822 1840 823 1844
rect 827 1840 828 1844
rect 822 1839 828 1840
rect 910 1844 916 1845
rect 910 1840 911 1844
rect 915 1840 916 1844
rect 910 1839 916 1840
rect 990 1844 996 1845
rect 990 1840 991 1844
rect 995 1840 996 1844
rect 990 1839 996 1840
rect 1062 1844 1068 1845
rect 1062 1840 1063 1844
rect 1067 1840 1068 1844
rect 1062 1839 1068 1840
rect 1134 1844 1140 1845
rect 1134 1840 1135 1844
rect 1139 1840 1140 1844
rect 1134 1839 1140 1840
rect 1190 1844 1196 1845
rect 1190 1840 1191 1844
rect 1195 1840 1196 1844
rect 1190 1839 1196 1840
rect 1240 1838 1242 1845
rect 1280 1841 1282 1873
rect 1312 1864 1314 1873
rect 1360 1864 1362 1873
rect 1416 1864 1418 1873
rect 1480 1864 1482 1873
rect 1544 1864 1546 1873
rect 1616 1864 1618 1873
rect 1688 1864 1690 1873
rect 1768 1864 1770 1873
rect 1864 1864 1866 1873
rect 1976 1864 1978 1873
rect 2096 1864 2098 1873
rect 2224 1864 2226 1873
rect 2360 1864 2362 1873
rect 1310 1863 1316 1864
rect 1310 1859 1311 1863
rect 1315 1859 1316 1863
rect 1310 1858 1316 1859
rect 1358 1863 1364 1864
rect 1358 1859 1359 1863
rect 1363 1859 1364 1863
rect 1358 1858 1364 1859
rect 1414 1863 1420 1864
rect 1414 1859 1415 1863
rect 1419 1859 1420 1863
rect 1414 1858 1420 1859
rect 1478 1863 1484 1864
rect 1478 1859 1479 1863
rect 1483 1859 1484 1863
rect 1478 1858 1484 1859
rect 1542 1863 1548 1864
rect 1542 1859 1543 1863
rect 1547 1859 1548 1863
rect 1542 1858 1548 1859
rect 1614 1863 1620 1864
rect 1614 1859 1615 1863
rect 1619 1859 1620 1863
rect 1614 1858 1620 1859
rect 1686 1863 1692 1864
rect 1686 1859 1687 1863
rect 1691 1859 1692 1863
rect 1686 1858 1692 1859
rect 1766 1863 1772 1864
rect 1766 1859 1767 1863
rect 1771 1859 1772 1863
rect 1766 1858 1772 1859
rect 1862 1863 1868 1864
rect 1862 1859 1863 1863
rect 1867 1859 1868 1863
rect 1862 1858 1868 1859
rect 1974 1863 1980 1864
rect 1974 1859 1975 1863
rect 1979 1859 1980 1863
rect 1974 1858 1980 1859
rect 2094 1863 2100 1864
rect 2094 1859 2095 1863
rect 2099 1859 2100 1863
rect 2094 1858 2100 1859
rect 2222 1863 2228 1864
rect 2222 1859 2223 1863
rect 2227 1859 2228 1863
rect 2222 1858 2228 1859
rect 2358 1863 2364 1864
rect 2358 1859 2359 1863
rect 2363 1859 2364 1863
rect 2358 1858 2364 1859
rect 2408 1841 2410 1873
rect 1278 1840 1284 1841
rect 110 1837 116 1838
rect 110 1833 111 1837
rect 115 1833 116 1837
rect 110 1832 116 1833
rect 1238 1837 1244 1838
rect 1238 1833 1239 1837
rect 1243 1833 1244 1837
rect 1278 1836 1279 1840
rect 1283 1836 1284 1840
rect 1278 1835 1284 1836
rect 2406 1840 2412 1841
rect 2406 1836 2407 1840
rect 2411 1836 2412 1840
rect 2406 1835 2412 1836
rect 1238 1832 1244 1833
rect 1278 1823 1284 1824
rect 110 1820 116 1821
rect 110 1816 111 1820
rect 115 1816 116 1820
rect 110 1815 116 1816
rect 1238 1820 1244 1821
rect 1238 1816 1239 1820
rect 1243 1816 1244 1820
rect 1278 1819 1279 1823
rect 1283 1819 1284 1823
rect 1278 1818 1284 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 1238 1815 1244 1816
rect 112 1783 114 1815
rect 134 1797 140 1798
rect 134 1793 135 1797
rect 139 1793 140 1797
rect 134 1792 140 1793
rect 174 1797 180 1798
rect 174 1793 175 1797
rect 179 1793 180 1797
rect 174 1792 180 1793
rect 214 1797 220 1798
rect 214 1793 215 1797
rect 219 1793 220 1797
rect 214 1792 220 1793
rect 270 1797 276 1798
rect 270 1793 271 1797
rect 275 1793 276 1797
rect 270 1792 276 1793
rect 350 1797 356 1798
rect 350 1793 351 1797
rect 355 1793 356 1797
rect 350 1792 356 1793
rect 438 1797 444 1798
rect 438 1793 439 1797
rect 443 1793 444 1797
rect 438 1792 444 1793
rect 534 1797 540 1798
rect 534 1793 535 1797
rect 539 1793 540 1797
rect 534 1792 540 1793
rect 630 1797 636 1798
rect 630 1793 631 1797
rect 635 1793 636 1797
rect 630 1792 636 1793
rect 726 1797 732 1798
rect 726 1793 727 1797
rect 731 1793 732 1797
rect 726 1792 732 1793
rect 822 1797 828 1798
rect 822 1793 823 1797
rect 827 1793 828 1797
rect 822 1792 828 1793
rect 910 1797 916 1798
rect 910 1793 911 1797
rect 915 1793 916 1797
rect 910 1792 916 1793
rect 990 1797 996 1798
rect 990 1793 991 1797
rect 995 1793 996 1797
rect 990 1792 996 1793
rect 1062 1797 1068 1798
rect 1062 1793 1063 1797
rect 1067 1793 1068 1797
rect 1062 1792 1068 1793
rect 1134 1797 1140 1798
rect 1134 1793 1135 1797
rect 1139 1793 1140 1797
rect 1134 1792 1140 1793
rect 1190 1797 1196 1798
rect 1190 1793 1191 1797
rect 1195 1793 1196 1797
rect 1190 1792 1196 1793
rect 136 1783 138 1792
rect 176 1783 178 1792
rect 216 1783 218 1792
rect 272 1783 274 1792
rect 352 1783 354 1792
rect 440 1783 442 1792
rect 536 1783 538 1792
rect 632 1783 634 1792
rect 728 1783 730 1792
rect 824 1783 826 1792
rect 912 1783 914 1792
rect 992 1783 994 1792
rect 1064 1783 1066 1792
rect 1136 1783 1138 1792
rect 1192 1783 1194 1792
rect 1240 1783 1242 1815
rect 1280 1807 1282 1818
rect 1310 1816 1316 1817
rect 1310 1812 1311 1816
rect 1315 1812 1316 1816
rect 1310 1811 1316 1812
rect 1358 1816 1364 1817
rect 1358 1812 1359 1816
rect 1363 1812 1364 1816
rect 1358 1811 1364 1812
rect 1414 1816 1420 1817
rect 1414 1812 1415 1816
rect 1419 1812 1420 1816
rect 1414 1811 1420 1812
rect 1478 1816 1484 1817
rect 1478 1812 1479 1816
rect 1483 1812 1484 1816
rect 1478 1811 1484 1812
rect 1542 1816 1548 1817
rect 1542 1812 1543 1816
rect 1547 1812 1548 1816
rect 1542 1811 1548 1812
rect 1614 1816 1620 1817
rect 1614 1812 1615 1816
rect 1619 1812 1620 1816
rect 1614 1811 1620 1812
rect 1686 1816 1692 1817
rect 1686 1812 1687 1816
rect 1691 1812 1692 1816
rect 1686 1811 1692 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1862 1816 1868 1817
rect 1862 1812 1863 1816
rect 1867 1812 1868 1816
rect 1862 1811 1868 1812
rect 1974 1816 1980 1817
rect 1974 1812 1975 1816
rect 1979 1812 1980 1816
rect 1974 1811 1980 1812
rect 2094 1816 2100 1817
rect 2094 1812 2095 1816
rect 2099 1812 2100 1816
rect 2094 1811 2100 1812
rect 2222 1816 2228 1817
rect 2222 1812 2223 1816
rect 2227 1812 2228 1816
rect 2222 1811 2228 1812
rect 2358 1816 2364 1817
rect 2358 1812 2359 1816
rect 2363 1812 2364 1816
rect 2358 1811 2364 1812
rect 1312 1807 1314 1811
rect 1360 1807 1362 1811
rect 1416 1807 1418 1811
rect 1480 1807 1482 1811
rect 1544 1807 1546 1811
rect 1616 1807 1618 1811
rect 1688 1807 1690 1811
rect 1768 1807 1770 1811
rect 1864 1807 1866 1811
rect 1976 1807 1978 1811
rect 2096 1807 2098 1811
rect 2224 1807 2226 1811
rect 2360 1807 2362 1811
rect 2408 1807 2410 1818
rect 1279 1806 1283 1807
rect 1279 1801 1283 1802
rect 1311 1806 1315 1807
rect 1311 1801 1315 1802
rect 1359 1806 1363 1807
rect 1359 1801 1363 1802
rect 1407 1806 1411 1807
rect 1407 1801 1411 1802
rect 1415 1806 1419 1807
rect 1415 1801 1419 1802
rect 1471 1806 1475 1807
rect 1471 1801 1475 1802
rect 1479 1806 1483 1807
rect 1479 1801 1483 1802
rect 1535 1806 1539 1807
rect 1535 1801 1539 1802
rect 1543 1806 1547 1807
rect 1543 1801 1547 1802
rect 1599 1806 1603 1807
rect 1599 1801 1603 1802
rect 1615 1806 1619 1807
rect 1615 1801 1619 1802
rect 1663 1806 1667 1807
rect 1663 1801 1667 1802
rect 1687 1806 1691 1807
rect 1687 1801 1691 1802
rect 1727 1806 1731 1807
rect 1727 1801 1731 1802
rect 1767 1806 1771 1807
rect 1767 1801 1771 1802
rect 1783 1806 1787 1807
rect 1783 1801 1787 1802
rect 1839 1806 1843 1807
rect 1839 1801 1843 1802
rect 1863 1806 1867 1807
rect 1863 1801 1867 1802
rect 1895 1806 1899 1807
rect 1895 1801 1899 1802
rect 1959 1806 1963 1807
rect 1959 1801 1963 1802
rect 1975 1806 1979 1807
rect 1975 1801 1979 1802
rect 2095 1806 2099 1807
rect 2095 1801 2099 1802
rect 2223 1806 2227 1807
rect 2223 1801 2227 1802
rect 2359 1806 2363 1807
rect 2359 1801 2363 1802
rect 2407 1806 2411 1807
rect 2407 1801 2411 1802
rect 1280 1794 1282 1801
rect 1406 1800 1412 1801
rect 1406 1796 1407 1800
rect 1411 1796 1412 1800
rect 1406 1795 1412 1796
rect 1470 1800 1476 1801
rect 1470 1796 1471 1800
rect 1475 1796 1476 1800
rect 1470 1795 1476 1796
rect 1534 1800 1540 1801
rect 1534 1796 1535 1800
rect 1539 1796 1540 1800
rect 1534 1795 1540 1796
rect 1598 1800 1604 1801
rect 1598 1796 1599 1800
rect 1603 1796 1604 1800
rect 1598 1795 1604 1796
rect 1662 1800 1668 1801
rect 1662 1796 1663 1800
rect 1667 1796 1668 1800
rect 1662 1795 1668 1796
rect 1726 1800 1732 1801
rect 1726 1796 1727 1800
rect 1731 1796 1732 1800
rect 1726 1795 1732 1796
rect 1782 1800 1788 1801
rect 1782 1796 1783 1800
rect 1787 1796 1788 1800
rect 1782 1795 1788 1796
rect 1838 1800 1844 1801
rect 1838 1796 1839 1800
rect 1843 1796 1844 1800
rect 1838 1795 1844 1796
rect 1894 1800 1900 1801
rect 1894 1796 1895 1800
rect 1899 1796 1900 1800
rect 1894 1795 1900 1796
rect 1958 1800 1964 1801
rect 1958 1796 1959 1800
rect 1963 1796 1964 1800
rect 1958 1795 1964 1796
rect 2408 1794 2410 1801
rect 1278 1793 1284 1794
rect 1278 1789 1279 1793
rect 1283 1789 1284 1793
rect 1278 1788 1284 1789
rect 2406 1793 2412 1794
rect 2406 1789 2407 1793
rect 2411 1789 2412 1793
rect 2406 1788 2412 1789
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 135 1782 139 1783
rect 135 1777 139 1778
rect 175 1782 179 1783
rect 175 1777 179 1778
rect 215 1782 219 1783
rect 215 1777 219 1778
rect 271 1782 275 1783
rect 271 1777 275 1778
rect 287 1782 291 1783
rect 287 1777 291 1778
rect 351 1782 355 1783
rect 351 1777 355 1778
rect 375 1782 379 1783
rect 375 1777 379 1778
rect 439 1782 443 1783
rect 439 1777 443 1778
rect 471 1782 475 1783
rect 471 1777 475 1778
rect 535 1782 539 1783
rect 535 1777 539 1778
rect 567 1782 571 1783
rect 567 1777 571 1778
rect 631 1782 635 1783
rect 631 1777 635 1778
rect 663 1782 667 1783
rect 663 1777 667 1778
rect 727 1782 731 1783
rect 727 1777 731 1778
rect 751 1782 755 1783
rect 751 1777 755 1778
rect 823 1782 827 1783
rect 823 1777 827 1778
rect 831 1782 835 1783
rect 831 1777 835 1778
rect 903 1782 907 1783
rect 903 1777 907 1778
rect 911 1782 915 1783
rect 911 1777 915 1778
rect 967 1782 971 1783
rect 967 1777 971 1778
rect 991 1782 995 1783
rect 991 1777 995 1778
rect 1031 1782 1035 1783
rect 1031 1777 1035 1778
rect 1063 1782 1067 1783
rect 1063 1777 1067 1778
rect 1087 1782 1091 1783
rect 1087 1777 1091 1778
rect 1135 1782 1139 1783
rect 1135 1777 1139 1778
rect 1151 1782 1155 1783
rect 1151 1777 1155 1778
rect 1191 1782 1195 1783
rect 1191 1777 1195 1778
rect 1239 1782 1243 1783
rect 1239 1777 1243 1778
rect 112 1745 114 1777
rect 136 1768 138 1777
rect 176 1768 178 1777
rect 216 1768 218 1777
rect 288 1768 290 1777
rect 376 1768 378 1777
rect 472 1768 474 1777
rect 568 1768 570 1777
rect 664 1768 666 1777
rect 752 1768 754 1777
rect 832 1768 834 1777
rect 904 1768 906 1777
rect 968 1768 970 1777
rect 1032 1768 1034 1777
rect 1088 1768 1090 1777
rect 1152 1768 1154 1777
rect 1192 1768 1194 1777
rect 134 1767 140 1768
rect 134 1763 135 1767
rect 139 1763 140 1767
rect 134 1762 140 1763
rect 174 1767 180 1768
rect 174 1763 175 1767
rect 179 1763 180 1767
rect 174 1762 180 1763
rect 214 1767 220 1768
rect 214 1763 215 1767
rect 219 1763 220 1767
rect 214 1762 220 1763
rect 286 1767 292 1768
rect 286 1763 287 1767
rect 291 1763 292 1767
rect 286 1762 292 1763
rect 374 1767 380 1768
rect 374 1763 375 1767
rect 379 1763 380 1767
rect 374 1762 380 1763
rect 470 1767 476 1768
rect 470 1763 471 1767
rect 475 1763 476 1767
rect 470 1762 476 1763
rect 566 1767 572 1768
rect 566 1763 567 1767
rect 571 1763 572 1767
rect 566 1762 572 1763
rect 662 1767 668 1768
rect 662 1763 663 1767
rect 667 1763 668 1767
rect 662 1762 668 1763
rect 750 1767 756 1768
rect 750 1763 751 1767
rect 755 1763 756 1767
rect 750 1762 756 1763
rect 830 1767 836 1768
rect 830 1763 831 1767
rect 835 1763 836 1767
rect 830 1762 836 1763
rect 902 1767 908 1768
rect 902 1763 903 1767
rect 907 1763 908 1767
rect 902 1762 908 1763
rect 966 1767 972 1768
rect 966 1763 967 1767
rect 971 1763 972 1767
rect 966 1762 972 1763
rect 1030 1767 1036 1768
rect 1030 1763 1031 1767
rect 1035 1763 1036 1767
rect 1030 1762 1036 1763
rect 1086 1767 1092 1768
rect 1086 1763 1087 1767
rect 1091 1763 1092 1767
rect 1086 1762 1092 1763
rect 1150 1767 1156 1768
rect 1150 1763 1151 1767
rect 1155 1763 1156 1767
rect 1150 1762 1156 1763
rect 1190 1767 1196 1768
rect 1190 1763 1191 1767
rect 1195 1763 1196 1767
rect 1190 1762 1196 1763
rect 1240 1745 1242 1777
rect 1278 1776 1284 1777
rect 1278 1772 1279 1776
rect 1283 1772 1284 1776
rect 1278 1771 1284 1772
rect 2406 1776 2412 1777
rect 2406 1772 2407 1776
rect 2411 1772 2412 1776
rect 2406 1771 2412 1772
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 110 1739 116 1740
rect 1238 1744 1244 1745
rect 1238 1740 1239 1744
rect 1243 1740 1244 1744
rect 1238 1739 1244 1740
rect 1280 1739 1282 1771
rect 1406 1753 1412 1754
rect 1406 1749 1407 1753
rect 1411 1749 1412 1753
rect 1406 1748 1412 1749
rect 1470 1753 1476 1754
rect 1470 1749 1471 1753
rect 1475 1749 1476 1753
rect 1470 1748 1476 1749
rect 1534 1753 1540 1754
rect 1534 1749 1535 1753
rect 1539 1749 1540 1753
rect 1534 1748 1540 1749
rect 1598 1753 1604 1754
rect 1598 1749 1599 1753
rect 1603 1749 1604 1753
rect 1598 1748 1604 1749
rect 1662 1753 1668 1754
rect 1662 1749 1663 1753
rect 1667 1749 1668 1753
rect 1662 1748 1668 1749
rect 1726 1753 1732 1754
rect 1726 1749 1727 1753
rect 1731 1749 1732 1753
rect 1726 1748 1732 1749
rect 1782 1753 1788 1754
rect 1782 1749 1783 1753
rect 1787 1749 1788 1753
rect 1782 1748 1788 1749
rect 1838 1753 1844 1754
rect 1838 1749 1839 1753
rect 1843 1749 1844 1753
rect 1838 1748 1844 1749
rect 1894 1753 1900 1754
rect 1894 1749 1895 1753
rect 1899 1749 1900 1753
rect 1894 1748 1900 1749
rect 1958 1753 1964 1754
rect 1958 1749 1959 1753
rect 1963 1749 1964 1753
rect 1958 1748 1964 1749
rect 1408 1739 1410 1748
rect 1472 1739 1474 1748
rect 1536 1739 1538 1748
rect 1600 1739 1602 1748
rect 1664 1739 1666 1748
rect 1728 1739 1730 1748
rect 1784 1739 1786 1748
rect 1840 1739 1842 1748
rect 1896 1739 1898 1748
rect 1960 1739 1962 1748
rect 2408 1739 2410 1771
rect 1279 1738 1283 1739
rect 1279 1733 1283 1734
rect 1303 1738 1307 1739
rect 1303 1733 1307 1734
rect 1351 1738 1355 1739
rect 1351 1733 1355 1734
rect 1407 1738 1411 1739
rect 1407 1733 1411 1734
rect 1423 1738 1427 1739
rect 1423 1733 1427 1734
rect 1471 1738 1475 1739
rect 1471 1733 1475 1734
rect 1503 1738 1507 1739
rect 1503 1733 1507 1734
rect 1535 1738 1539 1739
rect 1535 1733 1539 1734
rect 1583 1738 1587 1739
rect 1583 1733 1587 1734
rect 1599 1738 1603 1739
rect 1599 1733 1603 1734
rect 1663 1738 1667 1739
rect 1663 1733 1667 1734
rect 1727 1738 1731 1739
rect 1727 1733 1731 1734
rect 1735 1738 1739 1739
rect 1735 1733 1739 1734
rect 1783 1738 1787 1739
rect 1783 1733 1787 1734
rect 1807 1738 1811 1739
rect 1807 1733 1811 1734
rect 1839 1738 1843 1739
rect 1839 1733 1843 1734
rect 1871 1738 1875 1739
rect 1871 1733 1875 1734
rect 1895 1738 1899 1739
rect 1895 1733 1899 1734
rect 1935 1738 1939 1739
rect 1935 1733 1939 1734
rect 1959 1738 1963 1739
rect 1959 1733 1963 1734
rect 1999 1738 2003 1739
rect 1999 1733 2003 1734
rect 2063 1738 2067 1739
rect 2063 1733 2067 1734
rect 2407 1738 2411 1739
rect 2407 1733 2411 1734
rect 110 1727 116 1728
rect 110 1723 111 1727
rect 115 1723 116 1727
rect 110 1722 116 1723
rect 1238 1727 1244 1728
rect 1238 1723 1239 1727
rect 1243 1723 1244 1727
rect 1238 1722 1244 1723
rect 112 1711 114 1722
rect 134 1720 140 1721
rect 134 1716 135 1720
rect 139 1716 140 1720
rect 134 1715 140 1716
rect 174 1720 180 1721
rect 174 1716 175 1720
rect 179 1716 180 1720
rect 174 1715 180 1716
rect 214 1720 220 1721
rect 214 1716 215 1720
rect 219 1716 220 1720
rect 214 1715 220 1716
rect 286 1720 292 1721
rect 286 1716 287 1720
rect 291 1716 292 1720
rect 286 1715 292 1716
rect 374 1720 380 1721
rect 374 1716 375 1720
rect 379 1716 380 1720
rect 374 1715 380 1716
rect 470 1720 476 1721
rect 470 1716 471 1720
rect 475 1716 476 1720
rect 470 1715 476 1716
rect 566 1720 572 1721
rect 566 1716 567 1720
rect 571 1716 572 1720
rect 566 1715 572 1716
rect 662 1720 668 1721
rect 662 1716 663 1720
rect 667 1716 668 1720
rect 662 1715 668 1716
rect 750 1720 756 1721
rect 750 1716 751 1720
rect 755 1716 756 1720
rect 750 1715 756 1716
rect 830 1720 836 1721
rect 830 1716 831 1720
rect 835 1716 836 1720
rect 830 1715 836 1716
rect 902 1720 908 1721
rect 902 1716 903 1720
rect 907 1716 908 1720
rect 902 1715 908 1716
rect 966 1720 972 1721
rect 966 1716 967 1720
rect 971 1716 972 1720
rect 966 1715 972 1716
rect 1030 1720 1036 1721
rect 1030 1716 1031 1720
rect 1035 1716 1036 1720
rect 1030 1715 1036 1716
rect 1086 1720 1092 1721
rect 1086 1716 1087 1720
rect 1091 1716 1092 1720
rect 1086 1715 1092 1716
rect 1150 1720 1156 1721
rect 1150 1716 1151 1720
rect 1155 1716 1156 1720
rect 1150 1715 1156 1716
rect 1190 1720 1196 1721
rect 1190 1716 1191 1720
rect 1195 1716 1196 1720
rect 1190 1715 1196 1716
rect 136 1711 138 1715
rect 176 1711 178 1715
rect 216 1711 218 1715
rect 288 1711 290 1715
rect 376 1711 378 1715
rect 472 1711 474 1715
rect 568 1711 570 1715
rect 664 1711 666 1715
rect 752 1711 754 1715
rect 832 1711 834 1715
rect 904 1711 906 1715
rect 968 1711 970 1715
rect 1032 1711 1034 1715
rect 1088 1711 1090 1715
rect 1152 1711 1154 1715
rect 1192 1711 1194 1715
rect 1240 1711 1242 1722
rect 111 1710 115 1711
rect 111 1705 115 1706
rect 135 1710 139 1711
rect 135 1705 139 1706
rect 175 1710 179 1711
rect 175 1705 179 1706
rect 215 1710 219 1711
rect 215 1705 219 1706
rect 239 1710 243 1711
rect 239 1705 243 1706
rect 287 1710 291 1711
rect 287 1705 291 1706
rect 319 1710 323 1711
rect 319 1705 323 1706
rect 375 1710 379 1711
rect 375 1705 379 1706
rect 415 1710 419 1711
rect 415 1705 419 1706
rect 471 1710 475 1711
rect 471 1705 475 1706
rect 511 1710 515 1711
rect 511 1705 515 1706
rect 567 1710 571 1711
rect 567 1705 571 1706
rect 615 1710 619 1711
rect 615 1705 619 1706
rect 663 1710 667 1711
rect 663 1705 667 1706
rect 711 1710 715 1711
rect 711 1705 715 1706
rect 751 1710 755 1711
rect 751 1705 755 1706
rect 799 1710 803 1711
rect 799 1705 803 1706
rect 831 1710 835 1711
rect 831 1705 835 1706
rect 879 1710 883 1711
rect 879 1705 883 1706
rect 903 1710 907 1711
rect 903 1705 907 1706
rect 951 1710 955 1711
rect 951 1705 955 1706
rect 967 1710 971 1711
rect 967 1705 971 1706
rect 1015 1710 1019 1711
rect 1015 1705 1019 1706
rect 1031 1710 1035 1711
rect 1031 1705 1035 1706
rect 1087 1710 1091 1711
rect 1087 1705 1091 1706
rect 1151 1710 1155 1711
rect 1151 1705 1155 1706
rect 1159 1710 1163 1711
rect 1159 1705 1163 1706
rect 1191 1710 1195 1711
rect 1191 1705 1195 1706
rect 1239 1710 1243 1711
rect 1239 1705 1243 1706
rect 112 1698 114 1705
rect 134 1704 140 1705
rect 134 1700 135 1704
rect 139 1700 140 1704
rect 134 1699 140 1700
rect 174 1704 180 1705
rect 174 1700 175 1704
rect 179 1700 180 1704
rect 174 1699 180 1700
rect 238 1704 244 1705
rect 238 1700 239 1704
rect 243 1700 244 1704
rect 238 1699 244 1700
rect 318 1704 324 1705
rect 318 1700 319 1704
rect 323 1700 324 1704
rect 318 1699 324 1700
rect 414 1704 420 1705
rect 414 1700 415 1704
rect 419 1700 420 1704
rect 414 1699 420 1700
rect 510 1704 516 1705
rect 510 1700 511 1704
rect 515 1700 516 1704
rect 510 1699 516 1700
rect 614 1704 620 1705
rect 614 1700 615 1704
rect 619 1700 620 1704
rect 614 1699 620 1700
rect 710 1704 716 1705
rect 710 1700 711 1704
rect 715 1700 716 1704
rect 710 1699 716 1700
rect 798 1704 804 1705
rect 798 1700 799 1704
rect 803 1700 804 1704
rect 798 1699 804 1700
rect 878 1704 884 1705
rect 878 1700 879 1704
rect 883 1700 884 1704
rect 878 1699 884 1700
rect 950 1704 956 1705
rect 950 1700 951 1704
rect 955 1700 956 1704
rect 950 1699 956 1700
rect 1014 1704 1020 1705
rect 1014 1700 1015 1704
rect 1019 1700 1020 1704
rect 1014 1699 1020 1700
rect 1086 1704 1092 1705
rect 1086 1700 1087 1704
rect 1091 1700 1092 1704
rect 1086 1699 1092 1700
rect 1158 1704 1164 1705
rect 1158 1700 1159 1704
rect 1163 1700 1164 1704
rect 1158 1699 1164 1700
rect 1240 1698 1242 1705
rect 1280 1701 1282 1733
rect 1304 1724 1306 1733
rect 1352 1724 1354 1733
rect 1424 1724 1426 1733
rect 1504 1724 1506 1733
rect 1584 1724 1586 1733
rect 1664 1724 1666 1733
rect 1736 1724 1738 1733
rect 1808 1724 1810 1733
rect 1872 1724 1874 1733
rect 1936 1724 1938 1733
rect 2000 1724 2002 1733
rect 2064 1724 2066 1733
rect 1302 1723 1308 1724
rect 1302 1719 1303 1723
rect 1307 1719 1308 1723
rect 1302 1718 1308 1719
rect 1350 1723 1356 1724
rect 1350 1719 1351 1723
rect 1355 1719 1356 1723
rect 1350 1718 1356 1719
rect 1422 1723 1428 1724
rect 1422 1719 1423 1723
rect 1427 1719 1428 1723
rect 1422 1718 1428 1719
rect 1502 1723 1508 1724
rect 1502 1719 1503 1723
rect 1507 1719 1508 1723
rect 1502 1718 1508 1719
rect 1582 1723 1588 1724
rect 1582 1719 1583 1723
rect 1587 1719 1588 1723
rect 1582 1718 1588 1719
rect 1662 1723 1668 1724
rect 1662 1719 1663 1723
rect 1667 1719 1668 1723
rect 1662 1718 1668 1719
rect 1734 1723 1740 1724
rect 1734 1719 1735 1723
rect 1739 1719 1740 1723
rect 1734 1718 1740 1719
rect 1806 1723 1812 1724
rect 1806 1719 1807 1723
rect 1811 1719 1812 1723
rect 1806 1718 1812 1719
rect 1870 1723 1876 1724
rect 1870 1719 1871 1723
rect 1875 1719 1876 1723
rect 1870 1718 1876 1719
rect 1934 1723 1940 1724
rect 1934 1719 1935 1723
rect 1939 1719 1940 1723
rect 1934 1718 1940 1719
rect 1998 1723 2004 1724
rect 1998 1719 1999 1723
rect 2003 1719 2004 1723
rect 1998 1718 2004 1719
rect 2062 1723 2068 1724
rect 2062 1719 2063 1723
rect 2067 1719 2068 1723
rect 2062 1718 2068 1719
rect 2408 1701 2410 1733
rect 1278 1700 1284 1701
rect 110 1697 116 1698
rect 110 1693 111 1697
rect 115 1693 116 1697
rect 110 1692 116 1693
rect 1238 1697 1244 1698
rect 1238 1693 1239 1697
rect 1243 1693 1244 1697
rect 1278 1696 1279 1700
rect 1283 1696 1284 1700
rect 1278 1695 1284 1696
rect 2406 1700 2412 1701
rect 2406 1696 2407 1700
rect 2411 1696 2412 1700
rect 2406 1695 2412 1696
rect 1238 1692 1244 1693
rect 1278 1683 1284 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 110 1675 116 1676
rect 1238 1680 1244 1681
rect 1238 1676 1239 1680
rect 1243 1676 1244 1680
rect 1278 1679 1279 1683
rect 1283 1679 1284 1683
rect 1278 1678 1284 1679
rect 2406 1683 2412 1684
rect 2406 1679 2407 1683
rect 2411 1679 2412 1683
rect 2406 1678 2412 1679
rect 1238 1675 1244 1676
rect 112 1639 114 1675
rect 134 1657 140 1658
rect 134 1653 135 1657
rect 139 1653 140 1657
rect 134 1652 140 1653
rect 174 1657 180 1658
rect 174 1653 175 1657
rect 179 1653 180 1657
rect 174 1652 180 1653
rect 238 1657 244 1658
rect 238 1653 239 1657
rect 243 1653 244 1657
rect 238 1652 244 1653
rect 318 1657 324 1658
rect 318 1653 319 1657
rect 323 1653 324 1657
rect 318 1652 324 1653
rect 414 1657 420 1658
rect 414 1653 415 1657
rect 419 1653 420 1657
rect 414 1652 420 1653
rect 510 1657 516 1658
rect 510 1653 511 1657
rect 515 1653 516 1657
rect 510 1652 516 1653
rect 614 1657 620 1658
rect 614 1653 615 1657
rect 619 1653 620 1657
rect 614 1652 620 1653
rect 710 1657 716 1658
rect 710 1653 711 1657
rect 715 1653 716 1657
rect 710 1652 716 1653
rect 798 1657 804 1658
rect 798 1653 799 1657
rect 803 1653 804 1657
rect 798 1652 804 1653
rect 878 1657 884 1658
rect 878 1653 879 1657
rect 883 1653 884 1657
rect 878 1652 884 1653
rect 950 1657 956 1658
rect 950 1653 951 1657
rect 955 1653 956 1657
rect 950 1652 956 1653
rect 1014 1657 1020 1658
rect 1014 1653 1015 1657
rect 1019 1653 1020 1657
rect 1014 1652 1020 1653
rect 1086 1657 1092 1658
rect 1086 1653 1087 1657
rect 1091 1653 1092 1657
rect 1086 1652 1092 1653
rect 1158 1657 1164 1658
rect 1158 1653 1159 1657
rect 1163 1653 1164 1657
rect 1158 1652 1164 1653
rect 136 1639 138 1652
rect 176 1639 178 1652
rect 240 1639 242 1652
rect 320 1639 322 1652
rect 416 1639 418 1652
rect 512 1639 514 1652
rect 616 1639 618 1652
rect 712 1639 714 1652
rect 800 1639 802 1652
rect 880 1639 882 1652
rect 952 1639 954 1652
rect 1016 1639 1018 1652
rect 1088 1639 1090 1652
rect 1160 1639 1162 1652
rect 1240 1639 1242 1675
rect 1280 1671 1282 1678
rect 1302 1676 1308 1677
rect 1302 1672 1303 1676
rect 1307 1672 1308 1676
rect 1302 1671 1308 1672
rect 1350 1676 1356 1677
rect 1350 1672 1351 1676
rect 1355 1672 1356 1676
rect 1350 1671 1356 1672
rect 1422 1676 1428 1677
rect 1422 1672 1423 1676
rect 1427 1672 1428 1676
rect 1422 1671 1428 1672
rect 1502 1676 1508 1677
rect 1502 1672 1503 1676
rect 1507 1672 1508 1676
rect 1502 1671 1508 1672
rect 1582 1676 1588 1677
rect 1582 1672 1583 1676
rect 1587 1672 1588 1676
rect 1582 1671 1588 1672
rect 1662 1676 1668 1677
rect 1662 1672 1663 1676
rect 1667 1672 1668 1676
rect 1662 1671 1668 1672
rect 1734 1676 1740 1677
rect 1734 1672 1735 1676
rect 1739 1672 1740 1676
rect 1734 1671 1740 1672
rect 1806 1676 1812 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1870 1676 1876 1677
rect 1870 1672 1871 1676
rect 1875 1672 1876 1676
rect 1870 1671 1876 1672
rect 1934 1676 1940 1677
rect 1934 1672 1935 1676
rect 1939 1672 1940 1676
rect 1934 1671 1940 1672
rect 1998 1676 2004 1677
rect 1998 1672 1999 1676
rect 2003 1672 2004 1676
rect 1998 1671 2004 1672
rect 2062 1676 2068 1677
rect 2062 1672 2063 1676
rect 2067 1672 2068 1676
rect 2062 1671 2068 1672
rect 2408 1671 2410 1678
rect 1279 1670 1283 1671
rect 1279 1665 1283 1666
rect 1303 1670 1307 1671
rect 1303 1665 1307 1666
rect 1351 1670 1355 1671
rect 1351 1665 1355 1666
rect 1359 1670 1363 1671
rect 1359 1665 1363 1666
rect 1423 1670 1427 1671
rect 1423 1665 1427 1666
rect 1447 1670 1451 1671
rect 1447 1665 1451 1666
rect 1503 1670 1507 1671
rect 1503 1665 1507 1666
rect 1543 1670 1547 1671
rect 1543 1665 1547 1666
rect 1583 1670 1587 1671
rect 1583 1665 1587 1666
rect 1639 1670 1643 1671
rect 1639 1665 1643 1666
rect 1663 1670 1667 1671
rect 1663 1665 1667 1666
rect 1727 1670 1731 1671
rect 1727 1665 1731 1666
rect 1735 1670 1739 1671
rect 1735 1665 1739 1666
rect 1807 1670 1811 1671
rect 1807 1665 1811 1666
rect 1815 1670 1819 1671
rect 1815 1665 1819 1666
rect 1871 1670 1875 1671
rect 1871 1665 1875 1666
rect 1895 1670 1899 1671
rect 1895 1665 1899 1666
rect 1935 1670 1939 1671
rect 1935 1665 1939 1666
rect 1967 1670 1971 1671
rect 1967 1665 1971 1666
rect 1999 1670 2003 1671
rect 1999 1665 2003 1666
rect 2031 1670 2035 1671
rect 2031 1665 2035 1666
rect 2063 1670 2067 1671
rect 2063 1665 2067 1666
rect 2095 1670 2099 1671
rect 2095 1665 2099 1666
rect 2159 1670 2163 1671
rect 2159 1665 2163 1666
rect 2223 1670 2227 1671
rect 2223 1665 2227 1666
rect 2407 1670 2411 1671
rect 2407 1665 2411 1666
rect 1280 1658 1282 1665
rect 1302 1664 1308 1665
rect 1302 1660 1303 1664
rect 1307 1660 1308 1664
rect 1302 1659 1308 1660
rect 1358 1664 1364 1665
rect 1358 1660 1359 1664
rect 1363 1660 1364 1664
rect 1358 1659 1364 1660
rect 1446 1664 1452 1665
rect 1446 1660 1447 1664
rect 1451 1660 1452 1664
rect 1446 1659 1452 1660
rect 1542 1664 1548 1665
rect 1542 1660 1543 1664
rect 1547 1660 1548 1664
rect 1542 1659 1548 1660
rect 1638 1664 1644 1665
rect 1638 1660 1639 1664
rect 1643 1660 1644 1664
rect 1638 1659 1644 1660
rect 1726 1664 1732 1665
rect 1726 1660 1727 1664
rect 1731 1660 1732 1664
rect 1726 1659 1732 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1894 1664 1900 1665
rect 1894 1660 1895 1664
rect 1899 1660 1900 1664
rect 1894 1659 1900 1660
rect 1966 1664 1972 1665
rect 1966 1660 1967 1664
rect 1971 1660 1972 1664
rect 1966 1659 1972 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2094 1664 2100 1665
rect 2094 1660 2095 1664
rect 2099 1660 2100 1664
rect 2094 1659 2100 1660
rect 2158 1664 2164 1665
rect 2158 1660 2159 1664
rect 2163 1660 2164 1664
rect 2158 1659 2164 1660
rect 2222 1664 2228 1665
rect 2222 1660 2223 1664
rect 2227 1660 2228 1664
rect 2222 1659 2228 1660
rect 2408 1658 2410 1665
rect 1278 1657 1284 1658
rect 1278 1653 1279 1657
rect 1283 1653 1284 1657
rect 1278 1652 1284 1653
rect 2406 1657 2412 1658
rect 2406 1653 2407 1657
rect 2411 1653 2412 1657
rect 2406 1652 2412 1653
rect 1278 1640 1284 1641
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 175 1638 179 1639
rect 175 1633 179 1634
rect 239 1638 243 1639
rect 239 1633 243 1634
rect 271 1638 275 1639
rect 271 1633 275 1634
rect 311 1638 315 1639
rect 311 1633 315 1634
rect 319 1638 323 1639
rect 319 1633 323 1634
rect 359 1638 363 1639
rect 359 1633 363 1634
rect 415 1638 419 1639
rect 415 1633 419 1634
rect 471 1638 475 1639
rect 471 1633 475 1634
rect 511 1638 515 1639
rect 511 1633 515 1634
rect 535 1638 539 1639
rect 535 1633 539 1634
rect 599 1638 603 1639
rect 599 1633 603 1634
rect 615 1638 619 1639
rect 615 1633 619 1634
rect 663 1638 667 1639
rect 663 1633 667 1634
rect 711 1638 715 1639
rect 711 1633 715 1634
rect 719 1638 723 1639
rect 719 1633 723 1634
rect 775 1638 779 1639
rect 775 1633 779 1634
rect 799 1638 803 1639
rect 799 1633 803 1634
rect 831 1638 835 1639
rect 831 1633 835 1634
rect 879 1638 883 1639
rect 879 1633 883 1634
rect 887 1638 891 1639
rect 887 1633 891 1634
rect 943 1638 947 1639
rect 943 1633 947 1634
rect 951 1638 955 1639
rect 951 1633 955 1634
rect 999 1638 1003 1639
rect 999 1633 1003 1634
rect 1015 1638 1019 1639
rect 1015 1633 1019 1634
rect 1087 1638 1091 1639
rect 1087 1633 1091 1634
rect 1159 1638 1163 1639
rect 1159 1633 1163 1634
rect 1239 1638 1243 1639
rect 1278 1636 1279 1640
rect 1283 1636 1284 1640
rect 1278 1635 1284 1636
rect 2406 1640 2412 1641
rect 2406 1636 2407 1640
rect 2411 1636 2412 1640
rect 2406 1635 2412 1636
rect 1239 1633 1243 1634
rect 112 1601 114 1633
rect 272 1624 274 1633
rect 312 1624 314 1633
rect 360 1624 362 1633
rect 416 1624 418 1633
rect 472 1624 474 1633
rect 536 1624 538 1633
rect 600 1624 602 1633
rect 664 1624 666 1633
rect 720 1624 722 1633
rect 776 1624 778 1633
rect 832 1624 834 1633
rect 888 1624 890 1633
rect 944 1624 946 1633
rect 1000 1624 1002 1633
rect 270 1623 276 1624
rect 270 1619 271 1623
rect 275 1619 276 1623
rect 270 1618 276 1619
rect 310 1623 316 1624
rect 310 1619 311 1623
rect 315 1619 316 1623
rect 310 1618 316 1619
rect 358 1623 364 1624
rect 358 1619 359 1623
rect 363 1619 364 1623
rect 358 1618 364 1619
rect 414 1623 420 1624
rect 414 1619 415 1623
rect 419 1619 420 1623
rect 414 1618 420 1619
rect 470 1623 476 1624
rect 470 1619 471 1623
rect 475 1619 476 1623
rect 470 1618 476 1619
rect 534 1623 540 1624
rect 534 1619 535 1623
rect 539 1619 540 1623
rect 534 1618 540 1619
rect 598 1623 604 1624
rect 598 1619 599 1623
rect 603 1619 604 1623
rect 598 1618 604 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 718 1623 724 1624
rect 718 1619 719 1623
rect 723 1619 724 1623
rect 718 1618 724 1619
rect 774 1623 780 1624
rect 774 1619 775 1623
rect 779 1619 780 1623
rect 774 1618 780 1619
rect 830 1623 836 1624
rect 830 1619 831 1623
rect 835 1619 836 1623
rect 830 1618 836 1619
rect 886 1623 892 1624
rect 886 1619 887 1623
rect 891 1619 892 1623
rect 886 1618 892 1619
rect 942 1623 948 1624
rect 942 1619 943 1623
rect 947 1619 948 1623
rect 942 1618 948 1619
rect 998 1623 1004 1624
rect 998 1619 999 1623
rect 1003 1619 1004 1623
rect 998 1618 1004 1619
rect 1240 1601 1242 1633
rect 1280 1603 1282 1635
rect 1302 1617 1308 1618
rect 1302 1613 1303 1617
rect 1307 1613 1308 1617
rect 1302 1612 1308 1613
rect 1358 1617 1364 1618
rect 1358 1613 1359 1617
rect 1363 1613 1364 1617
rect 1358 1612 1364 1613
rect 1446 1617 1452 1618
rect 1446 1613 1447 1617
rect 1451 1613 1452 1617
rect 1446 1612 1452 1613
rect 1542 1617 1548 1618
rect 1542 1613 1543 1617
rect 1547 1613 1548 1617
rect 1542 1612 1548 1613
rect 1638 1617 1644 1618
rect 1638 1613 1639 1617
rect 1643 1613 1644 1617
rect 1638 1612 1644 1613
rect 1726 1617 1732 1618
rect 1726 1613 1727 1617
rect 1731 1613 1732 1617
rect 1726 1612 1732 1613
rect 1814 1617 1820 1618
rect 1814 1613 1815 1617
rect 1819 1613 1820 1617
rect 1814 1612 1820 1613
rect 1894 1617 1900 1618
rect 1894 1613 1895 1617
rect 1899 1613 1900 1617
rect 1894 1612 1900 1613
rect 1966 1617 1972 1618
rect 1966 1613 1967 1617
rect 1971 1613 1972 1617
rect 1966 1612 1972 1613
rect 2030 1617 2036 1618
rect 2030 1613 2031 1617
rect 2035 1613 2036 1617
rect 2030 1612 2036 1613
rect 2094 1617 2100 1618
rect 2094 1613 2095 1617
rect 2099 1613 2100 1617
rect 2094 1612 2100 1613
rect 2158 1617 2164 1618
rect 2158 1613 2159 1617
rect 2163 1613 2164 1617
rect 2158 1612 2164 1613
rect 2222 1617 2228 1618
rect 2222 1613 2223 1617
rect 2227 1613 2228 1617
rect 2222 1612 2228 1613
rect 1304 1603 1306 1612
rect 1360 1603 1362 1612
rect 1448 1603 1450 1612
rect 1544 1603 1546 1612
rect 1640 1603 1642 1612
rect 1728 1603 1730 1612
rect 1816 1603 1818 1612
rect 1896 1603 1898 1612
rect 1968 1603 1970 1612
rect 2032 1603 2034 1612
rect 2096 1603 2098 1612
rect 2160 1603 2162 1612
rect 2224 1603 2226 1612
rect 2408 1603 2410 1635
rect 1279 1602 1283 1603
rect 110 1600 116 1601
rect 110 1596 111 1600
rect 115 1596 116 1600
rect 110 1595 116 1596
rect 1238 1600 1244 1601
rect 1238 1596 1239 1600
rect 1243 1596 1244 1600
rect 1279 1597 1283 1598
rect 1303 1602 1307 1603
rect 1303 1597 1307 1598
rect 1327 1602 1331 1603
rect 1327 1597 1331 1598
rect 1359 1602 1363 1603
rect 1359 1597 1363 1598
rect 1399 1602 1403 1603
rect 1399 1597 1403 1598
rect 1447 1602 1451 1603
rect 1447 1597 1451 1598
rect 1479 1602 1483 1603
rect 1479 1597 1483 1598
rect 1543 1602 1547 1603
rect 1543 1597 1547 1598
rect 1567 1602 1571 1603
rect 1567 1597 1571 1598
rect 1639 1602 1643 1603
rect 1639 1597 1643 1598
rect 1655 1602 1659 1603
rect 1655 1597 1659 1598
rect 1727 1602 1731 1603
rect 1727 1597 1731 1598
rect 1743 1602 1747 1603
rect 1743 1597 1747 1598
rect 1815 1602 1819 1603
rect 1815 1597 1819 1598
rect 1831 1602 1835 1603
rect 1831 1597 1835 1598
rect 1895 1602 1899 1603
rect 1895 1597 1899 1598
rect 1911 1602 1915 1603
rect 1911 1597 1915 1598
rect 1967 1602 1971 1603
rect 1967 1597 1971 1598
rect 1983 1602 1987 1603
rect 1983 1597 1987 1598
rect 2031 1602 2035 1603
rect 2031 1597 2035 1598
rect 2047 1602 2051 1603
rect 2047 1597 2051 1598
rect 2095 1602 2099 1603
rect 2095 1597 2099 1598
rect 2111 1602 2115 1603
rect 2111 1597 2115 1598
rect 2159 1602 2163 1603
rect 2159 1597 2163 1598
rect 2167 1602 2171 1603
rect 2167 1597 2171 1598
rect 2215 1602 2219 1603
rect 2215 1597 2219 1598
rect 2223 1602 2227 1603
rect 2223 1597 2227 1598
rect 2271 1602 2275 1603
rect 2271 1597 2275 1598
rect 2319 1602 2323 1603
rect 2319 1597 2323 1598
rect 2359 1602 2363 1603
rect 2359 1597 2363 1598
rect 2407 1602 2411 1603
rect 2407 1597 2411 1598
rect 1238 1595 1244 1596
rect 110 1583 116 1584
rect 110 1579 111 1583
rect 115 1579 116 1583
rect 110 1578 116 1579
rect 1238 1583 1244 1584
rect 1238 1579 1239 1583
rect 1243 1579 1244 1583
rect 1238 1578 1244 1579
rect 112 1563 114 1578
rect 270 1576 276 1577
rect 270 1572 271 1576
rect 275 1572 276 1576
rect 270 1571 276 1572
rect 310 1576 316 1577
rect 310 1572 311 1576
rect 315 1572 316 1576
rect 310 1571 316 1572
rect 358 1576 364 1577
rect 358 1572 359 1576
rect 363 1572 364 1576
rect 358 1571 364 1572
rect 414 1576 420 1577
rect 414 1572 415 1576
rect 419 1572 420 1576
rect 414 1571 420 1572
rect 470 1576 476 1577
rect 470 1572 471 1576
rect 475 1572 476 1576
rect 470 1571 476 1572
rect 534 1576 540 1577
rect 534 1572 535 1576
rect 539 1572 540 1576
rect 534 1571 540 1572
rect 598 1576 604 1577
rect 598 1572 599 1576
rect 603 1572 604 1576
rect 598 1571 604 1572
rect 662 1576 668 1577
rect 662 1572 663 1576
rect 667 1572 668 1576
rect 662 1571 668 1572
rect 718 1576 724 1577
rect 718 1572 719 1576
rect 723 1572 724 1576
rect 718 1571 724 1572
rect 774 1576 780 1577
rect 774 1572 775 1576
rect 779 1572 780 1576
rect 774 1571 780 1572
rect 830 1576 836 1577
rect 830 1572 831 1576
rect 835 1572 836 1576
rect 830 1571 836 1572
rect 886 1576 892 1577
rect 886 1572 887 1576
rect 891 1572 892 1576
rect 886 1571 892 1572
rect 942 1576 948 1577
rect 942 1572 943 1576
rect 947 1572 948 1576
rect 942 1571 948 1572
rect 998 1576 1004 1577
rect 998 1572 999 1576
rect 1003 1572 1004 1576
rect 998 1571 1004 1572
rect 272 1563 274 1571
rect 312 1563 314 1571
rect 360 1563 362 1571
rect 416 1563 418 1571
rect 472 1563 474 1571
rect 536 1563 538 1571
rect 600 1563 602 1571
rect 664 1563 666 1571
rect 720 1563 722 1571
rect 776 1563 778 1571
rect 832 1563 834 1571
rect 888 1563 890 1571
rect 944 1563 946 1571
rect 1000 1563 1002 1571
rect 1240 1563 1242 1578
rect 1280 1565 1282 1597
rect 1328 1588 1330 1597
rect 1400 1588 1402 1597
rect 1480 1588 1482 1597
rect 1568 1588 1570 1597
rect 1656 1588 1658 1597
rect 1744 1588 1746 1597
rect 1832 1588 1834 1597
rect 1912 1588 1914 1597
rect 1984 1588 1986 1597
rect 2048 1588 2050 1597
rect 2112 1588 2114 1597
rect 2168 1588 2170 1597
rect 2216 1588 2218 1597
rect 2272 1588 2274 1597
rect 2320 1588 2322 1597
rect 2360 1588 2362 1597
rect 1326 1587 1332 1588
rect 1326 1583 1327 1587
rect 1331 1583 1332 1587
rect 1326 1582 1332 1583
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1583 1404 1587
rect 1398 1582 1404 1583
rect 1478 1587 1484 1588
rect 1478 1583 1479 1587
rect 1483 1583 1484 1587
rect 1478 1582 1484 1583
rect 1566 1587 1572 1588
rect 1566 1583 1567 1587
rect 1571 1583 1572 1587
rect 1566 1582 1572 1583
rect 1654 1587 1660 1588
rect 1654 1583 1655 1587
rect 1659 1583 1660 1587
rect 1654 1582 1660 1583
rect 1742 1587 1748 1588
rect 1742 1583 1743 1587
rect 1747 1583 1748 1587
rect 1742 1582 1748 1583
rect 1830 1587 1836 1588
rect 1830 1583 1831 1587
rect 1835 1583 1836 1587
rect 1830 1582 1836 1583
rect 1910 1587 1916 1588
rect 1910 1583 1911 1587
rect 1915 1583 1916 1587
rect 1910 1582 1916 1583
rect 1982 1587 1988 1588
rect 1982 1583 1983 1587
rect 1987 1583 1988 1587
rect 1982 1582 1988 1583
rect 2046 1587 2052 1588
rect 2046 1583 2047 1587
rect 2051 1583 2052 1587
rect 2046 1582 2052 1583
rect 2110 1587 2116 1588
rect 2110 1583 2111 1587
rect 2115 1583 2116 1587
rect 2110 1582 2116 1583
rect 2166 1587 2172 1588
rect 2166 1583 2167 1587
rect 2171 1583 2172 1587
rect 2166 1582 2172 1583
rect 2214 1587 2220 1588
rect 2214 1583 2215 1587
rect 2219 1583 2220 1587
rect 2214 1582 2220 1583
rect 2270 1587 2276 1588
rect 2270 1583 2271 1587
rect 2275 1583 2276 1587
rect 2270 1582 2276 1583
rect 2318 1587 2324 1588
rect 2318 1583 2319 1587
rect 2323 1583 2324 1587
rect 2318 1582 2324 1583
rect 2358 1587 2364 1588
rect 2358 1583 2359 1587
rect 2363 1583 2364 1587
rect 2358 1582 2364 1583
rect 2408 1565 2410 1597
rect 1278 1564 1284 1565
rect 111 1562 115 1563
rect 111 1557 115 1558
rect 271 1562 275 1563
rect 271 1557 275 1558
rect 311 1562 315 1563
rect 311 1557 315 1558
rect 327 1562 331 1563
rect 327 1557 331 1558
rect 359 1562 363 1563
rect 359 1557 363 1558
rect 367 1562 371 1563
rect 367 1557 371 1558
rect 407 1562 411 1563
rect 407 1557 411 1558
rect 415 1562 419 1563
rect 415 1557 419 1558
rect 447 1562 451 1563
rect 447 1557 451 1558
rect 471 1562 475 1563
rect 471 1557 475 1558
rect 487 1562 491 1563
rect 487 1557 491 1558
rect 527 1562 531 1563
rect 527 1557 531 1558
rect 535 1562 539 1563
rect 535 1557 539 1558
rect 567 1562 571 1563
rect 567 1557 571 1558
rect 599 1562 603 1563
rect 599 1557 603 1558
rect 607 1562 611 1563
rect 607 1557 611 1558
rect 647 1562 651 1563
rect 647 1557 651 1558
rect 663 1562 667 1563
rect 663 1557 667 1558
rect 687 1562 691 1563
rect 687 1557 691 1558
rect 719 1562 723 1563
rect 719 1557 723 1558
rect 727 1562 731 1563
rect 727 1557 731 1558
rect 767 1562 771 1563
rect 767 1557 771 1558
rect 775 1562 779 1563
rect 775 1557 779 1558
rect 807 1562 811 1563
rect 807 1557 811 1558
rect 831 1562 835 1563
rect 831 1557 835 1558
rect 847 1562 851 1563
rect 847 1557 851 1558
rect 887 1562 891 1563
rect 887 1557 891 1558
rect 927 1562 931 1563
rect 927 1557 931 1558
rect 943 1562 947 1563
rect 943 1557 947 1558
rect 999 1562 1003 1563
rect 999 1557 1003 1558
rect 1239 1562 1243 1563
rect 1278 1560 1279 1564
rect 1283 1560 1284 1564
rect 1278 1559 1284 1560
rect 2406 1564 2412 1565
rect 2406 1560 2407 1564
rect 2411 1560 2412 1564
rect 2406 1559 2412 1560
rect 1239 1557 1243 1558
rect 112 1550 114 1557
rect 326 1556 332 1557
rect 326 1552 327 1556
rect 331 1552 332 1556
rect 326 1551 332 1552
rect 366 1556 372 1557
rect 366 1552 367 1556
rect 371 1552 372 1556
rect 366 1551 372 1552
rect 406 1556 412 1557
rect 406 1552 407 1556
rect 411 1552 412 1556
rect 406 1551 412 1552
rect 446 1556 452 1557
rect 446 1552 447 1556
rect 451 1552 452 1556
rect 446 1551 452 1552
rect 486 1556 492 1557
rect 486 1552 487 1556
rect 491 1552 492 1556
rect 486 1551 492 1552
rect 526 1556 532 1557
rect 526 1552 527 1556
rect 531 1552 532 1556
rect 526 1551 532 1552
rect 566 1556 572 1557
rect 566 1552 567 1556
rect 571 1552 572 1556
rect 566 1551 572 1552
rect 606 1556 612 1557
rect 606 1552 607 1556
rect 611 1552 612 1556
rect 606 1551 612 1552
rect 646 1556 652 1557
rect 646 1552 647 1556
rect 651 1552 652 1556
rect 646 1551 652 1552
rect 686 1556 692 1557
rect 686 1552 687 1556
rect 691 1552 692 1556
rect 686 1551 692 1552
rect 726 1556 732 1557
rect 726 1552 727 1556
rect 731 1552 732 1556
rect 726 1551 732 1552
rect 766 1556 772 1557
rect 766 1552 767 1556
rect 771 1552 772 1556
rect 766 1551 772 1552
rect 806 1556 812 1557
rect 806 1552 807 1556
rect 811 1552 812 1556
rect 806 1551 812 1552
rect 846 1556 852 1557
rect 846 1552 847 1556
rect 851 1552 852 1556
rect 846 1551 852 1552
rect 886 1556 892 1557
rect 886 1552 887 1556
rect 891 1552 892 1556
rect 886 1551 892 1552
rect 926 1556 932 1557
rect 926 1552 927 1556
rect 931 1552 932 1556
rect 926 1551 932 1552
rect 1240 1550 1242 1557
rect 110 1549 116 1550
rect 110 1545 111 1549
rect 115 1545 116 1549
rect 110 1544 116 1545
rect 1238 1549 1244 1550
rect 1238 1545 1239 1549
rect 1243 1545 1244 1549
rect 1238 1544 1244 1545
rect 1278 1547 1284 1548
rect 1278 1543 1279 1547
rect 1283 1543 1284 1547
rect 1278 1542 1284 1543
rect 2406 1547 2412 1548
rect 2406 1543 2407 1547
rect 2411 1543 2412 1547
rect 2406 1542 2412 1543
rect 110 1532 116 1533
rect 110 1528 111 1532
rect 115 1528 116 1532
rect 110 1527 116 1528
rect 1238 1532 1244 1533
rect 1238 1528 1239 1532
rect 1243 1528 1244 1532
rect 1280 1531 1282 1542
rect 1326 1540 1332 1541
rect 1326 1536 1327 1540
rect 1331 1536 1332 1540
rect 1326 1535 1332 1536
rect 1398 1540 1404 1541
rect 1398 1536 1399 1540
rect 1403 1536 1404 1540
rect 1398 1535 1404 1536
rect 1478 1540 1484 1541
rect 1478 1536 1479 1540
rect 1483 1536 1484 1540
rect 1478 1535 1484 1536
rect 1566 1540 1572 1541
rect 1566 1536 1567 1540
rect 1571 1536 1572 1540
rect 1566 1535 1572 1536
rect 1654 1540 1660 1541
rect 1654 1536 1655 1540
rect 1659 1536 1660 1540
rect 1654 1535 1660 1536
rect 1742 1540 1748 1541
rect 1742 1536 1743 1540
rect 1747 1536 1748 1540
rect 1742 1535 1748 1536
rect 1830 1540 1836 1541
rect 1830 1536 1831 1540
rect 1835 1536 1836 1540
rect 1830 1535 1836 1536
rect 1910 1540 1916 1541
rect 1910 1536 1911 1540
rect 1915 1536 1916 1540
rect 1910 1535 1916 1536
rect 1982 1540 1988 1541
rect 1982 1536 1983 1540
rect 1987 1536 1988 1540
rect 1982 1535 1988 1536
rect 2046 1540 2052 1541
rect 2046 1536 2047 1540
rect 2051 1536 2052 1540
rect 2046 1535 2052 1536
rect 2110 1540 2116 1541
rect 2110 1536 2111 1540
rect 2115 1536 2116 1540
rect 2110 1535 2116 1536
rect 2166 1540 2172 1541
rect 2166 1536 2167 1540
rect 2171 1536 2172 1540
rect 2166 1535 2172 1536
rect 2214 1540 2220 1541
rect 2214 1536 2215 1540
rect 2219 1536 2220 1540
rect 2214 1535 2220 1536
rect 2270 1540 2276 1541
rect 2270 1536 2271 1540
rect 2275 1536 2276 1540
rect 2270 1535 2276 1536
rect 2318 1540 2324 1541
rect 2318 1536 2319 1540
rect 2323 1536 2324 1540
rect 2318 1535 2324 1536
rect 2358 1540 2364 1541
rect 2358 1536 2359 1540
rect 2363 1536 2364 1540
rect 2358 1535 2364 1536
rect 1328 1531 1330 1535
rect 1400 1531 1402 1535
rect 1480 1531 1482 1535
rect 1568 1531 1570 1535
rect 1656 1531 1658 1535
rect 1744 1531 1746 1535
rect 1832 1531 1834 1535
rect 1912 1531 1914 1535
rect 1984 1531 1986 1535
rect 2048 1531 2050 1535
rect 2112 1531 2114 1535
rect 2168 1531 2170 1535
rect 2216 1531 2218 1535
rect 2272 1531 2274 1535
rect 2320 1531 2322 1535
rect 2360 1531 2362 1535
rect 2408 1531 2410 1542
rect 1238 1527 1244 1528
rect 1279 1530 1283 1531
rect 112 1455 114 1527
rect 326 1509 332 1510
rect 326 1505 327 1509
rect 331 1505 332 1509
rect 326 1504 332 1505
rect 366 1509 372 1510
rect 366 1505 367 1509
rect 371 1505 372 1509
rect 366 1504 372 1505
rect 406 1509 412 1510
rect 406 1505 407 1509
rect 411 1505 412 1509
rect 406 1504 412 1505
rect 446 1509 452 1510
rect 446 1505 447 1509
rect 451 1505 452 1509
rect 446 1504 452 1505
rect 486 1509 492 1510
rect 486 1505 487 1509
rect 491 1505 492 1509
rect 486 1504 492 1505
rect 526 1509 532 1510
rect 526 1505 527 1509
rect 531 1505 532 1509
rect 526 1504 532 1505
rect 566 1509 572 1510
rect 566 1505 567 1509
rect 571 1505 572 1509
rect 566 1504 572 1505
rect 606 1509 612 1510
rect 606 1505 607 1509
rect 611 1505 612 1509
rect 606 1504 612 1505
rect 646 1509 652 1510
rect 646 1505 647 1509
rect 651 1505 652 1509
rect 646 1504 652 1505
rect 686 1509 692 1510
rect 686 1505 687 1509
rect 691 1505 692 1509
rect 686 1504 692 1505
rect 726 1509 732 1510
rect 726 1505 727 1509
rect 731 1505 732 1509
rect 726 1504 732 1505
rect 766 1509 772 1510
rect 766 1505 767 1509
rect 771 1505 772 1509
rect 766 1504 772 1505
rect 806 1509 812 1510
rect 806 1505 807 1509
rect 811 1505 812 1509
rect 806 1504 812 1505
rect 846 1509 852 1510
rect 846 1505 847 1509
rect 851 1505 852 1509
rect 846 1504 852 1505
rect 886 1509 892 1510
rect 886 1505 887 1509
rect 891 1505 892 1509
rect 886 1504 892 1505
rect 926 1509 932 1510
rect 926 1505 927 1509
rect 931 1505 932 1509
rect 926 1504 932 1505
rect 328 1455 330 1504
rect 368 1455 370 1504
rect 408 1455 410 1504
rect 448 1455 450 1504
rect 488 1455 490 1504
rect 528 1455 530 1504
rect 568 1455 570 1504
rect 608 1455 610 1504
rect 648 1455 650 1504
rect 688 1455 690 1504
rect 728 1455 730 1504
rect 768 1455 770 1504
rect 808 1455 810 1504
rect 848 1455 850 1504
rect 888 1455 890 1504
rect 928 1455 930 1504
rect 1240 1455 1242 1527
rect 1279 1525 1283 1526
rect 1327 1530 1331 1531
rect 1327 1525 1331 1526
rect 1335 1530 1339 1531
rect 1335 1525 1339 1526
rect 1399 1530 1403 1531
rect 1399 1525 1403 1526
rect 1415 1530 1419 1531
rect 1415 1525 1419 1526
rect 1479 1530 1483 1531
rect 1479 1525 1483 1526
rect 1503 1530 1507 1531
rect 1503 1525 1507 1526
rect 1567 1530 1571 1531
rect 1567 1525 1571 1526
rect 1615 1530 1619 1531
rect 1615 1525 1619 1526
rect 1655 1530 1659 1531
rect 1655 1525 1659 1526
rect 1743 1530 1747 1531
rect 1743 1525 1747 1526
rect 1831 1530 1835 1531
rect 1831 1525 1835 1526
rect 1887 1530 1891 1531
rect 1887 1525 1891 1526
rect 1911 1530 1915 1531
rect 1911 1525 1915 1526
rect 1983 1530 1987 1531
rect 1983 1525 1987 1526
rect 2047 1530 2051 1531
rect 2047 1525 2051 1526
rect 2111 1530 2115 1531
rect 2111 1525 2115 1526
rect 2167 1530 2171 1531
rect 2167 1525 2171 1526
rect 2215 1530 2219 1531
rect 2215 1525 2219 1526
rect 2271 1530 2275 1531
rect 2271 1525 2275 1526
rect 2319 1530 2323 1531
rect 2319 1525 2323 1526
rect 2359 1530 2363 1531
rect 2359 1525 2363 1526
rect 2407 1530 2411 1531
rect 2407 1525 2411 1526
rect 1280 1518 1282 1525
rect 1334 1524 1340 1525
rect 1334 1520 1335 1524
rect 1339 1520 1340 1524
rect 1334 1519 1340 1520
rect 1414 1524 1420 1525
rect 1414 1520 1415 1524
rect 1419 1520 1420 1524
rect 1414 1519 1420 1520
rect 1502 1524 1508 1525
rect 1502 1520 1503 1524
rect 1507 1520 1508 1524
rect 1502 1519 1508 1520
rect 1614 1524 1620 1525
rect 1614 1520 1615 1524
rect 1619 1520 1620 1524
rect 1614 1519 1620 1520
rect 1742 1524 1748 1525
rect 1742 1520 1743 1524
rect 1747 1520 1748 1524
rect 1742 1519 1748 1520
rect 1886 1524 1892 1525
rect 1886 1520 1887 1524
rect 1891 1520 1892 1524
rect 1886 1519 1892 1520
rect 2046 1524 2052 1525
rect 2046 1520 2047 1524
rect 2051 1520 2052 1524
rect 2046 1519 2052 1520
rect 2214 1524 2220 1525
rect 2214 1520 2215 1524
rect 2219 1520 2220 1524
rect 2214 1519 2220 1520
rect 2358 1524 2364 1525
rect 2358 1520 2359 1524
rect 2363 1520 2364 1524
rect 2358 1519 2364 1520
rect 2408 1518 2410 1525
rect 1278 1517 1284 1518
rect 1278 1513 1279 1517
rect 1283 1513 1284 1517
rect 1278 1512 1284 1513
rect 2406 1517 2412 1518
rect 2406 1513 2407 1517
rect 2411 1513 2412 1517
rect 2406 1512 2412 1513
rect 1278 1500 1284 1501
rect 1278 1496 1279 1500
rect 1283 1496 1284 1500
rect 1278 1495 1284 1496
rect 2406 1500 2412 1501
rect 2406 1496 2407 1500
rect 2411 1496 2412 1500
rect 2406 1495 2412 1496
rect 1280 1463 1282 1495
rect 1334 1477 1340 1478
rect 1334 1473 1335 1477
rect 1339 1473 1340 1477
rect 1334 1472 1340 1473
rect 1414 1477 1420 1478
rect 1414 1473 1415 1477
rect 1419 1473 1420 1477
rect 1414 1472 1420 1473
rect 1502 1477 1508 1478
rect 1502 1473 1503 1477
rect 1507 1473 1508 1477
rect 1502 1472 1508 1473
rect 1614 1477 1620 1478
rect 1614 1473 1615 1477
rect 1619 1473 1620 1477
rect 1614 1472 1620 1473
rect 1742 1477 1748 1478
rect 1742 1473 1743 1477
rect 1747 1473 1748 1477
rect 1742 1472 1748 1473
rect 1886 1477 1892 1478
rect 1886 1473 1887 1477
rect 1891 1473 1892 1477
rect 1886 1472 1892 1473
rect 2046 1477 2052 1478
rect 2046 1473 2047 1477
rect 2051 1473 2052 1477
rect 2046 1472 2052 1473
rect 2214 1477 2220 1478
rect 2214 1473 2215 1477
rect 2219 1473 2220 1477
rect 2214 1472 2220 1473
rect 2358 1477 2364 1478
rect 2358 1473 2359 1477
rect 2363 1473 2364 1477
rect 2358 1472 2364 1473
rect 1336 1463 1338 1472
rect 1416 1463 1418 1472
rect 1504 1463 1506 1472
rect 1616 1463 1618 1472
rect 1744 1463 1746 1472
rect 1888 1463 1890 1472
rect 2048 1463 2050 1472
rect 2216 1463 2218 1472
rect 2360 1463 2362 1472
rect 2408 1463 2410 1495
rect 1279 1462 1283 1463
rect 1279 1457 1283 1458
rect 1335 1462 1339 1463
rect 1335 1457 1339 1458
rect 1375 1462 1379 1463
rect 1375 1457 1379 1458
rect 1415 1462 1419 1463
rect 1415 1457 1419 1458
rect 1463 1462 1467 1463
rect 1463 1457 1467 1458
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1551 1462 1555 1463
rect 1551 1457 1555 1458
rect 1615 1462 1619 1463
rect 1615 1457 1619 1458
rect 1639 1462 1643 1463
rect 1639 1457 1643 1458
rect 1727 1462 1731 1463
rect 1727 1457 1731 1458
rect 1743 1462 1747 1463
rect 1743 1457 1747 1458
rect 1807 1462 1811 1463
rect 1807 1457 1811 1458
rect 1879 1462 1883 1463
rect 1879 1457 1883 1458
rect 1887 1462 1891 1463
rect 1887 1457 1891 1458
rect 1943 1462 1947 1463
rect 1943 1457 1947 1458
rect 1999 1462 2003 1463
rect 1999 1457 2003 1458
rect 2047 1462 2051 1463
rect 2047 1457 2051 1458
rect 2095 1462 2099 1463
rect 2095 1457 2099 1458
rect 2143 1462 2147 1463
rect 2143 1457 2147 1458
rect 2191 1462 2195 1463
rect 2191 1457 2195 1458
rect 2215 1462 2219 1463
rect 2215 1457 2219 1458
rect 2239 1462 2243 1463
rect 2239 1457 2243 1458
rect 2279 1462 2283 1463
rect 2279 1457 2283 1458
rect 2319 1462 2323 1463
rect 2319 1457 2323 1458
rect 2359 1462 2363 1463
rect 2359 1457 2363 1458
rect 2407 1462 2411 1463
rect 2407 1457 2411 1458
rect 111 1454 115 1455
rect 111 1449 115 1450
rect 143 1454 147 1455
rect 143 1449 147 1450
rect 183 1454 187 1455
rect 183 1449 187 1450
rect 223 1454 227 1455
rect 223 1449 227 1450
rect 263 1454 267 1455
rect 263 1449 267 1450
rect 319 1454 323 1455
rect 319 1449 323 1450
rect 327 1454 331 1455
rect 327 1449 331 1450
rect 367 1454 371 1455
rect 367 1449 371 1450
rect 391 1454 395 1455
rect 391 1449 395 1450
rect 407 1454 411 1455
rect 407 1449 411 1450
rect 447 1454 451 1455
rect 447 1449 451 1450
rect 471 1454 475 1455
rect 471 1449 475 1450
rect 487 1454 491 1455
rect 487 1449 491 1450
rect 527 1454 531 1455
rect 527 1449 531 1450
rect 559 1454 563 1455
rect 559 1449 563 1450
rect 567 1454 571 1455
rect 567 1449 571 1450
rect 607 1454 611 1455
rect 607 1449 611 1450
rect 647 1454 651 1455
rect 647 1449 651 1450
rect 687 1454 691 1455
rect 687 1449 691 1450
rect 727 1454 731 1455
rect 727 1449 731 1450
rect 767 1454 771 1455
rect 767 1449 771 1450
rect 807 1454 811 1455
rect 807 1449 811 1450
rect 847 1454 851 1455
rect 847 1449 851 1450
rect 879 1454 883 1455
rect 879 1449 883 1450
rect 887 1454 891 1455
rect 887 1449 891 1450
rect 927 1454 931 1455
rect 927 1449 931 1450
rect 943 1454 947 1455
rect 943 1449 947 1450
rect 999 1454 1003 1455
rect 999 1449 1003 1450
rect 1047 1454 1051 1455
rect 1047 1449 1051 1450
rect 1103 1454 1107 1455
rect 1103 1449 1107 1450
rect 1151 1454 1155 1455
rect 1151 1449 1155 1450
rect 1191 1454 1195 1455
rect 1191 1449 1195 1450
rect 1239 1454 1243 1455
rect 1239 1449 1243 1450
rect 112 1417 114 1449
rect 144 1440 146 1449
rect 184 1440 186 1449
rect 224 1440 226 1449
rect 264 1440 266 1449
rect 320 1440 322 1449
rect 392 1440 394 1449
rect 472 1440 474 1449
rect 560 1440 562 1449
rect 648 1440 650 1449
rect 728 1440 730 1449
rect 808 1440 810 1449
rect 880 1440 882 1449
rect 944 1440 946 1449
rect 1000 1440 1002 1449
rect 1048 1440 1050 1449
rect 1104 1440 1106 1449
rect 1152 1440 1154 1449
rect 1192 1440 1194 1449
rect 142 1439 148 1440
rect 142 1435 143 1439
rect 147 1435 148 1439
rect 142 1434 148 1435
rect 182 1439 188 1440
rect 182 1435 183 1439
rect 187 1435 188 1439
rect 182 1434 188 1435
rect 222 1439 228 1440
rect 222 1435 223 1439
rect 227 1435 228 1439
rect 222 1434 228 1435
rect 262 1439 268 1440
rect 262 1435 263 1439
rect 267 1435 268 1439
rect 262 1434 268 1435
rect 318 1439 324 1440
rect 318 1435 319 1439
rect 323 1435 324 1439
rect 318 1434 324 1435
rect 390 1439 396 1440
rect 390 1435 391 1439
rect 395 1435 396 1439
rect 390 1434 396 1435
rect 470 1439 476 1440
rect 470 1435 471 1439
rect 475 1435 476 1439
rect 470 1434 476 1435
rect 558 1439 564 1440
rect 558 1435 559 1439
rect 563 1435 564 1439
rect 558 1434 564 1435
rect 646 1439 652 1440
rect 646 1435 647 1439
rect 651 1435 652 1439
rect 646 1434 652 1435
rect 726 1439 732 1440
rect 726 1435 727 1439
rect 731 1435 732 1439
rect 726 1434 732 1435
rect 806 1439 812 1440
rect 806 1435 807 1439
rect 811 1435 812 1439
rect 806 1434 812 1435
rect 878 1439 884 1440
rect 878 1435 879 1439
rect 883 1435 884 1439
rect 878 1434 884 1435
rect 942 1439 948 1440
rect 942 1435 943 1439
rect 947 1435 948 1439
rect 942 1434 948 1435
rect 998 1439 1004 1440
rect 998 1435 999 1439
rect 1003 1435 1004 1439
rect 998 1434 1004 1435
rect 1046 1439 1052 1440
rect 1046 1435 1047 1439
rect 1051 1435 1052 1439
rect 1046 1434 1052 1435
rect 1102 1439 1108 1440
rect 1102 1435 1103 1439
rect 1107 1435 1108 1439
rect 1102 1434 1108 1435
rect 1150 1439 1156 1440
rect 1150 1435 1151 1439
rect 1155 1435 1156 1439
rect 1150 1434 1156 1435
rect 1190 1439 1196 1440
rect 1190 1435 1191 1439
rect 1195 1435 1196 1439
rect 1190 1434 1196 1435
rect 1240 1417 1242 1449
rect 1280 1425 1282 1457
rect 1376 1448 1378 1457
rect 1464 1448 1466 1457
rect 1552 1448 1554 1457
rect 1640 1448 1642 1457
rect 1728 1448 1730 1457
rect 1808 1448 1810 1457
rect 1880 1448 1882 1457
rect 1944 1448 1946 1457
rect 2000 1448 2002 1457
rect 2048 1448 2050 1457
rect 2096 1448 2098 1457
rect 2144 1448 2146 1457
rect 2192 1448 2194 1457
rect 2240 1448 2242 1457
rect 2280 1448 2282 1457
rect 2320 1448 2322 1457
rect 2360 1448 2362 1457
rect 1374 1447 1380 1448
rect 1374 1443 1375 1447
rect 1379 1443 1380 1447
rect 1374 1442 1380 1443
rect 1462 1447 1468 1448
rect 1462 1443 1463 1447
rect 1467 1443 1468 1447
rect 1462 1442 1468 1443
rect 1550 1447 1556 1448
rect 1550 1443 1551 1447
rect 1555 1443 1556 1447
rect 1550 1442 1556 1443
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1726 1447 1732 1448
rect 1726 1443 1727 1447
rect 1731 1443 1732 1447
rect 1726 1442 1732 1443
rect 1806 1447 1812 1448
rect 1806 1443 1807 1447
rect 1811 1443 1812 1447
rect 1806 1442 1812 1443
rect 1878 1447 1884 1448
rect 1878 1443 1879 1447
rect 1883 1443 1884 1447
rect 1878 1442 1884 1443
rect 1942 1447 1948 1448
rect 1942 1443 1943 1447
rect 1947 1443 1948 1447
rect 1942 1442 1948 1443
rect 1998 1447 2004 1448
rect 1998 1443 1999 1447
rect 2003 1443 2004 1447
rect 1998 1442 2004 1443
rect 2046 1447 2052 1448
rect 2046 1443 2047 1447
rect 2051 1443 2052 1447
rect 2046 1442 2052 1443
rect 2094 1447 2100 1448
rect 2094 1443 2095 1447
rect 2099 1443 2100 1447
rect 2094 1442 2100 1443
rect 2142 1447 2148 1448
rect 2142 1443 2143 1447
rect 2147 1443 2148 1447
rect 2142 1442 2148 1443
rect 2190 1447 2196 1448
rect 2190 1443 2191 1447
rect 2195 1443 2196 1447
rect 2190 1442 2196 1443
rect 2238 1447 2244 1448
rect 2238 1443 2239 1447
rect 2243 1443 2244 1447
rect 2238 1442 2244 1443
rect 2278 1447 2284 1448
rect 2278 1443 2279 1447
rect 2283 1443 2284 1447
rect 2278 1442 2284 1443
rect 2318 1447 2324 1448
rect 2318 1443 2319 1447
rect 2323 1443 2324 1447
rect 2318 1442 2324 1443
rect 2358 1447 2364 1448
rect 2358 1443 2359 1447
rect 2363 1443 2364 1447
rect 2358 1442 2364 1443
rect 2408 1425 2410 1457
rect 1278 1424 1284 1425
rect 1278 1420 1279 1424
rect 1283 1420 1284 1424
rect 1278 1419 1284 1420
rect 2406 1424 2412 1425
rect 2406 1420 2407 1424
rect 2411 1420 2412 1424
rect 2406 1419 2412 1420
rect 110 1416 116 1417
rect 110 1412 111 1416
rect 115 1412 116 1416
rect 110 1411 116 1412
rect 1238 1416 1244 1417
rect 1238 1412 1239 1416
rect 1243 1412 1244 1416
rect 1238 1411 1244 1412
rect 1278 1407 1284 1408
rect 1278 1403 1279 1407
rect 1283 1403 1284 1407
rect 1278 1402 1284 1403
rect 2406 1407 2412 1408
rect 2406 1403 2407 1407
rect 2411 1403 2412 1407
rect 2406 1402 2412 1403
rect 110 1399 116 1400
rect 110 1395 111 1399
rect 115 1395 116 1399
rect 110 1394 116 1395
rect 1238 1399 1244 1400
rect 1238 1395 1239 1399
rect 1243 1395 1244 1399
rect 1238 1394 1244 1395
rect 112 1387 114 1394
rect 142 1392 148 1393
rect 142 1388 143 1392
rect 147 1388 148 1392
rect 142 1387 148 1388
rect 182 1392 188 1393
rect 182 1388 183 1392
rect 187 1388 188 1392
rect 182 1387 188 1388
rect 222 1392 228 1393
rect 222 1388 223 1392
rect 227 1388 228 1392
rect 222 1387 228 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 318 1392 324 1393
rect 318 1388 319 1392
rect 323 1388 324 1392
rect 318 1387 324 1388
rect 390 1392 396 1393
rect 390 1388 391 1392
rect 395 1388 396 1392
rect 390 1387 396 1388
rect 470 1392 476 1393
rect 470 1388 471 1392
rect 475 1388 476 1392
rect 470 1387 476 1388
rect 558 1392 564 1393
rect 558 1388 559 1392
rect 563 1388 564 1392
rect 558 1387 564 1388
rect 646 1392 652 1393
rect 646 1388 647 1392
rect 651 1388 652 1392
rect 646 1387 652 1388
rect 726 1392 732 1393
rect 726 1388 727 1392
rect 731 1388 732 1392
rect 726 1387 732 1388
rect 806 1392 812 1393
rect 806 1388 807 1392
rect 811 1388 812 1392
rect 806 1387 812 1388
rect 878 1392 884 1393
rect 878 1388 879 1392
rect 883 1388 884 1392
rect 878 1387 884 1388
rect 942 1392 948 1393
rect 942 1388 943 1392
rect 947 1388 948 1392
rect 942 1387 948 1388
rect 998 1392 1004 1393
rect 998 1388 999 1392
rect 1003 1388 1004 1392
rect 998 1387 1004 1388
rect 1046 1392 1052 1393
rect 1046 1388 1047 1392
rect 1051 1388 1052 1392
rect 1046 1387 1052 1388
rect 1102 1392 1108 1393
rect 1102 1388 1103 1392
rect 1107 1388 1108 1392
rect 1102 1387 1108 1388
rect 1150 1392 1156 1393
rect 1150 1388 1151 1392
rect 1155 1388 1156 1392
rect 1150 1387 1156 1388
rect 1190 1392 1196 1393
rect 1190 1388 1191 1392
rect 1195 1388 1196 1392
rect 1190 1387 1196 1388
rect 1240 1387 1242 1394
rect 1280 1387 1282 1402
rect 1374 1400 1380 1401
rect 1374 1396 1375 1400
rect 1379 1396 1380 1400
rect 1374 1395 1380 1396
rect 1462 1400 1468 1401
rect 1462 1396 1463 1400
rect 1467 1396 1468 1400
rect 1462 1395 1468 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1806 1400 1812 1401
rect 1806 1396 1807 1400
rect 1811 1396 1812 1400
rect 1806 1395 1812 1396
rect 1878 1400 1884 1401
rect 1878 1396 1879 1400
rect 1883 1396 1884 1400
rect 1878 1395 1884 1396
rect 1942 1400 1948 1401
rect 1942 1396 1943 1400
rect 1947 1396 1948 1400
rect 1942 1395 1948 1396
rect 1998 1400 2004 1401
rect 1998 1396 1999 1400
rect 2003 1396 2004 1400
rect 1998 1395 2004 1396
rect 2046 1400 2052 1401
rect 2046 1396 2047 1400
rect 2051 1396 2052 1400
rect 2046 1395 2052 1396
rect 2094 1400 2100 1401
rect 2094 1396 2095 1400
rect 2099 1396 2100 1400
rect 2094 1395 2100 1396
rect 2142 1400 2148 1401
rect 2142 1396 2143 1400
rect 2147 1396 2148 1400
rect 2142 1395 2148 1396
rect 2190 1400 2196 1401
rect 2190 1396 2191 1400
rect 2195 1396 2196 1400
rect 2190 1395 2196 1396
rect 2238 1400 2244 1401
rect 2238 1396 2239 1400
rect 2243 1396 2244 1400
rect 2238 1395 2244 1396
rect 2278 1400 2284 1401
rect 2278 1396 2279 1400
rect 2283 1396 2284 1400
rect 2278 1395 2284 1396
rect 2318 1400 2324 1401
rect 2318 1396 2319 1400
rect 2323 1396 2324 1400
rect 2318 1395 2324 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 1376 1387 1378 1395
rect 1464 1387 1466 1395
rect 1552 1387 1554 1395
rect 1640 1387 1642 1395
rect 1728 1387 1730 1395
rect 1808 1387 1810 1395
rect 1880 1387 1882 1395
rect 1944 1387 1946 1395
rect 2000 1387 2002 1395
rect 2048 1387 2050 1395
rect 2096 1387 2098 1395
rect 2144 1387 2146 1395
rect 2192 1387 2194 1395
rect 2240 1387 2242 1395
rect 2280 1387 2282 1395
rect 2320 1387 2322 1395
rect 2360 1387 2362 1395
rect 2408 1387 2410 1402
rect 111 1386 115 1387
rect 111 1381 115 1382
rect 143 1386 147 1387
rect 143 1381 147 1382
rect 167 1386 171 1387
rect 167 1381 171 1382
rect 183 1386 187 1387
rect 183 1381 187 1382
rect 207 1386 211 1387
rect 207 1381 211 1382
rect 223 1386 227 1387
rect 223 1381 227 1382
rect 247 1386 251 1387
rect 247 1381 251 1382
rect 263 1386 267 1387
rect 263 1381 267 1382
rect 303 1386 307 1387
rect 303 1381 307 1382
rect 319 1386 323 1387
rect 319 1381 323 1382
rect 367 1386 371 1387
rect 367 1381 371 1382
rect 391 1386 395 1387
rect 391 1381 395 1382
rect 439 1386 443 1387
rect 439 1381 443 1382
rect 471 1386 475 1387
rect 471 1381 475 1382
rect 519 1386 523 1387
rect 519 1381 523 1382
rect 559 1386 563 1387
rect 559 1381 563 1382
rect 599 1386 603 1387
rect 599 1381 603 1382
rect 647 1386 651 1387
rect 647 1381 651 1382
rect 679 1386 683 1387
rect 679 1381 683 1382
rect 727 1386 731 1387
rect 727 1381 731 1382
rect 751 1386 755 1387
rect 751 1381 755 1382
rect 807 1386 811 1387
rect 807 1381 811 1382
rect 823 1386 827 1387
rect 823 1381 827 1382
rect 879 1386 883 1387
rect 879 1381 883 1382
rect 887 1386 891 1387
rect 887 1381 891 1382
rect 943 1386 947 1387
rect 943 1381 947 1382
rect 951 1386 955 1387
rect 951 1381 955 1382
rect 999 1386 1003 1387
rect 999 1381 1003 1382
rect 1015 1386 1019 1387
rect 1015 1381 1019 1382
rect 1047 1386 1051 1387
rect 1047 1381 1051 1382
rect 1079 1386 1083 1387
rect 1079 1381 1083 1382
rect 1103 1386 1107 1387
rect 1103 1381 1107 1382
rect 1143 1386 1147 1387
rect 1143 1381 1147 1382
rect 1151 1386 1155 1387
rect 1151 1381 1155 1382
rect 1191 1386 1195 1387
rect 1191 1381 1195 1382
rect 1239 1386 1243 1387
rect 1239 1381 1243 1382
rect 1279 1386 1283 1387
rect 1279 1381 1283 1382
rect 1303 1386 1307 1387
rect 1303 1381 1307 1382
rect 1343 1386 1347 1387
rect 1343 1381 1347 1382
rect 1375 1386 1379 1387
rect 1375 1381 1379 1382
rect 1399 1386 1403 1387
rect 1399 1381 1403 1382
rect 1463 1386 1467 1387
rect 1463 1381 1467 1382
rect 1535 1386 1539 1387
rect 1535 1381 1539 1382
rect 1551 1386 1555 1387
rect 1551 1381 1555 1382
rect 1607 1386 1611 1387
rect 1607 1381 1611 1382
rect 1639 1386 1643 1387
rect 1639 1381 1643 1382
rect 1687 1386 1691 1387
rect 1687 1381 1691 1382
rect 1727 1386 1731 1387
rect 1727 1381 1731 1382
rect 1767 1386 1771 1387
rect 1767 1381 1771 1382
rect 1807 1386 1811 1387
rect 1807 1381 1811 1382
rect 1847 1386 1851 1387
rect 1847 1381 1851 1382
rect 1879 1386 1883 1387
rect 1879 1381 1883 1382
rect 1935 1386 1939 1387
rect 1935 1381 1939 1382
rect 1943 1386 1947 1387
rect 1943 1381 1947 1382
rect 1999 1386 2003 1387
rect 1999 1381 2003 1382
rect 2023 1386 2027 1387
rect 2023 1381 2027 1382
rect 2047 1386 2051 1387
rect 2047 1381 2051 1382
rect 2095 1386 2099 1387
rect 2095 1381 2099 1382
rect 2111 1386 2115 1387
rect 2111 1381 2115 1382
rect 2143 1386 2147 1387
rect 2143 1381 2147 1382
rect 2191 1386 2195 1387
rect 2191 1381 2195 1382
rect 2199 1386 2203 1387
rect 2199 1381 2203 1382
rect 2239 1386 2243 1387
rect 2239 1381 2243 1382
rect 2279 1386 2283 1387
rect 2279 1381 2283 1382
rect 2287 1386 2291 1387
rect 2287 1381 2291 1382
rect 2319 1386 2323 1387
rect 2319 1381 2323 1382
rect 2359 1386 2363 1387
rect 2359 1381 2363 1382
rect 2407 1386 2411 1387
rect 2407 1381 2411 1382
rect 112 1374 114 1381
rect 166 1380 172 1381
rect 166 1376 167 1380
rect 171 1376 172 1380
rect 166 1375 172 1376
rect 206 1380 212 1381
rect 206 1376 207 1380
rect 211 1376 212 1380
rect 206 1375 212 1376
rect 246 1380 252 1381
rect 246 1376 247 1380
rect 251 1376 252 1380
rect 246 1375 252 1376
rect 302 1380 308 1381
rect 302 1376 303 1380
rect 307 1376 308 1380
rect 302 1375 308 1376
rect 366 1380 372 1381
rect 366 1376 367 1380
rect 371 1376 372 1380
rect 366 1375 372 1376
rect 438 1380 444 1381
rect 438 1376 439 1380
rect 443 1376 444 1380
rect 438 1375 444 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 598 1380 604 1381
rect 598 1376 599 1380
rect 603 1376 604 1380
rect 598 1375 604 1376
rect 678 1380 684 1381
rect 678 1376 679 1380
rect 683 1376 684 1380
rect 678 1375 684 1376
rect 750 1380 756 1381
rect 750 1376 751 1380
rect 755 1376 756 1380
rect 750 1375 756 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 886 1380 892 1381
rect 886 1376 887 1380
rect 891 1376 892 1380
rect 886 1375 892 1376
rect 950 1380 956 1381
rect 950 1376 951 1380
rect 955 1376 956 1380
rect 950 1375 956 1376
rect 1014 1380 1020 1381
rect 1014 1376 1015 1380
rect 1019 1376 1020 1380
rect 1014 1375 1020 1376
rect 1078 1380 1084 1381
rect 1078 1376 1079 1380
rect 1083 1376 1084 1380
rect 1078 1375 1084 1376
rect 1142 1380 1148 1381
rect 1142 1376 1143 1380
rect 1147 1376 1148 1380
rect 1142 1375 1148 1376
rect 1190 1380 1196 1381
rect 1190 1376 1191 1380
rect 1195 1376 1196 1380
rect 1190 1375 1196 1376
rect 1240 1374 1242 1381
rect 1280 1374 1282 1381
rect 1302 1380 1308 1381
rect 1302 1376 1303 1380
rect 1307 1376 1308 1380
rect 1302 1375 1308 1376
rect 1342 1380 1348 1381
rect 1342 1376 1343 1380
rect 1347 1376 1348 1380
rect 1342 1375 1348 1376
rect 1398 1380 1404 1381
rect 1398 1376 1399 1380
rect 1403 1376 1404 1380
rect 1398 1375 1404 1376
rect 1462 1380 1468 1381
rect 1462 1376 1463 1380
rect 1467 1376 1468 1380
rect 1462 1375 1468 1376
rect 1534 1380 1540 1381
rect 1534 1376 1535 1380
rect 1539 1376 1540 1380
rect 1534 1375 1540 1376
rect 1606 1380 1612 1381
rect 1606 1376 1607 1380
rect 1611 1376 1612 1380
rect 1606 1375 1612 1376
rect 1686 1380 1692 1381
rect 1686 1376 1687 1380
rect 1691 1376 1692 1380
rect 1686 1375 1692 1376
rect 1766 1380 1772 1381
rect 1766 1376 1767 1380
rect 1771 1376 1772 1380
rect 1766 1375 1772 1376
rect 1846 1380 1852 1381
rect 1846 1376 1847 1380
rect 1851 1376 1852 1380
rect 1846 1375 1852 1376
rect 1934 1380 1940 1381
rect 1934 1376 1935 1380
rect 1939 1376 1940 1380
rect 1934 1375 1940 1376
rect 2022 1380 2028 1381
rect 2022 1376 2023 1380
rect 2027 1376 2028 1380
rect 2022 1375 2028 1376
rect 2110 1380 2116 1381
rect 2110 1376 2111 1380
rect 2115 1376 2116 1380
rect 2110 1375 2116 1376
rect 2198 1380 2204 1381
rect 2198 1376 2199 1380
rect 2203 1376 2204 1380
rect 2198 1375 2204 1376
rect 2286 1380 2292 1381
rect 2286 1376 2287 1380
rect 2291 1376 2292 1380
rect 2286 1375 2292 1376
rect 2358 1380 2364 1381
rect 2358 1376 2359 1380
rect 2363 1376 2364 1380
rect 2358 1375 2364 1376
rect 2408 1374 2410 1381
rect 110 1373 116 1374
rect 110 1369 111 1373
rect 115 1369 116 1373
rect 110 1368 116 1369
rect 1238 1373 1244 1374
rect 1238 1369 1239 1373
rect 1243 1369 1244 1373
rect 1238 1368 1244 1369
rect 1278 1373 1284 1374
rect 1278 1369 1279 1373
rect 1283 1369 1284 1373
rect 1278 1368 1284 1369
rect 2406 1373 2412 1374
rect 2406 1369 2407 1373
rect 2411 1369 2412 1373
rect 2406 1368 2412 1369
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 110 1351 116 1352
rect 1238 1356 1244 1357
rect 1238 1352 1239 1356
rect 1243 1352 1244 1356
rect 1238 1351 1244 1352
rect 1278 1356 1284 1357
rect 1278 1352 1279 1356
rect 1283 1352 1284 1356
rect 1278 1351 1284 1352
rect 2406 1356 2412 1357
rect 2406 1352 2407 1356
rect 2411 1352 2412 1356
rect 2406 1351 2412 1352
rect 112 1315 114 1351
rect 166 1333 172 1334
rect 166 1329 167 1333
rect 171 1329 172 1333
rect 166 1328 172 1329
rect 206 1333 212 1334
rect 206 1329 207 1333
rect 211 1329 212 1333
rect 206 1328 212 1329
rect 246 1333 252 1334
rect 246 1329 247 1333
rect 251 1329 252 1333
rect 246 1328 252 1329
rect 302 1333 308 1334
rect 302 1329 303 1333
rect 307 1329 308 1333
rect 302 1328 308 1329
rect 366 1333 372 1334
rect 366 1329 367 1333
rect 371 1329 372 1333
rect 366 1328 372 1329
rect 438 1333 444 1334
rect 438 1329 439 1333
rect 443 1329 444 1333
rect 438 1328 444 1329
rect 518 1333 524 1334
rect 518 1329 519 1333
rect 523 1329 524 1333
rect 518 1328 524 1329
rect 598 1333 604 1334
rect 598 1329 599 1333
rect 603 1329 604 1333
rect 598 1328 604 1329
rect 678 1333 684 1334
rect 678 1329 679 1333
rect 683 1329 684 1333
rect 678 1328 684 1329
rect 750 1333 756 1334
rect 750 1329 751 1333
rect 755 1329 756 1333
rect 750 1328 756 1329
rect 822 1333 828 1334
rect 822 1329 823 1333
rect 827 1329 828 1333
rect 822 1328 828 1329
rect 886 1333 892 1334
rect 886 1329 887 1333
rect 891 1329 892 1333
rect 886 1328 892 1329
rect 950 1333 956 1334
rect 950 1329 951 1333
rect 955 1329 956 1333
rect 950 1328 956 1329
rect 1014 1333 1020 1334
rect 1014 1329 1015 1333
rect 1019 1329 1020 1333
rect 1014 1328 1020 1329
rect 1078 1333 1084 1334
rect 1078 1329 1079 1333
rect 1083 1329 1084 1333
rect 1078 1328 1084 1329
rect 1142 1333 1148 1334
rect 1142 1329 1143 1333
rect 1147 1329 1148 1333
rect 1142 1328 1148 1329
rect 1190 1333 1196 1334
rect 1190 1329 1191 1333
rect 1195 1329 1196 1333
rect 1190 1328 1196 1329
rect 168 1315 170 1328
rect 208 1315 210 1328
rect 248 1315 250 1328
rect 304 1315 306 1328
rect 368 1315 370 1328
rect 440 1315 442 1328
rect 520 1315 522 1328
rect 600 1315 602 1328
rect 680 1315 682 1328
rect 752 1315 754 1328
rect 824 1315 826 1328
rect 888 1315 890 1328
rect 952 1315 954 1328
rect 1016 1315 1018 1328
rect 1080 1315 1082 1328
rect 1144 1315 1146 1328
rect 1192 1315 1194 1328
rect 1240 1315 1242 1351
rect 1280 1319 1282 1351
rect 1302 1333 1308 1334
rect 1302 1329 1303 1333
rect 1307 1329 1308 1333
rect 1302 1328 1308 1329
rect 1342 1333 1348 1334
rect 1342 1329 1343 1333
rect 1347 1329 1348 1333
rect 1342 1328 1348 1329
rect 1398 1333 1404 1334
rect 1398 1329 1399 1333
rect 1403 1329 1404 1333
rect 1398 1328 1404 1329
rect 1462 1333 1468 1334
rect 1462 1329 1463 1333
rect 1467 1329 1468 1333
rect 1462 1328 1468 1329
rect 1534 1333 1540 1334
rect 1534 1329 1535 1333
rect 1539 1329 1540 1333
rect 1534 1328 1540 1329
rect 1606 1333 1612 1334
rect 1606 1329 1607 1333
rect 1611 1329 1612 1333
rect 1606 1328 1612 1329
rect 1686 1333 1692 1334
rect 1686 1329 1687 1333
rect 1691 1329 1692 1333
rect 1686 1328 1692 1329
rect 1766 1333 1772 1334
rect 1766 1329 1767 1333
rect 1771 1329 1772 1333
rect 1766 1328 1772 1329
rect 1846 1333 1852 1334
rect 1846 1329 1847 1333
rect 1851 1329 1852 1333
rect 1846 1328 1852 1329
rect 1934 1333 1940 1334
rect 1934 1329 1935 1333
rect 1939 1329 1940 1333
rect 1934 1328 1940 1329
rect 2022 1333 2028 1334
rect 2022 1329 2023 1333
rect 2027 1329 2028 1333
rect 2022 1328 2028 1329
rect 2110 1333 2116 1334
rect 2110 1329 2111 1333
rect 2115 1329 2116 1333
rect 2110 1328 2116 1329
rect 2198 1333 2204 1334
rect 2198 1329 2199 1333
rect 2203 1329 2204 1333
rect 2198 1328 2204 1329
rect 2286 1333 2292 1334
rect 2286 1329 2287 1333
rect 2291 1329 2292 1333
rect 2286 1328 2292 1329
rect 2358 1333 2364 1334
rect 2358 1329 2359 1333
rect 2363 1329 2364 1333
rect 2358 1328 2364 1329
rect 1304 1319 1306 1328
rect 1344 1319 1346 1328
rect 1400 1319 1402 1328
rect 1464 1319 1466 1328
rect 1536 1319 1538 1328
rect 1608 1319 1610 1328
rect 1688 1319 1690 1328
rect 1768 1319 1770 1328
rect 1848 1319 1850 1328
rect 1936 1319 1938 1328
rect 2024 1319 2026 1328
rect 2112 1319 2114 1328
rect 2200 1319 2202 1328
rect 2288 1319 2290 1328
rect 2360 1319 2362 1328
rect 2408 1319 2410 1351
rect 1279 1318 1283 1319
rect 111 1314 115 1315
rect 111 1309 115 1310
rect 167 1314 171 1315
rect 167 1309 171 1310
rect 183 1314 187 1315
rect 183 1309 187 1310
rect 207 1314 211 1315
rect 207 1309 211 1310
rect 231 1314 235 1315
rect 231 1309 235 1310
rect 247 1314 251 1315
rect 247 1309 251 1310
rect 287 1314 291 1315
rect 287 1309 291 1310
rect 303 1314 307 1315
rect 303 1309 307 1310
rect 351 1314 355 1315
rect 351 1309 355 1310
rect 367 1314 371 1315
rect 367 1309 371 1310
rect 423 1314 427 1315
rect 423 1309 427 1310
rect 439 1314 443 1315
rect 439 1309 443 1310
rect 495 1314 499 1315
rect 495 1309 499 1310
rect 519 1314 523 1315
rect 519 1309 523 1310
rect 567 1314 571 1315
rect 567 1309 571 1310
rect 599 1314 603 1315
rect 599 1309 603 1310
rect 639 1314 643 1315
rect 639 1309 643 1310
rect 679 1314 683 1315
rect 679 1309 683 1310
rect 703 1314 707 1315
rect 703 1309 707 1310
rect 751 1314 755 1315
rect 751 1309 755 1310
rect 767 1314 771 1315
rect 767 1309 771 1310
rect 823 1314 827 1315
rect 823 1309 827 1310
rect 879 1314 883 1315
rect 879 1309 883 1310
rect 887 1314 891 1315
rect 887 1309 891 1310
rect 935 1314 939 1315
rect 935 1309 939 1310
rect 951 1314 955 1315
rect 951 1309 955 1310
rect 999 1314 1003 1315
rect 999 1309 1003 1310
rect 1015 1314 1019 1315
rect 1015 1309 1019 1310
rect 1079 1314 1083 1315
rect 1079 1309 1083 1310
rect 1143 1314 1147 1315
rect 1143 1309 1147 1310
rect 1191 1314 1195 1315
rect 1191 1309 1195 1310
rect 1239 1314 1243 1315
rect 1279 1313 1283 1314
rect 1303 1318 1307 1319
rect 1303 1313 1307 1314
rect 1343 1318 1347 1319
rect 1343 1313 1347 1314
rect 1383 1318 1387 1319
rect 1383 1313 1387 1314
rect 1399 1318 1403 1319
rect 1399 1313 1403 1314
rect 1423 1318 1427 1319
rect 1423 1313 1427 1314
rect 1463 1318 1467 1319
rect 1463 1313 1467 1314
rect 1503 1318 1507 1319
rect 1503 1313 1507 1314
rect 1535 1318 1539 1319
rect 1535 1313 1539 1314
rect 1543 1318 1547 1319
rect 1543 1313 1547 1314
rect 1583 1318 1587 1319
rect 1583 1313 1587 1314
rect 1607 1318 1611 1319
rect 1607 1313 1611 1314
rect 1623 1318 1627 1319
rect 1623 1313 1627 1314
rect 1679 1318 1683 1319
rect 1679 1313 1683 1314
rect 1687 1318 1691 1319
rect 1687 1313 1691 1314
rect 1735 1318 1739 1319
rect 1735 1313 1739 1314
rect 1767 1318 1771 1319
rect 1767 1313 1771 1314
rect 1791 1318 1795 1319
rect 1791 1313 1795 1314
rect 1847 1318 1851 1319
rect 1847 1313 1851 1314
rect 1903 1318 1907 1319
rect 1903 1313 1907 1314
rect 1935 1318 1939 1319
rect 1935 1313 1939 1314
rect 1967 1318 1971 1319
rect 1967 1313 1971 1314
rect 2023 1318 2027 1319
rect 2023 1313 2027 1314
rect 2039 1318 2043 1319
rect 2039 1313 2043 1314
rect 2111 1318 2115 1319
rect 2111 1313 2115 1314
rect 2119 1318 2123 1319
rect 2119 1313 2123 1314
rect 2199 1318 2203 1319
rect 2199 1313 2203 1314
rect 2287 1318 2291 1319
rect 2287 1313 2291 1314
rect 2359 1318 2363 1319
rect 2359 1313 2363 1314
rect 2407 1318 2411 1319
rect 2407 1313 2411 1314
rect 1239 1309 1243 1310
rect 112 1277 114 1309
rect 184 1300 186 1309
rect 232 1300 234 1309
rect 288 1300 290 1309
rect 352 1300 354 1309
rect 424 1300 426 1309
rect 496 1300 498 1309
rect 568 1300 570 1309
rect 640 1300 642 1309
rect 704 1300 706 1309
rect 768 1300 770 1309
rect 824 1300 826 1309
rect 880 1300 882 1309
rect 936 1300 938 1309
rect 1000 1300 1002 1309
rect 182 1299 188 1300
rect 182 1295 183 1299
rect 187 1295 188 1299
rect 182 1294 188 1295
rect 230 1299 236 1300
rect 230 1295 231 1299
rect 235 1295 236 1299
rect 230 1294 236 1295
rect 286 1299 292 1300
rect 286 1295 287 1299
rect 291 1295 292 1299
rect 286 1294 292 1295
rect 350 1299 356 1300
rect 350 1295 351 1299
rect 355 1295 356 1299
rect 350 1294 356 1295
rect 422 1299 428 1300
rect 422 1295 423 1299
rect 427 1295 428 1299
rect 422 1294 428 1295
rect 494 1299 500 1300
rect 494 1295 495 1299
rect 499 1295 500 1299
rect 494 1294 500 1295
rect 566 1299 572 1300
rect 566 1295 567 1299
rect 571 1295 572 1299
rect 566 1294 572 1295
rect 638 1299 644 1300
rect 638 1295 639 1299
rect 643 1295 644 1299
rect 638 1294 644 1295
rect 702 1299 708 1300
rect 702 1295 703 1299
rect 707 1295 708 1299
rect 702 1294 708 1295
rect 766 1299 772 1300
rect 766 1295 767 1299
rect 771 1295 772 1299
rect 766 1294 772 1295
rect 822 1299 828 1300
rect 822 1295 823 1299
rect 827 1295 828 1299
rect 822 1294 828 1295
rect 878 1299 884 1300
rect 878 1295 879 1299
rect 883 1295 884 1299
rect 878 1294 884 1295
rect 934 1299 940 1300
rect 934 1295 935 1299
rect 939 1295 940 1299
rect 934 1294 940 1295
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1295 1004 1299
rect 998 1294 1004 1295
rect 1240 1277 1242 1309
rect 1280 1281 1282 1313
rect 1304 1304 1306 1313
rect 1344 1304 1346 1313
rect 1384 1304 1386 1313
rect 1424 1304 1426 1313
rect 1464 1304 1466 1313
rect 1504 1304 1506 1313
rect 1544 1304 1546 1313
rect 1584 1304 1586 1313
rect 1624 1304 1626 1313
rect 1680 1304 1682 1313
rect 1736 1304 1738 1313
rect 1792 1304 1794 1313
rect 1848 1304 1850 1313
rect 1904 1304 1906 1313
rect 1968 1304 1970 1313
rect 2040 1304 2042 1313
rect 2120 1304 2122 1313
rect 2200 1304 2202 1313
rect 2288 1304 2290 1313
rect 2360 1304 2362 1313
rect 1302 1303 1308 1304
rect 1302 1299 1303 1303
rect 1307 1299 1308 1303
rect 1302 1298 1308 1299
rect 1342 1303 1348 1304
rect 1342 1299 1343 1303
rect 1347 1299 1348 1303
rect 1342 1298 1348 1299
rect 1382 1303 1388 1304
rect 1382 1299 1383 1303
rect 1387 1299 1388 1303
rect 1382 1298 1388 1299
rect 1422 1303 1428 1304
rect 1422 1299 1423 1303
rect 1427 1299 1428 1303
rect 1422 1298 1428 1299
rect 1462 1303 1468 1304
rect 1462 1299 1463 1303
rect 1467 1299 1468 1303
rect 1462 1298 1468 1299
rect 1502 1303 1508 1304
rect 1502 1299 1503 1303
rect 1507 1299 1508 1303
rect 1502 1298 1508 1299
rect 1542 1303 1548 1304
rect 1542 1299 1543 1303
rect 1547 1299 1548 1303
rect 1542 1298 1548 1299
rect 1582 1303 1588 1304
rect 1582 1299 1583 1303
rect 1587 1299 1588 1303
rect 1582 1298 1588 1299
rect 1622 1303 1628 1304
rect 1622 1299 1623 1303
rect 1627 1299 1628 1303
rect 1622 1298 1628 1299
rect 1678 1303 1684 1304
rect 1678 1299 1679 1303
rect 1683 1299 1684 1303
rect 1678 1298 1684 1299
rect 1734 1303 1740 1304
rect 1734 1299 1735 1303
rect 1739 1299 1740 1303
rect 1734 1298 1740 1299
rect 1790 1303 1796 1304
rect 1790 1299 1791 1303
rect 1795 1299 1796 1303
rect 1790 1298 1796 1299
rect 1846 1303 1852 1304
rect 1846 1299 1847 1303
rect 1851 1299 1852 1303
rect 1846 1298 1852 1299
rect 1902 1303 1908 1304
rect 1902 1299 1903 1303
rect 1907 1299 1908 1303
rect 1902 1298 1908 1299
rect 1966 1303 1972 1304
rect 1966 1299 1967 1303
rect 1971 1299 1972 1303
rect 1966 1298 1972 1299
rect 2038 1303 2044 1304
rect 2038 1299 2039 1303
rect 2043 1299 2044 1303
rect 2038 1298 2044 1299
rect 2118 1303 2124 1304
rect 2118 1299 2119 1303
rect 2123 1299 2124 1303
rect 2118 1298 2124 1299
rect 2198 1303 2204 1304
rect 2198 1299 2199 1303
rect 2203 1299 2204 1303
rect 2198 1298 2204 1299
rect 2286 1303 2292 1304
rect 2286 1299 2287 1303
rect 2291 1299 2292 1303
rect 2286 1298 2292 1299
rect 2358 1303 2364 1304
rect 2358 1299 2359 1303
rect 2363 1299 2364 1303
rect 2358 1298 2364 1299
rect 2408 1281 2410 1313
rect 1278 1280 1284 1281
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 110 1271 116 1272
rect 1238 1276 1244 1277
rect 1238 1272 1239 1276
rect 1243 1272 1244 1276
rect 1278 1276 1279 1280
rect 1283 1276 1284 1280
rect 1278 1275 1284 1276
rect 2406 1280 2412 1281
rect 2406 1276 2407 1280
rect 2411 1276 2412 1280
rect 2406 1275 2412 1276
rect 1238 1271 1244 1272
rect 1278 1263 1284 1264
rect 110 1259 116 1260
rect 110 1255 111 1259
rect 115 1255 116 1259
rect 110 1254 116 1255
rect 1238 1259 1244 1260
rect 1238 1255 1239 1259
rect 1243 1255 1244 1259
rect 1278 1259 1279 1263
rect 1283 1259 1284 1263
rect 1278 1258 1284 1259
rect 2406 1263 2412 1264
rect 2406 1259 2407 1263
rect 2411 1259 2412 1263
rect 2406 1258 2412 1259
rect 1238 1254 1244 1255
rect 112 1243 114 1254
rect 182 1252 188 1253
rect 182 1248 183 1252
rect 187 1248 188 1252
rect 182 1247 188 1248
rect 230 1252 236 1253
rect 230 1248 231 1252
rect 235 1248 236 1252
rect 230 1247 236 1248
rect 286 1252 292 1253
rect 286 1248 287 1252
rect 291 1248 292 1252
rect 286 1247 292 1248
rect 350 1252 356 1253
rect 350 1248 351 1252
rect 355 1248 356 1252
rect 350 1247 356 1248
rect 422 1252 428 1253
rect 422 1248 423 1252
rect 427 1248 428 1252
rect 422 1247 428 1248
rect 494 1252 500 1253
rect 494 1248 495 1252
rect 499 1248 500 1252
rect 494 1247 500 1248
rect 566 1252 572 1253
rect 566 1248 567 1252
rect 571 1248 572 1252
rect 566 1247 572 1248
rect 638 1252 644 1253
rect 638 1248 639 1252
rect 643 1248 644 1252
rect 638 1247 644 1248
rect 702 1252 708 1253
rect 702 1248 703 1252
rect 707 1248 708 1252
rect 702 1247 708 1248
rect 766 1252 772 1253
rect 766 1248 767 1252
rect 771 1248 772 1252
rect 766 1247 772 1248
rect 822 1252 828 1253
rect 822 1248 823 1252
rect 827 1248 828 1252
rect 822 1247 828 1248
rect 878 1252 884 1253
rect 878 1248 879 1252
rect 883 1248 884 1252
rect 878 1247 884 1248
rect 934 1252 940 1253
rect 934 1248 935 1252
rect 939 1248 940 1252
rect 934 1247 940 1248
rect 998 1252 1004 1253
rect 998 1248 999 1252
rect 1003 1248 1004 1252
rect 998 1247 1004 1248
rect 184 1243 186 1247
rect 232 1243 234 1247
rect 288 1243 290 1247
rect 352 1243 354 1247
rect 424 1243 426 1247
rect 496 1243 498 1247
rect 568 1243 570 1247
rect 640 1243 642 1247
rect 704 1243 706 1247
rect 768 1243 770 1247
rect 824 1243 826 1247
rect 880 1243 882 1247
rect 936 1243 938 1247
rect 1000 1243 1002 1247
rect 1240 1243 1242 1254
rect 1280 1243 1282 1258
rect 1302 1256 1308 1257
rect 1302 1252 1303 1256
rect 1307 1252 1308 1256
rect 1302 1251 1308 1252
rect 1342 1256 1348 1257
rect 1342 1252 1343 1256
rect 1347 1252 1348 1256
rect 1342 1251 1348 1252
rect 1382 1256 1388 1257
rect 1382 1252 1383 1256
rect 1387 1252 1388 1256
rect 1382 1251 1388 1252
rect 1422 1256 1428 1257
rect 1422 1252 1423 1256
rect 1427 1252 1428 1256
rect 1422 1251 1428 1252
rect 1462 1256 1468 1257
rect 1462 1252 1463 1256
rect 1467 1252 1468 1256
rect 1462 1251 1468 1252
rect 1502 1256 1508 1257
rect 1502 1252 1503 1256
rect 1507 1252 1508 1256
rect 1502 1251 1508 1252
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1582 1256 1588 1257
rect 1582 1252 1583 1256
rect 1587 1252 1588 1256
rect 1582 1251 1588 1252
rect 1622 1256 1628 1257
rect 1622 1252 1623 1256
rect 1627 1252 1628 1256
rect 1622 1251 1628 1252
rect 1678 1256 1684 1257
rect 1678 1252 1679 1256
rect 1683 1252 1684 1256
rect 1678 1251 1684 1252
rect 1734 1256 1740 1257
rect 1734 1252 1735 1256
rect 1739 1252 1740 1256
rect 1734 1251 1740 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1846 1256 1852 1257
rect 1846 1252 1847 1256
rect 1851 1252 1852 1256
rect 1846 1251 1852 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2198 1256 2204 1257
rect 2198 1252 2199 1256
rect 2203 1252 2204 1256
rect 2198 1251 2204 1252
rect 2286 1256 2292 1257
rect 2286 1252 2287 1256
rect 2291 1252 2292 1256
rect 2286 1251 2292 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 1304 1243 1306 1251
rect 1344 1243 1346 1251
rect 1384 1243 1386 1251
rect 1424 1243 1426 1251
rect 1464 1243 1466 1251
rect 1504 1243 1506 1251
rect 1544 1243 1546 1251
rect 1584 1243 1586 1251
rect 1624 1243 1626 1251
rect 1680 1243 1682 1251
rect 1736 1243 1738 1251
rect 1792 1243 1794 1251
rect 1848 1243 1850 1251
rect 1904 1243 1906 1251
rect 1968 1243 1970 1251
rect 2040 1243 2042 1251
rect 2120 1243 2122 1251
rect 2200 1243 2202 1251
rect 2288 1243 2290 1251
rect 2360 1243 2362 1251
rect 2408 1243 2410 1258
rect 111 1242 115 1243
rect 111 1237 115 1238
rect 135 1242 139 1243
rect 135 1237 139 1238
rect 175 1242 179 1243
rect 175 1237 179 1238
rect 183 1242 187 1243
rect 183 1237 187 1238
rect 231 1242 235 1243
rect 231 1237 235 1238
rect 287 1242 291 1243
rect 287 1237 291 1238
rect 311 1242 315 1243
rect 311 1237 315 1238
rect 351 1242 355 1243
rect 351 1237 355 1238
rect 399 1242 403 1243
rect 399 1237 403 1238
rect 423 1242 427 1243
rect 423 1237 427 1238
rect 487 1242 491 1243
rect 487 1237 491 1238
rect 495 1242 499 1243
rect 495 1237 499 1238
rect 567 1242 571 1243
rect 567 1237 571 1238
rect 575 1242 579 1243
rect 575 1237 579 1238
rect 639 1242 643 1243
rect 639 1237 643 1238
rect 663 1242 667 1243
rect 663 1237 667 1238
rect 703 1242 707 1243
rect 703 1237 707 1238
rect 743 1242 747 1243
rect 743 1237 747 1238
rect 767 1242 771 1243
rect 767 1237 771 1238
rect 815 1242 819 1243
rect 815 1237 819 1238
rect 823 1242 827 1243
rect 823 1237 827 1238
rect 879 1242 883 1243
rect 879 1237 883 1238
rect 935 1242 939 1243
rect 935 1237 939 1238
rect 943 1242 947 1243
rect 943 1237 947 1238
rect 999 1242 1003 1243
rect 999 1237 1003 1238
rect 1007 1242 1011 1243
rect 1007 1237 1011 1238
rect 1071 1242 1075 1243
rect 1071 1237 1075 1238
rect 1239 1242 1243 1243
rect 1239 1237 1243 1238
rect 1279 1242 1283 1243
rect 1279 1237 1283 1238
rect 1303 1242 1307 1243
rect 1303 1237 1307 1238
rect 1343 1242 1347 1243
rect 1343 1237 1347 1238
rect 1375 1242 1379 1243
rect 1375 1237 1379 1238
rect 1383 1242 1387 1243
rect 1383 1237 1387 1238
rect 1423 1242 1427 1243
rect 1423 1237 1427 1238
rect 1463 1242 1467 1243
rect 1463 1237 1467 1238
rect 1479 1242 1483 1243
rect 1479 1237 1483 1238
rect 1503 1242 1507 1243
rect 1503 1237 1507 1238
rect 1543 1242 1547 1243
rect 1543 1237 1547 1238
rect 1583 1242 1587 1243
rect 1583 1237 1587 1238
rect 1623 1242 1627 1243
rect 1623 1237 1627 1238
rect 1679 1242 1683 1243
rect 1679 1237 1683 1238
rect 1687 1242 1691 1243
rect 1687 1237 1691 1238
rect 1735 1242 1739 1243
rect 1735 1237 1739 1238
rect 1791 1242 1795 1243
rect 1791 1237 1795 1238
rect 1847 1242 1851 1243
rect 1847 1237 1851 1238
rect 1887 1242 1891 1243
rect 1887 1237 1891 1238
rect 1903 1242 1907 1243
rect 1903 1237 1907 1238
rect 1967 1242 1971 1243
rect 1967 1237 1971 1238
rect 1983 1242 1987 1243
rect 1983 1237 1987 1238
rect 2039 1242 2043 1243
rect 2039 1237 2043 1238
rect 2071 1242 2075 1243
rect 2071 1237 2075 1238
rect 2119 1242 2123 1243
rect 2119 1237 2123 1238
rect 2151 1242 2155 1243
rect 2151 1237 2155 1238
rect 2199 1242 2203 1243
rect 2199 1237 2203 1238
rect 2223 1242 2227 1243
rect 2223 1237 2227 1238
rect 2287 1242 2291 1243
rect 2287 1237 2291 1238
rect 2303 1242 2307 1243
rect 2303 1237 2307 1238
rect 2359 1242 2363 1243
rect 2359 1237 2363 1238
rect 2407 1242 2411 1243
rect 2407 1237 2411 1238
rect 112 1230 114 1237
rect 134 1236 140 1237
rect 134 1232 135 1236
rect 139 1232 140 1236
rect 134 1231 140 1232
rect 174 1236 180 1237
rect 174 1232 175 1236
rect 179 1232 180 1236
rect 174 1231 180 1232
rect 230 1236 236 1237
rect 230 1232 231 1236
rect 235 1232 236 1236
rect 230 1231 236 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 398 1236 404 1237
rect 398 1232 399 1236
rect 403 1232 404 1236
rect 398 1231 404 1232
rect 486 1236 492 1237
rect 486 1232 487 1236
rect 491 1232 492 1236
rect 486 1231 492 1232
rect 574 1236 580 1237
rect 574 1232 575 1236
rect 579 1232 580 1236
rect 574 1231 580 1232
rect 662 1236 668 1237
rect 662 1232 663 1236
rect 667 1232 668 1236
rect 662 1231 668 1232
rect 742 1236 748 1237
rect 742 1232 743 1236
rect 747 1232 748 1236
rect 742 1231 748 1232
rect 814 1236 820 1237
rect 814 1232 815 1236
rect 819 1232 820 1236
rect 814 1231 820 1232
rect 878 1236 884 1237
rect 878 1232 879 1236
rect 883 1232 884 1236
rect 878 1231 884 1232
rect 942 1236 948 1237
rect 942 1232 943 1236
rect 947 1232 948 1236
rect 942 1231 948 1232
rect 1006 1236 1012 1237
rect 1006 1232 1007 1236
rect 1011 1232 1012 1236
rect 1006 1231 1012 1232
rect 1070 1236 1076 1237
rect 1070 1232 1071 1236
rect 1075 1232 1076 1236
rect 1070 1231 1076 1232
rect 1240 1230 1242 1237
rect 1280 1230 1282 1237
rect 1302 1236 1308 1237
rect 1302 1232 1303 1236
rect 1307 1232 1308 1236
rect 1302 1231 1308 1232
rect 1374 1236 1380 1237
rect 1374 1232 1375 1236
rect 1379 1232 1380 1236
rect 1374 1231 1380 1232
rect 1478 1236 1484 1237
rect 1478 1232 1479 1236
rect 1483 1232 1484 1236
rect 1478 1231 1484 1232
rect 1582 1236 1588 1237
rect 1582 1232 1583 1236
rect 1587 1232 1588 1236
rect 1582 1231 1588 1232
rect 1686 1236 1692 1237
rect 1686 1232 1687 1236
rect 1691 1232 1692 1236
rect 1686 1231 1692 1232
rect 1790 1236 1796 1237
rect 1790 1232 1791 1236
rect 1795 1232 1796 1236
rect 1790 1231 1796 1232
rect 1886 1236 1892 1237
rect 1886 1232 1887 1236
rect 1891 1232 1892 1236
rect 1886 1231 1892 1232
rect 1982 1236 1988 1237
rect 1982 1232 1983 1236
rect 1987 1232 1988 1236
rect 1982 1231 1988 1232
rect 2070 1236 2076 1237
rect 2070 1232 2071 1236
rect 2075 1232 2076 1236
rect 2070 1231 2076 1232
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2222 1236 2228 1237
rect 2222 1232 2223 1236
rect 2227 1232 2228 1236
rect 2222 1231 2228 1232
rect 2302 1236 2308 1237
rect 2302 1232 2303 1236
rect 2307 1232 2308 1236
rect 2302 1231 2308 1232
rect 2358 1236 2364 1237
rect 2358 1232 2359 1236
rect 2363 1232 2364 1236
rect 2358 1231 2364 1232
rect 2408 1230 2410 1237
rect 110 1229 116 1230
rect 110 1225 111 1229
rect 115 1225 116 1229
rect 110 1224 116 1225
rect 1238 1229 1244 1230
rect 1238 1225 1239 1229
rect 1243 1225 1244 1229
rect 1238 1224 1244 1225
rect 1278 1229 1284 1230
rect 1278 1225 1279 1229
rect 1283 1225 1284 1229
rect 1278 1224 1284 1225
rect 2406 1229 2412 1230
rect 2406 1225 2407 1229
rect 2411 1225 2412 1229
rect 2406 1224 2412 1225
rect 110 1212 116 1213
rect 110 1208 111 1212
rect 115 1208 116 1212
rect 110 1207 116 1208
rect 1238 1212 1244 1213
rect 1238 1208 1239 1212
rect 1243 1208 1244 1212
rect 1238 1207 1244 1208
rect 1278 1212 1284 1213
rect 1278 1208 1279 1212
rect 1283 1208 1284 1212
rect 1278 1207 1284 1208
rect 2406 1212 2412 1213
rect 2406 1208 2407 1212
rect 2411 1208 2412 1212
rect 2406 1207 2412 1208
rect 112 1175 114 1207
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 174 1189 180 1190
rect 174 1185 175 1189
rect 179 1185 180 1189
rect 174 1184 180 1185
rect 230 1189 236 1190
rect 230 1185 231 1189
rect 235 1185 236 1189
rect 230 1184 236 1185
rect 310 1189 316 1190
rect 310 1185 311 1189
rect 315 1185 316 1189
rect 310 1184 316 1185
rect 398 1189 404 1190
rect 398 1185 399 1189
rect 403 1185 404 1189
rect 398 1184 404 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 574 1189 580 1190
rect 574 1185 575 1189
rect 579 1185 580 1189
rect 574 1184 580 1185
rect 662 1189 668 1190
rect 662 1185 663 1189
rect 667 1185 668 1189
rect 662 1184 668 1185
rect 742 1189 748 1190
rect 742 1185 743 1189
rect 747 1185 748 1189
rect 742 1184 748 1185
rect 814 1189 820 1190
rect 814 1185 815 1189
rect 819 1185 820 1189
rect 814 1184 820 1185
rect 878 1189 884 1190
rect 878 1185 879 1189
rect 883 1185 884 1189
rect 878 1184 884 1185
rect 942 1189 948 1190
rect 942 1185 943 1189
rect 947 1185 948 1189
rect 942 1184 948 1185
rect 1006 1189 1012 1190
rect 1006 1185 1007 1189
rect 1011 1185 1012 1189
rect 1006 1184 1012 1185
rect 1070 1189 1076 1190
rect 1070 1185 1071 1189
rect 1075 1185 1076 1189
rect 1070 1184 1076 1185
rect 136 1175 138 1184
rect 176 1175 178 1184
rect 232 1175 234 1184
rect 312 1175 314 1184
rect 400 1175 402 1184
rect 488 1175 490 1184
rect 576 1175 578 1184
rect 664 1175 666 1184
rect 744 1175 746 1184
rect 816 1175 818 1184
rect 880 1175 882 1184
rect 944 1175 946 1184
rect 1008 1175 1010 1184
rect 1072 1175 1074 1184
rect 1240 1175 1242 1207
rect 1280 1175 1282 1207
rect 1302 1189 1308 1190
rect 1302 1185 1303 1189
rect 1307 1185 1308 1189
rect 1302 1184 1308 1185
rect 1374 1189 1380 1190
rect 1374 1185 1375 1189
rect 1379 1185 1380 1189
rect 1374 1184 1380 1185
rect 1478 1189 1484 1190
rect 1478 1185 1479 1189
rect 1483 1185 1484 1189
rect 1478 1184 1484 1185
rect 1582 1189 1588 1190
rect 1582 1185 1583 1189
rect 1587 1185 1588 1189
rect 1582 1184 1588 1185
rect 1686 1189 1692 1190
rect 1686 1185 1687 1189
rect 1691 1185 1692 1189
rect 1686 1184 1692 1185
rect 1790 1189 1796 1190
rect 1790 1185 1791 1189
rect 1795 1185 1796 1189
rect 1790 1184 1796 1185
rect 1886 1189 1892 1190
rect 1886 1185 1887 1189
rect 1891 1185 1892 1189
rect 1886 1184 1892 1185
rect 1982 1189 1988 1190
rect 1982 1185 1983 1189
rect 1987 1185 1988 1189
rect 1982 1184 1988 1185
rect 2070 1189 2076 1190
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 2150 1189 2156 1190
rect 2150 1185 2151 1189
rect 2155 1185 2156 1189
rect 2150 1184 2156 1185
rect 2222 1189 2228 1190
rect 2222 1185 2223 1189
rect 2227 1185 2228 1189
rect 2222 1184 2228 1185
rect 2302 1189 2308 1190
rect 2302 1185 2303 1189
rect 2307 1185 2308 1189
rect 2302 1184 2308 1185
rect 2358 1189 2364 1190
rect 2358 1185 2359 1189
rect 2363 1185 2364 1189
rect 2358 1184 2364 1185
rect 1304 1175 1306 1184
rect 1376 1175 1378 1184
rect 1480 1175 1482 1184
rect 1584 1175 1586 1184
rect 1688 1175 1690 1184
rect 1792 1175 1794 1184
rect 1888 1175 1890 1184
rect 1984 1175 1986 1184
rect 2072 1175 2074 1184
rect 2152 1175 2154 1184
rect 2224 1175 2226 1184
rect 2304 1175 2306 1184
rect 2360 1175 2362 1184
rect 2408 1175 2410 1207
rect 111 1174 115 1175
rect 111 1169 115 1170
rect 135 1174 139 1175
rect 135 1169 139 1170
rect 175 1174 179 1175
rect 175 1169 179 1170
rect 231 1174 235 1175
rect 231 1169 235 1170
rect 239 1174 243 1175
rect 239 1169 243 1170
rect 311 1174 315 1175
rect 311 1169 315 1170
rect 327 1174 331 1175
rect 327 1169 331 1170
rect 399 1174 403 1175
rect 399 1169 403 1170
rect 431 1174 435 1175
rect 431 1169 435 1170
rect 487 1174 491 1175
rect 487 1169 491 1170
rect 535 1174 539 1175
rect 535 1169 539 1170
rect 575 1174 579 1175
rect 575 1169 579 1170
rect 639 1174 643 1175
rect 639 1169 643 1170
rect 663 1174 667 1175
rect 663 1169 667 1170
rect 743 1174 747 1175
rect 743 1169 747 1170
rect 815 1174 819 1175
rect 815 1169 819 1170
rect 839 1174 843 1175
rect 839 1169 843 1170
rect 879 1174 883 1175
rect 879 1169 883 1170
rect 919 1174 923 1175
rect 919 1169 923 1170
rect 943 1174 947 1175
rect 943 1169 947 1170
rect 999 1174 1003 1175
rect 999 1169 1003 1170
rect 1007 1174 1011 1175
rect 1007 1169 1011 1170
rect 1071 1174 1075 1175
rect 1071 1169 1075 1170
rect 1143 1174 1147 1175
rect 1143 1169 1147 1170
rect 1191 1174 1195 1175
rect 1191 1169 1195 1170
rect 1239 1174 1243 1175
rect 1239 1169 1243 1170
rect 1279 1174 1283 1175
rect 1279 1169 1283 1170
rect 1303 1174 1307 1175
rect 1303 1169 1307 1170
rect 1343 1174 1347 1175
rect 1343 1169 1347 1170
rect 1375 1174 1379 1175
rect 1375 1169 1379 1170
rect 1407 1174 1411 1175
rect 1407 1169 1411 1170
rect 1479 1174 1483 1175
rect 1479 1169 1483 1170
rect 1487 1174 1491 1175
rect 1487 1169 1491 1170
rect 1583 1174 1587 1175
rect 1583 1169 1587 1170
rect 1687 1174 1691 1175
rect 1687 1169 1691 1170
rect 1791 1174 1795 1175
rect 1791 1169 1795 1170
rect 1799 1174 1803 1175
rect 1799 1169 1803 1170
rect 1887 1174 1891 1175
rect 1887 1169 1891 1170
rect 1903 1174 1907 1175
rect 1903 1169 1907 1170
rect 1983 1174 1987 1175
rect 1983 1169 1987 1170
rect 1999 1174 2003 1175
rect 1999 1169 2003 1170
rect 2071 1174 2075 1175
rect 2071 1169 2075 1170
rect 2079 1174 2083 1175
rect 2079 1169 2083 1170
rect 2151 1174 2155 1175
rect 2151 1169 2155 1170
rect 2159 1174 2163 1175
rect 2159 1169 2163 1170
rect 2223 1174 2227 1175
rect 2223 1169 2227 1170
rect 2231 1174 2235 1175
rect 2231 1169 2235 1170
rect 2303 1174 2307 1175
rect 2303 1169 2307 1170
rect 2359 1174 2363 1175
rect 2359 1169 2363 1170
rect 2407 1174 2411 1175
rect 2407 1169 2411 1170
rect 112 1137 114 1169
rect 136 1160 138 1169
rect 176 1160 178 1169
rect 240 1160 242 1169
rect 328 1160 330 1169
rect 432 1160 434 1169
rect 536 1160 538 1169
rect 640 1160 642 1169
rect 744 1160 746 1169
rect 840 1160 842 1169
rect 920 1160 922 1169
rect 1000 1160 1002 1169
rect 1072 1160 1074 1169
rect 1144 1160 1146 1169
rect 1192 1160 1194 1169
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1155 140 1159
rect 134 1154 140 1155
rect 174 1159 180 1160
rect 174 1155 175 1159
rect 179 1155 180 1159
rect 174 1154 180 1155
rect 238 1159 244 1160
rect 238 1155 239 1159
rect 243 1155 244 1159
rect 238 1154 244 1155
rect 326 1159 332 1160
rect 326 1155 327 1159
rect 331 1155 332 1159
rect 326 1154 332 1155
rect 430 1159 436 1160
rect 430 1155 431 1159
rect 435 1155 436 1159
rect 430 1154 436 1155
rect 534 1159 540 1160
rect 534 1155 535 1159
rect 539 1155 540 1159
rect 534 1154 540 1155
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1155 644 1159
rect 638 1154 644 1155
rect 742 1159 748 1160
rect 742 1155 743 1159
rect 747 1155 748 1159
rect 742 1154 748 1155
rect 838 1159 844 1160
rect 838 1155 839 1159
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 918 1159 924 1160
rect 918 1155 919 1159
rect 923 1155 924 1159
rect 918 1154 924 1155
rect 998 1159 1004 1160
rect 998 1155 999 1159
rect 1003 1155 1004 1159
rect 998 1154 1004 1155
rect 1070 1159 1076 1160
rect 1070 1155 1071 1159
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 1142 1159 1148 1160
rect 1142 1155 1143 1159
rect 1147 1155 1148 1159
rect 1142 1154 1148 1155
rect 1190 1159 1196 1160
rect 1190 1155 1191 1159
rect 1195 1155 1196 1159
rect 1190 1154 1196 1155
rect 1240 1137 1242 1169
rect 1280 1137 1282 1169
rect 1304 1160 1306 1169
rect 1344 1160 1346 1169
rect 1408 1160 1410 1169
rect 1488 1160 1490 1169
rect 1584 1160 1586 1169
rect 1688 1160 1690 1169
rect 1800 1160 1802 1169
rect 1904 1160 1906 1169
rect 2000 1160 2002 1169
rect 2080 1160 2082 1169
rect 2160 1160 2162 1169
rect 2232 1160 2234 1169
rect 2304 1160 2306 1169
rect 2360 1160 2362 1169
rect 1302 1159 1308 1160
rect 1302 1155 1303 1159
rect 1307 1155 1308 1159
rect 1302 1154 1308 1155
rect 1342 1159 1348 1160
rect 1342 1155 1343 1159
rect 1347 1155 1348 1159
rect 1342 1154 1348 1155
rect 1406 1159 1412 1160
rect 1406 1155 1407 1159
rect 1411 1155 1412 1159
rect 1406 1154 1412 1155
rect 1486 1159 1492 1160
rect 1486 1155 1487 1159
rect 1491 1155 1492 1159
rect 1486 1154 1492 1155
rect 1582 1159 1588 1160
rect 1582 1155 1583 1159
rect 1587 1155 1588 1159
rect 1582 1154 1588 1155
rect 1686 1159 1692 1160
rect 1686 1155 1687 1159
rect 1691 1155 1692 1159
rect 1686 1154 1692 1155
rect 1798 1159 1804 1160
rect 1798 1155 1799 1159
rect 1803 1155 1804 1159
rect 1798 1154 1804 1155
rect 1902 1159 1908 1160
rect 1902 1155 1903 1159
rect 1907 1155 1908 1159
rect 1902 1154 1908 1155
rect 1998 1159 2004 1160
rect 1998 1155 1999 1159
rect 2003 1155 2004 1159
rect 1998 1154 2004 1155
rect 2078 1159 2084 1160
rect 2078 1155 2079 1159
rect 2083 1155 2084 1159
rect 2078 1154 2084 1155
rect 2158 1159 2164 1160
rect 2158 1155 2159 1159
rect 2163 1155 2164 1159
rect 2158 1154 2164 1155
rect 2230 1159 2236 1160
rect 2230 1155 2231 1159
rect 2235 1155 2236 1159
rect 2230 1154 2236 1155
rect 2302 1159 2308 1160
rect 2302 1155 2303 1159
rect 2307 1155 2308 1159
rect 2302 1154 2308 1155
rect 2358 1159 2364 1160
rect 2358 1155 2359 1159
rect 2363 1155 2364 1159
rect 2358 1154 2364 1155
rect 2408 1137 2410 1169
rect 110 1136 116 1137
rect 110 1132 111 1136
rect 115 1132 116 1136
rect 110 1131 116 1132
rect 1238 1136 1244 1137
rect 1238 1132 1239 1136
rect 1243 1132 1244 1136
rect 1238 1131 1244 1132
rect 1278 1136 1284 1137
rect 1278 1132 1279 1136
rect 1283 1132 1284 1136
rect 1278 1131 1284 1132
rect 2406 1136 2412 1137
rect 2406 1132 2407 1136
rect 2411 1132 2412 1136
rect 2406 1131 2412 1132
rect 110 1119 116 1120
rect 110 1115 111 1119
rect 115 1115 116 1119
rect 110 1114 116 1115
rect 1238 1119 1244 1120
rect 1238 1115 1239 1119
rect 1243 1115 1244 1119
rect 1238 1114 1244 1115
rect 1278 1119 1284 1120
rect 1278 1115 1279 1119
rect 1283 1115 1284 1119
rect 1278 1114 1284 1115
rect 2406 1119 2412 1120
rect 2406 1115 2407 1119
rect 2411 1115 2412 1119
rect 2406 1114 2412 1115
rect 112 1103 114 1114
rect 134 1112 140 1113
rect 134 1108 135 1112
rect 139 1108 140 1112
rect 134 1107 140 1108
rect 174 1112 180 1113
rect 174 1108 175 1112
rect 179 1108 180 1112
rect 174 1107 180 1108
rect 238 1112 244 1113
rect 238 1108 239 1112
rect 243 1108 244 1112
rect 238 1107 244 1108
rect 326 1112 332 1113
rect 326 1108 327 1112
rect 331 1108 332 1112
rect 326 1107 332 1108
rect 430 1112 436 1113
rect 430 1108 431 1112
rect 435 1108 436 1112
rect 430 1107 436 1108
rect 534 1112 540 1113
rect 534 1108 535 1112
rect 539 1108 540 1112
rect 534 1107 540 1108
rect 638 1112 644 1113
rect 638 1108 639 1112
rect 643 1108 644 1112
rect 638 1107 644 1108
rect 742 1112 748 1113
rect 742 1108 743 1112
rect 747 1108 748 1112
rect 742 1107 748 1108
rect 838 1112 844 1113
rect 838 1108 839 1112
rect 843 1108 844 1112
rect 838 1107 844 1108
rect 918 1112 924 1113
rect 918 1108 919 1112
rect 923 1108 924 1112
rect 918 1107 924 1108
rect 998 1112 1004 1113
rect 998 1108 999 1112
rect 1003 1108 1004 1112
rect 998 1107 1004 1108
rect 1070 1112 1076 1113
rect 1070 1108 1071 1112
rect 1075 1108 1076 1112
rect 1070 1107 1076 1108
rect 1142 1112 1148 1113
rect 1142 1108 1143 1112
rect 1147 1108 1148 1112
rect 1142 1107 1148 1108
rect 1190 1112 1196 1113
rect 1190 1108 1191 1112
rect 1195 1108 1196 1112
rect 1190 1107 1196 1108
rect 136 1103 138 1107
rect 176 1103 178 1107
rect 240 1103 242 1107
rect 328 1103 330 1107
rect 432 1103 434 1107
rect 536 1103 538 1107
rect 640 1103 642 1107
rect 744 1103 746 1107
rect 840 1103 842 1107
rect 920 1103 922 1107
rect 1000 1103 1002 1107
rect 1072 1103 1074 1107
rect 1144 1103 1146 1107
rect 1192 1103 1194 1107
rect 1240 1103 1242 1114
rect 1280 1107 1282 1114
rect 1302 1112 1308 1113
rect 1302 1108 1303 1112
rect 1307 1108 1308 1112
rect 1302 1107 1308 1108
rect 1342 1112 1348 1113
rect 1342 1108 1343 1112
rect 1347 1108 1348 1112
rect 1342 1107 1348 1108
rect 1406 1112 1412 1113
rect 1406 1108 1407 1112
rect 1411 1108 1412 1112
rect 1406 1107 1412 1108
rect 1486 1112 1492 1113
rect 1486 1108 1487 1112
rect 1491 1108 1492 1112
rect 1486 1107 1492 1108
rect 1582 1112 1588 1113
rect 1582 1108 1583 1112
rect 1587 1108 1588 1112
rect 1582 1107 1588 1108
rect 1686 1112 1692 1113
rect 1686 1108 1687 1112
rect 1691 1108 1692 1112
rect 1686 1107 1692 1108
rect 1798 1112 1804 1113
rect 1798 1108 1799 1112
rect 1803 1108 1804 1112
rect 1798 1107 1804 1108
rect 1902 1112 1908 1113
rect 1902 1108 1903 1112
rect 1907 1108 1908 1112
rect 1902 1107 1908 1108
rect 1998 1112 2004 1113
rect 1998 1108 1999 1112
rect 2003 1108 2004 1112
rect 1998 1107 2004 1108
rect 2078 1112 2084 1113
rect 2078 1108 2079 1112
rect 2083 1108 2084 1112
rect 2078 1107 2084 1108
rect 2158 1112 2164 1113
rect 2158 1108 2159 1112
rect 2163 1108 2164 1112
rect 2158 1107 2164 1108
rect 2230 1112 2236 1113
rect 2230 1108 2231 1112
rect 2235 1108 2236 1112
rect 2230 1107 2236 1108
rect 2302 1112 2308 1113
rect 2302 1108 2303 1112
rect 2307 1108 2308 1112
rect 2302 1107 2308 1108
rect 2358 1112 2364 1113
rect 2358 1108 2359 1112
rect 2363 1108 2364 1112
rect 2358 1107 2364 1108
rect 2408 1107 2410 1114
rect 1279 1106 1283 1107
rect 111 1102 115 1103
rect 111 1097 115 1098
rect 135 1102 139 1103
rect 135 1097 139 1098
rect 175 1102 179 1103
rect 175 1097 179 1098
rect 239 1102 243 1103
rect 239 1097 243 1098
rect 247 1102 251 1103
rect 247 1097 251 1098
rect 327 1102 331 1103
rect 327 1097 331 1098
rect 415 1102 419 1103
rect 415 1097 419 1098
rect 431 1102 435 1103
rect 431 1097 435 1098
rect 503 1102 507 1103
rect 503 1097 507 1098
rect 535 1102 539 1103
rect 535 1097 539 1098
rect 583 1102 587 1103
rect 583 1097 587 1098
rect 639 1102 643 1103
rect 639 1097 643 1098
rect 663 1102 667 1103
rect 663 1097 667 1098
rect 735 1102 739 1103
rect 735 1097 739 1098
rect 743 1102 747 1103
rect 743 1097 747 1098
rect 799 1102 803 1103
rect 799 1097 803 1098
rect 839 1102 843 1103
rect 839 1097 843 1098
rect 863 1102 867 1103
rect 863 1097 867 1098
rect 919 1102 923 1103
rect 919 1097 923 1098
rect 983 1102 987 1103
rect 983 1097 987 1098
rect 999 1102 1003 1103
rect 999 1097 1003 1098
rect 1047 1102 1051 1103
rect 1047 1097 1051 1098
rect 1071 1102 1075 1103
rect 1071 1097 1075 1098
rect 1143 1102 1147 1103
rect 1143 1097 1147 1098
rect 1191 1102 1195 1103
rect 1191 1097 1195 1098
rect 1239 1102 1243 1103
rect 1279 1101 1283 1102
rect 1303 1106 1307 1107
rect 1303 1101 1307 1102
rect 1343 1106 1347 1107
rect 1343 1101 1347 1102
rect 1407 1106 1411 1107
rect 1407 1101 1411 1102
rect 1431 1106 1435 1107
rect 1431 1101 1435 1102
rect 1471 1106 1475 1107
rect 1471 1101 1475 1102
rect 1487 1106 1491 1107
rect 1487 1101 1491 1102
rect 1511 1106 1515 1107
rect 1511 1101 1515 1102
rect 1559 1106 1563 1107
rect 1559 1101 1563 1102
rect 1583 1106 1587 1107
rect 1583 1101 1587 1102
rect 1615 1106 1619 1107
rect 1615 1101 1619 1102
rect 1671 1106 1675 1107
rect 1671 1101 1675 1102
rect 1687 1106 1691 1107
rect 1687 1101 1691 1102
rect 1727 1106 1731 1107
rect 1727 1101 1731 1102
rect 1775 1106 1779 1107
rect 1775 1101 1779 1102
rect 1799 1106 1803 1107
rect 1799 1101 1803 1102
rect 1823 1106 1827 1107
rect 1823 1101 1827 1102
rect 1871 1106 1875 1107
rect 1871 1101 1875 1102
rect 1903 1106 1907 1107
rect 1903 1101 1907 1102
rect 1919 1106 1923 1107
rect 1919 1101 1923 1102
rect 1967 1106 1971 1107
rect 1967 1101 1971 1102
rect 1999 1106 2003 1107
rect 1999 1101 2003 1102
rect 2015 1106 2019 1107
rect 2015 1101 2019 1102
rect 2063 1106 2067 1107
rect 2063 1101 2067 1102
rect 2079 1106 2083 1107
rect 2079 1101 2083 1102
rect 2119 1106 2123 1107
rect 2119 1101 2123 1102
rect 2159 1106 2163 1107
rect 2159 1101 2163 1102
rect 2175 1106 2179 1107
rect 2175 1101 2179 1102
rect 2231 1106 2235 1107
rect 2231 1101 2235 1102
rect 2303 1106 2307 1107
rect 2303 1101 2307 1102
rect 2359 1106 2363 1107
rect 2359 1101 2363 1102
rect 2407 1106 2411 1107
rect 2407 1101 2411 1102
rect 1239 1097 1243 1098
rect 112 1090 114 1097
rect 134 1096 140 1097
rect 134 1092 135 1096
rect 139 1092 140 1096
rect 134 1091 140 1092
rect 174 1096 180 1097
rect 174 1092 175 1096
rect 179 1092 180 1096
rect 174 1091 180 1092
rect 246 1096 252 1097
rect 246 1092 247 1096
rect 251 1092 252 1096
rect 246 1091 252 1092
rect 326 1096 332 1097
rect 326 1092 327 1096
rect 331 1092 332 1096
rect 326 1091 332 1092
rect 414 1096 420 1097
rect 414 1092 415 1096
rect 419 1092 420 1096
rect 414 1091 420 1092
rect 502 1096 508 1097
rect 502 1092 503 1096
rect 507 1092 508 1096
rect 502 1091 508 1092
rect 582 1096 588 1097
rect 582 1092 583 1096
rect 587 1092 588 1096
rect 582 1091 588 1092
rect 662 1096 668 1097
rect 662 1092 663 1096
rect 667 1092 668 1096
rect 662 1091 668 1092
rect 734 1096 740 1097
rect 734 1092 735 1096
rect 739 1092 740 1096
rect 734 1091 740 1092
rect 798 1096 804 1097
rect 798 1092 799 1096
rect 803 1092 804 1096
rect 798 1091 804 1092
rect 862 1096 868 1097
rect 862 1092 863 1096
rect 867 1092 868 1096
rect 862 1091 868 1092
rect 918 1096 924 1097
rect 918 1092 919 1096
rect 923 1092 924 1096
rect 918 1091 924 1092
rect 982 1096 988 1097
rect 982 1092 983 1096
rect 987 1092 988 1096
rect 982 1091 988 1092
rect 1046 1096 1052 1097
rect 1046 1092 1047 1096
rect 1051 1092 1052 1096
rect 1046 1091 1052 1092
rect 1240 1090 1242 1097
rect 1280 1094 1282 1101
rect 1430 1100 1436 1101
rect 1430 1096 1431 1100
rect 1435 1096 1436 1100
rect 1430 1095 1436 1096
rect 1470 1100 1476 1101
rect 1470 1096 1471 1100
rect 1475 1096 1476 1100
rect 1470 1095 1476 1096
rect 1510 1100 1516 1101
rect 1510 1096 1511 1100
rect 1515 1096 1516 1100
rect 1510 1095 1516 1096
rect 1558 1100 1564 1101
rect 1558 1096 1559 1100
rect 1563 1096 1564 1100
rect 1558 1095 1564 1096
rect 1614 1100 1620 1101
rect 1614 1096 1615 1100
rect 1619 1096 1620 1100
rect 1614 1095 1620 1096
rect 1670 1100 1676 1101
rect 1670 1096 1671 1100
rect 1675 1096 1676 1100
rect 1670 1095 1676 1096
rect 1726 1100 1732 1101
rect 1726 1096 1727 1100
rect 1731 1096 1732 1100
rect 1726 1095 1732 1096
rect 1774 1100 1780 1101
rect 1774 1096 1775 1100
rect 1779 1096 1780 1100
rect 1774 1095 1780 1096
rect 1822 1100 1828 1101
rect 1822 1096 1823 1100
rect 1827 1096 1828 1100
rect 1822 1095 1828 1096
rect 1870 1100 1876 1101
rect 1870 1096 1871 1100
rect 1875 1096 1876 1100
rect 1870 1095 1876 1096
rect 1918 1100 1924 1101
rect 1918 1096 1919 1100
rect 1923 1096 1924 1100
rect 1918 1095 1924 1096
rect 1966 1100 1972 1101
rect 1966 1096 1967 1100
rect 1971 1096 1972 1100
rect 1966 1095 1972 1096
rect 2014 1100 2020 1101
rect 2014 1096 2015 1100
rect 2019 1096 2020 1100
rect 2014 1095 2020 1096
rect 2062 1100 2068 1101
rect 2062 1096 2063 1100
rect 2067 1096 2068 1100
rect 2062 1095 2068 1096
rect 2118 1100 2124 1101
rect 2118 1096 2119 1100
rect 2123 1096 2124 1100
rect 2118 1095 2124 1096
rect 2174 1100 2180 1101
rect 2174 1096 2175 1100
rect 2179 1096 2180 1100
rect 2174 1095 2180 1096
rect 2230 1100 2236 1101
rect 2230 1096 2231 1100
rect 2235 1096 2236 1100
rect 2230 1095 2236 1096
rect 2408 1094 2410 1101
rect 1278 1093 1284 1094
rect 110 1089 116 1090
rect 110 1085 111 1089
rect 115 1085 116 1089
rect 110 1084 116 1085
rect 1238 1089 1244 1090
rect 1238 1085 1239 1089
rect 1243 1085 1244 1089
rect 1278 1089 1279 1093
rect 1283 1089 1284 1093
rect 1278 1088 1284 1089
rect 2406 1093 2412 1094
rect 2406 1089 2407 1093
rect 2411 1089 2412 1093
rect 2406 1088 2412 1089
rect 1238 1084 1244 1085
rect 1278 1076 1284 1077
rect 110 1072 116 1073
rect 110 1068 111 1072
rect 115 1068 116 1072
rect 110 1067 116 1068
rect 1238 1072 1244 1073
rect 1238 1068 1239 1072
rect 1243 1068 1244 1072
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 2406 1076 2412 1077
rect 2406 1072 2407 1076
rect 2411 1072 2412 1076
rect 2406 1071 2412 1072
rect 1238 1067 1244 1068
rect 112 1035 114 1067
rect 134 1049 140 1050
rect 134 1045 135 1049
rect 139 1045 140 1049
rect 134 1044 140 1045
rect 174 1049 180 1050
rect 174 1045 175 1049
rect 179 1045 180 1049
rect 174 1044 180 1045
rect 246 1049 252 1050
rect 246 1045 247 1049
rect 251 1045 252 1049
rect 246 1044 252 1045
rect 326 1049 332 1050
rect 326 1045 327 1049
rect 331 1045 332 1049
rect 326 1044 332 1045
rect 414 1049 420 1050
rect 414 1045 415 1049
rect 419 1045 420 1049
rect 414 1044 420 1045
rect 502 1049 508 1050
rect 502 1045 503 1049
rect 507 1045 508 1049
rect 502 1044 508 1045
rect 582 1049 588 1050
rect 582 1045 583 1049
rect 587 1045 588 1049
rect 582 1044 588 1045
rect 662 1049 668 1050
rect 662 1045 663 1049
rect 667 1045 668 1049
rect 662 1044 668 1045
rect 734 1049 740 1050
rect 734 1045 735 1049
rect 739 1045 740 1049
rect 734 1044 740 1045
rect 798 1049 804 1050
rect 798 1045 799 1049
rect 803 1045 804 1049
rect 798 1044 804 1045
rect 862 1049 868 1050
rect 862 1045 863 1049
rect 867 1045 868 1049
rect 862 1044 868 1045
rect 918 1049 924 1050
rect 918 1045 919 1049
rect 923 1045 924 1049
rect 918 1044 924 1045
rect 982 1049 988 1050
rect 982 1045 983 1049
rect 987 1045 988 1049
rect 982 1044 988 1045
rect 1046 1049 1052 1050
rect 1046 1045 1047 1049
rect 1051 1045 1052 1049
rect 1046 1044 1052 1045
rect 136 1035 138 1044
rect 176 1035 178 1044
rect 248 1035 250 1044
rect 328 1035 330 1044
rect 416 1035 418 1044
rect 504 1035 506 1044
rect 584 1035 586 1044
rect 664 1035 666 1044
rect 736 1035 738 1044
rect 800 1035 802 1044
rect 864 1035 866 1044
rect 920 1035 922 1044
rect 984 1035 986 1044
rect 1048 1035 1050 1044
rect 1240 1035 1242 1067
rect 1280 1039 1282 1071
rect 1430 1053 1436 1054
rect 1430 1049 1431 1053
rect 1435 1049 1436 1053
rect 1430 1048 1436 1049
rect 1470 1053 1476 1054
rect 1470 1049 1471 1053
rect 1475 1049 1476 1053
rect 1470 1048 1476 1049
rect 1510 1053 1516 1054
rect 1510 1049 1511 1053
rect 1515 1049 1516 1053
rect 1510 1048 1516 1049
rect 1558 1053 1564 1054
rect 1558 1049 1559 1053
rect 1563 1049 1564 1053
rect 1558 1048 1564 1049
rect 1614 1053 1620 1054
rect 1614 1049 1615 1053
rect 1619 1049 1620 1053
rect 1614 1048 1620 1049
rect 1670 1053 1676 1054
rect 1670 1049 1671 1053
rect 1675 1049 1676 1053
rect 1670 1048 1676 1049
rect 1726 1053 1732 1054
rect 1726 1049 1727 1053
rect 1731 1049 1732 1053
rect 1726 1048 1732 1049
rect 1774 1053 1780 1054
rect 1774 1049 1775 1053
rect 1779 1049 1780 1053
rect 1774 1048 1780 1049
rect 1822 1053 1828 1054
rect 1822 1049 1823 1053
rect 1827 1049 1828 1053
rect 1822 1048 1828 1049
rect 1870 1053 1876 1054
rect 1870 1049 1871 1053
rect 1875 1049 1876 1053
rect 1870 1048 1876 1049
rect 1918 1053 1924 1054
rect 1918 1049 1919 1053
rect 1923 1049 1924 1053
rect 1918 1048 1924 1049
rect 1966 1053 1972 1054
rect 1966 1049 1967 1053
rect 1971 1049 1972 1053
rect 1966 1048 1972 1049
rect 2014 1053 2020 1054
rect 2014 1049 2015 1053
rect 2019 1049 2020 1053
rect 2014 1048 2020 1049
rect 2062 1053 2068 1054
rect 2062 1049 2063 1053
rect 2067 1049 2068 1053
rect 2062 1048 2068 1049
rect 2118 1053 2124 1054
rect 2118 1049 2119 1053
rect 2123 1049 2124 1053
rect 2118 1048 2124 1049
rect 2174 1053 2180 1054
rect 2174 1049 2175 1053
rect 2179 1049 2180 1053
rect 2174 1048 2180 1049
rect 2230 1053 2236 1054
rect 2230 1049 2231 1053
rect 2235 1049 2236 1053
rect 2230 1048 2236 1049
rect 1432 1039 1434 1048
rect 1472 1039 1474 1048
rect 1512 1039 1514 1048
rect 1560 1039 1562 1048
rect 1616 1039 1618 1048
rect 1672 1039 1674 1048
rect 1728 1039 1730 1048
rect 1776 1039 1778 1048
rect 1824 1039 1826 1048
rect 1872 1039 1874 1048
rect 1920 1039 1922 1048
rect 1968 1039 1970 1048
rect 2016 1039 2018 1048
rect 2064 1039 2066 1048
rect 2120 1039 2122 1048
rect 2176 1039 2178 1048
rect 2232 1039 2234 1048
rect 2408 1039 2410 1071
rect 1279 1038 1283 1039
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 135 1034 139 1035
rect 135 1029 139 1030
rect 175 1034 179 1035
rect 175 1029 179 1030
rect 247 1034 251 1035
rect 247 1029 251 1030
rect 255 1034 259 1035
rect 255 1029 259 1030
rect 327 1034 331 1035
rect 327 1029 331 1030
rect 399 1034 403 1035
rect 399 1029 403 1030
rect 415 1034 419 1035
rect 415 1029 419 1030
rect 463 1034 467 1035
rect 463 1029 467 1030
rect 503 1034 507 1035
rect 503 1029 507 1030
rect 519 1034 523 1035
rect 519 1029 523 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 583 1034 587 1035
rect 583 1029 587 1030
rect 623 1034 627 1035
rect 623 1029 627 1030
rect 663 1034 667 1035
rect 663 1029 667 1030
rect 671 1034 675 1035
rect 671 1029 675 1030
rect 735 1034 739 1035
rect 735 1029 739 1030
rect 799 1034 803 1035
rect 799 1029 803 1030
rect 807 1034 811 1035
rect 807 1029 811 1030
rect 863 1034 867 1035
rect 863 1029 867 1030
rect 895 1034 899 1035
rect 895 1029 899 1030
rect 919 1034 923 1035
rect 919 1029 923 1030
rect 983 1034 987 1035
rect 983 1029 987 1030
rect 999 1034 1003 1035
rect 999 1029 1003 1030
rect 1047 1034 1051 1035
rect 1047 1029 1051 1030
rect 1103 1034 1107 1035
rect 1103 1029 1107 1030
rect 1191 1034 1195 1035
rect 1191 1029 1195 1030
rect 1239 1034 1243 1035
rect 1279 1033 1283 1034
rect 1431 1038 1435 1039
rect 1431 1033 1435 1034
rect 1471 1038 1475 1039
rect 1471 1033 1475 1034
rect 1511 1038 1515 1039
rect 1511 1033 1515 1034
rect 1559 1038 1563 1039
rect 1559 1033 1563 1034
rect 1575 1038 1579 1039
rect 1575 1033 1579 1034
rect 1615 1038 1619 1039
rect 1615 1033 1619 1034
rect 1655 1038 1659 1039
rect 1655 1033 1659 1034
rect 1671 1038 1675 1039
rect 1671 1033 1675 1034
rect 1695 1038 1699 1039
rect 1695 1033 1699 1034
rect 1727 1038 1731 1039
rect 1727 1033 1731 1034
rect 1735 1038 1739 1039
rect 1735 1033 1739 1034
rect 1775 1038 1779 1039
rect 1775 1033 1779 1034
rect 1823 1038 1827 1039
rect 1823 1033 1827 1034
rect 1871 1038 1875 1039
rect 1871 1033 1875 1034
rect 1879 1038 1883 1039
rect 1879 1033 1883 1034
rect 1919 1038 1923 1039
rect 1919 1033 1923 1034
rect 1943 1038 1947 1039
rect 1943 1033 1947 1034
rect 1967 1038 1971 1039
rect 1967 1033 1971 1034
rect 2015 1038 2019 1039
rect 2015 1033 2019 1034
rect 2063 1038 2067 1039
rect 2063 1033 2067 1034
rect 2095 1038 2099 1039
rect 2095 1033 2099 1034
rect 2119 1038 2123 1039
rect 2119 1033 2123 1034
rect 2175 1038 2179 1039
rect 2175 1033 2179 1034
rect 2231 1038 2235 1039
rect 2231 1033 2235 1034
rect 2255 1038 2259 1039
rect 2255 1033 2259 1034
rect 2407 1038 2411 1039
rect 2407 1033 2411 1034
rect 1239 1029 1243 1030
rect 112 997 114 1029
rect 176 1020 178 1029
rect 256 1020 258 1029
rect 328 1020 330 1029
rect 400 1020 402 1029
rect 464 1020 466 1029
rect 520 1020 522 1029
rect 576 1020 578 1029
rect 624 1020 626 1029
rect 672 1020 674 1029
rect 736 1020 738 1029
rect 808 1020 810 1029
rect 896 1020 898 1029
rect 1000 1020 1002 1029
rect 1104 1020 1106 1029
rect 1192 1020 1194 1029
rect 174 1019 180 1020
rect 174 1015 175 1019
rect 179 1015 180 1019
rect 174 1014 180 1015
rect 254 1019 260 1020
rect 254 1015 255 1019
rect 259 1015 260 1019
rect 254 1014 260 1015
rect 326 1019 332 1020
rect 326 1015 327 1019
rect 331 1015 332 1019
rect 326 1014 332 1015
rect 398 1019 404 1020
rect 398 1015 399 1019
rect 403 1015 404 1019
rect 398 1014 404 1015
rect 462 1019 468 1020
rect 462 1015 463 1019
rect 467 1015 468 1019
rect 462 1014 468 1015
rect 518 1019 524 1020
rect 518 1015 519 1019
rect 523 1015 524 1019
rect 518 1014 524 1015
rect 574 1019 580 1020
rect 574 1015 575 1019
rect 579 1015 580 1019
rect 574 1014 580 1015
rect 622 1019 628 1020
rect 622 1015 623 1019
rect 627 1015 628 1019
rect 622 1014 628 1015
rect 670 1019 676 1020
rect 670 1015 671 1019
rect 675 1015 676 1019
rect 670 1014 676 1015
rect 734 1019 740 1020
rect 734 1015 735 1019
rect 739 1015 740 1019
rect 734 1014 740 1015
rect 806 1019 812 1020
rect 806 1015 807 1019
rect 811 1015 812 1019
rect 806 1014 812 1015
rect 894 1019 900 1020
rect 894 1015 895 1019
rect 899 1015 900 1019
rect 894 1014 900 1015
rect 998 1019 1004 1020
rect 998 1015 999 1019
rect 1003 1015 1004 1019
rect 998 1014 1004 1015
rect 1102 1019 1108 1020
rect 1102 1015 1103 1019
rect 1107 1015 1108 1019
rect 1102 1014 1108 1015
rect 1190 1019 1196 1020
rect 1190 1015 1191 1019
rect 1195 1015 1196 1019
rect 1190 1014 1196 1015
rect 1240 997 1242 1029
rect 1280 1001 1282 1033
rect 1576 1024 1578 1033
rect 1616 1024 1618 1033
rect 1656 1024 1658 1033
rect 1696 1024 1698 1033
rect 1736 1024 1738 1033
rect 1776 1024 1778 1033
rect 1824 1024 1826 1033
rect 1880 1024 1882 1033
rect 1944 1024 1946 1033
rect 2016 1024 2018 1033
rect 2096 1024 2098 1033
rect 2176 1024 2178 1033
rect 2256 1024 2258 1033
rect 1574 1023 1580 1024
rect 1574 1019 1575 1023
rect 1579 1019 1580 1023
rect 1574 1018 1580 1019
rect 1614 1023 1620 1024
rect 1614 1019 1615 1023
rect 1619 1019 1620 1023
rect 1614 1018 1620 1019
rect 1654 1023 1660 1024
rect 1654 1019 1655 1023
rect 1659 1019 1660 1023
rect 1654 1018 1660 1019
rect 1694 1023 1700 1024
rect 1694 1019 1695 1023
rect 1699 1019 1700 1023
rect 1694 1018 1700 1019
rect 1734 1023 1740 1024
rect 1734 1019 1735 1023
rect 1739 1019 1740 1023
rect 1734 1018 1740 1019
rect 1774 1023 1780 1024
rect 1774 1019 1775 1023
rect 1779 1019 1780 1023
rect 1774 1018 1780 1019
rect 1822 1023 1828 1024
rect 1822 1019 1823 1023
rect 1827 1019 1828 1023
rect 1822 1018 1828 1019
rect 1878 1023 1884 1024
rect 1878 1019 1879 1023
rect 1883 1019 1884 1023
rect 1878 1018 1884 1019
rect 1942 1023 1948 1024
rect 1942 1019 1943 1023
rect 1947 1019 1948 1023
rect 1942 1018 1948 1019
rect 2014 1023 2020 1024
rect 2014 1019 2015 1023
rect 2019 1019 2020 1023
rect 2014 1018 2020 1019
rect 2094 1023 2100 1024
rect 2094 1019 2095 1023
rect 2099 1019 2100 1023
rect 2094 1018 2100 1019
rect 2174 1023 2180 1024
rect 2174 1019 2175 1023
rect 2179 1019 2180 1023
rect 2174 1018 2180 1019
rect 2254 1023 2260 1024
rect 2254 1019 2255 1023
rect 2259 1019 2260 1023
rect 2254 1018 2260 1019
rect 2408 1001 2410 1033
rect 1278 1000 1284 1001
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 1238 996 1244 997
rect 1238 992 1239 996
rect 1243 992 1244 996
rect 1278 996 1279 1000
rect 1283 996 1284 1000
rect 1278 995 1284 996
rect 2406 1000 2412 1001
rect 2406 996 2407 1000
rect 2411 996 2412 1000
rect 2406 995 2412 996
rect 1238 991 1244 992
rect 1278 983 1284 984
rect 110 979 116 980
rect 110 975 111 979
rect 115 975 116 979
rect 110 974 116 975
rect 1238 979 1244 980
rect 1238 975 1239 979
rect 1243 975 1244 979
rect 1278 979 1279 983
rect 1283 979 1284 983
rect 1278 978 1284 979
rect 2406 983 2412 984
rect 2406 979 2407 983
rect 2411 979 2412 983
rect 2406 978 2412 979
rect 1238 974 1244 975
rect 112 967 114 974
rect 174 972 180 973
rect 174 968 175 972
rect 179 968 180 972
rect 174 967 180 968
rect 254 972 260 973
rect 254 968 255 972
rect 259 968 260 972
rect 254 967 260 968
rect 326 972 332 973
rect 326 968 327 972
rect 331 968 332 972
rect 326 967 332 968
rect 398 972 404 973
rect 398 968 399 972
rect 403 968 404 972
rect 398 967 404 968
rect 462 972 468 973
rect 462 968 463 972
rect 467 968 468 972
rect 462 967 468 968
rect 518 972 524 973
rect 518 968 519 972
rect 523 968 524 972
rect 518 967 524 968
rect 574 972 580 973
rect 574 968 575 972
rect 579 968 580 972
rect 574 967 580 968
rect 622 972 628 973
rect 622 968 623 972
rect 627 968 628 972
rect 622 967 628 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 806 972 812 973
rect 806 968 807 972
rect 811 968 812 972
rect 806 967 812 968
rect 894 972 900 973
rect 894 968 895 972
rect 899 968 900 972
rect 894 967 900 968
rect 998 972 1004 973
rect 998 968 999 972
rect 1003 968 1004 972
rect 998 967 1004 968
rect 1102 972 1108 973
rect 1102 968 1103 972
rect 1107 968 1108 972
rect 1102 967 1108 968
rect 1190 972 1196 973
rect 1190 968 1191 972
rect 1195 968 1196 972
rect 1190 967 1196 968
rect 1240 967 1242 974
rect 111 966 115 967
rect 111 961 115 962
rect 175 966 179 967
rect 175 961 179 962
rect 215 966 219 967
rect 215 961 219 962
rect 255 966 259 967
rect 255 961 259 962
rect 303 966 307 967
rect 303 961 307 962
rect 327 966 331 967
rect 327 961 331 962
rect 359 966 363 967
rect 359 961 363 962
rect 399 966 403 967
rect 399 961 403 962
rect 415 966 419 967
rect 415 961 419 962
rect 463 966 467 967
rect 463 961 467 962
rect 519 966 523 967
rect 519 961 523 962
rect 575 966 579 967
rect 575 961 579 962
rect 623 966 627 967
rect 623 961 627 962
rect 639 966 643 967
rect 639 961 643 962
rect 671 966 675 967
rect 671 961 675 962
rect 711 966 715 967
rect 711 961 715 962
rect 735 966 739 967
rect 735 961 739 962
rect 783 966 787 967
rect 783 961 787 962
rect 807 966 811 967
rect 807 961 811 962
rect 855 966 859 967
rect 855 961 859 962
rect 895 966 899 967
rect 895 961 899 962
rect 927 966 931 967
rect 927 961 931 962
rect 999 966 1003 967
rect 999 961 1003 962
rect 1071 966 1075 967
rect 1071 961 1075 962
rect 1103 966 1107 967
rect 1103 961 1107 962
rect 1143 966 1147 967
rect 1143 961 1147 962
rect 1191 966 1195 967
rect 1191 961 1195 962
rect 1239 966 1243 967
rect 1280 963 1282 978
rect 1574 976 1580 977
rect 1574 972 1575 976
rect 1579 972 1580 976
rect 1574 971 1580 972
rect 1614 976 1620 977
rect 1614 972 1615 976
rect 1619 972 1620 976
rect 1614 971 1620 972
rect 1654 976 1660 977
rect 1654 972 1655 976
rect 1659 972 1660 976
rect 1654 971 1660 972
rect 1694 976 1700 977
rect 1694 972 1695 976
rect 1699 972 1700 976
rect 1694 971 1700 972
rect 1734 976 1740 977
rect 1734 972 1735 976
rect 1739 972 1740 976
rect 1734 971 1740 972
rect 1774 976 1780 977
rect 1774 972 1775 976
rect 1779 972 1780 976
rect 1774 971 1780 972
rect 1822 976 1828 977
rect 1822 972 1823 976
rect 1827 972 1828 976
rect 1822 971 1828 972
rect 1878 976 1884 977
rect 1878 972 1879 976
rect 1883 972 1884 976
rect 1878 971 1884 972
rect 1942 976 1948 977
rect 1942 972 1943 976
rect 1947 972 1948 976
rect 1942 971 1948 972
rect 2014 976 2020 977
rect 2014 972 2015 976
rect 2019 972 2020 976
rect 2014 971 2020 972
rect 2094 976 2100 977
rect 2094 972 2095 976
rect 2099 972 2100 976
rect 2094 971 2100 972
rect 2174 976 2180 977
rect 2174 972 2175 976
rect 2179 972 2180 976
rect 2174 971 2180 972
rect 2254 976 2260 977
rect 2254 972 2255 976
rect 2259 972 2260 976
rect 2254 971 2260 972
rect 1576 963 1578 971
rect 1616 963 1618 971
rect 1656 963 1658 971
rect 1696 963 1698 971
rect 1736 963 1738 971
rect 1776 963 1778 971
rect 1824 963 1826 971
rect 1880 963 1882 971
rect 1944 963 1946 971
rect 2016 963 2018 971
rect 2096 963 2098 971
rect 2176 963 2178 971
rect 2256 963 2258 971
rect 2408 963 2410 978
rect 1239 961 1243 962
rect 1279 962 1283 963
rect 112 954 114 961
rect 214 960 220 961
rect 214 956 215 960
rect 219 956 220 960
rect 214 955 220 956
rect 254 960 260 961
rect 254 956 255 960
rect 259 956 260 960
rect 254 955 260 956
rect 302 960 308 961
rect 302 956 303 960
rect 307 956 308 960
rect 302 955 308 956
rect 358 960 364 961
rect 358 956 359 960
rect 363 956 364 960
rect 358 955 364 956
rect 414 960 420 961
rect 414 956 415 960
rect 419 956 420 960
rect 414 955 420 956
rect 462 960 468 961
rect 462 956 463 960
rect 467 956 468 960
rect 462 955 468 956
rect 518 960 524 961
rect 518 956 519 960
rect 523 956 524 960
rect 518 955 524 956
rect 574 960 580 961
rect 574 956 575 960
rect 579 956 580 960
rect 574 955 580 956
rect 638 960 644 961
rect 638 956 639 960
rect 643 956 644 960
rect 638 955 644 956
rect 710 960 716 961
rect 710 956 711 960
rect 715 956 716 960
rect 710 955 716 956
rect 782 960 788 961
rect 782 956 783 960
rect 787 956 788 960
rect 782 955 788 956
rect 854 960 860 961
rect 854 956 855 960
rect 859 956 860 960
rect 854 955 860 956
rect 926 960 932 961
rect 926 956 927 960
rect 931 956 932 960
rect 926 955 932 956
rect 998 960 1004 961
rect 998 956 999 960
rect 1003 956 1004 960
rect 998 955 1004 956
rect 1070 960 1076 961
rect 1070 956 1071 960
rect 1075 956 1076 960
rect 1070 955 1076 956
rect 1142 960 1148 961
rect 1142 956 1143 960
rect 1147 956 1148 960
rect 1142 955 1148 956
rect 1190 960 1196 961
rect 1190 956 1191 960
rect 1195 956 1196 960
rect 1190 955 1196 956
rect 1240 954 1242 961
rect 1279 957 1283 958
rect 1303 962 1307 963
rect 1303 957 1307 958
rect 1351 962 1355 963
rect 1351 957 1355 958
rect 1431 962 1435 963
rect 1431 957 1435 958
rect 1511 962 1515 963
rect 1511 957 1515 958
rect 1575 962 1579 963
rect 1575 957 1579 958
rect 1591 962 1595 963
rect 1591 957 1595 958
rect 1615 962 1619 963
rect 1615 957 1619 958
rect 1655 962 1659 963
rect 1655 957 1659 958
rect 1679 962 1683 963
rect 1679 957 1683 958
rect 1695 962 1699 963
rect 1695 957 1699 958
rect 1735 962 1739 963
rect 1735 957 1739 958
rect 1767 962 1771 963
rect 1767 957 1771 958
rect 1775 962 1779 963
rect 1775 957 1779 958
rect 1823 962 1827 963
rect 1823 957 1827 958
rect 1855 962 1859 963
rect 1855 957 1859 958
rect 1879 962 1883 963
rect 1879 957 1883 958
rect 1943 962 1947 963
rect 1943 957 1947 958
rect 2015 962 2019 963
rect 2015 957 2019 958
rect 2023 962 2027 963
rect 2023 957 2027 958
rect 2095 962 2099 963
rect 2095 957 2099 958
rect 2103 962 2107 963
rect 2103 957 2107 958
rect 2175 962 2179 963
rect 2175 957 2179 958
rect 2183 962 2187 963
rect 2183 957 2187 958
rect 2255 962 2259 963
rect 2255 957 2259 958
rect 2271 962 2275 963
rect 2271 957 2275 958
rect 2407 962 2411 963
rect 2407 957 2411 958
rect 110 953 116 954
rect 110 949 111 953
rect 115 949 116 953
rect 110 948 116 949
rect 1238 953 1244 954
rect 1238 949 1239 953
rect 1243 949 1244 953
rect 1280 950 1282 957
rect 1302 956 1308 957
rect 1302 952 1303 956
rect 1307 952 1308 956
rect 1302 951 1308 952
rect 1350 956 1356 957
rect 1350 952 1351 956
rect 1355 952 1356 956
rect 1350 951 1356 952
rect 1430 956 1436 957
rect 1430 952 1431 956
rect 1435 952 1436 956
rect 1430 951 1436 952
rect 1510 956 1516 957
rect 1510 952 1511 956
rect 1515 952 1516 956
rect 1510 951 1516 952
rect 1590 956 1596 957
rect 1590 952 1591 956
rect 1595 952 1596 956
rect 1590 951 1596 952
rect 1678 956 1684 957
rect 1678 952 1679 956
rect 1683 952 1684 956
rect 1678 951 1684 952
rect 1766 956 1772 957
rect 1766 952 1767 956
rect 1771 952 1772 956
rect 1766 951 1772 952
rect 1854 956 1860 957
rect 1854 952 1855 956
rect 1859 952 1860 956
rect 1854 951 1860 952
rect 1942 956 1948 957
rect 1942 952 1943 956
rect 1947 952 1948 956
rect 1942 951 1948 952
rect 2022 956 2028 957
rect 2022 952 2023 956
rect 2027 952 2028 956
rect 2022 951 2028 952
rect 2102 956 2108 957
rect 2102 952 2103 956
rect 2107 952 2108 956
rect 2102 951 2108 952
rect 2182 956 2188 957
rect 2182 952 2183 956
rect 2187 952 2188 956
rect 2182 951 2188 952
rect 2270 956 2276 957
rect 2270 952 2271 956
rect 2275 952 2276 956
rect 2270 951 2276 952
rect 2408 950 2410 957
rect 1238 948 1244 949
rect 1278 949 1284 950
rect 1278 945 1279 949
rect 1283 945 1284 949
rect 1278 944 1284 945
rect 2406 949 2412 950
rect 2406 945 2407 949
rect 2411 945 2412 949
rect 2406 944 2412 945
rect 110 936 116 937
rect 110 932 111 936
rect 115 932 116 936
rect 110 931 116 932
rect 1238 936 1244 937
rect 1238 932 1239 936
rect 1243 932 1244 936
rect 1238 931 1244 932
rect 1278 932 1284 933
rect 112 891 114 931
rect 214 913 220 914
rect 214 909 215 913
rect 219 909 220 913
rect 214 908 220 909
rect 254 913 260 914
rect 254 909 255 913
rect 259 909 260 913
rect 254 908 260 909
rect 302 913 308 914
rect 302 909 303 913
rect 307 909 308 913
rect 302 908 308 909
rect 358 913 364 914
rect 358 909 359 913
rect 363 909 364 913
rect 358 908 364 909
rect 414 913 420 914
rect 414 909 415 913
rect 419 909 420 913
rect 414 908 420 909
rect 462 913 468 914
rect 462 909 463 913
rect 467 909 468 913
rect 462 908 468 909
rect 518 913 524 914
rect 518 909 519 913
rect 523 909 524 913
rect 518 908 524 909
rect 574 913 580 914
rect 574 909 575 913
rect 579 909 580 913
rect 574 908 580 909
rect 638 913 644 914
rect 638 909 639 913
rect 643 909 644 913
rect 638 908 644 909
rect 710 913 716 914
rect 710 909 711 913
rect 715 909 716 913
rect 710 908 716 909
rect 782 913 788 914
rect 782 909 783 913
rect 787 909 788 913
rect 782 908 788 909
rect 854 913 860 914
rect 854 909 855 913
rect 859 909 860 913
rect 854 908 860 909
rect 926 913 932 914
rect 926 909 927 913
rect 931 909 932 913
rect 926 908 932 909
rect 998 913 1004 914
rect 998 909 999 913
rect 1003 909 1004 913
rect 998 908 1004 909
rect 1070 913 1076 914
rect 1070 909 1071 913
rect 1075 909 1076 913
rect 1070 908 1076 909
rect 1142 913 1148 914
rect 1142 909 1143 913
rect 1147 909 1148 913
rect 1142 908 1148 909
rect 1190 913 1196 914
rect 1190 909 1191 913
rect 1195 909 1196 913
rect 1190 908 1196 909
rect 216 891 218 908
rect 256 891 258 908
rect 304 891 306 908
rect 360 891 362 908
rect 416 891 418 908
rect 464 891 466 908
rect 520 891 522 908
rect 576 891 578 908
rect 640 891 642 908
rect 712 891 714 908
rect 784 891 786 908
rect 856 891 858 908
rect 928 891 930 908
rect 1000 891 1002 908
rect 1072 891 1074 908
rect 1144 891 1146 908
rect 1192 891 1194 908
rect 1240 891 1242 931
rect 1278 928 1279 932
rect 1283 928 1284 932
rect 1278 927 1284 928
rect 2406 932 2412 933
rect 2406 928 2407 932
rect 2411 928 2412 932
rect 2406 927 2412 928
rect 1280 895 1282 927
rect 1302 909 1308 910
rect 1302 905 1303 909
rect 1307 905 1308 909
rect 1302 904 1308 905
rect 1350 909 1356 910
rect 1350 905 1351 909
rect 1355 905 1356 909
rect 1350 904 1356 905
rect 1430 909 1436 910
rect 1430 905 1431 909
rect 1435 905 1436 909
rect 1430 904 1436 905
rect 1510 909 1516 910
rect 1510 905 1511 909
rect 1515 905 1516 909
rect 1510 904 1516 905
rect 1590 909 1596 910
rect 1590 905 1591 909
rect 1595 905 1596 909
rect 1590 904 1596 905
rect 1678 909 1684 910
rect 1678 905 1679 909
rect 1683 905 1684 909
rect 1678 904 1684 905
rect 1766 909 1772 910
rect 1766 905 1767 909
rect 1771 905 1772 909
rect 1766 904 1772 905
rect 1854 909 1860 910
rect 1854 905 1855 909
rect 1859 905 1860 909
rect 1854 904 1860 905
rect 1942 909 1948 910
rect 1942 905 1943 909
rect 1947 905 1948 909
rect 1942 904 1948 905
rect 2022 909 2028 910
rect 2022 905 2023 909
rect 2027 905 2028 909
rect 2022 904 2028 905
rect 2102 909 2108 910
rect 2102 905 2103 909
rect 2107 905 2108 909
rect 2102 904 2108 905
rect 2182 909 2188 910
rect 2182 905 2183 909
rect 2187 905 2188 909
rect 2182 904 2188 905
rect 2270 909 2276 910
rect 2270 905 2271 909
rect 2275 905 2276 909
rect 2270 904 2276 905
rect 1304 895 1306 904
rect 1352 895 1354 904
rect 1432 895 1434 904
rect 1512 895 1514 904
rect 1592 895 1594 904
rect 1680 895 1682 904
rect 1768 895 1770 904
rect 1856 895 1858 904
rect 1944 895 1946 904
rect 2024 895 2026 904
rect 2104 895 2106 904
rect 2184 895 2186 904
rect 2272 895 2274 904
rect 2408 895 2410 927
rect 1279 894 1283 895
rect 111 890 115 891
rect 111 885 115 886
rect 191 890 195 891
rect 191 885 195 886
rect 215 890 219 891
rect 215 885 219 886
rect 231 890 235 891
rect 231 885 235 886
rect 255 890 259 891
rect 255 885 259 886
rect 287 890 291 891
rect 287 885 291 886
rect 303 890 307 891
rect 303 885 307 886
rect 359 890 363 891
rect 359 885 363 886
rect 415 890 419 891
rect 415 885 419 886
rect 447 890 451 891
rect 447 885 451 886
rect 463 890 467 891
rect 463 885 467 886
rect 519 890 523 891
rect 519 885 523 886
rect 543 890 547 891
rect 543 885 547 886
rect 575 890 579 891
rect 575 885 579 886
rect 639 890 643 891
rect 639 885 643 886
rect 711 890 715 891
rect 711 885 715 886
rect 727 890 731 891
rect 727 885 731 886
rect 783 890 787 891
rect 783 885 787 886
rect 807 890 811 891
rect 807 885 811 886
rect 855 890 859 891
rect 855 885 859 886
rect 887 890 891 891
rect 887 885 891 886
rect 927 890 931 891
rect 927 885 931 886
rect 959 890 963 891
rect 959 885 963 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 1023 890 1027 891
rect 1023 885 1027 886
rect 1071 890 1075 891
rect 1071 885 1075 886
rect 1087 890 1091 891
rect 1087 885 1091 886
rect 1143 890 1147 891
rect 1143 885 1147 886
rect 1159 890 1163 891
rect 1159 885 1163 886
rect 1191 890 1195 891
rect 1191 885 1195 886
rect 1239 890 1243 891
rect 1279 889 1283 890
rect 1303 894 1307 895
rect 1303 889 1307 890
rect 1351 894 1355 895
rect 1351 889 1355 890
rect 1431 894 1435 895
rect 1431 889 1435 890
rect 1439 894 1443 895
rect 1439 889 1443 890
rect 1479 894 1483 895
rect 1479 889 1483 890
rect 1511 894 1515 895
rect 1511 889 1515 890
rect 1519 894 1523 895
rect 1519 889 1523 890
rect 1559 894 1563 895
rect 1559 889 1563 890
rect 1591 894 1595 895
rect 1591 889 1595 890
rect 1607 894 1611 895
rect 1607 889 1611 890
rect 1655 894 1659 895
rect 1655 889 1659 890
rect 1679 894 1683 895
rect 1679 889 1683 890
rect 1711 894 1715 895
rect 1711 889 1715 890
rect 1767 894 1771 895
rect 1767 889 1771 890
rect 1775 894 1779 895
rect 1775 889 1779 890
rect 1847 894 1851 895
rect 1847 889 1851 890
rect 1855 894 1859 895
rect 1855 889 1859 890
rect 1919 894 1923 895
rect 1919 889 1923 890
rect 1943 894 1947 895
rect 1943 889 1947 890
rect 1991 894 1995 895
rect 1991 889 1995 890
rect 2023 894 2027 895
rect 2023 889 2027 890
rect 2063 894 2067 895
rect 2063 889 2067 890
rect 2103 894 2107 895
rect 2103 889 2107 890
rect 2135 894 2139 895
rect 2135 889 2139 890
rect 2183 894 2187 895
rect 2183 889 2187 890
rect 2215 894 2219 895
rect 2215 889 2219 890
rect 2271 894 2275 895
rect 2271 889 2275 890
rect 2295 894 2299 895
rect 2295 889 2299 890
rect 2407 894 2411 895
rect 2407 889 2411 890
rect 1239 885 1243 886
rect 112 853 114 885
rect 192 876 194 885
rect 232 876 234 885
rect 288 876 290 885
rect 360 876 362 885
rect 448 876 450 885
rect 544 876 546 885
rect 640 876 642 885
rect 728 876 730 885
rect 808 876 810 885
rect 888 876 890 885
rect 960 876 962 885
rect 1024 876 1026 885
rect 1088 876 1090 885
rect 1160 876 1162 885
rect 190 875 196 876
rect 190 871 191 875
rect 195 871 196 875
rect 190 870 196 871
rect 230 875 236 876
rect 230 871 231 875
rect 235 871 236 875
rect 230 870 236 871
rect 286 875 292 876
rect 286 871 287 875
rect 291 871 292 875
rect 286 870 292 871
rect 358 875 364 876
rect 358 871 359 875
rect 363 871 364 875
rect 358 870 364 871
rect 446 875 452 876
rect 446 871 447 875
rect 451 871 452 875
rect 446 870 452 871
rect 542 875 548 876
rect 542 871 543 875
rect 547 871 548 875
rect 542 870 548 871
rect 638 875 644 876
rect 638 871 639 875
rect 643 871 644 875
rect 638 870 644 871
rect 726 875 732 876
rect 726 871 727 875
rect 731 871 732 875
rect 726 870 732 871
rect 806 875 812 876
rect 806 871 807 875
rect 811 871 812 875
rect 806 870 812 871
rect 886 875 892 876
rect 886 871 887 875
rect 891 871 892 875
rect 886 870 892 871
rect 958 875 964 876
rect 958 871 959 875
rect 963 871 964 875
rect 958 870 964 871
rect 1022 875 1028 876
rect 1022 871 1023 875
rect 1027 871 1028 875
rect 1022 870 1028 871
rect 1086 875 1092 876
rect 1086 871 1087 875
rect 1091 871 1092 875
rect 1086 870 1092 871
rect 1158 875 1164 876
rect 1158 871 1159 875
rect 1163 871 1164 875
rect 1158 870 1164 871
rect 1240 853 1242 885
rect 1280 857 1282 889
rect 1440 880 1442 889
rect 1480 880 1482 889
rect 1520 880 1522 889
rect 1560 880 1562 889
rect 1608 880 1610 889
rect 1656 880 1658 889
rect 1712 880 1714 889
rect 1776 880 1778 889
rect 1848 880 1850 889
rect 1920 880 1922 889
rect 1992 880 1994 889
rect 2064 880 2066 889
rect 2136 880 2138 889
rect 2216 880 2218 889
rect 2296 880 2298 889
rect 1438 879 1444 880
rect 1438 875 1439 879
rect 1443 875 1444 879
rect 1438 874 1444 875
rect 1478 879 1484 880
rect 1478 875 1479 879
rect 1483 875 1484 879
rect 1478 874 1484 875
rect 1518 879 1524 880
rect 1518 875 1519 879
rect 1523 875 1524 879
rect 1518 874 1524 875
rect 1558 879 1564 880
rect 1558 875 1559 879
rect 1563 875 1564 879
rect 1558 874 1564 875
rect 1606 879 1612 880
rect 1606 875 1607 879
rect 1611 875 1612 879
rect 1606 874 1612 875
rect 1654 879 1660 880
rect 1654 875 1655 879
rect 1659 875 1660 879
rect 1654 874 1660 875
rect 1710 879 1716 880
rect 1710 875 1711 879
rect 1715 875 1716 879
rect 1710 874 1716 875
rect 1774 879 1780 880
rect 1774 875 1775 879
rect 1779 875 1780 879
rect 1774 874 1780 875
rect 1846 879 1852 880
rect 1846 875 1847 879
rect 1851 875 1852 879
rect 1846 874 1852 875
rect 1918 879 1924 880
rect 1918 875 1919 879
rect 1923 875 1924 879
rect 1918 874 1924 875
rect 1990 879 1996 880
rect 1990 875 1991 879
rect 1995 875 1996 879
rect 1990 874 1996 875
rect 2062 879 2068 880
rect 2062 875 2063 879
rect 2067 875 2068 879
rect 2062 874 2068 875
rect 2134 879 2140 880
rect 2134 875 2135 879
rect 2139 875 2140 879
rect 2134 874 2140 875
rect 2214 879 2220 880
rect 2214 875 2215 879
rect 2219 875 2220 879
rect 2214 874 2220 875
rect 2294 879 2300 880
rect 2294 875 2295 879
rect 2299 875 2300 879
rect 2294 874 2300 875
rect 2408 857 2410 889
rect 1278 856 1284 857
rect 110 852 116 853
rect 110 848 111 852
rect 115 848 116 852
rect 110 847 116 848
rect 1238 852 1244 853
rect 1238 848 1239 852
rect 1243 848 1244 852
rect 1278 852 1279 856
rect 1283 852 1284 856
rect 1278 851 1284 852
rect 2406 856 2412 857
rect 2406 852 2407 856
rect 2411 852 2412 856
rect 2406 851 2412 852
rect 1238 847 1244 848
rect 1278 839 1284 840
rect 110 835 116 836
rect 110 831 111 835
rect 115 831 116 835
rect 110 830 116 831
rect 1238 835 1244 836
rect 1238 831 1239 835
rect 1243 831 1244 835
rect 1278 835 1279 839
rect 1283 835 1284 839
rect 1278 834 1284 835
rect 2406 839 2412 840
rect 2406 835 2407 839
rect 2411 835 2412 839
rect 2406 834 2412 835
rect 1238 830 1244 831
rect 112 823 114 830
rect 190 828 196 829
rect 190 824 191 828
rect 195 824 196 828
rect 190 823 196 824
rect 230 828 236 829
rect 230 824 231 828
rect 235 824 236 828
rect 230 823 236 824
rect 286 828 292 829
rect 286 824 287 828
rect 291 824 292 828
rect 286 823 292 824
rect 358 828 364 829
rect 358 824 359 828
rect 363 824 364 828
rect 358 823 364 824
rect 446 828 452 829
rect 446 824 447 828
rect 451 824 452 828
rect 446 823 452 824
rect 542 828 548 829
rect 542 824 543 828
rect 547 824 548 828
rect 542 823 548 824
rect 638 828 644 829
rect 638 824 639 828
rect 643 824 644 828
rect 638 823 644 824
rect 726 828 732 829
rect 726 824 727 828
rect 731 824 732 828
rect 726 823 732 824
rect 806 828 812 829
rect 806 824 807 828
rect 811 824 812 828
rect 806 823 812 824
rect 886 828 892 829
rect 886 824 887 828
rect 891 824 892 828
rect 886 823 892 824
rect 958 828 964 829
rect 958 824 959 828
rect 963 824 964 828
rect 958 823 964 824
rect 1022 828 1028 829
rect 1022 824 1023 828
rect 1027 824 1028 828
rect 1022 823 1028 824
rect 1086 828 1092 829
rect 1086 824 1087 828
rect 1091 824 1092 828
rect 1086 823 1092 824
rect 1158 828 1164 829
rect 1158 824 1159 828
rect 1163 824 1164 828
rect 1158 823 1164 824
rect 1240 823 1242 830
rect 111 822 115 823
rect 111 817 115 818
rect 135 822 139 823
rect 135 817 139 818
rect 175 822 179 823
rect 175 817 179 818
rect 191 822 195 823
rect 191 817 195 818
rect 231 822 235 823
rect 231 817 235 818
rect 239 822 243 823
rect 239 817 243 818
rect 287 822 291 823
rect 287 817 291 818
rect 327 822 331 823
rect 327 817 331 818
rect 359 822 363 823
rect 359 817 363 818
rect 415 822 419 823
rect 415 817 419 818
rect 447 822 451 823
rect 447 817 451 818
rect 503 822 507 823
rect 503 817 507 818
rect 543 822 547 823
rect 543 817 547 818
rect 591 822 595 823
rect 591 817 595 818
rect 639 822 643 823
rect 639 817 643 818
rect 671 822 675 823
rect 671 817 675 818
rect 727 822 731 823
rect 727 817 731 818
rect 743 822 747 823
rect 743 817 747 818
rect 807 822 811 823
rect 807 817 811 818
rect 815 822 819 823
rect 815 817 819 818
rect 879 822 883 823
rect 879 817 883 818
rect 887 822 891 823
rect 887 817 891 818
rect 943 822 947 823
rect 943 817 947 818
rect 959 822 963 823
rect 959 817 963 818
rect 1015 822 1019 823
rect 1015 817 1019 818
rect 1023 822 1027 823
rect 1023 817 1027 818
rect 1087 822 1091 823
rect 1087 817 1091 818
rect 1159 822 1163 823
rect 1159 817 1163 818
rect 1239 822 1243 823
rect 1239 817 1243 818
rect 112 810 114 817
rect 134 816 140 817
rect 134 812 135 816
rect 139 812 140 816
rect 134 811 140 812
rect 174 816 180 817
rect 174 812 175 816
rect 179 812 180 816
rect 174 811 180 812
rect 238 816 244 817
rect 238 812 239 816
rect 243 812 244 816
rect 238 811 244 812
rect 326 816 332 817
rect 326 812 327 816
rect 331 812 332 816
rect 326 811 332 812
rect 414 816 420 817
rect 414 812 415 816
rect 419 812 420 816
rect 414 811 420 812
rect 502 816 508 817
rect 502 812 503 816
rect 507 812 508 816
rect 502 811 508 812
rect 590 816 596 817
rect 590 812 591 816
rect 595 812 596 816
rect 590 811 596 812
rect 670 816 676 817
rect 670 812 671 816
rect 675 812 676 816
rect 670 811 676 812
rect 742 816 748 817
rect 742 812 743 816
rect 747 812 748 816
rect 742 811 748 812
rect 814 816 820 817
rect 814 812 815 816
rect 819 812 820 816
rect 814 811 820 812
rect 878 816 884 817
rect 878 812 879 816
rect 883 812 884 816
rect 878 811 884 812
rect 942 816 948 817
rect 942 812 943 816
rect 947 812 948 816
rect 942 811 948 812
rect 1014 816 1020 817
rect 1014 812 1015 816
rect 1019 812 1020 816
rect 1014 811 1020 812
rect 1240 810 1242 817
rect 1280 815 1282 834
rect 1438 832 1444 833
rect 1438 828 1439 832
rect 1443 828 1444 832
rect 1438 827 1444 828
rect 1478 832 1484 833
rect 1478 828 1479 832
rect 1483 828 1484 832
rect 1478 827 1484 828
rect 1518 832 1524 833
rect 1518 828 1519 832
rect 1523 828 1524 832
rect 1518 827 1524 828
rect 1558 832 1564 833
rect 1558 828 1559 832
rect 1563 828 1564 832
rect 1558 827 1564 828
rect 1606 832 1612 833
rect 1606 828 1607 832
rect 1611 828 1612 832
rect 1606 827 1612 828
rect 1654 832 1660 833
rect 1654 828 1655 832
rect 1659 828 1660 832
rect 1654 827 1660 828
rect 1710 832 1716 833
rect 1710 828 1711 832
rect 1715 828 1716 832
rect 1710 827 1716 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1846 832 1852 833
rect 1846 828 1847 832
rect 1851 828 1852 832
rect 1846 827 1852 828
rect 1918 832 1924 833
rect 1918 828 1919 832
rect 1923 828 1924 832
rect 1918 827 1924 828
rect 1990 832 1996 833
rect 1990 828 1991 832
rect 1995 828 1996 832
rect 1990 827 1996 828
rect 2062 832 2068 833
rect 2062 828 2063 832
rect 2067 828 2068 832
rect 2062 827 2068 828
rect 2134 832 2140 833
rect 2134 828 2135 832
rect 2139 828 2140 832
rect 2134 827 2140 828
rect 2214 832 2220 833
rect 2214 828 2215 832
rect 2219 828 2220 832
rect 2214 827 2220 828
rect 2294 832 2300 833
rect 2294 828 2295 832
rect 2299 828 2300 832
rect 2294 827 2300 828
rect 1440 815 1442 827
rect 1480 815 1482 827
rect 1520 815 1522 827
rect 1560 815 1562 827
rect 1608 815 1610 827
rect 1656 815 1658 827
rect 1712 815 1714 827
rect 1776 815 1778 827
rect 1848 815 1850 827
rect 1920 815 1922 827
rect 1992 815 1994 827
rect 2064 815 2066 827
rect 2136 815 2138 827
rect 2216 815 2218 827
rect 2296 815 2298 827
rect 2408 815 2410 834
rect 1279 814 1283 815
rect 110 809 116 810
rect 110 805 111 809
rect 115 805 116 809
rect 110 804 116 805
rect 1238 809 1244 810
rect 1279 809 1283 810
rect 1359 814 1363 815
rect 1359 809 1363 810
rect 1415 814 1419 815
rect 1415 809 1419 810
rect 1439 814 1443 815
rect 1439 809 1443 810
rect 1471 814 1475 815
rect 1471 809 1475 810
rect 1479 814 1483 815
rect 1479 809 1483 810
rect 1519 814 1523 815
rect 1519 809 1523 810
rect 1535 814 1539 815
rect 1535 809 1539 810
rect 1559 814 1563 815
rect 1559 809 1563 810
rect 1591 814 1595 815
rect 1591 809 1595 810
rect 1607 814 1611 815
rect 1607 809 1611 810
rect 1647 814 1651 815
rect 1647 809 1651 810
rect 1655 814 1659 815
rect 1655 809 1659 810
rect 1703 814 1707 815
rect 1703 809 1707 810
rect 1711 814 1715 815
rect 1711 809 1715 810
rect 1759 814 1763 815
rect 1759 809 1763 810
rect 1775 814 1779 815
rect 1775 809 1779 810
rect 1815 814 1819 815
rect 1815 809 1819 810
rect 1847 814 1851 815
rect 1847 809 1851 810
rect 1871 814 1875 815
rect 1871 809 1875 810
rect 1919 814 1923 815
rect 1919 809 1923 810
rect 1935 814 1939 815
rect 1935 809 1939 810
rect 1991 814 1995 815
rect 1991 809 1995 810
rect 1999 814 2003 815
rect 1999 809 2003 810
rect 2063 814 2067 815
rect 2063 809 2067 810
rect 2071 814 2075 815
rect 2071 809 2075 810
rect 2135 814 2139 815
rect 2135 809 2139 810
rect 2143 814 2147 815
rect 2143 809 2147 810
rect 2215 814 2219 815
rect 2215 809 2219 810
rect 2223 814 2227 815
rect 2223 809 2227 810
rect 2295 814 2299 815
rect 2295 809 2299 810
rect 2303 814 2307 815
rect 2303 809 2307 810
rect 2359 814 2363 815
rect 2359 809 2363 810
rect 2407 814 2411 815
rect 2407 809 2411 810
rect 1238 805 1239 809
rect 1243 805 1244 809
rect 1238 804 1244 805
rect 1280 802 1282 809
rect 1358 808 1364 809
rect 1358 804 1359 808
rect 1363 804 1364 808
rect 1358 803 1364 804
rect 1414 808 1420 809
rect 1414 804 1415 808
rect 1419 804 1420 808
rect 1414 803 1420 804
rect 1470 808 1476 809
rect 1470 804 1471 808
rect 1475 804 1476 808
rect 1470 803 1476 804
rect 1534 808 1540 809
rect 1534 804 1535 808
rect 1539 804 1540 808
rect 1534 803 1540 804
rect 1590 808 1596 809
rect 1590 804 1591 808
rect 1595 804 1596 808
rect 1590 803 1596 804
rect 1646 808 1652 809
rect 1646 804 1647 808
rect 1651 804 1652 808
rect 1646 803 1652 804
rect 1702 808 1708 809
rect 1702 804 1703 808
rect 1707 804 1708 808
rect 1702 803 1708 804
rect 1758 808 1764 809
rect 1758 804 1759 808
rect 1763 804 1764 808
rect 1758 803 1764 804
rect 1814 808 1820 809
rect 1814 804 1815 808
rect 1819 804 1820 808
rect 1814 803 1820 804
rect 1870 808 1876 809
rect 1870 804 1871 808
rect 1875 804 1876 808
rect 1870 803 1876 804
rect 1934 808 1940 809
rect 1934 804 1935 808
rect 1939 804 1940 808
rect 1934 803 1940 804
rect 1998 808 2004 809
rect 1998 804 1999 808
rect 2003 804 2004 808
rect 1998 803 2004 804
rect 2070 808 2076 809
rect 2070 804 2071 808
rect 2075 804 2076 808
rect 2070 803 2076 804
rect 2142 808 2148 809
rect 2142 804 2143 808
rect 2147 804 2148 808
rect 2142 803 2148 804
rect 2222 808 2228 809
rect 2222 804 2223 808
rect 2227 804 2228 808
rect 2222 803 2228 804
rect 2302 808 2308 809
rect 2302 804 2303 808
rect 2307 804 2308 808
rect 2302 803 2308 804
rect 2358 808 2364 809
rect 2358 804 2359 808
rect 2363 804 2364 808
rect 2358 803 2364 804
rect 2408 802 2410 809
rect 1278 801 1284 802
rect 1278 797 1279 801
rect 1283 797 1284 801
rect 1278 796 1284 797
rect 2406 801 2412 802
rect 2406 797 2407 801
rect 2411 797 2412 801
rect 2406 796 2412 797
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 110 787 116 788
rect 1238 792 1244 793
rect 1238 788 1239 792
rect 1243 788 1244 792
rect 1238 787 1244 788
rect 112 751 114 787
rect 134 769 140 770
rect 134 765 135 769
rect 139 765 140 769
rect 134 764 140 765
rect 174 769 180 770
rect 174 765 175 769
rect 179 765 180 769
rect 174 764 180 765
rect 238 769 244 770
rect 238 765 239 769
rect 243 765 244 769
rect 238 764 244 765
rect 326 769 332 770
rect 326 765 327 769
rect 331 765 332 769
rect 326 764 332 765
rect 414 769 420 770
rect 414 765 415 769
rect 419 765 420 769
rect 414 764 420 765
rect 502 769 508 770
rect 502 765 503 769
rect 507 765 508 769
rect 502 764 508 765
rect 590 769 596 770
rect 590 765 591 769
rect 595 765 596 769
rect 590 764 596 765
rect 670 769 676 770
rect 670 765 671 769
rect 675 765 676 769
rect 670 764 676 765
rect 742 769 748 770
rect 742 765 743 769
rect 747 765 748 769
rect 742 764 748 765
rect 814 769 820 770
rect 814 765 815 769
rect 819 765 820 769
rect 814 764 820 765
rect 878 769 884 770
rect 878 765 879 769
rect 883 765 884 769
rect 878 764 884 765
rect 942 769 948 770
rect 942 765 943 769
rect 947 765 948 769
rect 942 764 948 765
rect 1014 769 1020 770
rect 1014 765 1015 769
rect 1019 765 1020 769
rect 1014 764 1020 765
rect 136 751 138 764
rect 176 751 178 764
rect 240 751 242 764
rect 328 751 330 764
rect 416 751 418 764
rect 504 751 506 764
rect 592 751 594 764
rect 672 751 674 764
rect 744 751 746 764
rect 816 751 818 764
rect 880 751 882 764
rect 944 751 946 764
rect 1016 751 1018 764
rect 1240 751 1242 787
rect 1278 784 1284 785
rect 1278 780 1279 784
rect 1283 780 1284 784
rect 1278 779 1284 780
rect 2406 784 2412 785
rect 2406 780 2407 784
rect 2411 780 2412 784
rect 2406 779 2412 780
rect 111 750 115 751
rect 111 745 115 746
rect 135 750 139 751
rect 135 745 139 746
rect 175 750 179 751
rect 175 745 179 746
rect 191 750 195 751
rect 191 745 195 746
rect 239 750 243 751
rect 239 745 243 746
rect 263 750 267 751
rect 263 745 267 746
rect 327 750 331 751
rect 327 745 331 746
rect 335 750 339 751
rect 335 745 339 746
rect 399 750 403 751
rect 399 745 403 746
rect 415 750 419 751
rect 415 745 419 746
rect 455 750 459 751
rect 455 745 459 746
rect 503 750 507 751
rect 503 745 507 746
rect 543 750 547 751
rect 543 745 547 746
rect 583 750 587 751
rect 583 745 587 746
rect 591 750 595 751
rect 591 745 595 746
rect 623 750 627 751
rect 623 745 627 746
rect 671 750 675 751
rect 671 745 675 746
rect 719 750 723 751
rect 719 745 723 746
rect 743 750 747 751
rect 743 745 747 746
rect 767 750 771 751
rect 767 745 771 746
rect 815 750 819 751
rect 815 745 819 746
rect 863 750 867 751
rect 863 745 867 746
rect 879 750 883 751
rect 879 745 883 746
rect 911 750 915 751
rect 911 745 915 746
rect 943 750 947 751
rect 943 745 947 746
rect 1015 750 1019 751
rect 1015 745 1019 746
rect 1239 750 1243 751
rect 1280 747 1282 779
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1534 761 1540 762
rect 1534 757 1535 761
rect 1539 757 1540 761
rect 1534 756 1540 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1590 756 1596 757
rect 1646 761 1652 762
rect 1646 757 1647 761
rect 1651 757 1652 761
rect 1646 756 1652 757
rect 1702 761 1708 762
rect 1702 757 1703 761
rect 1707 757 1708 761
rect 1702 756 1708 757
rect 1758 761 1764 762
rect 1758 757 1759 761
rect 1763 757 1764 761
rect 1758 756 1764 757
rect 1814 761 1820 762
rect 1814 757 1815 761
rect 1819 757 1820 761
rect 1814 756 1820 757
rect 1870 761 1876 762
rect 1870 757 1871 761
rect 1875 757 1876 761
rect 1870 756 1876 757
rect 1934 761 1940 762
rect 1934 757 1935 761
rect 1939 757 1940 761
rect 1934 756 1940 757
rect 1998 761 2004 762
rect 1998 757 1999 761
rect 2003 757 2004 761
rect 1998 756 2004 757
rect 2070 761 2076 762
rect 2070 757 2071 761
rect 2075 757 2076 761
rect 2070 756 2076 757
rect 2142 761 2148 762
rect 2142 757 2143 761
rect 2147 757 2148 761
rect 2142 756 2148 757
rect 2222 761 2228 762
rect 2222 757 2223 761
rect 2227 757 2228 761
rect 2222 756 2228 757
rect 2302 761 2308 762
rect 2302 757 2303 761
rect 2307 757 2308 761
rect 2302 756 2308 757
rect 2358 761 2364 762
rect 2358 757 2359 761
rect 2363 757 2364 761
rect 2358 756 2364 757
rect 1360 747 1362 756
rect 1416 747 1418 756
rect 1472 747 1474 756
rect 1536 747 1538 756
rect 1592 747 1594 756
rect 1648 747 1650 756
rect 1704 747 1706 756
rect 1760 747 1762 756
rect 1816 747 1818 756
rect 1872 747 1874 756
rect 1936 747 1938 756
rect 2000 747 2002 756
rect 2072 747 2074 756
rect 2144 747 2146 756
rect 2224 747 2226 756
rect 2304 747 2306 756
rect 2360 747 2362 756
rect 2408 747 2410 779
rect 1239 745 1243 746
rect 1279 746 1283 747
rect 112 713 114 745
rect 136 736 138 745
rect 192 736 194 745
rect 264 736 266 745
rect 336 736 338 745
rect 400 736 402 745
rect 456 736 458 745
rect 504 736 506 745
rect 544 736 546 745
rect 584 736 586 745
rect 624 736 626 745
rect 672 736 674 745
rect 720 736 722 745
rect 768 736 770 745
rect 816 736 818 745
rect 864 736 866 745
rect 912 736 914 745
rect 134 735 140 736
rect 134 731 135 735
rect 139 731 140 735
rect 134 730 140 731
rect 190 735 196 736
rect 190 731 191 735
rect 195 731 196 735
rect 190 730 196 731
rect 262 735 268 736
rect 262 731 263 735
rect 267 731 268 735
rect 262 730 268 731
rect 334 735 340 736
rect 334 731 335 735
rect 339 731 340 735
rect 334 730 340 731
rect 398 735 404 736
rect 398 731 399 735
rect 403 731 404 735
rect 398 730 404 731
rect 454 735 460 736
rect 454 731 455 735
rect 459 731 460 735
rect 454 730 460 731
rect 502 735 508 736
rect 502 731 503 735
rect 507 731 508 735
rect 502 730 508 731
rect 542 735 548 736
rect 542 731 543 735
rect 547 731 548 735
rect 542 730 548 731
rect 582 735 588 736
rect 582 731 583 735
rect 587 731 588 735
rect 582 730 588 731
rect 622 735 628 736
rect 622 731 623 735
rect 627 731 628 735
rect 622 730 628 731
rect 670 735 676 736
rect 670 731 671 735
rect 675 731 676 735
rect 670 730 676 731
rect 718 735 724 736
rect 718 731 719 735
rect 723 731 724 735
rect 718 730 724 731
rect 766 735 772 736
rect 766 731 767 735
rect 771 731 772 735
rect 766 730 772 731
rect 814 735 820 736
rect 814 731 815 735
rect 819 731 820 735
rect 814 730 820 731
rect 862 735 868 736
rect 862 731 863 735
rect 867 731 868 735
rect 862 730 868 731
rect 910 735 916 736
rect 910 731 911 735
rect 915 731 916 735
rect 910 730 916 731
rect 1240 713 1242 745
rect 1279 741 1283 742
rect 1303 746 1307 747
rect 1303 741 1307 742
rect 1343 746 1347 747
rect 1343 741 1347 742
rect 1359 746 1363 747
rect 1359 741 1363 742
rect 1407 746 1411 747
rect 1407 741 1411 742
rect 1415 746 1419 747
rect 1415 741 1419 742
rect 1471 746 1475 747
rect 1471 741 1475 742
rect 1487 746 1491 747
rect 1487 741 1491 742
rect 1535 746 1539 747
rect 1535 741 1539 742
rect 1575 746 1579 747
rect 1575 741 1579 742
rect 1591 746 1595 747
rect 1591 741 1595 742
rect 1647 746 1651 747
rect 1647 741 1651 742
rect 1663 746 1667 747
rect 1663 741 1667 742
rect 1703 746 1707 747
rect 1703 741 1707 742
rect 1751 746 1755 747
rect 1751 741 1755 742
rect 1759 746 1763 747
rect 1759 741 1763 742
rect 1815 746 1819 747
rect 1815 741 1819 742
rect 1831 746 1835 747
rect 1831 741 1835 742
rect 1871 746 1875 747
rect 1871 741 1875 742
rect 1911 746 1915 747
rect 1911 741 1915 742
rect 1935 746 1939 747
rect 1935 741 1939 742
rect 1991 746 1995 747
rect 1991 741 1995 742
rect 1999 746 2003 747
rect 1999 741 2003 742
rect 2071 746 2075 747
rect 2071 741 2075 742
rect 2079 746 2083 747
rect 2079 741 2083 742
rect 2143 746 2147 747
rect 2143 741 2147 742
rect 2175 746 2179 747
rect 2175 741 2179 742
rect 2223 746 2227 747
rect 2223 741 2227 742
rect 2279 746 2283 747
rect 2279 741 2283 742
rect 2303 746 2307 747
rect 2303 741 2307 742
rect 2359 746 2363 747
rect 2359 741 2363 742
rect 2407 746 2411 747
rect 2407 741 2411 742
rect 110 712 116 713
rect 110 708 111 712
rect 115 708 116 712
rect 110 707 116 708
rect 1238 712 1244 713
rect 1238 708 1239 712
rect 1243 708 1244 712
rect 1280 709 1282 741
rect 1304 732 1306 741
rect 1344 732 1346 741
rect 1408 732 1410 741
rect 1488 732 1490 741
rect 1576 732 1578 741
rect 1664 732 1666 741
rect 1752 732 1754 741
rect 1832 732 1834 741
rect 1912 732 1914 741
rect 1992 732 1994 741
rect 2080 732 2082 741
rect 2176 732 2178 741
rect 2280 732 2282 741
rect 2360 732 2362 741
rect 1302 731 1308 732
rect 1302 727 1303 731
rect 1307 727 1308 731
rect 1302 726 1308 727
rect 1342 731 1348 732
rect 1342 727 1343 731
rect 1347 727 1348 731
rect 1342 726 1348 727
rect 1406 731 1412 732
rect 1406 727 1407 731
rect 1411 727 1412 731
rect 1406 726 1412 727
rect 1486 731 1492 732
rect 1486 727 1487 731
rect 1491 727 1492 731
rect 1486 726 1492 727
rect 1574 731 1580 732
rect 1574 727 1575 731
rect 1579 727 1580 731
rect 1574 726 1580 727
rect 1662 731 1668 732
rect 1662 727 1663 731
rect 1667 727 1668 731
rect 1662 726 1668 727
rect 1750 731 1756 732
rect 1750 727 1751 731
rect 1755 727 1756 731
rect 1750 726 1756 727
rect 1830 731 1836 732
rect 1830 727 1831 731
rect 1835 727 1836 731
rect 1830 726 1836 727
rect 1910 731 1916 732
rect 1910 727 1911 731
rect 1915 727 1916 731
rect 1910 726 1916 727
rect 1990 731 1996 732
rect 1990 727 1991 731
rect 1995 727 1996 731
rect 1990 726 1996 727
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 727 2084 731
rect 2078 726 2084 727
rect 2174 731 2180 732
rect 2174 727 2175 731
rect 2179 727 2180 731
rect 2174 726 2180 727
rect 2278 731 2284 732
rect 2278 727 2279 731
rect 2283 727 2284 731
rect 2278 726 2284 727
rect 2358 731 2364 732
rect 2358 727 2359 731
rect 2363 727 2364 731
rect 2358 726 2364 727
rect 2408 709 2410 741
rect 1238 707 1244 708
rect 1278 708 1284 709
rect 1278 704 1279 708
rect 1283 704 1284 708
rect 1278 703 1284 704
rect 2406 708 2412 709
rect 2406 704 2407 708
rect 2411 704 2412 708
rect 2406 703 2412 704
rect 110 695 116 696
rect 110 691 111 695
rect 115 691 116 695
rect 110 690 116 691
rect 1238 695 1244 696
rect 1238 691 1239 695
rect 1243 691 1244 695
rect 1238 690 1244 691
rect 1278 691 1284 692
rect 112 679 114 690
rect 134 688 140 689
rect 134 684 135 688
rect 139 684 140 688
rect 134 683 140 684
rect 190 688 196 689
rect 190 684 191 688
rect 195 684 196 688
rect 190 683 196 684
rect 262 688 268 689
rect 262 684 263 688
rect 267 684 268 688
rect 262 683 268 684
rect 334 688 340 689
rect 334 684 335 688
rect 339 684 340 688
rect 334 683 340 684
rect 398 688 404 689
rect 398 684 399 688
rect 403 684 404 688
rect 398 683 404 684
rect 454 688 460 689
rect 454 684 455 688
rect 459 684 460 688
rect 454 683 460 684
rect 502 688 508 689
rect 502 684 503 688
rect 507 684 508 688
rect 502 683 508 684
rect 542 688 548 689
rect 542 684 543 688
rect 547 684 548 688
rect 542 683 548 684
rect 582 688 588 689
rect 582 684 583 688
rect 587 684 588 688
rect 582 683 588 684
rect 622 688 628 689
rect 622 684 623 688
rect 627 684 628 688
rect 622 683 628 684
rect 670 688 676 689
rect 670 684 671 688
rect 675 684 676 688
rect 670 683 676 684
rect 718 688 724 689
rect 718 684 719 688
rect 723 684 724 688
rect 718 683 724 684
rect 766 688 772 689
rect 766 684 767 688
rect 771 684 772 688
rect 766 683 772 684
rect 814 688 820 689
rect 814 684 815 688
rect 819 684 820 688
rect 814 683 820 684
rect 862 688 868 689
rect 862 684 863 688
rect 867 684 868 688
rect 862 683 868 684
rect 910 688 916 689
rect 910 684 911 688
rect 915 684 916 688
rect 910 683 916 684
rect 136 679 138 683
rect 192 679 194 683
rect 264 679 266 683
rect 336 679 338 683
rect 400 679 402 683
rect 456 679 458 683
rect 504 679 506 683
rect 544 679 546 683
rect 584 679 586 683
rect 624 679 626 683
rect 672 679 674 683
rect 720 679 722 683
rect 768 679 770 683
rect 816 679 818 683
rect 864 679 866 683
rect 912 679 914 683
rect 1240 679 1242 690
rect 1278 687 1279 691
rect 1283 687 1284 691
rect 1278 686 1284 687
rect 2406 691 2412 692
rect 2406 687 2407 691
rect 2411 687 2412 691
rect 2406 686 2412 687
rect 111 678 115 679
rect 111 673 115 674
rect 135 678 139 679
rect 135 673 139 674
rect 191 678 195 679
rect 191 673 195 674
rect 199 678 203 679
rect 199 673 203 674
rect 263 678 267 679
rect 263 673 267 674
rect 279 678 283 679
rect 279 673 283 674
rect 335 678 339 679
rect 335 673 339 674
rect 351 678 355 679
rect 351 673 355 674
rect 399 678 403 679
rect 399 673 403 674
rect 415 678 419 679
rect 415 673 419 674
rect 455 678 459 679
rect 455 673 459 674
rect 487 678 491 679
rect 487 673 491 674
rect 503 678 507 679
rect 503 673 507 674
rect 543 678 547 679
rect 543 673 547 674
rect 559 678 563 679
rect 559 673 563 674
rect 583 678 587 679
rect 583 673 587 674
rect 623 678 627 679
rect 623 673 627 674
rect 639 678 643 679
rect 639 673 643 674
rect 671 678 675 679
rect 671 673 675 674
rect 711 678 715 679
rect 711 673 715 674
rect 719 678 723 679
rect 719 673 723 674
rect 767 678 771 679
rect 767 673 771 674
rect 783 678 787 679
rect 783 673 787 674
rect 815 678 819 679
rect 815 673 819 674
rect 855 678 859 679
rect 855 673 859 674
rect 863 678 867 679
rect 863 673 867 674
rect 911 678 915 679
rect 911 673 915 674
rect 919 678 923 679
rect 919 673 923 674
rect 983 678 987 679
rect 983 673 987 674
rect 1039 678 1043 679
rect 1039 673 1043 674
rect 1095 678 1099 679
rect 1095 673 1099 674
rect 1151 678 1155 679
rect 1151 673 1155 674
rect 1191 678 1195 679
rect 1191 673 1195 674
rect 1239 678 1243 679
rect 1280 675 1282 686
rect 1302 684 1308 685
rect 1302 680 1303 684
rect 1307 680 1308 684
rect 1302 679 1308 680
rect 1342 684 1348 685
rect 1342 680 1343 684
rect 1347 680 1348 684
rect 1342 679 1348 680
rect 1406 684 1412 685
rect 1406 680 1407 684
rect 1411 680 1412 684
rect 1406 679 1412 680
rect 1486 684 1492 685
rect 1486 680 1487 684
rect 1491 680 1492 684
rect 1486 679 1492 680
rect 1574 684 1580 685
rect 1574 680 1575 684
rect 1579 680 1580 684
rect 1574 679 1580 680
rect 1662 684 1668 685
rect 1662 680 1663 684
rect 1667 680 1668 684
rect 1662 679 1668 680
rect 1750 684 1756 685
rect 1750 680 1751 684
rect 1755 680 1756 684
rect 1750 679 1756 680
rect 1830 684 1836 685
rect 1830 680 1831 684
rect 1835 680 1836 684
rect 1830 679 1836 680
rect 1910 684 1916 685
rect 1910 680 1911 684
rect 1915 680 1916 684
rect 1910 679 1916 680
rect 1990 684 1996 685
rect 1990 680 1991 684
rect 1995 680 1996 684
rect 1990 679 1996 680
rect 2078 684 2084 685
rect 2078 680 2079 684
rect 2083 680 2084 684
rect 2078 679 2084 680
rect 2174 684 2180 685
rect 2174 680 2175 684
rect 2179 680 2180 684
rect 2174 679 2180 680
rect 2278 684 2284 685
rect 2278 680 2279 684
rect 2283 680 2284 684
rect 2278 679 2284 680
rect 2358 684 2364 685
rect 2358 680 2359 684
rect 2363 680 2364 684
rect 2358 679 2364 680
rect 1304 675 1306 679
rect 1344 675 1346 679
rect 1408 675 1410 679
rect 1488 675 1490 679
rect 1576 675 1578 679
rect 1664 675 1666 679
rect 1752 675 1754 679
rect 1832 675 1834 679
rect 1912 675 1914 679
rect 1992 675 1994 679
rect 2080 675 2082 679
rect 2176 675 2178 679
rect 2280 675 2282 679
rect 2360 675 2362 679
rect 2408 675 2410 686
rect 1239 673 1243 674
rect 1279 674 1283 675
rect 112 666 114 673
rect 134 672 140 673
rect 134 668 135 672
rect 139 668 140 672
rect 134 667 140 668
rect 198 672 204 673
rect 198 668 199 672
rect 203 668 204 672
rect 198 667 204 668
rect 278 672 284 673
rect 278 668 279 672
rect 283 668 284 672
rect 278 667 284 668
rect 350 672 356 673
rect 350 668 351 672
rect 355 668 356 672
rect 350 667 356 668
rect 414 672 420 673
rect 414 668 415 672
rect 419 668 420 672
rect 414 667 420 668
rect 486 672 492 673
rect 486 668 487 672
rect 491 668 492 672
rect 486 667 492 668
rect 558 672 564 673
rect 558 668 559 672
rect 563 668 564 672
rect 558 667 564 668
rect 638 672 644 673
rect 638 668 639 672
rect 643 668 644 672
rect 638 667 644 668
rect 710 672 716 673
rect 710 668 711 672
rect 715 668 716 672
rect 710 667 716 668
rect 782 672 788 673
rect 782 668 783 672
rect 787 668 788 672
rect 782 667 788 668
rect 854 672 860 673
rect 854 668 855 672
rect 859 668 860 672
rect 854 667 860 668
rect 918 672 924 673
rect 918 668 919 672
rect 923 668 924 672
rect 918 667 924 668
rect 982 672 988 673
rect 982 668 983 672
rect 987 668 988 672
rect 982 667 988 668
rect 1038 672 1044 673
rect 1038 668 1039 672
rect 1043 668 1044 672
rect 1038 667 1044 668
rect 1094 672 1100 673
rect 1094 668 1095 672
rect 1099 668 1100 672
rect 1094 667 1100 668
rect 1150 672 1156 673
rect 1150 668 1151 672
rect 1155 668 1156 672
rect 1150 667 1156 668
rect 1190 672 1196 673
rect 1190 668 1191 672
rect 1195 668 1196 672
rect 1190 667 1196 668
rect 1240 666 1242 673
rect 1279 669 1283 670
rect 1303 674 1307 675
rect 1303 669 1307 670
rect 1343 674 1347 675
rect 1343 669 1347 670
rect 1399 674 1403 675
rect 1399 669 1403 670
rect 1407 674 1411 675
rect 1407 669 1411 670
rect 1487 674 1491 675
rect 1487 669 1491 670
rect 1511 674 1515 675
rect 1511 669 1515 670
rect 1575 674 1579 675
rect 1575 669 1579 670
rect 1623 674 1627 675
rect 1623 669 1627 670
rect 1663 674 1667 675
rect 1663 669 1667 670
rect 1727 674 1731 675
rect 1727 669 1731 670
rect 1751 674 1755 675
rect 1751 669 1755 670
rect 1815 674 1819 675
rect 1815 669 1819 670
rect 1831 674 1835 675
rect 1831 669 1835 670
rect 1895 674 1899 675
rect 1895 669 1899 670
rect 1911 674 1915 675
rect 1911 669 1915 670
rect 1975 674 1979 675
rect 1975 669 1979 670
rect 1991 674 1995 675
rect 1991 669 1995 670
rect 2047 674 2051 675
rect 2047 669 2051 670
rect 2079 674 2083 675
rect 2079 669 2083 670
rect 2111 674 2115 675
rect 2111 669 2115 670
rect 2175 674 2179 675
rect 2175 669 2179 670
rect 2239 674 2243 675
rect 2239 669 2243 670
rect 2279 674 2283 675
rect 2279 669 2283 670
rect 2311 674 2315 675
rect 2311 669 2315 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2407 674 2411 675
rect 2407 669 2411 670
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 110 660 116 661
rect 1238 665 1244 666
rect 1238 661 1239 665
rect 1243 661 1244 665
rect 1280 662 1282 669
rect 1302 668 1308 669
rect 1302 664 1303 668
rect 1307 664 1308 668
rect 1302 663 1308 664
rect 1398 668 1404 669
rect 1398 664 1399 668
rect 1403 664 1404 668
rect 1398 663 1404 664
rect 1510 668 1516 669
rect 1510 664 1511 668
rect 1515 664 1516 668
rect 1510 663 1516 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1726 668 1732 669
rect 1726 664 1727 668
rect 1731 664 1732 668
rect 1726 663 1732 664
rect 1814 668 1820 669
rect 1814 664 1815 668
rect 1819 664 1820 668
rect 1814 663 1820 664
rect 1894 668 1900 669
rect 1894 664 1895 668
rect 1899 664 1900 668
rect 1894 663 1900 664
rect 1974 668 1980 669
rect 1974 664 1975 668
rect 1979 664 1980 668
rect 1974 663 1980 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2110 668 2116 669
rect 2110 664 2111 668
rect 2115 664 2116 668
rect 2110 663 2116 664
rect 2174 668 2180 669
rect 2174 664 2175 668
rect 2179 664 2180 668
rect 2174 663 2180 664
rect 2238 668 2244 669
rect 2238 664 2239 668
rect 2243 664 2244 668
rect 2238 663 2244 664
rect 2310 668 2316 669
rect 2310 664 2311 668
rect 2315 664 2316 668
rect 2310 663 2316 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 2408 662 2410 669
rect 1238 660 1244 661
rect 1278 661 1284 662
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 110 648 116 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 1238 648 1244 649
rect 1238 644 1239 648
rect 1243 644 1244 648
rect 1238 643 1244 644
rect 1278 644 1284 645
rect 112 603 114 643
rect 134 625 140 626
rect 134 621 135 625
rect 139 621 140 625
rect 134 620 140 621
rect 198 625 204 626
rect 198 621 199 625
rect 203 621 204 625
rect 198 620 204 621
rect 278 625 284 626
rect 278 621 279 625
rect 283 621 284 625
rect 278 620 284 621
rect 350 625 356 626
rect 350 621 351 625
rect 355 621 356 625
rect 350 620 356 621
rect 414 625 420 626
rect 414 621 415 625
rect 419 621 420 625
rect 414 620 420 621
rect 486 625 492 626
rect 486 621 487 625
rect 491 621 492 625
rect 486 620 492 621
rect 558 625 564 626
rect 558 621 559 625
rect 563 621 564 625
rect 558 620 564 621
rect 638 625 644 626
rect 638 621 639 625
rect 643 621 644 625
rect 638 620 644 621
rect 710 625 716 626
rect 710 621 711 625
rect 715 621 716 625
rect 710 620 716 621
rect 782 625 788 626
rect 782 621 783 625
rect 787 621 788 625
rect 782 620 788 621
rect 854 625 860 626
rect 854 621 855 625
rect 859 621 860 625
rect 854 620 860 621
rect 918 625 924 626
rect 918 621 919 625
rect 923 621 924 625
rect 918 620 924 621
rect 982 625 988 626
rect 982 621 983 625
rect 987 621 988 625
rect 982 620 988 621
rect 1038 625 1044 626
rect 1038 621 1039 625
rect 1043 621 1044 625
rect 1038 620 1044 621
rect 1094 625 1100 626
rect 1094 621 1095 625
rect 1099 621 1100 625
rect 1094 620 1100 621
rect 1150 625 1156 626
rect 1150 621 1151 625
rect 1155 621 1156 625
rect 1150 620 1156 621
rect 1190 625 1196 626
rect 1190 621 1191 625
rect 1195 621 1196 625
rect 1190 620 1196 621
rect 136 603 138 620
rect 200 603 202 620
rect 280 603 282 620
rect 352 603 354 620
rect 416 603 418 620
rect 488 603 490 620
rect 560 603 562 620
rect 640 603 642 620
rect 712 603 714 620
rect 784 603 786 620
rect 856 603 858 620
rect 920 603 922 620
rect 984 603 986 620
rect 1040 603 1042 620
rect 1096 603 1098 620
rect 1152 603 1154 620
rect 1192 603 1194 620
rect 1240 603 1242 643
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1278 639 1284 640
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 1280 603 1282 639
rect 1302 621 1308 622
rect 1302 617 1303 621
rect 1307 617 1308 621
rect 1302 616 1308 617
rect 1398 621 1404 622
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1398 616 1404 617
rect 1510 621 1516 622
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1622 621 1628 622
rect 1622 617 1623 621
rect 1627 617 1628 621
rect 1622 616 1628 617
rect 1726 621 1732 622
rect 1726 617 1727 621
rect 1731 617 1732 621
rect 1726 616 1732 617
rect 1814 621 1820 622
rect 1814 617 1815 621
rect 1819 617 1820 621
rect 1814 616 1820 617
rect 1894 621 1900 622
rect 1894 617 1895 621
rect 1899 617 1900 621
rect 1894 616 1900 617
rect 1974 621 1980 622
rect 1974 617 1975 621
rect 1979 617 1980 621
rect 1974 616 1980 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2110 621 2116 622
rect 2110 617 2111 621
rect 2115 617 2116 621
rect 2110 616 2116 617
rect 2174 621 2180 622
rect 2174 617 2175 621
rect 2179 617 2180 621
rect 2174 616 2180 617
rect 2238 621 2244 622
rect 2238 617 2239 621
rect 2243 617 2244 621
rect 2238 616 2244 617
rect 2310 621 2316 622
rect 2310 617 2311 621
rect 2315 617 2316 621
rect 2310 616 2316 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 1304 603 1306 616
rect 1400 603 1402 616
rect 1512 603 1514 616
rect 1624 603 1626 616
rect 1728 603 1730 616
rect 1816 603 1818 616
rect 1896 603 1898 616
rect 1976 603 1978 616
rect 2048 603 2050 616
rect 2112 603 2114 616
rect 2176 603 2178 616
rect 2240 603 2242 616
rect 2312 603 2314 616
rect 2360 603 2362 616
rect 2408 603 2410 639
rect 111 602 115 603
rect 111 597 115 598
rect 135 602 139 603
rect 135 597 139 598
rect 191 602 195 603
rect 191 597 195 598
rect 199 602 203 603
rect 199 597 203 598
rect 271 602 275 603
rect 271 597 275 598
rect 279 602 283 603
rect 279 597 283 598
rect 351 602 355 603
rect 351 597 355 598
rect 359 602 363 603
rect 359 597 363 598
rect 415 602 419 603
rect 415 597 419 598
rect 447 602 451 603
rect 447 597 451 598
rect 487 602 491 603
rect 487 597 491 598
rect 535 602 539 603
rect 535 597 539 598
rect 559 602 563 603
rect 559 597 563 598
rect 623 602 627 603
rect 623 597 627 598
rect 639 602 643 603
rect 639 597 643 598
rect 703 602 707 603
rect 703 597 707 598
rect 711 602 715 603
rect 711 597 715 598
rect 783 602 787 603
rect 783 597 787 598
rect 855 602 859 603
rect 855 597 859 598
rect 919 602 923 603
rect 919 597 923 598
rect 975 602 979 603
rect 975 597 979 598
rect 983 602 987 603
rect 983 597 987 598
rect 1023 602 1027 603
rect 1023 597 1027 598
rect 1039 602 1043 603
rect 1039 597 1043 598
rect 1079 602 1083 603
rect 1079 597 1083 598
rect 1095 602 1099 603
rect 1095 597 1099 598
rect 1135 602 1139 603
rect 1135 597 1139 598
rect 1151 602 1155 603
rect 1151 597 1155 598
rect 1191 602 1195 603
rect 1191 597 1195 598
rect 1239 602 1243 603
rect 1239 597 1243 598
rect 1279 602 1283 603
rect 1279 597 1283 598
rect 1303 602 1307 603
rect 1303 597 1307 598
rect 1399 602 1403 603
rect 1399 597 1403 598
rect 1415 602 1419 603
rect 1415 597 1419 598
rect 1455 602 1459 603
rect 1455 597 1459 598
rect 1495 602 1499 603
rect 1495 597 1499 598
rect 1511 602 1515 603
rect 1511 597 1515 598
rect 1543 602 1547 603
rect 1543 597 1547 598
rect 1599 602 1603 603
rect 1599 597 1603 598
rect 1623 602 1627 603
rect 1623 597 1627 598
rect 1663 602 1667 603
rect 1663 597 1667 598
rect 1727 602 1731 603
rect 1727 597 1731 598
rect 1791 602 1795 603
rect 1791 597 1795 598
rect 1815 602 1819 603
rect 1815 597 1819 598
rect 1847 602 1851 603
rect 1847 597 1851 598
rect 1895 602 1899 603
rect 1895 597 1899 598
rect 1911 602 1915 603
rect 1911 597 1915 598
rect 1975 602 1979 603
rect 1975 597 1979 598
rect 2047 602 2051 603
rect 2047 597 2051 598
rect 2111 602 2115 603
rect 2111 597 2115 598
rect 2119 602 2123 603
rect 2119 597 2123 598
rect 2175 602 2179 603
rect 2175 597 2179 598
rect 2199 602 2203 603
rect 2199 597 2203 598
rect 2239 602 2243 603
rect 2239 597 2243 598
rect 2287 602 2291 603
rect 2287 597 2291 598
rect 2311 602 2315 603
rect 2311 597 2315 598
rect 2359 602 2363 603
rect 2359 597 2363 598
rect 2407 602 2411 603
rect 2407 597 2411 598
rect 112 565 114 597
rect 136 588 138 597
rect 192 588 194 597
rect 272 588 274 597
rect 360 588 362 597
rect 448 588 450 597
rect 536 588 538 597
rect 624 588 626 597
rect 704 588 706 597
rect 784 588 786 597
rect 856 588 858 597
rect 920 588 922 597
rect 976 588 978 597
rect 1024 588 1026 597
rect 1080 588 1082 597
rect 1136 588 1138 597
rect 1192 588 1194 597
rect 134 587 140 588
rect 134 583 135 587
rect 139 583 140 587
rect 134 582 140 583
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 270 587 276 588
rect 270 583 271 587
rect 275 583 276 587
rect 270 582 276 583
rect 358 587 364 588
rect 358 583 359 587
rect 363 583 364 587
rect 358 582 364 583
rect 446 587 452 588
rect 446 583 447 587
rect 451 583 452 587
rect 446 582 452 583
rect 534 587 540 588
rect 534 583 535 587
rect 539 583 540 587
rect 534 582 540 583
rect 622 587 628 588
rect 622 583 623 587
rect 627 583 628 587
rect 622 582 628 583
rect 702 587 708 588
rect 702 583 703 587
rect 707 583 708 587
rect 702 582 708 583
rect 782 587 788 588
rect 782 583 783 587
rect 787 583 788 587
rect 782 582 788 583
rect 854 587 860 588
rect 854 583 855 587
rect 859 583 860 587
rect 854 582 860 583
rect 918 587 924 588
rect 918 583 919 587
rect 923 583 924 587
rect 918 582 924 583
rect 974 587 980 588
rect 974 583 975 587
rect 979 583 980 587
rect 974 582 980 583
rect 1022 587 1028 588
rect 1022 583 1023 587
rect 1027 583 1028 587
rect 1022 582 1028 583
rect 1078 587 1084 588
rect 1078 583 1079 587
rect 1083 583 1084 587
rect 1078 582 1084 583
rect 1134 587 1140 588
rect 1134 583 1135 587
rect 1139 583 1140 587
rect 1134 582 1140 583
rect 1190 587 1196 588
rect 1190 583 1191 587
rect 1195 583 1196 587
rect 1190 582 1196 583
rect 1240 565 1242 597
rect 1280 565 1282 597
rect 1416 588 1418 597
rect 1456 588 1458 597
rect 1496 588 1498 597
rect 1544 588 1546 597
rect 1600 588 1602 597
rect 1664 588 1666 597
rect 1728 588 1730 597
rect 1792 588 1794 597
rect 1848 588 1850 597
rect 1912 588 1914 597
rect 1976 588 1978 597
rect 2048 588 2050 597
rect 2120 588 2122 597
rect 2200 588 2202 597
rect 2288 588 2290 597
rect 2360 588 2362 597
rect 1414 587 1420 588
rect 1414 583 1415 587
rect 1419 583 1420 587
rect 1414 582 1420 583
rect 1454 587 1460 588
rect 1454 583 1455 587
rect 1459 583 1460 587
rect 1454 582 1460 583
rect 1494 587 1500 588
rect 1494 583 1495 587
rect 1499 583 1500 587
rect 1494 582 1500 583
rect 1542 587 1548 588
rect 1542 583 1543 587
rect 1547 583 1548 587
rect 1542 582 1548 583
rect 1598 587 1604 588
rect 1598 583 1599 587
rect 1603 583 1604 587
rect 1598 582 1604 583
rect 1662 587 1668 588
rect 1662 583 1663 587
rect 1667 583 1668 587
rect 1662 582 1668 583
rect 1726 587 1732 588
rect 1726 583 1727 587
rect 1731 583 1732 587
rect 1726 582 1732 583
rect 1790 587 1796 588
rect 1790 583 1791 587
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1846 587 1852 588
rect 1846 583 1847 587
rect 1851 583 1852 587
rect 1846 582 1852 583
rect 1910 587 1916 588
rect 1910 583 1911 587
rect 1915 583 1916 587
rect 1910 582 1916 583
rect 1974 587 1980 588
rect 1974 583 1975 587
rect 1979 583 1980 587
rect 1974 582 1980 583
rect 2046 587 2052 588
rect 2046 583 2047 587
rect 2051 583 2052 587
rect 2046 582 2052 583
rect 2118 587 2124 588
rect 2118 583 2119 587
rect 2123 583 2124 587
rect 2118 582 2124 583
rect 2198 587 2204 588
rect 2198 583 2199 587
rect 2203 583 2204 587
rect 2198 582 2204 583
rect 2286 587 2292 588
rect 2286 583 2287 587
rect 2291 583 2292 587
rect 2286 582 2292 583
rect 2358 587 2364 588
rect 2358 583 2359 587
rect 2363 583 2364 587
rect 2358 582 2364 583
rect 2408 565 2410 597
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 110 559 116 560
rect 1238 564 1244 565
rect 1238 560 1239 564
rect 1243 560 1244 564
rect 1238 559 1244 560
rect 1278 564 1284 565
rect 1278 560 1279 564
rect 1283 560 1284 564
rect 1278 559 1284 560
rect 2406 564 2412 565
rect 2406 560 2407 564
rect 2411 560 2412 564
rect 2406 559 2412 560
rect 110 547 116 548
rect 110 543 111 547
rect 115 543 116 547
rect 110 542 116 543
rect 1238 547 1244 548
rect 1238 543 1239 547
rect 1243 543 1244 547
rect 1238 542 1244 543
rect 1278 547 1284 548
rect 1278 543 1279 547
rect 1283 543 1284 547
rect 1278 542 1284 543
rect 2406 547 2412 548
rect 2406 543 2407 547
rect 2411 543 2412 547
rect 2406 542 2412 543
rect 112 527 114 542
rect 134 540 140 541
rect 134 536 135 540
rect 139 536 140 540
rect 134 535 140 536
rect 190 540 196 541
rect 190 536 191 540
rect 195 536 196 540
rect 190 535 196 536
rect 270 540 276 541
rect 270 536 271 540
rect 275 536 276 540
rect 270 535 276 536
rect 358 540 364 541
rect 358 536 359 540
rect 363 536 364 540
rect 358 535 364 536
rect 446 540 452 541
rect 446 536 447 540
rect 451 536 452 540
rect 446 535 452 536
rect 534 540 540 541
rect 534 536 535 540
rect 539 536 540 540
rect 534 535 540 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 702 540 708 541
rect 702 536 703 540
rect 707 536 708 540
rect 702 535 708 536
rect 782 540 788 541
rect 782 536 783 540
rect 787 536 788 540
rect 782 535 788 536
rect 854 540 860 541
rect 854 536 855 540
rect 859 536 860 540
rect 854 535 860 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 974 540 980 541
rect 974 536 975 540
rect 979 536 980 540
rect 974 535 980 536
rect 1022 540 1028 541
rect 1022 536 1023 540
rect 1027 536 1028 540
rect 1022 535 1028 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 1134 540 1140 541
rect 1134 536 1135 540
rect 1139 536 1140 540
rect 1134 535 1140 536
rect 1190 540 1196 541
rect 1190 536 1191 540
rect 1195 536 1196 540
rect 1190 535 1196 536
rect 136 527 138 535
rect 192 527 194 535
rect 272 527 274 535
rect 360 527 362 535
rect 448 527 450 535
rect 536 527 538 535
rect 624 527 626 535
rect 704 527 706 535
rect 784 527 786 535
rect 856 527 858 535
rect 920 527 922 535
rect 976 527 978 535
rect 1024 527 1026 535
rect 1080 527 1082 535
rect 1136 527 1138 535
rect 1192 527 1194 535
rect 1240 527 1242 542
rect 1280 535 1282 542
rect 1414 540 1420 541
rect 1414 536 1415 540
rect 1419 536 1420 540
rect 1414 535 1420 536
rect 1454 540 1460 541
rect 1454 536 1455 540
rect 1459 536 1460 540
rect 1454 535 1460 536
rect 1494 540 1500 541
rect 1494 536 1495 540
rect 1499 536 1500 540
rect 1494 535 1500 536
rect 1542 540 1548 541
rect 1542 536 1543 540
rect 1547 536 1548 540
rect 1542 535 1548 536
rect 1598 540 1604 541
rect 1598 536 1599 540
rect 1603 536 1604 540
rect 1598 535 1604 536
rect 1662 540 1668 541
rect 1662 536 1663 540
rect 1667 536 1668 540
rect 1662 535 1668 536
rect 1726 540 1732 541
rect 1726 536 1727 540
rect 1731 536 1732 540
rect 1726 535 1732 536
rect 1790 540 1796 541
rect 1790 536 1791 540
rect 1795 536 1796 540
rect 1790 535 1796 536
rect 1846 540 1852 541
rect 1846 536 1847 540
rect 1851 536 1852 540
rect 1846 535 1852 536
rect 1910 540 1916 541
rect 1910 536 1911 540
rect 1915 536 1916 540
rect 1910 535 1916 536
rect 1974 540 1980 541
rect 1974 536 1975 540
rect 1979 536 1980 540
rect 1974 535 1980 536
rect 2046 540 2052 541
rect 2046 536 2047 540
rect 2051 536 2052 540
rect 2046 535 2052 536
rect 2118 540 2124 541
rect 2118 536 2119 540
rect 2123 536 2124 540
rect 2118 535 2124 536
rect 2198 540 2204 541
rect 2198 536 2199 540
rect 2203 536 2204 540
rect 2198 535 2204 536
rect 2286 540 2292 541
rect 2286 536 2287 540
rect 2291 536 2292 540
rect 2286 535 2292 536
rect 2358 540 2364 541
rect 2358 536 2359 540
rect 2363 536 2364 540
rect 2358 535 2364 536
rect 2408 535 2410 542
rect 1279 534 1283 535
rect 1279 529 1283 530
rect 1303 534 1307 535
rect 1303 529 1307 530
rect 1375 534 1379 535
rect 1375 529 1379 530
rect 1415 534 1419 535
rect 1415 529 1419 530
rect 1455 534 1459 535
rect 1455 529 1459 530
rect 1479 534 1483 535
rect 1479 529 1483 530
rect 1495 534 1499 535
rect 1495 529 1499 530
rect 1543 534 1547 535
rect 1543 529 1547 530
rect 1583 534 1587 535
rect 1583 529 1587 530
rect 1599 534 1603 535
rect 1599 529 1603 530
rect 1663 534 1667 535
rect 1663 529 1667 530
rect 1695 534 1699 535
rect 1695 529 1699 530
rect 1727 534 1731 535
rect 1727 529 1731 530
rect 1791 534 1795 535
rect 1791 529 1795 530
rect 1799 534 1803 535
rect 1799 529 1803 530
rect 1847 534 1851 535
rect 1847 529 1851 530
rect 1903 534 1907 535
rect 1903 529 1907 530
rect 1911 534 1915 535
rect 1911 529 1915 530
rect 1975 534 1979 535
rect 1975 529 1979 530
rect 2007 534 2011 535
rect 2007 529 2011 530
rect 2047 534 2051 535
rect 2047 529 2051 530
rect 2103 534 2107 535
rect 2103 529 2107 530
rect 2119 534 2123 535
rect 2119 529 2123 530
rect 2191 534 2195 535
rect 2191 529 2195 530
rect 2199 534 2203 535
rect 2199 529 2203 530
rect 2287 534 2291 535
rect 2287 529 2291 530
rect 2359 534 2363 535
rect 2359 529 2363 530
rect 2407 534 2411 535
rect 2407 529 2411 530
rect 111 526 115 527
rect 111 521 115 522
rect 135 526 139 527
rect 135 521 139 522
rect 191 526 195 527
rect 191 521 195 522
rect 263 526 267 527
rect 263 521 267 522
rect 271 526 275 527
rect 271 521 275 522
rect 335 526 339 527
rect 335 521 339 522
rect 359 526 363 527
rect 359 521 363 522
rect 415 526 419 527
rect 415 521 419 522
rect 447 526 451 527
rect 447 521 451 522
rect 495 526 499 527
rect 495 521 499 522
rect 535 526 539 527
rect 535 521 539 522
rect 575 526 579 527
rect 575 521 579 522
rect 623 526 627 527
rect 623 521 627 522
rect 647 526 651 527
rect 647 521 651 522
rect 703 526 707 527
rect 703 521 707 522
rect 719 526 723 527
rect 719 521 723 522
rect 783 526 787 527
rect 783 521 787 522
rect 847 526 851 527
rect 847 521 851 522
rect 855 526 859 527
rect 855 521 859 522
rect 903 526 907 527
rect 903 521 907 522
rect 919 526 923 527
rect 919 521 923 522
rect 959 526 963 527
rect 959 521 963 522
rect 975 526 979 527
rect 975 521 979 522
rect 1023 526 1027 527
rect 1023 521 1027 522
rect 1079 526 1083 527
rect 1079 521 1083 522
rect 1087 526 1091 527
rect 1087 521 1091 522
rect 1135 526 1139 527
rect 1135 521 1139 522
rect 1151 526 1155 527
rect 1151 521 1155 522
rect 1191 526 1195 527
rect 1191 521 1195 522
rect 1239 526 1243 527
rect 1280 522 1282 529
rect 1302 528 1308 529
rect 1302 524 1303 528
rect 1307 524 1308 528
rect 1302 523 1308 524
rect 1374 528 1380 529
rect 1374 524 1375 528
rect 1379 524 1380 528
rect 1374 523 1380 524
rect 1478 528 1484 529
rect 1478 524 1479 528
rect 1483 524 1484 528
rect 1478 523 1484 524
rect 1582 528 1588 529
rect 1582 524 1583 528
rect 1587 524 1588 528
rect 1582 523 1588 524
rect 1694 528 1700 529
rect 1694 524 1695 528
rect 1699 524 1700 528
rect 1694 523 1700 524
rect 1798 528 1804 529
rect 1798 524 1799 528
rect 1803 524 1804 528
rect 1798 523 1804 524
rect 1902 528 1908 529
rect 1902 524 1903 528
rect 1907 524 1908 528
rect 1902 523 1908 524
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 2006 523 2012 524
rect 2102 528 2108 529
rect 2102 524 2103 528
rect 2107 524 2108 528
rect 2102 523 2108 524
rect 2190 528 2196 529
rect 2190 524 2191 528
rect 2195 524 2196 528
rect 2190 523 2196 524
rect 2286 528 2292 529
rect 2286 524 2287 528
rect 2291 524 2292 528
rect 2286 523 2292 524
rect 2358 528 2364 529
rect 2358 524 2359 528
rect 2363 524 2364 528
rect 2358 523 2364 524
rect 2408 522 2410 529
rect 1239 521 1243 522
rect 1278 521 1284 522
rect 112 514 114 521
rect 134 520 140 521
rect 134 516 135 520
rect 139 516 140 520
rect 134 515 140 516
rect 190 520 196 521
rect 190 516 191 520
rect 195 516 196 520
rect 190 515 196 516
rect 262 520 268 521
rect 262 516 263 520
rect 267 516 268 520
rect 262 515 268 516
rect 334 520 340 521
rect 334 516 335 520
rect 339 516 340 520
rect 334 515 340 516
rect 414 520 420 521
rect 414 516 415 520
rect 419 516 420 520
rect 414 515 420 516
rect 494 520 500 521
rect 494 516 495 520
rect 499 516 500 520
rect 494 515 500 516
rect 574 520 580 521
rect 574 516 575 520
rect 579 516 580 520
rect 574 515 580 516
rect 646 520 652 521
rect 646 516 647 520
rect 651 516 652 520
rect 646 515 652 516
rect 718 520 724 521
rect 718 516 719 520
rect 723 516 724 520
rect 718 515 724 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 846 520 852 521
rect 846 516 847 520
rect 851 516 852 520
rect 846 515 852 516
rect 902 520 908 521
rect 902 516 903 520
rect 907 516 908 520
rect 902 515 908 516
rect 958 520 964 521
rect 958 516 959 520
rect 963 516 964 520
rect 958 515 964 516
rect 1022 520 1028 521
rect 1022 516 1023 520
rect 1027 516 1028 520
rect 1022 515 1028 516
rect 1086 520 1092 521
rect 1086 516 1087 520
rect 1091 516 1092 520
rect 1086 515 1092 516
rect 1150 520 1156 521
rect 1150 516 1151 520
rect 1155 516 1156 520
rect 1150 515 1156 516
rect 1190 520 1196 521
rect 1190 516 1191 520
rect 1195 516 1196 520
rect 1190 515 1196 516
rect 1240 514 1242 521
rect 1278 517 1279 521
rect 1283 517 1284 521
rect 1278 516 1284 517
rect 2406 521 2412 522
rect 2406 517 2407 521
rect 2411 517 2412 521
rect 2406 516 2412 517
rect 110 513 116 514
rect 110 509 111 513
rect 115 509 116 513
rect 110 508 116 509
rect 1238 513 1244 514
rect 1238 509 1239 513
rect 1243 509 1244 513
rect 1238 508 1244 509
rect 1278 504 1284 505
rect 1278 500 1279 504
rect 1283 500 1284 504
rect 1278 499 1284 500
rect 2406 504 2412 505
rect 2406 500 2407 504
rect 2411 500 2412 504
rect 2406 499 2412 500
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 110 491 116 492
rect 1238 496 1244 497
rect 1238 492 1239 496
rect 1243 492 1244 496
rect 1238 491 1244 492
rect 112 459 114 491
rect 134 473 140 474
rect 134 469 135 473
rect 139 469 140 473
rect 134 468 140 469
rect 190 473 196 474
rect 190 469 191 473
rect 195 469 196 473
rect 190 468 196 469
rect 262 473 268 474
rect 262 469 263 473
rect 267 469 268 473
rect 262 468 268 469
rect 334 473 340 474
rect 334 469 335 473
rect 339 469 340 473
rect 334 468 340 469
rect 414 473 420 474
rect 414 469 415 473
rect 419 469 420 473
rect 414 468 420 469
rect 494 473 500 474
rect 494 469 495 473
rect 499 469 500 473
rect 494 468 500 469
rect 574 473 580 474
rect 574 469 575 473
rect 579 469 580 473
rect 574 468 580 469
rect 646 473 652 474
rect 646 469 647 473
rect 651 469 652 473
rect 646 468 652 469
rect 718 473 724 474
rect 718 469 719 473
rect 723 469 724 473
rect 718 468 724 469
rect 782 473 788 474
rect 782 469 783 473
rect 787 469 788 473
rect 782 468 788 469
rect 846 473 852 474
rect 846 469 847 473
rect 851 469 852 473
rect 846 468 852 469
rect 902 473 908 474
rect 902 469 903 473
rect 907 469 908 473
rect 902 468 908 469
rect 958 473 964 474
rect 958 469 959 473
rect 963 469 964 473
rect 958 468 964 469
rect 1022 473 1028 474
rect 1022 469 1023 473
rect 1027 469 1028 473
rect 1022 468 1028 469
rect 1086 473 1092 474
rect 1086 469 1087 473
rect 1091 469 1092 473
rect 1086 468 1092 469
rect 1150 473 1156 474
rect 1150 469 1151 473
rect 1155 469 1156 473
rect 1150 468 1156 469
rect 1190 473 1196 474
rect 1190 469 1191 473
rect 1195 469 1196 473
rect 1190 468 1196 469
rect 136 459 138 468
rect 192 459 194 468
rect 264 459 266 468
rect 336 459 338 468
rect 416 459 418 468
rect 496 459 498 468
rect 576 459 578 468
rect 648 459 650 468
rect 720 459 722 468
rect 784 459 786 468
rect 848 459 850 468
rect 904 459 906 468
rect 960 459 962 468
rect 1024 459 1026 468
rect 1088 459 1090 468
rect 1152 459 1154 468
rect 1192 459 1194 468
rect 1240 459 1242 491
rect 1280 463 1282 499
rect 1302 481 1308 482
rect 1302 477 1303 481
rect 1307 477 1308 481
rect 1302 476 1308 477
rect 1374 481 1380 482
rect 1374 477 1375 481
rect 1379 477 1380 481
rect 1374 476 1380 477
rect 1478 481 1484 482
rect 1478 477 1479 481
rect 1483 477 1484 481
rect 1478 476 1484 477
rect 1582 481 1588 482
rect 1582 477 1583 481
rect 1587 477 1588 481
rect 1582 476 1588 477
rect 1694 481 1700 482
rect 1694 477 1695 481
rect 1699 477 1700 481
rect 1694 476 1700 477
rect 1798 481 1804 482
rect 1798 477 1799 481
rect 1803 477 1804 481
rect 1798 476 1804 477
rect 1902 481 1908 482
rect 1902 477 1903 481
rect 1907 477 1908 481
rect 1902 476 1908 477
rect 2006 481 2012 482
rect 2006 477 2007 481
rect 2011 477 2012 481
rect 2006 476 2012 477
rect 2102 481 2108 482
rect 2102 477 2103 481
rect 2107 477 2108 481
rect 2102 476 2108 477
rect 2190 481 2196 482
rect 2190 477 2191 481
rect 2195 477 2196 481
rect 2190 476 2196 477
rect 2286 481 2292 482
rect 2286 477 2287 481
rect 2291 477 2292 481
rect 2286 476 2292 477
rect 2358 481 2364 482
rect 2358 477 2359 481
rect 2363 477 2364 481
rect 2358 476 2364 477
rect 1304 463 1306 476
rect 1376 463 1378 476
rect 1480 463 1482 476
rect 1584 463 1586 476
rect 1696 463 1698 476
rect 1800 463 1802 476
rect 1904 463 1906 476
rect 2008 463 2010 476
rect 2104 463 2106 476
rect 2192 463 2194 476
rect 2288 463 2290 476
rect 2360 463 2362 476
rect 2408 463 2410 499
rect 1279 462 1283 463
rect 111 458 115 459
rect 111 453 115 454
rect 135 458 139 459
rect 135 453 139 454
rect 183 458 187 459
rect 183 453 187 454
rect 191 458 195 459
rect 191 453 195 454
rect 223 458 227 459
rect 223 453 227 454
rect 263 458 267 459
rect 263 453 267 454
rect 311 458 315 459
rect 311 453 315 454
rect 335 458 339 459
rect 335 453 339 454
rect 367 458 371 459
rect 367 453 371 454
rect 415 458 419 459
rect 415 453 419 454
rect 431 458 435 459
rect 431 453 435 454
rect 495 458 499 459
rect 495 453 499 454
rect 559 458 563 459
rect 559 453 563 454
rect 575 458 579 459
rect 575 453 579 454
rect 615 458 619 459
rect 615 453 619 454
rect 647 458 651 459
rect 647 453 651 454
rect 671 458 675 459
rect 671 453 675 454
rect 719 458 723 459
rect 719 453 723 454
rect 775 458 779 459
rect 775 453 779 454
rect 783 458 787 459
rect 783 453 787 454
rect 831 458 835 459
rect 831 453 835 454
rect 847 458 851 459
rect 847 453 851 454
rect 887 458 891 459
rect 887 453 891 454
rect 903 458 907 459
rect 903 453 907 454
rect 959 458 963 459
rect 959 453 963 454
rect 1023 458 1027 459
rect 1023 453 1027 454
rect 1087 458 1091 459
rect 1087 453 1091 454
rect 1151 458 1155 459
rect 1151 453 1155 454
rect 1191 458 1195 459
rect 1191 453 1195 454
rect 1239 458 1243 459
rect 1279 457 1283 458
rect 1303 462 1307 463
rect 1303 457 1307 458
rect 1343 462 1347 463
rect 1343 457 1347 458
rect 1375 462 1379 463
rect 1375 457 1379 458
rect 1399 462 1403 463
rect 1399 457 1403 458
rect 1463 462 1467 463
rect 1463 457 1467 458
rect 1479 462 1483 463
rect 1479 457 1483 458
rect 1527 462 1531 463
rect 1527 457 1531 458
rect 1583 462 1587 463
rect 1583 457 1587 458
rect 1591 462 1595 463
rect 1591 457 1595 458
rect 1663 462 1667 463
rect 1663 457 1667 458
rect 1695 462 1699 463
rect 1695 457 1699 458
rect 1735 462 1739 463
rect 1735 457 1739 458
rect 1799 462 1803 463
rect 1799 457 1803 458
rect 1815 462 1819 463
rect 1815 457 1819 458
rect 1895 462 1899 463
rect 1895 457 1899 458
rect 1903 462 1907 463
rect 1903 457 1907 458
rect 1975 462 1979 463
rect 1975 457 1979 458
rect 2007 462 2011 463
rect 2007 457 2011 458
rect 2055 462 2059 463
rect 2055 457 2059 458
rect 2103 462 2107 463
rect 2103 457 2107 458
rect 2135 462 2139 463
rect 2135 457 2139 458
rect 2191 462 2195 463
rect 2191 457 2195 458
rect 2215 462 2219 463
rect 2215 457 2219 458
rect 2287 462 2291 463
rect 2287 457 2291 458
rect 2295 462 2299 463
rect 2295 457 2299 458
rect 2359 462 2363 463
rect 2359 457 2363 458
rect 2407 462 2411 463
rect 2407 457 2411 458
rect 1239 453 1243 454
rect 112 421 114 453
rect 184 444 186 453
rect 224 444 226 453
rect 264 444 266 453
rect 312 444 314 453
rect 368 444 370 453
rect 432 444 434 453
rect 496 444 498 453
rect 560 444 562 453
rect 616 444 618 453
rect 672 444 674 453
rect 720 444 722 453
rect 776 444 778 453
rect 832 444 834 453
rect 888 444 890 453
rect 182 443 188 444
rect 182 439 183 443
rect 187 439 188 443
rect 182 438 188 439
rect 222 443 228 444
rect 222 439 223 443
rect 227 439 228 443
rect 222 438 228 439
rect 262 443 268 444
rect 262 439 263 443
rect 267 439 268 443
rect 262 438 268 439
rect 310 443 316 444
rect 310 439 311 443
rect 315 439 316 443
rect 310 438 316 439
rect 366 443 372 444
rect 366 439 367 443
rect 371 439 372 443
rect 366 438 372 439
rect 430 443 436 444
rect 430 439 431 443
rect 435 439 436 443
rect 430 438 436 439
rect 494 443 500 444
rect 494 439 495 443
rect 499 439 500 443
rect 494 438 500 439
rect 558 443 564 444
rect 558 439 559 443
rect 563 439 564 443
rect 558 438 564 439
rect 614 443 620 444
rect 614 439 615 443
rect 619 439 620 443
rect 614 438 620 439
rect 670 443 676 444
rect 670 439 671 443
rect 675 439 676 443
rect 670 438 676 439
rect 718 443 724 444
rect 718 439 719 443
rect 723 439 724 443
rect 718 438 724 439
rect 774 443 780 444
rect 774 439 775 443
rect 779 439 780 443
rect 774 438 780 439
rect 830 443 836 444
rect 830 439 831 443
rect 835 439 836 443
rect 830 438 836 439
rect 886 443 892 444
rect 886 439 887 443
rect 891 439 892 443
rect 886 438 892 439
rect 1240 421 1242 453
rect 1280 425 1282 457
rect 1304 448 1306 457
rect 1344 448 1346 457
rect 1400 448 1402 457
rect 1464 448 1466 457
rect 1528 448 1530 457
rect 1592 448 1594 457
rect 1664 448 1666 457
rect 1736 448 1738 457
rect 1816 448 1818 457
rect 1896 448 1898 457
rect 1976 448 1978 457
rect 2056 448 2058 457
rect 2136 448 2138 457
rect 2216 448 2218 457
rect 2296 448 2298 457
rect 2360 448 2362 457
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1398 447 1404 448
rect 1398 443 1399 447
rect 1403 443 1404 447
rect 1398 442 1404 443
rect 1462 447 1468 448
rect 1462 443 1463 447
rect 1467 443 1468 447
rect 1462 442 1468 443
rect 1526 447 1532 448
rect 1526 443 1527 447
rect 1531 443 1532 447
rect 1526 442 1532 443
rect 1590 447 1596 448
rect 1590 443 1591 447
rect 1595 443 1596 447
rect 1590 442 1596 443
rect 1662 447 1668 448
rect 1662 443 1663 447
rect 1667 443 1668 447
rect 1662 442 1668 443
rect 1734 447 1740 448
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1734 442 1740 443
rect 1814 447 1820 448
rect 1814 443 1815 447
rect 1819 443 1820 447
rect 1814 442 1820 443
rect 1894 447 1900 448
rect 1894 443 1895 447
rect 1899 443 1900 447
rect 1894 442 1900 443
rect 1974 447 1980 448
rect 1974 443 1975 447
rect 1979 443 1980 447
rect 1974 442 1980 443
rect 2054 447 2060 448
rect 2054 443 2055 447
rect 2059 443 2060 447
rect 2054 442 2060 443
rect 2134 447 2140 448
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2134 442 2140 443
rect 2214 447 2220 448
rect 2214 443 2215 447
rect 2219 443 2220 447
rect 2214 442 2220 443
rect 2294 447 2300 448
rect 2294 443 2295 447
rect 2299 443 2300 447
rect 2294 442 2300 443
rect 2358 447 2364 448
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2358 442 2364 443
rect 2408 425 2410 457
rect 1278 424 1284 425
rect 110 420 116 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 1238 420 1244 421
rect 1238 416 1239 420
rect 1243 416 1244 420
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1278 419 1284 420
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2406 419 2412 420
rect 1238 415 1244 416
rect 1278 407 1284 408
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 110 398 116 399
rect 1238 403 1244 404
rect 1238 399 1239 403
rect 1243 399 1244 403
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1278 402 1284 403
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 1238 398 1244 399
rect 112 391 114 398
rect 182 396 188 397
rect 182 392 183 396
rect 187 392 188 396
rect 182 391 188 392
rect 222 396 228 397
rect 222 392 223 396
rect 227 392 228 396
rect 222 391 228 392
rect 262 396 268 397
rect 262 392 263 396
rect 267 392 268 396
rect 262 391 268 392
rect 310 396 316 397
rect 310 392 311 396
rect 315 392 316 396
rect 310 391 316 392
rect 366 396 372 397
rect 366 392 367 396
rect 371 392 372 396
rect 366 391 372 392
rect 430 396 436 397
rect 430 392 431 396
rect 435 392 436 396
rect 430 391 436 392
rect 494 396 500 397
rect 494 392 495 396
rect 499 392 500 396
rect 494 391 500 392
rect 558 396 564 397
rect 558 392 559 396
rect 563 392 564 396
rect 558 391 564 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 718 396 724 397
rect 718 392 719 396
rect 723 392 724 396
rect 718 391 724 392
rect 774 396 780 397
rect 774 392 775 396
rect 779 392 780 396
rect 774 391 780 392
rect 830 396 836 397
rect 830 392 831 396
rect 835 392 836 396
rect 830 391 836 392
rect 886 396 892 397
rect 886 392 887 396
rect 891 392 892 396
rect 886 391 892 392
rect 1240 391 1242 398
rect 1280 391 1282 402
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1398 400 1404 401
rect 1398 396 1399 400
rect 1403 396 1404 400
rect 1398 395 1404 396
rect 1462 400 1468 401
rect 1462 396 1463 400
rect 1467 396 1468 400
rect 1462 395 1468 396
rect 1526 400 1532 401
rect 1526 396 1527 400
rect 1531 396 1532 400
rect 1526 395 1532 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1662 400 1668 401
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1814 400 1820 401
rect 1814 396 1815 400
rect 1819 396 1820 400
rect 1814 395 1820 396
rect 1894 400 1900 401
rect 1894 396 1895 400
rect 1899 396 1900 400
rect 1894 395 1900 396
rect 1974 400 1980 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 2054 400 2060 401
rect 2054 396 2055 400
rect 2059 396 2060 400
rect 2054 395 2060 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2214 400 2220 401
rect 2214 396 2215 400
rect 2219 396 2220 400
rect 2214 395 2220 396
rect 2294 400 2300 401
rect 2294 396 2295 400
rect 2299 396 2300 400
rect 2294 395 2300 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 1304 391 1306 395
rect 1344 391 1346 395
rect 1400 391 1402 395
rect 1464 391 1466 395
rect 1528 391 1530 395
rect 1592 391 1594 395
rect 1664 391 1666 395
rect 1736 391 1738 395
rect 1816 391 1818 395
rect 1896 391 1898 395
rect 1976 391 1978 395
rect 2056 391 2058 395
rect 2136 391 2138 395
rect 2216 391 2218 395
rect 2296 391 2298 395
rect 2360 391 2362 395
rect 2408 391 2410 402
rect 111 390 115 391
rect 111 385 115 386
rect 135 390 139 391
rect 135 385 139 386
rect 175 390 179 391
rect 175 385 179 386
rect 183 390 187 391
rect 183 385 187 386
rect 223 390 227 391
rect 223 385 227 386
rect 231 390 235 391
rect 231 385 235 386
rect 263 390 267 391
rect 263 385 267 386
rect 287 390 291 391
rect 287 385 291 386
rect 311 390 315 391
rect 311 385 315 386
rect 343 390 347 391
rect 343 385 347 386
rect 367 390 371 391
rect 367 385 371 386
rect 391 390 395 391
rect 391 385 395 386
rect 431 390 435 391
rect 431 385 435 386
rect 439 390 443 391
rect 439 385 443 386
rect 487 390 491 391
rect 487 385 491 386
rect 495 390 499 391
rect 495 385 499 386
rect 535 390 539 391
rect 535 385 539 386
rect 559 390 563 391
rect 559 385 563 386
rect 583 390 587 391
rect 583 385 587 386
rect 615 390 619 391
rect 615 385 619 386
rect 631 390 635 391
rect 631 385 635 386
rect 671 390 675 391
rect 671 385 675 386
rect 679 390 683 391
rect 679 385 683 386
rect 719 390 723 391
rect 719 385 723 386
rect 727 390 731 391
rect 727 385 731 386
rect 775 390 779 391
rect 775 385 779 386
rect 831 390 835 391
rect 831 385 835 386
rect 887 390 891 391
rect 887 385 891 386
rect 1239 390 1243 391
rect 1239 385 1243 386
rect 1279 390 1283 391
rect 1279 385 1283 386
rect 1303 390 1307 391
rect 1303 385 1307 386
rect 1343 390 1347 391
rect 1343 385 1347 386
rect 1399 390 1403 391
rect 1399 385 1403 386
rect 1447 390 1451 391
rect 1447 385 1451 386
rect 1463 390 1467 391
rect 1463 385 1467 386
rect 1487 390 1491 391
rect 1487 385 1491 386
rect 1527 390 1531 391
rect 1527 385 1531 386
rect 1535 390 1539 391
rect 1535 385 1539 386
rect 1591 390 1595 391
rect 1591 385 1595 386
rect 1663 390 1667 391
rect 1663 385 1667 386
rect 1735 390 1739 391
rect 1735 385 1739 386
rect 1815 390 1819 391
rect 1815 385 1819 386
rect 1895 390 1899 391
rect 1895 385 1899 386
rect 1967 390 1971 391
rect 1967 385 1971 386
rect 1975 390 1979 391
rect 1975 385 1979 386
rect 2039 390 2043 391
rect 2039 385 2043 386
rect 2055 390 2059 391
rect 2055 385 2059 386
rect 2111 390 2115 391
rect 2111 385 2115 386
rect 2135 390 2139 391
rect 2135 385 2139 386
rect 2175 390 2179 391
rect 2175 385 2179 386
rect 2215 390 2219 391
rect 2215 385 2219 386
rect 2239 390 2243 391
rect 2239 385 2243 386
rect 2295 390 2299 391
rect 2295 385 2299 386
rect 2303 390 2307 391
rect 2303 385 2307 386
rect 2359 390 2363 391
rect 2359 385 2363 386
rect 2407 390 2411 391
rect 2407 385 2411 386
rect 112 378 114 385
rect 134 384 140 385
rect 134 380 135 384
rect 139 380 140 384
rect 134 379 140 380
rect 174 384 180 385
rect 174 380 175 384
rect 179 380 180 384
rect 174 379 180 380
rect 230 384 236 385
rect 230 380 231 384
rect 235 380 236 384
rect 230 379 236 380
rect 286 384 292 385
rect 286 380 287 384
rect 291 380 292 384
rect 286 379 292 380
rect 342 384 348 385
rect 342 380 343 384
rect 347 380 348 384
rect 342 379 348 380
rect 390 384 396 385
rect 390 380 391 384
rect 395 380 396 384
rect 390 379 396 380
rect 438 384 444 385
rect 438 380 439 384
rect 443 380 444 384
rect 438 379 444 380
rect 486 384 492 385
rect 486 380 487 384
rect 491 380 492 384
rect 486 379 492 380
rect 534 384 540 385
rect 534 380 535 384
rect 539 380 540 384
rect 534 379 540 380
rect 582 384 588 385
rect 582 380 583 384
rect 587 380 588 384
rect 582 379 588 380
rect 630 384 636 385
rect 630 380 631 384
rect 635 380 636 384
rect 630 379 636 380
rect 678 384 684 385
rect 678 380 679 384
rect 683 380 684 384
rect 678 379 684 380
rect 726 384 732 385
rect 726 380 727 384
rect 731 380 732 384
rect 726 379 732 380
rect 774 384 780 385
rect 774 380 775 384
rect 779 380 780 384
rect 774 379 780 380
rect 1240 378 1242 385
rect 1280 378 1282 385
rect 1446 384 1452 385
rect 1446 380 1447 384
rect 1451 380 1452 384
rect 1446 379 1452 380
rect 1486 384 1492 385
rect 1486 380 1487 384
rect 1491 380 1492 384
rect 1486 379 1492 380
rect 1534 384 1540 385
rect 1534 380 1535 384
rect 1539 380 1540 384
rect 1534 379 1540 380
rect 1590 384 1596 385
rect 1590 380 1591 384
rect 1595 380 1596 384
rect 1590 379 1596 380
rect 1662 384 1668 385
rect 1662 380 1663 384
rect 1667 380 1668 384
rect 1662 379 1668 380
rect 1734 384 1740 385
rect 1734 380 1735 384
rect 1739 380 1740 384
rect 1734 379 1740 380
rect 1814 384 1820 385
rect 1814 380 1815 384
rect 1819 380 1820 384
rect 1814 379 1820 380
rect 1894 384 1900 385
rect 1894 380 1895 384
rect 1899 380 1900 384
rect 1894 379 1900 380
rect 1966 384 1972 385
rect 1966 380 1967 384
rect 1971 380 1972 384
rect 1966 379 1972 380
rect 2038 384 2044 385
rect 2038 380 2039 384
rect 2043 380 2044 384
rect 2038 379 2044 380
rect 2110 384 2116 385
rect 2110 380 2111 384
rect 2115 380 2116 384
rect 2110 379 2116 380
rect 2174 384 2180 385
rect 2174 380 2175 384
rect 2179 380 2180 384
rect 2174 379 2180 380
rect 2238 384 2244 385
rect 2238 380 2239 384
rect 2243 380 2244 384
rect 2238 379 2244 380
rect 2302 384 2308 385
rect 2302 380 2303 384
rect 2307 380 2308 384
rect 2302 379 2308 380
rect 2358 384 2364 385
rect 2358 380 2359 384
rect 2363 380 2364 384
rect 2358 379 2364 380
rect 2408 378 2410 385
rect 110 377 116 378
rect 110 373 111 377
rect 115 373 116 377
rect 110 372 116 373
rect 1238 377 1244 378
rect 1238 373 1239 377
rect 1243 373 1244 377
rect 1238 372 1244 373
rect 1278 377 1284 378
rect 1278 373 1279 377
rect 1283 373 1284 377
rect 1278 372 1284 373
rect 2406 377 2412 378
rect 2406 373 2407 377
rect 2411 373 2412 377
rect 2406 372 2412 373
rect 110 360 116 361
rect 110 356 111 360
rect 115 356 116 360
rect 110 355 116 356
rect 1238 360 1244 361
rect 1238 356 1239 360
rect 1243 356 1244 360
rect 1238 355 1244 356
rect 1278 360 1284 361
rect 1278 356 1279 360
rect 1283 356 1284 360
rect 1278 355 1284 356
rect 2406 360 2412 361
rect 2406 356 2407 360
rect 2411 356 2412 360
rect 2406 355 2412 356
rect 112 319 114 355
rect 134 337 140 338
rect 134 333 135 337
rect 139 333 140 337
rect 134 332 140 333
rect 174 337 180 338
rect 174 333 175 337
rect 179 333 180 337
rect 174 332 180 333
rect 230 337 236 338
rect 230 333 231 337
rect 235 333 236 337
rect 230 332 236 333
rect 286 337 292 338
rect 286 333 287 337
rect 291 333 292 337
rect 286 332 292 333
rect 342 337 348 338
rect 342 333 343 337
rect 347 333 348 337
rect 342 332 348 333
rect 390 337 396 338
rect 390 333 391 337
rect 395 333 396 337
rect 390 332 396 333
rect 438 337 444 338
rect 438 333 439 337
rect 443 333 444 337
rect 438 332 444 333
rect 486 337 492 338
rect 486 333 487 337
rect 491 333 492 337
rect 486 332 492 333
rect 534 337 540 338
rect 534 333 535 337
rect 539 333 540 337
rect 534 332 540 333
rect 582 337 588 338
rect 582 333 583 337
rect 587 333 588 337
rect 582 332 588 333
rect 630 337 636 338
rect 630 333 631 337
rect 635 333 636 337
rect 630 332 636 333
rect 678 337 684 338
rect 678 333 679 337
rect 683 333 684 337
rect 678 332 684 333
rect 726 337 732 338
rect 726 333 727 337
rect 731 333 732 337
rect 726 332 732 333
rect 774 337 780 338
rect 774 333 775 337
rect 779 333 780 337
rect 774 332 780 333
rect 136 319 138 332
rect 176 319 178 332
rect 232 319 234 332
rect 288 319 290 332
rect 344 319 346 332
rect 392 319 394 332
rect 440 319 442 332
rect 488 319 490 332
rect 536 319 538 332
rect 584 319 586 332
rect 632 319 634 332
rect 680 319 682 332
rect 728 319 730 332
rect 776 319 778 332
rect 1240 319 1242 355
rect 1280 319 1282 355
rect 1446 337 1452 338
rect 1446 333 1447 337
rect 1451 333 1452 337
rect 1446 332 1452 333
rect 1486 337 1492 338
rect 1486 333 1487 337
rect 1491 333 1492 337
rect 1486 332 1492 333
rect 1534 337 1540 338
rect 1534 333 1535 337
rect 1539 333 1540 337
rect 1534 332 1540 333
rect 1590 337 1596 338
rect 1590 333 1591 337
rect 1595 333 1596 337
rect 1590 332 1596 333
rect 1662 337 1668 338
rect 1662 333 1663 337
rect 1667 333 1668 337
rect 1662 332 1668 333
rect 1734 337 1740 338
rect 1734 333 1735 337
rect 1739 333 1740 337
rect 1734 332 1740 333
rect 1814 337 1820 338
rect 1814 333 1815 337
rect 1819 333 1820 337
rect 1814 332 1820 333
rect 1894 337 1900 338
rect 1894 333 1895 337
rect 1899 333 1900 337
rect 1894 332 1900 333
rect 1966 337 1972 338
rect 1966 333 1967 337
rect 1971 333 1972 337
rect 1966 332 1972 333
rect 2038 337 2044 338
rect 2038 333 2039 337
rect 2043 333 2044 337
rect 2038 332 2044 333
rect 2110 337 2116 338
rect 2110 333 2111 337
rect 2115 333 2116 337
rect 2110 332 2116 333
rect 2174 337 2180 338
rect 2174 333 2175 337
rect 2179 333 2180 337
rect 2174 332 2180 333
rect 2238 337 2244 338
rect 2238 333 2239 337
rect 2243 333 2244 337
rect 2238 332 2244 333
rect 2302 337 2308 338
rect 2302 333 2303 337
rect 2307 333 2308 337
rect 2302 332 2308 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 1448 319 1450 332
rect 1488 319 1490 332
rect 1536 319 1538 332
rect 1592 319 1594 332
rect 1664 319 1666 332
rect 1736 319 1738 332
rect 1816 319 1818 332
rect 1896 319 1898 332
rect 1968 319 1970 332
rect 2040 319 2042 332
rect 2112 319 2114 332
rect 2176 319 2178 332
rect 2240 319 2242 332
rect 2304 319 2306 332
rect 2360 319 2362 332
rect 2408 319 2410 355
rect 111 318 115 319
rect 111 313 115 314
rect 135 318 139 319
rect 135 313 139 314
rect 175 318 179 319
rect 175 313 179 314
rect 183 318 187 319
rect 183 313 187 314
rect 231 318 235 319
rect 231 313 235 314
rect 255 318 259 319
rect 255 313 259 314
rect 287 318 291 319
rect 287 313 291 314
rect 327 318 331 319
rect 327 313 331 314
rect 343 318 347 319
rect 343 313 347 314
rect 391 318 395 319
rect 391 313 395 314
rect 439 318 443 319
rect 439 313 443 314
rect 447 318 451 319
rect 447 313 451 314
rect 487 318 491 319
rect 487 313 491 314
rect 503 318 507 319
rect 503 313 507 314
rect 535 318 539 319
rect 535 313 539 314
rect 551 318 555 319
rect 551 313 555 314
rect 583 318 587 319
rect 583 313 587 314
rect 591 318 595 319
rect 591 313 595 314
rect 631 318 635 319
rect 631 313 635 314
rect 679 318 683 319
rect 679 313 683 314
rect 727 318 731 319
rect 727 313 731 314
rect 775 318 779 319
rect 775 313 779 314
rect 823 318 827 319
rect 823 313 827 314
rect 871 318 875 319
rect 871 313 875 314
rect 919 318 923 319
rect 919 313 923 314
rect 1239 318 1243 319
rect 1239 313 1243 314
rect 1279 318 1283 319
rect 1279 313 1283 314
rect 1447 318 1451 319
rect 1447 313 1451 314
rect 1487 318 1491 319
rect 1487 313 1491 314
rect 1495 318 1499 319
rect 1495 313 1499 314
rect 1535 318 1539 319
rect 1535 313 1539 314
rect 1575 318 1579 319
rect 1575 313 1579 314
rect 1591 318 1595 319
rect 1591 313 1595 314
rect 1615 318 1619 319
rect 1615 313 1619 314
rect 1655 318 1659 319
rect 1655 313 1659 314
rect 1663 318 1667 319
rect 1663 313 1667 314
rect 1695 318 1699 319
rect 1695 313 1699 314
rect 1735 318 1739 319
rect 1735 313 1739 314
rect 1743 318 1747 319
rect 1743 313 1747 314
rect 1799 318 1803 319
rect 1799 313 1803 314
rect 1815 318 1819 319
rect 1815 313 1819 314
rect 1863 318 1867 319
rect 1863 313 1867 314
rect 1895 318 1899 319
rect 1895 313 1899 314
rect 1935 318 1939 319
rect 1935 313 1939 314
rect 1967 318 1971 319
rect 1967 313 1971 314
rect 2007 318 2011 319
rect 2007 313 2011 314
rect 2039 318 2043 319
rect 2039 313 2043 314
rect 2071 318 2075 319
rect 2071 313 2075 314
rect 2111 318 2115 319
rect 2111 313 2115 314
rect 2135 318 2139 319
rect 2135 313 2139 314
rect 2175 318 2179 319
rect 2175 313 2179 314
rect 2191 318 2195 319
rect 2191 313 2195 314
rect 2239 318 2243 319
rect 2239 313 2243 314
rect 2255 318 2259 319
rect 2255 313 2259 314
rect 2303 318 2307 319
rect 2303 313 2307 314
rect 2319 318 2323 319
rect 2319 313 2323 314
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 112 281 114 313
rect 136 304 138 313
rect 184 304 186 313
rect 256 304 258 313
rect 328 304 330 313
rect 392 304 394 313
rect 448 304 450 313
rect 504 304 506 313
rect 552 304 554 313
rect 592 304 594 313
rect 632 304 634 313
rect 680 304 682 313
rect 728 304 730 313
rect 776 304 778 313
rect 824 304 826 313
rect 872 304 874 313
rect 920 304 922 313
rect 134 303 140 304
rect 134 299 135 303
rect 139 299 140 303
rect 134 298 140 299
rect 182 303 188 304
rect 182 299 183 303
rect 187 299 188 303
rect 182 298 188 299
rect 254 303 260 304
rect 254 299 255 303
rect 259 299 260 303
rect 254 298 260 299
rect 326 303 332 304
rect 326 299 327 303
rect 331 299 332 303
rect 326 298 332 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 446 303 452 304
rect 446 299 447 303
rect 451 299 452 303
rect 446 298 452 299
rect 502 303 508 304
rect 502 299 503 303
rect 507 299 508 303
rect 502 298 508 299
rect 550 303 556 304
rect 550 299 551 303
rect 555 299 556 303
rect 550 298 556 299
rect 590 303 596 304
rect 590 299 591 303
rect 595 299 596 303
rect 590 298 596 299
rect 630 303 636 304
rect 630 299 631 303
rect 635 299 636 303
rect 630 298 636 299
rect 678 303 684 304
rect 678 299 679 303
rect 683 299 684 303
rect 678 298 684 299
rect 726 303 732 304
rect 726 299 727 303
rect 731 299 732 303
rect 726 298 732 299
rect 774 303 780 304
rect 774 299 775 303
rect 779 299 780 303
rect 774 298 780 299
rect 822 303 828 304
rect 822 299 823 303
rect 827 299 828 303
rect 822 298 828 299
rect 870 303 876 304
rect 870 299 871 303
rect 875 299 876 303
rect 870 298 876 299
rect 918 303 924 304
rect 918 299 919 303
rect 923 299 924 303
rect 918 298 924 299
rect 1240 281 1242 313
rect 1280 281 1282 313
rect 1496 304 1498 313
rect 1536 304 1538 313
rect 1576 304 1578 313
rect 1616 304 1618 313
rect 1656 304 1658 313
rect 1696 304 1698 313
rect 1744 304 1746 313
rect 1800 304 1802 313
rect 1864 304 1866 313
rect 1936 304 1938 313
rect 2008 304 2010 313
rect 2072 304 2074 313
rect 2136 304 2138 313
rect 2192 304 2194 313
rect 2256 304 2258 313
rect 2320 304 2322 313
rect 2360 304 2362 313
rect 1494 303 1500 304
rect 1494 299 1495 303
rect 1499 299 1500 303
rect 1494 298 1500 299
rect 1534 303 1540 304
rect 1534 299 1535 303
rect 1539 299 1540 303
rect 1534 298 1540 299
rect 1574 303 1580 304
rect 1574 299 1575 303
rect 1579 299 1580 303
rect 1574 298 1580 299
rect 1614 303 1620 304
rect 1614 299 1615 303
rect 1619 299 1620 303
rect 1614 298 1620 299
rect 1654 303 1660 304
rect 1654 299 1655 303
rect 1659 299 1660 303
rect 1654 298 1660 299
rect 1694 303 1700 304
rect 1694 299 1695 303
rect 1699 299 1700 303
rect 1694 298 1700 299
rect 1742 303 1748 304
rect 1742 299 1743 303
rect 1747 299 1748 303
rect 1742 298 1748 299
rect 1798 303 1804 304
rect 1798 299 1799 303
rect 1803 299 1804 303
rect 1798 298 1804 299
rect 1862 303 1868 304
rect 1862 299 1863 303
rect 1867 299 1868 303
rect 1862 298 1868 299
rect 1934 303 1940 304
rect 1934 299 1935 303
rect 1939 299 1940 303
rect 1934 298 1940 299
rect 2006 303 2012 304
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2070 303 2076 304
rect 2070 299 2071 303
rect 2075 299 2076 303
rect 2070 298 2076 299
rect 2134 303 2140 304
rect 2134 299 2135 303
rect 2139 299 2140 303
rect 2134 298 2140 299
rect 2190 303 2196 304
rect 2190 299 2191 303
rect 2195 299 2196 303
rect 2190 298 2196 299
rect 2254 303 2260 304
rect 2254 299 2255 303
rect 2259 299 2260 303
rect 2254 298 2260 299
rect 2318 303 2324 304
rect 2318 299 2319 303
rect 2323 299 2324 303
rect 2318 298 2324 299
rect 2358 303 2364 304
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2358 298 2364 299
rect 2408 281 2410 313
rect 110 280 116 281
rect 110 276 111 280
rect 115 276 116 280
rect 110 275 116 276
rect 1238 280 1244 281
rect 1238 276 1239 280
rect 1243 276 1244 280
rect 1238 275 1244 276
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 1278 275 1284 276
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2406 275 2412 276
rect 110 263 116 264
rect 110 259 111 263
rect 115 259 116 263
rect 110 258 116 259
rect 1238 263 1244 264
rect 1238 259 1239 263
rect 1243 259 1244 263
rect 1238 258 1244 259
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1278 258 1284 259
rect 2406 263 2412 264
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 112 243 114 258
rect 134 256 140 257
rect 134 252 135 256
rect 139 252 140 256
rect 134 251 140 252
rect 182 256 188 257
rect 182 252 183 256
rect 187 252 188 256
rect 182 251 188 252
rect 254 256 260 257
rect 254 252 255 256
rect 259 252 260 256
rect 254 251 260 252
rect 326 256 332 257
rect 326 252 327 256
rect 331 252 332 256
rect 326 251 332 252
rect 390 256 396 257
rect 390 252 391 256
rect 395 252 396 256
rect 390 251 396 252
rect 446 256 452 257
rect 446 252 447 256
rect 451 252 452 256
rect 446 251 452 252
rect 502 256 508 257
rect 502 252 503 256
rect 507 252 508 256
rect 502 251 508 252
rect 550 256 556 257
rect 550 252 551 256
rect 555 252 556 256
rect 550 251 556 252
rect 590 256 596 257
rect 590 252 591 256
rect 595 252 596 256
rect 590 251 596 252
rect 630 256 636 257
rect 630 252 631 256
rect 635 252 636 256
rect 630 251 636 252
rect 678 256 684 257
rect 678 252 679 256
rect 683 252 684 256
rect 678 251 684 252
rect 726 256 732 257
rect 726 252 727 256
rect 731 252 732 256
rect 726 251 732 252
rect 774 256 780 257
rect 774 252 775 256
rect 779 252 780 256
rect 774 251 780 252
rect 822 256 828 257
rect 822 252 823 256
rect 827 252 828 256
rect 822 251 828 252
rect 870 256 876 257
rect 870 252 871 256
rect 875 252 876 256
rect 870 251 876 252
rect 918 256 924 257
rect 918 252 919 256
rect 923 252 924 256
rect 918 251 924 252
rect 136 243 138 251
rect 184 243 186 251
rect 256 243 258 251
rect 328 243 330 251
rect 392 243 394 251
rect 448 243 450 251
rect 504 243 506 251
rect 552 243 554 251
rect 592 243 594 251
rect 632 243 634 251
rect 680 243 682 251
rect 728 243 730 251
rect 776 243 778 251
rect 824 243 826 251
rect 872 243 874 251
rect 920 243 922 251
rect 1240 243 1242 258
rect 1280 247 1282 258
rect 1494 256 1500 257
rect 1494 252 1495 256
rect 1499 252 1500 256
rect 1494 251 1500 252
rect 1534 256 1540 257
rect 1534 252 1535 256
rect 1539 252 1540 256
rect 1534 251 1540 252
rect 1574 256 1580 257
rect 1574 252 1575 256
rect 1579 252 1580 256
rect 1574 251 1580 252
rect 1614 256 1620 257
rect 1614 252 1615 256
rect 1619 252 1620 256
rect 1614 251 1620 252
rect 1654 256 1660 257
rect 1654 252 1655 256
rect 1659 252 1660 256
rect 1654 251 1660 252
rect 1694 256 1700 257
rect 1694 252 1695 256
rect 1699 252 1700 256
rect 1694 251 1700 252
rect 1742 256 1748 257
rect 1742 252 1743 256
rect 1747 252 1748 256
rect 1742 251 1748 252
rect 1798 256 1804 257
rect 1798 252 1799 256
rect 1803 252 1804 256
rect 1798 251 1804 252
rect 1862 256 1868 257
rect 1862 252 1863 256
rect 1867 252 1868 256
rect 1862 251 1868 252
rect 1934 256 1940 257
rect 1934 252 1935 256
rect 1939 252 1940 256
rect 1934 251 1940 252
rect 2006 256 2012 257
rect 2006 252 2007 256
rect 2011 252 2012 256
rect 2006 251 2012 252
rect 2070 256 2076 257
rect 2070 252 2071 256
rect 2075 252 2076 256
rect 2070 251 2076 252
rect 2134 256 2140 257
rect 2134 252 2135 256
rect 2139 252 2140 256
rect 2134 251 2140 252
rect 2190 256 2196 257
rect 2190 252 2191 256
rect 2195 252 2196 256
rect 2190 251 2196 252
rect 2254 256 2260 257
rect 2254 252 2255 256
rect 2259 252 2260 256
rect 2254 251 2260 252
rect 2318 256 2324 257
rect 2318 252 2319 256
rect 2323 252 2324 256
rect 2318 251 2324 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 1496 247 1498 251
rect 1536 247 1538 251
rect 1576 247 1578 251
rect 1616 247 1618 251
rect 1656 247 1658 251
rect 1696 247 1698 251
rect 1744 247 1746 251
rect 1800 247 1802 251
rect 1864 247 1866 251
rect 1936 247 1938 251
rect 2008 247 2010 251
rect 2072 247 2074 251
rect 2136 247 2138 251
rect 2192 247 2194 251
rect 2256 247 2258 251
rect 2320 247 2322 251
rect 2360 247 2362 251
rect 2408 247 2410 258
rect 1279 246 1283 247
rect 111 242 115 243
rect 111 237 115 238
rect 135 242 139 243
rect 135 237 139 238
rect 175 242 179 243
rect 175 237 179 238
rect 183 242 187 243
rect 183 237 187 238
rect 247 242 251 243
rect 247 237 251 238
rect 255 242 259 243
rect 255 237 259 238
rect 327 242 331 243
rect 327 237 331 238
rect 391 242 395 243
rect 391 237 395 238
rect 415 242 419 243
rect 415 237 419 238
rect 447 242 451 243
rect 447 237 451 238
rect 495 242 499 243
rect 495 237 499 238
rect 503 242 507 243
rect 503 237 507 238
rect 551 242 555 243
rect 551 237 555 238
rect 575 242 579 243
rect 575 237 579 238
rect 591 242 595 243
rect 591 237 595 238
rect 631 242 635 243
rect 631 237 635 238
rect 655 242 659 243
rect 655 237 659 238
rect 679 242 683 243
rect 679 237 683 238
rect 727 242 731 243
rect 727 237 731 238
rect 775 242 779 243
rect 775 237 779 238
rect 791 242 795 243
rect 791 237 795 238
rect 823 242 827 243
rect 823 237 827 238
rect 847 242 851 243
rect 847 237 851 238
rect 871 242 875 243
rect 871 237 875 238
rect 903 242 907 243
rect 903 237 907 238
rect 919 242 923 243
rect 919 237 923 238
rect 959 242 963 243
rect 959 237 963 238
rect 1023 242 1027 243
rect 1023 237 1027 238
rect 1239 242 1243 243
rect 1279 241 1283 242
rect 1367 246 1371 247
rect 1367 241 1371 242
rect 1407 246 1411 247
rect 1407 241 1411 242
rect 1447 246 1451 247
rect 1447 241 1451 242
rect 1495 246 1499 247
rect 1495 241 1499 242
rect 1535 246 1539 247
rect 1535 241 1539 242
rect 1551 246 1555 247
rect 1551 241 1555 242
rect 1575 246 1579 247
rect 1575 241 1579 242
rect 1607 246 1611 247
rect 1607 241 1611 242
rect 1615 246 1619 247
rect 1615 241 1619 242
rect 1655 246 1659 247
rect 1655 241 1659 242
rect 1671 246 1675 247
rect 1671 241 1675 242
rect 1695 246 1699 247
rect 1695 241 1699 242
rect 1735 246 1739 247
rect 1735 241 1739 242
rect 1743 246 1747 247
rect 1743 241 1747 242
rect 1799 246 1803 247
rect 1799 241 1803 242
rect 1807 246 1811 247
rect 1807 241 1811 242
rect 1863 246 1867 247
rect 1863 241 1867 242
rect 1887 246 1891 247
rect 1887 241 1891 242
rect 1935 246 1939 247
rect 1935 241 1939 242
rect 1975 246 1979 247
rect 1975 241 1979 242
rect 2007 246 2011 247
rect 2007 241 2011 242
rect 2071 246 2075 247
rect 2071 241 2075 242
rect 2135 246 2139 247
rect 2135 241 2139 242
rect 2167 246 2171 247
rect 2167 241 2171 242
rect 2191 246 2195 247
rect 2191 241 2195 242
rect 2255 246 2259 247
rect 2255 241 2259 242
rect 2271 246 2275 247
rect 2271 241 2275 242
rect 2319 246 2323 247
rect 2319 241 2323 242
rect 2359 246 2363 247
rect 2359 241 2363 242
rect 2407 246 2411 247
rect 2407 241 2411 242
rect 1239 237 1243 238
rect 112 230 114 237
rect 134 236 140 237
rect 134 232 135 236
rect 139 232 140 236
rect 134 231 140 232
rect 174 236 180 237
rect 174 232 175 236
rect 179 232 180 236
rect 174 231 180 232
rect 246 236 252 237
rect 246 232 247 236
rect 251 232 252 236
rect 246 231 252 232
rect 326 236 332 237
rect 326 232 327 236
rect 331 232 332 236
rect 326 231 332 232
rect 414 236 420 237
rect 414 232 415 236
rect 419 232 420 236
rect 414 231 420 232
rect 494 236 500 237
rect 494 232 495 236
rect 499 232 500 236
rect 494 231 500 232
rect 574 236 580 237
rect 574 232 575 236
rect 579 232 580 236
rect 574 231 580 232
rect 654 236 660 237
rect 654 232 655 236
rect 659 232 660 236
rect 654 231 660 232
rect 726 236 732 237
rect 726 232 727 236
rect 731 232 732 236
rect 726 231 732 232
rect 790 236 796 237
rect 790 232 791 236
rect 795 232 796 236
rect 790 231 796 232
rect 846 236 852 237
rect 846 232 847 236
rect 851 232 852 236
rect 846 231 852 232
rect 902 236 908 237
rect 902 232 903 236
rect 907 232 908 236
rect 902 231 908 232
rect 958 236 964 237
rect 958 232 959 236
rect 963 232 964 236
rect 958 231 964 232
rect 1022 236 1028 237
rect 1022 232 1023 236
rect 1027 232 1028 236
rect 1022 231 1028 232
rect 1240 230 1242 237
rect 1280 234 1282 241
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1446 240 1452 241
rect 1446 236 1447 240
rect 1451 236 1452 240
rect 1446 235 1452 236
rect 1494 240 1500 241
rect 1494 236 1495 240
rect 1499 236 1500 240
rect 1494 235 1500 236
rect 1550 240 1556 241
rect 1550 236 1551 240
rect 1555 236 1556 240
rect 1550 235 1556 236
rect 1606 240 1612 241
rect 1606 236 1607 240
rect 1611 236 1612 240
rect 1606 235 1612 236
rect 1670 240 1676 241
rect 1670 236 1671 240
rect 1675 236 1676 240
rect 1670 235 1676 236
rect 1734 240 1740 241
rect 1734 236 1735 240
rect 1739 236 1740 240
rect 1734 235 1740 236
rect 1806 240 1812 241
rect 1806 236 1807 240
rect 1811 236 1812 240
rect 1806 235 1812 236
rect 1886 240 1892 241
rect 1886 236 1887 240
rect 1891 236 1892 240
rect 1886 235 1892 236
rect 1974 240 1980 241
rect 1974 236 1975 240
rect 1979 236 1980 240
rect 1974 235 1980 236
rect 2070 240 2076 241
rect 2070 236 2071 240
rect 2075 236 2076 240
rect 2070 235 2076 236
rect 2166 240 2172 241
rect 2166 236 2167 240
rect 2171 236 2172 240
rect 2166 235 2172 236
rect 2270 240 2276 241
rect 2270 236 2271 240
rect 2275 236 2276 240
rect 2270 235 2276 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 2408 234 2410 241
rect 1278 233 1284 234
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 110 224 116 225
rect 1238 229 1244 230
rect 1238 225 1239 229
rect 1243 225 1244 229
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 1238 224 1244 225
rect 1278 216 1284 217
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 110 207 116 208
rect 1238 212 1244 213
rect 1238 208 1239 212
rect 1243 208 1244 212
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1278 211 1284 212
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 1238 207 1244 208
rect 112 155 114 207
rect 134 189 140 190
rect 134 185 135 189
rect 139 185 140 189
rect 134 184 140 185
rect 174 189 180 190
rect 174 185 175 189
rect 179 185 180 189
rect 174 184 180 185
rect 246 189 252 190
rect 246 185 247 189
rect 251 185 252 189
rect 246 184 252 185
rect 326 189 332 190
rect 326 185 327 189
rect 331 185 332 189
rect 326 184 332 185
rect 414 189 420 190
rect 414 185 415 189
rect 419 185 420 189
rect 414 184 420 185
rect 494 189 500 190
rect 494 185 495 189
rect 499 185 500 189
rect 494 184 500 185
rect 574 189 580 190
rect 574 185 575 189
rect 579 185 580 189
rect 574 184 580 185
rect 654 189 660 190
rect 654 185 655 189
rect 659 185 660 189
rect 654 184 660 185
rect 726 189 732 190
rect 726 185 727 189
rect 731 185 732 189
rect 726 184 732 185
rect 790 189 796 190
rect 790 185 791 189
rect 795 185 796 189
rect 790 184 796 185
rect 846 189 852 190
rect 846 185 847 189
rect 851 185 852 189
rect 846 184 852 185
rect 902 189 908 190
rect 902 185 903 189
rect 907 185 908 189
rect 902 184 908 185
rect 958 189 964 190
rect 958 185 959 189
rect 963 185 964 189
rect 958 184 964 185
rect 1022 189 1028 190
rect 1022 185 1023 189
rect 1027 185 1028 189
rect 1022 184 1028 185
rect 136 155 138 184
rect 176 155 178 184
rect 248 155 250 184
rect 328 155 330 184
rect 416 155 418 184
rect 496 155 498 184
rect 576 155 578 184
rect 656 155 658 184
rect 728 155 730 184
rect 792 155 794 184
rect 848 155 850 184
rect 904 155 906 184
rect 960 155 962 184
rect 1024 155 1026 184
rect 1240 155 1242 207
rect 1280 163 1282 211
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1446 193 1452 194
rect 1446 189 1447 193
rect 1451 189 1452 193
rect 1446 188 1452 189
rect 1494 193 1500 194
rect 1494 189 1495 193
rect 1499 189 1500 193
rect 1494 188 1500 189
rect 1550 193 1556 194
rect 1550 189 1551 193
rect 1555 189 1556 193
rect 1550 188 1556 189
rect 1606 193 1612 194
rect 1606 189 1607 193
rect 1611 189 1612 193
rect 1606 188 1612 189
rect 1670 193 1676 194
rect 1670 189 1671 193
rect 1675 189 1676 193
rect 1670 188 1676 189
rect 1734 193 1740 194
rect 1734 189 1735 193
rect 1739 189 1740 193
rect 1734 188 1740 189
rect 1806 193 1812 194
rect 1806 189 1807 193
rect 1811 189 1812 193
rect 1806 188 1812 189
rect 1886 193 1892 194
rect 1886 189 1887 193
rect 1891 189 1892 193
rect 1886 188 1892 189
rect 1974 193 1980 194
rect 1974 189 1975 193
rect 1979 189 1980 193
rect 1974 188 1980 189
rect 2070 193 2076 194
rect 2070 189 2071 193
rect 2075 189 2076 193
rect 2070 188 2076 189
rect 2166 193 2172 194
rect 2166 189 2167 193
rect 2171 189 2172 193
rect 2166 188 2172 189
rect 2270 193 2276 194
rect 2270 189 2271 193
rect 2275 189 2276 193
rect 2270 188 2276 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1368 163 1370 188
rect 1408 163 1410 188
rect 1448 163 1450 188
rect 1496 163 1498 188
rect 1552 163 1554 188
rect 1608 163 1610 188
rect 1672 163 1674 188
rect 1736 163 1738 188
rect 1808 163 1810 188
rect 1888 163 1890 188
rect 1976 163 1978 188
rect 2072 163 2074 188
rect 2168 163 2170 188
rect 2272 163 2274 188
rect 2360 163 2362 188
rect 2408 163 2410 211
rect 1279 162 1283 163
rect 1279 157 1283 158
rect 1303 162 1307 163
rect 1303 157 1307 158
rect 1343 162 1347 163
rect 1343 157 1347 158
rect 1367 162 1371 163
rect 1367 157 1371 158
rect 1383 162 1387 163
rect 1383 157 1387 158
rect 1407 162 1411 163
rect 1407 157 1411 158
rect 1423 162 1427 163
rect 1423 157 1427 158
rect 1447 162 1451 163
rect 1447 157 1451 158
rect 1463 162 1467 163
rect 1463 157 1467 158
rect 1495 162 1499 163
rect 1495 157 1499 158
rect 1519 162 1523 163
rect 1519 157 1523 158
rect 1551 162 1555 163
rect 1551 157 1555 158
rect 1583 162 1587 163
rect 1583 157 1587 158
rect 1607 162 1611 163
rect 1607 157 1611 158
rect 1647 162 1651 163
rect 1647 157 1651 158
rect 1671 162 1675 163
rect 1671 157 1675 158
rect 1711 162 1715 163
rect 1711 157 1715 158
rect 1735 162 1739 163
rect 1735 157 1739 158
rect 1767 162 1771 163
rect 1767 157 1771 158
rect 1807 162 1811 163
rect 1807 157 1811 158
rect 1823 162 1827 163
rect 1823 157 1827 158
rect 1871 162 1875 163
rect 1871 157 1875 158
rect 1887 162 1891 163
rect 1887 157 1891 158
rect 1919 162 1923 163
rect 1919 157 1923 158
rect 1967 162 1971 163
rect 1967 157 1971 158
rect 1975 162 1979 163
rect 1975 157 1979 158
rect 2015 162 2019 163
rect 2015 157 2019 158
rect 2063 162 2067 163
rect 2063 157 2067 158
rect 2071 162 2075 163
rect 2071 157 2075 158
rect 2111 162 2115 163
rect 2111 157 2115 158
rect 2159 162 2163 163
rect 2159 157 2163 158
rect 2167 162 2171 163
rect 2167 157 2171 158
rect 2215 162 2219 163
rect 2215 157 2219 158
rect 2271 162 2275 163
rect 2271 157 2275 158
rect 2319 162 2323 163
rect 2319 157 2323 158
rect 2359 162 2363 163
rect 2359 157 2363 158
rect 2407 162 2411 163
rect 2407 157 2411 158
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 175 154 179 155
rect 175 149 179 150
rect 215 154 219 155
rect 215 149 219 150
rect 247 154 251 155
rect 247 149 251 150
rect 255 154 259 155
rect 255 149 259 150
rect 295 154 299 155
rect 295 149 299 150
rect 327 154 331 155
rect 327 149 331 150
rect 335 154 339 155
rect 335 149 339 150
rect 375 154 379 155
rect 375 149 379 150
rect 415 154 419 155
rect 415 149 419 150
rect 423 154 427 155
rect 423 149 427 150
rect 471 154 475 155
rect 471 149 475 150
rect 495 154 499 155
rect 495 149 499 150
rect 527 154 531 155
rect 527 149 531 150
rect 575 154 579 155
rect 575 149 579 150
rect 583 154 587 155
rect 583 149 587 150
rect 631 154 635 155
rect 631 149 635 150
rect 655 154 659 155
rect 655 149 659 150
rect 679 154 683 155
rect 679 149 683 150
rect 727 154 731 155
rect 727 149 731 150
rect 767 154 771 155
rect 767 149 771 150
rect 791 154 795 155
rect 791 149 795 150
rect 807 154 811 155
rect 807 149 811 150
rect 847 154 851 155
rect 847 149 851 150
rect 887 154 891 155
rect 887 149 891 150
rect 903 154 907 155
rect 903 149 907 150
rect 927 154 931 155
rect 927 149 931 150
rect 959 154 963 155
rect 959 149 963 150
rect 975 154 979 155
rect 975 149 979 150
rect 1023 154 1027 155
rect 1023 149 1027 150
rect 1071 154 1075 155
rect 1071 149 1075 150
rect 1111 154 1115 155
rect 1111 149 1115 150
rect 1151 154 1155 155
rect 1151 149 1155 150
rect 1191 154 1195 155
rect 1191 149 1195 150
rect 1239 154 1243 155
rect 1239 149 1243 150
rect 112 117 114 149
rect 136 140 138 149
rect 176 140 178 149
rect 216 140 218 149
rect 256 140 258 149
rect 296 140 298 149
rect 336 140 338 149
rect 376 140 378 149
rect 424 140 426 149
rect 472 140 474 149
rect 528 140 530 149
rect 584 140 586 149
rect 632 140 634 149
rect 680 140 682 149
rect 728 140 730 149
rect 768 140 770 149
rect 808 140 810 149
rect 848 140 850 149
rect 888 140 890 149
rect 928 140 930 149
rect 976 140 978 149
rect 1024 140 1026 149
rect 1072 140 1074 149
rect 1112 140 1114 149
rect 1152 140 1154 149
rect 1192 140 1194 149
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 174 139 180 140
rect 174 135 175 139
rect 179 135 180 139
rect 174 134 180 135
rect 214 139 220 140
rect 214 135 215 139
rect 219 135 220 139
rect 214 134 220 135
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 294 139 300 140
rect 294 135 295 139
rect 299 135 300 139
rect 294 134 300 135
rect 334 139 340 140
rect 334 135 335 139
rect 339 135 340 139
rect 334 134 340 135
rect 374 139 380 140
rect 374 135 375 139
rect 379 135 380 139
rect 374 134 380 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 470 139 476 140
rect 470 135 471 139
rect 475 135 476 139
rect 470 134 476 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 582 139 588 140
rect 582 135 583 139
rect 587 135 588 139
rect 582 134 588 135
rect 630 139 636 140
rect 630 135 631 139
rect 635 135 636 139
rect 630 134 636 135
rect 678 139 684 140
rect 678 135 679 139
rect 683 135 684 139
rect 678 134 684 135
rect 726 139 732 140
rect 726 135 727 139
rect 731 135 732 139
rect 726 134 732 135
rect 766 139 772 140
rect 766 135 767 139
rect 771 135 772 139
rect 766 134 772 135
rect 806 139 812 140
rect 806 135 807 139
rect 811 135 812 139
rect 806 134 812 135
rect 846 139 852 140
rect 846 135 847 139
rect 851 135 852 139
rect 846 134 852 135
rect 886 139 892 140
rect 886 135 887 139
rect 891 135 892 139
rect 886 134 892 135
rect 926 139 932 140
rect 926 135 927 139
rect 931 135 932 139
rect 926 134 932 135
rect 974 139 980 140
rect 974 135 975 139
rect 979 135 980 139
rect 974 134 980 135
rect 1022 139 1028 140
rect 1022 135 1023 139
rect 1027 135 1028 139
rect 1022 134 1028 135
rect 1070 139 1076 140
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1070 134 1076 135
rect 1110 139 1116 140
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1240 117 1242 149
rect 1280 125 1282 157
rect 1304 148 1306 157
rect 1344 148 1346 157
rect 1384 148 1386 157
rect 1424 148 1426 157
rect 1464 148 1466 157
rect 1520 148 1522 157
rect 1584 148 1586 157
rect 1648 148 1650 157
rect 1712 148 1714 157
rect 1768 148 1770 157
rect 1824 148 1826 157
rect 1872 148 1874 157
rect 1920 148 1922 157
rect 1968 148 1970 157
rect 2016 148 2018 157
rect 2064 148 2066 157
rect 2112 148 2114 157
rect 2160 148 2162 157
rect 2216 148 2218 157
rect 2272 148 2274 157
rect 2320 148 2322 157
rect 2360 148 2362 157
rect 1302 147 1308 148
rect 1302 143 1303 147
rect 1307 143 1308 147
rect 1302 142 1308 143
rect 1342 147 1348 148
rect 1342 143 1343 147
rect 1347 143 1348 147
rect 1342 142 1348 143
rect 1382 147 1388 148
rect 1382 143 1383 147
rect 1387 143 1388 147
rect 1382 142 1388 143
rect 1422 147 1428 148
rect 1422 143 1423 147
rect 1427 143 1428 147
rect 1422 142 1428 143
rect 1462 147 1468 148
rect 1462 143 1463 147
rect 1467 143 1468 147
rect 1462 142 1468 143
rect 1518 147 1524 148
rect 1518 143 1519 147
rect 1523 143 1524 147
rect 1518 142 1524 143
rect 1582 147 1588 148
rect 1582 143 1583 147
rect 1587 143 1588 147
rect 1582 142 1588 143
rect 1646 147 1652 148
rect 1646 143 1647 147
rect 1651 143 1652 147
rect 1646 142 1652 143
rect 1710 147 1716 148
rect 1710 143 1711 147
rect 1715 143 1716 147
rect 1710 142 1716 143
rect 1766 147 1772 148
rect 1766 143 1767 147
rect 1771 143 1772 147
rect 1766 142 1772 143
rect 1822 147 1828 148
rect 1822 143 1823 147
rect 1827 143 1828 147
rect 1822 142 1828 143
rect 1870 147 1876 148
rect 1870 143 1871 147
rect 1875 143 1876 147
rect 1870 142 1876 143
rect 1918 147 1924 148
rect 1918 143 1919 147
rect 1923 143 1924 147
rect 1918 142 1924 143
rect 1966 147 1972 148
rect 1966 143 1967 147
rect 1971 143 1972 147
rect 1966 142 1972 143
rect 2014 147 2020 148
rect 2014 143 2015 147
rect 2019 143 2020 147
rect 2014 142 2020 143
rect 2062 147 2068 148
rect 2062 143 2063 147
rect 2067 143 2068 147
rect 2062 142 2068 143
rect 2110 147 2116 148
rect 2110 143 2111 147
rect 2115 143 2116 147
rect 2110 142 2116 143
rect 2158 147 2164 148
rect 2158 143 2159 147
rect 2163 143 2164 147
rect 2158 142 2164 143
rect 2214 147 2220 148
rect 2214 143 2215 147
rect 2219 143 2220 147
rect 2214 142 2220 143
rect 2270 147 2276 148
rect 2270 143 2271 147
rect 2275 143 2276 147
rect 2270 142 2276 143
rect 2318 147 2324 148
rect 2318 143 2319 147
rect 2323 143 2324 147
rect 2318 142 2324 143
rect 2358 147 2364 148
rect 2358 143 2359 147
rect 2363 143 2364 147
rect 2358 142 2364 143
rect 2408 125 2410 157
rect 1278 124 1284 125
rect 1278 120 1279 124
rect 1283 120 1284 124
rect 1278 119 1284 120
rect 2406 124 2412 125
rect 2406 120 2407 124
rect 2411 120 2412 124
rect 2406 119 2412 120
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 110 111 116 112
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1238 111 1244 112
rect 1278 107 1284 108
rect 1278 103 1279 107
rect 1283 103 1284 107
rect 1278 102 1284 103
rect 2406 107 2412 108
rect 2406 103 2407 107
rect 2411 103 2412 107
rect 2406 102 2412 103
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1280 95 1282 102
rect 1302 100 1308 101
rect 1302 96 1303 100
rect 1307 96 1308 100
rect 1302 95 1308 96
rect 1342 100 1348 101
rect 1342 96 1343 100
rect 1347 96 1348 100
rect 1342 95 1348 96
rect 1382 100 1388 101
rect 1382 96 1383 100
rect 1387 96 1388 100
rect 1382 95 1388 96
rect 1422 100 1428 101
rect 1422 96 1423 100
rect 1427 96 1428 100
rect 1422 95 1428 96
rect 1462 100 1468 101
rect 1462 96 1463 100
rect 1467 96 1468 100
rect 1462 95 1468 96
rect 1518 100 1524 101
rect 1518 96 1519 100
rect 1523 96 1524 100
rect 1518 95 1524 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1646 100 1652 101
rect 1646 96 1647 100
rect 1651 96 1652 100
rect 1646 95 1652 96
rect 1710 100 1716 101
rect 1710 96 1711 100
rect 1715 96 1716 100
rect 1710 95 1716 96
rect 1766 100 1772 101
rect 1766 96 1767 100
rect 1771 96 1772 100
rect 1766 95 1772 96
rect 1822 100 1828 101
rect 1822 96 1823 100
rect 1827 96 1828 100
rect 1822 95 1828 96
rect 1870 100 1876 101
rect 1870 96 1871 100
rect 1875 96 1876 100
rect 1870 95 1876 96
rect 1918 100 1924 101
rect 1918 96 1919 100
rect 1923 96 1924 100
rect 1918 95 1924 96
rect 1966 100 1972 101
rect 1966 96 1967 100
rect 1971 96 1972 100
rect 1966 95 1972 96
rect 2014 100 2020 101
rect 2014 96 2015 100
rect 2019 96 2020 100
rect 2014 95 2020 96
rect 2062 100 2068 101
rect 2062 96 2063 100
rect 2067 96 2068 100
rect 2062 95 2068 96
rect 2110 100 2116 101
rect 2110 96 2111 100
rect 2115 96 2116 100
rect 2110 95 2116 96
rect 2158 100 2164 101
rect 2158 96 2159 100
rect 2163 96 2164 100
rect 2158 95 2164 96
rect 2214 100 2220 101
rect 2214 96 2215 100
rect 2219 96 2220 100
rect 2214 95 2220 96
rect 2270 100 2276 101
rect 2270 96 2271 100
rect 2275 96 2276 100
rect 2270 95 2276 96
rect 2318 100 2324 101
rect 2318 96 2319 100
rect 2323 96 2324 100
rect 2318 95 2324 96
rect 2358 100 2364 101
rect 2358 96 2359 100
rect 2363 96 2364 100
rect 2358 95 2364 96
rect 2408 95 2410 102
rect 1238 94 1244 95
rect 1279 94 1283 95
rect 112 87 114 94
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 174 92 180 93
rect 174 88 175 92
rect 179 88 180 92
rect 174 87 180 88
rect 214 92 220 93
rect 214 88 215 92
rect 219 88 220 92
rect 214 87 220 88
rect 254 92 260 93
rect 254 88 255 92
rect 259 88 260 92
rect 254 87 260 88
rect 294 92 300 93
rect 294 88 295 92
rect 299 88 300 92
rect 294 87 300 88
rect 334 92 340 93
rect 334 88 335 92
rect 339 88 340 92
rect 334 87 340 88
rect 374 92 380 93
rect 374 88 375 92
rect 379 88 380 92
rect 374 87 380 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 526 92 532 93
rect 526 88 527 92
rect 531 88 532 92
rect 526 87 532 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 678 92 684 93
rect 678 88 679 92
rect 683 88 684 92
rect 678 87 684 88
rect 726 92 732 93
rect 726 88 727 92
rect 731 88 732 92
rect 726 87 732 88
rect 766 92 772 93
rect 766 88 767 92
rect 771 88 772 92
rect 766 87 772 88
rect 806 92 812 93
rect 806 88 807 92
rect 811 88 812 92
rect 806 87 812 88
rect 846 92 852 93
rect 846 88 847 92
rect 851 88 852 92
rect 846 87 852 88
rect 886 92 892 93
rect 886 88 887 92
rect 891 88 892 92
rect 886 87 892 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 974 92 980 93
rect 974 88 975 92
rect 979 88 980 92
rect 974 87 980 88
rect 1022 92 1028 93
rect 1022 88 1023 92
rect 1027 88 1028 92
rect 1022 87 1028 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
rect 1240 87 1242 94
rect 1279 89 1283 90
rect 1303 94 1307 95
rect 1303 89 1307 90
rect 1343 94 1347 95
rect 1343 89 1347 90
rect 1383 94 1387 95
rect 1383 89 1387 90
rect 1423 94 1427 95
rect 1423 89 1427 90
rect 1463 94 1467 95
rect 1463 89 1467 90
rect 1519 94 1523 95
rect 1519 89 1523 90
rect 1583 94 1587 95
rect 1583 89 1587 90
rect 1647 94 1651 95
rect 1647 89 1651 90
rect 1711 94 1715 95
rect 1711 89 1715 90
rect 1767 94 1771 95
rect 1767 89 1771 90
rect 1823 94 1827 95
rect 1823 89 1827 90
rect 1871 94 1875 95
rect 1871 89 1875 90
rect 1919 94 1923 95
rect 1919 89 1923 90
rect 1967 94 1971 95
rect 1967 89 1971 90
rect 2015 94 2019 95
rect 2015 89 2019 90
rect 2063 94 2067 95
rect 2063 89 2067 90
rect 2111 94 2115 95
rect 2111 89 2115 90
rect 2159 94 2163 95
rect 2159 89 2163 90
rect 2215 94 2219 95
rect 2215 89 2219 90
rect 2271 94 2275 95
rect 2271 89 2275 90
rect 2319 94 2323 95
rect 2319 89 2323 90
rect 2359 94 2363 95
rect 2359 89 2363 90
rect 2407 94 2411 95
rect 2407 89 2411 90
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 175 86 179 87
rect 175 81 179 82
rect 215 86 219 87
rect 215 81 219 82
rect 255 86 259 87
rect 255 81 259 82
rect 295 86 299 87
rect 295 81 299 82
rect 335 86 339 87
rect 335 81 339 82
rect 375 86 379 87
rect 375 81 379 82
rect 423 86 427 87
rect 423 81 427 82
rect 471 86 475 87
rect 471 81 475 82
rect 527 86 531 87
rect 527 81 531 82
rect 583 86 587 87
rect 583 81 587 82
rect 631 86 635 87
rect 631 81 635 82
rect 679 86 683 87
rect 679 81 683 82
rect 727 86 731 87
rect 727 81 731 82
rect 767 86 771 87
rect 767 81 771 82
rect 807 86 811 87
rect 807 81 811 82
rect 847 86 851 87
rect 847 81 851 82
rect 887 86 891 87
rect 887 81 891 82
rect 927 86 931 87
rect 927 81 931 82
rect 975 86 979 87
rect 975 81 979 82
rect 1023 86 1027 87
rect 1023 81 1027 82
rect 1071 86 1075 87
rect 1071 81 1075 82
rect 1111 86 1115 87
rect 1111 81 1115 82
rect 1151 86 1155 87
rect 1151 81 1155 82
rect 1191 86 1195 87
rect 1191 81 1195 82
rect 1239 86 1243 87
rect 1239 81 1243 82
<< m4c >>
rect 1279 2510 1283 2514
rect 1535 2510 1539 2514
rect 1575 2510 1579 2514
rect 1615 2510 1619 2514
rect 1655 2510 1659 2514
rect 1695 2510 1699 2514
rect 1735 2510 1739 2514
rect 1775 2510 1779 2514
rect 1815 2510 1819 2514
rect 1855 2510 1859 2514
rect 1895 2510 1899 2514
rect 1935 2510 1939 2514
rect 1975 2510 1979 2514
rect 2407 2510 2411 2514
rect 111 2498 115 2502
rect 135 2498 139 2502
rect 175 2498 179 2502
rect 215 2498 219 2502
rect 255 2498 259 2502
rect 311 2498 315 2502
rect 391 2498 395 2502
rect 479 2498 483 2502
rect 567 2498 571 2502
rect 655 2498 659 2502
rect 743 2498 747 2502
rect 831 2498 835 2502
rect 927 2498 931 2502
rect 1239 2498 1243 2502
rect 1279 2442 1283 2446
rect 1359 2442 1363 2446
rect 1399 2442 1403 2446
rect 1455 2442 1459 2446
rect 1519 2442 1523 2446
rect 1535 2442 1539 2446
rect 1575 2442 1579 2446
rect 1599 2442 1603 2446
rect 1615 2442 1619 2446
rect 1655 2442 1659 2446
rect 1679 2442 1683 2446
rect 1695 2442 1699 2446
rect 1735 2442 1739 2446
rect 1759 2442 1763 2446
rect 1775 2442 1779 2446
rect 1815 2442 1819 2446
rect 1839 2442 1843 2446
rect 1855 2442 1859 2446
rect 1895 2442 1899 2446
rect 1919 2442 1923 2446
rect 1935 2442 1939 2446
rect 1975 2442 1979 2446
rect 1999 2442 2003 2446
rect 2079 2442 2083 2446
rect 2159 2442 2163 2446
rect 2247 2442 2251 2446
rect 2335 2442 2339 2446
rect 2407 2442 2411 2446
rect 111 2430 115 2434
rect 135 2430 139 2434
rect 175 2430 179 2434
rect 183 2430 187 2434
rect 215 2430 219 2434
rect 247 2430 251 2434
rect 255 2430 259 2434
rect 311 2430 315 2434
rect 319 2430 323 2434
rect 391 2430 395 2434
rect 471 2430 475 2434
rect 479 2430 483 2434
rect 543 2430 547 2434
rect 567 2430 571 2434
rect 615 2430 619 2434
rect 655 2430 659 2434
rect 679 2430 683 2434
rect 735 2430 739 2434
rect 743 2430 747 2434
rect 791 2430 795 2434
rect 831 2430 835 2434
rect 839 2430 843 2434
rect 887 2430 891 2434
rect 927 2430 931 2434
rect 935 2430 939 2434
rect 991 2430 995 2434
rect 1047 2430 1051 2434
rect 1239 2430 1243 2434
rect 1279 2374 1283 2378
rect 1359 2374 1363 2378
rect 1399 2374 1403 2378
rect 1407 2374 1411 2378
rect 1455 2374 1459 2378
rect 1471 2374 1475 2378
rect 1519 2374 1523 2378
rect 1543 2374 1547 2378
rect 1599 2374 1603 2378
rect 1615 2374 1619 2378
rect 1679 2374 1683 2378
rect 1695 2374 1699 2378
rect 1759 2374 1763 2378
rect 1775 2374 1779 2378
rect 1839 2374 1843 2378
rect 1855 2374 1859 2378
rect 1919 2374 1923 2378
rect 1927 2374 1931 2378
rect 1999 2374 2003 2378
rect 2071 2374 2075 2378
rect 2079 2374 2083 2378
rect 2143 2374 2147 2378
rect 2159 2374 2163 2378
rect 2223 2374 2227 2378
rect 2247 2374 2251 2378
rect 2303 2374 2307 2378
rect 2335 2374 2339 2378
rect 2359 2374 2363 2378
rect 2407 2374 2411 2378
rect 111 2354 115 2358
rect 135 2354 139 2358
rect 175 2354 179 2358
rect 183 2354 187 2358
rect 215 2354 219 2358
rect 247 2354 251 2358
rect 271 2354 275 2358
rect 319 2354 323 2358
rect 351 2354 355 2358
rect 391 2354 395 2358
rect 431 2354 435 2358
rect 471 2354 475 2358
rect 519 2354 523 2358
rect 543 2354 547 2358
rect 599 2354 603 2358
rect 615 2354 619 2358
rect 679 2354 683 2358
rect 735 2354 739 2358
rect 751 2354 755 2358
rect 791 2354 795 2358
rect 823 2354 827 2358
rect 839 2354 843 2358
rect 887 2354 891 2358
rect 935 2354 939 2358
rect 959 2354 963 2358
rect 991 2354 995 2358
rect 1031 2354 1035 2358
rect 1047 2354 1051 2358
rect 1239 2354 1243 2358
rect 1279 2302 1283 2306
rect 1359 2302 1363 2306
rect 1407 2302 1411 2306
rect 1471 2302 1475 2306
rect 1503 2302 1507 2306
rect 1543 2302 1547 2306
rect 1583 2302 1587 2306
rect 1615 2302 1619 2306
rect 1623 2302 1627 2306
rect 1663 2302 1667 2306
rect 1695 2302 1699 2306
rect 1703 2302 1707 2306
rect 1759 2302 1763 2306
rect 1775 2302 1779 2306
rect 1823 2302 1827 2306
rect 1855 2302 1859 2306
rect 1895 2302 1899 2306
rect 1927 2302 1931 2306
rect 1967 2302 1971 2306
rect 1999 2302 2003 2306
rect 2047 2302 2051 2306
rect 2071 2302 2075 2306
rect 2127 2302 2131 2306
rect 2143 2302 2147 2306
rect 2207 2302 2211 2306
rect 2223 2302 2227 2306
rect 2295 2302 2299 2306
rect 2303 2302 2307 2306
rect 2359 2302 2363 2306
rect 2407 2302 2411 2306
rect 111 2282 115 2286
rect 135 2282 139 2286
rect 175 2282 179 2286
rect 215 2282 219 2286
rect 231 2282 235 2286
rect 271 2282 275 2286
rect 303 2282 307 2286
rect 351 2282 355 2286
rect 375 2282 379 2286
rect 431 2282 435 2286
rect 455 2282 459 2286
rect 519 2282 523 2286
rect 535 2282 539 2286
rect 599 2282 603 2286
rect 615 2282 619 2286
rect 679 2282 683 2286
rect 687 2282 691 2286
rect 751 2282 755 2286
rect 759 2282 763 2286
rect 823 2282 827 2286
rect 831 2282 835 2286
rect 887 2282 891 2286
rect 911 2282 915 2286
rect 959 2282 963 2286
rect 991 2282 995 2286
rect 1031 2282 1035 2286
rect 1239 2282 1243 2286
rect 1279 2226 1283 2230
rect 1303 2226 1307 2230
rect 1343 2226 1347 2230
rect 1383 2226 1387 2230
rect 1431 2226 1435 2230
rect 1495 2226 1499 2230
rect 1503 2226 1507 2230
rect 1543 2226 1547 2230
rect 1567 2226 1571 2230
rect 1583 2226 1587 2230
rect 1623 2226 1627 2230
rect 1639 2226 1643 2230
rect 1663 2226 1667 2230
rect 1703 2226 1707 2230
rect 1711 2226 1715 2230
rect 1759 2226 1763 2230
rect 1783 2226 1787 2230
rect 1823 2226 1827 2230
rect 1855 2226 1859 2230
rect 1895 2226 1899 2230
rect 1935 2226 1939 2230
rect 1967 2226 1971 2230
rect 2015 2226 2019 2230
rect 2047 2226 2051 2230
rect 2095 2226 2099 2230
rect 2127 2226 2131 2230
rect 2183 2226 2187 2230
rect 2207 2226 2211 2230
rect 2279 2226 2283 2230
rect 2295 2226 2299 2230
rect 2359 2226 2363 2230
rect 2407 2226 2411 2230
rect 111 2214 115 2218
rect 135 2214 139 2218
rect 175 2214 179 2218
rect 231 2214 235 2218
rect 247 2214 251 2218
rect 287 2214 291 2218
rect 303 2214 307 2218
rect 327 2214 331 2218
rect 375 2214 379 2218
rect 431 2214 435 2218
rect 455 2214 459 2218
rect 495 2214 499 2218
rect 535 2214 539 2218
rect 551 2214 555 2218
rect 607 2214 611 2218
rect 615 2214 619 2218
rect 663 2214 667 2218
rect 687 2214 691 2218
rect 719 2214 723 2218
rect 759 2214 763 2218
rect 783 2214 787 2218
rect 831 2214 835 2218
rect 847 2214 851 2218
rect 911 2214 915 2218
rect 991 2214 995 2218
rect 1239 2214 1243 2218
rect 1279 2158 1283 2162
rect 1303 2158 1307 2162
rect 1343 2158 1347 2162
rect 1351 2158 1355 2162
rect 1383 2158 1387 2162
rect 1431 2158 1435 2162
rect 1439 2158 1443 2162
rect 1495 2158 1499 2162
rect 1535 2158 1539 2162
rect 1567 2158 1571 2162
rect 1631 2158 1635 2162
rect 1639 2158 1643 2162
rect 1711 2158 1715 2162
rect 1727 2158 1731 2162
rect 1783 2158 1787 2162
rect 1815 2158 1819 2162
rect 1855 2158 1859 2162
rect 1895 2158 1899 2162
rect 1935 2158 1939 2162
rect 1975 2158 1979 2162
rect 2015 2158 2019 2162
rect 2047 2158 2051 2162
rect 2095 2158 2099 2162
rect 2111 2158 2115 2162
rect 2175 2158 2179 2162
rect 2183 2158 2187 2162
rect 2239 2158 2243 2162
rect 2279 2158 2283 2162
rect 2311 2158 2315 2162
rect 2359 2158 2363 2162
rect 2407 2158 2411 2162
rect 111 2138 115 2142
rect 247 2138 251 2142
rect 287 2138 291 2142
rect 327 2138 331 2142
rect 375 2138 379 2142
rect 383 2138 387 2142
rect 423 2138 427 2142
rect 431 2138 435 2142
rect 463 2138 467 2142
rect 495 2138 499 2142
rect 503 2138 507 2142
rect 551 2138 555 2142
rect 607 2138 611 2142
rect 663 2138 667 2142
rect 719 2138 723 2142
rect 727 2138 731 2142
rect 783 2138 787 2142
rect 791 2138 795 2142
rect 847 2138 851 2142
rect 855 2138 859 2142
rect 911 2138 915 2142
rect 967 2138 971 2142
rect 1023 2138 1027 2142
rect 1079 2138 1083 2142
rect 1143 2138 1147 2142
rect 1239 2138 1243 2142
rect 1279 2086 1283 2090
rect 1303 2086 1307 2090
rect 1343 2086 1347 2090
rect 1351 2086 1355 2090
rect 1399 2086 1403 2090
rect 1439 2086 1443 2090
rect 1479 2086 1483 2090
rect 1535 2086 1539 2090
rect 1567 2086 1571 2090
rect 1631 2086 1635 2090
rect 1663 2086 1667 2090
rect 1727 2086 1731 2090
rect 1759 2086 1763 2090
rect 1815 2086 1819 2090
rect 1847 2086 1851 2090
rect 1895 2086 1899 2090
rect 1935 2086 1939 2090
rect 1975 2086 1979 2090
rect 2015 2086 2019 2090
rect 2047 2086 2051 2090
rect 2095 2086 2099 2090
rect 2111 2086 2115 2090
rect 2167 2086 2171 2090
rect 2175 2086 2179 2090
rect 2239 2086 2243 2090
rect 2311 2086 2315 2090
rect 2359 2086 2363 2090
rect 2407 2086 2411 2090
rect 111 2070 115 2074
rect 383 2070 387 2074
rect 423 2070 427 2074
rect 463 2070 467 2074
rect 503 2070 507 2074
rect 543 2070 547 2074
rect 551 2070 555 2074
rect 583 2070 587 2074
rect 607 2070 611 2074
rect 631 2070 635 2074
rect 663 2070 667 2074
rect 687 2070 691 2074
rect 727 2070 731 2074
rect 743 2070 747 2074
rect 791 2070 795 2074
rect 799 2070 803 2074
rect 847 2070 851 2074
rect 855 2070 859 2074
rect 903 2070 907 2074
rect 911 2070 915 2074
rect 959 2070 963 2074
rect 967 2070 971 2074
rect 1015 2070 1019 2074
rect 1023 2070 1027 2074
rect 1071 2070 1075 2074
rect 1079 2070 1083 2074
rect 1143 2070 1147 2074
rect 1239 2070 1243 2074
rect 1279 2010 1283 2014
rect 1303 2010 1307 2014
rect 1343 2010 1347 2014
rect 1351 2010 1355 2014
rect 1399 2010 1403 2014
rect 1423 2010 1427 2014
rect 1479 2010 1483 2014
rect 1495 2010 1499 2014
rect 1567 2010 1571 2014
rect 1575 2010 1579 2014
rect 1663 2010 1667 2014
rect 1751 2010 1755 2014
rect 1759 2010 1763 2014
rect 1839 2010 1843 2014
rect 1847 2010 1851 2014
rect 1919 2010 1923 2014
rect 1935 2010 1939 2014
rect 1999 2010 2003 2014
rect 2015 2010 2019 2014
rect 2071 2010 2075 2014
rect 2095 2010 2099 2014
rect 2135 2010 2139 2014
rect 2167 2010 2171 2014
rect 2191 2010 2195 2014
rect 2239 2010 2243 2014
rect 2255 2010 2259 2014
rect 2311 2010 2315 2014
rect 2319 2010 2323 2014
rect 2359 2010 2363 2014
rect 2407 2010 2411 2014
rect 111 1994 115 1998
rect 367 1994 371 1998
rect 383 1994 387 1998
rect 407 1994 411 1998
rect 423 1994 427 1998
rect 455 1994 459 1998
rect 463 1994 467 1998
rect 503 1994 507 1998
rect 511 1994 515 1998
rect 543 1994 547 1998
rect 567 1994 571 1998
rect 583 1994 587 1998
rect 631 1994 635 1998
rect 687 1994 691 1998
rect 695 1994 699 1998
rect 743 1994 747 1998
rect 759 1994 763 1998
rect 799 1994 803 1998
rect 815 1994 819 1998
rect 847 1994 851 1998
rect 871 1994 875 1998
rect 903 1994 907 1998
rect 935 1994 939 1998
rect 959 1994 963 1998
rect 999 1994 1003 1998
rect 1015 1994 1019 1998
rect 1063 1994 1067 1998
rect 1071 1994 1075 1998
rect 1239 1994 1243 1998
rect 1279 1942 1283 1946
rect 1303 1942 1307 1946
rect 1351 1942 1355 1946
rect 1359 1942 1363 1946
rect 1423 1942 1427 1946
rect 1447 1942 1451 1946
rect 1495 1942 1499 1946
rect 1535 1942 1539 1946
rect 1575 1942 1579 1946
rect 1623 1942 1627 1946
rect 1663 1942 1667 1946
rect 1711 1942 1715 1946
rect 1751 1942 1755 1946
rect 1791 1942 1795 1946
rect 1839 1942 1843 1946
rect 1863 1942 1867 1946
rect 1919 1942 1923 1946
rect 1935 1942 1939 1946
rect 1999 1942 2003 1946
rect 2007 1942 2011 1946
rect 2071 1942 2075 1946
rect 2079 1942 2083 1946
rect 2135 1942 2139 1946
rect 2151 1942 2155 1946
rect 2191 1942 2195 1946
rect 2223 1942 2227 1946
rect 2255 1942 2259 1946
rect 2303 1942 2307 1946
rect 2319 1942 2323 1946
rect 2359 1942 2363 1946
rect 2407 1942 2411 1946
rect 111 1922 115 1926
rect 175 1922 179 1926
rect 215 1922 219 1926
rect 263 1922 267 1926
rect 319 1922 323 1926
rect 367 1922 371 1926
rect 391 1922 395 1926
rect 407 1922 411 1926
rect 455 1922 459 1926
rect 471 1922 475 1926
rect 511 1922 515 1926
rect 551 1922 555 1926
rect 567 1922 571 1926
rect 631 1922 635 1926
rect 639 1922 643 1926
rect 695 1922 699 1926
rect 719 1922 723 1926
rect 759 1922 763 1926
rect 799 1922 803 1926
rect 815 1922 819 1926
rect 871 1922 875 1926
rect 879 1922 883 1926
rect 935 1922 939 1926
rect 959 1922 963 1926
rect 999 1922 1003 1926
rect 1039 1922 1043 1926
rect 1063 1922 1067 1926
rect 1119 1922 1123 1926
rect 1239 1922 1243 1926
rect 1279 1874 1283 1878
rect 1303 1874 1307 1878
rect 1311 1874 1315 1878
rect 1359 1874 1363 1878
rect 1415 1874 1419 1878
rect 1447 1874 1451 1878
rect 1479 1874 1483 1878
rect 1535 1874 1539 1878
rect 1543 1874 1547 1878
rect 1615 1874 1619 1878
rect 1623 1874 1627 1878
rect 1687 1874 1691 1878
rect 1711 1874 1715 1878
rect 1767 1874 1771 1878
rect 1791 1874 1795 1878
rect 1863 1874 1867 1878
rect 1935 1874 1939 1878
rect 1975 1874 1979 1878
rect 2007 1874 2011 1878
rect 2079 1874 2083 1878
rect 2095 1874 2099 1878
rect 2151 1874 2155 1878
rect 2223 1874 2227 1878
rect 2303 1874 2307 1878
rect 2359 1874 2363 1878
rect 2407 1874 2411 1878
rect 111 1846 115 1850
rect 135 1846 139 1850
rect 175 1846 179 1850
rect 215 1846 219 1850
rect 263 1846 267 1850
rect 271 1846 275 1850
rect 319 1846 323 1850
rect 351 1846 355 1850
rect 391 1846 395 1850
rect 439 1846 443 1850
rect 471 1846 475 1850
rect 535 1846 539 1850
rect 551 1846 555 1850
rect 631 1846 635 1850
rect 639 1846 643 1850
rect 719 1846 723 1850
rect 727 1846 731 1850
rect 799 1846 803 1850
rect 823 1846 827 1850
rect 879 1846 883 1850
rect 911 1846 915 1850
rect 959 1846 963 1850
rect 991 1846 995 1850
rect 1039 1846 1043 1850
rect 1063 1846 1067 1850
rect 1119 1846 1123 1850
rect 1135 1846 1139 1850
rect 1191 1846 1195 1850
rect 1239 1846 1243 1850
rect 1279 1802 1283 1806
rect 1311 1802 1315 1806
rect 1359 1802 1363 1806
rect 1407 1802 1411 1806
rect 1415 1802 1419 1806
rect 1471 1802 1475 1806
rect 1479 1802 1483 1806
rect 1535 1802 1539 1806
rect 1543 1802 1547 1806
rect 1599 1802 1603 1806
rect 1615 1802 1619 1806
rect 1663 1802 1667 1806
rect 1687 1802 1691 1806
rect 1727 1802 1731 1806
rect 1767 1802 1771 1806
rect 1783 1802 1787 1806
rect 1839 1802 1843 1806
rect 1863 1802 1867 1806
rect 1895 1802 1899 1806
rect 1959 1802 1963 1806
rect 1975 1802 1979 1806
rect 2095 1802 2099 1806
rect 2223 1802 2227 1806
rect 2359 1802 2363 1806
rect 2407 1802 2411 1806
rect 111 1778 115 1782
rect 135 1778 139 1782
rect 175 1778 179 1782
rect 215 1778 219 1782
rect 271 1778 275 1782
rect 287 1778 291 1782
rect 351 1778 355 1782
rect 375 1778 379 1782
rect 439 1778 443 1782
rect 471 1778 475 1782
rect 535 1778 539 1782
rect 567 1778 571 1782
rect 631 1778 635 1782
rect 663 1778 667 1782
rect 727 1778 731 1782
rect 751 1778 755 1782
rect 823 1778 827 1782
rect 831 1778 835 1782
rect 903 1778 907 1782
rect 911 1778 915 1782
rect 967 1778 971 1782
rect 991 1778 995 1782
rect 1031 1778 1035 1782
rect 1063 1778 1067 1782
rect 1087 1778 1091 1782
rect 1135 1778 1139 1782
rect 1151 1778 1155 1782
rect 1191 1778 1195 1782
rect 1239 1778 1243 1782
rect 1279 1734 1283 1738
rect 1303 1734 1307 1738
rect 1351 1734 1355 1738
rect 1407 1734 1411 1738
rect 1423 1734 1427 1738
rect 1471 1734 1475 1738
rect 1503 1734 1507 1738
rect 1535 1734 1539 1738
rect 1583 1734 1587 1738
rect 1599 1734 1603 1738
rect 1663 1734 1667 1738
rect 1727 1734 1731 1738
rect 1735 1734 1739 1738
rect 1783 1734 1787 1738
rect 1807 1734 1811 1738
rect 1839 1734 1843 1738
rect 1871 1734 1875 1738
rect 1895 1734 1899 1738
rect 1935 1734 1939 1738
rect 1959 1734 1963 1738
rect 1999 1734 2003 1738
rect 2063 1734 2067 1738
rect 2407 1734 2411 1738
rect 111 1706 115 1710
rect 135 1706 139 1710
rect 175 1706 179 1710
rect 215 1706 219 1710
rect 239 1706 243 1710
rect 287 1706 291 1710
rect 319 1706 323 1710
rect 375 1706 379 1710
rect 415 1706 419 1710
rect 471 1706 475 1710
rect 511 1706 515 1710
rect 567 1706 571 1710
rect 615 1706 619 1710
rect 663 1706 667 1710
rect 711 1706 715 1710
rect 751 1706 755 1710
rect 799 1706 803 1710
rect 831 1706 835 1710
rect 879 1706 883 1710
rect 903 1706 907 1710
rect 951 1706 955 1710
rect 967 1706 971 1710
rect 1015 1706 1019 1710
rect 1031 1706 1035 1710
rect 1087 1706 1091 1710
rect 1151 1706 1155 1710
rect 1159 1706 1163 1710
rect 1191 1706 1195 1710
rect 1239 1706 1243 1710
rect 1279 1666 1283 1670
rect 1303 1666 1307 1670
rect 1351 1666 1355 1670
rect 1359 1666 1363 1670
rect 1423 1666 1427 1670
rect 1447 1666 1451 1670
rect 1503 1666 1507 1670
rect 1543 1666 1547 1670
rect 1583 1666 1587 1670
rect 1639 1666 1643 1670
rect 1663 1666 1667 1670
rect 1727 1666 1731 1670
rect 1735 1666 1739 1670
rect 1807 1666 1811 1670
rect 1815 1666 1819 1670
rect 1871 1666 1875 1670
rect 1895 1666 1899 1670
rect 1935 1666 1939 1670
rect 1967 1666 1971 1670
rect 1999 1666 2003 1670
rect 2031 1666 2035 1670
rect 2063 1666 2067 1670
rect 2095 1666 2099 1670
rect 2159 1666 2163 1670
rect 2223 1666 2227 1670
rect 2407 1666 2411 1670
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 175 1634 179 1638
rect 239 1634 243 1638
rect 271 1634 275 1638
rect 311 1634 315 1638
rect 319 1634 323 1638
rect 359 1634 363 1638
rect 415 1634 419 1638
rect 471 1634 475 1638
rect 511 1634 515 1638
rect 535 1634 539 1638
rect 599 1634 603 1638
rect 615 1634 619 1638
rect 663 1634 667 1638
rect 711 1634 715 1638
rect 719 1634 723 1638
rect 775 1634 779 1638
rect 799 1634 803 1638
rect 831 1634 835 1638
rect 879 1634 883 1638
rect 887 1634 891 1638
rect 943 1634 947 1638
rect 951 1634 955 1638
rect 999 1634 1003 1638
rect 1015 1634 1019 1638
rect 1087 1634 1091 1638
rect 1159 1634 1163 1638
rect 1239 1634 1243 1638
rect 1279 1598 1283 1602
rect 1303 1598 1307 1602
rect 1327 1598 1331 1602
rect 1359 1598 1363 1602
rect 1399 1598 1403 1602
rect 1447 1598 1451 1602
rect 1479 1598 1483 1602
rect 1543 1598 1547 1602
rect 1567 1598 1571 1602
rect 1639 1598 1643 1602
rect 1655 1598 1659 1602
rect 1727 1598 1731 1602
rect 1743 1598 1747 1602
rect 1815 1598 1819 1602
rect 1831 1598 1835 1602
rect 1895 1598 1899 1602
rect 1911 1598 1915 1602
rect 1967 1598 1971 1602
rect 1983 1598 1987 1602
rect 2031 1598 2035 1602
rect 2047 1598 2051 1602
rect 2095 1598 2099 1602
rect 2111 1598 2115 1602
rect 2159 1598 2163 1602
rect 2167 1598 2171 1602
rect 2215 1598 2219 1602
rect 2223 1598 2227 1602
rect 2271 1598 2275 1602
rect 2319 1598 2323 1602
rect 2359 1598 2363 1602
rect 2407 1598 2411 1602
rect 111 1558 115 1562
rect 271 1558 275 1562
rect 311 1558 315 1562
rect 327 1558 331 1562
rect 359 1558 363 1562
rect 367 1558 371 1562
rect 407 1558 411 1562
rect 415 1558 419 1562
rect 447 1558 451 1562
rect 471 1558 475 1562
rect 487 1558 491 1562
rect 527 1558 531 1562
rect 535 1558 539 1562
rect 567 1558 571 1562
rect 599 1558 603 1562
rect 607 1558 611 1562
rect 647 1558 651 1562
rect 663 1558 667 1562
rect 687 1558 691 1562
rect 719 1558 723 1562
rect 727 1558 731 1562
rect 767 1558 771 1562
rect 775 1558 779 1562
rect 807 1558 811 1562
rect 831 1558 835 1562
rect 847 1558 851 1562
rect 887 1558 891 1562
rect 927 1558 931 1562
rect 943 1558 947 1562
rect 999 1558 1003 1562
rect 1239 1558 1243 1562
rect 1279 1526 1283 1530
rect 1327 1526 1331 1530
rect 1335 1526 1339 1530
rect 1399 1526 1403 1530
rect 1415 1526 1419 1530
rect 1479 1526 1483 1530
rect 1503 1526 1507 1530
rect 1567 1526 1571 1530
rect 1615 1526 1619 1530
rect 1655 1526 1659 1530
rect 1743 1526 1747 1530
rect 1831 1526 1835 1530
rect 1887 1526 1891 1530
rect 1911 1526 1915 1530
rect 1983 1526 1987 1530
rect 2047 1526 2051 1530
rect 2111 1526 2115 1530
rect 2167 1526 2171 1530
rect 2215 1526 2219 1530
rect 2271 1526 2275 1530
rect 2319 1526 2323 1530
rect 2359 1526 2363 1530
rect 2407 1526 2411 1530
rect 1279 1458 1283 1462
rect 1335 1458 1339 1462
rect 1375 1458 1379 1462
rect 1415 1458 1419 1462
rect 1463 1458 1467 1462
rect 1503 1458 1507 1462
rect 1551 1458 1555 1462
rect 1615 1458 1619 1462
rect 1639 1458 1643 1462
rect 1727 1458 1731 1462
rect 1743 1458 1747 1462
rect 1807 1458 1811 1462
rect 1879 1458 1883 1462
rect 1887 1458 1891 1462
rect 1943 1458 1947 1462
rect 1999 1458 2003 1462
rect 2047 1458 2051 1462
rect 2095 1458 2099 1462
rect 2143 1458 2147 1462
rect 2191 1458 2195 1462
rect 2215 1458 2219 1462
rect 2239 1458 2243 1462
rect 2279 1458 2283 1462
rect 2319 1458 2323 1462
rect 2359 1458 2363 1462
rect 2407 1458 2411 1462
rect 111 1450 115 1454
rect 143 1450 147 1454
rect 183 1450 187 1454
rect 223 1450 227 1454
rect 263 1450 267 1454
rect 319 1450 323 1454
rect 327 1450 331 1454
rect 367 1450 371 1454
rect 391 1450 395 1454
rect 407 1450 411 1454
rect 447 1450 451 1454
rect 471 1450 475 1454
rect 487 1450 491 1454
rect 527 1450 531 1454
rect 559 1450 563 1454
rect 567 1450 571 1454
rect 607 1450 611 1454
rect 647 1450 651 1454
rect 687 1450 691 1454
rect 727 1450 731 1454
rect 767 1450 771 1454
rect 807 1450 811 1454
rect 847 1450 851 1454
rect 879 1450 883 1454
rect 887 1450 891 1454
rect 927 1450 931 1454
rect 943 1450 947 1454
rect 999 1450 1003 1454
rect 1047 1450 1051 1454
rect 1103 1450 1107 1454
rect 1151 1450 1155 1454
rect 1191 1450 1195 1454
rect 1239 1450 1243 1454
rect 111 1382 115 1386
rect 143 1382 147 1386
rect 167 1382 171 1386
rect 183 1382 187 1386
rect 207 1382 211 1386
rect 223 1382 227 1386
rect 247 1382 251 1386
rect 263 1382 267 1386
rect 303 1382 307 1386
rect 319 1382 323 1386
rect 367 1382 371 1386
rect 391 1382 395 1386
rect 439 1382 443 1386
rect 471 1382 475 1386
rect 519 1382 523 1386
rect 559 1382 563 1386
rect 599 1382 603 1386
rect 647 1382 651 1386
rect 679 1382 683 1386
rect 727 1382 731 1386
rect 751 1382 755 1386
rect 807 1382 811 1386
rect 823 1382 827 1386
rect 879 1382 883 1386
rect 887 1382 891 1386
rect 943 1382 947 1386
rect 951 1382 955 1386
rect 999 1382 1003 1386
rect 1015 1382 1019 1386
rect 1047 1382 1051 1386
rect 1079 1382 1083 1386
rect 1103 1382 1107 1386
rect 1143 1382 1147 1386
rect 1151 1382 1155 1386
rect 1191 1382 1195 1386
rect 1239 1382 1243 1386
rect 1279 1382 1283 1386
rect 1303 1382 1307 1386
rect 1343 1382 1347 1386
rect 1375 1382 1379 1386
rect 1399 1382 1403 1386
rect 1463 1382 1467 1386
rect 1535 1382 1539 1386
rect 1551 1382 1555 1386
rect 1607 1382 1611 1386
rect 1639 1382 1643 1386
rect 1687 1382 1691 1386
rect 1727 1382 1731 1386
rect 1767 1382 1771 1386
rect 1807 1382 1811 1386
rect 1847 1382 1851 1386
rect 1879 1382 1883 1386
rect 1935 1382 1939 1386
rect 1943 1382 1947 1386
rect 1999 1382 2003 1386
rect 2023 1382 2027 1386
rect 2047 1382 2051 1386
rect 2095 1382 2099 1386
rect 2111 1382 2115 1386
rect 2143 1382 2147 1386
rect 2191 1382 2195 1386
rect 2199 1382 2203 1386
rect 2239 1382 2243 1386
rect 2279 1382 2283 1386
rect 2287 1382 2291 1386
rect 2319 1382 2323 1386
rect 2359 1382 2363 1386
rect 2407 1382 2411 1386
rect 111 1310 115 1314
rect 167 1310 171 1314
rect 183 1310 187 1314
rect 207 1310 211 1314
rect 231 1310 235 1314
rect 247 1310 251 1314
rect 287 1310 291 1314
rect 303 1310 307 1314
rect 351 1310 355 1314
rect 367 1310 371 1314
rect 423 1310 427 1314
rect 439 1310 443 1314
rect 495 1310 499 1314
rect 519 1310 523 1314
rect 567 1310 571 1314
rect 599 1310 603 1314
rect 639 1310 643 1314
rect 679 1310 683 1314
rect 703 1310 707 1314
rect 751 1310 755 1314
rect 767 1310 771 1314
rect 823 1310 827 1314
rect 879 1310 883 1314
rect 887 1310 891 1314
rect 935 1310 939 1314
rect 951 1310 955 1314
rect 999 1310 1003 1314
rect 1015 1310 1019 1314
rect 1079 1310 1083 1314
rect 1143 1310 1147 1314
rect 1191 1310 1195 1314
rect 1239 1310 1243 1314
rect 1279 1314 1283 1318
rect 1303 1314 1307 1318
rect 1343 1314 1347 1318
rect 1383 1314 1387 1318
rect 1399 1314 1403 1318
rect 1423 1314 1427 1318
rect 1463 1314 1467 1318
rect 1503 1314 1507 1318
rect 1535 1314 1539 1318
rect 1543 1314 1547 1318
rect 1583 1314 1587 1318
rect 1607 1314 1611 1318
rect 1623 1314 1627 1318
rect 1679 1314 1683 1318
rect 1687 1314 1691 1318
rect 1735 1314 1739 1318
rect 1767 1314 1771 1318
rect 1791 1314 1795 1318
rect 1847 1314 1851 1318
rect 1903 1314 1907 1318
rect 1935 1314 1939 1318
rect 1967 1314 1971 1318
rect 2023 1314 2027 1318
rect 2039 1314 2043 1318
rect 2111 1314 2115 1318
rect 2119 1314 2123 1318
rect 2199 1314 2203 1318
rect 2287 1314 2291 1318
rect 2359 1314 2363 1318
rect 2407 1314 2411 1318
rect 111 1238 115 1242
rect 135 1238 139 1242
rect 175 1238 179 1242
rect 183 1238 187 1242
rect 231 1238 235 1242
rect 287 1238 291 1242
rect 311 1238 315 1242
rect 351 1238 355 1242
rect 399 1238 403 1242
rect 423 1238 427 1242
rect 487 1238 491 1242
rect 495 1238 499 1242
rect 567 1238 571 1242
rect 575 1238 579 1242
rect 639 1238 643 1242
rect 663 1238 667 1242
rect 703 1238 707 1242
rect 743 1238 747 1242
rect 767 1238 771 1242
rect 815 1238 819 1242
rect 823 1238 827 1242
rect 879 1238 883 1242
rect 935 1238 939 1242
rect 943 1238 947 1242
rect 999 1238 1003 1242
rect 1007 1238 1011 1242
rect 1071 1238 1075 1242
rect 1239 1238 1243 1242
rect 1279 1238 1283 1242
rect 1303 1238 1307 1242
rect 1343 1238 1347 1242
rect 1375 1238 1379 1242
rect 1383 1238 1387 1242
rect 1423 1238 1427 1242
rect 1463 1238 1467 1242
rect 1479 1238 1483 1242
rect 1503 1238 1507 1242
rect 1543 1238 1547 1242
rect 1583 1238 1587 1242
rect 1623 1238 1627 1242
rect 1679 1238 1683 1242
rect 1687 1238 1691 1242
rect 1735 1238 1739 1242
rect 1791 1238 1795 1242
rect 1847 1238 1851 1242
rect 1887 1238 1891 1242
rect 1903 1238 1907 1242
rect 1967 1238 1971 1242
rect 1983 1238 1987 1242
rect 2039 1238 2043 1242
rect 2071 1238 2075 1242
rect 2119 1238 2123 1242
rect 2151 1238 2155 1242
rect 2199 1238 2203 1242
rect 2223 1238 2227 1242
rect 2287 1238 2291 1242
rect 2303 1238 2307 1242
rect 2359 1238 2363 1242
rect 2407 1238 2411 1242
rect 111 1170 115 1174
rect 135 1170 139 1174
rect 175 1170 179 1174
rect 231 1170 235 1174
rect 239 1170 243 1174
rect 311 1170 315 1174
rect 327 1170 331 1174
rect 399 1170 403 1174
rect 431 1170 435 1174
rect 487 1170 491 1174
rect 535 1170 539 1174
rect 575 1170 579 1174
rect 639 1170 643 1174
rect 663 1170 667 1174
rect 743 1170 747 1174
rect 815 1170 819 1174
rect 839 1170 843 1174
rect 879 1170 883 1174
rect 919 1170 923 1174
rect 943 1170 947 1174
rect 999 1170 1003 1174
rect 1007 1170 1011 1174
rect 1071 1170 1075 1174
rect 1143 1170 1147 1174
rect 1191 1170 1195 1174
rect 1239 1170 1243 1174
rect 1279 1170 1283 1174
rect 1303 1170 1307 1174
rect 1343 1170 1347 1174
rect 1375 1170 1379 1174
rect 1407 1170 1411 1174
rect 1479 1170 1483 1174
rect 1487 1170 1491 1174
rect 1583 1170 1587 1174
rect 1687 1170 1691 1174
rect 1791 1170 1795 1174
rect 1799 1170 1803 1174
rect 1887 1170 1891 1174
rect 1903 1170 1907 1174
rect 1983 1170 1987 1174
rect 1999 1170 2003 1174
rect 2071 1170 2075 1174
rect 2079 1170 2083 1174
rect 2151 1170 2155 1174
rect 2159 1170 2163 1174
rect 2223 1170 2227 1174
rect 2231 1170 2235 1174
rect 2303 1170 2307 1174
rect 2359 1170 2363 1174
rect 2407 1170 2411 1174
rect 111 1098 115 1102
rect 135 1098 139 1102
rect 175 1098 179 1102
rect 239 1098 243 1102
rect 247 1098 251 1102
rect 327 1098 331 1102
rect 415 1098 419 1102
rect 431 1098 435 1102
rect 503 1098 507 1102
rect 535 1098 539 1102
rect 583 1098 587 1102
rect 639 1098 643 1102
rect 663 1098 667 1102
rect 735 1098 739 1102
rect 743 1098 747 1102
rect 799 1098 803 1102
rect 839 1098 843 1102
rect 863 1098 867 1102
rect 919 1098 923 1102
rect 983 1098 987 1102
rect 999 1098 1003 1102
rect 1047 1098 1051 1102
rect 1071 1098 1075 1102
rect 1143 1098 1147 1102
rect 1191 1098 1195 1102
rect 1239 1098 1243 1102
rect 1279 1102 1283 1106
rect 1303 1102 1307 1106
rect 1343 1102 1347 1106
rect 1407 1102 1411 1106
rect 1431 1102 1435 1106
rect 1471 1102 1475 1106
rect 1487 1102 1491 1106
rect 1511 1102 1515 1106
rect 1559 1102 1563 1106
rect 1583 1102 1587 1106
rect 1615 1102 1619 1106
rect 1671 1102 1675 1106
rect 1687 1102 1691 1106
rect 1727 1102 1731 1106
rect 1775 1102 1779 1106
rect 1799 1102 1803 1106
rect 1823 1102 1827 1106
rect 1871 1102 1875 1106
rect 1903 1102 1907 1106
rect 1919 1102 1923 1106
rect 1967 1102 1971 1106
rect 1999 1102 2003 1106
rect 2015 1102 2019 1106
rect 2063 1102 2067 1106
rect 2079 1102 2083 1106
rect 2119 1102 2123 1106
rect 2159 1102 2163 1106
rect 2175 1102 2179 1106
rect 2231 1102 2235 1106
rect 2303 1102 2307 1106
rect 2359 1102 2363 1106
rect 2407 1102 2411 1106
rect 111 1030 115 1034
rect 135 1030 139 1034
rect 175 1030 179 1034
rect 247 1030 251 1034
rect 255 1030 259 1034
rect 327 1030 331 1034
rect 399 1030 403 1034
rect 415 1030 419 1034
rect 463 1030 467 1034
rect 503 1030 507 1034
rect 519 1030 523 1034
rect 575 1030 579 1034
rect 583 1030 587 1034
rect 623 1030 627 1034
rect 663 1030 667 1034
rect 671 1030 675 1034
rect 735 1030 739 1034
rect 799 1030 803 1034
rect 807 1030 811 1034
rect 863 1030 867 1034
rect 895 1030 899 1034
rect 919 1030 923 1034
rect 983 1030 987 1034
rect 999 1030 1003 1034
rect 1047 1030 1051 1034
rect 1103 1030 1107 1034
rect 1191 1030 1195 1034
rect 1239 1030 1243 1034
rect 1279 1034 1283 1038
rect 1431 1034 1435 1038
rect 1471 1034 1475 1038
rect 1511 1034 1515 1038
rect 1559 1034 1563 1038
rect 1575 1034 1579 1038
rect 1615 1034 1619 1038
rect 1655 1034 1659 1038
rect 1671 1034 1675 1038
rect 1695 1034 1699 1038
rect 1727 1034 1731 1038
rect 1735 1034 1739 1038
rect 1775 1034 1779 1038
rect 1823 1034 1827 1038
rect 1871 1034 1875 1038
rect 1879 1034 1883 1038
rect 1919 1034 1923 1038
rect 1943 1034 1947 1038
rect 1967 1034 1971 1038
rect 2015 1034 2019 1038
rect 2063 1034 2067 1038
rect 2095 1034 2099 1038
rect 2119 1034 2123 1038
rect 2175 1034 2179 1038
rect 2231 1034 2235 1038
rect 2255 1034 2259 1038
rect 2407 1034 2411 1038
rect 111 962 115 966
rect 175 962 179 966
rect 215 962 219 966
rect 255 962 259 966
rect 303 962 307 966
rect 327 962 331 966
rect 359 962 363 966
rect 399 962 403 966
rect 415 962 419 966
rect 463 962 467 966
rect 519 962 523 966
rect 575 962 579 966
rect 623 962 627 966
rect 639 962 643 966
rect 671 962 675 966
rect 711 962 715 966
rect 735 962 739 966
rect 783 962 787 966
rect 807 962 811 966
rect 855 962 859 966
rect 895 962 899 966
rect 927 962 931 966
rect 999 962 1003 966
rect 1071 962 1075 966
rect 1103 962 1107 966
rect 1143 962 1147 966
rect 1191 962 1195 966
rect 1239 962 1243 966
rect 1279 958 1283 962
rect 1303 958 1307 962
rect 1351 958 1355 962
rect 1431 958 1435 962
rect 1511 958 1515 962
rect 1575 958 1579 962
rect 1591 958 1595 962
rect 1615 958 1619 962
rect 1655 958 1659 962
rect 1679 958 1683 962
rect 1695 958 1699 962
rect 1735 958 1739 962
rect 1767 958 1771 962
rect 1775 958 1779 962
rect 1823 958 1827 962
rect 1855 958 1859 962
rect 1879 958 1883 962
rect 1943 958 1947 962
rect 2015 958 2019 962
rect 2023 958 2027 962
rect 2095 958 2099 962
rect 2103 958 2107 962
rect 2175 958 2179 962
rect 2183 958 2187 962
rect 2255 958 2259 962
rect 2271 958 2275 962
rect 2407 958 2411 962
rect 111 886 115 890
rect 191 886 195 890
rect 215 886 219 890
rect 231 886 235 890
rect 255 886 259 890
rect 287 886 291 890
rect 303 886 307 890
rect 359 886 363 890
rect 415 886 419 890
rect 447 886 451 890
rect 463 886 467 890
rect 519 886 523 890
rect 543 886 547 890
rect 575 886 579 890
rect 639 886 643 890
rect 711 886 715 890
rect 727 886 731 890
rect 783 886 787 890
rect 807 886 811 890
rect 855 886 859 890
rect 887 886 891 890
rect 927 886 931 890
rect 959 886 963 890
rect 999 886 1003 890
rect 1023 886 1027 890
rect 1071 886 1075 890
rect 1087 886 1091 890
rect 1143 886 1147 890
rect 1159 886 1163 890
rect 1191 886 1195 890
rect 1239 886 1243 890
rect 1279 890 1283 894
rect 1303 890 1307 894
rect 1351 890 1355 894
rect 1431 890 1435 894
rect 1439 890 1443 894
rect 1479 890 1483 894
rect 1511 890 1515 894
rect 1519 890 1523 894
rect 1559 890 1563 894
rect 1591 890 1595 894
rect 1607 890 1611 894
rect 1655 890 1659 894
rect 1679 890 1683 894
rect 1711 890 1715 894
rect 1767 890 1771 894
rect 1775 890 1779 894
rect 1847 890 1851 894
rect 1855 890 1859 894
rect 1919 890 1923 894
rect 1943 890 1947 894
rect 1991 890 1995 894
rect 2023 890 2027 894
rect 2063 890 2067 894
rect 2103 890 2107 894
rect 2135 890 2139 894
rect 2183 890 2187 894
rect 2215 890 2219 894
rect 2271 890 2275 894
rect 2295 890 2299 894
rect 2407 890 2411 894
rect 111 818 115 822
rect 135 818 139 822
rect 175 818 179 822
rect 191 818 195 822
rect 231 818 235 822
rect 239 818 243 822
rect 287 818 291 822
rect 327 818 331 822
rect 359 818 363 822
rect 415 818 419 822
rect 447 818 451 822
rect 503 818 507 822
rect 543 818 547 822
rect 591 818 595 822
rect 639 818 643 822
rect 671 818 675 822
rect 727 818 731 822
rect 743 818 747 822
rect 807 818 811 822
rect 815 818 819 822
rect 879 818 883 822
rect 887 818 891 822
rect 943 818 947 822
rect 959 818 963 822
rect 1015 818 1019 822
rect 1023 818 1027 822
rect 1087 818 1091 822
rect 1159 818 1163 822
rect 1239 818 1243 822
rect 1279 810 1283 814
rect 1359 810 1363 814
rect 1415 810 1419 814
rect 1439 810 1443 814
rect 1471 810 1475 814
rect 1479 810 1483 814
rect 1519 810 1523 814
rect 1535 810 1539 814
rect 1559 810 1563 814
rect 1591 810 1595 814
rect 1607 810 1611 814
rect 1647 810 1651 814
rect 1655 810 1659 814
rect 1703 810 1707 814
rect 1711 810 1715 814
rect 1759 810 1763 814
rect 1775 810 1779 814
rect 1815 810 1819 814
rect 1847 810 1851 814
rect 1871 810 1875 814
rect 1919 810 1923 814
rect 1935 810 1939 814
rect 1991 810 1995 814
rect 1999 810 2003 814
rect 2063 810 2067 814
rect 2071 810 2075 814
rect 2135 810 2139 814
rect 2143 810 2147 814
rect 2215 810 2219 814
rect 2223 810 2227 814
rect 2295 810 2299 814
rect 2303 810 2307 814
rect 2359 810 2363 814
rect 2407 810 2411 814
rect 111 746 115 750
rect 135 746 139 750
rect 175 746 179 750
rect 191 746 195 750
rect 239 746 243 750
rect 263 746 267 750
rect 327 746 331 750
rect 335 746 339 750
rect 399 746 403 750
rect 415 746 419 750
rect 455 746 459 750
rect 503 746 507 750
rect 543 746 547 750
rect 583 746 587 750
rect 591 746 595 750
rect 623 746 627 750
rect 671 746 675 750
rect 719 746 723 750
rect 743 746 747 750
rect 767 746 771 750
rect 815 746 819 750
rect 863 746 867 750
rect 879 746 883 750
rect 911 746 915 750
rect 943 746 947 750
rect 1015 746 1019 750
rect 1239 746 1243 750
rect 1279 742 1283 746
rect 1303 742 1307 746
rect 1343 742 1347 746
rect 1359 742 1363 746
rect 1407 742 1411 746
rect 1415 742 1419 746
rect 1471 742 1475 746
rect 1487 742 1491 746
rect 1535 742 1539 746
rect 1575 742 1579 746
rect 1591 742 1595 746
rect 1647 742 1651 746
rect 1663 742 1667 746
rect 1703 742 1707 746
rect 1751 742 1755 746
rect 1759 742 1763 746
rect 1815 742 1819 746
rect 1831 742 1835 746
rect 1871 742 1875 746
rect 1911 742 1915 746
rect 1935 742 1939 746
rect 1991 742 1995 746
rect 1999 742 2003 746
rect 2071 742 2075 746
rect 2079 742 2083 746
rect 2143 742 2147 746
rect 2175 742 2179 746
rect 2223 742 2227 746
rect 2279 742 2283 746
rect 2303 742 2307 746
rect 2359 742 2363 746
rect 2407 742 2411 746
rect 111 674 115 678
rect 135 674 139 678
rect 191 674 195 678
rect 199 674 203 678
rect 263 674 267 678
rect 279 674 283 678
rect 335 674 339 678
rect 351 674 355 678
rect 399 674 403 678
rect 415 674 419 678
rect 455 674 459 678
rect 487 674 491 678
rect 503 674 507 678
rect 543 674 547 678
rect 559 674 563 678
rect 583 674 587 678
rect 623 674 627 678
rect 639 674 643 678
rect 671 674 675 678
rect 711 674 715 678
rect 719 674 723 678
rect 767 674 771 678
rect 783 674 787 678
rect 815 674 819 678
rect 855 674 859 678
rect 863 674 867 678
rect 911 674 915 678
rect 919 674 923 678
rect 983 674 987 678
rect 1039 674 1043 678
rect 1095 674 1099 678
rect 1151 674 1155 678
rect 1191 674 1195 678
rect 1239 674 1243 678
rect 1279 670 1283 674
rect 1303 670 1307 674
rect 1343 670 1347 674
rect 1399 670 1403 674
rect 1407 670 1411 674
rect 1487 670 1491 674
rect 1511 670 1515 674
rect 1575 670 1579 674
rect 1623 670 1627 674
rect 1663 670 1667 674
rect 1727 670 1731 674
rect 1751 670 1755 674
rect 1815 670 1819 674
rect 1831 670 1835 674
rect 1895 670 1899 674
rect 1911 670 1915 674
rect 1975 670 1979 674
rect 1991 670 1995 674
rect 2047 670 2051 674
rect 2079 670 2083 674
rect 2111 670 2115 674
rect 2175 670 2179 674
rect 2239 670 2243 674
rect 2279 670 2283 674
rect 2311 670 2315 674
rect 2359 670 2363 674
rect 2407 670 2411 674
rect 111 598 115 602
rect 135 598 139 602
rect 191 598 195 602
rect 199 598 203 602
rect 271 598 275 602
rect 279 598 283 602
rect 351 598 355 602
rect 359 598 363 602
rect 415 598 419 602
rect 447 598 451 602
rect 487 598 491 602
rect 535 598 539 602
rect 559 598 563 602
rect 623 598 627 602
rect 639 598 643 602
rect 703 598 707 602
rect 711 598 715 602
rect 783 598 787 602
rect 855 598 859 602
rect 919 598 923 602
rect 975 598 979 602
rect 983 598 987 602
rect 1023 598 1027 602
rect 1039 598 1043 602
rect 1079 598 1083 602
rect 1095 598 1099 602
rect 1135 598 1139 602
rect 1151 598 1155 602
rect 1191 598 1195 602
rect 1239 598 1243 602
rect 1279 598 1283 602
rect 1303 598 1307 602
rect 1399 598 1403 602
rect 1415 598 1419 602
rect 1455 598 1459 602
rect 1495 598 1499 602
rect 1511 598 1515 602
rect 1543 598 1547 602
rect 1599 598 1603 602
rect 1623 598 1627 602
rect 1663 598 1667 602
rect 1727 598 1731 602
rect 1791 598 1795 602
rect 1815 598 1819 602
rect 1847 598 1851 602
rect 1895 598 1899 602
rect 1911 598 1915 602
rect 1975 598 1979 602
rect 2047 598 2051 602
rect 2111 598 2115 602
rect 2119 598 2123 602
rect 2175 598 2179 602
rect 2199 598 2203 602
rect 2239 598 2243 602
rect 2287 598 2291 602
rect 2311 598 2315 602
rect 2359 598 2363 602
rect 2407 598 2411 602
rect 1279 530 1283 534
rect 1303 530 1307 534
rect 1375 530 1379 534
rect 1415 530 1419 534
rect 1455 530 1459 534
rect 1479 530 1483 534
rect 1495 530 1499 534
rect 1543 530 1547 534
rect 1583 530 1587 534
rect 1599 530 1603 534
rect 1663 530 1667 534
rect 1695 530 1699 534
rect 1727 530 1731 534
rect 1791 530 1795 534
rect 1799 530 1803 534
rect 1847 530 1851 534
rect 1903 530 1907 534
rect 1911 530 1915 534
rect 1975 530 1979 534
rect 2007 530 2011 534
rect 2047 530 2051 534
rect 2103 530 2107 534
rect 2119 530 2123 534
rect 2191 530 2195 534
rect 2199 530 2203 534
rect 2287 530 2291 534
rect 2359 530 2363 534
rect 2407 530 2411 534
rect 111 522 115 526
rect 135 522 139 526
rect 191 522 195 526
rect 263 522 267 526
rect 271 522 275 526
rect 335 522 339 526
rect 359 522 363 526
rect 415 522 419 526
rect 447 522 451 526
rect 495 522 499 526
rect 535 522 539 526
rect 575 522 579 526
rect 623 522 627 526
rect 647 522 651 526
rect 703 522 707 526
rect 719 522 723 526
rect 783 522 787 526
rect 847 522 851 526
rect 855 522 859 526
rect 903 522 907 526
rect 919 522 923 526
rect 959 522 963 526
rect 975 522 979 526
rect 1023 522 1027 526
rect 1079 522 1083 526
rect 1087 522 1091 526
rect 1135 522 1139 526
rect 1151 522 1155 526
rect 1191 522 1195 526
rect 1239 522 1243 526
rect 111 454 115 458
rect 135 454 139 458
rect 183 454 187 458
rect 191 454 195 458
rect 223 454 227 458
rect 263 454 267 458
rect 311 454 315 458
rect 335 454 339 458
rect 367 454 371 458
rect 415 454 419 458
rect 431 454 435 458
rect 495 454 499 458
rect 559 454 563 458
rect 575 454 579 458
rect 615 454 619 458
rect 647 454 651 458
rect 671 454 675 458
rect 719 454 723 458
rect 775 454 779 458
rect 783 454 787 458
rect 831 454 835 458
rect 847 454 851 458
rect 887 454 891 458
rect 903 454 907 458
rect 959 454 963 458
rect 1023 454 1027 458
rect 1087 454 1091 458
rect 1151 454 1155 458
rect 1191 454 1195 458
rect 1239 454 1243 458
rect 1279 458 1283 462
rect 1303 458 1307 462
rect 1343 458 1347 462
rect 1375 458 1379 462
rect 1399 458 1403 462
rect 1463 458 1467 462
rect 1479 458 1483 462
rect 1527 458 1531 462
rect 1583 458 1587 462
rect 1591 458 1595 462
rect 1663 458 1667 462
rect 1695 458 1699 462
rect 1735 458 1739 462
rect 1799 458 1803 462
rect 1815 458 1819 462
rect 1895 458 1899 462
rect 1903 458 1907 462
rect 1975 458 1979 462
rect 2007 458 2011 462
rect 2055 458 2059 462
rect 2103 458 2107 462
rect 2135 458 2139 462
rect 2191 458 2195 462
rect 2215 458 2219 462
rect 2287 458 2291 462
rect 2295 458 2299 462
rect 2359 458 2363 462
rect 2407 458 2411 462
rect 111 386 115 390
rect 135 386 139 390
rect 175 386 179 390
rect 183 386 187 390
rect 223 386 227 390
rect 231 386 235 390
rect 263 386 267 390
rect 287 386 291 390
rect 311 386 315 390
rect 343 386 347 390
rect 367 386 371 390
rect 391 386 395 390
rect 431 386 435 390
rect 439 386 443 390
rect 487 386 491 390
rect 495 386 499 390
rect 535 386 539 390
rect 559 386 563 390
rect 583 386 587 390
rect 615 386 619 390
rect 631 386 635 390
rect 671 386 675 390
rect 679 386 683 390
rect 719 386 723 390
rect 727 386 731 390
rect 775 386 779 390
rect 831 386 835 390
rect 887 386 891 390
rect 1239 386 1243 390
rect 1279 386 1283 390
rect 1303 386 1307 390
rect 1343 386 1347 390
rect 1399 386 1403 390
rect 1447 386 1451 390
rect 1463 386 1467 390
rect 1487 386 1491 390
rect 1527 386 1531 390
rect 1535 386 1539 390
rect 1591 386 1595 390
rect 1663 386 1667 390
rect 1735 386 1739 390
rect 1815 386 1819 390
rect 1895 386 1899 390
rect 1967 386 1971 390
rect 1975 386 1979 390
rect 2039 386 2043 390
rect 2055 386 2059 390
rect 2111 386 2115 390
rect 2135 386 2139 390
rect 2175 386 2179 390
rect 2215 386 2219 390
rect 2239 386 2243 390
rect 2295 386 2299 390
rect 2303 386 2307 390
rect 2359 386 2363 390
rect 2407 386 2411 390
rect 111 314 115 318
rect 135 314 139 318
rect 175 314 179 318
rect 183 314 187 318
rect 231 314 235 318
rect 255 314 259 318
rect 287 314 291 318
rect 327 314 331 318
rect 343 314 347 318
rect 391 314 395 318
rect 439 314 443 318
rect 447 314 451 318
rect 487 314 491 318
rect 503 314 507 318
rect 535 314 539 318
rect 551 314 555 318
rect 583 314 587 318
rect 591 314 595 318
rect 631 314 635 318
rect 679 314 683 318
rect 727 314 731 318
rect 775 314 779 318
rect 823 314 827 318
rect 871 314 875 318
rect 919 314 923 318
rect 1239 314 1243 318
rect 1279 314 1283 318
rect 1447 314 1451 318
rect 1487 314 1491 318
rect 1495 314 1499 318
rect 1535 314 1539 318
rect 1575 314 1579 318
rect 1591 314 1595 318
rect 1615 314 1619 318
rect 1655 314 1659 318
rect 1663 314 1667 318
rect 1695 314 1699 318
rect 1735 314 1739 318
rect 1743 314 1747 318
rect 1799 314 1803 318
rect 1815 314 1819 318
rect 1863 314 1867 318
rect 1895 314 1899 318
rect 1935 314 1939 318
rect 1967 314 1971 318
rect 2007 314 2011 318
rect 2039 314 2043 318
rect 2071 314 2075 318
rect 2111 314 2115 318
rect 2135 314 2139 318
rect 2175 314 2179 318
rect 2191 314 2195 318
rect 2239 314 2243 318
rect 2255 314 2259 318
rect 2303 314 2307 318
rect 2319 314 2323 318
rect 2359 314 2363 318
rect 2407 314 2411 318
rect 111 238 115 242
rect 135 238 139 242
rect 175 238 179 242
rect 183 238 187 242
rect 247 238 251 242
rect 255 238 259 242
rect 327 238 331 242
rect 391 238 395 242
rect 415 238 419 242
rect 447 238 451 242
rect 495 238 499 242
rect 503 238 507 242
rect 551 238 555 242
rect 575 238 579 242
rect 591 238 595 242
rect 631 238 635 242
rect 655 238 659 242
rect 679 238 683 242
rect 727 238 731 242
rect 775 238 779 242
rect 791 238 795 242
rect 823 238 827 242
rect 847 238 851 242
rect 871 238 875 242
rect 903 238 907 242
rect 919 238 923 242
rect 959 238 963 242
rect 1023 238 1027 242
rect 1239 238 1243 242
rect 1279 242 1283 246
rect 1367 242 1371 246
rect 1407 242 1411 246
rect 1447 242 1451 246
rect 1495 242 1499 246
rect 1535 242 1539 246
rect 1551 242 1555 246
rect 1575 242 1579 246
rect 1607 242 1611 246
rect 1615 242 1619 246
rect 1655 242 1659 246
rect 1671 242 1675 246
rect 1695 242 1699 246
rect 1735 242 1739 246
rect 1743 242 1747 246
rect 1799 242 1803 246
rect 1807 242 1811 246
rect 1863 242 1867 246
rect 1887 242 1891 246
rect 1935 242 1939 246
rect 1975 242 1979 246
rect 2007 242 2011 246
rect 2071 242 2075 246
rect 2135 242 2139 246
rect 2167 242 2171 246
rect 2191 242 2195 246
rect 2255 242 2259 246
rect 2271 242 2275 246
rect 2319 242 2323 246
rect 2359 242 2363 246
rect 2407 242 2411 246
rect 1279 158 1283 162
rect 1303 158 1307 162
rect 1343 158 1347 162
rect 1367 158 1371 162
rect 1383 158 1387 162
rect 1407 158 1411 162
rect 1423 158 1427 162
rect 1447 158 1451 162
rect 1463 158 1467 162
rect 1495 158 1499 162
rect 1519 158 1523 162
rect 1551 158 1555 162
rect 1583 158 1587 162
rect 1607 158 1611 162
rect 1647 158 1651 162
rect 1671 158 1675 162
rect 1711 158 1715 162
rect 1735 158 1739 162
rect 1767 158 1771 162
rect 1807 158 1811 162
rect 1823 158 1827 162
rect 1871 158 1875 162
rect 1887 158 1891 162
rect 1919 158 1923 162
rect 1967 158 1971 162
rect 1975 158 1979 162
rect 2015 158 2019 162
rect 2063 158 2067 162
rect 2071 158 2075 162
rect 2111 158 2115 162
rect 2159 158 2163 162
rect 2167 158 2171 162
rect 2215 158 2219 162
rect 2271 158 2275 162
rect 2319 158 2323 162
rect 2359 158 2363 162
rect 2407 158 2411 162
rect 111 150 115 154
rect 135 150 139 154
rect 175 150 179 154
rect 215 150 219 154
rect 247 150 251 154
rect 255 150 259 154
rect 295 150 299 154
rect 327 150 331 154
rect 335 150 339 154
rect 375 150 379 154
rect 415 150 419 154
rect 423 150 427 154
rect 471 150 475 154
rect 495 150 499 154
rect 527 150 531 154
rect 575 150 579 154
rect 583 150 587 154
rect 631 150 635 154
rect 655 150 659 154
rect 679 150 683 154
rect 727 150 731 154
rect 767 150 771 154
rect 791 150 795 154
rect 807 150 811 154
rect 847 150 851 154
rect 887 150 891 154
rect 903 150 907 154
rect 927 150 931 154
rect 959 150 963 154
rect 975 150 979 154
rect 1023 150 1027 154
rect 1071 150 1075 154
rect 1111 150 1115 154
rect 1151 150 1155 154
rect 1191 150 1195 154
rect 1239 150 1243 154
rect 1279 90 1283 94
rect 1303 90 1307 94
rect 1343 90 1347 94
rect 1383 90 1387 94
rect 1423 90 1427 94
rect 1463 90 1467 94
rect 1519 90 1523 94
rect 1583 90 1587 94
rect 1647 90 1651 94
rect 1711 90 1715 94
rect 1767 90 1771 94
rect 1823 90 1827 94
rect 1871 90 1875 94
rect 1919 90 1923 94
rect 1967 90 1971 94
rect 2015 90 2019 94
rect 2063 90 2067 94
rect 2111 90 2115 94
rect 2159 90 2163 94
rect 2215 90 2219 94
rect 2271 90 2275 94
rect 2319 90 2323 94
rect 2359 90 2363 94
rect 2407 90 2411 94
rect 111 82 115 86
rect 135 82 139 86
rect 175 82 179 86
rect 215 82 219 86
rect 255 82 259 86
rect 295 82 299 86
rect 335 82 339 86
rect 375 82 379 86
rect 423 82 427 86
rect 471 82 475 86
rect 527 82 531 86
rect 583 82 587 86
rect 631 82 635 86
rect 679 82 683 86
rect 727 82 731 86
rect 767 82 771 86
rect 807 82 811 86
rect 847 82 851 86
rect 887 82 891 86
rect 927 82 931 86
rect 975 82 979 86
rect 1023 82 1027 86
rect 1071 82 1075 86
rect 1111 82 1115 86
rect 1151 82 1155 86
rect 1191 82 1195 86
rect 1239 82 1243 86
<< m4 >>
rect 1250 2509 1251 2515
rect 1257 2514 2435 2515
rect 1257 2510 1279 2514
rect 1283 2510 1535 2514
rect 1539 2510 1575 2514
rect 1579 2510 1615 2514
rect 1619 2510 1655 2514
rect 1659 2510 1695 2514
rect 1699 2510 1735 2514
rect 1739 2510 1775 2514
rect 1779 2510 1815 2514
rect 1819 2510 1855 2514
rect 1859 2510 1895 2514
rect 1899 2510 1935 2514
rect 1939 2510 1975 2514
rect 1979 2510 2407 2514
rect 2411 2510 2435 2514
rect 1257 2509 2435 2510
rect 2441 2509 2442 2515
rect 96 2497 97 2503
rect 103 2502 1263 2503
rect 103 2498 111 2502
rect 115 2498 135 2502
rect 139 2498 175 2502
rect 179 2498 215 2502
rect 219 2498 255 2502
rect 259 2498 311 2502
rect 315 2498 391 2502
rect 395 2498 479 2502
rect 483 2498 567 2502
rect 571 2498 655 2502
rect 659 2498 743 2502
rect 747 2498 831 2502
rect 835 2498 927 2502
rect 931 2498 1239 2502
rect 1243 2498 1263 2502
rect 103 2497 1263 2498
rect 1269 2497 1270 2503
rect 1262 2441 1263 2447
rect 1269 2446 2447 2447
rect 1269 2442 1279 2446
rect 1283 2442 1359 2446
rect 1363 2442 1399 2446
rect 1403 2442 1455 2446
rect 1459 2442 1519 2446
rect 1523 2442 1535 2446
rect 1539 2442 1575 2446
rect 1579 2442 1599 2446
rect 1603 2442 1615 2446
rect 1619 2442 1655 2446
rect 1659 2442 1679 2446
rect 1683 2442 1695 2446
rect 1699 2442 1735 2446
rect 1739 2442 1759 2446
rect 1763 2442 1775 2446
rect 1779 2442 1815 2446
rect 1819 2442 1839 2446
rect 1843 2442 1855 2446
rect 1859 2442 1895 2446
rect 1899 2442 1919 2446
rect 1923 2442 1935 2446
rect 1939 2442 1975 2446
rect 1979 2442 1999 2446
rect 2003 2442 2079 2446
rect 2083 2442 2159 2446
rect 2163 2442 2247 2446
rect 2251 2442 2335 2446
rect 2339 2442 2407 2446
rect 2411 2442 2447 2446
rect 1269 2441 2447 2442
rect 2453 2441 2454 2447
rect 84 2429 85 2435
rect 91 2434 1251 2435
rect 91 2430 111 2434
rect 115 2430 135 2434
rect 139 2430 175 2434
rect 179 2430 183 2434
rect 187 2430 215 2434
rect 219 2430 247 2434
rect 251 2430 255 2434
rect 259 2430 311 2434
rect 315 2430 319 2434
rect 323 2430 391 2434
rect 395 2430 471 2434
rect 475 2430 479 2434
rect 483 2430 543 2434
rect 547 2430 567 2434
rect 571 2430 615 2434
rect 619 2430 655 2434
rect 659 2430 679 2434
rect 683 2430 735 2434
rect 739 2430 743 2434
rect 747 2430 791 2434
rect 795 2430 831 2434
rect 835 2430 839 2434
rect 843 2430 887 2434
rect 891 2430 927 2434
rect 931 2430 935 2434
rect 939 2430 991 2434
rect 995 2430 1047 2434
rect 1051 2430 1239 2434
rect 1243 2430 1251 2434
rect 91 2429 1251 2430
rect 1257 2429 1258 2435
rect 1250 2373 1251 2379
rect 1257 2378 2435 2379
rect 1257 2374 1279 2378
rect 1283 2374 1359 2378
rect 1363 2374 1399 2378
rect 1403 2374 1407 2378
rect 1411 2374 1455 2378
rect 1459 2374 1471 2378
rect 1475 2374 1519 2378
rect 1523 2374 1543 2378
rect 1547 2374 1599 2378
rect 1603 2374 1615 2378
rect 1619 2374 1679 2378
rect 1683 2374 1695 2378
rect 1699 2374 1759 2378
rect 1763 2374 1775 2378
rect 1779 2374 1839 2378
rect 1843 2374 1855 2378
rect 1859 2374 1919 2378
rect 1923 2374 1927 2378
rect 1931 2374 1999 2378
rect 2003 2374 2071 2378
rect 2075 2374 2079 2378
rect 2083 2374 2143 2378
rect 2147 2374 2159 2378
rect 2163 2374 2223 2378
rect 2227 2374 2247 2378
rect 2251 2374 2303 2378
rect 2307 2374 2335 2378
rect 2339 2374 2359 2378
rect 2363 2374 2407 2378
rect 2411 2374 2435 2378
rect 1257 2373 2435 2374
rect 2441 2373 2442 2379
rect 96 2353 97 2359
rect 103 2358 1263 2359
rect 103 2354 111 2358
rect 115 2354 135 2358
rect 139 2354 175 2358
rect 179 2354 183 2358
rect 187 2354 215 2358
rect 219 2354 247 2358
rect 251 2354 271 2358
rect 275 2354 319 2358
rect 323 2354 351 2358
rect 355 2354 391 2358
rect 395 2354 431 2358
rect 435 2354 471 2358
rect 475 2354 519 2358
rect 523 2354 543 2358
rect 547 2354 599 2358
rect 603 2354 615 2358
rect 619 2354 679 2358
rect 683 2354 735 2358
rect 739 2354 751 2358
rect 755 2354 791 2358
rect 795 2354 823 2358
rect 827 2354 839 2358
rect 843 2354 887 2358
rect 891 2354 935 2358
rect 939 2354 959 2358
rect 963 2354 991 2358
rect 995 2354 1031 2358
rect 1035 2354 1047 2358
rect 1051 2354 1239 2358
rect 1243 2354 1263 2358
rect 103 2353 1263 2354
rect 1269 2353 1270 2359
rect 1262 2301 1263 2307
rect 1269 2306 2447 2307
rect 1269 2302 1279 2306
rect 1283 2302 1359 2306
rect 1363 2302 1407 2306
rect 1411 2302 1471 2306
rect 1475 2302 1503 2306
rect 1507 2302 1543 2306
rect 1547 2302 1583 2306
rect 1587 2302 1615 2306
rect 1619 2302 1623 2306
rect 1627 2302 1663 2306
rect 1667 2302 1695 2306
rect 1699 2302 1703 2306
rect 1707 2302 1759 2306
rect 1763 2302 1775 2306
rect 1779 2302 1823 2306
rect 1827 2302 1855 2306
rect 1859 2302 1895 2306
rect 1899 2302 1927 2306
rect 1931 2302 1967 2306
rect 1971 2302 1999 2306
rect 2003 2302 2047 2306
rect 2051 2302 2071 2306
rect 2075 2302 2127 2306
rect 2131 2302 2143 2306
rect 2147 2302 2207 2306
rect 2211 2302 2223 2306
rect 2227 2302 2295 2306
rect 2299 2302 2303 2306
rect 2307 2302 2359 2306
rect 2363 2302 2407 2306
rect 2411 2302 2447 2306
rect 1269 2301 2447 2302
rect 2453 2301 2454 2307
rect 84 2281 85 2287
rect 91 2286 1251 2287
rect 91 2282 111 2286
rect 115 2282 135 2286
rect 139 2282 175 2286
rect 179 2282 215 2286
rect 219 2282 231 2286
rect 235 2282 271 2286
rect 275 2282 303 2286
rect 307 2282 351 2286
rect 355 2282 375 2286
rect 379 2282 431 2286
rect 435 2282 455 2286
rect 459 2282 519 2286
rect 523 2282 535 2286
rect 539 2282 599 2286
rect 603 2282 615 2286
rect 619 2282 679 2286
rect 683 2282 687 2286
rect 691 2282 751 2286
rect 755 2282 759 2286
rect 763 2282 823 2286
rect 827 2282 831 2286
rect 835 2282 887 2286
rect 891 2282 911 2286
rect 915 2282 959 2286
rect 963 2282 991 2286
rect 995 2282 1031 2286
rect 1035 2282 1239 2286
rect 1243 2282 1251 2286
rect 91 2281 1251 2282
rect 1257 2281 1258 2287
rect 1250 2225 1251 2231
rect 1257 2230 2435 2231
rect 1257 2226 1279 2230
rect 1283 2226 1303 2230
rect 1307 2226 1343 2230
rect 1347 2226 1383 2230
rect 1387 2226 1431 2230
rect 1435 2226 1495 2230
rect 1499 2226 1503 2230
rect 1507 2226 1543 2230
rect 1547 2226 1567 2230
rect 1571 2226 1583 2230
rect 1587 2226 1623 2230
rect 1627 2226 1639 2230
rect 1643 2226 1663 2230
rect 1667 2226 1703 2230
rect 1707 2226 1711 2230
rect 1715 2226 1759 2230
rect 1763 2226 1783 2230
rect 1787 2226 1823 2230
rect 1827 2226 1855 2230
rect 1859 2226 1895 2230
rect 1899 2226 1935 2230
rect 1939 2226 1967 2230
rect 1971 2226 2015 2230
rect 2019 2226 2047 2230
rect 2051 2226 2095 2230
rect 2099 2226 2127 2230
rect 2131 2226 2183 2230
rect 2187 2226 2207 2230
rect 2211 2226 2279 2230
rect 2283 2226 2295 2230
rect 2299 2226 2359 2230
rect 2363 2226 2407 2230
rect 2411 2226 2435 2230
rect 1257 2225 2435 2226
rect 2441 2225 2442 2231
rect 96 2213 97 2219
rect 103 2218 1263 2219
rect 103 2214 111 2218
rect 115 2214 135 2218
rect 139 2214 175 2218
rect 179 2214 231 2218
rect 235 2214 247 2218
rect 251 2214 287 2218
rect 291 2214 303 2218
rect 307 2214 327 2218
rect 331 2214 375 2218
rect 379 2214 431 2218
rect 435 2214 455 2218
rect 459 2214 495 2218
rect 499 2214 535 2218
rect 539 2214 551 2218
rect 555 2214 607 2218
rect 611 2214 615 2218
rect 619 2214 663 2218
rect 667 2214 687 2218
rect 691 2214 719 2218
rect 723 2214 759 2218
rect 763 2214 783 2218
rect 787 2214 831 2218
rect 835 2214 847 2218
rect 851 2214 911 2218
rect 915 2214 991 2218
rect 995 2214 1239 2218
rect 1243 2214 1263 2218
rect 103 2213 1263 2214
rect 1269 2213 1270 2219
rect 1262 2157 1263 2163
rect 1269 2162 2447 2163
rect 1269 2158 1279 2162
rect 1283 2158 1303 2162
rect 1307 2158 1343 2162
rect 1347 2158 1351 2162
rect 1355 2158 1383 2162
rect 1387 2158 1431 2162
rect 1435 2158 1439 2162
rect 1443 2158 1495 2162
rect 1499 2158 1535 2162
rect 1539 2158 1567 2162
rect 1571 2158 1631 2162
rect 1635 2158 1639 2162
rect 1643 2158 1711 2162
rect 1715 2158 1727 2162
rect 1731 2158 1783 2162
rect 1787 2158 1815 2162
rect 1819 2158 1855 2162
rect 1859 2158 1895 2162
rect 1899 2158 1935 2162
rect 1939 2158 1975 2162
rect 1979 2158 2015 2162
rect 2019 2158 2047 2162
rect 2051 2158 2095 2162
rect 2099 2158 2111 2162
rect 2115 2158 2175 2162
rect 2179 2158 2183 2162
rect 2187 2158 2239 2162
rect 2243 2158 2279 2162
rect 2283 2158 2311 2162
rect 2315 2158 2359 2162
rect 2363 2158 2407 2162
rect 2411 2158 2447 2162
rect 1269 2157 2447 2158
rect 2453 2157 2454 2163
rect 84 2137 85 2143
rect 91 2142 1251 2143
rect 91 2138 111 2142
rect 115 2138 247 2142
rect 251 2138 287 2142
rect 291 2138 327 2142
rect 331 2138 375 2142
rect 379 2138 383 2142
rect 387 2138 423 2142
rect 427 2138 431 2142
rect 435 2138 463 2142
rect 467 2138 495 2142
rect 499 2138 503 2142
rect 507 2138 551 2142
rect 555 2138 607 2142
rect 611 2138 663 2142
rect 667 2138 719 2142
rect 723 2138 727 2142
rect 731 2138 783 2142
rect 787 2138 791 2142
rect 795 2138 847 2142
rect 851 2138 855 2142
rect 859 2138 911 2142
rect 915 2138 967 2142
rect 971 2138 1023 2142
rect 1027 2138 1079 2142
rect 1083 2138 1143 2142
rect 1147 2138 1239 2142
rect 1243 2138 1251 2142
rect 91 2137 1251 2138
rect 1257 2137 1258 2143
rect 1250 2085 1251 2091
rect 1257 2090 2435 2091
rect 1257 2086 1279 2090
rect 1283 2086 1303 2090
rect 1307 2086 1343 2090
rect 1347 2086 1351 2090
rect 1355 2086 1399 2090
rect 1403 2086 1439 2090
rect 1443 2086 1479 2090
rect 1483 2086 1535 2090
rect 1539 2086 1567 2090
rect 1571 2086 1631 2090
rect 1635 2086 1663 2090
rect 1667 2086 1727 2090
rect 1731 2086 1759 2090
rect 1763 2086 1815 2090
rect 1819 2086 1847 2090
rect 1851 2086 1895 2090
rect 1899 2086 1935 2090
rect 1939 2086 1975 2090
rect 1979 2086 2015 2090
rect 2019 2086 2047 2090
rect 2051 2086 2095 2090
rect 2099 2086 2111 2090
rect 2115 2086 2167 2090
rect 2171 2086 2175 2090
rect 2179 2086 2239 2090
rect 2243 2086 2311 2090
rect 2315 2086 2359 2090
rect 2363 2086 2407 2090
rect 2411 2086 2435 2090
rect 1257 2085 2435 2086
rect 2441 2085 2442 2091
rect 96 2069 97 2075
rect 103 2074 1263 2075
rect 103 2070 111 2074
rect 115 2070 383 2074
rect 387 2070 423 2074
rect 427 2070 463 2074
rect 467 2070 503 2074
rect 507 2070 543 2074
rect 547 2070 551 2074
rect 555 2070 583 2074
rect 587 2070 607 2074
rect 611 2070 631 2074
rect 635 2070 663 2074
rect 667 2070 687 2074
rect 691 2070 727 2074
rect 731 2070 743 2074
rect 747 2070 791 2074
rect 795 2070 799 2074
rect 803 2070 847 2074
rect 851 2070 855 2074
rect 859 2070 903 2074
rect 907 2070 911 2074
rect 915 2070 959 2074
rect 963 2070 967 2074
rect 971 2070 1015 2074
rect 1019 2070 1023 2074
rect 1027 2070 1071 2074
rect 1075 2070 1079 2074
rect 1083 2070 1143 2074
rect 1147 2070 1239 2074
rect 1243 2070 1263 2074
rect 103 2069 1263 2070
rect 1269 2069 1270 2075
rect 1262 2009 1263 2015
rect 1269 2014 2447 2015
rect 1269 2010 1279 2014
rect 1283 2010 1303 2014
rect 1307 2010 1343 2014
rect 1347 2010 1351 2014
rect 1355 2010 1399 2014
rect 1403 2010 1423 2014
rect 1427 2010 1479 2014
rect 1483 2010 1495 2014
rect 1499 2010 1567 2014
rect 1571 2010 1575 2014
rect 1579 2010 1663 2014
rect 1667 2010 1751 2014
rect 1755 2010 1759 2014
rect 1763 2010 1839 2014
rect 1843 2010 1847 2014
rect 1851 2010 1919 2014
rect 1923 2010 1935 2014
rect 1939 2010 1999 2014
rect 2003 2010 2015 2014
rect 2019 2010 2071 2014
rect 2075 2010 2095 2014
rect 2099 2010 2135 2014
rect 2139 2010 2167 2014
rect 2171 2010 2191 2014
rect 2195 2010 2239 2014
rect 2243 2010 2255 2014
rect 2259 2010 2311 2014
rect 2315 2010 2319 2014
rect 2323 2010 2359 2014
rect 2363 2010 2407 2014
rect 2411 2010 2447 2014
rect 1269 2009 2447 2010
rect 2453 2009 2454 2015
rect 84 1993 85 1999
rect 91 1998 1251 1999
rect 91 1994 111 1998
rect 115 1994 367 1998
rect 371 1994 383 1998
rect 387 1994 407 1998
rect 411 1994 423 1998
rect 427 1994 455 1998
rect 459 1994 463 1998
rect 467 1994 503 1998
rect 507 1994 511 1998
rect 515 1994 543 1998
rect 547 1994 567 1998
rect 571 1994 583 1998
rect 587 1994 631 1998
rect 635 1994 687 1998
rect 691 1994 695 1998
rect 699 1994 743 1998
rect 747 1994 759 1998
rect 763 1994 799 1998
rect 803 1994 815 1998
rect 819 1994 847 1998
rect 851 1994 871 1998
rect 875 1994 903 1998
rect 907 1994 935 1998
rect 939 1994 959 1998
rect 963 1994 999 1998
rect 1003 1994 1015 1998
rect 1019 1994 1063 1998
rect 1067 1994 1071 1998
rect 1075 1994 1239 1998
rect 1243 1994 1251 1998
rect 91 1993 1251 1994
rect 1257 1993 1258 1999
rect 1250 1941 1251 1947
rect 1257 1946 2435 1947
rect 1257 1942 1279 1946
rect 1283 1942 1303 1946
rect 1307 1942 1351 1946
rect 1355 1942 1359 1946
rect 1363 1942 1423 1946
rect 1427 1942 1447 1946
rect 1451 1942 1495 1946
rect 1499 1942 1535 1946
rect 1539 1942 1575 1946
rect 1579 1942 1623 1946
rect 1627 1942 1663 1946
rect 1667 1942 1711 1946
rect 1715 1942 1751 1946
rect 1755 1942 1791 1946
rect 1795 1942 1839 1946
rect 1843 1942 1863 1946
rect 1867 1942 1919 1946
rect 1923 1942 1935 1946
rect 1939 1942 1999 1946
rect 2003 1942 2007 1946
rect 2011 1942 2071 1946
rect 2075 1942 2079 1946
rect 2083 1942 2135 1946
rect 2139 1942 2151 1946
rect 2155 1942 2191 1946
rect 2195 1942 2223 1946
rect 2227 1942 2255 1946
rect 2259 1942 2303 1946
rect 2307 1942 2319 1946
rect 2323 1942 2359 1946
rect 2363 1942 2407 1946
rect 2411 1942 2435 1946
rect 1257 1941 2435 1942
rect 2441 1941 2442 1947
rect 96 1921 97 1927
rect 103 1926 1263 1927
rect 103 1922 111 1926
rect 115 1922 175 1926
rect 179 1922 215 1926
rect 219 1922 263 1926
rect 267 1922 319 1926
rect 323 1922 367 1926
rect 371 1922 391 1926
rect 395 1922 407 1926
rect 411 1922 455 1926
rect 459 1922 471 1926
rect 475 1922 511 1926
rect 515 1922 551 1926
rect 555 1922 567 1926
rect 571 1922 631 1926
rect 635 1922 639 1926
rect 643 1922 695 1926
rect 699 1922 719 1926
rect 723 1922 759 1926
rect 763 1922 799 1926
rect 803 1922 815 1926
rect 819 1922 871 1926
rect 875 1922 879 1926
rect 883 1922 935 1926
rect 939 1922 959 1926
rect 963 1922 999 1926
rect 1003 1922 1039 1926
rect 1043 1922 1063 1926
rect 1067 1922 1119 1926
rect 1123 1922 1239 1926
rect 1243 1922 1263 1926
rect 103 1921 1263 1922
rect 1269 1921 1270 1927
rect 1262 1873 1263 1879
rect 1269 1878 2447 1879
rect 1269 1874 1279 1878
rect 1283 1874 1303 1878
rect 1307 1874 1311 1878
rect 1315 1874 1359 1878
rect 1363 1874 1415 1878
rect 1419 1874 1447 1878
rect 1451 1874 1479 1878
rect 1483 1874 1535 1878
rect 1539 1874 1543 1878
rect 1547 1874 1615 1878
rect 1619 1874 1623 1878
rect 1627 1874 1687 1878
rect 1691 1874 1711 1878
rect 1715 1874 1767 1878
rect 1771 1874 1791 1878
rect 1795 1874 1863 1878
rect 1867 1874 1935 1878
rect 1939 1874 1975 1878
rect 1979 1874 2007 1878
rect 2011 1874 2079 1878
rect 2083 1874 2095 1878
rect 2099 1874 2151 1878
rect 2155 1874 2223 1878
rect 2227 1874 2303 1878
rect 2307 1874 2359 1878
rect 2363 1874 2407 1878
rect 2411 1874 2447 1878
rect 1269 1873 2447 1874
rect 2453 1873 2454 1879
rect 84 1845 85 1851
rect 91 1850 1251 1851
rect 91 1846 111 1850
rect 115 1846 135 1850
rect 139 1846 175 1850
rect 179 1846 215 1850
rect 219 1846 263 1850
rect 267 1846 271 1850
rect 275 1846 319 1850
rect 323 1846 351 1850
rect 355 1846 391 1850
rect 395 1846 439 1850
rect 443 1846 471 1850
rect 475 1846 535 1850
rect 539 1846 551 1850
rect 555 1846 631 1850
rect 635 1846 639 1850
rect 643 1846 719 1850
rect 723 1846 727 1850
rect 731 1846 799 1850
rect 803 1846 823 1850
rect 827 1846 879 1850
rect 883 1846 911 1850
rect 915 1846 959 1850
rect 963 1846 991 1850
rect 995 1846 1039 1850
rect 1043 1846 1063 1850
rect 1067 1846 1119 1850
rect 1123 1846 1135 1850
rect 1139 1846 1191 1850
rect 1195 1846 1239 1850
rect 1243 1846 1251 1850
rect 91 1845 1251 1846
rect 1257 1845 1258 1851
rect 1250 1801 1251 1807
rect 1257 1806 2435 1807
rect 1257 1802 1279 1806
rect 1283 1802 1311 1806
rect 1315 1802 1359 1806
rect 1363 1802 1407 1806
rect 1411 1802 1415 1806
rect 1419 1802 1471 1806
rect 1475 1802 1479 1806
rect 1483 1802 1535 1806
rect 1539 1802 1543 1806
rect 1547 1802 1599 1806
rect 1603 1802 1615 1806
rect 1619 1802 1663 1806
rect 1667 1802 1687 1806
rect 1691 1802 1727 1806
rect 1731 1802 1767 1806
rect 1771 1802 1783 1806
rect 1787 1802 1839 1806
rect 1843 1802 1863 1806
rect 1867 1802 1895 1806
rect 1899 1802 1959 1806
rect 1963 1802 1975 1806
rect 1979 1802 2095 1806
rect 2099 1802 2223 1806
rect 2227 1802 2359 1806
rect 2363 1802 2407 1806
rect 2411 1802 2435 1806
rect 1257 1801 2435 1802
rect 2441 1801 2442 1807
rect 96 1777 97 1783
rect 103 1782 1263 1783
rect 103 1778 111 1782
rect 115 1778 135 1782
rect 139 1778 175 1782
rect 179 1778 215 1782
rect 219 1778 271 1782
rect 275 1778 287 1782
rect 291 1778 351 1782
rect 355 1778 375 1782
rect 379 1778 439 1782
rect 443 1778 471 1782
rect 475 1778 535 1782
rect 539 1778 567 1782
rect 571 1778 631 1782
rect 635 1778 663 1782
rect 667 1778 727 1782
rect 731 1778 751 1782
rect 755 1778 823 1782
rect 827 1778 831 1782
rect 835 1778 903 1782
rect 907 1778 911 1782
rect 915 1778 967 1782
rect 971 1778 991 1782
rect 995 1778 1031 1782
rect 1035 1778 1063 1782
rect 1067 1778 1087 1782
rect 1091 1778 1135 1782
rect 1139 1778 1151 1782
rect 1155 1778 1191 1782
rect 1195 1778 1239 1782
rect 1243 1778 1263 1782
rect 103 1777 1263 1778
rect 1269 1777 1270 1783
rect 1262 1733 1263 1739
rect 1269 1738 2447 1739
rect 1269 1734 1279 1738
rect 1283 1734 1303 1738
rect 1307 1734 1351 1738
rect 1355 1734 1407 1738
rect 1411 1734 1423 1738
rect 1427 1734 1471 1738
rect 1475 1734 1503 1738
rect 1507 1734 1535 1738
rect 1539 1734 1583 1738
rect 1587 1734 1599 1738
rect 1603 1734 1663 1738
rect 1667 1734 1727 1738
rect 1731 1734 1735 1738
rect 1739 1734 1783 1738
rect 1787 1734 1807 1738
rect 1811 1734 1839 1738
rect 1843 1734 1871 1738
rect 1875 1734 1895 1738
rect 1899 1734 1935 1738
rect 1939 1734 1959 1738
rect 1963 1734 1999 1738
rect 2003 1734 2063 1738
rect 2067 1734 2407 1738
rect 2411 1734 2447 1738
rect 1269 1733 2447 1734
rect 2453 1733 2454 1739
rect 84 1705 85 1711
rect 91 1710 1251 1711
rect 91 1706 111 1710
rect 115 1706 135 1710
rect 139 1706 175 1710
rect 179 1706 215 1710
rect 219 1706 239 1710
rect 243 1706 287 1710
rect 291 1706 319 1710
rect 323 1706 375 1710
rect 379 1706 415 1710
rect 419 1706 471 1710
rect 475 1706 511 1710
rect 515 1706 567 1710
rect 571 1706 615 1710
rect 619 1706 663 1710
rect 667 1706 711 1710
rect 715 1706 751 1710
rect 755 1706 799 1710
rect 803 1706 831 1710
rect 835 1706 879 1710
rect 883 1706 903 1710
rect 907 1706 951 1710
rect 955 1706 967 1710
rect 971 1706 1015 1710
rect 1019 1706 1031 1710
rect 1035 1706 1087 1710
rect 1091 1706 1151 1710
rect 1155 1706 1159 1710
rect 1163 1706 1191 1710
rect 1195 1706 1239 1710
rect 1243 1706 1251 1710
rect 91 1705 1251 1706
rect 1257 1705 1258 1711
rect 1250 1665 1251 1671
rect 1257 1670 2435 1671
rect 1257 1666 1279 1670
rect 1283 1666 1303 1670
rect 1307 1666 1351 1670
rect 1355 1666 1359 1670
rect 1363 1666 1423 1670
rect 1427 1666 1447 1670
rect 1451 1666 1503 1670
rect 1507 1666 1543 1670
rect 1547 1666 1583 1670
rect 1587 1666 1639 1670
rect 1643 1666 1663 1670
rect 1667 1666 1727 1670
rect 1731 1666 1735 1670
rect 1739 1666 1807 1670
rect 1811 1666 1815 1670
rect 1819 1666 1871 1670
rect 1875 1666 1895 1670
rect 1899 1666 1935 1670
rect 1939 1666 1967 1670
rect 1971 1666 1999 1670
rect 2003 1666 2031 1670
rect 2035 1666 2063 1670
rect 2067 1666 2095 1670
rect 2099 1666 2159 1670
rect 2163 1666 2223 1670
rect 2227 1666 2407 1670
rect 2411 1666 2435 1670
rect 1257 1665 2435 1666
rect 2441 1665 2442 1671
rect 96 1633 97 1639
rect 103 1638 1263 1639
rect 103 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 175 1638
rect 179 1634 239 1638
rect 243 1634 271 1638
rect 275 1634 311 1638
rect 315 1634 319 1638
rect 323 1634 359 1638
rect 363 1634 415 1638
rect 419 1634 471 1638
rect 475 1634 511 1638
rect 515 1634 535 1638
rect 539 1634 599 1638
rect 603 1634 615 1638
rect 619 1634 663 1638
rect 667 1634 711 1638
rect 715 1634 719 1638
rect 723 1634 775 1638
rect 779 1634 799 1638
rect 803 1634 831 1638
rect 835 1634 879 1638
rect 883 1634 887 1638
rect 891 1634 943 1638
rect 947 1634 951 1638
rect 955 1634 999 1638
rect 1003 1634 1015 1638
rect 1019 1634 1087 1638
rect 1091 1634 1159 1638
rect 1163 1634 1239 1638
rect 1243 1634 1263 1638
rect 103 1633 1263 1634
rect 1269 1633 1270 1639
rect 1262 1597 1263 1603
rect 1269 1602 2447 1603
rect 1269 1598 1279 1602
rect 1283 1598 1303 1602
rect 1307 1598 1327 1602
rect 1331 1598 1359 1602
rect 1363 1598 1399 1602
rect 1403 1598 1447 1602
rect 1451 1598 1479 1602
rect 1483 1598 1543 1602
rect 1547 1598 1567 1602
rect 1571 1598 1639 1602
rect 1643 1598 1655 1602
rect 1659 1598 1727 1602
rect 1731 1598 1743 1602
rect 1747 1598 1815 1602
rect 1819 1598 1831 1602
rect 1835 1598 1895 1602
rect 1899 1598 1911 1602
rect 1915 1598 1967 1602
rect 1971 1598 1983 1602
rect 1987 1598 2031 1602
rect 2035 1598 2047 1602
rect 2051 1598 2095 1602
rect 2099 1598 2111 1602
rect 2115 1598 2159 1602
rect 2163 1598 2167 1602
rect 2171 1598 2215 1602
rect 2219 1598 2223 1602
rect 2227 1598 2271 1602
rect 2275 1598 2319 1602
rect 2323 1598 2359 1602
rect 2363 1598 2407 1602
rect 2411 1598 2447 1602
rect 1269 1597 2447 1598
rect 2453 1597 2454 1603
rect 84 1557 85 1563
rect 91 1562 1251 1563
rect 91 1558 111 1562
rect 115 1558 271 1562
rect 275 1558 311 1562
rect 315 1558 327 1562
rect 331 1558 359 1562
rect 363 1558 367 1562
rect 371 1558 407 1562
rect 411 1558 415 1562
rect 419 1558 447 1562
rect 451 1558 471 1562
rect 475 1558 487 1562
rect 491 1558 527 1562
rect 531 1558 535 1562
rect 539 1558 567 1562
rect 571 1558 599 1562
rect 603 1558 607 1562
rect 611 1558 647 1562
rect 651 1558 663 1562
rect 667 1558 687 1562
rect 691 1558 719 1562
rect 723 1558 727 1562
rect 731 1558 767 1562
rect 771 1558 775 1562
rect 779 1558 807 1562
rect 811 1558 831 1562
rect 835 1558 847 1562
rect 851 1558 887 1562
rect 891 1558 927 1562
rect 931 1558 943 1562
rect 947 1558 999 1562
rect 1003 1558 1239 1562
rect 1243 1558 1251 1562
rect 91 1557 1251 1558
rect 1257 1557 1258 1563
rect 1250 1525 1251 1531
rect 1257 1530 2435 1531
rect 1257 1526 1279 1530
rect 1283 1526 1327 1530
rect 1331 1526 1335 1530
rect 1339 1526 1399 1530
rect 1403 1526 1415 1530
rect 1419 1526 1479 1530
rect 1483 1526 1503 1530
rect 1507 1526 1567 1530
rect 1571 1526 1615 1530
rect 1619 1526 1655 1530
rect 1659 1526 1743 1530
rect 1747 1526 1831 1530
rect 1835 1526 1887 1530
rect 1891 1526 1911 1530
rect 1915 1526 1983 1530
rect 1987 1526 2047 1530
rect 2051 1526 2111 1530
rect 2115 1526 2167 1530
rect 2171 1526 2215 1530
rect 2219 1526 2271 1530
rect 2275 1526 2319 1530
rect 2323 1526 2359 1530
rect 2363 1526 2407 1530
rect 2411 1526 2435 1530
rect 1257 1525 2435 1526
rect 2441 1525 2442 1531
rect 1262 1457 1263 1463
rect 1269 1462 2447 1463
rect 1269 1458 1279 1462
rect 1283 1458 1335 1462
rect 1339 1458 1375 1462
rect 1379 1458 1415 1462
rect 1419 1458 1463 1462
rect 1467 1458 1503 1462
rect 1507 1458 1551 1462
rect 1555 1458 1615 1462
rect 1619 1458 1639 1462
rect 1643 1458 1727 1462
rect 1731 1458 1743 1462
rect 1747 1458 1807 1462
rect 1811 1458 1879 1462
rect 1883 1458 1887 1462
rect 1891 1458 1943 1462
rect 1947 1458 1999 1462
rect 2003 1458 2047 1462
rect 2051 1458 2095 1462
rect 2099 1458 2143 1462
rect 2147 1458 2191 1462
rect 2195 1458 2215 1462
rect 2219 1458 2239 1462
rect 2243 1458 2279 1462
rect 2283 1458 2319 1462
rect 2323 1458 2359 1462
rect 2363 1458 2407 1462
rect 2411 1458 2447 1462
rect 1269 1457 2447 1458
rect 2453 1457 2454 1463
rect 1262 1455 1270 1457
rect 96 1449 97 1455
rect 103 1454 1263 1455
rect 103 1450 111 1454
rect 115 1450 143 1454
rect 147 1450 183 1454
rect 187 1450 223 1454
rect 227 1450 263 1454
rect 267 1450 319 1454
rect 323 1450 327 1454
rect 331 1450 367 1454
rect 371 1450 391 1454
rect 395 1450 407 1454
rect 411 1450 447 1454
rect 451 1450 471 1454
rect 475 1450 487 1454
rect 491 1450 527 1454
rect 531 1450 559 1454
rect 563 1450 567 1454
rect 571 1450 607 1454
rect 611 1450 647 1454
rect 651 1450 687 1454
rect 691 1450 727 1454
rect 731 1450 767 1454
rect 771 1450 807 1454
rect 811 1450 847 1454
rect 851 1450 879 1454
rect 883 1450 887 1454
rect 891 1450 927 1454
rect 931 1450 943 1454
rect 947 1450 999 1454
rect 1003 1450 1047 1454
rect 1051 1450 1103 1454
rect 1107 1450 1151 1454
rect 1155 1450 1191 1454
rect 1195 1450 1239 1454
rect 1243 1450 1263 1454
rect 103 1449 1263 1450
rect 1269 1449 1270 1455
rect 84 1381 85 1387
rect 91 1386 1251 1387
rect 91 1382 111 1386
rect 115 1382 143 1386
rect 147 1382 167 1386
rect 171 1382 183 1386
rect 187 1382 207 1386
rect 211 1382 223 1386
rect 227 1382 247 1386
rect 251 1382 263 1386
rect 267 1382 303 1386
rect 307 1382 319 1386
rect 323 1382 367 1386
rect 371 1382 391 1386
rect 395 1382 439 1386
rect 443 1382 471 1386
rect 475 1382 519 1386
rect 523 1382 559 1386
rect 563 1382 599 1386
rect 603 1382 647 1386
rect 651 1382 679 1386
rect 683 1382 727 1386
rect 731 1382 751 1386
rect 755 1382 807 1386
rect 811 1382 823 1386
rect 827 1382 879 1386
rect 883 1382 887 1386
rect 891 1382 943 1386
rect 947 1382 951 1386
rect 955 1382 999 1386
rect 1003 1382 1015 1386
rect 1019 1382 1047 1386
rect 1051 1382 1079 1386
rect 1083 1382 1103 1386
rect 1107 1382 1143 1386
rect 1147 1382 1151 1386
rect 1155 1382 1191 1386
rect 1195 1382 1239 1386
rect 1243 1382 1251 1386
rect 91 1381 1251 1382
rect 1257 1386 2442 1387
rect 1257 1382 1279 1386
rect 1283 1382 1303 1386
rect 1307 1382 1343 1386
rect 1347 1382 1375 1386
rect 1379 1382 1399 1386
rect 1403 1382 1463 1386
rect 1467 1382 1535 1386
rect 1539 1382 1551 1386
rect 1555 1382 1607 1386
rect 1611 1382 1639 1386
rect 1643 1382 1687 1386
rect 1691 1382 1727 1386
rect 1731 1382 1767 1386
rect 1771 1382 1807 1386
rect 1811 1382 1847 1386
rect 1851 1382 1879 1386
rect 1883 1382 1935 1386
rect 1939 1382 1943 1386
rect 1947 1382 1999 1386
rect 2003 1382 2023 1386
rect 2027 1382 2047 1386
rect 2051 1382 2095 1386
rect 2099 1382 2111 1386
rect 2115 1382 2143 1386
rect 2147 1382 2191 1386
rect 2195 1382 2199 1386
rect 2203 1382 2239 1386
rect 2243 1382 2279 1386
rect 2283 1382 2287 1386
rect 2291 1382 2319 1386
rect 2323 1382 2359 1386
rect 2363 1382 2407 1386
rect 2411 1382 2442 1386
rect 1257 1381 2442 1382
rect 1262 1318 2454 1319
rect 1262 1315 1279 1318
rect 96 1309 97 1315
rect 103 1314 1263 1315
rect 103 1310 111 1314
rect 115 1310 167 1314
rect 171 1310 183 1314
rect 187 1310 207 1314
rect 211 1310 231 1314
rect 235 1310 247 1314
rect 251 1310 287 1314
rect 291 1310 303 1314
rect 307 1310 351 1314
rect 355 1310 367 1314
rect 371 1310 423 1314
rect 427 1310 439 1314
rect 443 1310 495 1314
rect 499 1310 519 1314
rect 523 1310 567 1314
rect 571 1310 599 1314
rect 603 1310 639 1314
rect 643 1310 679 1314
rect 683 1310 703 1314
rect 707 1310 751 1314
rect 755 1310 767 1314
rect 771 1310 823 1314
rect 827 1310 879 1314
rect 883 1310 887 1314
rect 891 1310 935 1314
rect 939 1310 951 1314
rect 955 1310 999 1314
rect 1003 1310 1015 1314
rect 1019 1310 1079 1314
rect 1083 1310 1143 1314
rect 1147 1310 1191 1314
rect 1195 1310 1239 1314
rect 1243 1310 1263 1314
rect 103 1309 1263 1310
rect 1269 1314 1279 1315
rect 1283 1314 1303 1318
rect 1307 1314 1343 1318
rect 1347 1314 1383 1318
rect 1387 1314 1399 1318
rect 1403 1314 1423 1318
rect 1427 1314 1463 1318
rect 1467 1314 1503 1318
rect 1507 1314 1535 1318
rect 1539 1314 1543 1318
rect 1547 1314 1583 1318
rect 1587 1314 1607 1318
rect 1611 1314 1623 1318
rect 1627 1314 1679 1318
rect 1683 1314 1687 1318
rect 1691 1314 1735 1318
rect 1739 1314 1767 1318
rect 1771 1314 1791 1318
rect 1795 1314 1847 1318
rect 1851 1314 1903 1318
rect 1907 1314 1935 1318
rect 1939 1314 1967 1318
rect 1971 1314 2023 1318
rect 2027 1314 2039 1318
rect 2043 1314 2111 1318
rect 2115 1314 2119 1318
rect 2123 1314 2199 1318
rect 2203 1314 2287 1318
rect 2291 1314 2359 1318
rect 2363 1314 2407 1318
rect 2411 1314 2454 1318
rect 1269 1313 2454 1314
rect 1269 1309 1270 1313
rect 84 1237 85 1243
rect 91 1242 1251 1243
rect 91 1238 111 1242
rect 115 1238 135 1242
rect 139 1238 175 1242
rect 179 1238 183 1242
rect 187 1238 231 1242
rect 235 1238 287 1242
rect 291 1238 311 1242
rect 315 1238 351 1242
rect 355 1238 399 1242
rect 403 1238 423 1242
rect 427 1238 487 1242
rect 491 1238 495 1242
rect 499 1238 567 1242
rect 571 1238 575 1242
rect 579 1238 639 1242
rect 643 1238 663 1242
rect 667 1238 703 1242
rect 707 1238 743 1242
rect 747 1238 767 1242
rect 771 1238 815 1242
rect 819 1238 823 1242
rect 827 1238 879 1242
rect 883 1238 935 1242
rect 939 1238 943 1242
rect 947 1238 999 1242
rect 1003 1238 1007 1242
rect 1011 1238 1071 1242
rect 1075 1238 1239 1242
rect 1243 1238 1251 1242
rect 91 1237 1251 1238
rect 1257 1242 2442 1243
rect 1257 1238 1279 1242
rect 1283 1238 1303 1242
rect 1307 1238 1343 1242
rect 1347 1238 1375 1242
rect 1379 1238 1383 1242
rect 1387 1238 1423 1242
rect 1427 1238 1463 1242
rect 1467 1238 1479 1242
rect 1483 1238 1503 1242
rect 1507 1238 1543 1242
rect 1547 1238 1583 1242
rect 1587 1238 1623 1242
rect 1627 1238 1679 1242
rect 1683 1238 1687 1242
rect 1691 1238 1735 1242
rect 1739 1238 1791 1242
rect 1795 1238 1847 1242
rect 1851 1238 1887 1242
rect 1891 1238 1903 1242
rect 1907 1238 1967 1242
rect 1971 1238 1983 1242
rect 1987 1238 2039 1242
rect 2043 1238 2071 1242
rect 2075 1238 2119 1242
rect 2123 1238 2151 1242
rect 2155 1238 2199 1242
rect 2203 1238 2223 1242
rect 2227 1238 2287 1242
rect 2291 1238 2303 1242
rect 2307 1238 2359 1242
rect 2363 1238 2407 1242
rect 2411 1238 2442 1242
rect 1257 1237 2442 1238
rect 96 1169 97 1175
rect 103 1174 1263 1175
rect 103 1170 111 1174
rect 115 1170 135 1174
rect 139 1170 175 1174
rect 179 1170 231 1174
rect 235 1170 239 1174
rect 243 1170 311 1174
rect 315 1170 327 1174
rect 331 1170 399 1174
rect 403 1170 431 1174
rect 435 1170 487 1174
rect 491 1170 535 1174
rect 539 1170 575 1174
rect 579 1170 639 1174
rect 643 1170 663 1174
rect 667 1170 743 1174
rect 747 1170 815 1174
rect 819 1170 839 1174
rect 843 1170 879 1174
rect 883 1170 919 1174
rect 923 1170 943 1174
rect 947 1170 999 1174
rect 1003 1170 1007 1174
rect 1011 1170 1071 1174
rect 1075 1170 1143 1174
rect 1147 1170 1191 1174
rect 1195 1170 1239 1174
rect 1243 1170 1263 1174
rect 103 1169 1263 1170
rect 1269 1174 2454 1175
rect 1269 1170 1279 1174
rect 1283 1170 1303 1174
rect 1307 1170 1343 1174
rect 1347 1170 1375 1174
rect 1379 1170 1407 1174
rect 1411 1170 1479 1174
rect 1483 1170 1487 1174
rect 1491 1170 1583 1174
rect 1587 1170 1687 1174
rect 1691 1170 1791 1174
rect 1795 1170 1799 1174
rect 1803 1170 1887 1174
rect 1891 1170 1903 1174
rect 1907 1170 1983 1174
rect 1987 1170 1999 1174
rect 2003 1170 2071 1174
rect 2075 1170 2079 1174
rect 2083 1170 2151 1174
rect 2155 1170 2159 1174
rect 2163 1170 2223 1174
rect 2227 1170 2231 1174
rect 2235 1170 2303 1174
rect 2307 1170 2359 1174
rect 2363 1170 2407 1174
rect 2411 1170 2454 1174
rect 1269 1169 2454 1170
rect 1250 1106 2442 1107
rect 1250 1103 1279 1106
rect 84 1097 85 1103
rect 91 1102 1251 1103
rect 91 1098 111 1102
rect 115 1098 135 1102
rect 139 1098 175 1102
rect 179 1098 239 1102
rect 243 1098 247 1102
rect 251 1098 327 1102
rect 331 1098 415 1102
rect 419 1098 431 1102
rect 435 1098 503 1102
rect 507 1098 535 1102
rect 539 1098 583 1102
rect 587 1098 639 1102
rect 643 1098 663 1102
rect 667 1098 735 1102
rect 739 1098 743 1102
rect 747 1098 799 1102
rect 803 1098 839 1102
rect 843 1098 863 1102
rect 867 1098 919 1102
rect 923 1098 983 1102
rect 987 1098 999 1102
rect 1003 1098 1047 1102
rect 1051 1098 1071 1102
rect 1075 1098 1143 1102
rect 1147 1098 1191 1102
rect 1195 1098 1239 1102
rect 1243 1098 1251 1102
rect 91 1097 1251 1098
rect 1257 1102 1279 1103
rect 1283 1102 1303 1106
rect 1307 1102 1343 1106
rect 1347 1102 1407 1106
rect 1411 1102 1431 1106
rect 1435 1102 1471 1106
rect 1475 1102 1487 1106
rect 1491 1102 1511 1106
rect 1515 1102 1559 1106
rect 1563 1102 1583 1106
rect 1587 1102 1615 1106
rect 1619 1102 1671 1106
rect 1675 1102 1687 1106
rect 1691 1102 1727 1106
rect 1731 1102 1775 1106
rect 1779 1102 1799 1106
rect 1803 1102 1823 1106
rect 1827 1102 1871 1106
rect 1875 1102 1903 1106
rect 1907 1102 1919 1106
rect 1923 1102 1967 1106
rect 1971 1102 1999 1106
rect 2003 1102 2015 1106
rect 2019 1102 2063 1106
rect 2067 1102 2079 1106
rect 2083 1102 2119 1106
rect 2123 1102 2159 1106
rect 2163 1102 2175 1106
rect 2179 1102 2231 1106
rect 2235 1102 2303 1106
rect 2307 1102 2359 1106
rect 2363 1102 2407 1106
rect 2411 1102 2442 1106
rect 1257 1101 2442 1102
rect 1257 1097 1258 1101
rect 1262 1038 2454 1039
rect 1262 1035 1279 1038
rect 96 1029 97 1035
rect 103 1034 1263 1035
rect 103 1030 111 1034
rect 115 1030 135 1034
rect 139 1030 175 1034
rect 179 1030 247 1034
rect 251 1030 255 1034
rect 259 1030 327 1034
rect 331 1030 399 1034
rect 403 1030 415 1034
rect 419 1030 463 1034
rect 467 1030 503 1034
rect 507 1030 519 1034
rect 523 1030 575 1034
rect 579 1030 583 1034
rect 587 1030 623 1034
rect 627 1030 663 1034
rect 667 1030 671 1034
rect 675 1030 735 1034
rect 739 1030 799 1034
rect 803 1030 807 1034
rect 811 1030 863 1034
rect 867 1030 895 1034
rect 899 1030 919 1034
rect 923 1030 983 1034
rect 987 1030 999 1034
rect 1003 1030 1047 1034
rect 1051 1030 1103 1034
rect 1107 1030 1191 1034
rect 1195 1030 1239 1034
rect 1243 1030 1263 1034
rect 103 1029 1263 1030
rect 1269 1034 1279 1035
rect 1283 1034 1431 1038
rect 1435 1034 1471 1038
rect 1475 1034 1511 1038
rect 1515 1034 1559 1038
rect 1563 1034 1575 1038
rect 1579 1034 1615 1038
rect 1619 1034 1655 1038
rect 1659 1034 1671 1038
rect 1675 1034 1695 1038
rect 1699 1034 1727 1038
rect 1731 1034 1735 1038
rect 1739 1034 1775 1038
rect 1779 1034 1823 1038
rect 1827 1034 1871 1038
rect 1875 1034 1879 1038
rect 1883 1034 1919 1038
rect 1923 1034 1943 1038
rect 1947 1034 1967 1038
rect 1971 1034 2015 1038
rect 2019 1034 2063 1038
rect 2067 1034 2095 1038
rect 2099 1034 2119 1038
rect 2123 1034 2175 1038
rect 2179 1034 2231 1038
rect 2235 1034 2255 1038
rect 2259 1034 2407 1038
rect 2411 1034 2454 1038
rect 1269 1033 2454 1034
rect 1269 1029 1270 1033
rect 84 961 85 967
rect 91 966 1251 967
rect 91 962 111 966
rect 115 962 175 966
rect 179 962 215 966
rect 219 962 255 966
rect 259 962 303 966
rect 307 962 327 966
rect 331 962 359 966
rect 363 962 399 966
rect 403 962 415 966
rect 419 962 463 966
rect 467 962 519 966
rect 523 962 575 966
rect 579 962 623 966
rect 627 962 639 966
rect 643 962 671 966
rect 675 962 711 966
rect 715 962 735 966
rect 739 962 783 966
rect 787 962 807 966
rect 811 962 855 966
rect 859 962 895 966
rect 899 962 927 966
rect 931 962 999 966
rect 1003 962 1071 966
rect 1075 962 1103 966
rect 1107 962 1143 966
rect 1147 962 1191 966
rect 1195 962 1239 966
rect 1243 962 1251 966
rect 91 961 1251 962
rect 1257 963 1258 967
rect 1257 962 2442 963
rect 1257 961 1279 962
rect 1250 958 1279 961
rect 1283 958 1303 962
rect 1307 958 1351 962
rect 1355 958 1431 962
rect 1435 958 1511 962
rect 1515 958 1575 962
rect 1579 958 1591 962
rect 1595 958 1615 962
rect 1619 958 1655 962
rect 1659 958 1679 962
rect 1683 958 1695 962
rect 1699 958 1735 962
rect 1739 958 1767 962
rect 1771 958 1775 962
rect 1779 958 1823 962
rect 1827 958 1855 962
rect 1859 958 1879 962
rect 1883 958 1943 962
rect 1947 958 2015 962
rect 2019 958 2023 962
rect 2027 958 2095 962
rect 2099 958 2103 962
rect 2107 958 2175 962
rect 2179 958 2183 962
rect 2187 958 2255 962
rect 2259 958 2271 962
rect 2275 958 2407 962
rect 2411 958 2442 962
rect 1250 957 2442 958
rect 1262 894 2454 895
rect 1262 891 1279 894
rect 96 885 97 891
rect 103 890 1263 891
rect 103 886 111 890
rect 115 886 191 890
rect 195 886 215 890
rect 219 886 231 890
rect 235 886 255 890
rect 259 886 287 890
rect 291 886 303 890
rect 307 886 359 890
rect 363 886 415 890
rect 419 886 447 890
rect 451 886 463 890
rect 467 886 519 890
rect 523 886 543 890
rect 547 886 575 890
rect 579 886 639 890
rect 643 886 711 890
rect 715 886 727 890
rect 731 886 783 890
rect 787 886 807 890
rect 811 886 855 890
rect 859 886 887 890
rect 891 886 927 890
rect 931 886 959 890
rect 963 886 999 890
rect 1003 886 1023 890
rect 1027 886 1071 890
rect 1075 886 1087 890
rect 1091 886 1143 890
rect 1147 886 1159 890
rect 1163 886 1191 890
rect 1195 886 1239 890
rect 1243 886 1263 890
rect 103 885 1263 886
rect 1269 890 1279 891
rect 1283 890 1303 894
rect 1307 890 1351 894
rect 1355 890 1431 894
rect 1435 890 1439 894
rect 1443 890 1479 894
rect 1483 890 1511 894
rect 1515 890 1519 894
rect 1523 890 1559 894
rect 1563 890 1591 894
rect 1595 890 1607 894
rect 1611 890 1655 894
rect 1659 890 1679 894
rect 1683 890 1711 894
rect 1715 890 1767 894
rect 1771 890 1775 894
rect 1779 890 1847 894
rect 1851 890 1855 894
rect 1859 890 1919 894
rect 1923 890 1943 894
rect 1947 890 1991 894
rect 1995 890 2023 894
rect 2027 890 2063 894
rect 2067 890 2103 894
rect 2107 890 2135 894
rect 2139 890 2183 894
rect 2187 890 2215 894
rect 2219 890 2271 894
rect 2275 890 2295 894
rect 2299 890 2407 894
rect 2411 890 2454 894
rect 1269 889 2454 890
rect 1269 885 1270 889
rect 84 817 85 823
rect 91 822 1251 823
rect 91 818 111 822
rect 115 818 135 822
rect 139 818 175 822
rect 179 818 191 822
rect 195 818 231 822
rect 235 818 239 822
rect 243 818 287 822
rect 291 818 327 822
rect 331 818 359 822
rect 363 818 415 822
rect 419 818 447 822
rect 451 818 503 822
rect 507 818 543 822
rect 547 818 591 822
rect 595 818 639 822
rect 643 818 671 822
rect 675 818 727 822
rect 731 818 743 822
rect 747 818 807 822
rect 811 818 815 822
rect 819 818 879 822
rect 883 818 887 822
rect 891 818 943 822
rect 947 818 959 822
rect 963 818 1015 822
rect 1019 818 1023 822
rect 1027 818 1087 822
rect 1091 818 1159 822
rect 1163 818 1239 822
rect 1243 818 1251 822
rect 91 817 1251 818
rect 1257 817 1258 823
rect 1250 815 1258 817
rect 1250 809 1251 815
rect 1257 814 2435 815
rect 1257 810 1279 814
rect 1283 810 1359 814
rect 1363 810 1415 814
rect 1419 810 1439 814
rect 1443 810 1471 814
rect 1475 810 1479 814
rect 1483 810 1519 814
rect 1523 810 1535 814
rect 1539 810 1559 814
rect 1563 810 1591 814
rect 1595 810 1607 814
rect 1611 810 1647 814
rect 1651 810 1655 814
rect 1659 810 1703 814
rect 1707 810 1711 814
rect 1715 810 1759 814
rect 1763 810 1775 814
rect 1779 810 1815 814
rect 1819 810 1847 814
rect 1851 810 1871 814
rect 1875 810 1919 814
rect 1923 810 1935 814
rect 1939 810 1991 814
rect 1995 810 1999 814
rect 2003 810 2063 814
rect 2067 810 2071 814
rect 2075 810 2135 814
rect 2139 810 2143 814
rect 2147 810 2215 814
rect 2219 810 2223 814
rect 2227 810 2295 814
rect 2299 810 2303 814
rect 2307 810 2359 814
rect 2363 810 2407 814
rect 2411 810 2435 814
rect 1257 809 2435 810
rect 2441 809 2442 815
rect 96 745 97 751
rect 103 750 1263 751
rect 103 746 111 750
rect 115 746 135 750
rect 139 746 175 750
rect 179 746 191 750
rect 195 746 239 750
rect 243 746 263 750
rect 267 746 327 750
rect 331 746 335 750
rect 339 746 399 750
rect 403 746 415 750
rect 419 746 455 750
rect 459 746 503 750
rect 507 746 543 750
rect 547 746 583 750
rect 587 746 591 750
rect 595 746 623 750
rect 627 746 671 750
rect 675 746 719 750
rect 723 746 743 750
rect 747 746 767 750
rect 771 746 815 750
rect 819 746 863 750
rect 867 746 879 750
rect 883 746 911 750
rect 915 746 943 750
rect 947 746 1015 750
rect 1019 746 1239 750
rect 1243 746 1263 750
rect 103 745 1263 746
rect 1269 747 1270 751
rect 1269 746 2454 747
rect 1269 745 1279 746
rect 1262 742 1279 745
rect 1283 742 1303 746
rect 1307 742 1343 746
rect 1347 742 1359 746
rect 1363 742 1407 746
rect 1411 742 1415 746
rect 1419 742 1471 746
rect 1475 742 1487 746
rect 1491 742 1535 746
rect 1539 742 1575 746
rect 1579 742 1591 746
rect 1595 742 1647 746
rect 1651 742 1663 746
rect 1667 742 1703 746
rect 1707 742 1751 746
rect 1755 742 1759 746
rect 1763 742 1815 746
rect 1819 742 1831 746
rect 1835 742 1871 746
rect 1875 742 1911 746
rect 1915 742 1935 746
rect 1939 742 1991 746
rect 1995 742 1999 746
rect 2003 742 2071 746
rect 2075 742 2079 746
rect 2083 742 2143 746
rect 2147 742 2175 746
rect 2179 742 2223 746
rect 2227 742 2279 746
rect 2283 742 2303 746
rect 2307 742 2359 746
rect 2363 742 2407 746
rect 2411 742 2454 746
rect 1262 741 2454 742
rect 84 673 85 679
rect 91 678 1251 679
rect 91 674 111 678
rect 115 674 135 678
rect 139 674 191 678
rect 195 674 199 678
rect 203 674 263 678
rect 267 674 279 678
rect 283 674 335 678
rect 339 674 351 678
rect 355 674 399 678
rect 403 674 415 678
rect 419 674 455 678
rect 459 674 487 678
rect 491 674 503 678
rect 507 674 543 678
rect 547 674 559 678
rect 563 674 583 678
rect 587 674 623 678
rect 627 674 639 678
rect 643 674 671 678
rect 675 674 711 678
rect 715 674 719 678
rect 723 674 767 678
rect 771 674 783 678
rect 787 674 815 678
rect 819 674 855 678
rect 859 674 863 678
rect 867 674 911 678
rect 915 674 919 678
rect 923 674 983 678
rect 987 674 1039 678
rect 1043 674 1095 678
rect 1099 674 1151 678
rect 1155 674 1191 678
rect 1195 674 1239 678
rect 1243 674 1251 678
rect 91 673 1251 674
rect 1257 675 1258 679
rect 1257 674 2442 675
rect 1257 673 1279 674
rect 1250 670 1279 673
rect 1283 670 1303 674
rect 1307 670 1343 674
rect 1347 670 1399 674
rect 1403 670 1407 674
rect 1411 670 1487 674
rect 1491 670 1511 674
rect 1515 670 1575 674
rect 1579 670 1623 674
rect 1627 670 1663 674
rect 1667 670 1727 674
rect 1731 670 1751 674
rect 1755 670 1815 674
rect 1819 670 1831 674
rect 1835 670 1895 674
rect 1899 670 1911 674
rect 1915 670 1975 674
rect 1979 670 1991 674
rect 1995 670 2047 674
rect 2051 670 2079 674
rect 2083 670 2111 674
rect 2115 670 2175 674
rect 2179 670 2239 674
rect 2243 670 2279 674
rect 2283 670 2311 674
rect 2315 670 2359 674
rect 2363 670 2407 674
rect 2411 670 2442 674
rect 1250 669 2442 670
rect 96 597 97 603
rect 103 602 1263 603
rect 103 598 111 602
rect 115 598 135 602
rect 139 598 191 602
rect 195 598 199 602
rect 203 598 271 602
rect 275 598 279 602
rect 283 598 351 602
rect 355 598 359 602
rect 363 598 415 602
rect 419 598 447 602
rect 451 598 487 602
rect 491 598 535 602
rect 539 598 559 602
rect 563 598 623 602
rect 627 598 639 602
rect 643 598 703 602
rect 707 598 711 602
rect 715 598 783 602
rect 787 598 855 602
rect 859 598 919 602
rect 923 598 975 602
rect 979 598 983 602
rect 987 598 1023 602
rect 1027 598 1039 602
rect 1043 598 1079 602
rect 1083 598 1095 602
rect 1099 598 1135 602
rect 1139 598 1151 602
rect 1155 598 1191 602
rect 1195 598 1239 602
rect 1243 598 1263 602
rect 103 597 1263 598
rect 1269 602 2454 603
rect 1269 598 1279 602
rect 1283 598 1303 602
rect 1307 598 1399 602
rect 1403 598 1415 602
rect 1419 598 1455 602
rect 1459 598 1495 602
rect 1499 598 1511 602
rect 1515 598 1543 602
rect 1547 598 1599 602
rect 1603 598 1623 602
rect 1627 598 1663 602
rect 1667 598 1727 602
rect 1731 598 1791 602
rect 1795 598 1815 602
rect 1819 598 1847 602
rect 1851 598 1895 602
rect 1899 598 1911 602
rect 1915 598 1975 602
rect 1979 598 2047 602
rect 2051 598 2111 602
rect 2115 598 2119 602
rect 2123 598 2175 602
rect 2179 598 2199 602
rect 2203 598 2239 602
rect 2243 598 2287 602
rect 2291 598 2311 602
rect 2315 598 2359 602
rect 2363 598 2407 602
rect 2411 598 2454 602
rect 1269 597 2454 598
rect 1250 529 1251 535
rect 1257 534 2435 535
rect 1257 530 1279 534
rect 1283 530 1303 534
rect 1307 530 1375 534
rect 1379 530 1415 534
rect 1419 530 1455 534
rect 1459 530 1479 534
rect 1483 530 1495 534
rect 1499 530 1543 534
rect 1547 530 1583 534
rect 1587 530 1599 534
rect 1603 530 1663 534
rect 1667 530 1695 534
rect 1699 530 1727 534
rect 1731 530 1791 534
rect 1795 530 1799 534
rect 1803 530 1847 534
rect 1851 530 1903 534
rect 1907 530 1911 534
rect 1915 530 1975 534
rect 1979 530 2007 534
rect 2011 530 2047 534
rect 2051 530 2103 534
rect 2107 530 2119 534
rect 2123 530 2191 534
rect 2195 530 2199 534
rect 2203 530 2287 534
rect 2291 530 2359 534
rect 2363 530 2407 534
rect 2411 530 2435 534
rect 1257 529 2435 530
rect 2441 529 2442 535
rect 1250 527 1258 529
rect 84 521 85 527
rect 91 526 1251 527
rect 91 522 111 526
rect 115 522 135 526
rect 139 522 191 526
rect 195 522 263 526
rect 267 522 271 526
rect 275 522 335 526
rect 339 522 359 526
rect 363 522 415 526
rect 419 522 447 526
rect 451 522 495 526
rect 499 522 535 526
rect 539 522 575 526
rect 579 522 623 526
rect 627 522 647 526
rect 651 522 703 526
rect 707 522 719 526
rect 723 522 783 526
rect 787 522 847 526
rect 851 522 855 526
rect 859 522 903 526
rect 907 522 919 526
rect 923 522 959 526
rect 963 522 975 526
rect 979 522 1023 526
rect 1027 522 1079 526
rect 1083 522 1087 526
rect 1091 522 1135 526
rect 1139 522 1151 526
rect 1155 522 1191 526
rect 1195 522 1239 526
rect 1243 522 1251 526
rect 91 521 1251 522
rect 1257 521 1258 527
rect 1262 462 2454 463
rect 1262 459 1279 462
rect 96 453 97 459
rect 103 458 1263 459
rect 103 454 111 458
rect 115 454 135 458
rect 139 454 183 458
rect 187 454 191 458
rect 195 454 223 458
rect 227 454 263 458
rect 267 454 311 458
rect 315 454 335 458
rect 339 454 367 458
rect 371 454 415 458
rect 419 454 431 458
rect 435 454 495 458
rect 499 454 559 458
rect 563 454 575 458
rect 579 454 615 458
rect 619 454 647 458
rect 651 454 671 458
rect 675 454 719 458
rect 723 454 775 458
rect 779 454 783 458
rect 787 454 831 458
rect 835 454 847 458
rect 851 454 887 458
rect 891 454 903 458
rect 907 454 959 458
rect 963 454 1023 458
rect 1027 454 1087 458
rect 1091 454 1151 458
rect 1155 454 1191 458
rect 1195 454 1239 458
rect 1243 454 1263 458
rect 103 453 1263 454
rect 1269 458 1279 459
rect 1283 458 1303 462
rect 1307 458 1343 462
rect 1347 458 1375 462
rect 1379 458 1399 462
rect 1403 458 1463 462
rect 1467 458 1479 462
rect 1483 458 1527 462
rect 1531 458 1583 462
rect 1587 458 1591 462
rect 1595 458 1663 462
rect 1667 458 1695 462
rect 1699 458 1735 462
rect 1739 458 1799 462
rect 1803 458 1815 462
rect 1819 458 1895 462
rect 1899 458 1903 462
rect 1907 458 1975 462
rect 1979 458 2007 462
rect 2011 458 2055 462
rect 2059 458 2103 462
rect 2107 458 2135 462
rect 2139 458 2191 462
rect 2195 458 2215 462
rect 2219 458 2287 462
rect 2291 458 2295 462
rect 2299 458 2359 462
rect 2363 458 2407 462
rect 2411 458 2454 462
rect 1269 457 2454 458
rect 1269 453 1270 457
rect 84 385 85 391
rect 91 390 1251 391
rect 91 386 111 390
rect 115 386 135 390
rect 139 386 175 390
rect 179 386 183 390
rect 187 386 223 390
rect 227 386 231 390
rect 235 386 263 390
rect 267 386 287 390
rect 291 386 311 390
rect 315 386 343 390
rect 347 386 367 390
rect 371 386 391 390
rect 395 386 431 390
rect 435 386 439 390
rect 443 386 487 390
rect 491 386 495 390
rect 499 386 535 390
rect 539 386 559 390
rect 563 386 583 390
rect 587 386 615 390
rect 619 386 631 390
rect 635 386 671 390
rect 675 386 679 390
rect 683 386 719 390
rect 723 386 727 390
rect 731 386 775 390
rect 779 386 831 390
rect 835 386 887 390
rect 891 386 1239 390
rect 1243 386 1251 390
rect 91 385 1251 386
rect 1257 390 2442 391
rect 1257 386 1279 390
rect 1283 386 1303 390
rect 1307 386 1343 390
rect 1347 386 1399 390
rect 1403 386 1447 390
rect 1451 386 1463 390
rect 1467 386 1487 390
rect 1491 386 1527 390
rect 1531 386 1535 390
rect 1539 386 1591 390
rect 1595 386 1663 390
rect 1667 386 1735 390
rect 1739 386 1815 390
rect 1819 386 1895 390
rect 1899 386 1967 390
rect 1971 386 1975 390
rect 1979 386 2039 390
rect 2043 386 2055 390
rect 2059 386 2111 390
rect 2115 386 2135 390
rect 2139 386 2175 390
rect 2179 386 2215 390
rect 2219 386 2239 390
rect 2243 386 2295 390
rect 2299 386 2303 390
rect 2307 386 2359 390
rect 2363 386 2407 390
rect 2411 386 2442 390
rect 1257 385 2442 386
rect 96 313 97 319
rect 103 318 1263 319
rect 103 314 111 318
rect 115 314 135 318
rect 139 314 175 318
rect 179 314 183 318
rect 187 314 231 318
rect 235 314 255 318
rect 259 314 287 318
rect 291 314 327 318
rect 331 314 343 318
rect 347 314 391 318
rect 395 314 439 318
rect 443 314 447 318
rect 451 314 487 318
rect 491 314 503 318
rect 507 314 535 318
rect 539 314 551 318
rect 555 314 583 318
rect 587 314 591 318
rect 595 314 631 318
rect 635 314 679 318
rect 683 314 727 318
rect 731 314 775 318
rect 779 314 823 318
rect 827 314 871 318
rect 875 314 919 318
rect 923 314 1239 318
rect 1243 314 1263 318
rect 103 313 1263 314
rect 1269 318 2454 319
rect 1269 314 1279 318
rect 1283 314 1447 318
rect 1451 314 1487 318
rect 1491 314 1495 318
rect 1499 314 1535 318
rect 1539 314 1575 318
rect 1579 314 1591 318
rect 1595 314 1615 318
rect 1619 314 1655 318
rect 1659 314 1663 318
rect 1667 314 1695 318
rect 1699 314 1735 318
rect 1739 314 1743 318
rect 1747 314 1799 318
rect 1803 314 1815 318
rect 1819 314 1863 318
rect 1867 314 1895 318
rect 1899 314 1935 318
rect 1939 314 1967 318
rect 1971 314 2007 318
rect 2011 314 2039 318
rect 2043 314 2071 318
rect 2075 314 2111 318
rect 2115 314 2135 318
rect 2139 314 2175 318
rect 2179 314 2191 318
rect 2195 314 2239 318
rect 2243 314 2255 318
rect 2259 314 2303 318
rect 2307 314 2319 318
rect 2323 314 2359 318
rect 2363 314 2407 318
rect 2411 314 2454 318
rect 1269 313 2454 314
rect 1250 246 2442 247
rect 1250 243 1279 246
rect 84 237 85 243
rect 91 242 1251 243
rect 91 238 111 242
rect 115 238 135 242
rect 139 238 175 242
rect 179 238 183 242
rect 187 238 247 242
rect 251 238 255 242
rect 259 238 327 242
rect 331 238 391 242
rect 395 238 415 242
rect 419 238 447 242
rect 451 238 495 242
rect 499 238 503 242
rect 507 238 551 242
rect 555 238 575 242
rect 579 238 591 242
rect 595 238 631 242
rect 635 238 655 242
rect 659 238 679 242
rect 683 238 727 242
rect 731 238 775 242
rect 779 238 791 242
rect 795 238 823 242
rect 827 238 847 242
rect 851 238 871 242
rect 875 238 903 242
rect 907 238 919 242
rect 923 238 959 242
rect 963 238 1023 242
rect 1027 238 1239 242
rect 1243 238 1251 242
rect 91 237 1251 238
rect 1257 242 1279 243
rect 1283 242 1367 246
rect 1371 242 1407 246
rect 1411 242 1447 246
rect 1451 242 1495 246
rect 1499 242 1535 246
rect 1539 242 1551 246
rect 1555 242 1575 246
rect 1579 242 1607 246
rect 1611 242 1615 246
rect 1619 242 1655 246
rect 1659 242 1671 246
rect 1675 242 1695 246
rect 1699 242 1735 246
rect 1739 242 1743 246
rect 1747 242 1799 246
rect 1803 242 1807 246
rect 1811 242 1863 246
rect 1867 242 1887 246
rect 1891 242 1935 246
rect 1939 242 1975 246
rect 1979 242 2007 246
rect 2011 242 2071 246
rect 2075 242 2135 246
rect 2139 242 2167 246
rect 2171 242 2191 246
rect 2195 242 2255 246
rect 2259 242 2271 246
rect 2275 242 2319 246
rect 2323 242 2359 246
rect 2363 242 2407 246
rect 2411 242 2442 246
rect 1257 241 2442 242
rect 1257 237 1258 241
rect 1262 157 1263 163
rect 1269 162 2447 163
rect 1269 158 1279 162
rect 1283 158 1303 162
rect 1307 158 1343 162
rect 1347 158 1367 162
rect 1371 158 1383 162
rect 1387 158 1407 162
rect 1411 158 1423 162
rect 1427 158 1447 162
rect 1451 158 1463 162
rect 1467 158 1495 162
rect 1499 158 1519 162
rect 1523 158 1551 162
rect 1555 158 1583 162
rect 1587 158 1607 162
rect 1611 158 1647 162
rect 1651 158 1671 162
rect 1675 158 1711 162
rect 1715 158 1735 162
rect 1739 158 1767 162
rect 1771 158 1807 162
rect 1811 158 1823 162
rect 1827 158 1871 162
rect 1875 158 1887 162
rect 1891 158 1919 162
rect 1923 158 1967 162
rect 1971 158 1975 162
rect 1979 158 2015 162
rect 2019 158 2063 162
rect 2067 158 2071 162
rect 2075 158 2111 162
rect 2115 158 2159 162
rect 2163 158 2167 162
rect 2171 158 2215 162
rect 2219 158 2271 162
rect 2275 158 2319 162
rect 2323 158 2359 162
rect 2363 158 2407 162
rect 2411 158 2447 162
rect 1269 157 2447 158
rect 2453 157 2454 163
rect 1262 155 1270 157
rect 96 149 97 155
rect 103 154 1263 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 175 154
rect 179 150 215 154
rect 219 150 247 154
rect 251 150 255 154
rect 259 150 295 154
rect 299 150 327 154
rect 331 150 335 154
rect 339 150 375 154
rect 379 150 415 154
rect 419 150 423 154
rect 427 150 471 154
rect 475 150 495 154
rect 499 150 527 154
rect 531 150 575 154
rect 579 150 583 154
rect 587 150 631 154
rect 635 150 655 154
rect 659 150 679 154
rect 683 150 727 154
rect 731 150 767 154
rect 771 150 791 154
rect 795 150 807 154
rect 811 150 847 154
rect 851 150 887 154
rect 891 150 903 154
rect 907 150 927 154
rect 931 150 959 154
rect 963 150 975 154
rect 979 150 1023 154
rect 1027 150 1071 154
rect 1075 150 1111 154
rect 1115 150 1151 154
rect 1155 150 1191 154
rect 1195 150 1239 154
rect 1243 150 1263 154
rect 103 149 1263 150
rect 1269 149 1270 155
rect 1250 89 1251 95
rect 1257 94 2435 95
rect 1257 90 1279 94
rect 1283 90 1303 94
rect 1307 90 1343 94
rect 1347 90 1383 94
rect 1387 90 1423 94
rect 1427 90 1463 94
rect 1467 90 1519 94
rect 1523 90 1583 94
rect 1587 90 1647 94
rect 1651 90 1711 94
rect 1715 90 1767 94
rect 1771 90 1823 94
rect 1827 90 1871 94
rect 1875 90 1919 94
rect 1923 90 1967 94
rect 1971 90 2015 94
rect 2019 90 2063 94
rect 2067 90 2111 94
rect 2115 90 2159 94
rect 2163 90 2215 94
rect 2219 90 2271 94
rect 2275 90 2319 94
rect 2323 90 2359 94
rect 2363 90 2407 94
rect 2411 90 2435 94
rect 1257 89 2435 90
rect 2441 89 2442 95
rect 1250 87 1258 89
rect 84 81 85 87
rect 91 86 1251 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 175 86
rect 179 82 215 86
rect 219 82 255 86
rect 259 82 295 86
rect 299 82 335 86
rect 339 82 375 86
rect 379 82 423 86
rect 427 82 471 86
rect 475 82 527 86
rect 531 82 583 86
rect 587 82 631 86
rect 635 82 679 86
rect 683 82 727 86
rect 731 82 767 86
rect 771 82 807 86
rect 811 82 847 86
rect 851 82 887 86
rect 891 82 927 86
rect 931 82 975 86
rect 979 82 1023 86
rect 1027 82 1071 86
rect 1075 82 1111 86
rect 1115 82 1151 86
rect 1155 82 1191 86
rect 1195 82 1239 86
rect 1243 82 1251 86
rect 91 81 1251 82
rect 1257 81 1258 87
<< m5c >>
rect 1251 2509 1257 2515
rect 2435 2509 2441 2515
rect 97 2497 103 2503
rect 1263 2497 1269 2503
rect 1263 2441 1269 2447
rect 2447 2441 2453 2447
rect 85 2429 91 2435
rect 1251 2429 1257 2435
rect 1251 2373 1257 2379
rect 2435 2373 2441 2379
rect 97 2353 103 2359
rect 1263 2353 1269 2359
rect 1263 2301 1269 2307
rect 2447 2301 2453 2307
rect 85 2281 91 2287
rect 1251 2281 1257 2287
rect 1251 2225 1257 2231
rect 2435 2225 2441 2231
rect 97 2213 103 2219
rect 1263 2213 1269 2219
rect 1263 2157 1269 2163
rect 2447 2157 2453 2163
rect 85 2137 91 2143
rect 1251 2137 1257 2143
rect 1251 2085 1257 2091
rect 2435 2085 2441 2091
rect 97 2069 103 2075
rect 1263 2069 1269 2075
rect 1263 2009 1269 2015
rect 2447 2009 2453 2015
rect 85 1993 91 1999
rect 1251 1993 1257 1999
rect 1251 1941 1257 1947
rect 2435 1941 2441 1947
rect 97 1921 103 1927
rect 1263 1921 1269 1927
rect 1263 1873 1269 1879
rect 2447 1873 2453 1879
rect 85 1845 91 1851
rect 1251 1845 1257 1851
rect 1251 1801 1257 1807
rect 2435 1801 2441 1807
rect 97 1777 103 1783
rect 1263 1777 1269 1783
rect 1263 1733 1269 1739
rect 2447 1733 2453 1739
rect 85 1705 91 1711
rect 1251 1705 1257 1711
rect 1251 1665 1257 1671
rect 2435 1665 2441 1671
rect 97 1633 103 1639
rect 1263 1633 1269 1639
rect 1263 1597 1269 1603
rect 2447 1597 2453 1603
rect 85 1557 91 1563
rect 1251 1557 1257 1563
rect 1251 1525 1257 1531
rect 2435 1525 2441 1531
rect 1263 1457 1269 1463
rect 2447 1457 2453 1463
rect 97 1449 103 1455
rect 1263 1449 1269 1455
rect 85 1381 91 1387
rect 1251 1381 1257 1387
rect 97 1309 103 1315
rect 1263 1309 1269 1315
rect 85 1237 91 1243
rect 1251 1237 1257 1243
rect 97 1169 103 1175
rect 1263 1169 1269 1175
rect 85 1097 91 1103
rect 1251 1097 1257 1103
rect 97 1029 103 1035
rect 1263 1029 1269 1035
rect 85 961 91 967
rect 1251 961 1257 967
rect 97 885 103 891
rect 1263 885 1269 891
rect 85 817 91 823
rect 1251 817 1257 823
rect 1251 809 1257 815
rect 2435 809 2441 815
rect 97 745 103 751
rect 1263 745 1269 751
rect 85 673 91 679
rect 1251 673 1257 679
rect 97 597 103 603
rect 1263 597 1269 603
rect 1251 529 1257 535
rect 2435 529 2441 535
rect 85 521 91 527
rect 1251 521 1257 527
rect 97 453 103 459
rect 1263 453 1269 459
rect 85 385 91 391
rect 1251 385 1257 391
rect 97 313 103 319
rect 1263 313 1269 319
rect 85 237 91 243
rect 1251 237 1257 243
rect 1263 157 1269 163
rect 2447 157 2453 163
rect 97 149 103 155
rect 1263 149 1269 155
rect 1251 89 1257 95
rect 2435 89 2441 95
rect 85 81 91 87
rect 1251 81 1257 87
<< m5 >>
rect 84 2435 92 2520
rect 84 2429 85 2435
rect 91 2429 92 2435
rect 84 2287 92 2429
rect 84 2281 85 2287
rect 91 2281 92 2287
rect 84 2143 92 2281
rect 84 2137 85 2143
rect 91 2137 92 2143
rect 84 1999 92 2137
rect 84 1993 85 1999
rect 91 1993 92 1999
rect 84 1851 92 1993
rect 84 1845 85 1851
rect 91 1845 92 1851
rect 84 1711 92 1845
rect 84 1705 85 1711
rect 91 1705 92 1711
rect 84 1563 92 1705
rect 84 1557 85 1563
rect 91 1557 92 1563
rect 84 1387 92 1557
rect 84 1381 85 1387
rect 91 1381 92 1387
rect 84 1243 92 1381
rect 84 1237 85 1243
rect 91 1237 92 1243
rect 84 1103 92 1237
rect 84 1097 85 1103
rect 91 1097 92 1103
rect 84 967 92 1097
rect 84 961 85 967
rect 91 961 92 967
rect 84 823 92 961
rect 84 817 85 823
rect 91 817 92 823
rect 84 679 92 817
rect 84 673 85 679
rect 91 673 92 679
rect 84 527 92 673
rect 84 521 85 527
rect 91 521 92 527
rect 84 391 92 521
rect 84 385 85 391
rect 91 385 92 391
rect 84 243 92 385
rect 84 237 85 243
rect 91 237 92 243
rect 84 87 92 237
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2503 104 2520
rect 96 2497 97 2503
rect 103 2497 104 2503
rect 96 2359 104 2497
rect 96 2353 97 2359
rect 103 2353 104 2359
rect 96 2219 104 2353
rect 96 2213 97 2219
rect 103 2213 104 2219
rect 96 2075 104 2213
rect 96 2069 97 2075
rect 103 2069 104 2075
rect 96 1927 104 2069
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1783 104 1921
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1639 104 1777
rect 96 1633 97 1639
rect 103 1633 104 1639
rect 96 1455 104 1633
rect 96 1449 97 1455
rect 103 1449 104 1455
rect 96 1315 104 1449
rect 96 1309 97 1315
rect 103 1309 104 1315
rect 96 1175 104 1309
rect 96 1169 97 1175
rect 103 1169 104 1175
rect 96 1035 104 1169
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 891 104 1029
rect 96 885 97 891
rect 103 885 104 891
rect 96 751 104 885
rect 96 745 97 751
rect 103 745 104 751
rect 96 603 104 745
rect 96 597 97 603
rect 103 597 104 603
rect 96 459 104 597
rect 96 453 97 459
rect 103 453 104 459
rect 96 319 104 453
rect 96 313 97 319
rect 103 313 104 319
rect 96 155 104 313
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1250 2515 1258 2520
rect 1250 2509 1251 2515
rect 1257 2509 1258 2515
rect 1250 2435 1258 2509
rect 1250 2429 1251 2435
rect 1257 2429 1258 2435
rect 1250 2379 1258 2429
rect 1250 2373 1251 2379
rect 1257 2373 1258 2379
rect 1250 2287 1258 2373
rect 1250 2281 1251 2287
rect 1257 2281 1258 2287
rect 1250 2231 1258 2281
rect 1250 2225 1251 2231
rect 1257 2225 1258 2231
rect 1250 2143 1258 2225
rect 1250 2137 1251 2143
rect 1257 2137 1258 2143
rect 1250 2091 1258 2137
rect 1250 2085 1251 2091
rect 1257 2085 1258 2091
rect 1250 1999 1258 2085
rect 1250 1993 1251 1999
rect 1257 1993 1258 1999
rect 1250 1947 1258 1993
rect 1250 1941 1251 1947
rect 1257 1941 1258 1947
rect 1250 1851 1258 1941
rect 1250 1845 1251 1851
rect 1257 1845 1258 1851
rect 1250 1807 1258 1845
rect 1250 1801 1251 1807
rect 1257 1801 1258 1807
rect 1250 1711 1258 1801
rect 1250 1705 1251 1711
rect 1257 1705 1258 1711
rect 1250 1671 1258 1705
rect 1250 1665 1251 1671
rect 1257 1665 1258 1671
rect 1250 1563 1258 1665
rect 1250 1557 1251 1563
rect 1257 1557 1258 1563
rect 1250 1531 1258 1557
rect 1250 1525 1251 1531
rect 1257 1525 1258 1531
rect 1250 1387 1258 1525
rect 1250 1381 1251 1387
rect 1257 1381 1258 1387
rect 1250 1243 1258 1381
rect 1250 1237 1251 1243
rect 1257 1237 1258 1243
rect 1250 1103 1258 1237
rect 1250 1097 1251 1103
rect 1257 1097 1258 1103
rect 1250 967 1258 1097
rect 1250 961 1251 967
rect 1257 961 1258 967
rect 1250 823 1258 961
rect 1250 817 1251 823
rect 1257 817 1258 823
rect 1250 815 1258 817
rect 1250 809 1251 815
rect 1257 809 1258 815
rect 1250 679 1258 809
rect 1250 673 1251 679
rect 1257 673 1258 679
rect 1250 535 1258 673
rect 1250 529 1251 535
rect 1257 529 1258 535
rect 1250 527 1258 529
rect 1250 521 1251 527
rect 1257 521 1258 527
rect 1250 391 1258 521
rect 1250 385 1251 391
rect 1257 385 1258 391
rect 1250 243 1258 385
rect 1250 237 1251 243
rect 1257 237 1258 243
rect 1250 95 1258 237
rect 1250 89 1251 95
rect 1257 89 1258 95
rect 1250 87 1258 89
rect 1250 81 1251 87
rect 1257 81 1258 87
rect 1250 72 1258 81
rect 1262 2503 1270 2520
rect 1262 2497 1263 2503
rect 1269 2497 1270 2503
rect 1262 2447 1270 2497
rect 1262 2441 1263 2447
rect 1269 2441 1270 2447
rect 1262 2359 1270 2441
rect 1262 2353 1263 2359
rect 1269 2353 1270 2359
rect 1262 2307 1270 2353
rect 1262 2301 1263 2307
rect 1269 2301 1270 2307
rect 1262 2219 1270 2301
rect 1262 2213 1263 2219
rect 1269 2213 1270 2219
rect 1262 2163 1270 2213
rect 1262 2157 1263 2163
rect 1269 2157 1270 2163
rect 1262 2075 1270 2157
rect 1262 2069 1263 2075
rect 1269 2069 1270 2075
rect 1262 2015 1270 2069
rect 1262 2009 1263 2015
rect 1269 2009 1270 2015
rect 1262 1927 1270 2009
rect 1262 1921 1263 1927
rect 1269 1921 1270 1927
rect 1262 1879 1270 1921
rect 1262 1873 1263 1879
rect 1269 1873 1270 1879
rect 1262 1783 1270 1873
rect 1262 1777 1263 1783
rect 1269 1777 1270 1783
rect 1262 1739 1270 1777
rect 1262 1733 1263 1739
rect 1269 1733 1270 1739
rect 1262 1639 1270 1733
rect 1262 1633 1263 1639
rect 1269 1633 1270 1639
rect 1262 1603 1270 1633
rect 1262 1597 1263 1603
rect 1269 1597 1270 1603
rect 1262 1463 1270 1597
rect 1262 1457 1263 1463
rect 1269 1457 1270 1463
rect 1262 1455 1270 1457
rect 1262 1449 1263 1455
rect 1269 1449 1270 1455
rect 1262 1315 1270 1449
rect 1262 1309 1263 1315
rect 1269 1309 1270 1315
rect 1262 1175 1270 1309
rect 1262 1169 1263 1175
rect 1269 1169 1270 1175
rect 1262 1035 1270 1169
rect 1262 1029 1263 1035
rect 1269 1029 1270 1035
rect 1262 891 1270 1029
rect 1262 885 1263 891
rect 1269 885 1270 891
rect 1262 751 1270 885
rect 1262 745 1263 751
rect 1269 745 1270 751
rect 1262 603 1270 745
rect 1262 597 1263 603
rect 1269 597 1270 603
rect 1262 459 1270 597
rect 1262 453 1263 459
rect 1269 453 1270 459
rect 1262 319 1270 453
rect 1262 313 1263 319
rect 1269 313 1270 319
rect 1262 163 1270 313
rect 1262 157 1263 163
rect 1269 157 1270 163
rect 1262 155 1270 157
rect 1262 149 1263 155
rect 1269 149 1270 155
rect 1262 72 1270 149
rect 2434 2515 2442 2520
rect 2434 2509 2435 2515
rect 2441 2509 2442 2515
rect 2434 2379 2442 2509
rect 2434 2373 2435 2379
rect 2441 2373 2442 2379
rect 2434 2231 2442 2373
rect 2434 2225 2435 2231
rect 2441 2225 2442 2231
rect 2434 2091 2442 2225
rect 2434 2085 2435 2091
rect 2441 2085 2442 2091
rect 2434 1947 2442 2085
rect 2434 1941 2435 1947
rect 2441 1941 2442 1947
rect 2434 1807 2442 1941
rect 2434 1801 2435 1807
rect 2441 1801 2442 1807
rect 2434 1671 2442 1801
rect 2434 1665 2435 1671
rect 2441 1665 2442 1671
rect 2434 1531 2442 1665
rect 2434 1525 2435 1531
rect 2441 1525 2442 1531
rect 2434 815 2442 1525
rect 2434 809 2435 815
rect 2441 809 2442 815
rect 2434 535 2442 809
rect 2434 529 2435 535
rect 2441 529 2442 535
rect 2434 95 2442 529
rect 2434 89 2435 95
rect 2441 89 2442 95
rect 2434 72 2442 89
rect 2446 2447 2454 2520
rect 2446 2441 2447 2447
rect 2453 2441 2454 2447
rect 2446 2307 2454 2441
rect 2446 2301 2447 2307
rect 2453 2301 2454 2307
rect 2446 2163 2454 2301
rect 2446 2157 2447 2163
rect 2453 2157 2454 2163
rect 2446 2015 2454 2157
rect 2446 2009 2447 2015
rect 2453 2009 2454 2015
rect 2446 1879 2454 2009
rect 2446 1873 2447 1879
rect 2453 1873 2454 1879
rect 2446 1739 2454 1873
rect 2446 1733 2447 1739
rect 2453 1733 2454 1739
rect 2446 1603 2454 1733
rect 2446 1597 2447 1603
rect 2453 1597 2454 1603
rect 2446 1463 2454 1597
rect 2446 1457 2447 1463
rect 2453 1457 2454 1463
rect 2446 163 2454 1457
rect 2446 157 2447 163
rect 2453 157 2454 163
rect 2446 72 2454 157
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__133
timestamp 1731220636
transform 1 0 2400 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220636
transform 1 0 1272 0 -1 2504
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220636
transform 1 0 2400 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220636
transform 1 0 1272 0 1 2384
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220636
transform 1 0 2400 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220636
transform 1 0 1272 0 -1 2368
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220636
transform 1 0 2400 0 1 2244
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220636
transform 1 0 1272 0 1 2244
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220636
transform 1 0 2400 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220636
transform 1 0 1272 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220636
transform 1 0 2400 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220636
transform 1 0 1272 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220636
transform 1 0 2400 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220636
transform 1 0 1272 0 -1 2080
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220636
transform 1 0 2400 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220636
transform 1 0 1272 0 1 1952
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220636
transform 1 0 2400 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220636
transform 1 0 1272 0 -1 1936
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220636
transform 1 0 2400 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220636
transform 1 0 1272 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220636
transform 1 0 2400 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220636
transform 1 0 1272 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220636
transform 1 0 2400 0 1 1676
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220636
transform 1 0 1272 0 1 1676
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220636
transform 1 0 2400 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220636
transform 1 0 1272 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220636
transform 1 0 2400 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220636
transform 1 0 1272 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220636
transform 1 0 2400 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220636
transform 1 0 1272 0 -1 1520
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220636
transform 1 0 2400 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220636
transform 1 0 1272 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220636
transform 1 0 2400 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220636
transform 1 0 1272 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220636
transform 1 0 2400 0 1 1256
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220636
transform 1 0 1272 0 1 1256
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220636
transform 1 0 2400 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220636
transform 1 0 1272 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220636
transform 1 0 2400 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220636
transform 1 0 1272 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220636
transform 1 0 2400 0 -1 1096
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220636
transform 1 0 1272 0 -1 1096
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220636
transform 1 0 2400 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220636
transform 1 0 1272 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220636
transform 1 0 2400 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220636
transform 1 0 1272 0 -1 952
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220636
transform 1 0 2400 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220636
transform 1 0 1272 0 1 832
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220636
transform 1 0 2400 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220636
transform 1 0 1272 0 -1 804
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220636
transform 1 0 2400 0 1 684
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220636
transform 1 0 1272 0 1 684
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220636
transform 1 0 2400 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220636
transform 1 0 1272 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220636
transform 1 0 2400 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220636
transform 1 0 1272 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220636
transform 1 0 2400 0 -1 524
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220636
transform 1 0 1272 0 -1 524
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220636
transform 1 0 2400 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220636
transform 1 0 1272 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220636
transform 1 0 2400 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220636
transform 1 0 1272 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220636
transform 1 0 2400 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220636
transform 1 0 1272 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220636
transform 1 0 2400 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220636
transform 1 0 1272 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220636
transform 1 0 2400 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220636
transform 1 0 1272 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220636
transform 1 0 1232 0 1 2440
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220636
transform 1 0 104 0 1 2440
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220636
transform 1 0 1232 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220636
transform 1 0 104 0 -1 2424
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220636
transform 1 0 1232 0 1 2296
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220636
transform 1 0 104 0 1 2296
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220636
transform 1 0 1232 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220636
transform 1 0 104 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220636
transform 1 0 1232 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220636
transform 1 0 104 0 1 2156
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220636
transform 1 0 1232 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220636
transform 1 0 104 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220636
transform 1 0 1232 0 1 2012
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220636
transform 1 0 104 0 1 2012
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220636
transform 1 0 1232 0 -1 1988
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220636
transform 1 0 104 0 -1 1988
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220636
transform 1 0 1232 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220636
transform 1 0 104 0 1 1864
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220636
transform 1 0 1232 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220636
transform 1 0 104 0 -1 1840
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220636
transform 1 0 1232 0 1 1720
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220636
transform 1 0 104 0 1 1720
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220636
transform 1 0 1232 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220636
transform 1 0 104 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220636
transform 1 0 1232 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220636
transform 1 0 104 0 1 1576
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220636
transform 1 0 1232 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220636
transform 1 0 104 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220636
transform 1 0 1232 0 1 1392
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220636
transform 1 0 104 0 1 1392
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220636
transform 1 0 1232 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220636
transform 1 0 104 0 -1 1376
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220636
transform 1 0 1232 0 1 1252
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220636
transform 1 0 104 0 1 1252
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220636
transform 1 0 1232 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220636
transform 1 0 104 0 -1 1232
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220636
transform 1 0 1232 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220636
transform 1 0 104 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220636
transform 1 0 1232 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220636
transform 1 0 104 0 -1 1092
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220636
transform 1 0 1232 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220636
transform 1 0 104 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220636
transform 1 0 1232 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220636
transform 1 0 104 0 -1 956
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220636
transform 1 0 1232 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220636
transform 1 0 104 0 1 828
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220636
transform 1 0 1232 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220636
transform 1 0 104 0 -1 812
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220636
transform 1 0 1232 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220636
transform 1 0 104 0 1 688
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220636
transform 1 0 1232 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220636
transform 1 0 104 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220636
transform 1 0 1232 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220636
transform 1 0 104 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220636
transform 1 0 1232 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220636
transform 1 0 104 0 -1 516
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220636
transform 1 0 1232 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220636
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220636
transform 1 0 1232 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220636
transform 1 0 104 0 -1 380
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220636
transform 1 0 1232 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220636
transform 1 0 104 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220636
transform 1 0 1232 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220636
transform 1 0 104 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220636
transform 1 0 1232 0 1 92
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220636
transform 1 0 104 0 1 92
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X2  tst_5999_6
timestamp 1731220636
transform 1 0 2264 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5998_6
timestamp 1731220636
transform 1 0 2312 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5997_6
timestamp 1731220636
transform 1 0 2352 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5996_6
timestamp 1731220636
transform 1 0 2352 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5995_6
timestamp 1731220636
transform 1 0 2352 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5994_6
timestamp 1731220636
transform 1 0 2312 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5993_6
timestamp 1731220636
transform 1 0 2352 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5992_6
timestamp 1731220636
transform 1 0 2288 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5991_6
timestamp 1731220636
transform 1 0 2352 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5990_6
timestamp 1731220636
transform 1 0 2352 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5989_6
timestamp 1731220636
transform 1 0 2352 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5988_6
timestamp 1731220636
transform 1 0 2352 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5987_6
timestamp 1731220636
transform 1 0 2352 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5986_6
timestamp 1731220636
transform 1 0 2352 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5985_6
timestamp 1731220636
transform 1 0 2296 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5984_6
timestamp 1731220636
transform 1 0 2216 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5983_6
timestamp 1731220636
transform 1 0 2304 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5982_6
timestamp 1731220636
transform 1 0 2280 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5981_6
timestamp 1731220636
transform 1 0 2280 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5980_6
timestamp 1731220636
transform 1 0 2184 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5979_6
timestamp 1731220636
transform 1 0 2096 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5978_6
timestamp 1731220636
transform 1 0 2208 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5977_6
timestamp 1731220636
transform 1 0 2128 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5976_6
timestamp 1731220636
transform 1 0 2048 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5975_6
timestamp 1731220636
transform 1 0 2032 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5974_6
timestamp 1731220636
transform 1 0 1960 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5973_6
timestamp 1731220636
transform 1 0 2104 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5972_6
timestamp 1731220636
transform 1 0 2168 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5971_6
timestamp 1731220636
transform 1 0 2232 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5970_6
timestamp 1731220636
transform 1 0 2296 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5969_6
timestamp 1731220636
transform 1 0 2248 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5968_6
timestamp 1731220636
transform 1 0 2184 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5967_6
timestamp 1731220636
transform 1 0 2128 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5966_6
timestamp 1731220636
transform 1 0 2064 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5965_6
timestamp 1731220636
transform 1 0 2064 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5964_6
timestamp 1731220636
transform 1 0 2160 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5963_6
timestamp 1731220636
transform 1 0 2264 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5962_6
timestamp 1731220636
transform 1 0 2208 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5961_6
timestamp 1731220636
transform 1 0 2152 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5960_6
timestamp 1731220636
transform 1 0 2104 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5959_6
timestamp 1731220636
transform 1 0 2056 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5958_6
timestamp 1731220636
transform 1 0 2008 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5957_6
timestamp 1731220636
transform 1 0 1960 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5956_6
timestamp 1731220636
transform 1 0 1912 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5955_6
timestamp 1731220636
transform 1 0 1864 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5954_6
timestamp 1731220636
transform 1 0 1816 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5953_6
timestamp 1731220636
transform 1 0 1760 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5952_6
timestamp 1731220636
transform 1 0 1704 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5951_6
timestamp 1731220636
transform 1 0 1968 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5950_6
timestamp 1731220636
transform 1 0 1880 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5949_6
timestamp 1731220636
transform 1 0 1800 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5948_6
timestamp 1731220636
transform 1 0 1728 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5947_6
timestamp 1731220636
transform 1 0 2000 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5946_6
timestamp 1731220636
transform 1 0 1928 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5945_6
timestamp 1731220636
transform 1 0 1856 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5944_6
timestamp 1731220636
transform 1 0 1792 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5943_6
timestamp 1731220636
transform 1 0 1808 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5942_6
timestamp 1731220636
transform 1 0 1728 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5941_6
timestamp 1731220636
transform 1 0 1656 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5940_6
timestamp 1731220636
transform 1 0 1584 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5939_6
timestamp 1731220636
transform 1 0 1656 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5938_6
timestamp 1731220636
transform 1 0 1888 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5937_6
timestamp 1731220636
transform 1 0 1968 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5936_6
timestamp 1731220636
transform 1 0 1888 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5935_6
timestamp 1731220636
transform 1 0 1808 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5934_6
timestamp 1731220636
transform 1 0 1728 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5933_6
timestamp 1731220636
transform 1 0 1688 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5932_6
timestamp 1731220636
transform 1 0 1792 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5931_6
timestamp 1731220636
transform 1 0 2000 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5930_6
timestamp 1731220636
transform 1 0 1896 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5929_6
timestamp 1731220636
transform 1 0 1840 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5928_6
timestamp 1731220636
transform 1 0 1784 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5927_6
timestamp 1731220636
transform 1 0 1904 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5926_6
timestamp 1731220636
transform 1 0 1968 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5925_6
timestamp 1731220636
transform 1 0 2192 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5924_6
timestamp 1731220636
transform 1 0 2112 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5923_6
timestamp 1731220636
transform 1 0 2040 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5922_6
timestamp 1731220636
transform 1 0 1968 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5921_6
timestamp 1731220636
transform 1 0 1888 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5920_6
timestamp 1731220636
transform 1 0 1808 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5919_6
timestamp 1731220636
transform 1 0 2040 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5918_6
timestamp 1731220636
transform 1 0 2104 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5917_6
timestamp 1731220636
transform 1 0 2168 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5916_6
timestamp 1731220636
transform 1 0 2232 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5915_6
timestamp 1731220636
transform 1 0 2272 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5914_6
timestamp 1731220636
transform 1 0 2168 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5913_6
timestamp 1731220636
transform 1 0 2072 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5912_6
timestamp 1731220636
transform 1 0 1984 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5911_6
timestamp 1731220636
transform 1 0 1904 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5910_6
timestamp 1731220636
transform 1 0 1824 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5909_6
timestamp 1731220636
transform 1 0 2136 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5908_6
timestamp 1731220636
transform 1 0 2064 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5907_6
timestamp 1731220636
transform 1 0 1992 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5906_6
timestamp 1731220636
transform 1 0 1928 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5905_6
timestamp 1731220636
transform 1 0 1864 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5904_6
timestamp 1731220636
transform 1 0 1808 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5903_6
timestamp 1731220636
transform 1 0 1752 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5902_6
timestamp 1731220636
transform 1 0 1984 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5901_6
timestamp 1731220636
transform 1 0 1912 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5900_6
timestamp 1731220636
transform 1 0 1840 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5899_6
timestamp 1731220636
transform 1 0 1768 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5898_6
timestamp 1731220636
transform 1 0 1760 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5897_6
timestamp 1731220636
transform 1 0 1848 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5896_6
timestamp 1731220636
transform 1 0 1936 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5895_6
timestamp 1731220636
transform 1 0 2008 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5894_6
timestamp 1731220636
transform 1 0 1936 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5893_6
timestamp 1731220636
transform 1 0 1872 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5892_6
timestamp 1731220636
transform 1 0 1816 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5891_6
timestamp 1731220636
transform 1 0 1768 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5890_6
timestamp 1731220636
transform 1 0 1816 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5889_6
timestamp 1731220636
transform 1 0 1864 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5888_6
timestamp 1731220636
transform 1 0 1912 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5887_6
timestamp 1731220636
transform 1 0 1960 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5886_6
timestamp 1731220636
transform 1 0 2008 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5885_6
timestamp 1731220636
transform 1 0 2056 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5884_6
timestamp 1731220636
transform 1 0 2112 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5883_6
timestamp 1731220636
transform 1 0 2088 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5882_6
timestamp 1731220636
transform 1 0 2096 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5881_6
timestamp 1731220636
transform 1 0 2016 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5880_6
timestamp 1731220636
transform 1 0 2056 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5879_6
timestamp 1731220636
transform 1 0 2128 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5878_6
timestamp 1731220636
transform 1 0 2208 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5877_6
timestamp 1731220636
transform 1 0 2288 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5876_6
timestamp 1731220636
transform 1 0 2264 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5875_6
timestamp 1731220636
transform 1 0 2176 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5874_6
timestamp 1731220636
transform 1 0 2168 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5873_6
timestamp 1731220636
transform 1 0 2248 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5872_6
timestamp 1731220636
transform 1 0 2224 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5871_6
timestamp 1731220636
transform 1 0 2168 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5870_6
timestamp 1731220636
transform 1 0 2072 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5869_6
timestamp 1731220636
transform 1 0 1992 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5868_6
timestamp 1731220636
transform 1 0 1896 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5867_6
timestamp 1731220636
transform 1 0 2144 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5866_6
timestamp 1731220636
transform 1 0 2064 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5865_6
timestamp 1731220636
transform 1 0 1976 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5864_6
timestamp 1731220636
transform 1 0 1880 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5863_6
timestamp 1731220636
transform 1 0 1784 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5862_6
timestamp 1731220636
transform 1 0 2192 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5861_6
timestamp 1731220636
transform 1 0 2112 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5860_6
timestamp 1731220636
transform 1 0 2032 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5859_6
timestamp 1731220636
transform 1 0 1960 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5858_6
timestamp 1731220636
transform 1 0 1896 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5857_6
timestamp 1731220636
transform 1 0 1840 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5856_6
timestamp 1731220636
transform 1 0 1784 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5855_6
timestamp 1731220636
transform 1 0 1760 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5854_6
timestamp 1731220636
transform 1 0 1840 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5853_6
timestamp 1731220636
transform 1 0 1928 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5852_6
timestamp 1731220636
transform 1 0 2104 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5851_6
timestamp 1731220636
transform 1 0 2016 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5850_6
timestamp 1731220636
transform 1 0 1936 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5849_6
timestamp 1731220636
transform 1 0 1872 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5848_6
timestamp 1731220636
transform 1 0 1800 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5847_6
timestamp 1731220636
transform 1 0 1992 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5846_6
timestamp 1731220636
transform 1 0 2040 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5845_6
timestamp 1731220636
transform 1 0 2088 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5844_6
timestamp 1731220636
transform 1 0 2136 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5843_6
timestamp 1731220636
transform 1 0 2184 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5842_6
timestamp 1731220636
transform 1 0 2232 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5841_6
timestamp 1731220636
transform 1 0 2272 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5840_6
timestamp 1731220636
transform 1 0 2312 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5839_6
timestamp 1731220636
transform 1 0 2280 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5838_6
timestamp 1731220636
transform 1 0 2192 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5837_6
timestamp 1731220636
transform 1 0 2280 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5836_6
timestamp 1731220636
transform 1 0 2216 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5835_6
timestamp 1731220636
transform 1 0 2152 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5834_6
timestamp 1731220636
transform 1 0 2224 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5833_6
timestamp 1731220636
transform 1 0 2296 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5832_6
timestamp 1731220636
transform 1 0 2352 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5831_6
timestamp 1731220636
transform 1 0 2296 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5830_6
timestamp 1731220636
transform 1 0 2352 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5829_6
timestamp 1731220636
transform 1 0 2352 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5828_6
timestamp 1731220636
transform 1 0 2352 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5827_6
timestamp 1731220636
transform 1 0 2352 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5826_6
timestamp 1731220636
transform 1 0 2352 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5825_6
timestamp 1731220636
transform 1 0 2208 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5824_6
timestamp 1731220636
transform 1 0 2352 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5823_6
timestamp 1731220636
transform 1 0 2312 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5822_6
timestamp 1731220636
transform 1 0 2264 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5821_6
timestamp 1731220636
transform 1 0 2208 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5820_6
timestamp 1731220636
transform 1 0 2160 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5819_6
timestamp 1731220636
transform 1 0 2104 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5818_6
timestamp 1731220636
transform 1 0 2040 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5817_6
timestamp 1731220636
transform 1 0 1976 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5816_6
timestamp 1731220636
transform 1 0 1904 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5815_6
timestamp 1731220636
transform 1 0 2216 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5814_6
timestamp 1731220636
transform 1 0 2152 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5813_6
timestamp 1731220636
transform 1 0 2088 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5812_6
timestamp 1731220636
transform 1 0 2024 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5811_6
timestamp 1731220636
transform 1 0 1960 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5810_6
timestamp 1731220636
transform 1 0 1888 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5809_6
timestamp 1731220636
transform 1 0 1808 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5808_6
timestamp 1731220636
transform 1 0 2056 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5807_6
timestamp 1731220636
transform 1 0 1992 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5806_6
timestamp 1731220636
transform 1 0 1928 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5805_6
timestamp 1731220636
transform 1 0 1864 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5804_6
timestamp 1731220636
transform 1 0 1800 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5803_6
timestamp 1731220636
transform 1 0 1728 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5802_6
timestamp 1731220636
transform 1 0 1952 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5801_6
timestamp 1731220636
transform 1 0 1888 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5800_6
timestamp 1731220636
transform 1 0 1832 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5799_6
timestamp 1731220636
transform 1 0 1776 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5798_6
timestamp 1731220636
transform 1 0 1720 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5797_6
timestamp 1731220636
transform 1 0 1656 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5796_6
timestamp 1731220636
transform 1 0 1680 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5795_6
timestamp 1731220636
transform 1 0 1760 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5794_6
timestamp 1731220636
transform 1 0 1856 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5793_6
timestamp 1731220636
transform 1 0 2216 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5792_6
timestamp 1731220636
transform 1 0 2088 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5791_6
timestamp 1731220636
transform 1 0 1968 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5790_6
timestamp 1731220636
transform 1 0 1928 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5789_6
timestamp 1731220636
transform 1 0 1856 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5788_6
timestamp 1731220636
transform 1 0 1784 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5787_6
timestamp 1731220636
transform 1 0 2000 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5786_6
timestamp 1731220636
transform 1 0 2144 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5785_6
timestamp 1731220636
transform 1 0 2072 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5784_6
timestamp 1731220636
transform 1 0 1992 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5783_6
timestamp 1731220636
transform 1 0 1912 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5782_6
timestamp 1731220636
transform 1 0 2064 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5781_6
timestamp 1731220636
transform 1 0 2128 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5780_6
timestamp 1731220636
transform 1 0 2184 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5779_6
timestamp 1731220636
transform 1 0 2160 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5778_6
timestamp 1731220636
transform 1 0 2088 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5777_6
timestamp 1731220636
transform 1 0 2232 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5776_6
timestamp 1731220636
transform 1 0 2304 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5775_6
timestamp 1731220636
transform 1 0 2312 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5774_6
timestamp 1731220636
transform 1 0 2352 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5773_6
timestamp 1731220636
transform 1 0 2352 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5772_6
timestamp 1731220636
transform 1 0 2352 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5771_6
timestamp 1731220636
transform 1 0 2296 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5770_6
timestamp 1731220636
transform 1 0 2216 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5769_6
timestamp 1731220636
transform 1 0 2248 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5768_6
timestamp 1731220636
transform 1 0 2352 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5767_6
timestamp 1731220636
transform 1 0 2352 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5766_6
timestamp 1731220636
transform 1 0 2304 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5765_6
timestamp 1731220636
transform 1 0 2352 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5764_6
timestamp 1731220636
transform 1 0 2352 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5763_6
timestamp 1731220636
transform 1 0 2288 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5762_6
timestamp 1731220636
transform 1 0 2296 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5761_6
timestamp 1731220636
transform 1 0 2352 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5760_6
timestamp 1731220636
transform 1 0 2328 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5759_6
timestamp 1731220636
transform 1 0 2216 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5758_6
timestamp 1731220636
transform 1 0 2200 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5757_6
timestamp 1731220636
transform 1 0 2120 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5756_6
timestamp 1731220636
transform 1 0 2176 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5755_6
timestamp 1731220636
transform 1 0 2272 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5754_6
timestamp 1731220636
transform 1 0 2232 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5753_6
timestamp 1731220636
transform 1 0 2168 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5752_6
timestamp 1731220636
transform 1 0 2104 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5751_6
timestamp 1731220636
transform 1 0 2008 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5750_6
timestamp 1731220636
transform 1 0 1928 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5749_6
timestamp 1731220636
transform 1 0 2040 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5748_6
timestamp 1731220636
transform 1 0 1968 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5747_6
timestamp 1731220636
transform 1 0 1888 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5746_6
timestamp 1731220636
transform 1 0 1808 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5745_6
timestamp 1731220636
transform 1 0 2088 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5744_6
timestamp 1731220636
transform 1 0 2008 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5743_6
timestamp 1731220636
transform 1 0 1928 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5742_6
timestamp 1731220636
transform 1 0 1848 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5741_6
timestamp 1731220636
transform 1 0 1776 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5740_6
timestamp 1731220636
transform 1 0 2040 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5739_6
timestamp 1731220636
transform 1 0 1960 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5738_6
timestamp 1731220636
transform 1 0 1888 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5737_6
timestamp 1731220636
transform 1 0 1816 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5736_6
timestamp 1731220636
transform 1 0 1752 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5735_6
timestamp 1731220636
transform 1 0 1768 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5734_6
timestamp 1731220636
transform 1 0 1848 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5733_6
timestamp 1731220636
transform 1 0 1920 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5732_6
timestamp 1731220636
transform 1 0 1992 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5731_6
timestamp 1731220636
transform 1 0 2064 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5730_6
timestamp 1731220636
transform 1 0 2136 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5729_6
timestamp 1731220636
transform 1 0 2240 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5728_6
timestamp 1731220636
transform 1 0 2152 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5727_6
timestamp 1731220636
transform 1 0 2072 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5726_6
timestamp 1731220636
transform 1 0 1992 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5725_6
timestamp 1731220636
transform 1 0 1912 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5724_6
timestamp 1731220636
transform 1 0 1832 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5723_6
timestamp 1731220636
transform 1 0 1968 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5722_6
timestamp 1731220636
transform 1 0 1928 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5721_6
timestamp 1731220636
transform 1 0 1888 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5720_6
timestamp 1731220636
transform 1 0 1848 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5719_6
timestamp 1731220636
transform 1 0 1808 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5718_6
timestamp 1731220636
transform 1 0 1768 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5717_6
timestamp 1731220636
transform 1 0 1728 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5716_6
timestamp 1731220636
transform 1 0 1688 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5715_6
timestamp 1731220636
transform 1 0 1648 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5714_6
timestamp 1731220636
transform 1 0 1608 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5713_6
timestamp 1731220636
transform 1 0 1568 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5712_6
timestamp 1731220636
transform 1 0 1528 0 -1 2512
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5711_6
timestamp 1731220636
transform 1 0 1752 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5710_6
timestamp 1731220636
transform 1 0 1672 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5709_6
timestamp 1731220636
transform 1 0 1592 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5708_6
timestamp 1731220636
transform 1 0 1512 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5707_6
timestamp 1731220636
transform 1 0 1448 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5706_6
timestamp 1731220636
transform 1 0 1392 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5705_6
timestamp 1731220636
transform 1 0 1352 0 1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5704_6
timestamp 1731220636
transform 1 0 1352 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5703_6
timestamp 1731220636
transform 1 0 1400 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5702_6
timestamp 1731220636
transform 1 0 1464 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5701_6
timestamp 1731220636
transform 1 0 1536 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5700_6
timestamp 1731220636
transform 1 0 1688 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5699_6
timestamp 1731220636
transform 1 0 1608 0 -1 2376
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5698_6
timestamp 1731220636
transform 1 0 1576 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5697_6
timestamp 1731220636
transform 1 0 1536 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5696_6
timestamp 1731220636
transform 1 0 1496 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5695_6
timestamp 1731220636
transform 1 0 1616 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5694_6
timestamp 1731220636
transform 1 0 1696 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5693_6
timestamp 1731220636
transform 1 0 1656 0 1 2236
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5692_6
timestamp 1731220636
transform 1 0 1632 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5691_6
timestamp 1731220636
transform 1 0 1704 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5690_6
timestamp 1731220636
transform 1 0 1720 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5689_6
timestamp 1731220636
transform 1 0 1752 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5688_6
timestamp 1731220636
transform 1 0 1840 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5687_6
timestamp 1731220636
transform 1 0 1832 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5686_6
timestamp 1731220636
transform 1 0 1744 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5685_6
timestamp 1731220636
transform 1 0 1656 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5684_6
timestamp 1731220636
transform 1 0 1704 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5683_6
timestamp 1731220636
transform 1 0 1616 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5682_6
timestamp 1731220636
transform 1 0 1528 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5681_6
timestamp 1731220636
transform 1 0 1488 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5680_6
timestamp 1731220636
transform 1 0 1416 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5679_6
timestamp 1731220636
transform 1 0 1568 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5678_6
timestamp 1731220636
transform 1 0 1656 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5677_6
timestamp 1731220636
transform 1 0 1560 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5676_6
timestamp 1731220636
transform 1 0 1472 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5675_6
timestamp 1731220636
transform 1 0 1392 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5674_6
timestamp 1731220636
transform 1 0 1432 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5673_6
timestamp 1731220636
transform 1 0 1528 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5672_6
timestamp 1731220636
transform 1 0 1624 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5671_6
timestamp 1731220636
transform 1 0 1560 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5670_6
timestamp 1731220636
transform 1 0 1488 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5669_6
timestamp 1731220636
transform 1 0 1424 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5668_6
timestamp 1731220636
transform 1 0 1376 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5667_6
timestamp 1731220636
transform 1 0 1336 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5666_6
timestamp 1731220636
transform 1 0 1296 0 -1 2228
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5665_6
timestamp 1731220636
transform 1 0 1344 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5664_6
timestamp 1731220636
transform 1 0 1296 0 1 2092
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5663_6
timestamp 1731220636
transform 1 0 1296 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5662_6
timestamp 1731220636
transform 1 0 1336 0 -1 2088
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5661_6
timestamp 1731220636
transform 1 0 1344 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5660_6
timestamp 1731220636
transform 1 0 1296 0 1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5659_6
timestamp 1731220636
transform 1 0 1296 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5658_6
timestamp 1731220636
transform 1 0 1352 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5657_6
timestamp 1731220636
transform 1 0 1440 0 -1 1944
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5656_6
timestamp 1731220636
transform 1 0 1408 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5655_6
timestamp 1731220636
transform 1 0 1352 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5654_6
timestamp 1731220636
transform 1 0 1304 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5653_6
timestamp 1731220636
transform 1 0 1472 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5652_6
timestamp 1731220636
transform 1 0 1536 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5651_6
timestamp 1731220636
transform 1 0 1608 0 1 1808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5650_6
timestamp 1731220636
transform 1 0 1592 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5649_6
timestamp 1731220636
transform 1 0 1528 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5648_6
timestamp 1731220636
transform 1 0 1464 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5647_6
timestamp 1731220636
transform 1 0 1400 0 -1 1804
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5646_6
timestamp 1731220636
transform 1 0 1416 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5645_6
timestamp 1731220636
transform 1 0 1496 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5644_6
timestamp 1731220636
transform 1 0 1576 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5643_6
timestamp 1731220636
transform 1 0 1656 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5642_6
timestamp 1731220636
transform 1 0 1720 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5641_6
timestamp 1731220636
transform 1 0 1632 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5640_6
timestamp 1731220636
transform 1 0 1536 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5639_6
timestamp 1731220636
transform 1 0 1472 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5638_6
timestamp 1731220636
transform 1 0 1560 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5637_6
timestamp 1731220636
transform 1 0 1648 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5636_6
timestamp 1731220636
transform 1 0 1736 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5635_6
timestamp 1731220636
transform 1 0 1824 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5634_6
timestamp 1731220636
transform 1 0 2040 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5633_6
timestamp 1731220636
transform 1 0 1880 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5632_6
timestamp 1731220636
transform 1 0 1736 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5631_6
timestamp 1731220636
transform 1 0 1608 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5630_6
timestamp 1731220636
transform 1 0 1720 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5629_6
timestamp 1731220636
transform 1 0 1632 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5628_6
timestamp 1731220636
transform 1 0 1544 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5627_6
timestamp 1731220636
transform 1 0 1528 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5626_6
timestamp 1731220636
transform 1 0 1600 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5625_6
timestamp 1731220636
transform 1 0 1680 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5624_6
timestamp 1731220636
transform 1 0 1728 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5623_6
timestamp 1731220636
transform 1 0 1672 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5622_6
timestamp 1731220636
transform 1 0 1616 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5621_6
timestamp 1731220636
transform 1 0 1576 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5620_6
timestamp 1731220636
transform 1 0 1456 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5619_6
timestamp 1731220636
transform 1 0 1416 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5618_6
timestamp 1731220636
transform 1 0 1376 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5617_6
timestamp 1731220636
transform 1 0 1336 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5616_6
timestamp 1731220636
transform 1 0 1296 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5615_6
timestamp 1731220636
transform 1 0 1296 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5614_6
timestamp 1731220636
transform 1 0 1184 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5613_6
timestamp 1731220636
transform 1 0 1136 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5612_6
timestamp 1731220636
transform 1 0 1072 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5611_6
timestamp 1731220636
transform 1 0 1184 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5610_6
timestamp 1731220636
transform 1 0 1144 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5609_6
timestamp 1731220636
transform 1 0 1096 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5608_6
timestamp 1731220636
transform 1 0 1040 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5607_6
timestamp 1731220636
transform 1 0 992 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5606_6
timestamp 1731220636
transform 1 0 936 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5605_6
timestamp 1731220636
transform 1 0 872 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5604_6
timestamp 1731220636
transform 1 0 800 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5603_6
timestamp 1731220636
transform 1 0 720 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5602_6
timestamp 1731220636
transform 1 0 1008 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5601_6
timestamp 1731220636
transform 1 0 944 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5600_6
timestamp 1731220636
transform 1 0 880 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5599_6
timestamp 1731220636
transform 1 0 816 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5598_6
timestamp 1731220636
transform 1 0 744 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5597_6
timestamp 1731220636
transform 1 0 672 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5596_6
timestamp 1731220636
transform 1 0 992 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5595_6
timestamp 1731220636
transform 1 0 928 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5594_6
timestamp 1731220636
transform 1 0 872 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5593_6
timestamp 1731220636
transform 1 0 816 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5592_6
timestamp 1731220636
transform 1 0 760 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5591_6
timestamp 1731220636
transform 1 0 696 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5590_6
timestamp 1731220636
transform 1 0 632 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5589_6
timestamp 1731220636
transform 1 0 656 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5588_6
timestamp 1731220636
transform 1 0 736 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5587_6
timestamp 1731220636
transform 1 0 808 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5586_6
timestamp 1731220636
transform 1 0 872 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5585_6
timestamp 1731220636
transform 1 0 936 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5584_6
timestamp 1731220636
transform 1 0 1000 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5583_6
timestamp 1731220636
transform 1 0 1064 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5582_6
timestamp 1731220636
transform 1 0 1184 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5581_6
timestamp 1731220636
transform 1 0 1136 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5580_6
timestamp 1731220636
transform 1 0 1064 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5579_6
timestamp 1731220636
transform 1 0 992 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5578_6
timestamp 1731220636
transform 1 0 912 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5577_6
timestamp 1731220636
transform 1 0 832 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5576_6
timestamp 1731220636
transform 1 0 736 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5575_6
timestamp 1731220636
transform 1 0 1040 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5574_6
timestamp 1731220636
transform 1 0 976 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5573_6
timestamp 1731220636
transform 1 0 912 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5572_6
timestamp 1731220636
transform 1 0 856 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5571_6
timestamp 1731220636
transform 1 0 792 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5570_6
timestamp 1731220636
transform 1 0 728 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5569_6
timestamp 1731220636
transform 1 0 656 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5568_6
timestamp 1731220636
transform 1 0 1096 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5567_6
timestamp 1731220636
transform 1 0 992 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5566_6
timestamp 1731220636
transform 1 0 888 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5565_6
timestamp 1731220636
transform 1 0 800 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5564_6
timestamp 1731220636
transform 1 0 728 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5563_6
timestamp 1731220636
transform 1 0 664 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5562_6
timestamp 1731220636
transform 1 0 616 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5561_6
timestamp 1731220636
transform 1 0 848 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5560_6
timestamp 1731220636
transform 1 0 776 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5559_6
timestamp 1731220636
transform 1 0 704 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5558_6
timestamp 1731220636
transform 1 0 632 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5557_6
timestamp 1731220636
transform 1 0 568 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5556_6
timestamp 1731220636
transform 1 0 512 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5555_6
timestamp 1731220636
transform 1 0 456 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5554_6
timestamp 1731220636
transform 1 0 568 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5553_6
timestamp 1731220636
transform 1 0 512 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5552_6
timestamp 1731220636
transform 1 0 456 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5551_6
timestamp 1731220636
transform 1 0 392 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5550_6
timestamp 1731220636
transform 1 0 320 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5549_6
timestamp 1731220636
transform 1 0 576 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5548_6
timestamp 1731220636
transform 1 0 496 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5547_6
timestamp 1731220636
transform 1 0 408 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5546_6
timestamp 1731220636
transform 1 0 320 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5545_6
timestamp 1731220636
transform 1 0 632 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5544_6
timestamp 1731220636
transform 1 0 528 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5543_6
timestamp 1731220636
transform 1 0 424 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5542_6
timestamp 1731220636
transform 1 0 320 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5541_6
timestamp 1731220636
transform 1 0 232 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5540_6
timestamp 1731220636
transform 1 0 304 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5539_6
timestamp 1731220636
transform 1 0 392 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5538_6
timestamp 1731220636
transform 1 0 480 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5537_6
timestamp 1731220636
transform 1 0 568 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5536_6
timestamp 1731220636
transform 1 0 560 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5535_6
timestamp 1731220636
transform 1 0 488 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5534_6
timestamp 1731220636
transform 1 0 416 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5533_6
timestamp 1731220636
transform 1 0 344 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5532_6
timestamp 1731220636
transform 1 0 280 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5531_6
timestamp 1731220636
transform 1 0 592 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5530_6
timestamp 1731220636
transform 1 0 512 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5529_6
timestamp 1731220636
transform 1 0 432 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5528_6
timestamp 1731220636
transform 1 0 360 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5527_6
timestamp 1731220636
transform 1 0 640 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5526_6
timestamp 1731220636
transform 1 0 552 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5525_6
timestamp 1731220636
transform 1 0 464 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5524_6
timestamp 1731220636
transform 1 0 384 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5523_6
timestamp 1731220636
transform 1 0 312 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5522_6
timestamp 1731220636
transform 1 0 256 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5521_6
timestamp 1731220636
transform 1 0 216 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5520_6
timestamp 1731220636
transform 1 0 176 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5519_6
timestamp 1731220636
transform 1 0 136 0 1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5518_6
timestamp 1731220636
transform 1 0 296 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5517_6
timestamp 1731220636
transform 1 0 240 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5516_6
timestamp 1731220636
transform 1 0 200 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5515_6
timestamp 1731220636
transform 1 0 160 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5514_6
timestamp 1731220636
transform 1 0 176 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5513_6
timestamp 1731220636
transform 1 0 224 0 1 1244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5512_6
timestamp 1731220636
transform 1 0 224 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5511_6
timestamp 1731220636
transform 1 0 168 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5510_6
timestamp 1731220636
transform 1 0 128 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5509_6
timestamp 1731220636
transform 1 0 128 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5508_6
timestamp 1731220636
transform 1 0 168 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5507_6
timestamp 1731220636
transform 1 0 128 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5506_6
timestamp 1731220636
transform 1 0 240 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5505_6
timestamp 1731220636
transform 1 0 168 0 -1 1100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5504_6
timestamp 1731220636
transform 1 0 168 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5503_6
timestamp 1731220636
transform 1 0 248 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5502_6
timestamp 1731220636
transform 1 0 248 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5501_6
timestamp 1731220636
transform 1 0 208 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5500_6
timestamp 1731220636
transform 1 0 296 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5499_6
timestamp 1731220636
transform 1 0 352 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5498_6
timestamp 1731220636
transform 1 0 408 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5497_6
timestamp 1731220636
transform 1 0 632 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5496_6
timestamp 1731220636
transform 1 0 536 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5495_6
timestamp 1731220636
transform 1 0 440 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5494_6
timestamp 1731220636
transform 1 0 352 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5493_6
timestamp 1731220636
transform 1 0 280 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5492_6
timestamp 1731220636
transform 1 0 224 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5491_6
timestamp 1731220636
transform 1 0 184 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5490_6
timestamp 1731220636
transform 1 0 496 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5489_6
timestamp 1731220636
transform 1 0 408 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5488_6
timestamp 1731220636
transform 1 0 320 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5487_6
timestamp 1731220636
transform 1 0 232 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5486_6
timestamp 1731220636
transform 1 0 168 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5485_6
timestamp 1731220636
transform 1 0 128 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5484_6
timestamp 1731220636
transform 1 0 128 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5483_6
timestamp 1731220636
transform 1 0 184 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5482_6
timestamp 1731220636
transform 1 0 192 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5481_6
timestamp 1731220636
transform 1 0 128 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5480_6
timestamp 1731220636
transform 1 0 128 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5479_6
timestamp 1731220636
transform 1 0 184 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5478_6
timestamp 1731220636
transform 1 0 264 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5477_6
timestamp 1731220636
transform 1 0 256 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5476_6
timestamp 1731220636
transform 1 0 184 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5475_6
timestamp 1731220636
transform 1 0 128 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5474_6
timestamp 1731220636
transform 1 0 176 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5473_6
timestamp 1731220636
transform 1 0 216 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5472_6
timestamp 1731220636
transform 1 0 256 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5471_6
timestamp 1731220636
transform 1 0 280 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5470_6
timestamp 1731220636
transform 1 0 224 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5469_6
timestamp 1731220636
transform 1 0 168 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5468_6
timestamp 1731220636
transform 1 0 128 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5467_6
timestamp 1731220636
transform 1 0 248 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5466_6
timestamp 1731220636
transform 1 0 176 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5465_6
timestamp 1731220636
transform 1 0 128 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5464_6
timestamp 1731220636
transform 1 0 128 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5463_6
timestamp 1731220636
transform 1 0 168 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5462_6
timestamp 1731220636
transform 1 0 320 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5461_6
timestamp 1731220636
transform 1 0 240 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5460_6
timestamp 1731220636
transform 1 0 208 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5459_6
timestamp 1731220636
transform 1 0 168 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5458_6
timestamp 1731220636
transform 1 0 128 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5457_6
timestamp 1731220636
transform 1 0 248 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5456_6
timestamp 1731220636
transform 1 0 288 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5455_6
timestamp 1731220636
transform 1 0 328 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5454_6
timestamp 1731220636
transform 1 0 368 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5453_6
timestamp 1731220636
transform 1 0 416 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5452_6
timestamp 1731220636
transform 1 0 464 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5451_6
timestamp 1731220636
transform 1 0 576 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5450_6
timestamp 1731220636
transform 1 0 520 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5449_6
timestamp 1731220636
transform 1 0 488 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5448_6
timestamp 1731220636
transform 1 0 408 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5447_6
timestamp 1731220636
transform 1 0 568 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5446_6
timestamp 1731220636
transform 1 0 544 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5445_6
timestamp 1731220636
transform 1 0 496 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5444_6
timestamp 1731220636
transform 1 0 440 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5443_6
timestamp 1731220636
transform 1 0 384 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5442_6
timestamp 1731220636
transform 1 0 320 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5441_6
timestamp 1731220636
transform 1 0 336 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5440_6
timestamp 1731220636
transform 1 0 384 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5439_6
timestamp 1731220636
transform 1 0 432 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5438_6
timestamp 1731220636
transform 1 0 488 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5437_6
timestamp 1731220636
transform 1 0 424 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5436_6
timestamp 1731220636
transform 1 0 360 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5435_6
timestamp 1731220636
transform 1 0 304 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5434_6
timestamp 1731220636
transform 1 0 328 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5433_6
timestamp 1731220636
transform 1 0 408 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5432_6
timestamp 1731220636
transform 1 0 488 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5431_6
timestamp 1731220636
transform 1 0 568 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5430_6
timestamp 1731220636
transform 1 0 528 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5429_6
timestamp 1731220636
transform 1 0 440 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5428_6
timestamp 1731220636
transform 1 0 352 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5427_6
timestamp 1731220636
transform 1 0 696 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5426_6
timestamp 1731220636
transform 1 0 616 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5425_6
timestamp 1731220636
transform 1 0 552 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5424_6
timestamp 1731220636
transform 1 0 480 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5423_6
timestamp 1731220636
transform 1 0 408 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5422_6
timestamp 1731220636
transform 1 0 344 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5421_6
timestamp 1731220636
transform 1 0 272 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5420_6
timestamp 1731220636
transform 1 0 256 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5419_6
timestamp 1731220636
transform 1 0 328 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5418_6
timestamp 1731220636
transform 1 0 392 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5417_6
timestamp 1731220636
transform 1 0 448 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5416_6
timestamp 1731220636
transform 1 0 496 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5415_6
timestamp 1731220636
transform 1 0 536 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5414_6
timestamp 1731220636
transform 1 0 576 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5413_6
timestamp 1731220636
transform 1 0 616 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5412_6
timestamp 1731220636
transform 1 0 632 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5411_6
timestamp 1731220636
transform 1 0 704 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5410_6
timestamp 1731220636
transform 1 0 776 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5409_6
timestamp 1731220636
transform 1 0 760 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5408_6
timestamp 1731220636
transform 1 0 712 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5407_6
timestamp 1731220636
transform 1 0 664 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5406_6
timestamp 1731220636
transform 1 0 904 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5405_6
timestamp 1731220636
transform 1 0 856 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5404_6
timestamp 1731220636
transform 1 0 808 0 1 680
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5403_6
timestamp 1731220636
transform 1 0 736 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5402_6
timestamp 1731220636
transform 1 0 664 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5401_6
timestamp 1731220636
transform 1 0 584 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5400_6
timestamp 1731220636
transform 1 0 808 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5399_6
timestamp 1731220636
transform 1 0 1008 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5398_6
timestamp 1731220636
transform 1 0 936 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5397_6
timestamp 1731220636
transform 1 0 872 0 -1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5396_6
timestamp 1731220636
transform 1 0 800 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5395_6
timestamp 1731220636
transform 1 0 720 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5394_6
timestamp 1731220636
transform 1 0 880 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5393_6
timestamp 1731220636
transform 1 0 952 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5392_6
timestamp 1731220636
transform 1 0 1152 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5391_6
timestamp 1731220636
transform 1 0 1080 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5390_6
timestamp 1731220636
transform 1 0 1016 0 1 820
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5389_6
timestamp 1731220636
transform 1 0 992 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5388_6
timestamp 1731220636
transform 1 0 920 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5387_6
timestamp 1731220636
transform 1 0 1064 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5386_6
timestamp 1731220636
transform 1 0 1136 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5385_6
timestamp 1731220636
transform 1 0 1184 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5384_6
timestamp 1731220636
transform 1 0 1184 0 -1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5383_6
timestamp 1731220636
transform 1 0 1296 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5382_6
timestamp 1731220636
transform 1 0 1344 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5381_6
timestamp 1731220636
transform 1 0 1424 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5380_6
timestamp 1731220636
transform 1 0 1504 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5379_6
timestamp 1731220636
transform 1 0 1600 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5378_6
timestamp 1731220636
transform 1 0 1552 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5377_6
timestamp 1731220636
transform 1 0 1512 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5376_6
timestamp 1731220636
transform 1 0 1472 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5375_6
timestamp 1731220636
transform 1 0 1432 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5374_6
timestamp 1731220636
transform 1 0 1528 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5373_6
timestamp 1731220636
transform 1 0 1464 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5372_6
timestamp 1731220636
transform 1 0 1408 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5371_6
timestamp 1731220636
transform 1 0 1352 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5370_6
timestamp 1731220636
transform 1 0 1568 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5369_6
timestamp 1731220636
transform 1 0 1480 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5368_6
timestamp 1731220636
transform 1 0 1400 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5367_6
timestamp 1731220636
transform 1 0 1336 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5366_6
timestamp 1731220636
transform 1 0 1296 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5365_6
timestamp 1731220636
transform 1 0 1296 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5364_6
timestamp 1731220636
transform 1 0 1184 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5363_6
timestamp 1731220636
transform 1 0 1144 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5362_6
timestamp 1731220636
transform 1 0 1088 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5361_6
timestamp 1731220636
transform 1 0 1032 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5360_6
timestamp 1731220636
transform 1 0 976 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5359_6
timestamp 1731220636
transform 1 0 912 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5358_6
timestamp 1731220636
transform 1 0 848 0 -1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5357_6
timestamp 1731220636
transform 1 0 1184 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5356_6
timestamp 1731220636
transform 1 0 1128 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5355_6
timestamp 1731220636
transform 1 0 1072 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5354_6
timestamp 1731220636
transform 1 0 1016 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5353_6
timestamp 1731220636
transform 1 0 968 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5352_6
timestamp 1731220636
transform 1 0 912 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5351_6
timestamp 1731220636
transform 1 0 848 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5350_6
timestamp 1731220636
transform 1 0 776 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5349_6
timestamp 1731220636
transform 1 0 1016 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5348_6
timestamp 1731220636
transform 1 0 952 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5347_6
timestamp 1731220636
transform 1 0 896 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5346_6
timestamp 1731220636
transform 1 0 840 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5345_6
timestamp 1731220636
transform 1 0 776 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5344_6
timestamp 1731220636
transform 1 0 712 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5343_6
timestamp 1731220636
transform 1 0 640 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5342_6
timestamp 1731220636
transform 1 0 880 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5341_6
timestamp 1731220636
transform 1 0 824 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5340_6
timestamp 1731220636
transform 1 0 768 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5339_6
timestamp 1731220636
transform 1 0 712 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5338_6
timestamp 1731220636
transform 1 0 664 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5337_6
timestamp 1731220636
transform 1 0 608 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5336_6
timestamp 1731220636
transform 1 0 552 0 1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5335_6
timestamp 1731220636
transform 1 0 768 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5334_6
timestamp 1731220636
transform 1 0 720 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5333_6
timestamp 1731220636
transform 1 0 672 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5332_6
timestamp 1731220636
transform 1 0 624 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5331_6
timestamp 1731220636
transform 1 0 576 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5330_6
timestamp 1731220636
transform 1 0 528 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5329_6
timestamp 1731220636
transform 1 0 480 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5328_6
timestamp 1731220636
transform 1 0 584 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5327_6
timestamp 1731220636
transform 1 0 624 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5326_6
timestamp 1731220636
transform 1 0 672 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5325_6
timestamp 1731220636
transform 1 0 720 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5324_6
timestamp 1731220636
transform 1 0 768 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5323_6
timestamp 1731220636
transform 1 0 912 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5322_6
timestamp 1731220636
transform 1 0 864 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5321_6
timestamp 1731220636
transform 1 0 816 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5320_6
timestamp 1731220636
transform 1 0 784 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5319_6
timestamp 1731220636
transform 1 0 720 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5318_6
timestamp 1731220636
transform 1 0 648 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5317_6
timestamp 1731220636
transform 1 0 840 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5316_6
timestamp 1731220636
transform 1 0 1016 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5315_6
timestamp 1731220636
transform 1 0 952 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5314_6
timestamp 1731220636
transform 1 0 896 0 -1 240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5313_6
timestamp 1731220636
transform 1 0 720 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5312_6
timestamp 1731220636
transform 1 0 672 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5311_6
timestamp 1731220636
transform 1 0 624 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5310_6
timestamp 1731220636
transform 1 0 760 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5309_6
timestamp 1731220636
transform 1 0 800 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5308_6
timestamp 1731220636
transform 1 0 840 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5307_6
timestamp 1731220636
transform 1 0 880 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5306_6
timestamp 1731220636
transform 1 0 920 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5305_6
timestamp 1731220636
transform 1 0 968 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5304_6
timestamp 1731220636
transform 1 0 1016 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5303_6
timestamp 1731220636
transform 1 0 1064 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5302_6
timestamp 1731220636
transform 1 0 1104 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5301_6
timestamp 1731220636
transform 1 0 1144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5300_6
timestamp 1731220636
transform 1 0 1184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5299_6
timestamp 1731220636
transform 1 0 1296 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5298_6
timestamp 1731220636
transform 1 0 1336 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5297_6
timestamp 1731220636
transform 1 0 1376 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5296_6
timestamp 1731220636
transform 1 0 1416 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5295_6
timestamp 1731220636
transform 1 0 1456 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5294_6
timestamp 1731220636
transform 1 0 1640 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5293_6
timestamp 1731220636
transform 1 0 1576 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5292_6
timestamp 1731220636
transform 1 0 1512 0 1 92
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5291_6
timestamp 1731220636
transform 1 0 1440 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5290_6
timestamp 1731220636
transform 1 0 1400 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5289_6
timestamp 1731220636
transform 1 0 1360 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5288_6
timestamp 1731220636
transform 1 0 1488 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5287_6
timestamp 1731220636
transform 1 0 1544 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5286_6
timestamp 1731220636
transform 1 0 1600 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5285_6
timestamp 1731220636
transform 1 0 1664 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5284_6
timestamp 1731220636
transform 1 0 1736 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5283_6
timestamp 1731220636
transform 1 0 1688 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5282_6
timestamp 1731220636
transform 1 0 1648 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5281_6
timestamp 1731220636
transform 1 0 1608 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5280_6
timestamp 1731220636
transform 1 0 1568 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5279_6
timestamp 1731220636
transform 1 0 1528 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5278_6
timestamp 1731220636
transform 1 0 1488 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5277_6
timestamp 1731220636
transform 1 0 1584 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5276_6
timestamp 1731220636
transform 1 0 1528 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5275_6
timestamp 1731220636
transform 1 0 1480 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5274_6
timestamp 1731220636
transform 1 0 1440 0 -1 388
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5273_6
timestamp 1731220636
transform 1 0 1520 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5272_6
timestamp 1731220636
transform 1 0 1456 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5271_6
timestamp 1731220636
transform 1 0 1392 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5270_6
timestamp 1731220636
transform 1 0 1336 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5269_6
timestamp 1731220636
transform 1 0 1296 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5268_6
timestamp 1731220636
transform 1 0 1296 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5267_6
timestamp 1731220636
transform 1 0 1184 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5266_6
timestamp 1731220636
transform 1 0 1144 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5265_6
timestamp 1731220636
transform 1 0 1080 0 -1 524
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5264_6
timestamp 1731220636
transform 1 0 1368 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5263_6
timestamp 1731220636
transform 1 0 1472 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5262_6
timestamp 1731220636
transform 1 0 1576 0 -1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5261_6
timestamp 1731220636
transform 1 0 1488 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5260_6
timestamp 1731220636
transform 1 0 1448 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5259_6
timestamp 1731220636
transform 1 0 1408 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5258_6
timestamp 1731220636
transform 1 0 1536 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5257_6
timestamp 1731220636
transform 1 0 1720 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5256_6
timestamp 1731220636
transform 1 0 1656 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5255_6
timestamp 1731220636
transform 1 0 1592 0 1 532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5254_6
timestamp 1731220636
transform 1 0 1504 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5253_6
timestamp 1731220636
transform 1 0 1392 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5252_6
timestamp 1731220636
transform 1 0 1616 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5251_6
timestamp 1731220636
transform 1 0 1720 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5250_6
timestamp 1731220636
transform 1 0 1744 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5249_6
timestamp 1731220636
transform 1 0 1656 0 1 676
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5248_6
timestamp 1731220636
transform 1 0 1640 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5247_6
timestamp 1731220636
transform 1 0 1584 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5246_6
timestamp 1731220636
transform 1 0 1696 0 -1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5245_6
timestamp 1731220636
transform 1 0 1704 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5244_6
timestamp 1731220636
transform 1 0 1648 0 1 824
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5243_6
timestamp 1731220636
transform 1 0 1584 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5242_6
timestamp 1731220636
transform 1 0 1672 0 -1 960
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5241_6
timestamp 1731220636
transform 1 0 1768 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5240_6
timestamp 1731220636
transform 1 0 1728 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5239_6
timestamp 1731220636
transform 1 0 1688 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5238_6
timestamp 1731220636
transform 1 0 1648 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5237_6
timestamp 1731220636
transform 1 0 1608 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5236_6
timestamp 1731220636
transform 1 0 1568 0 1 968
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5235_6
timestamp 1731220636
transform 1 0 1720 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5234_6
timestamp 1731220636
transform 1 0 1664 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5233_6
timestamp 1731220636
transform 1 0 1608 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5232_6
timestamp 1731220636
transform 1 0 1552 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5231_6
timestamp 1731220636
transform 1 0 1504 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5230_6
timestamp 1731220636
transform 1 0 1464 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5229_6
timestamp 1731220636
transform 1 0 1424 0 -1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5228_6
timestamp 1731220636
transform 1 0 1792 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5227_6
timestamp 1731220636
transform 1 0 1680 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5226_6
timestamp 1731220636
transform 1 0 1576 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5225_6
timestamp 1731220636
transform 1 0 1480 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5224_6
timestamp 1731220636
transform 1 0 1400 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5223_6
timestamp 1731220636
transform 1 0 1336 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5222_6
timestamp 1731220636
transform 1 0 1296 0 1 1104
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5221_6
timestamp 1731220636
transform 1 0 1296 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5220_6
timestamp 1731220636
transform 1 0 1368 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5219_6
timestamp 1731220636
transform 1 0 1472 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5218_6
timestamp 1731220636
transform 1 0 1680 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5217_6
timestamp 1731220636
transform 1 0 1576 0 -1 1240
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5216_6
timestamp 1731220636
transform 1 0 1536 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5215_6
timestamp 1731220636
transform 1 0 1496 0 1 1248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5214_6
timestamp 1731220636
transform 1 0 1456 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5213_6
timestamp 1731220636
transform 1 0 1392 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5212_6
timestamp 1731220636
transform 1 0 1336 0 -1 1384
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5211_6
timestamp 1731220636
transform 1 0 1368 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5210_6
timestamp 1731220636
transform 1 0 1456 0 1 1392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5209_6
timestamp 1731220636
transform 1 0 1496 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5208_6
timestamp 1731220636
transform 1 0 1408 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5207_6
timestamp 1731220636
transform 1 0 1328 0 -1 1528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5206_6
timestamp 1731220636
transform 1 0 1320 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5205_6
timestamp 1731220636
transform 1 0 1392 0 1 1532
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5204_6
timestamp 1731220636
transform 1 0 1440 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5203_6
timestamp 1731220636
transform 1 0 1352 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5202_6
timestamp 1731220636
transform 1 0 1296 0 -1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5201_6
timestamp 1731220636
transform 1 0 1344 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5200_6
timestamp 1731220636
transform 1 0 1296 0 1 1668
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5199_6
timestamp 1731220636
transform 1 0 1184 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5198_6
timestamp 1731220636
transform 1 0 1144 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5197_6
timestamp 1731220636
transform 1 0 1080 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5196_6
timestamp 1731220636
transform 1 0 1024 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5195_6
timestamp 1731220636
transform 1 0 1184 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5194_6
timestamp 1731220636
transform 1 0 1128 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5193_6
timestamp 1731220636
transform 1 0 1056 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5192_6
timestamp 1731220636
transform 1 0 984 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5191_6
timestamp 1731220636
transform 1 0 904 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5190_6
timestamp 1731220636
transform 1 0 1112 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5189_6
timestamp 1731220636
transform 1 0 1032 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5188_6
timestamp 1731220636
transform 1 0 952 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5187_6
timestamp 1731220636
transform 1 0 872 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5186_6
timestamp 1731220636
transform 1 0 1056 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5185_6
timestamp 1731220636
transform 1 0 992 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5184_6
timestamp 1731220636
transform 1 0 928 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5183_6
timestamp 1731220636
transform 1 0 864 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5182_6
timestamp 1731220636
transform 1 0 952 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5181_6
timestamp 1731220636
transform 1 0 1008 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5180_6
timestamp 1731220636
transform 1 0 1064 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5179_6
timestamp 1731220636
transform 1 0 1136 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5178_6
timestamp 1731220636
transform 1 0 1072 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5177_6
timestamp 1731220636
transform 1 0 1016 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5176_6
timestamp 1731220636
transform 1 0 960 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5175_6
timestamp 1731220636
transform 1 0 904 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5174_6
timestamp 1731220636
transform 1 0 848 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5173_6
timestamp 1731220636
transform 1 0 896 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5172_6
timestamp 1731220636
transform 1 0 840 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5171_6
timestamp 1731220636
transform 1 0 792 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5170_6
timestamp 1731220636
transform 1 0 752 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5169_6
timestamp 1731220636
transform 1 0 688 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5168_6
timestamp 1731220636
transform 1 0 808 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5167_6
timestamp 1731220636
transform 1 0 792 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5166_6
timestamp 1731220636
transform 1 0 712 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5165_6
timestamp 1731220636
transform 1 0 632 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5164_6
timestamp 1731220636
transform 1 0 624 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5163_6
timestamp 1731220636
transform 1 0 720 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5162_6
timestamp 1731220636
transform 1 0 816 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5161_6
timestamp 1731220636
transform 1 0 744 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5160_6
timestamp 1731220636
transform 1 0 656 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5159_6
timestamp 1731220636
transform 1 0 824 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5158_6
timestamp 1731220636
transform 1 0 896 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5157_6
timestamp 1731220636
transform 1 0 960 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5156_6
timestamp 1731220636
transform 1 0 1152 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5155_6
timestamp 1731220636
transform 1 0 1080 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5154_6
timestamp 1731220636
transform 1 0 1008 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5153_6
timestamp 1731220636
transform 1 0 944 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5152_6
timestamp 1731220636
transform 1 0 872 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5151_6
timestamp 1731220636
transform 1 0 792 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5150_6
timestamp 1731220636
transform 1 0 704 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5149_6
timestamp 1731220636
transform 1 0 992 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5148_6
timestamp 1731220636
transform 1 0 936 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5147_6
timestamp 1731220636
transform 1 0 880 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5146_6
timestamp 1731220636
transform 1 0 824 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5145_6
timestamp 1731220636
transform 1 0 768 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5144_6
timestamp 1731220636
transform 1 0 712 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5143_6
timestamp 1731220636
transform 1 0 656 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5142_6
timestamp 1731220636
transform 1 0 920 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5141_6
timestamp 1731220636
transform 1 0 880 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5140_6
timestamp 1731220636
transform 1 0 840 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5139_6
timestamp 1731220636
transform 1 0 800 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5138_6
timestamp 1731220636
transform 1 0 760 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5137_6
timestamp 1731220636
transform 1 0 720 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5136_6
timestamp 1731220636
transform 1 0 680 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5135_6
timestamp 1731220636
transform 1 0 640 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5134_6
timestamp 1731220636
transform 1 0 600 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5133_6
timestamp 1731220636
transform 1 0 560 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5132_6
timestamp 1731220636
transform 1 0 520 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5131_6
timestamp 1731220636
transform 1 0 480 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5130_6
timestamp 1731220636
transform 1 0 440 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5129_6
timestamp 1731220636
transform 1 0 400 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5128_6
timestamp 1731220636
transform 1 0 360 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5127_6
timestamp 1731220636
transform 1 0 320 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5126_6
timestamp 1731220636
transform 1 0 592 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5125_6
timestamp 1731220636
transform 1 0 528 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5124_6
timestamp 1731220636
transform 1 0 464 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5123_6
timestamp 1731220636
transform 1 0 408 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5122_6
timestamp 1731220636
transform 1 0 352 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5121_6
timestamp 1731220636
transform 1 0 304 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5120_6
timestamp 1731220636
transform 1 0 264 0 1 1568
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5119_6
timestamp 1731220636
transform 1 0 608 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5118_6
timestamp 1731220636
transform 1 0 504 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5117_6
timestamp 1731220636
transform 1 0 408 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5116_6
timestamp 1731220636
transform 1 0 312 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5115_6
timestamp 1731220636
transform 1 0 232 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5114_6
timestamp 1731220636
transform 1 0 168 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5113_6
timestamp 1731220636
transform 1 0 128 0 -1 1708
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5112_6
timestamp 1731220636
transform 1 0 560 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5111_6
timestamp 1731220636
transform 1 0 464 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5110_6
timestamp 1731220636
transform 1 0 368 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5109_6
timestamp 1731220636
transform 1 0 280 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5108_6
timestamp 1731220636
transform 1 0 208 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5107_6
timestamp 1731220636
transform 1 0 168 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5106_6
timestamp 1731220636
transform 1 0 128 0 1 1712
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5105_6
timestamp 1731220636
transform 1 0 128 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5104_6
timestamp 1731220636
transform 1 0 168 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5103_6
timestamp 1731220636
transform 1 0 208 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5102_6
timestamp 1731220636
transform 1 0 264 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5101_6
timestamp 1731220636
transform 1 0 528 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5100_6
timestamp 1731220636
transform 1 0 432 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_599_6
timestamp 1731220636
transform 1 0 344 0 -1 1848
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_598_6
timestamp 1731220636
transform 1 0 256 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_597_6
timestamp 1731220636
transform 1 0 208 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_596_6
timestamp 1731220636
transform 1 0 168 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_595_6
timestamp 1731220636
transform 1 0 312 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_594_6
timestamp 1731220636
transform 1 0 384 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_593_6
timestamp 1731220636
transform 1 0 544 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_592_6
timestamp 1731220636
transform 1 0 464 0 1 1856
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_591_6
timestamp 1731220636
transform 1 0 448 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_590_6
timestamp 1731220636
transform 1 0 400 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_589_6
timestamp 1731220636
transform 1 0 360 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_588_6
timestamp 1731220636
transform 1 0 504 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_587_6
timestamp 1731220636
transform 1 0 560 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_586_6
timestamp 1731220636
transform 1 0 624 0 -1 1996
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_585_6
timestamp 1731220636
transform 1 0 680 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_584_6
timestamp 1731220636
transform 1 0 736 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_583_6
timestamp 1731220636
transform 1 0 720 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_582_6
timestamp 1731220636
transform 1 0 784 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_581_6
timestamp 1731220636
transform 1 0 776 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_580_6
timestamp 1731220636
transform 1 0 712 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_579_6
timestamp 1731220636
transform 1 0 904 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_578_6
timestamp 1731220636
transform 1 0 840 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_577_6
timestamp 1731220636
transform 1 0 824 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_576_6
timestamp 1731220636
transform 1 0 904 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_575_6
timestamp 1731220636
transform 1 0 984 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_574_6
timestamp 1731220636
transform 1 0 1024 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_573_6
timestamp 1731220636
transform 1 0 952 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_572_6
timestamp 1731220636
transform 1 0 880 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_571_6
timestamp 1731220636
transform 1 0 816 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_570_6
timestamp 1731220636
transform 1 0 1040 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_569_6
timestamp 1731220636
transform 1 0 984 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_568_6
timestamp 1731220636
transform 1 0 928 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_567_6
timestamp 1731220636
transform 1 0 880 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_566_6
timestamp 1731220636
transform 1 0 832 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_565_6
timestamp 1731220636
transform 1 0 920 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_564_6
timestamp 1731220636
transform 1 0 824 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_563_6
timestamp 1731220636
transform 1 0 736 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_562_6
timestamp 1731220636
transform 1 0 648 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_561_6
timestamp 1731220636
transform 1 0 784 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_560_6
timestamp 1731220636
transform 1 0 728 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_559_6
timestamp 1731220636
transform 1 0 672 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_558_6
timestamp 1731220636
transform 1 0 608 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_557_6
timestamp 1731220636
transform 1 0 536 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_556_6
timestamp 1731220636
transform 1 0 592 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_555_6
timestamp 1731220636
transform 1 0 672 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_554_6
timestamp 1731220636
transform 1 0 744 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_553_6
timestamp 1731220636
transform 1 0 752 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_552_6
timestamp 1731220636
transform 1 0 680 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_551_6
timestamp 1731220636
transform 1 0 608 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_550_6
timestamp 1731220636
transform 1 0 528 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_549_6
timestamp 1731220636
transform 1 0 656 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_548_6
timestamp 1731220636
transform 1 0 600 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_547_6
timestamp 1731220636
transform 1 0 544 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_546_6
timestamp 1731220636
transform 1 0 544 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_545_6
timestamp 1731220636
transform 1 0 600 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_544_6
timestamp 1731220636
transform 1 0 656 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_543_6
timestamp 1731220636
transform 1 0 624 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_542_6
timestamp 1731220636
transform 1 0 576 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_541_6
timestamp 1731220636
transform 1 0 536 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_540_6
timestamp 1731220636
transform 1 0 496 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_539_6
timestamp 1731220636
transform 1 0 456 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_538_6
timestamp 1731220636
transform 1 0 416 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_537_6
timestamp 1731220636
transform 1 0 376 0 1 2004
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_536_6
timestamp 1731220636
transform 1 0 496 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_535_6
timestamp 1731220636
transform 1 0 456 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_534_6
timestamp 1731220636
transform 1 0 416 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_533_6
timestamp 1731220636
transform 1 0 376 0 -1 2140
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_532_6
timestamp 1731220636
transform 1 0 488 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_531_6
timestamp 1731220636
transform 1 0 424 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_530_6
timestamp 1731220636
transform 1 0 368 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_529_6
timestamp 1731220636
transform 1 0 320 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_528_6
timestamp 1731220636
transform 1 0 280 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_527_6
timestamp 1731220636
transform 1 0 240 0 1 2148
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_526_6
timestamp 1731220636
transform 1 0 448 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_525_6
timestamp 1731220636
transform 1 0 368 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_524_6
timestamp 1731220636
transform 1 0 296 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_523_6
timestamp 1731220636
transform 1 0 224 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_522_6
timestamp 1731220636
transform 1 0 168 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_521_6
timestamp 1731220636
transform 1 0 128 0 -1 2284
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_520_6
timestamp 1731220636
transform 1 0 264 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_519_6
timestamp 1731220636
transform 1 0 208 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_518_6
timestamp 1731220636
transform 1 0 168 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_517_6
timestamp 1731220636
transform 1 0 128 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_516_6
timestamp 1731220636
transform 1 0 344 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_515_6
timestamp 1731220636
transform 1 0 424 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_514_6
timestamp 1731220636
transform 1 0 512 0 1 2288
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_513_6
timestamp 1731220636
transform 1 0 464 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_512_6
timestamp 1731220636
transform 1 0 384 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_511_6
timestamp 1731220636
transform 1 0 312 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_510_6
timestamp 1731220636
transform 1 0 240 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_59_6
timestamp 1731220636
transform 1 0 176 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_58_6
timestamp 1731220636
transform 1 0 128 0 -1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_57_6
timestamp 1731220636
transform 1 0 560 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_56_6
timestamp 1731220636
transform 1 0 472 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_55_6
timestamp 1731220636
transform 1 0 384 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_54_6
timestamp 1731220636
transform 1 0 304 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_53_6
timestamp 1731220636
transform 1 0 248 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_52_6
timestamp 1731220636
transform 1 0 208 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_51_6
timestamp 1731220636
transform 1 0 168 0 1 2432
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_50_6
timestamp 1731220636
transform 1 0 128 0 1 2432
box 4 6 36 64
<< end >>
