magic
tech sky130l
timestamp 1730421221
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 26 13 27
rect 8 23 9 26
rect 12 23 13 26
rect 8 19 13 23
rect 15 23 20 27
rect 15 20 16 23
rect 19 20 20 23
rect 15 19 20 20
<< pdc >>
rect 9 23 12 26
rect 16 20 19 23
<< ptransistor >>
rect 13 19 15 27
<< polysilicon >>
rect 13 34 20 35
rect 13 31 16 34
rect 19 31 20 34
rect 13 30 20 31
rect 13 27 15 30
rect 13 12 15 19
rect 13 4 15 6
<< pc >>
rect 16 31 19 34
<< m1 >>
rect 16 34 20 35
rect 8 31 12 32
rect 8 28 9 31
rect 19 31 20 34
rect 16 28 20 31
rect 8 26 12 28
rect 8 23 9 26
rect 8 22 12 23
rect 16 23 20 24
rect 19 20 20 23
rect 16 11 20 20
rect 8 10 12 11
rect 8 7 9 10
rect 8 4 12 7
rect 19 8 20 11
rect 16 4 20 8
<< m2c >>
rect 9 28 12 31
rect 9 7 12 10
<< m2 >>
rect 8 31 13 32
rect 8 28 9 31
rect 12 28 13 31
rect 8 27 13 28
rect 8 10 13 11
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
<< labels >>
rlabel m1 s 19 31 20 34 6 A
port 1 nsew signal input
rlabel m1 s 16 28 20 31 6 A
port 1 nsew signal input
rlabel m1 s 16 31 19 34 6 A
port 1 nsew signal input
rlabel m1 s 16 34 20 35 6 A
port 1 nsew signal input
rlabel m1 s 19 8 20 11 6 Y
port 2 nsew signal output
rlabel m1 s 19 20 20 23 6 Y
port 2 nsew signal output
rlabel m1 s 16 8 19 11 6 Y
port 2 nsew signal output
rlabel m1 s 16 11 20 20 6 Y
port 2 nsew signal output
rlabel m1 s 16 20 19 23 6 Y
port 2 nsew signal output
rlabel m1 s 16 23 20 24 6 Y
port 2 nsew signal output
rlabel m1 s 16 4 20 8 6 Y
port 2 nsew signal output
rlabel m2 s 12 28 13 31 6 Vdd
port 3 nsew power input
rlabel m2 s 9 28 12 31 6 Vdd
port 3 nsew power input
rlabel m2 s 8 27 13 28 6 Vdd
port 3 nsew power input
rlabel m2 s 8 28 9 31 6 Vdd
port 3 nsew power input
rlabel m2 s 8 31 13 32 6 Vdd
port 3 nsew power input
rlabel m2c s 9 28 12 31 6 Vdd
port 3 nsew power input
rlabel m1 s 9 23 12 26 6 Vdd
port 3 nsew power input
rlabel m1 s 9 28 12 31 6 Vdd
port 3 nsew power input
rlabel m1 s 8 22 12 23 6 Vdd
port 3 nsew power input
rlabel m1 s 8 23 9 26 6 Vdd
port 3 nsew power input
rlabel m1 s 8 26 12 28 6 Vdd
port 3 nsew power input
rlabel m1 s 8 28 9 31 6 Vdd
port 3 nsew power input
rlabel m1 s 8 31 12 32 6 Vdd
port 3 nsew power input
rlabel m2 s 12 7 13 10 6 GND
port 4 nsew ground input
rlabel m2 s 9 7 12 10 6 GND
port 4 nsew ground input
rlabel m2 s 8 6 13 7 6 GND
port 4 nsew ground input
rlabel m2 s 8 7 9 10 6 GND
port 4 nsew ground input
rlabel m2 s 8 10 13 11 6 GND
port 4 nsew ground input
rlabel m2c s 9 7 12 10 6 GND
port 4 nsew ground input
rlabel m1 s 9 7 12 10 6 GND
port 4 nsew ground input
rlabel m1 s 8 4 12 7 6 GND
port 4 nsew ground input
rlabel m1 s 8 7 9 10 6 GND
port 4 nsew ground input
rlabel m1 s 8 10 12 11 6 GND
port 4 nsew ground input
rlabel space 0 0 24 40 3 prboundary
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 16 9 16 9 3 Y
rlabel ndiffusion 16 12 16 12 3 Y
rlabel pdiffusion 16 20 16 20 3 Y
rlabel pdiffusion 16 21 16 21 3 Y
rlabel pdiffusion 16 24 16 24 3 Y
rlabel pdiffusion 13 24 13 24 3 Vdd
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 13 14 13 3 A
rlabel ptransistor 14 20 14 20 3 A
rlabel polysilicon 14 28 14 28 3 A
rlabel polysilicon 14 31 14 31 3 A
rlabel polysilicon 14 32 14 32 3 A
rlabel polysilicon 14 35 14 35 3 A
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 20 9 20 9 3 Y
port 2 e default output
rlabel m1 20 21 20 21 3 Y
port 2 e default output
rlabel m1 20 32 20 32 3 A
port 1 e default input
rlabel ndc 17 9 17 9 3 Y
port 2 e default output
rlabel m1 17 12 17 12 3 Y
port 2 e default output
rlabel pdc 17 21 17 21 3 Y
port 2 e default output
rlabel m1 17 24 17 24 3 Y
port 2 e default output
rlabel m1 17 29 17 29 3 A
port 1 e default input
rlabel pc 17 32 17 32 3 A
port 1 e
rlabel m1 17 35 17 35 3 A
port 1 e
rlabel m1 17 5 17 5 3 Y
port 2 e
rlabel pdc 10 24 10 24 3 Vdd
rlabel m1 9 5 9 5 3 GND
rlabel m1 9 23 9 23 3 Vdd
rlabel m1 9 24 9 24 3 Vdd
rlabel m1 9 27 9 27 3 Vdd
rlabel m2 13 8 13 8 3 GND
rlabel m2 13 29 13 29 3 Vdd
rlabel m2c 10 8 10 8 3 GND
rlabel m2c 10 29 10 29 3 Vdd
rlabel m2 9 7 9 7 3 GND
rlabel m2 9 8 9 8 3 GND
rlabel m2 9 11 9 11 3 GND
rlabel m2 9 28 9 28 3 Vdd
rlabel m2 9 29 9 29 3 Vdd
rlabel m2 9 32 9 32 3 Vdd
<< properties >>
string LEFclass CORE
string LEFsite CoreSite
string FIXED_BBOX 0 0 24 40
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
