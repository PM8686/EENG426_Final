magic
tech sky130l
timestamp 1731220429
<< m2 >>
rect 110 5693 116 5694
rect 1934 5693 1940 5694
rect 110 5689 111 5693
rect 115 5689 116 5693
rect 110 5688 116 5689
rect 158 5692 164 5693
rect 158 5688 159 5692
rect 163 5688 164 5692
rect 158 5687 164 5688
rect 302 5692 308 5693
rect 302 5688 303 5692
rect 307 5688 308 5692
rect 302 5687 308 5688
rect 502 5692 508 5693
rect 502 5688 503 5692
rect 507 5688 508 5692
rect 502 5687 508 5688
rect 726 5692 732 5693
rect 726 5688 727 5692
rect 731 5688 732 5692
rect 726 5687 732 5688
rect 982 5692 988 5693
rect 982 5688 983 5692
rect 987 5688 988 5692
rect 982 5687 988 5688
rect 1254 5692 1260 5693
rect 1254 5688 1255 5692
rect 1259 5688 1260 5692
rect 1254 5687 1260 5688
rect 1542 5692 1548 5693
rect 1542 5688 1543 5692
rect 1547 5688 1548 5692
rect 1542 5687 1548 5688
rect 1814 5692 1820 5693
rect 1814 5688 1815 5692
rect 1819 5688 1820 5692
rect 1934 5689 1935 5693
rect 1939 5689 1940 5693
rect 1934 5688 1940 5689
rect 1814 5687 1820 5688
rect 130 5677 136 5678
rect 110 5676 116 5677
rect 110 5672 111 5676
rect 115 5672 116 5676
rect 130 5673 131 5677
rect 135 5673 136 5677
rect 130 5672 136 5673
rect 274 5677 280 5678
rect 274 5673 275 5677
rect 279 5673 280 5677
rect 274 5672 280 5673
rect 474 5677 480 5678
rect 474 5673 475 5677
rect 479 5673 480 5677
rect 474 5672 480 5673
rect 698 5677 704 5678
rect 698 5673 699 5677
rect 703 5673 704 5677
rect 698 5672 704 5673
rect 954 5677 960 5678
rect 954 5673 955 5677
rect 959 5673 960 5677
rect 954 5672 960 5673
rect 1226 5677 1232 5678
rect 1226 5673 1227 5677
rect 1231 5673 1232 5677
rect 1226 5672 1232 5673
rect 1514 5677 1520 5678
rect 1514 5673 1515 5677
rect 1519 5673 1520 5677
rect 1514 5672 1520 5673
rect 1786 5677 1792 5678
rect 1786 5673 1787 5677
rect 1791 5673 1792 5677
rect 1786 5672 1792 5673
rect 1934 5676 1940 5677
rect 1934 5672 1935 5676
rect 1939 5672 1940 5676
rect 110 5671 116 5672
rect 1934 5671 1940 5672
rect 1974 5628 1980 5629
rect 3798 5628 3804 5629
rect 1974 5624 1975 5628
rect 1979 5624 1980 5628
rect 1974 5623 1980 5624
rect 1994 5627 2000 5628
rect 1994 5623 1995 5627
rect 1999 5623 2000 5627
rect 1994 5622 2000 5623
rect 2178 5627 2184 5628
rect 2178 5623 2179 5627
rect 2183 5623 2184 5627
rect 2178 5622 2184 5623
rect 2386 5627 2392 5628
rect 2386 5623 2387 5627
rect 2391 5623 2392 5627
rect 2386 5622 2392 5623
rect 2586 5627 2592 5628
rect 2586 5623 2587 5627
rect 2591 5623 2592 5627
rect 2586 5622 2592 5623
rect 2778 5627 2784 5628
rect 2778 5623 2779 5627
rect 2783 5623 2784 5627
rect 2778 5622 2784 5623
rect 2962 5627 2968 5628
rect 2962 5623 2963 5627
rect 2967 5623 2968 5627
rect 2962 5622 2968 5623
rect 3146 5627 3152 5628
rect 3146 5623 3147 5627
rect 3151 5623 3152 5627
rect 3146 5622 3152 5623
rect 3322 5627 3328 5628
rect 3322 5623 3323 5627
rect 3327 5623 3328 5627
rect 3322 5622 3328 5623
rect 3498 5627 3504 5628
rect 3498 5623 3499 5627
rect 3503 5623 3504 5627
rect 3498 5622 3504 5623
rect 3650 5627 3656 5628
rect 3650 5623 3651 5627
rect 3655 5623 3656 5627
rect 3798 5624 3799 5628
rect 3803 5624 3804 5628
rect 3798 5623 3804 5624
rect 3650 5622 3656 5623
rect 2022 5612 2028 5613
rect 1974 5611 1980 5612
rect 1974 5607 1975 5611
rect 1979 5607 1980 5611
rect 2022 5608 2023 5612
rect 2027 5608 2028 5612
rect 2022 5607 2028 5608
rect 2206 5612 2212 5613
rect 2206 5608 2207 5612
rect 2211 5608 2212 5612
rect 2206 5607 2212 5608
rect 2414 5612 2420 5613
rect 2414 5608 2415 5612
rect 2419 5608 2420 5612
rect 2414 5607 2420 5608
rect 2614 5612 2620 5613
rect 2614 5608 2615 5612
rect 2619 5608 2620 5612
rect 2614 5607 2620 5608
rect 2806 5612 2812 5613
rect 2806 5608 2807 5612
rect 2811 5608 2812 5612
rect 2806 5607 2812 5608
rect 2990 5612 2996 5613
rect 2990 5608 2991 5612
rect 2995 5608 2996 5612
rect 2990 5607 2996 5608
rect 3174 5612 3180 5613
rect 3174 5608 3175 5612
rect 3179 5608 3180 5612
rect 3174 5607 3180 5608
rect 3350 5612 3356 5613
rect 3350 5608 3351 5612
rect 3355 5608 3356 5612
rect 3350 5607 3356 5608
rect 3526 5612 3532 5613
rect 3526 5608 3527 5612
rect 3531 5608 3532 5612
rect 3526 5607 3532 5608
rect 3678 5612 3684 5613
rect 3678 5608 3679 5612
rect 3683 5608 3684 5612
rect 3678 5607 3684 5608
rect 3798 5611 3804 5612
rect 3798 5607 3799 5611
rect 3803 5607 3804 5611
rect 1974 5606 1980 5607
rect 3798 5606 3804 5607
rect 3838 5584 3844 5585
rect 5662 5584 5668 5585
rect 3838 5580 3839 5584
rect 3843 5580 3844 5584
rect 3838 5579 3844 5580
rect 4290 5583 4296 5584
rect 4290 5579 4291 5583
rect 4295 5579 4296 5583
rect 4290 5578 4296 5579
rect 4426 5583 4432 5584
rect 4426 5579 4427 5583
rect 4431 5579 4432 5583
rect 4426 5578 4432 5579
rect 4562 5583 4568 5584
rect 4562 5579 4563 5583
rect 4567 5579 4568 5583
rect 4562 5578 4568 5579
rect 4698 5583 4704 5584
rect 4698 5579 4699 5583
rect 4703 5579 4704 5583
rect 4698 5578 4704 5579
rect 4834 5583 4840 5584
rect 4834 5579 4835 5583
rect 4839 5579 4840 5583
rect 4834 5578 4840 5579
rect 4970 5583 4976 5584
rect 4970 5579 4971 5583
rect 4975 5579 4976 5583
rect 4970 5578 4976 5579
rect 5106 5583 5112 5584
rect 5106 5579 5107 5583
rect 5111 5579 5112 5583
rect 5662 5580 5663 5584
rect 5667 5580 5668 5584
rect 5662 5579 5668 5580
rect 5106 5578 5112 5579
rect 4318 5568 4324 5569
rect 3838 5567 3844 5568
rect 3838 5563 3839 5567
rect 3843 5563 3844 5567
rect 4318 5564 4319 5568
rect 4323 5564 4324 5568
rect 4318 5563 4324 5564
rect 4454 5568 4460 5569
rect 4454 5564 4455 5568
rect 4459 5564 4460 5568
rect 4454 5563 4460 5564
rect 4590 5568 4596 5569
rect 4590 5564 4591 5568
rect 4595 5564 4596 5568
rect 4590 5563 4596 5564
rect 4726 5568 4732 5569
rect 4726 5564 4727 5568
rect 4731 5564 4732 5568
rect 4726 5563 4732 5564
rect 4862 5568 4868 5569
rect 4862 5564 4863 5568
rect 4867 5564 4868 5568
rect 4862 5563 4868 5564
rect 4998 5568 5004 5569
rect 4998 5564 4999 5568
rect 5003 5564 5004 5568
rect 4998 5563 5004 5564
rect 5134 5568 5140 5569
rect 5134 5564 5135 5568
rect 5139 5564 5140 5568
rect 5134 5563 5140 5564
rect 5662 5567 5668 5568
rect 5662 5563 5663 5567
rect 5667 5563 5668 5567
rect 3838 5562 3844 5563
rect 5662 5562 5668 5563
rect 1974 5553 1980 5554
rect 3798 5553 3804 5554
rect 1974 5549 1975 5553
rect 1979 5549 1980 5553
rect 1974 5548 1980 5549
rect 2262 5552 2268 5553
rect 2262 5548 2263 5552
rect 2267 5548 2268 5552
rect 2262 5547 2268 5548
rect 2502 5552 2508 5553
rect 2502 5548 2503 5552
rect 2507 5548 2508 5552
rect 2502 5547 2508 5548
rect 2742 5552 2748 5553
rect 2742 5548 2743 5552
rect 2747 5548 2748 5552
rect 2742 5547 2748 5548
rect 2982 5552 2988 5553
rect 2982 5548 2983 5552
rect 2987 5548 2988 5552
rect 2982 5547 2988 5548
rect 3222 5552 3228 5553
rect 3222 5548 3223 5552
rect 3227 5548 3228 5552
rect 3222 5547 3228 5548
rect 3462 5552 3468 5553
rect 3462 5548 3463 5552
rect 3467 5548 3468 5552
rect 3462 5547 3468 5548
rect 3678 5552 3684 5553
rect 3678 5548 3679 5552
rect 3683 5548 3684 5552
rect 3798 5549 3799 5553
rect 3803 5549 3804 5553
rect 3798 5548 3804 5549
rect 3678 5547 3684 5548
rect 110 5540 116 5541
rect 1934 5540 1940 5541
rect 110 5536 111 5540
rect 115 5536 116 5540
rect 110 5535 116 5536
rect 562 5539 568 5540
rect 562 5535 563 5539
rect 567 5535 568 5539
rect 562 5534 568 5535
rect 722 5539 728 5540
rect 722 5535 723 5539
rect 727 5535 728 5539
rect 722 5534 728 5535
rect 882 5539 888 5540
rect 882 5535 883 5539
rect 887 5535 888 5539
rect 882 5534 888 5535
rect 1050 5539 1056 5540
rect 1050 5535 1051 5539
rect 1055 5535 1056 5539
rect 1050 5534 1056 5535
rect 1226 5539 1232 5540
rect 1226 5535 1227 5539
rect 1231 5535 1232 5539
rect 1226 5534 1232 5535
rect 1402 5539 1408 5540
rect 1402 5535 1403 5539
rect 1407 5535 1408 5539
rect 1402 5534 1408 5535
rect 1578 5539 1584 5540
rect 1578 5535 1579 5539
rect 1583 5535 1584 5539
rect 1578 5534 1584 5535
rect 1762 5539 1768 5540
rect 1762 5535 1763 5539
rect 1767 5535 1768 5539
rect 1934 5536 1935 5540
rect 1939 5536 1940 5540
rect 2234 5537 2240 5538
rect 1934 5535 1940 5536
rect 1974 5536 1980 5537
rect 1762 5534 1768 5535
rect 1974 5532 1975 5536
rect 1979 5532 1980 5536
rect 2234 5533 2235 5537
rect 2239 5533 2240 5537
rect 2234 5532 2240 5533
rect 2474 5537 2480 5538
rect 2474 5533 2475 5537
rect 2479 5533 2480 5537
rect 2474 5532 2480 5533
rect 2714 5537 2720 5538
rect 2714 5533 2715 5537
rect 2719 5533 2720 5537
rect 2714 5532 2720 5533
rect 2954 5537 2960 5538
rect 2954 5533 2955 5537
rect 2959 5533 2960 5537
rect 2954 5532 2960 5533
rect 3194 5537 3200 5538
rect 3194 5533 3195 5537
rect 3199 5533 3200 5537
rect 3194 5532 3200 5533
rect 3434 5537 3440 5538
rect 3434 5533 3435 5537
rect 3439 5533 3440 5537
rect 3434 5532 3440 5533
rect 3650 5537 3656 5538
rect 3650 5533 3651 5537
rect 3655 5533 3656 5537
rect 3650 5532 3656 5533
rect 3798 5536 3804 5537
rect 3798 5532 3799 5536
rect 3803 5532 3804 5536
rect 1974 5531 1980 5532
rect 3798 5531 3804 5532
rect 590 5524 596 5525
rect 110 5523 116 5524
rect 110 5519 111 5523
rect 115 5519 116 5523
rect 590 5520 591 5524
rect 595 5520 596 5524
rect 590 5519 596 5520
rect 750 5524 756 5525
rect 750 5520 751 5524
rect 755 5520 756 5524
rect 750 5519 756 5520
rect 910 5524 916 5525
rect 910 5520 911 5524
rect 915 5520 916 5524
rect 910 5519 916 5520
rect 1078 5524 1084 5525
rect 1078 5520 1079 5524
rect 1083 5520 1084 5524
rect 1078 5519 1084 5520
rect 1254 5524 1260 5525
rect 1254 5520 1255 5524
rect 1259 5520 1260 5524
rect 1254 5519 1260 5520
rect 1430 5524 1436 5525
rect 1430 5520 1431 5524
rect 1435 5520 1436 5524
rect 1430 5519 1436 5520
rect 1606 5524 1612 5525
rect 1606 5520 1607 5524
rect 1611 5520 1612 5524
rect 1606 5519 1612 5520
rect 1790 5524 1796 5525
rect 1790 5520 1791 5524
rect 1795 5520 1796 5524
rect 1790 5519 1796 5520
rect 1934 5523 1940 5524
rect 1934 5519 1935 5523
rect 1939 5519 1940 5523
rect 110 5518 116 5519
rect 1934 5518 1940 5519
rect 3838 5509 3844 5510
rect 5662 5509 5668 5510
rect 3838 5505 3839 5509
rect 3843 5505 3844 5509
rect 3838 5504 3844 5505
rect 3886 5508 3892 5509
rect 3886 5504 3887 5508
rect 3891 5504 3892 5508
rect 3886 5503 3892 5504
rect 4126 5508 4132 5509
rect 4126 5504 4127 5508
rect 4131 5504 4132 5508
rect 4126 5503 4132 5504
rect 4374 5508 4380 5509
rect 4374 5504 4375 5508
rect 4379 5504 4380 5508
rect 4374 5503 4380 5504
rect 4614 5508 4620 5509
rect 4614 5504 4615 5508
rect 4619 5504 4620 5508
rect 4614 5503 4620 5504
rect 4846 5508 4852 5509
rect 4846 5504 4847 5508
rect 4851 5504 4852 5508
rect 4846 5503 4852 5504
rect 5078 5508 5084 5509
rect 5078 5504 5079 5508
rect 5083 5504 5084 5508
rect 5078 5503 5084 5504
rect 5310 5508 5316 5509
rect 5310 5504 5311 5508
rect 5315 5504 5316 5508
rect 5662 5505 5663 5509
rect 5667 5505 5668 5509
rect 5662 5504 5668 5505
rect 5310 5503 5316 5504
rect 3858 5493 3864 5494
rect 3838 5492 3844 5493
rect 3838 5488 3839 5492
rect 3843 5488 3844 5492
rect 3858 5489 3859 5493
rect 3863 5489 3864 5493
rect 3858 5488 3864 5489
rect 4098 5493 4104 5494
rect 4098 5489 4099 5493
rect 4103 5489 4104 5493
rect 4098 5488 4104 5489
rect 4346 5493 4352 5494
rect 4346 5489 4347 5493
rect 4351 5489 4352 5493
rect 4346 5488 4352 5489
rect 4586 5493 4592 5494
rect 4586 5489 4587 5493
rect 4591 5489 4592 5493
rect 4586 5488 4592 5489
rect 4818 5493 4824 5494
rect 4818 5489 4819 5493
rect 4823 5489 4824 5493
rect 4818 5488 4824 5489
rect 5050 5493 5056 5494
rect 5050 5489 5051 5493
rect 5055 5489 5056 5493
rect 5050 5488 5056 5489
rect 5282 5493 5288 5494
rect 5282 5489 5283 5493
rect 5287 5489 5288 5493
rect 5282 5488 5288 5489
rect 5662 5492 5668 5493
rect 5662 5488 5663 5492
rect 5667 5488 5668 5492
rect 3838 5487 3844 5488
rect 5662 5487 5668 5488
rect 110 5453 116 5454
rect 1934 5453 1940 5454
rect 110 5449 111 5453
rect 115 5449 116 5453
rect 110 5448 116 5449
rect 590 5452 596 5453
rect 590 5448 591 5452
rect 595 5448 596 5452
rect 590 5447 596 5448
rect 726 5452 732 5453
rect 726 5448 727 5452
rect 731 5448 732 5452
rect 726 5447 732 5448
rect 862 5452 868 5453
rect 862 5448 863 5452
rect 867 5448 868 5452
rect 862 5447 868 5448
rect 998 5452 1004 5453
rect 998 5448 999 5452
rect 1003 5448 1004 5452
rect 998 5447 1004 5448
rect 1134 5452 1140 5453
rect 1134 5448 1135 5452
rect 1139 5448 1140 5452
rect 1134 5447 1140 5448
rect 1270 5452 1276 5453
rect 1270 5448 1271 5452
rect 1275 5448 1276 5452
rect 1270 5447 1276 5448
rect 1406 5452 1412 5453
rect 1406 5448 1407 5452
rect 1411 5448 1412 5452
rect 1406 5447 1412 5448
rect 1542 5452 1548 5453
rect 1542 5448 1543 5452
rect 1547 5448 1548 5452
rect 1542 5447 1548 5448
rect 1678 5452 1684 5453
rect 1678 5448 1679 5452
rect 1683 5448 1684 5452
rect 1678 5447 1684 5448
rect 1814 5452 1820 5453
rect 1814 5448 1815 5452
rect 1819 5448 1820 5452
rect 1934 5449 1935 5453
rect 1939 5449 1940 5453
rect 1934 5448 1940 5449
rect 1814 5447 1820 5448
rect 562 5437 568 5438
rect 110 5436 116 5437
rect 110 5432 111 5436
rect 115 5432 116 5436
rect 562 5433 563 5437
rect 567 5433 568 5437
rect 562 5432 568 5433
rect 698 5437 704 5438
rect 698 5433 699 5437
rect 703 5433 704 5437
rect 698 5432 704 5433
rect 834 5437 840 5438
rect 834 5433 835 5437
rect 839 5433 840 5437
rect 834 5432 840 5433
rect 970 5437 976 5438
rect 970 5433 971 5437
rect 975 5433 976 5437
rect 970 5432 976 5433
rect 1106 5437 1112 5438
rect 1106 5433 1107 5437
rect 1111 5433 1112 5437
rect 1106 5432 1112 5433
rect 1242 5437 1248 5438
rect 1242 5433 1243 5437
rect 1247 5433 1248 5437
rect 1242 5432 1248 5433
rect 1378 5437 1384 5438
rect 1378 5433 1379 5437
rect 1383 5433 1384 5437
rect 1378 5432 1384 5433
rect 1514 5437 1520 5438
rect 1514 5433 1515 5437
rect 1519 5433 1520 5437
rect 1514 5432 1520 5433
rect 1650 5437 1656 5438
rect 1650 5433 1651 5437
rect 1655 5433 1656 5437
rect 1650 5432 1656 5433
rect 1786 5437 1792 5438
rect 1786 5433 1787 5437
rect 1791 5433 1792 5437
rect 1786 5432 1792 5433
rect 1934 5436 1940 5437
rect 1934 5432 1935 5436
rect 1939 5432 1940 5436
rect 110 5431 116 5432
rect 1934 5431 1940 5432
rect 1974 5396 1980 5397
rect 3798 5396 3804 5397
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 2426 5395 2432 5396
rect 2426 5391 2427 5395
rect 2431 5391 2432 5395
rect 2426 5390 2432 5391
rect 2642 5395 2648 5396
rect 2642 5391 2643 5395
rect 2647 5391 2648 5395
rect 2642 5390 2648 5391
rect 2858 5395 2864 5396
rect 2858 5391 2859 5395
rect 2863 5391 2864 5395
rect 2858 5390 2864 5391
rect 3074 5395 3080 5396
rect 3074 5391 3075 5395
rect 3079 5391 3080 5395
rect 3074 5390 3080 5391
rect 3290 5395 3296 5396
rect 3290 5391 3291 5395
rect 3295 5391 3296 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3290 5390 3296 5391
rect 2454 5380 2460 5381
rect 1974 5379 1980 5380
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 2454 5376 2455 5380
rect 2459 5376 2460 5380
rect 2454 5375 2460 5376
rect 2670 5380 2676 5381
rect 2670 5376 2671 5380
rect 2675 5376 2676 5380
rect 2670 5375 2676 5376
rect 2886 5380 2892 5381
rect 2886 5376 2887 5380
rect 2891 5376 2892 5380
rect 2886 5375 2892 5376
rect 3102 5380 3108 5381
rect 3102 5376 3103 5380
rect 3107 5376 3108 5380
rect 3102 5375 3108 5376
rect 3318 5380 3324 5381
rect 3318 5376 3319 5380
rect 3323 5376 3324 5380
rect 3318 5375 3324 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 1974 5374 1980 5375
rect 3798 5374 3804 5375
rect 3838 5356 3844 5357
rect 5662 5356 5668 5357
rect 3838 5352 3839 5356
rect 3843 5352 3844 5356
rect 3838 5351 3844 5352
rect 3858 5355 3864 5356
rect 3858 5351 3859 5355
rect 3863 5351 3864 5355
rect 3858 5350 3864 5351
rect 4074 5355 4080 5356
rect 4074 5351 4075 5355
rect 4079 5351 4080 5355
rect 4074 5350 4080 5351
rect 4306 5355 4312 5356
rect 4306 5351 4307 5355
rect 4311 5351 4312 5355
rect 4306 5350 4312 5351
rect 4530 5355 4536 5356
rect 4530 5351 4531 5355
rect 4535 5351 4536 5355
rect 4530 5350 4536 5351
rect 4738 5355 4744 5356
rect 4738 5351 4739 5355
rect 4743 5351 4744 5355
rect 4738 5350 4744 5351
rect 4938 5355 4944 5356
rect 4938 5351 4939 5355
rect 4943 5351 4944 5355
rect 4938 5350 4944 5351
rect 5138 5355 5144 5356
rect 5138 5351 5139 5355
rect 5143 5351 5144 5355
rect 5138 5350 5144 5351
rect 5338 5355 5344 5356
rect 5338 5351 5339 5355
rect 5343 5351 5344 5355
rect 5338 5350 5344 5351
rect 5514 5355 5520 5356
rect 5514 5351 5515 5355
rect 5519 5351 5520 5355
rect 5662 5352 5663 5356
rect 5667 5352 5668 5356
rect 5662 5351 5668 5352
rect 5514 5350 5520 5351
rect 3886 5340 3892 5341
rect 3838 5339 3844 5340
rect 3838 5335 3839 5339
rect 3843 5335 3844 5339
rect 3886 5336 3887 5340
rect 3891 5336 3892 5340
rect 3886 5335 3892 5336
rect 4102 5340 4108 5341
rect 4102 5336 4103 5340
rect 4107 5336 4108 5340
rect 4102 5335 4108 5336
rect 4334 5340 4340 5341
rect 4334 5336 4335 5340
rect 4339 5336 4340 5340
rect 4334 5335 4340 5336
rect 4558 5340 4564 5341
rect 4558 5336 4559 5340
rect 4563 5336 4564 5340
rect 4558 5335 4564 5336
rect 4766 5340 4772 5341
rect 4766 5336 4767 5340
rect 4771 5336 4772 5340
rect 4766 5335 4772 5336
rect 4966 5340 4972 5341
rect 4966 5336 4967 5340
rect 4971 5336 4972 5340
rect 4966 5335 4972 5336
rect 5166 5340 5172 5341
rect 5166 5336 5167 5340
rect 5171 5336 5172 5340
rect 5166 5335 5172 5336
rect 5366 5340 5372 5341
rect 5366 5336 5367 5340
rect 5371 5336 5372 5340
rect 5366 5335 5372 5336
rect 5542 5340 5548 5341
rect 5542 5336 5543 5340
rect 5547 5336 5548 5340
rect 5542 5335 5548 5336
rect 5662 5339 5668 5340
rect 5662 5335 5663 5339
rect 5667 5335 5668 5339
rect 3838 5334 3844 5335
rect 5662 5334 5668 5335
rect 1974 5321 1980 5322
rect 3798 5321 3804 5322
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2446 5320 2452 5321
rect 2446 5316 2447 5320
rect 2451 5316 2452 5320
rect 2446 5315 2452 5316
rect 2582 5320 2588 5321
rect 2582 5316 2583 5320
rect 2587 5316 2588 5320
rect 2582 5315 2588 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2854 5320 2860 5321
rect 2854 5316 2855 5320
rect 2859 5316 2860 5320
rect 2854 5315 2860 5316
rect 2990 5320 2996 5321
rect 2990 5316 2991 5320
rect 2995 5316 2996 5320
rect 2990 5315 2996 5316
rect 3134 5320 3140 5321
rect 3134 5316 3135 5320
rect 3139 5316 3140 5320
rect 3134 5315 3140 5316
rect 3286 5320 3292 5321
rect 3286 5316 3287 5320
rect 3291 5316 3292 5320
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3286 5315 3292 5316
rect 2418 5305 2424 5306
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2418 5301 2419 5305
rect 2423 5301 2424 5305
rect 2418 5300 2424 5301
rect 2554 5305 2560 5306
rect 2554 5301 2555 5305
rect 2559 5301 2560 5305
rect 2554 5300 2560 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2826 5305 2832 5306
rect 2826 5301 2827 5305
rect 2831 5301 2832 5305
rect 2826 5300 2832 5301
rect 2962 5305 2968 5306
rect 2962 5301 2963 5305
rect 2967 5301 2968 5305
rect 2962 5300 2968 5301
rect 3106 5305 3112 5306
rect 3106 5301 3107 5305
rect 3111 5301 3112 5305
rect 3106 5300 3112 5301
rect 3258 5305 3264 5306
rect 3258 5301 3259 5305
rect 3263 5301 3264 5305
rect 3258 5300 3264 5301
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 1974 5299 1980 5300
rect 3798 5299 3804 5300
rect 3838 5265 3844 5266
rect 5662 5265 5668 5266
rect 3838 5261 3839 5265
rect 3843 5261 3844 5265
rect 3838 5260 3844 5261
rect 3886 5264 3892 5265
rect 3886 5260 3887 5264
rect 3891 5260 3892 5264
rect 3886 5259 3892 5260
rect 4094 5264 4100 5265
rect 4094 5260 4095 5264
rect 4099 5260 4100 5264
rect 4094 5259 4100 5260
rect 4342 5264 4348 5265
rect 4342 5260 4343 5264
rect 4347 5260 4348 5264
rect 4342 5259 4348 5260
rect 4614 5264 4620 5265
rect 4614 5260 4615 5264
rect 4619 5260 4620 5264
rect 4614 5259 4620 5260
rect 4910 5264 4916 5265
rect 4910 5260 4911 5264
rect 4915 5260 4916 5264
rect 4910 5259 4916 5260
rect 5214 5264 5220 5265
rect 5214 5260 5215 5264
rect 5219 5260 5220 5264
rect 5214 5259 5220 5260
rect 5526 5264 5532 5265
rect 5526 5260 5527 5264
rect 5531 5260 5532 5264
rect 5662 5261 5663 5265
rect 5667 5261 5668 5265
rect 5662 5260 5668 5261
rect 5526 5259 5532 5260
rect 3858 5249 3864 5250
rect 3838 5248 3844 5249
rect 3838 5244 3839 5248
rect 3843 5244 3844 5248
rect 3858 5245 3859 5249
rect 3863 5245 3864 5249
rect 3858 5244 3864 5245
rect 4066 5249 4072 5250
rect 4066 5245 4067 5249
rect 4071 5245 4072 5249
rect 4066 5244 4072 5245
rect 4314 5249 4320 5250
rect 4314 5245 4315 5249
rect 4319 5245 4320 5249
rect 4314 5244 4320 5245
rect 4586 5249 4592 5250
rect 4586 5245 4587 5249
rect 4591 5245 4592 5249
rect 4586 5244 4592 5245
rect 4882 5249 4888 5250
rect 4882 5245 4883 5249
rect 4887 5245 4888 5249
rect 4882 5244 4888 5245
rect 5186 5249 5192 5250
rect 5186 5245 5187 5249
rect 5191 5245 5192 5249
rect 5186 5244 5192 5245
rect 5498 5249 5504 5250
rect 5498 5245 5499 5249
rect 5503 5245 5504 5249
rect 5498 5244 5504 5245
rect 5662 5248 5668 5249
rect 5662 5244 5663 5248
rect 5667 5244 5668 5248
rect 3838 5243 3844 5244
rect 5662 5243 5668 5244
rect 110 5200 116 5201
rect 1934 5200 1940 5201
rect 110 5196 111 5200
rect 115 5196 116 5200
rect 110 5195 116 5196
rect 458 5199 464 5200
rect 458 5195 459 5199
rect 463 5195 464 5199
rect 458 5194 464 5195
rect 594 5199 600 5200
rect 594 5195 595 5199
rect 599 5195 600 5199
rect 594 5194 600 5195
rect 730 5199 736 5200
rect 730 5195 731 5199
rect 735 5195 736 5199
rect 730 5194 736 5195
rect 866 5199 872 5200
rect 866 5195 867 5199
rect 871 5195 872 5199
rect 866 5194 872 5195
rect 1002 5199 1008 5200
rect 1002 5195 1003 5199
rect 1007 5195 1008 5199
rect 1002 5194 1008 5195
rect 1138 5199 1144 5200
rect 1138 5195 1139 5199
rect 1143 5195 1144 5199
rect 1138 5194 1144 5195
rect 1274 5199 1280 5200
rect 1274 5195 1275 5199
rect 1279 5195 1280 5199
rect 1274 5194 1280 5195
rect 1410 5199 1416 5200
rect 1410 5195 1411 5199
rect 1415 5195 1416 5199
rect 1410 5194 1416 5195
rect 1546 5199 1552 5200
rect 1546 5195 1547 5199
rect 1551 5195 1552 5199
rect 1934 5196 1935 5200
rect 1939 5196 1940 5200
rect 1934 5195 1940 5196
rect 1546 5194 1552 5195
rect 486 5184 492 5185
rect 110 5183 116 5184
rect 110 5179 111 5183
rect 115 5179 116 5183
rect 486 5180 487 5184
rect 491 5180 492 5184
rect 486 5179 492 5180
rect 622 5184 628 5185
rect 622 5180 623 5184
rect 627 5180 628 5184
rect 622 5179 628 5180
rect 758 5184 764 5185
rect 758 5180 759 5184
rect 763 5180 764 5184
rect 758 5179 764 5180
rect 894 5184 900 5185
rect 894 5180 895 5184
rect 899 5180 900 5184
rect 894 5179 900 5180
rect 1030 5184 1036 5185
rect 1030 5180 1031 5184
rect 1035 5180 1036 5184
rect 1030 5179 1036 5180
rect 1166 5184 1172 5185
rect 1166 5180 1167 5184
rect 1171 5180 1172 5184
rect 1166 5179 1172 5180
rect 1302 5184 1308 5185
rect 1302 5180 1303 5184
rect 1307 5180 1308 5184
rect 1302 5179 1308 5180
rect 1438 5184 1444 5185
rect 1438 5180 1439 5184
rect 1443 5180 1444 5184
rect 1438 5179 1444 5180
rect 1574 5184 1580 5185
rect 1574 5180 1575 5184
rect 1579 5180 1580 5184
rect 1574 5179 1580 5180
rect 1934 5183 1940 5184
rect 1934 5179 1935 5183
rect 1939 5179 1940 5183
rect 110 5178 116 5179
rect 1934 5178 1940 5179
rect 1974 5172 1980 5173
rect 3798 5172 3804 5173
rect 1974 5168 1975 5172
rect 1979 5168 1980 5172
rect 1974 5167 1980 5168
rect 2098 5171 2104 5172
rect 2098 5167 2099 5171
rect 2103 5167 2104 5171
rect 2098 5166 2104 5167
rect 2234 5171 2240 5172
rect 2234 5167 2235 5171
rect 2239 5167 2240 5171
rect 2234 5166 2240 5167
rect 2378 5171 2384 5172
rect 2378 5167 2379 5171
rect 2383 5167 2384 5171
rect 2378 5166 2384 5167
rect 2530 5171 2536 5172
rect 2530 5167 2531 5171
rect 2535 5167 2536 5171
rect 2530 5166 2536 5167
rect 2698 5171 2704 5172
rect 2698 5167 2699 5171
rect 2703 5167 2704 5171
rect 2698 5166 2704 5167
rect 2882 5171 2888 5172
rect 2882 5167 2883 5171
rect 2887 5167 2888 5171
rect 2882 5166 2888 5167
rect 3066 5171 3072 5172
rect 3066 5167 3067 5171
rect 3071 5167 3072 5171
rect 3066 5166 3072 5167
rect 3258 5171 3264 5172
rect 3258 5167 3259 5171
rect 3263 5167 3264 5171
rect 3798 5168 3799 5172
rect 3803 5168 3804 5172
rect 3798 5167 3804 5168
rect 3258 5166 3264 5167
rect 2126 5156 2132 5157
rect 1974 5155 1980 5156
rect 1974 5151 1975 5155
rect 1979 5151 1980 5155
rect 2126 5152 2127 5156
rect 2131 5152 2132 5156
rect 2126 5151 2132 5152
rect 2262 5156 2268 5157
rect 2262 5152 2263 5156
rect 2267 5152 2268 5156
rect 2262 5151 2268 5152
rect 2406 5156 2412 5157
rect 2406 5152 2407 5156
rect 2411 5152 2412 5156
rect 2406 5151 2412 5152
rect 2558 5156 2564 5157
rect 2558 5152 2559 5156
rect 2563 5152 2564 5156
rect 2558 5151 2564 5152
rect 2726 5156 2732 5157
rect 2726 5152 2727 5156
rect 2731 5152 2732 5156
rect 2726 5151 2732 5152
rect 2910 5156 2916 5157
rect 2910 5152 2911 5156
rect 2915 5152 2916 5156
rect 2910 5151 2916 5152
rect 3094 5156 3100 5157
rect 3094 5152 3095 5156
rect 3099 5152 3100 5156
rect 3094 5151 3100 5152
rect 3286 5156 3292 5157
rect 3286 5152 3287 5156
rect 3291 5152 3292 5156
rect 3286 5151 3292 5152
rect 3798 5155 3804 5156
rect 3798 5151 3799 5155
rect 3803 5151 3804 5155
rect 1974 5150 1980 5151
rect 3798 5150 3804 5151
rect 110 5109 116 5110
rect 1934 5109 1940 5110
rect 110 5105 111 5109
rect 115 5105 116 5109
rect 110 5104 116 5105
rect 318 5108 324 5109
rect 318 5104 319 5108
rect 323 5104 324 5108
rect 318 5103 324 5104
rect 502 5108 508 5109
rect 502 5104 503 5108
rect 507 5104 508 5108
rect 502 5103 508 5104
rect 702 5108 708 5109
rect 702 5104 703 5108
rect 707 5104 708 5108
rect 702 5103 708 5104
rect 918 5108 924 5109
rect 918 5104 919 5108
rect 923 5104 924 5108
rect 918 5103 924 5104
rect 1150 5108 1156 5109
rect 1150 5104 1151 5108
rect 1155 5104 1156 5108
rect 1150 5103 1156 5104
rect 1390 5108 1396 5109
rect 1390 5104 1391 5108
rect 1395 5104 1396 5108
rect 1390 5103 1396 5104
rect 1630 5108 1636 5109
rect 1630 5104 1631 5108
rect 1635 5104 1636 5108
rect 1934 5105 1935 5109
rect 1939 5105 1940 5109
rect 1934 5104 1940 5105
rect 3838 5108 3844 5109
rect 5662 5108 5668 5109
rect 3838 5104 3839 5108
rect 3843 5104 3844 5108
rect 1630 5103 1636 5104
rect 3838 5103 3844 5104
rect 3858 5107 3864 5108
rect 3858 5103 3859 5107
rect 3863 5103 3864 5107
rect 3858 5102 3864 5103
rect 3994 5107 4000 5108
rect 3994 5103 3995 5107
rect 3999 5103 4000 5107
rect 3994 5102 4000 5103
rect 4154 5107 4160 5108
rect 4154 5103 4155 5107
rect 4159 5103 4160 5107
rect 4154 5102 4160 5103
rect 4362 5107 4368 5108
rect 4362 5103 4363 5107
rect 4367 5103 4368 5107
rect 4362 5102 4368 5103
rect 4610 5107 4616 5108
rect 4610 5103 4611 5107
rect 4615 5103 4616 5107
rect 4610 5102 4616 5103
rect 4882 5107 4888 5108
rect 4882 5103 4883 5107
rect 4887 5103 4888 5107
rect 4882 5102 4888 5103
rect 5170 5107 5176 5108
rect 5170 5103 5171 5107
rect 5175 5103 5176 5107
rect 5170 5102 5176 5103
rect 5466 5107 5472 5108
rect 5466 5103 5467 5107
rect 5471 5103 5472 5107
rect 5662 5104 5663 5108
rect 5667 5104 5668 5108
rect 5662 5103 5668 5104
rect 5466 5102 5472 5103
rect 290 5093 296 5094
rect 110 5092 116 5093
rect 110 5088 111 5092
rect 115 5088 116 5092
rect 290 5089 291 5093
rect 295 5089 296 5093
rect 290 5088 296 5089
rect 474 5093 480 5094
rect 474 5089 475 5093
rect 479 5089 480 5093
rect 474 5088 480 5089
rect 674 5093 680 5094
rect 674 5089 675 5093
rect 679 5089 680 5093
rect 674 5088 680 5089
rect 890 5093 896 5094
rect 890 5089 891 5093
rect 895 5089 896 5093
rect 890 5088 896 5089
rect 1122 5093 1128 5094
rect 1122 5089 1123 5093
rect 1127 5089 1128 5093
rect 1122 5088 1128 5089
rect 1362 5093 1368 5094
rect 1362 5089 1363 5093
rect 1367 5089 1368 5093
rect 1362 5088 1368 5089
rect 1602 5093 1608 5094
rect 1602 5089 1603 5093
rect 1607 5089 1608 5093
rect 1602 5088 1608 5089
rect 1934 5092 1940 5093
rect 3886 5092 3892 5093
rect 1934 5088 1935 5092
rect 1939 5088 1940 5092
rect 110 5087 116 5088
rect 1934 5087 1940 5088
rect 3838 5091 3844 5092
rect 3838 5087 3839 5091
rect 3843 5087 3844 5091
rect 3886 5088 3887 5092
rect 3891 5088 3892 5092
rect 3886 5087 3892 5088
rect 4022 5092 4028 5093
rect 4022 5088 4023 5092
rect 4027 5088 4028 5092
rect 4022 5087 4028 5088
rect 4182 5092 4188 5093
rect 4182 5088 4183 5092
rect 4187 5088 4188 5092
rect 4182 5087 4188 5088
rect 4390 5092 4396 5093
rect 4390 5088 4391 5092
rect 4395 5088 4396 5092
rect 4390 5087 4396 5088
rect 4638 5092 4644 5093
rect 4638 5088 4639 5092
rect 4643 5088 4644 5092
rect 4638 5087 4644 5088
rect 4910 5092 4916 5093
rect 4910 5088 4911 5092
rect 4915 5088 4916 5092
rect 4910 5087 4916 5088
rect 5198 5092 5204 5093
rect 5198 5088 5199 5092
rect 5203 5088 5204 5092
rect 5198 5087 5204 5088
rect 5494 5092 5500 5093
rect 5494 5088 5495 5092
rect 5499 5088 5500 5092
rect 5494 5087 5500 5088
rect 5662 5091 5668 5092
rect 5662 5087 5663 5091
rect 5667 5087 5668 5091
rect 3838 5086 3844 5087
rect 5662 5086 5668 5087
rect 1974 5073 1980 5074
rect 3798 5073 3804 5074
rect 1974 5069 1975 5073
rect 1979 5069 1980 5073
rect 1974 5068 1980 5069
rect 2078 5072 2084 5073
rect 2078 5068 2079 5072
rect 2083 5068 2084 5072
rect 2078 5067 2084 5068
rect 2358 5072 2364 5073
rect 2358 5068 2359 5072
rect 2363 5068 2364 5072
rect 2358 5067 2364 5068
rect 2638 5072 2644 5073
rect 2638 5068 2639 5072
rect 2643 5068 2644 5072
rect 2638 5067 2644 5068
rect 2910 5072 2916 5073
rect 2910 5068 2911 5072
rect 2915 5068 2916 5072
rect 2910 5067 2916 5068
rect 3174 5072 3180 5073
rect 3174 5068 3175 5072
rect 3179 5068 3180 5072
rect 3174 5067 3180 5068
rect 3438 5072 3444 5073
rect 3438 5068 3439 5072
rect 3443 5068 3444 5072
rect 3438 5067 3444 5068
rect 3678 5072 3684 5073
rect 3678 5068 3679 5072
rect 3683 5068 3684 5072
rect 3798 5069 3799 5073
rect 3803 5069 3804 5073
rect 3798 5068 3804 5069
rect 3678 5067 3684 5068
rect 2050 5057 2056 5058
rect 1974 5056 1980 5057
rect 1974 5052 1975 5056
rect 1979 5052 1980 5056
rect 2050 5053 2051 5057
rect 2055 5053 2056 5057
rect 2050 5052 2056 5053
rect 2330 5057 2336 5058
rect 2330 5053 2331 5057
rect 2335 5053 2336 5057
rect 2330 5052 2336 5053
rect 2610 5057 2616 5058
rect 2610 5053 2611 5057
rect 2615 5053 2616 5057
rect 2610 5052 2616 5053
rect 2882 5057 2888 5058
rect 2882 5053 2883 5057
rect 2887 5053 2888 5057
rect 2882 5052 2888 5053
rect 3146 5057 3152 5058
rect 3146 5053 3147 5057
rect 3151 5053 3152 5057
rect 3146 5052 3152 5053
rect 3410 5057 3416 5058
rect 3410 5053 3411 5057
rect 3415 5053 3416 5057
rect 3410 5052 3416 5053
rect 3650 5057 3656 5058
rect 3650 5053 3651 5057
rect 3655 5053 3656 5057
rect 3650 5052 3656 5053
rect 3798 5056 3804 5057
rect 3798 5052 3799 5056
rect 3803 5052 3804 5056
rect 1974 5051 1980 5052
rect 3798 5051 3804 5052
rect 3838 5017 3844 5018
rect 5662 5017 5668 5018
rect 3838 5013 3839 5017
rect 3843 5013 3844 5017
rect 3838 5012 3844 5013
rect 4446 5016 4452 5017
rect 4446 5012 4447 5016
rect 4451 5012 4452 5016
rect 4446 5011 4452 5012
rect 4630 5016 4636 5017
rect 4630 5012 4631 5016
rect 4635 5012 4636 5016
rect 4630 5011 4636 5012
rect 4830 5016 4836 5017
rect 4830 5012 4831 5016
rect 4835 5012 4836 5016
rect 4830 5011 4836 5012
rect 5046 5016 5052 5017
rect 5046 5012 5047 5016
rect 5051 5012 5052 5016
rect 5046 5011 5052 5012
rect 5278 5016 5284 5017
rect 5278 5012 5279 5016
rect 5283 5012 5284 5016
rect 5278 5011 5284 5012
rect 5510 5016 5516 5017
rect 5510 5012 5511 5016
rect 5515 5012 5516 5016
rect 5662 5013 5663 5017
rect 5667 5013 5668 5017
rect 5662 5012 5668 5013
rect 5510 5011 5516 5012
rect 4418 5001 4424 5002
rect 3838 5000 3844 5001
rect 3838 4996 3839 5000
rect 3843 4996 3844 5000
rect 4418 4997 4419 5001
rect 4423 4997 4424 5001
rect 4418 4996 4424 4997
rect 4602 5001 4608 5002
rect 4602 4997 4603 5001
rect 4607 4997 4608 5001
rect 4602 4996 4608 4997
rect 4802 5001 4808 5002
rect 4802 4997 4803 5001
rect 4807 4997 4808 5001
rect 4802 4996 4808 4997
rect 5018 5001 5024 5002
rect 5018 4997 5019 5001
rect 5023 4997 5024 5001
rect 5018 4996 5024 4997
rect 5250 5001 5256 5002
rect 5250 4997 5251 5001
rect 5255 4997 5256 5001
rect 5250 4996 5256 4997
rect 5482 5001 5488 5002
rect 5482 4997 5483 5001
rect 5487 4997 5488 5001
rect 5482 4996 5488 4997
rect 5662 5000 5668 5001
rect 5662 4996 5663 5000
rect 5667 4996 5668 5000
rect 3838 4995 3844 4996
rect 5662 4995 5668 4996
rect 110 4960 116 4961
rect 1934 4960 1940 4961
rect 110 4956 111 4960
rect 115 4956 116 4960
rect 110 4955 116 4956
rect 138 4959 144 4960
rect 138 4955 139 4959
rect 143 4955 144 4959
rect 138 4954 144 4955
rect 410 4959 416 4960
rect 410 4955 411 4959
rect 415 4955 416 4959
rect 410 4954 416 4955
rect 682 4959 688 4960
rect 682 4955 683 4959
rect 687 4955 688 4959
rect 682 4954 688 4955
rect 962 4959 968 4960
rect 962 4955 963 4959
rect 967 4955 968 4959
rect 962 4954 968 4955
rect 1242 4959 1248 4960
rect 1242 4955 1243 4959
rect 1247 4955 1248 4959
rect 1242 4954 1248 4955
rect 1522 4959 1528 4960
rect 1522 4955 1523 4959
rect 1527 4955 1528 4959
rect 1522 4954 1528 4955
rect 1786 4959 1792 4960
rect 1786 4955 1787 4959
rect 1791 4955 1792 4959
rect 1934 4956 1935 4960
rect 1939 4956 1940 4960
rect 1934 4955 1940 4956
rect 1786 4954 1792 4955
rect 166 4944 172 4945
rect 110 4943 116 4944
rect 110 4939 111 4943
rect 115 4939 116 4943
rect 166 4940 167 4944
rect 171 4940 172 4944
rect 166 4939 172 4940
rect 438 4944 444 4945
rect 438 4940 439 4944
rect 443 4940 444 4944
rect 438 4939 444 4940
rect 710 4944 716 4945
rect 710 4940 711 4944
rect 715 4940 716 4944
rect 710 4939 716 4940
rect 990 4944 996 4945
rect 990 4940 991 4944
rect 995 4940 996 4944
rect 990 4939 996 4940
rect 1270 4944 1276 4945
rect 1270 4940 1271 4944
rect 1275 4940 1276 4944
rect 1270 4939 1276 4940
rect 1550 4944 1556 4945
rect 1550 4940 1551 4944
rect 1555 4940 1556 4944
rect 1550 4939 1556 4940
rect 1814 4944 1820 4945
rect 1814 4940 1815 4944
rect 1819 4940 1820 4944
rect 1814 4939 1820 4940
rect 1934 4943 1940 4944
rect 1934 4939 1935 4943
rect 1939 4939 1940 4943
rect 110 4938 116 4939
rect 1934 4938 1940 4939
rect 1974 4904 1980 4905
rect 3798 4904 3804 4905
rect 1974 4900 1975 4904
rect 1979 4900 1980 4904
rect 1974 4899 1980 4900
rect 1994 4903 2000 4904
rect 1994 4899 1995 4903
rect 1999 4899 2000 4903
rect 1994 4898 2000 4899
rect 2130 4903 2136 4904
rect 2130 4899 2131 4903
rect 2135 4899 2136 4903
rect 2130 4898 2136 4899
rect 2298 4903 2304 4904
rect 2298 4899 2299 4903
rect 2303 4899 2304 4903
rect 2298 4898 2304 4899
rect 2466 4903 2472 4904
rect 2466 4899 2467 4903
rect 2471 4899 2472 4903
rect 2466 4898 2472 4899
rect 2642 4903 2648 4904
rect 2642 4899 2643 4903
rect 2647 4899 2648 4903
rect 2642 4898 2648 4899
rect 2818 4903 2824 4904
rect 2818 4899 2819 4903
rect 2823 4899 2824 4903
rect 2818 4898 2824 4899
rect 2986 4903 2992 4904
rect 2986 4899 2987 4903
rect 2991 4899 2992 4903
rect 2986 4898 2992 4899
rect 3154 4903 3160 4904
rect 3154 4899 3155 4903
rect 3159 4899 3160 4903
rect 3154 4898 3160 4899
rect 3322 4903 3328 4904
rect 3322 4899 3323 4903
rect 3327 4899 3328 4903
rect 3322 4898 3328 4899
rect 3498 4903 3504 4904
rect 3498 4899 3499 4903
rect 3503 4899 3504 4903
rect 3498 4898 3504 4899
rect 3650 4903 3656 4904
rect 3650 4899 3651 4903
rect 3655 4899 3656 4903
rect 3798 4900 3799 4904
rect 3803 4900 3804 4904
rect 3798 4899 3804 4900
rect 3650 4898 3656 4899
rect 2022 4888 2028 4889
rect 1974 4887 1980 4888
rect 110 4885 116 4886
rect 1934 4885 1940 4886
rect 110 4881 111 4885
rect 115 4881 116 4885
rect 110 4880 116 4881
rect 158 4884 164 4885
rect 158 4880 159 4884
rect 163 4880 164 4884
rect 158 4879 164 4880
rect 414 4884 420 4885
rect 414 4880 415 4884
rect 419 4880 420 4884
rect 414 4879 420 4880
rect 734 4884 740 4885
rect 734 4880 735 4884
rect 739 4880 740 4884
rect 734 4879 740 4880
rect 1086 4884 1092 4885
rect 1086 4880 1087 4884
rect 1091 4880 1092 4884
rect 1086 4879 1092 4880
rect 1462 4884 1468 4885
rect 1462 4880 1463 4884
rect 1467 4880 1468 4884
rect 1462 4879 1468 4880
rect 1814 4884 1820 4885
rect 1814 4880 1815 4884
rect 1819 4880 1820 4884
rect 1934 4881 1935 4885
rect 1939 4881 1940 4885
rect 1974 4883 1975 4887
rect 1979 4883 1980 4887
rect 2022 4884 2023 4888
rect 2027 4884 2028 4888
rect 2022 4883 2028 4884
rect 2158 4888 2164 4889
rect 2158 4884 2159 4888
rect 2163 4884 2164 4888
rect 2158 4883 2164 4884
rect 2326 4888 2332 4889
rect 2326 4884 2327 4888
rect 2331 4884 2332 4888
rect 2326 4883 2332 4884
rect 2494 4888 2500 4889
rect 2494 4884 2495 4888
rect 2499 4884 2500 4888
rect 2494 4883 2500 4884
rect 2670 4888 2676 4889
rect 2670 4884 2671 4888
rect 2675 4884 2676 4888
rect 2670 4883 2676 4884
rect 2846 4888 2852 4889
rect 2846 4884 2847 4888
rect 2851 4884 2852 4888
rect 2846 4883 2852 4884
rect 3014 4888 3020 4889
rect 3014 4884 3015 4888
rect 3019 4884 3020 4888
rect 3014 4883 3020 4884
rect 3182 4888 3188 4889
rect 3182 4884 3183 4888
rect 3187 4884 3188 4888
rect 3182 4883 3188 4884
rect 3350 4888 3356 4889
rect 3350 4884 3351 4888
rect 3355 4884 3356 4888
rect 3350 4883 3356 4884
rect 3526 4888 3532 4889
rect 3526 4884 3527 4888
rect 3531 4884 3532 4888
rect 3526 4883 3532 4884
rect 3678 4888 3684 4889
rect 3678 4884 3679 4888
rect 3683 4884 3684 4888
rect 3678 4883 3684 4884
rect 3798 4887 3804 4888
rect 3798 4883 3799 4887
rect 3803 4883 3804 4887
rect 1974 4882 1980 4883
rect 3798 4882 3804 4883
rect 1934 4880 1940 4881
rect 1814 4879 1820 4880
rect 130 4869 136 4870
rect 110 4868 116 4869
rect 110 4864 111 4868
rect 115 4864 116 4868
rect 130 4865 131 4869
rect 135 4865 136 4869
rect 130 4864 136 4865
rect 386 4869 392 4870
rect 386 4865 387 4869
rect 391 4865 392 4869
rect 386 4864 392 4865
rect 706 4869 712 4870
rect 706 4865 707 4869
rect 711 4865 712 4869
rect 706 4864 712 4865
rect 1058 4869 1064 4870
rect 1058 4865 1059 4869
rect 1063 4865 1064 4869
rect 1058 4864 1064 4865
rect 1434 4869 1440 4870
rect 1434 4865 1435 4869
rect 1439 4865 1440 4869
rect 1434 4864 1440 4865
rect 1786 4869 1792 4870
rect 1786 4865 1787 4869
rect 1791 4865 1792 4869
rect 1786 4864 1792 4865
rect 1934 4868 1940 4869
rect 1934 4864 1935 4868
rect 1939 4864 1940 4868
rect 110 4863 116 4864
rect 1934 4863 1940 4864
rect 3838 4852 3844 4853
rect 5662 4852 5668 4853
rect 3838 4848 3839 4852
rect 3843 4848 3844 4852
rect 3838 4847 3844 4848
rect 4674 4851 4680 4852
rect 4674 4847 4675 4851
rect 4679 4847 4680 4851
rect 4674 4846 4680 4847
rect 4826 4851 4832 4852
rect 4826 4847 4827 4851
rect 4831 4847 4832 4851
rect 4826 4846 4832 4847
rect 4986 4851 4992 4852
rect 4986 4847 4987 4851
rect 4991 4847 4992 4851
rect 4986 4846 4992 4847
rect 5154 4851 5160 4852
rect 5154 4847 5155 4851
rect 5159 4847 5160 4851
rect 5154 4846 5160 4847
rect 5322 4851 5328 4852
rect 5322 4847 5323 4851
rect 5327 4847 5328 4851
rect 5322 4846 5328 4847
rect 5498 4851 5504 4852
rect 5498 4847 5499 4851
rect 5503 4847 5504 4851
rect 5662 4848 5663 4852
rect 5667 4848 5668 4852
rect 5662 4847 5668 4848
rect 5498 4846 5504 4847
rect 4702 4836 4708 4837
rect 3838 4835 3844 4836
rect 3838 4831 3839 4835
rect 3843 4831 3844 4835
rect 4702 4832 4703 4836
rect 4707 4832 4708 4836
rect 4702 4831 4708 4832
rect 4854 4836 4860 4837
rect 4854 4832 4855 4836
rect 4859 4832 4860 4836
rect 4854 4831 4860 4832
rect 5014 4836 5020 4837
rect 5014 4832 5015 4836
rect 5019 4832 5020 4836
rect 5014 4831 5020 4832
rect 5182 4836 5188 4837
rect 5182 4832 5183 4836
rect 5187 4832 5188 4836
rect 5182 4831 5188 4832
rect 5350 4836 5356 4837
rect 5350 4832 5351 4836
rect 5355 4832 5356 4836
rect 5350 4831 5356 4832
rect 5526 4836 5532 4837
rect 5526 4832 5527 4836
rect 5531 4832 5532 4836
rect 5526 4831 5532 4832
rect 5662 4835 5668 4836
rect 5662 4831 5663 4835
rect 5667 4831 5668 4835
rect 3838 4830 3844 4831
rect 5662 4830 5668 4831
rect 1974 4801 1980 4802
rect 3798 4801 3804 4802
rect 1974 4797 1975 4801
rect 1979 4797 1980 4801
rect 1974 4796 1980 4797
rect 2390 4800 2396 4801
rect 2390 4796 2391 4800
rect 2395 4796 2396 4800
rect 2390 4795 2396 4796
rect 2526 4800 2532 4801
rect 2526 4796 2527 4800
rect 2531 4796 2532 4800
rect 2526 4795 2532 4796
rect 2662 4800 2668 4801
rect 2662 4796 2663 4800
rect 2667 4796 2668 4800
rect 2662 4795 2668 4796
rect 2806 4800 2812 4801
rect 2806 4796 2807 4800
rect 2811 4796 2812 4800
rect 2806 4795 2812 4796
rect 2950 4800 2956 4801
rect 2950 4796 2951 4800
rect 2955 4796 2956 4800
rect 2950 4795 2956 4796
rect 3094 4800 3100 4801
rect 3094 4796 3095 4800
rect 3099 4796 3100 4800
rect 3094 4795 3100 4796
rect 3238 4800 3244 4801
rect 3238 4796 3239 4800
rect 3243 4796 3244 4800
rect 3238 4795 3244 4796
rect 3382 4800 3388 4801
rect 3382 4796 3383 4800
rect 3387 4796 3388 4800
rect 3382 4795 3388 4796
rect 3526 4800 3532 4801
rect 3526 4796 3527 4800
rect 3531 4796 3532 4800
rect 3798 4797 3799 4801
rect 3803 4797 3804 4801
rect 3798 4796 3804 4797
rect 3526 4795 3532 4796
rect 2362 4785 2368 4786
rect 1974 4784 1980 4785
rect 1974 4780 1975 4784
rect 1979 4780 1980 4784
rect 2362 4781 2363 4785
rect 2367 4781 2368 4785
rect 2362 4780 2368 4781
rect 2498 4785 2504 4786
rect 2498 4781 2499 4785
rect 2503 4781 2504 4785
rect 2498 4780 2504 4781
rect 2634 4785 2640 4786
rect 2634 4781 2635 4785
rect 2639 4781 2640 4785
rect 2634 4780 2640 4781
rect 2778 4785 2784 4786
rect 2778 4781 2779 4785
rect 2783 4781 2784 4785
rect 2778 4780 2784 4781
rect 2922 4785 2928 4786
rect 2922 4781 2923 4785
rect 2927 4781 2928 4785
rect 2922 4780 2928 4781
rect 3066 4785 3072 4786
rect 3066 4781 3067 4785
rect 3071 4781 3072 4785
rect 3066 4780 3072 4781
rect 3210 4785 3216 4786
rect 3210 4781 3211 4785
rect 3215 4781 3216 4785
rect 3210 4780 3216 4781
rect 3354 4785 3360 4786
rect 3354 4781 3355 4785
rect 3359 4781 3360 4785
rect 3354 4780 3360 4781
rect 3498 4785 3504 4786
rect 3498 4781 3499 4785
rect 3503 4781 3504 4785
rect 3498 4780 3504 4781
rect 3798 4784 3804 4785
rect 3798 4780 3799 4784
rect 3803 4780 3804 4784
rect 1974 4779 1980 4780
rect 3798 4779 3804 4780
rect 3838 4757 3844 4758
rect 5662 4757 5668 4758
rect 3838 4753 3839 4757
rect 3843 4753 3844 4757
rect 3838 4752 3844 4753
rect 4854 4756 4860 4757
rect 4854 4752 4855 4756
rect 4859 4752 4860 4756
rect 4854 4751 4860 4752
rect 4990 4756 4996 4757
rect 4990 4752 4991 4756
rect 4995 4752 4996 4756
rect 4990 4751 4996 4752
rect 5126 4756 5132 4757
rect 5126 4752 5127 4756
rect 5131 4752 5132 4756
rect 5126 4751 5132 4752
rect 5262 4756 5268 4757
rect 5262 4752 5263 4756
rect 5267 4752 5268 4756
rect 5262 4751 5268 4752
rect 5398 4756 5404 4757
rect 5398 4752 5399 4756
rect 5403 4752 5404 4756
rect 5398 4751 5404 4752
rect 5534 4756 5540 4757
rect 5534 4752 5535 4756
rect 5539 4752 5540 4756
rect 5662 4753 5663 4757
rect 5667 4753 5668 4757
rect 5662 4752 5668 4753
rect 5534 4751 5540 4752
rect 4826 4741 4832 4742
rect 3838 4740 3844 4741
rect 3838 4736 3839 4740
rect 3843 4736 3844 4740
rect 4826 4737 4827 4741
rect 4831 4737 4832 4741
rect 4826 4736 4832 4737
rect 4962 4741 4968 4742
rect 4962 4737 4963 4741
rect 4967 4737 4968 4741
rect 4962 4736 4968 4737
rect 5098 4741 5104 4742
rect 5098 4737 5099 4741
rect 5103 4737 5104 4741
rect 5098 4736 5104 4737
rect 5234 4741 5240 4742
rect 5234 4737 5235 4741
rect 5239 4737 5240 4741
rect 5234 4736 5240 4737
rect 5370 4741 5376 4742
rect 5370 4737 5371 4741
rect 5375 4737 5376 4741
rect 5370 4736 5376 4737
rect 5506 4741 5512 4742
rect 5506 4737 5507 4741
rect 5511 4737 5512 4741
rect 5506 4736 5512 4737
rect 5662 4740 5668 4741
rect 5662 4736 5663 4740
rect 5667 4736 5668 4740
rect 3838 4735 3844 4736
rect 5662 4735 5668 4736
rect 110 4724 116 4725
rect 1934 4724 1940 4725
rect 110 4720 111 4724
rect 115 4720 116 4724
rect 110 4719 116 4720
rect 130 4723 136 4724
rect 130 4719 131 4723
rect 135 4719 136 4723
rect 130 4718 136 4719
rect 266 4723 272 4724
rect 266 4719 267 4723
rect 271 4719 272 4723
rect 266 4718 272 4719
rect 402 4723 408 4724
rect 402 4719 403 4723
rect 407 4719 408 4723
rect 402 4718 408 4719
rect 538 4723 544 4724
rect 538 4719 539 4723
rect 543 4719 544 4723
rect 538 4718 544 4719
rect 674 4723 680 4724
rect 674 4719 675 4723
rect 679 4719 680 4723
rect 1934 4720 1935 4724
rect 1939 4720 1940 4724
rect 1934 4719 1940 4720
rect 674 4718 680 4719
rect 158 4708 164 4709
rect 110 4707 116 4708
rect 110 4703 111 4707
rect 115 4703 116 4707
rect 158 4704 159 4708
rect 163 4704 164 4708
rect 158 4703 164 4704
rect 294 4708 300 4709
rect 294 4704 295 4708
rect 299 4704 300 4708
rect 294 4703 300 4704
rect 430 4708 436 4709
rect 430 4704 431 4708
rect 435 4704 436 4708
rect 430 4703 436 4704
rect 566 4708 572 4709
rect 566 4704 567 4708
rect 571 4704 572 4708
rect 566 4703 572 4704
rect 702 4708 708 4709
rect 702 4704 703 4708
rect 707 4704 708 4708
rect 702 4703 708 4704
rect 1934 4707 1940 4708
rect 1934 4703 1935 4707
rect 1939 4703 1940 4707
rect 110 4702 116 4703
rect 1934 4702 1940 4703
rect 110 4645 116 4646
rect 1934 4645 1940 4646
rect 110 4641 111 4645
rect 115 4641 116 4645
rect 110 4640 116 4641
rect 158 4644 164 4645
rect 158 4640 159 4644
rect 163 4640 164 4644
rect 158 4639 164 4640
rect 294 4644 300 4645
rect 294 4640 295 4644
rect 299 4640 300 4644
rect 294 4639 300 4640
rect 430 4644 436 4645
rect 430 4640 431 4644
rect 435 4640 436 4644
rect 430 4639 436 4640
rect 566 4644 572 4645
rect 566 4640 567 4644
rect 571 4640 572 4644
rect 566 4639 572 4640
rect 702 4644 708 4645
rect 702 4640 703 4644
rect 707 4640 708 4644
rect 1934 4641 1935 4645
rect 1939 4641 1940 4645
rect 1934 4640 1940 4641
rect 1974 4644 1980 4645
rect 3798 4644 3804 4645
rect 1974 4640 1975 4644
rect 1979 4640 1980 4644
rect 702 4639 708 4640
rect 1974 4639 1980 4640
rect 1994 4643 2000 4644
rect 1994 4639 1995 4643
rect 1999 4639 2000 4643
rect 1994 4638 2000 4639
rect 2130 4643 2136 4644
rect 2130 4639 2131 4643
rect 2135 4639 2136 4643
rect 2130 4638 2136 4639
rect 2266 4643 2272 4644
rect 2266 4639 2267 4643
rect 2271 4639 2272 4643
rect 2266 4638 2272 4639
rect 2426 4643 2432 4644
rect 2426 4639 2427 4643
rect 2431 4639 2432 4643
rect 2426 4638 2432 4639
rect 2586 4643 2592 4644
rect 2586 4639 2587 4643
rect 2591 4639 2592 4643
rect 2586 4638 2592 4639
rect 2746 4643 2752 4644
rect 2746 4639 2747 4643
rect 2751 4639 2752 4643
rect 2746 4638 2752 4639
rect 2906 4643 2912 4644
rect 2906 4639 2907 4643
rect 2911 4639 2912 4643
rect 2906 4638 2912 4639
rect 3066 4643 3072 4644
rect 3066 4639 3067 4643
rect 3071 4639 3072 4643
rect 3066 4638 3072 4639
rect 3234 4643 3240 4644
rect 3234 4639 3235 4643
rect 3239 4639 3240 4643
rect 3798 4640 3799 4644
rect 3803 4640 3804 4644
rect 3798 4639 3804 4640
rect 3234 4638 3240 4639
rect 130 4629 136 4630
rect 110 4628 116 4629
rect 110 4624 111 4628
rect 115 4624 116 4628
rect 130 4625 131 4629
rect 135 4625 136 4629
rect 130 4624 136 4625
rect 266 4629 272 4630
rect 266 4625 267 4629
rect 271 4625 272 4629
rect 266 4624 272 4625
rect 402 4629 408 4630
rect 402 4625 403 4629
rect 407 4625 408 4629
rect 402 4624 408 4625
rect 538 4629 544 4630
rect 538 4625 539 4629
rect 543 4625 544 4629
rect 538 4624 544 4625
rect 674 4629 680 4630
rect 674 4625 675 4629
rect 679 4625 680 4629
rect 674 4624 680 4625
rect 1934 4628 1940 4629
rect 2022 4628 2028 4629
rect 1934 4624 1935 4628
rect 1939 4624 1940 4628
rect 110 4623 116 4624
rect 1934 4623 1940 4624
rect 1974 4627 1980 4628
rect 1974 4623 1975 4627
rect 1979 4623 1980 4627
rect 2022 4624 2023 4628
rect 2027 4624 2028 4628
rect 2022 4623 2028 4624
rect 2158 4628 2164 4629
rect 2158 4624 2159 4628
rect 2163 4624 2164 4628
rect 2158 4623 2164 4624
rect 2294 4628 2300 4629
rect 2294 4624 2295 4628
rect 2299 4624 2300 4628
rect 2294 4623 2300 4624
rect 2454 4628 2460 4629
rect 2454 4624 2455 4628
rect 2459 4624 2460 4628
rect 2454 4623 2460 4624
rect 2614 4628 2620 4629
rect 2614 4624 2615 4628
rect 2619 4624 2620 4628
rect 2614 4623 2620 4624
rect 2774 4628 2780 4629
rect 2774 4624 2775 4628
rect 2779 4624 2780 4628
rect 2774 4623 2780 4624
rect 2934 4628 2940 4629
rect 2934 4624 2935 4628
rect 2939 4624 2940 4628
rect 2934 4623 2940 4624
rect 3094 4628 3100 4629
rect 3094 4624 3095 4628
rect 3099 4624 3100 4628
rect 3094 4623 3100 4624
rect 3262 4628 3268 4629
rect 3262 4624 3263 4628
rect 3267 4624 3268 4628
rect 3262 4623 3268 4624
rect 3798 4627 3804 4628
rect 3798 4623 3799 4627
rect 3803 4623 3804 4627
rect 1974 4622 1980 4623
rect 3798 4622 3804 4623
rect 3838 4588 3844 4589
rect 5662 4588 5668 4589
rect 3838 4584 3839 4588
rect 3843 4584 3844 4588
rect 3838 4583 3844 4584
rect 4714 4587 4720 4588
rect 4714 4583 4715 4587
rect 4719 4583 4720 4587
rect 4714 4582 4720 4583
rect 4858 4587 4864 4588
rect 4858 4583 4859 4587
rect 4863 4583 4864 4587
rect 4858 4582 4864 4583
rect 5010 4587 5016 4588
rect 5010 4583 5011 4587
rect 5015 4583 5016 4587
rect 5010 4582 5016 4583
rect 5170 4587 5176 4588
rect 5170 4583 5171 4587
rect 5175 4583 5176 4587
rect 5170 4582 5176 4583
rect 5338 4587 5344 4588
rect 5338 4583 5339 4587
rect 5343 4583 5344 4587
rect 5338 4582 5344 4583
rect 5514 4587 5520 4588
rect 5514 4583 5515 4587
rect 5519 4583 5520 4587
rect 5662 4584 5663 4588
rect 5667 4584 5668 4588
rect 5662 4583 5668 4584
rect 5514 4582 5520 4583
rect 4742 4572 4748 4573
rect 3838 4571 3844 4572
rect 1974 4569 1980 4570
rect 3798 4569 3804 4570
rect 1974 4565 1975 4569
rect 1979 4565 1980 4569
rect 1974 4564 1980 4565
rect 2022 4568 2028 4569
rect 2022 4564 2023 4568
rect 2027 4564 2028 4568
rect 2022 4563 2028 4564
rect 2174 4568 2180 4569
rect 2174 4564 2175 4568
rect 2179 4564 2180 4568
rect 2174 4563 2180 4564
rect 2350 4568 2356 4569
rect 2350 4564 2351 4568
rect 2355 4564 2356 4568
rect 2350 4563 2356 4564
rect 2526 4568 2532 4569
rect 2526 4564 2527 4568
rect 2531 4564 2532 4568
rect 2526 4563 2532 4564
rect 2694 4568 2700 4569
rect 2694 4564 2695 4568
rect 2699 4564 2700 4568
rect 2694 4563 2700 4564
rect 2870 4568 2876 4569
rect 2870 4564 2871 4568
rect 2875 4564 2876 4568
rect 2870 4563 2876 4564
rect 3046 4568 3052 4569
rect 3046 4564 3047 4568
rect 3051 4564 3052 4568
rect 3798 4565 3799 4569
rect 3803 4565 3804 4569
rect 3838 4567 3839 4571
rect 3843 4567 3844 4571
rect 4742 4568 4743 4572
rect 4747 4568 4748 4572
rect 4742 4567 4748 4568
rect 4886 4572 4892 4573
rect 4886 4568 4887 4572
rect 4891 4568 4892 4572
rect 4886 4567 4892 4568
rect 5038 4572 5044 4573
rect 5038 4568 5039 4572
rect 5043 4568 5044 4572
rect 5038 4567 5044 4568
rect 5198 4572 5204 4573
rect 5198 4568 5199 4572
rect 5203 4568 5204 4572
rect 5198 4567 5204 4568
rect 5366 4572 5372 4573
rect 5366 4568 5367 4572
rect 5371 4568 5372 4572
rect 5366 4567 5372 4568
rect 5542 4572 5548 4573
rect 5542 4568 5543 4572
rect 5547 4568 5548 4572
rect 5542 4567 5548 4568
rect 5662 4571 5668 4572
rect 5662 4567 5663 4571
rect 5667 4567 5668 4571
rect 3838 4566 3844 4567
rect 5662 4566 5668 4567
rect 3798 4564 3804 4565
rect 3046 4563 3052 4564
rect 1994 4553 2000 4554
rect 1974 4552 1980 4553
rect 1974 4548 1975 4552
rect 1979 4548 1980 4552
rect 1994 4549 1995 4553
rect 1999 4549 2000 4553
rect 1994 4548 2000 4549
rect 2146 4553 2152 4554
rect 2146 4549 2147 4553
rect 2151 4549 2152 4553
rect 2146 4548 2152 4549
rect 2322 4553 2328 4554
rect 2322 4549 2323 4553
rect 2327 4549 2328 4553
rect 2322 4548 2328 4549
rect 2498 4553 2504 4554
rect 2498 4549 2499 4553
rect 2503 4549 2504 4553
rect 2498 4548 2504 4549
rect 2666 4553 2672 4554
rect 2666 4549 2667 4553
rect 2671 4549 2672 4553
rect 2666 4548 2672 4549
rect 2842 4553 2848 4554
rect 2842 4549 2843 4553
rect 2847 4549 2848 4553
rect 2842 4548 2848 4549
rect 3018 4553 3024 4554
rect 3018 4549 3019 4553
rect 3023 4549 3024 4553
rect 3018 4548 3024 4549
rect 3798 4552 3804 4553
rect 3798 4548 3799 4552
rect 3803 4548 3804 4552
rect 1974 4547 1980 4548
rect 3798 4547 3804 4548
rect 3838 4489 3844 4490
rect 5662 4489 5668 4490
rect 3838 4485 3839 4489
rect 3843 4485 3844 4489
rect 110 4484 116 4485
rect 1934 4484 1940 4485
rect 3838 4484 3844 4485
rect 3886 4488 3892 4489
rect 3886 4484 3887 4488
rect 3891 4484 3892 4488
rect 110 4480 111 4484
rect 115 4480 116 4484
rect 110 4479 116 4480
rect 298 4483 304 4484
rect 298 4479 299 4483
rect 303 4479 304 4483
rect 298 4478 304 4479
rect 490 4483 496 4484
rect 490 4479 491 4483
rect 495 4479 496 4483
rect 490 4478 496 4479
rect 690 4483 696 4484
rect 690 4479 691 4483
rect 695 4479 696 4483
rect 690 4478 696 4479
rect 906 4483 912 4484
rect 906 4479 907 4483
rect 911 4479 912 4483
rect 906 4478 912 4479
rect 1122 4483 1128 4484
rect 1122 4479 1123 4483
rect 1127 4479 1128 4483
rect 1122 4478 1128 4479
rect 1346 4483 1352 4484
rect 1346 4479 1347 4483
rect 1351 4479 1352 4483
rect 1346 4478 1352 4479
rect 1578 4483 1584 4484
rect 1578 4479 1579 4483
rect 1583 4479 1584 4483
rect 1578 4478 1584 4479
rect 1786 4483 1792 4484
rect 1786 4479 1787 4483
rect 1791 4479 1792 4483
rect 1934 4480 1935 4484
rect 1939 4480 1940 4484
rect 3886 4483 3892 4484
rect 4062 4488 4068 4489
rect 4062 4484 4063 4488
rect 4067 4484 4068 4488
rect 4062 4483 4068 4484
rect 4278 4488 4284 4489
rect 4278 4484 4279 4488
rect 4283 4484 4284 4488
rect 4278 4483 4284 4484
rect 4502 4488 4508 4489
rect 4502 4484 4503 4488
rect 4507 4484 4508 4488
rect 4502 4483 4508 4484
rect 4750 4488 4756 4489
rect 4750 4484 4751 4488
rect 4755 4484 4756 4488
rect 4750 4483 4756 4484
rect 5006 4488 5012 4489
rect 5006 4484 5007 4488
rect 5011 4484 5012 4488
rect 5006 4483 5012 4484
rect 5270 4488 5276 4489
rect 5270 4484 5271 4488
rect 5275 4484 5276 4488
rect 5270 4483 5276 4484
rect 5542 4488 5548 4489
rect 5542 4484 5543 4488
rect 5547 4484 5548 4488
rect 5662 4485 5663 4489
rect 5667 4485 5668 4489
rect 5662 4484 5668 4485
rect 5542 4483 5548 4484
rect 1934 4479 1940 4480
rect 1786 4478 1792 4479
rect 3858 4473 3864 4474
rect 3838 4472 3844 4473
rect 326 4468 332 4469
rect 110 4467 116 4468
rect 110 4463 111 4467
rect 115 4463 116 4467
rect 326 4464 327 4468
rect 331 4464 332 4468
rect 326 4463 332 4464
rect 518 4468 524 4469
rect 518 4464 519 4468
rect 523 4464 524 4468
rect 518 4463 524 4464
rect 718 4468 724 4469
rect 718 4464 719 4468
rect 723 4464 724 4468
rect 718 4463 724 4464
rect 934 4468 940 4469
rect 934 4464 935 4468
rect 939 4464 940 4468
rect 934 4463 940 4464
rect 1150 4468 1156 4469
rect 1150 4464 1151 4468
rect 1155 4464 1156 4468
rect 1150 4463 1156 4464
rect 1374 4468 1380 4469
rect 1374 4464 1375 4468
rect 1379 4464 1380 4468
rect 1374 4463 1380 4464
rect 1606 4468 1612 4469
rect 1606 4464 1607 4468
rect 1611 4464 1612 4468
rect 1606 4463 1612 4464
rect 1814 4468 1820 4469
rect 3838 4468 3839 4472
rect 3843 4468 3844 4472
rect 3858 4469 3859 4473
rect 3863 4469 3864 4473
rect 3858 4468 3864 4469
rect 4034 4473 4040 4474
rect 4034 4469 4035 4473
rect 4039 4469 4040 4473
rect 4034 4468 4040 4469
rect 4250 4473 4256 4474
rect 4250 4469 4251 4473
rect 4255 4469 4256 4473
rect 4250 4468 4256 4469
rect 4474 4473 4480 4474
rect 4474 4469 4475 4473
rect 4479 4469 4480 4473
rect 4474 4468 4480 4469
rect 4722 4473 4728 4474
rect 4722 4469 4723 4473
rect 4727 4469 4728 4473
rect 4722 4468 4728 4469
rect 4978 4473 4984 4474
rect 4978 4469 4979 4473
rect 4983 4469 4984 4473
rect 4978 4468 4984 4469
rect 5242 4473 5248 4474
rect 5242 4469 5243 4473
rect 5247 4469 5248 4473
rect 5242 4468 5248 4469
rect 5514 4473 5520 4474
rect 5514 4469 5515 4473
rect 5519 4469 5520 4473
rect 5514 4468 5520 4469
rect 5662 4472 5668 4473
rect 5662 4468 5663 4472
rect 5667 4468 5668 4472
rect 1814 4464 1815 4468
rect 1819 4464 1820 4468
rect 1814 4463 1820 4464
rect 1934 4467 1940 4468
rect 3838 4467 3844 4468
rect 5662 4467 5668 4468
rect 1934 4463 1935 4467
rect 1939 4463 1940 4467
rect 110 4462 116 4463
rect 1934 4462 1940 4463
rect 110 4409 116 4410
rect 1934 4409 1940 4410
rect 110 4405 111 4409
rect 115 4405 116 4409
rect 110 4404 116 4405
rect 558 4408 564 4409
rect 558 4404 559 4408
rect 563 4404 564 4408
rect 558 4403 564 4404
rect 718 4408 724 4409
rect 718 4404 719 4408
rect 723 4404 724 4408
rect 718 4403 724 4404
rect 886 4408 892 4409
rect 886 4404 887 4408
rect 891 4404 892 4408
rect 886 4403 892 4404
rect 1062 4408 1068 4409
rect 1062 4404 1063 4408
rect 1067 4404 1068 4408
rect 1062 4403 1068 4404
rect 1246 4408 1252 4409
rect 1246 4404 1247 4408
rect 1251 4404 1252 4408
rect 1246 4403 1252 4404
rect 1438 4408 1444 4409
rect 1438 4404 1439 4408
rect 1443 4404 1444 4408
rect 1438 4403 1444 4404
rect 1630 4408 1636 4409
rect 1630 4404 1631 4408
rect 1635 4404 1636 4408
rect 1630 4403 1636 4404
rect 1814 4408 1820 4409
rect 1814 4404 1815 4408
rect 1819 4404 1820 4408
rect 1934 4405 1935 4409
rect 1939 4405 1940 4409
rect 1934 4404 1940 4405
rect 1814 4403 1820 4404
rect 530 4393 536 4394
rect 110 4392 116 4393
rect 110 4388 111 4392
rect 115 4388 116 4392
rect 530 4389 531 4393
rect 535 4389 536 4393
rect 530 4388 536 4389
rect 690 4393 696 4394
rect 690 4389 691 4393
rect 695 4389 696 4393
rect 690 4388 696 4389
rect 858 4393 864 4394
rect 858 4389 859 4393
rect 863 4389 864 4393
rect 858 4388 864 4389
rect 1034 4393 1040 4394
rect 1034 4389 1035 4393
rect 1039 4389 1040 4393
rect 1034 4388 1040 4389
rect 1218 4393 1224 4394
rect 1218 4389 1219 4393
rect 1223 4389 1224 4393
rect 1218 4388 1224 4389
rect 1410 4393 1416 4394
rect 1410 4389 1411 4393
rect 1415 4389 1416 4393
rect 1410 4388 1416 4389
rect 1602 4393 1608 4394
rect 1602 4389 1603 4393
rect 1607 4389 1608 4393
rect 1602 4388 1608 4389
rect 1786 4393 1792 4394
rect 1786 4389 1787 4393
rect 1791 4389 1792 4393
rect 1786 4388 1792 4389
rect 1934 4392 1940 4393
rect 1934 4388 1935 4392
rect 1939 4388 1940 4392
rect 110 4387 116 4388
rect 1934 4387 1940 4388
rect 1974 4380 1980 4381
rect 3798 4380 3804 4381
rect 1974 4376 1975 4380
rect 1979 4376 1980 4380
rect 1974 4375 1980 4376
rect 2570 4379 2576 4380
rect 2570 4375 2571 4379
rect 2575 4375 2576 4379
rect 2570 4374 2576 4375
rect 3122 4379 3128 4380
rect 3122 4375 3123 4379
rect 3127 4375 3128 4379
rect 3122 4374 3128 4375
rect 3650 4379 3656 4380
rect 3650 4375 3651 4379
rect 3655 4375 3656 4379
rect 3798 4376 3799 4380
rect 3803 4376 3804 4380
rect 3798 4375 3804 4376
rect 3650 4374 3656 4375
rect 2598 4364 2604 4365
rect 1974 4363 1980 4364
rect 1974 4359 1975 4363
rect 1979 4359 1980 4363
rect 2598 4360 2599 4364
rect 2603 4360 2604 4364
rect 2598 4359 2604 4360
rect 3150 4364 3156 4365
rect 3150 4360 3151 4364
rect 3155 4360 3156 4364
rect 3150 4359 3156 4360
rect 3678 4364 3684 4365
rect 3678 4360 3679 4364
rect 3683 4360 3684 4364
rect 3678 4359 3684 4360
rect 3798 4363 3804 4364
rect 3798 4359 3799 4363
rect 3803 4359 3804 4363
rect 1974 4358 1980 4359
rect 3798 4358 3804 4359
rect 3838 4340 3844 4341
rect 5662 4340 5668 4341
rect 3838 4336 3839 4340
rect 3843 4336 3844 4340
rect 3838 4335 3844 4336
rect 3858 4339 3864 4340
rect 3858 4335 3859 4339
rect 3863 4335 3864 4339
rect 3858 4334 3864 4335
rect 3994 4339 4000 4340
rect 3994 4335 3995 4339
rect 3999 4335 4000 4339
rect 3994 4334 4000 4335
rect 4130 4339 4136 4340
rect 4130 4335 4131 4339
rect 4135 4335 4136 4339
rect 4130 4334 4136 4335
rect 4266 4339 4272 4340
rect 4266 4335 4267 4339
rect 4271 4335 4272 4339
rect 4266 4334 4272 4335
rect 4402 4339 4408 4340
rect 4402 4335 4403 4339
rect 4407 4335 4408 4339
rect 4402 4334 4408 4335
rect 4586 4339 4592 4340
rect 4586 4335 4587 4339
rect 4591 4335 4592 4339
rect 4586 4334 4592 4335
rect 4794 4339 4800 4340
rect 4794 4335 4795 4339
rect 4799 4335 4800 4339
rect 4794 4334 4800 4335
rect 5026 4339 5032 4340
rect 5026 4335 5027 4339
rect 5031 4335 5032 4339
rect 5026 4334 5032 4335
rect 5274 4339 5280 4340
rect 5274 4335 5275 4339
rect 5279 4335 5280 4339
rect 5274 4334 5280 4335
rect 5514 4339 5520 4340
rect 5514 4335 5515 4339
rect 5519 4335 5520 4339
rect 5662 4336 5663 4340
rect 5667 4336 5668 4340
rect 5662 4335 5668 4336
rect 5514 4334 5520 4335
rect 3886 4324 3892 4325
rect 3838 4323 3844 4324
rect 3838 4319 3839 4323
rect 3843 4319 3844 4323
rect 3886 4320 3887 4324
rect 3891 4320 3892 4324
rect 3886 4319 3892 4320
rect 4022 4324 4028 4325
rect 4022 4320 4023 4324
rect 4027 4320 4028 4324
rect 4022 4319 4028 4320
rect 4158 4324 4164 4325
rect 4158 4320 4159 4324
rect 4163 4320 4164 4324
rect 4158 4319 4164 4320
rect 4294 4324 4300 4325
rect 4294 4320 4295 4324
rect 4299 4320 4300 4324
rect 4294 4319 4300 4320
rect 4430 4324 4436 4325
rect 4430 4320 4431 4324
rect 4435 4320 4436 4324
rect 4430 4319 4436 4320
rect 4614 4324 4620 4325
rect 4614 4320 4615 4324
rect 4619 4320 4620 4324
rect 4614 4319 4620 4320
rect 4822 4324 4828 4325
rect 4822 4320 4823 4324
rect 4827 4320 4828 4324
rect 4822 4319 4828 4320
rect 5054 4324 5060 4325
rect 5054 4320 5055 4324
rect 5059 4320 5060 4324
rect 5054 4319 5060 4320
rect 5302 4324 5308 4325
rect 5302 4320 5303 4324
rect 5307 4320 5308 4324
rect 5302 4319 5308 4320
rect 5542 4324 5548 4325
rect 5542 4320 5543 4324
rect 5547 4320 5548 4324
rect 5542 4319 5548 4320
rect 5662 4323 5668 4324
rect 5662 4319 5663 4323
rect 5667 4319 5668 4323
rect 3838 4318 3844 4319
rect 5662 4318 5668 4319
rect 1974 4301 1980 4302
rect 3798 4301 3804 4302
rect 1974 4297 1975 4301
rect 1979 4297 1980 4301
rect 1974 4296 1980 4297
rect 2398 4300 2404 4301
rect 2398 4296 2399 4300
rect 2403 4296 2404 4300
rect 2398 4295 2404 4296
rect 2598 4300 2604 4301
rect 2598 4296 2599 4300
rect 2603 4296 2604 4300
rect 2598 4295 2604 4296
rect 2790 4300 2796 4301
rect 2790 4296 2791 4300
rect 2795 4296 2796 4300
rect 2790 4295 2796 4296
rect 2982 4300 2988 4301
rect 2982 4296 2983 4300
rect 2987 4296 2988 4300
rect 2982 4295 2988 4296
rect 3166 4300 3172 4301
rect 3166 4296 3167 4300
rect 3171 4296 3172 4300
rect 3166 4295 3172 4296
rect 3342 4300 3348 4301
rect 3342 4296 3343 4300
rect 3347 4296 3348 4300
rect 3342 4295 3348 4296
rect 3518 4300 3524 4301
rect 3518 4296 3519 4300
rect 3523 4296 3524 4300
rect 3518 4295 3524 4296
rect 3678 4300 3684 4301
rect 3678 4296 3679 4300
rect 3683 4296 3684 4300
rect 3798 4297 3799 4301
rect 3803 4297 3804 4301
rect 3798 4296 3804 4297
rect 3678 4295 3684 4296
rect 2370 4285 2376 4286
rect 1974 4284 1980 4285
rect 1974 4280 1975 4284
rect 1979 4280 1980 4284
rect 2370 4281 2371 4285
rect 2375 4281 2376 4285
rect 2370 4280 2376 4281
rect 2570 4285 2576 4286
rect 2570 4281 2571 4285
rect 2575 4281 2576 4285
rect 2570 4280 2576 4281
rect 2762 4285 2768 4286
rect 2762 4281 2763 4285
rect 2767 4281 2768 4285
rect 2762 4280 2768 4281
rect 2954 4285 2960 4286
rect 2954 4281 2955 4285
rect 2959 4281 2960 4285
rect 2954 4280 2960 4281
rect 3138 4285 3144 4286
rect 3138 4281 3139 4285
rect 3143 4281 3144 4285
rect 3138 4280 3144 4281
rect 3314 4285 3320 4286
rect 3314 4281 3315 4285
rect 3319 4281 3320 4285
rect 3314 4280 3320 4281
rect 3490 4285 3496 4286
rect 3490 4281 3491 4285
rect 3495 4281 3496 4285
rect 3490 4280 3496 4281
rect 3650 4285 3656 4286
rect 3650 4281 3651 4285
rect 3655 4281 3656 4285
rect 3650 4280 3656 4281
rect 3798 4284 3804 4285
rect 3798 4280 3799 4284
rect 3803 4280 3804 4284
rect 1974 4279 1980 4280
rect 3798 4279 3804 4280
rect 3838 4265 3844 4266
rect 5662 4265 5668 4266
rect 3838 4261 3839 4265
rect 3843 4261 3844 4265
rect 3838 4260 3844 4261
rect 4046 4264 4052 4265
rect 4046 4260 4047 4264
rect 4051 4260 4052 4264
rect 4046 4259 4052 4260
rect 4222 4264 4228 4265
rect 4222 4260 4223 4264
rect 4227 4260 4228 4264
rect 4222 4259 4228 4260
rect 4430 4264 4436 4265
rect 4430 4260 4431 4264
rect 4435 4260 4436 4264
rect 4430 4259 4436 4260
rect 4678 4264 4684 4265
rect 4678 4260 4679 4264
rect 4683 4260 4684 4264
rect 4678 4259 4684 4260
rect 4958 4264 4964 4265
rect 4958 4260 4959 4264
rect 4963 4260 4964 4264
rect 4958 4259 4964 4260
rect 5254 4264 5260 4265
rect 5254 4260 5255 4264
rect 5259 4260 5260 4264
rect 5254 4259 5260 4260
rect 5542 4264 5548 4265
rect 5542 4260 5543 4264
rect 5547 4260 5548 4264
rect 5662 4261 5663 4265
rect 5667 4261 5668 4265
rect 5662 4260 5668 4261
rect 5542 4259 5548 4260
rect 110 4252 116 4253
rect 1934 4252 1940 4253
rect 110 4248 111 4252
rect 115 4248 116 4252
rect 110 4247 116 4248
rect 746 4251 752 4252
rect 746 4247 747 4251
rect 751 4247 752 4251
rect 746 4246 752 4247
rect 882 4251 888 4252
rect 882 4247 883 4251
rect 887 4247 888 4251
rect 882 4246 888 4247
rect 1018 4251 1024 4252
rect 1018 4247 1019 4251
rect 1023 4247 1024 4251
rect 1018 4246 1024 4247
rect 1154 4251 1160 4252
rect 1154 4247 1155 4251
rect 1159 4247 1160 4251
rect 1154 4246 1160 4247
rect 1290 4251 1296 4252
rect 1290 4247 1291 4251
rect 1295 4247 1296 4251
rect 1290 4246 1296 4247
rect 1426 4251 1432 4252
rect 1426 4247 1427 4251
rect 1431 4247 1432 4251
rect 1426 4246 1432 4247
rect 1562 4251 1568 4252
rect 1562 4247 1563 4251
rect 1567 4247 1568 4251
rect 1562 4246 1568 4247
rect 1698 4251 1704 4252
rect 1698 4247 1699 4251
rect 1703 4247 1704 4251
rect 1934 4248 1935 4252
rect 1939 4248 1940 4252
rect 4018 4249 4024 4250
rect 1934 4247 1940 4248
rect 3838 4248 3844 4249
rect 1698 4246 1704 4247
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 4018 4245 4019 4249
rect 4023 4245 4024 4249
rect 4018 4244 4024 4245
rect 4194 4249 4200 4250
rect 4194 4245 4195 4249
rect 4199 4245 4200 4249
rect 4194 4244 4200 4245
rect 4402 4249 4408 4250
rect 4402 4245 4403 4249
rect 4407 4245 4408 4249
rect 4402 4244 4408 4245
rect 4650 4249 4656 4250
rect 4650 4245 4651 4249
rect 4655 4245 4656 4249
rect 4650 4244 4656 4245
rect 4930 4249 4936 4250
rect 4930 4245 4931 4249
rect 4935 4245 4936 4249
rect 4930 4244 4936 4245
rect 5226 4249 5232 4250
rect 5226 4245 5227 4249
rect 5231 4245 5232 4249
rect 5226 4244 5232 4245
rect 5514 4249 5520 4250
rect 5514 4245 5515 4249
rect 5519 4245 5520 4249
rect 5514 4244 5520 4245
rect 5662 4248 5668 4249
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 3838 4243 3844 4244
rect 5662 4243 5668 4244
rect 774 4236 780 4237
rect 110 4235 116 4236
rect 110 4231 111 4235
rect 115 4231 116 4235
rect 774 4232 775 4236
rect 779 4232 780 4236
rect 774 4231 780 4232
rect 910 4236 916 4237
rect 910 4232 911 4236
rect 915 4232 916 4236
rect 910 4231 916 4232
rect 1046 4236 1052 4237
rect 1046 4232 1047 4236
rect 1051 4232 1052 4236
rect 1046 4231 1052 4232
rect 1182 4236 1188 4237
rect 1182 4232 1183 4236
rect 1187 4232 1188 4236
rect 1182 4231 1188 4232
rect 1318 4236 1324 4237
rect 1318 4232 1319 4236
rect 1323 4232 1324 4236
rect 1318 4231 1324 4232
rect 1454 4236 1460 4237
rect 1454 4232 1455 4236
rect 1459 4232 1460 4236
rect 1454 4231 1460 4232
rect 1590 4236 1596 4237
rect 1590 4232 1591 4236
rect 1595 4232 1596 4236
rect 1590 4231 1596 4232
rect 1726 4236 1732 4237
rect 1726 4232 1727 4236
rect 1731 4232 1732 4236
rect 1726 4231 1732 4232
rect 1934 4235 1940 4236
rect 1934 4231 1935 4235
rect 1939 4231 1940 4235
rect 110 4230 116 4231
rect 1934 4230 1940 4231
rect 110 4165 116 4166
rect 1934 4165 1940 4166
rect 110 4161 111 4165
rect 115 4161 116 4165
rect 110 4160 116 4161
rect 726 4164 732 4165
rect 726 4160 727 4164
rect 731 4160 732 4164
rect 726 4159 732 4160
rect 862 4164 868 4165
rect 862 4160 863 4164
rect 867 4160 868 4164
rect 862 4159 868 4160
rect 998 4164 1004 4165
rect 998 4160 999 4164
rect 1003 4160 1004 4164
rect 998 4159 1004 4160
rect 1134 4164 1140 4165
rect 1134 4160 1135 4164
rect 1139 4160 1140 4164
rect 1134 4159 1140 4160
rect 1270 4164 1276 4165
rect 1270 4160 1271 4164
rect 1275 4160 1276 4164
rect 1270 4159 1276 4160
rect 1406 4164 1412 4165
rect 1406 4160 1407 4164
rect 1411 4160 1412 4164
rect 1406 4159 1412 4160
rect 1542 4164 1548 4165
rect 1542 4160 1543 4164
rect 1547 4160 1548 4164
rect 1542 4159 1548 4160
rect 1678 4164 1684 4165
rect 1678 4160 1679 4164
rect 1683 4160 1684 4164
rect 1678 4159 1684 4160
rect 1814 4164 1820 4165
rect 1814 4160 1815 4164
rect 1819 4160 1820 4164
rect 1934 4161 1935 4165
rect 1939 4161 1940 4165
rect 1934 4160 1940 4161
rect 1814 4159 1820 4160
rect 698 4149 704 4150
rect 110 4148 116 4149
rect 110 4144 111 4148
rect 115 4144 116 4148
rect 698 4145 699 4149
rect 703 4145 704 4149
rect 698 4144 704 4145
rect 834 4149 840 4150
rect 834 4145 835 4149
rect 839 4145 840 4149
rect 834 4144 840 4145
rect 970 4149 976 4150
rect 970 4145 971 4149
rect 975 4145 976 4149
rect 970 4144 976 4145
rect 1106 4149 1112 4150
rect 1106 4145 1107 4149
rect 1111 4145 1112 4149
rect 1106 4144 1112 4145
rect 1242 4149 1248 4150
rect 1242 4145 1243 4149
rect 1247 4145 1248 4149
rect 1242 4144 1248 4145
rect 1378 4149 1384 4150
rect 1378 4145 1379 4149
rect 1383 4145 1384 4149
rect 1378 4144 1384 4145
rect 1514 4149 1520 4150
rect 1514 4145 1515 4149
rect 1519 4145 1520 4149
rect 1514 4144 1520 4145
rect 1650 4149 1656 4150
rect 1650 4145 1651 4149
rect 1655 4145 1656 4149
rect 1650 4144 1656 4145
rect 1786 4149 1792 4150
rect 1786 4145 1787 4149
rect 1791 4145 1792 4149
rect 1786 4144 1792 4145
rect 1934 4148 1940 4149
rect 1934 4144 1935 4148
rect 1939 4144 1940 4148
rect 110 4143 116 4144
rect 1934 4143 1940 4144
rect 1974 4140 1980 4141
rect 3798 4140 3804 4141
rect 1974 4136 1975 4140
rect 1979 4136 1980 4140
rect 1974 4135 1980 4136
rect 2370 4139 2376 4140
rect 2370 4135 2371 4139
rect 2375 4135 2376 4139
rect 2370 4134 2376 4135
rect 2610 4139 2616 4140
rect 2610 4135 2611 4139
rect 2615 4135 2616 4139
rect 2610 4134 2616 4135
rect 2834 4139 2840 4140
rect 2834 4135 2835 4139
rect 2839 4135 2840 4139
rect 2834 4134 2840 4135
rect 3050 4139 3056 4140
rect 3050 4135 3051 4139
rect 3055 4135 3056 4139
rect 3050 4134 3056 4135
rect 3258 4139 3264 4140
rect 3258 4135 3259 4139
rect 3263 4135 3264 4139
rect 3258 4134 3264 4135
rect 3466 4139 3472 4140
rect 3466 4135 3467 4139
rect 3471 4135 3472 4139
rect 3466 4134 3472 4135
rect 3650 4139 3656 4140
rect 3650 4135 3651 4139
rect 3655 4135 3656 4139
rect 3798 4136 3799 4140
rect 3803 4136 3804 4140
rect 3798 4135 3804 4136
rect 3650 4134 3656 4135
rect 2398 4124 2404 4125
rect 1974 4123 1980 4124
rect 1974 4119 1975 4123
rect 1979 4119 1980 4123
rect 2398 4120 2399 4124
rect 2403 4120 2404 4124
rect 2398 4119 2404 4120
rect 2638 4124 2644 4125
rect 2638 4120 2639 4124
rect 2643 4120 2644 4124
rect 2638 4119 2644 4120
rect 2862 4124 2868 4125
rect 2862 4120 2863 4124
rect 2867 4120 2868 4124
rect 2862 4119 2868 4120
rect 3078 4124 3084 4125
rect 3078 4120 3079 4124
rect 3083 4120 3084 4124
rect 3078 4119 3084 4120
rect 3286 4124 3292 4125
rect 3286 4120 3287 4124
rect 3291 4120 3292 4124
rect 3286 4119 3292 4120
rect 3494 4124 3500 4125
rect 3494 4120 3495 4124
rect 3499 4120 3500 4124
rect 3494 4119 3500 4120
rect 3678 4124 3684 4125
rect 3678 4120 3679 4124
rect 3683 4120 3684 4124
rect 3678 4119 3684 4120
rect 3798 4123 3804 4124
rect 3798 4119 3799 4123
rect 3803 4119 3804 4123
rect 1974 4118 1980 4119
rect 3798 4118 3804 4119
rect 1974 4061 1980 4062
rect 3798 4061 3804 4062
rect 1974 4057 1975 4061
rect 1979 4057 1980 4061
rect 1974 4056 1980 4057
rect 2374 4060 2380 4061
rect 2374 4056 2375 4060
rect 2379 4056 2380 4060
rect 2374 4055 2380 4056
rect 2622 4060 2628 4061
rect 2622 4056 2623 4060
rect 2627 4056 2628 4060
rect 2622 4055 2628 4056
rect 2854 4060 2860 4061
rect 2854 4056 2855 4060
rect 2859 4056 2860 4060
rect 2854 4055 2860 4056
rect 3070 4060 3076 4061
rect 3070 4056 3071 4060
rect 3075 4056 3076 4060
rect 3070 4055 3076 4056
rect 3278 4060 3284 4061
rect 3278 4056 3279 4060
rect 3283 4056 3284 4060
rect 3278 4055 3284 4056
rect 3486 4060 3492 4061
rect 3486 4056 3487 4060
rect 3491 4056 3492 4060
rect 3486 4055 3492 4056
rect 3678 4060 3684 4061
rect 3678 4056 3679 4060
rect 3683 4056 3684 4060
rect 3798 4057 3799 4061
rect 3803 4057 3804 4061
rect 3798 4056 3804 4057
rect 3678 4055 3684 4056
rect 2346 4045 2352 4046
rect 1974 4044 1980 4045
rect 1974 4040 1975 4044
rect 1979 4040 1980 4044
rect 2346 4041 2347 4045
rect 2351 4041 2352 4045
rect 2346 4040 2352 4041
rect 2594 4045 2600 4046
rect 2594 4041 2595 4045
rect 2599 4041 2600 4045
rect 2594 4040 2600 4041
rect 2826 4045 2832 4046
rect 2826 4041 2827 4045
rect 2831 4041 2832 4045
rect 2826 4040 2832 4041
rect 3042 4045 3048 4046
rect 3042 4041 3043 4045
rect 3047 4041 3048 4045
rect 3042 4040 3048 4041
rect 3250 4045 3256 4046
rect 3250 4041 3251 4045
rect 3255 4041 3256 4045
rect 3250 4040 3256 4041
rect 3458 4045 3464 4046
rect 3458 4041 3459 4045
rect 3463 4041 3464 4045
rect 3458 4040 3464 4041
rect 3650 4045 3656 4046
rect 3650 4041 3651 4045
rect 3655 4041 3656 4045
rect 3650 4040 3656 4041
rect 3798 4044 3804 4045
rect 3798 4040 3799 4044
rect 3803 4040 3804 4044
rect 1974 4039 1980 4040
rect 3798 4039 3804 4040
rect 3838 4032 3844 4033
rect 5662 4032 5668 4033
rect 3838 4028 3839 4032
rect 3843 4028 3844 4032
rect 3838 4027 3844 4028
rect 5514 4031 5520 4032
rect 5514 4027 5515 4031
rect 5519 4027 5520 4031
rect 5662 4028 5663 4032
rect 5667 4028 5668 4032
rect 5662 4027 5668 4028
rect 5514 4026 5520 4027
rect 5542 4016 5548 4017
rect 3838 4015 3844 4016
rect 3838 4011 3839 4015
rect 3843 4011 3844 4015
rect 5542 4012 5543 4016
rect 5547 4012 5548 4016
rect 5542 4011 5548 4012
rect 5662 4015 5668 4016
rect 5662 4011 5663 4015
rect 5667 4011 5668 4015
rect 3838 4010 3844 4011
rect 5662 4010 5668 4011
rect 110 4004 116 4005
rect 1934 4004 1940 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 626 4003 632 4004
rect 626 3999 627 4003
rect 631 3999 632 4003
rect 626 3998 632 3999
rect 762 4003 768 4004
rect 762 3999 763 4003
rect 767 3999 768 4003
rect 762 3998 768 3999
rect 898 4003 904 4004
rect 898 3999 899 4003
rect 903 3999 904 4003
rect 898 3998 904 3999
rect 1034 4003 1040 4004
rect 1034 3999 1035 4003
rect 1039 3999 1040 4003
rect 1034 3998 1040 3999
rect 1170 4003 1176 4004
rect 1170 3999 1171 4003
rect 1175 3999 1176 4003
rect 1170 3998 1176 3999
rect 1306 4003 1312 4004
rect 1306 3999 1307 4003
rect 1311 3999 1312 4003
rect 1306 3998 1312 3999
rect 1442 4003 1448 4004
rect 1442 3999 1443 4003
rect 1447 3999 1448 4003
rect 1442 3998 1448 3999
rect 1578 4003 1584 4004
rect 1578 3999 1579 4003
rect 1583 3999 1584 4003
rect 1578 3998 1584 3999
rect 1714 4003 1720 4004
rect 1714 3999 1715 4003
rect 1719 3999 1720 4003
rect 1934 4000 1935 4004
rect 1939 4000 1940 4004
rect 1934 3999 1940 4000
rect 1714 3998 1720 3999
rect 654 3988 660 3989
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 654 3984 655 3988
rect 659 3984 660 3988
rect 654 3983 660 3984
rect 790 3988 796 3989
rect 790 3984 791 3988
rect 795 3984 796 3988
rect 790 3983 796 3984
rect 926 3988 932 3989
rect 926 3984 927 3988
rect 931 3984 932 3988
rect 926 3983 932 3984
rect 1062 3988 1068 3989
rect 1062 3984 1063 3988
rect 1067 3984 1068 3988
rect 1062 3983 1068 3984
rect 1198 3988 1204 3989
rect 1198 3984 1199 3988
rect 1203 3984 1204 3988
rect 1198 3983 1204 3984
rect 1334 3988 1340 3989
rect 1334 3984 1335 3988
rect 1339 3984 1340 3988
rect 1334 3983 1340 3984
rect 1470 3988 1476 3989
rect 1470 3984 1471 3988
rect 1475 3984 1476 3988
rect 1470 3983 1476 3984
rect 1606 3988 1612 3989
rect 1606 3984 1607 3988
rect 1611 3984 1612 3988
rect 1606 3983 1612 3984
rect 1742 3988 1748 3989
rect 1742 3984 1743 3988
rect 1747 3984 1748 3988
rect 1742 3983 1748 3984
rect 1934 3987 1940 3988
rect 1934 3983 1935 3987
rect 1939 3983 1940 3987
rect 110 3982 116 3983
rect 1934 3982 1940 3983
rect 3838 3949 3844 3950
rect 5662 3949 5668 3950
rect 3838 3945 3839 3949
rect 3843 3945 3844 3949
rect 3838 3944 3844 3945
rect 4182 3948 4188 3949
rect 4182 3944 4183 3948
rect 4187 3944 4188 3948
rect 4182 3943 4188 3944
rect 4318 3948 4324 3949
rect 4318 3944 4319 3948
rect 4323 3944 4324 3948
rect 4318 3943 4324 3944
rect 4454 3948 4460 3949
rect 4454 3944 4455 3948
rect 4459 3944 4460 3948
rect 4454 3943 4460 3944
rect 4590 3948 4596 3949
rect 4590 3944 4591 3948
rect 4595 3944 4596 3948
rect 4590 3943 4596 3944
rect 4726 3948 4732 3949
rect 4726 3944 4727 3948
rect 4731 3944 4732 3948
rect 4726 3943 4732 3944
rect 4862 3948 4868 3949
rect 4862 3944 4863 3948
rect 4867 3944 4868 3948
rect 4862 3943 4868 3944
rect 4998 3948 5004 3949
rect 4998 3944 4999 3948
rect 5003 3944 5004 3948
rect 4998 3943 5004 3944
rect 5134 3948 5140 3949
rect 5134 3944 5135 3948
rect 5139 3944 5140 3948
rect 5134 3943 5140 3944
rect 5270 3948 5276 3949
rect 5270 3944 5271 3948
rect 5275 3944 5276 3948
rect 5270 3943 5276 3944
rect 5406 3948 5412 3949
rect 5406 3944 5407 3948
rect 5411 3944 5412 3948
rect 5406 3943 5412 3944
rect 5542 3948 5548 3949
rect 5542 3944 5543 3948
rect 5547 3944 5548 3948
rect 5662 3945 5663 3949
rect 5667 3945 5668 3949
rect 5662 3944 5668 3945
rect 5542 3943 5548 3944
rect 4154 3933 4160 3934
rect 3838 3932 3844 3933
rect 3838 3928 3839 3932
rect 3843 3928 3844 3932
rect 4154 3929 4155 3933
rect 4159 3929 4160 3933
rect 4154 3928 4160 3929
rect 4290 3933 4296 3934
rect 4290 3929 4291 3933
rect 4295 3929 4296 3933
rect 4290 3928 4296 3929
rect 4426 3933 4432 3934
rect 4426 3929 4427 3933
rect 4431 3929 4432 3933
rect 4426 3928 4432 3929
rect 4562 3933 4568 3934
rect 4562 3929 4563 3933
rect 4567 3929 4568 3933
rect 4562 3928 4568 3929
rect 4698 3933 4704 3934
rect 4698 3929 4699 3933
rect 4703 3929 4704 3933
rect 4698 3928 4704 3929
rect 4834 3933 4840 3934
rect 4834 3929 4835 3933
rect 4839 3929 4840 3933
rect 4834 3928 4840 3929
rect 4970 3933 4976 3934
rect 4970 3929 4971 3933
rect 4975 3929 4976 3933
rect 4970 3928 4976 3929
rect 5106 3933 5112 3934
rect 5106 3929 5107 3933
rect 5111 3929 5112 3933
rect 5106 3928 5112 3929
rect 5242 3933 5248 3934
rect 5242 3929 5243 3933
rect 5247 3929 5248 3933
rect 5242 3928 5248 3929
rect 5378 3933 5384 3934
rect 5378 3929 5379 3933
rect 5383 3929 5384 3933
rect 5378 3928 5384 3929
rect 5514 3933 5520 3934
rect 5514 3929 5515 3933
rect 5519 3929 5520 3933
rect 5514 3928 5520 3929
rect 5662 3932 5668 3933
rect 5662 3928 5663 3932
rect 5667 3928 5668 3932
rect 3838 3927 3844 3928
rect 5662 3927 5668 3928
rect 110 3917 116 3918
rect 1934 3917 1940 3918
rect 110 3913 111 3917
rect 115 3913 116 3917
rect 110 3912 116 3913
rect 598 3916 604 3917
rect 598 3912 599 3916
rect 603 3912 604 3916
rect 598 3911 604 3912
rect 742 3916 748 3917
rect 742 3912 743 3916
rect 747 3912 748 3916
rect 742 3911 748 3912
rect 894 3916 900 3917
rect 894 3912 895 3916
rect 899 3912 900 3916
rect 894 3911 900 3912
rect 1046 3916 1052 3917
rect 1046 3912 1047 3916
rect 1051 3912 1052 3916
rect 1046 3911 1052 3912
rect 1198 3916 1204 3917
rect 1198 3912 1199 3916
rect 1203 3912 1204 3916
rect 1198 3911 1204 3912
rect 1358 3916 1364 3917
rect 1358 3912 1359 3916
rect 1363 3912 1364 3916
rect 1358 3911 1364 3912
rect 1518 3916 1524 3917
rect 1518 3912 1519 3916
rect 1523 3912 1524 3916
rect 1518 3911 1524 3912
rect 1678 3916 1684 3917
rect 1678 3912 1679 3916
rect 1683 3912 1684 3916
rect 1934 3913 1935 3917
rect 1939 3913 1940 3917
rect 1934 3912 1940 3913
rect 1974 3912 1980 3913
rect 3798 3912 3804 3913
rect 1678 3911 1684 3912
rect 1974 3908 1975 3912
rect 1979 3908 1980 3912
rect 1974 3907 1980 3908
rect 2322 3911 2328 3912
rect 2322 3907 2323 3911
rect 2327 3907 2328 3911
rect 2322 3906 2328 3907
rect 2570 3911 2576 3912
rect 2570 3907 2571 3911
rect 2575 3907 2576 3911
rect 2570 3906 2576 3907
rect 2802 3911 2808 3912
rect 2802 3907 2803 3911
rect 2807 3907 2808 3911
rect 2802 3906 2808 3907
rect 3026 3911 3032 3912
rect 3026 3907 3027 3911
rect 3031 3907 3032 3911
rect 3026 3906 3032 3907
rect 3242 3911 3248 3912
rect 3242 3907 3243 3911
rect 3247 3907 3248 3911
rect 3242 3906 3248 3907
rect 3458 3911 3464 3912
rect 3458 3907 3459 3911
rect 3463 3907 3464 3911
rect 3458 3906 3464 3907
rect 3650 3911 3656 3912
rect 3650 3907 3651 3911
rect 3655 3907 3656 3911
rect 3798 3908 3799 3912
rect 3803 3908 3804 3912
rect 3798 3907 3804 3908
rect 3650 3906 3656 3907
rect 570 3901 576 3902
rect 110 3900 116 3901
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 570 3897 571 3901
rect 575 3897 576 3901
rect 570 3896 576 3897
rect 714 3901 720 3902
rect 714 3897 715 3901
rect 719 3897 720 3901
rect 714 3896 720 3897
rect 866 3901 872 3902
rect 866 3897 867 3901
rect 871 3897 872 3901
rect 866 3896 872 3897
rect 1018 3901 1024 3902
rect 1018 3897 1019 3901
rect 1023 3897 1024 3901
rect 1018 3896 1024 3897
rect 1170 3901 1176 3902
rect 1170 3897 1171 3901
rect 1175 3897 1176 3901
rect 1170 3896 1176 3897
rect 1330 3901 1336 3902
rect 1330 3897 1331 3901
rect 1335 3897 1336 3901
rect 1330 3896 1336 3897
rect 1490 3901 1496 3902
rect 1490 3897 1491 3901
rect 1495 3897 1496 3901
rect 1490 3896 1496 3897
rect 1650 3901 1656 3902
rect 1650 3897 1651 3901
rect 1655 3897 1656 3901
rect 1650 3896 1656 3897
rect 1934 3900 1940 3901
rect 1934 3896 1935 3900
rect 1939 3896 1940 3900
rect 2350 3896 2356 3897
rect 110 3895 116 3896
rect 1934 3895 1940 3896
rect 1974 3895 1980 3896
rect 1974 3891 1975 3895
rect 1979 3891 1980 3895
rect 2350 3892 2351 3896
rect 2355 3892 2356 3896
rect 2350 3891 2356 3892
rect 2598 3896 2604 3897
rect 2598 3892 2599 3896
rect 2603 3892 2604 3896
rect 2598 3891 2604 3892
rect 2830 3896 2836 3897
rect 2830 3892 2831 3896
rect 2835 3892 2836 3896
rect 2830 3891 2836 3892
rect 3054 3896 3060 3897
rect 3054 3892 3055 3896
rect 3059 3892 3060 3896
rect 3054 3891 3060 3892
rect 3270 3896 3276 3897
rect 3270 3892 3271 3896
rect 3275 3892 3276 3896
rect 3270 3891 3276 3892
rect 3486 3896 3492 3897
rect 3486 3892 3487 3896
rect 3491 3892 3492 3896
rect 3486 3891 3492 3892
rect 3678 3896 3684 3897
rect 3678 3892 3679 3896
rect 3683 3892 3684 3896
rect 3678 3891 3684 3892
rect 3798 3895 3804 3896
rect 3798 3891 3799 3895
rect 3803 3891 3804 3895
rect 1974 3890 1980 3891
rect 3798 3890 3804 3891
rect 1974 3833 1980 3834
rect 3798 3833 3804 3834
rect 1974 3829 1975 3833
rect 1979 3829 1980 3833
rect 1974 3828 1980 3829
rect 2238 3832 2244 3833
rect 2238 3828 2239 3832
rect 2243 3828 2244 3832
rect 2238 3827 2244 3828
rect 2478 3832 2484 3833
rect 2478 3828 2479 3832
rect 2483 3828 2484 3832
rect 2478 3827 2484 3828
rect 2702 3832 2708 3833
rect 2702 3828 2703 3832
rect 2707 3828 2708 3832
rect 2702 3827 2708 3828
rect 2918 3832 2924 3833
rect 2918 3828 2919 3832
rect 2923 3828 2924 3832
rect 2918 3827 2924 3828
rect 3118 3832 3124 3833
rect 3118 3828 3119 3832
rect 3123 3828 3124 3832
rect 3118 3827 3124 3828
rect 3310 3832 3316 3833
rect 3310 3828 3311 3832
rect 3315 3828 3316 3832
rect 3310 3827 3316 3828
rect 3502 3832 3508 3833
rect 3502 3828 3503 3832
rect 3507 3828 3508 3832
rect 3502 3827 3508 3828
rect 3678 3832 3684 3833
rect 3678 3828 3679 3832
rect 3683 3828 3684 3832
rect 3798 3829 3799 3833
rect 3803 3829 3804 3833
rect 3798 3828 3804 3829
rect 3678 3827 3684 3828
rect 2210 3817 2216 3818
rect 1974 3816 1980 3817
rect 1974 3812 1975 3816
rect 1979 3812 1980 3816
rect 2210 3813 2211 3817
rect 2215 3813 2216 3817
rect 2210 3812 2216 3813
rect 2450 3817 2456 3818
rect 2450 3813 2451 3817
rect 2455 3813 2456 3817
rect 2450 3812 2456 3813
rect 2674 3817 2680 3818
rect 2674 3813 2675 3817
rect 2679 3813 2680 3817
rect 2674 3812 2680 3813
rect 2890 3817 2896 3818
rect 2890 3813 2891 3817
rect 2895 3813 2896 3817
rect 2890 3812 2896 3813
rect 3090 3817 3096 3818
rect 3090 3813 3091 3817
rect 3095 3813 3096 3817
rect 3090 3812 3096 3813
rect 3282 3817 3288 3818
rect 3282 3813 3283 3817
rect 3287 3813 3288 3817
rect 3282 3812 3288 3813
rect 3474 3817 3480 3818
rect 3474 3813 3475 3817
rect 3479 3813 3480 3817
rect 3474 3812 3480 3813
rect 3650 3817 3656 3818
rect 3650 3813 3651 3817
rect 3655 3813 3656 3817
rect 3650 3812 3656 3813
rect 3798 3816 3804 3817
rect 3798 3812 3799 3816
rect 3803 3812 3804 3816
rect 1974 3811 1980 3812
rect 3798 3811 3804 3812
rect 3838 3768 3844 3769
rect 5662 3768 5668 3769
rect 3838 3764 3839 3768
rect 3843 3764 3844 3768
rect 3838 3763 3844 3764
rect 4138 3767 4144 3768
rect 4138 3763 4139 3767
rect 4143 3763 4144 3767
rect 4138 3762 4144 3763
rect 4322 3767 4328 3768
rect 4322 3763 4323 3767
rect 4327 3763 4328 3767
rect 4322 3762 4328 3763
rect 4530 3767 4536 3768
rect 4530 3763 4531 3767
rect 4535 3763 4536 3767
rect 4530 3762 4536 3763
rect 4762 3767 4768 3768
rect 4762 3763 4763 3767
rect 4767 3763 4768 3767
rect 4762 3762 4768 3763
rect 5010 3767 5016 3768
rect 5010 3763 5011 3767
rect 5015 3763 5016 3767
rect 5010 3762 5016 3763
rect 5274 3767 5280 3768
rect 5274 3763 5275 3767
rect 5279 3763 5280 3767
rect 5274 3762 5280 3763
rect 5514 3767 5520 3768
rect 5514 3763 5515 3767
rect 5519 3763 5520 3767
rect 5662 3764 5663 3768
rect 5667 3764 5668 3768
rect 5662 3763 5668 3764
rect 5514 3762 5520 3763
rect 110 3760 116 3761
rect 1934 3760 1940 3761
rect 110 3756 111 3760
rect 115 3756 116 3760
rect 110 3755 116 3756
rect 426 3759 432 3760
rect 426 3755 427 3759
rect 431 3755 432 3759
rect 426 3754 432 3755
rect 586 3759 592 3760
rect 586 3755 587 3759
rect 591 3755 592 3759
rect 586 3754 592 3755
rect 754 3759 760 3760
rect 754 3755 755 3759
rect 759 3755 760 3759
rect 754 3754 760 3755
rect 922 3759 928 3760
rect 922 3755 923 3759
rect 927 3755 928 3759
rect 922 3754 928 3755
rect 1098 3759 1104 3760
rect 1098 3755 1099 3759
rect 1103 3755 1104 3759
rect 1098 3754 1104 3755
rect 1274 3759 1280 3760
rect 1274 3755 1275 3759
rect 1279 3755 1280 3759
rect 1274 3754 1280 3755
rect 1458 3759 1464 3760
rect 1458 3755 1459 3759
rect 1463 3755 1464 3759
rect 1458 3754 1464 3755
rect 1642 3759 1648 3760
rect 1642 3755 1643 3759
rect 1647 3755 1648 3759
rect 1934 3756 1935 3760
rect 1939 3756 1940 3760
rect 1934 3755 1940 3756
rect 1642 3754 1648 3755
rect 4166 3752 4172 3753
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 4166 3748 4167 3752
rect 4171 3748 4172 3752
rect 4166 3747 4172 3748
rect 4350 3752 4356 3753
rect 4350 3748 4351 3752
rect 4355 3748 4356 3752
rect 4350 3747 4356 3748
rect 4558 3752 4564 3753
rect 4558 3748 4559 3752
rect 4563 3748 4564 3752
rect 4558 3747 4564 3748
rect 4790 3752 4796 3753
rect 4790 3748 4791 3752
rect 4795 3748 4796 3752
rect 4790 3747 4796 3748
rect 5038 3752 5044 3753
rect 5038 3748 5039 3752
rect 5043 3748 5044 3752
rect 5038 3747 5044 3748
rect 5302 3752 5308 3753
rect 5302 3748 5303 3752
rect 5307 3748 5308 3752
rect 5302 3747 5308 3748
rect 5542 3752 5548 3753
rect 5542 3748 5543 3752
rect 5547 3748 5548 3752
rect 5542 3747 5548 3748
rect 5662 3751 5668 3752
rect 5662 3747 5663 3751
rect 5667 3747 5668 3751
rect 3838 3746 3844 3747
rect 5662 3746 5668 3747
rect 454 3744 460 3745
rect 110 3743 116 3744
rect 110 3739 111 3743
rect 115 3739 116 3743
rect 454 3740 455 3744
rect 459 3740 460 3744
rect 454 3739 460 3740
rect 614 3744 620 3745
rect 614 3740 615 3744
rect 619 3740 620 3744
rect 614 3739 620 3740
rect 782 3744 788 3745
rect 782 3740 783 3744
rect 787 3740 788 3744
rect 782 3739 788 3740
rect 950 3744 956 3745
rect 950 3740 951 3744
rect 955 3740 956 3744
rect 950 3739 956 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1302 3744 1308 3745
rect 1302 3740 1303 3744
rect 1307 3740 1308 3744
rect 1302 3739 1308 3740
rect 1486 3744 1492 3745
rect 1486 3740 1487 3744
rect 1491 3740 1492 3744
rect 1486 3739 1492 3740
rect 1670 3744 1676 3745
rect 1670 3740 1671 3744
rect 1675 3740 1676 3744
rect 1670 3739 1676 3740
rect 1934 3743 1940 3744
rect 1934 3739 1935 3743
rect 1939 3739 1940 3743
rect 110 3738 116 3739
rect 1934 3738 1940 3739
rect 1974 3676 1980 3677
rect 3798 3676 3804 3677
rect 110 3673 116 3674
rect 1934 3673 1940 3674
rect 110 3669 111 3673
rect 115 3669 116 3673
rect 110 3668 116 3669
rect 326 3672 332 3673
rect 326 3668 327 3672
rect 331 3668 332 3672
rect 326 3667 332 3668
rect 494 3672 500 3673
rect 494 3668 495 3672
rect 499 3668 500 3672
rect 494 3667 500 3668
rect 678 3672 684 3673
rect 678 3668 679 3672
rect 683 3668 684 3672
rect 678 3667 684 3668
rect 862 3672 868 3673
rect 862 3668 863 3672
rect 867 3668 868 3672
rect 862 3667 868 3668
rect 1054 3672 1060 3673
rect 1054 3668 1055 3672
rect 1059 3668 1060 3672
rect 1054 3667 1060 3668
rect 1254 3672 1260 3673
rect 1254 3668 1255 3672
rect 1259 3668 1260 3672
rect 1254 3667 1260 3668
rect 1454 3672 1460 3673
rect 1454 3668 1455 3672
rect 1459 3668 1460 3672
rect 1454 3667 1460 3668
rect 1654 3672 1660 3673
rect 1654 3668 1655 3672
rect 1659 3668 1660 3672
rect 1934 3669 1935 3673
rect 1939 3669 1940 3673
rect 1974 3672 1975 3676
rect 1979 3672 1980 3676
rect 1974 3671 1980 3672
rect 2226 3675 2232 3676
rect 2226 3671 2227 3675
rect 2231 3671 2232 3675
rect 2226 3670 2232 3671
rect 2450 3675 2456 3676
rect 2450 3671 2451 3675
rect 2455 3671 2456 3675
rect 2450 3670 2456 3671
rect 2666 3675 2672 3676
rect 2666 3671 2667 3675
rect 2671 3671 2672 3675
rect 2666 3670 2672 3671
rect 2874 3675 2880 3676
rect 2874 3671 2875 3675
rect 2879 3671 2880 3675
rect 2874 3670 2880 3671
rect 3074 3675 3080 3676
rect 3074 3671 3075 3675
rect 3079 3671 3080 3675
rect 3074 3670 3080 3671
rect 3274 3675 3280 3676
rect 3274 3671 3275 3675
rect 3279 3671 3280 3675
rect 3274 3670 3280 3671
rect 3474 3675 3480 3676
rect 3474 3671 3475 3675
rect 3479 3671 3480 3675
rect 3798 3672 3799 3676
rect 3803 3672 3804 3676
rect 3798 3671 3804 3672
rect 3838 3673 3844 3674
rect 5662 3673 5668 3674
rect 3474 3670 3480 3671
rect 1934 3668 1940 3669
rect 3838 3669 3839 3673
rect 3843 3669 3844 3673
rect 3838 3668 3844 3669
rect 4302 3672 4308 3673
rect 4302 3668 4303 3672
rect 4307 3668 4308 3672
rect 1654 3667 1660 3668
rect 4302 3667 4308 3668
rect 4478 3672 4484 3673
rect 4478 3668 4479 3672
rect 4483 3668 4484 3672
rect 4478 3667 4484 3668
rect 4670 3672 4676 3673
rect 4670 3668 4671 3672
rect 4675 3668 4676 3672
rect 4670 3667 4676 3668
rect 4878 3672 4884 3673
rect 4878 3668 4879 3672
rect 4883 3668 4884 3672
rect 4878 3667 4884 3668
rect 5102 3672 5108 3673
rect 5102 3668 5103 3672
rect 5107 3668 5108 3672
rect 5102 3667 5108 3668
rect 5334 3672 5340 3673
rect 5334 3668 5335 3672
rect 5339 3668 5340 3672
rect 5334 3667 5340 3668
rect 5542 3672 5548 3673
rect 5542 3668 5543 3672
rect 5547 3668 5548 3672
rect 5662 3669 5663 3673
rect 5667 3669 5668 3673
rect 5662 3668 5668 3669
rect 5542 3667 5548 3668
rect 2254 3660 2260 3661
rect 1974 3659 1980 3660
rect 298 3657 304 3658
rect 110 3656 116 3657
rect 110 3652 111 3656
rect 115 3652 116 3656
rect 298 3653 299 3657
rect 303 3653 304 3657
rect 298 3652 304 3653
rect 466 3657 472 3658
rect 466 3653 467 3657
rect 471 3653 472 3657
rect 466 3652 472 3653
rect 650 3657 656 3658
rect 650 3653 651 3657
rect 655 3653 656 3657
rect 650 3652 656 3653
rect 834 3657 840 3658
rect 834 3653 835 3657
rect 839 3653 840 3657
rect 834 3652 840 3653
rect 1026 3657 1032 3658
rect 1026 3653 1027 3657
rect 1031 3653 1032 3657
rect 1026 3652 1032 3653
rect 1226 3657 1232 3658
rect 1226 3653 1227 3657
rect 1231 3653 1232 3657
rect 1226 3652 1232 3653
rect 1426 3657 1432 3658
rect 1426 3653 1427 3657
rect 1431 3653 1432 3657
rect 1426 3652 1432 3653
rect 1626 3657 1632 3658
rect 1626 3653 1627 3657
rect 1631 3653 1632 3657
rect 1626 3652 1632 3653
rect 1934 3656 1940 3657
rect 1934 3652 1935 3656
rect 1939 3652 1940 3656
rect 1974 3655 1975 3659
rect 1979 3655 1980 3659
rect 2254 3656 2255 3660
rect 2259 3656 2260 3660
rect 2254 3655 2260 3656
rect 2478 3660 2484 3661
rect 2478 3656 2479 3660
rect 2483 3656 2484 3660
rect 2478 3655 2484 3656
rect 2694 3660 2700 3661
rect 2694 3656 2695 3660
rect 2699 3656 2700 3660
rect 2694 3655 2700 3656
rect 2902 3660 2908 3661
rect 2902 3656 2903 3660
rect 2907 3656 2908 3660
rect 2902 3655 2908 3656
rect 3102 3660 3108 3661
rect 3102 3656 3103 3660
rect 3107 3656 3108 3660
rect 3102 3655 3108 3656
rect 3302 3660 3308 3661
rect 3302 3656 3303 3660
rect 3307 3656 3308 3660
rect 3302 3655 3308 3656
rect 3502 3660 3508 3661
rect 3502 3656 3503 3660
rect 3507 3656 3508 3660
rect 3502 3655 3508 3656
rect 3798 3659 3804 3660
rect 3798 3655 3799 3659
rect 3803 3655 3804 3659
rect 4274 3657 4280 3658
rect 1974 3654 1980 3655
rect 3798 3654 3804 3655
rect 3838 3656 3844 3657
rect 110 3651 116 3652
rect 1934 3651 1940 3652
rect 3838 3652 3839 3656
rect 3843 3652 3844 3656
rect 4274 3653 4275 3657
rect 4279 3653 4280 3657
rect 4274 3652 4280 3653
rect 4450 3657 4456 3658
rect 4450 3653 4451 3657
rect 4455 3653 4456 3657
rect 4450 3652 4456 3653
rect 4642 3657 4648 3658
rect 4642 3653 4643 3657
rect 4647 3653 4648 3657
rect 4642 3652 4648 3653
rect 4850 3657 4856 3658
rect 4850 3653 4851 3657
rect 4855 3653 4856 3657
rect 4850 3652 4856 3653
rect 5074 3657 5080 3658
rect 5074 3653 5075 3657
rect 5079 3653 5080 3657
rect 5074 3652 5080 3653
rect 5306 3657 5312 3658
rect 5306 3653 5307 3657
rect 5311 3653 5312 3657
rect 5306 3652 5312 3653
rect 5514 3657 5520 3658
rect 5514 3653 5515 3657
rect 5519 3653 5520 3657
rect 5514 3652 5520 3653
rect 5662 3656 5668 3657
rect 5662 3652 5663 3656
rect 5667 3652 5668 3656
rect 3838 3651 3844 3652
rect 5662 3651 5668 3652
rect 1974 3597 1980 3598
rect 3798 3597 3804 3598
rect 1974 3593 1975 3597
rect 1979 3593 1980 3597
rect 1974 3592 1980 3593
rect 2134 3596 2140 3597
rect 2134 3592 2135 3596
rect 2139 3592 2140 3596
rect 2134 3591 2140 3592
rect 2310 3596 2316 3597
rect 2310 3592 2311 3596
rect 2315 3592 2316 3596
rect 2310 3591 2316 3592
rect 2478 3596 2484 3597
rect 2478 3592 2479 3596
rect 2483 3592 2484 3596
rect 2478 3591 2484 3592
rect 2646 3596 2652 3597
rect 2646 3592 2647 3596
rect 2651 3592 2652 3596
rect 2646 3591 2652 3592
rect 2806 3596 2812 3597
rect 2806 3592 2807 3596
rect 2811 3592 2812 3596
rect 2806 3591 2812 3592
rect 2966 3596 2972 3597
rect 2966 3592 2967 3596
rect 2971 3592 2972 3596
rect 2966 3591 2972 3592
rect 3134 3596 3140 3597
rect 3134 3592 3135 3596
rect 3139 3592 3140 3596
rect 3134 3591 3140 3592
rect 3302 3596 3308 3597
rect 3302 3592 3303 3596
rect 3307 3592 3308 3596
rect 3798 3593 3799 3597
rect 3803 3593 3804 3597
rect 3798 3592 3804 3593
rect 3302 3591 3308 3592
rect 2106 3581 2112 3582
rect 1974 3580 1980 3581
rect 1974 3576 1975 3580
rect 1979 3576 1980 3580
rect 2106 3577 2107 3581
rect 2111 3577 2112 3581
rect 2106 3576 2112 3577
rect 2282 3581 2288 3582
rect 2282 3577 2283 3581
rect 2287 3577 2288 3581
rect 2282 3576 2288 3577
rect 2450 3581 2456 3582
rect 2450 3577 2451 3581
rect 2455 3577 2456 3581
rect 2450 3576 2456 3577
rect 2618 3581 2624 3582
rect 2618 3577 2619 3581
rect 2623 3577 2624 3581
rect 2618 3576 2624 3577
rect 2778 3581 2784 3582
rect 2778 3577 2779 3581
rect 2783 3577 2784 3581
rect 2778 3576 2784 3577
rect 2938 3581 2944 3582
rect 2938 3577 2939 3581
rect 2943 3577 2944 3581
rect 2938 3576 2944 3577
rect 3106 3581 3112 3582
rect 3106 3577 3107 3581
rect 3111 3577 3112 3581
rect 3106 3576 3112 3577
rect 3274 3581 3280 3582
rect 3274 3577 3275 3581
rect 3279 3577 3280 3581
rect 3274 3576 3280 3577
rect 3798 3580 3804 3581
rect 3798 3576 3799 3580
rect 3803 3576 3804 3580
rect 1974 3575 1980 3576
rect 3798 3575 3804 3576
rect 110 3504 116 3505
rect 1934 3504 1940 3505
rect 110 3500 111 3504
rect 115 3500 116 3504
rect 110 3499 116 3500
rect 202 3503 208 3504
rect 202 3499 203 3503
rect 207 3499 208 3503
rect 202 3498 208 3499
rect 378 3503 384 3504
rect 378 3499 379 3503
rect 383 3499 384 3503
rect 378 3498 384 3499
rect 562 3503 568 3504
rect 562 3499 563 3503
rect 567 3499 568 3503
rect 562 3498 568 3499
rect 754 3503 760 3504
rect 754 3499 755 3503
rect 759 3499 760 3503
rect 754 3498 760 3499
rect 954 3503 960 3504
rect 954 3499 955 3503
rect 959 3499 960 3503
rect 954 3498 960 3499
rect 1162 3503 1168 3504
rect 1162 3499 1163 3503
rect 1167 3499 1168 3503
rect 1162 3498 1168 3499
rect 1378 3503 1384 3504
rect 1378 3499 1379 3503
rect 1383 3499 1384 3503
rect 1378 3498 1384 3499
rect 1594 3503 1600 3504
rect 1594 3499 1595 3503
rect 1599 3499 1600 3503
rect 1934 3500 1935 3504
rect 1939 3500 1940 3504
rect 1934 3499 1940 3500
rect 1594 3498 1600 3499
rect 3838 3496 3844 3497
rect 5662 3496 5668 3497
rect 3838 3492 3839 3496
rect 3843 3492 3844 3496
rect 3838 3491 3844 3492
rect 4554 3495 4560 3496
rect 4554 3491 4555 3495
rect 4559 3491 4560 3495
rect 4554 3490 4560 3491
rect 4698 3495 4704 3496
rect 4698 3491 4699 3495
rect 4703 3491 4704 3495
rect 4698 3490 4704 3491
rect 4850 3495 4856 3496
rect 4850 3491 4851 3495
rect 4855 3491 4856 3495
rect 4850 3490 4856 3491
rect 5010 3495 5016 3496
rect 5010 3491 5011 3495
rect 5015 3491 5016 3495
rect 5010 3490 5016 3491
rect 5178 3495 5184 3496
rect 5178 3491 5179 3495
rect 5183 3491 5184 3495
rect 5178 3490 5184 3491
rect 5354 3495 5360 3496
rect 5354 3491 5355 3495
rect 5359 3491 5360 3495
rect 5354 3490 5360 3491
rect 5514 3495 5520 3496
rect 5514 3491 5515 3495
rect 5519 3491 5520 3495
rect 5662 3492 5663 3496
rect 5667 3492 5668 3496
rect 5662 3491 5668 3492
rect 5514 3490 5520 3491
rect 230 3488 236 3489
rect 110 3487 116 3488
rect 110 3483 111 3487
rect 115 3483 116 3487
rect 230 3484 231 3488
rect 235 3484 236 3488
rect 230 3483 236 3484
rect 406 3488 412 3489
rect 406 3484 407 3488
rect 411 3484 412 3488
rect 406 3483 412 3484
rect 590 3488 596 3489
rect 590 3484 591 3488
rect 595 3484 596 3488
rect 590 3483 596 3484
rect 782 3488 788 3489
rect 782 3484 783 3488
rect 787 3484 788 3488
rect 782 3483 788 3484
rect 982 3488 988 3489
rect 982 3484 983 3488
rect 987 3484 988 3488
rect 982 3483 988 3484
rect 1190 3488 1196 3489
rect 1190 3484 1191 3488
rect 1195 3484 1196 3488
rect 1190 3483 1196 3484
rect 1406 3488 1412 3489
rect 1406 3484 1407 3488
rect 1411 3484 1412 3488
rect 1406 3483 1412 3484
rect 1622 3488 1628 3489
rect 1622 3484 1623 3488
rect 1627 3484 1628 3488
rect 1622 3483 1628 3484
rect 1934 3487 1940 3488
rect 1934 3483 1935 3487
rect 1939 3483 1940 3487
rect 110 3482 116 3483
rect 1934 3482 1940 3483
rect 4582 3480 4588 3481
rect 3838 3479 3844 3480
rect 3838 3475 3839 3479
rect 3843 3475 3844 3479
rect 4582 3476 4583 3480
rect 4587 3476 4588 3480
rect 4582 3475 4588 3476
rect 4726 3480 4732 3481
rect 4726 3476 4727 3480
rect 4731 3476 4732 3480
rect 4726 3475 4732 3476
rect 4878 3480 4884 3481
rect 4878 3476 4879 3480
rect 4883 3476 4884 3480
rect 4878 3475 4884 3476
rect 5038 3480 5044 3481
rect 5038 3476 5039 3480
rect 5043 3476 5044 3480
rect 5038 3475 5044 3476
rect 5206 3480 5212 3481
rect 5206 3476 5207 3480
rect 5211 3476 5212 3480
rect 5206 3475 5212 3476
rect 5382 3480 5388 3481
rect 5382 3476 5383 3480
rect 5387 3476 5388 3480
rect 5382 3475 5388 3476
rect 5542 3480 5548 3481
rect 5542 3476 5543 3480
rect 5547 3476 5548 3480
rect 5542 3475 5548 3476
rect 5662 3479 5668 3480
rect 5662 3475 5663 3479
rect 5667 3475 5668 3479
rect 3838 3474 3844 3475
rect 5662 3474 5668 3475
rect 1974 3424 1980 3425
rect 3798 3424 3804 3425
rect 1974 3420 1975 3424
rect 1979 3420 1980 3424
rect 1974 3419 1980 3420
rect 2034 3423 2040 3424
rect 2034 3419 2035 3423
rect 2039 3419 2040 3423
rect 2034 3418 2040 3419
rect 2186 3423 2192 3424
rect 2186 3419 2187 3423
rect 2191 3419 2192 3423
rect 2186 3418 2192 3419
rect 2338 3423 2344 3424
rect 2338 3419 2339 3423
rect 2343 3419 2344 3423
rect 2338 3418 2344 3419
rect 2490 3423 2496 3424
rect 2490 3419 2491 3423
rect 2495 3419 2496 3423
rect 2490 3418 2496 3419
rect 2642 3423 2648 3424
rect 2642 3419 2643 3423
rect 2647 3419 2648 3423
rect 2642 3418 2648 3419
rect 2794 3423 2800 3424
rect 2794 3419 2795 3423
rect 2799 3419 2800 3423
rect 2794 3418 2800 3419
rect 2946 3423 2952 3424
rect 2946 3419 2947 3423
rect 2951 3419 2952 3423
rect 2946 3418 2952 3419
rect 3098 3423 3104 3424
rect 3098 3419 3099 3423
rect 3103 3419 3104 3423
rect 3798 3420 3799 3424
rect 3803 3420 3804 3424
rect 3798 3419 3804 3420
rect 3098 3418 3104 3419
rect 110 3409 116 3410
rect 1934 3409 1940 3410
rect 3838 3409 3844 3410
rect 5662 3409 5668 3410
rect 110 3405 111 3409
rect 115 3405 116 3409
rect 110 3404 116 3405
rect 254 3408 260 3409
rect 254 3404 255 3408
rect 259 3404 260 3408
rect 254 3403 260 3404
rect 470 3408 476 3409
rect 470 3404 471 3408
rect 475 3404 476 3408
rect 470 3403 476 3404
rect 694 3408 700 3409
rect 694 3404 695 3408
rect 699 3404 700 3408
rect 694 3403 700 3404
rect 918 3408 924 3409
rect 918 3404 919 3408
rect 923 3404 924 3408
rect 918 3403 924 3404
rect 1142 3408 1148 3409
rect 1142 3404 1143 3408
rect 1147 3404 1148 3408
rect 1142 3403 1148 3404
rect 1366 3408 1372 3409
rect 1366 3404 1367 3408
rect 1371 3404 1372 3408
rect 1366 3403 1372 3404
rect 1590 3408 1596 3409
rect 1590 3404 1591 3408
rect 1595 3404 1596 3408
rect 1934 3405 1935 3409
rect 1939 3405 1940 3409
rect 2062 3408 2068 3409
rect 1934 3404 1940 3405
rect 1974 3407 1980 3408
rect 1590 3403 1596 3404
rect 1974 3403 1975 3407
rect 1979 3403 1980 3407
rect 2062 3404 2063 3408
rect 2067 3404 2068 3408
rect 2062 3403 2068 3404
rect 2214 3408 2220 3409
rect 2214 3404 2215 3408
rect 2219 3404 2220 3408
rect 2214 3403 2220 3404
rect 2366 3408 2372 3409
rect 2366 3404 2367 3408
rect 2371 3404 2372 3408
rect 2366 3403 2372 3404
rect 2518 3408 2524 3409
rect 2518 3404 2519 3408
rect 2523 3404 2524 3408
rect 2518 3403 2524 3404
rect 2670 3408 2676 3409
rect 2670 3404 2671 3408
rect 2675 3404 2676 3408
rect 2670 3403 2676 3404
rect 2822 3408 2828 3409
rect 2822 3404 2823 3408
rect 2827 3404 2828 3408
rect 2822 3403 2828 3404
rect 2974 3408 2980 3409
rect 2974 3404 2975 3408
rect 2979 3404 2980 3408
rect 2974 3403 2980 3404
rect 3126 3408 3132 3409
rect 3126 3404 3127 3408
rect 3131 3404 3132 3408
rect 3126 3403 3132 3404
rect 3798 3407 3804 3408
rect 3798 3403 3799 3407
rect 3803 3403 3804 3407
rect 3838 3405 3839 3409
rect 3843 3405 3844 3409
rect 3838 3404 3844 3405
rect 4902 3408 4908 3409
rect 4902 3404 4903 3408
rect 4907 3404 4908 3408
rect 4902 3403 4908 3404
rect 5038 3408 5044 3409
rect 5038 3404 5039 3408
rect 5043 3404 5044 3408
rect 5038 3403 5044 3404
rect 5174 3408 5180 3409
rect 5174 3404 5175 3408
rect 5179 3404 5180 3408
rect 5174 3403 5180 3404
rect 5310 3408 5316 3409
rect 5310 3404 5311 3408
rect 5315 3404 5316 3408
rect 5310 3403 5316 3404
rect 5446 3408 5452 3409
rect 5446 3404 5447 3408
rect 5451 3404 5452 3408
rect 5662 3405 5663 3409
rect 5667 3405 5668 3409
rect 5662 3404 5668 3405
rect 5446 3403 5452 3404
rect 1974 3402 1980 3403
rect 3798 3402 3804 3403
rect 226 3393 232 3394
rect 110 3392 116 3393
rect 110 3388 111 3392
rect 115 3388 116 3392
rect 226 3389 227 3393
rect 231 3389 232 3393
rect 226 3388 232 3389
rect 442 3393 448 3394
rect 442 3389 443 3393
rect 447 3389 448 3393
rect 442 3388 448 3389
rect 666 3393 672 3394
rect 666 3389 667 3393
rect 671 3389 672 3393
rect 666 3388 672 3389
rect 890 3393 896 3394
rect 890 3389 891 3393
rect 895 3389 896 3393
rect 890 3388 896 3389
rect 1114 3393 1120 3394
rect 1114 3389 1115 3393
rect 1119 3389 1120 3393
rect 1114 3388 1120 3389
rect 1338 3393 1344 3394
rect 1338 3389 1339 3393
rect 1343 3389 1344 3393
rect 1338 3388 1344 3389
rect 1562 3393 1568 3394
rect 4874 3393 4880 3394
rect 1562 3389 1563 3393
rect 1567 3389 1568 3393
rect 1562 3388 1568 3389
rect 1934 3392 1940 3393
rect 1934 3388 1935 3392
rect 1939 3388 1940 3392
rect 110 3387 116 3388
rect 1934 3387 1940 3388
rect 3838 3392 3844 3393
rect 3838 3388 3839 3392
rect 3843 3388 3844 3392
rect 4874 3389 4875 3393
rect 4879 3389 4880 3393
rect 4874 3388 4880 3389
rect 5010 3393 5016 3394
rect 5010 3389 5011 3393
rect 5015 3389 5016 3393
rect 5010 3388 5016 3389
rect 5146 3393 5152 3394
rect 5146 3389 5147 3393
rect 5151 3389 5152 3393
rect 5146 3388 5152 3389
rect 5282 3393 5288 3394
rect 5282 3389 5283 3393
rect 5287 3389 5288 3393
rect 5282 3388 5288 3389
rect 5418 3393 5424 3394
rect 5418 3389 5419 3393
rect 5423 3389 5424 3393
rect 5418 3388 5424 3389
rect 5662 3392 5668 3393
rect 5662 3388 5663 3392
rect 5667 3388 5668 3392
rect 3838 3387 3844 3388
rect 5662 3387 5668 3388
rect 1974 3337 1980 3338
rect 3798 3337 3804 3338
rect 1974 3333 1975 3337
rect 1979 3333 1980 3337
rect 1974 3332 1980 3333
rect 2022 3336 2028 3337
rect 2022 3332 2023 3336
rect 2027 3332 2028 3336
rect 2022 3331 2028 3332
rect 2190 3336 2196 3337
rect 2190 3332 2191 3336
rect 2195 3332 2196 3336
rect 2190 3331 2196 3332
rect 2374 3336 2380 3337
rect 2374 3332 2375 3336
rect 2379 3332 2380 3336
rect 2374 3331 2380 3332
rect 2550 3336 2556 3337
rect 2550 3332 2551 3336
rect 2555 3332 2556 3336
rect 2550 3331 2556 3332
rect 2726 3336 2732 3337
rect 2726 3332 2727 3336
rect 2731 3332 2732 3336
rect 2726 3331 2732 3332
rect 2894 3336 2900 3337
rect 2894 3332 2895 3336
rect 2899 3332 2900 3336
rect 2894 3331 2900 3332
rect 3070 3336 3076 3337
rect 3070 3332 3071 3336
rect 3075 3332 3076 3336
rect 3070 3331 3076 3332
rect 3246 3336 3252 3337
rect 3246 3332 3247 3336
rect 3251 3332 3252 3336
rect 3798 3333 3799 3337
rect 3803 3333 3804 3337
rect 3798 3332 3804 3333
rect 3246 3331 3252 3332
rect 1994 3321 2000 3322
rect 1974 3320 1980 3321
rect 1974 3316 1975 3320
rect 1979 3316 1980 3320
rect 1994 3317 1995 3321
rect 1999 3317 2000 3321
rect 1994 3316 2000 3317
rect 2162 3321 2168 3322
rect 2162 3317 2163 3321
rect 2167 3317 2168 3321
rect 2162 3316 2168 3317
rect 2346 3321 2352 3322
rect 2346 3317 2347 3321
rect 2351 3317 2352 3321
rect 2346 3316 2352 3317
rect 2522 3321 2528 3322
rect 2522 3317 2523 3321
rect 2527 3317 2528 3321
rect 2522 3316 2528 3317
rect 2698 3321 2704 3322
rect 2698 3317 2699 3321
rect 2703 3317 2704 3321
rect 2698 3316 2704 3317
rect 2866 3321 2872 3322
rect 2866 3317 2867 3321
rect 2871 3317 2872 3321
rect 2866 3316 2872 3317
rect 3042 3321 3048 3322
rect 3042 3317 3043 3321
rect 3047 3317 3048 3321
rect 3042 3316 3048 3317
rect 3218 3321 3224 3322
rect 3218 3317 3219 3321
rect 3223 3317 3224 3321
rect 3218 3316 3224 3317
rect 3798 3320 3804 3321
rect 3798 3316 3799 3320
rect 3803 3316 3804 3320
rect 1974 3315 1980 3316
rect 3798 3315 3804 3316
rect 3838 3260 3844 3261
rect 5662 3260 5668 3261
rect 3838 3256 3839 3260
rect 3843 3256 3844 3260
rect 3838 3255 3844 3256
rect 4698 3259 4704 3260
rect 4698 3255 4699 3259
rect 4703 3255 4704 3259
rect 4698 3254 4704 3255
rect 4834 3259 4840 3260
rect 4834 3255 4835 3259
rect 4839 3255 4840 3259
rect 4834 3254 4840 3255
rect 4970 3259 4976 3260
rect 4970 3255 4971 3259
rect 4975 3255 4976 3259
rect 4970 3254 4976 3255
rect 5106 3259 5112 3260
rect 5106 3255 5107 3259
rect 5111 3255 5112 3259
rect 5106 3254 5112 3255
rect 5242 3259 5248 3260
rect 5242 3255 5243 3259
rect 5247 3255 5248 3259
rect 5242 3254 5248 3255
rect 5378 3259 5384 3260
rect 5378 3255 5379 3259
rect 5383 3255 5384 3259
rect 5378 3254 5384 3255
rect 5514 3259 5520 3260
rect 5514 3255 5515 3259
rect 5519 3255 5520 3259
rect 5662 3256 5663 3260
rect 5667 3256 5668 3260
rect 5662 3255 5668 3256
rect 5514 3254 5520 3255
rect 110 3244 116 3245
rect 1934 3244 1940 3245
rect 4726 3244 4732 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 110 3239 116 3240
rect 210 3243 216 3244
rect 210 3239 211 3243
rect 215 3239 216 3243
rect 210 3238 216 3239
rect 418 3243 424 3244
rect 418 3239 419 3243
rect 423 3239 424 3243
rect 418 3238 424 3239
rect 634 3243 640 3244
rect 634 3239 635 3243
rect 639 3239 640 3243
rect 634 3238 640 3239
rect 850 3243 856 3244
rect 850 3239 851 3243
rect 855 3239 856 3243
rect 850 3238 856 3239
rect 1074 3243 1080 3244
rect 1074 3239 1075 3243
rect 1079 3239 1080 3243
rect 1074 3238 1080 3239
rect 1298 3243 1304 3244
rect 1298 3239 1299 3243
rect 1303 3239 1304 3243
rect 1298 3238 1304 3239
rect 1522 3243 1528 3244
rect 1522 3239 1523 3243
rect 1527 3239 1528 3243
rect 1934 3240 1935 3244
rect 1939 3240 1940 3244
rect 1934 3239 1940 3240
rect 3838 3243 3844 3244
rect 3838 3239 3839 3243
rect 3843 3239 3844 3243
rect 4726 3240 4727 3244
rect 4731 3240 4732 3244
rect 4726 3239 4732 3240
rect 4862 3244 4868 3245
rect 4862 3240 4863 3244
rect 4867 3240 4868 3244
rect 4862 3239 4868 3240
rect 4998 3244 5004 3245
rect 4998 3240 4999 3244
rect 5003 3240 5004 3244
rect 4998 3239 5004 3240
rect 5134 3244 5140 3245
rect 5134 3240 5135 3244
rect 5139 3240 5140 3244
rect 5134 3239 5140 3240
rect 5270 3244 5276 3245
rect 5270 3240 5271 3244
rect 5275 3240 5276 3244
rect 5270 3239 5276 3240
rect 5406 3244 5412 3245
rect 5406 3240 5407 3244
rect 5411 3240 5412 3244
rect 5406 3239 5412 3240
rect 5542 3244 5548 3245
rect 5542 3240 5543 3244
rect 5547 3240 5548 3244
rect 5542 3239 5548 3240
rect 5662 3243 5668 3244
rect 5662 3239 5663 3243
rect 5667 3239 5668 3243
rect 1522 3238 1528 3239
rect 3838 3238 3844 3239
rect 5662 3238 5668 3239
rect 238 3228 244 3229
rect 110 3227 116 3228
rect 110 3223 111 3227
rect 115 3223 116 3227
rect 238 3224 239 3228
rect 243 3224 244 3228
rect 238 3223 244 3224
rect 446 3228 452 3229
rect 446 3224 447 3228
rect 451 3224 452 3228
rect 446 3223 452 3224
rect 662 3228 668 3229
rect 662 3224 663 3228
rect 667 3224 668 3228
rect 662 3223 668 3224
rect 878 3228 884 3229
rect 878 3224 879 3228
rect 883 3224 884 3228
rect 878 3223 884 3224
rect 1102 3228 1108 3229
rect 1102 3224 1103 3228
rect 1107 3224 1108 3228
rect 1102 3223 1108 3224
rect 1326 3228 1332 3229
rect 1326 3224 1327 3228
rect 1331 3224 1332 3228
rect 1326 3223 1332 3224
rect 1550 3228 1556 3229
rect 1550 3224 1551 3228
rect 1555 3224 1556 3228
rect 1550 3223 1556 3224
rect 1934 3227 1940 3228
rect 1934 3223 1935 3227
rect 1939 3223 1940 3227
rect 110 3222 116 3223
rect 1934 3222 1940 3223
rect 1974 3184 1980 3185
rect 3798 3184 3804 3185
rect 1974 3180 1975 3184
rect 1979 3180 1980 3184
rect 1974 3179 1980 3180
rect 1994 3183 2000 3184
rect 1994 3179 1995 3183
rect 1999 3179 2000 3183
rect 1994 3178 2000 3179
rect 2210 3183 2216 3184
rect 2210 3179 2211 3183
rect 2215 3179 2216 3183
rect 2210 3178 2216 3179
rect 2434 3183 2440 3184
rect 2434 3179 2435 3183
rect 2439 3179 2440 3183
rect 2434 3178 2440 3179
rect 2650 3183 2656 3184
rect 2650 3179 2651 3183
rect 2655 3179 2656 3183
rect 2650 3178 2656 3179
rect 2850 3183 2856 3184
rect 2850 3179 2851 3183
rect 2855 3179 2856 3183
rect 2850 3178 2856 3179
rect 3050 3183 3056 3184
rect 3050 3179 3051 3183
rect 3055 3179 3056 3183
rect 3050 3178 3056 3179
rect 3250 3183 3256 3184
rect 3250 3179 3251 3183
rect 3255 3179 3256 3183
rect 3250 3178 3256 3179
rect 3450 3183 3456 3184
rect 3450 3179 3451 3183
rect 3455 3179 3456 3183
rect 3798 3180 3799 3184
rect 3803 3180 3804 3184
rect 3798 3179 3804 3180
rect 3450 3178 3456 3179
rect 3838 3177 3844 3178
rect 5662 3177 5668 3178
rect 3838 3173 3839 3177
rect 3843 3173 3844 3177
rect 3838 3172 3844 3173
rect 4566 3176 4572 3177
rect 4566 3172 4567 3176
rect 4571 3172 4572 3176
rect 4566 3171 4572 3172
rect 4742 3176 4748 3177
rect 4742 3172 4743 3176
rect 4747 3172 4748 3176
rect 4742 3171 4748 3172
rect 4934 3176 4940 3177
rect 4934 3172 4935 3176
rect 4939 3172 4940 3176
rect 4934 3171 4940 3172
rect 5134 3176 5140 3177
rect 5134 3172 5135 3176
rect 5139 3172 5140 3176
rect 5134 3171 5140 3172
rect 5350 3176 5356 3177
rect 5350 3172 5351 3176
rect 5355 3172 5356 3176
rect 5350 3171 5356 3172
rect 5542 3176 5548 3177
rect 5542 3172 5543 3176
rect 5547 3172 5548 3176
rect 5662 3173 5663 3177
rect 5667 3173 5668 3177
rect 5662 3172 5668 3173
rect 5542 3171 5548 3172
rect 2022 3168 2028 3169
rect 1974 3167 1980 3168
rect 1974 3163 1975 3167
rect 1979 3163 1980 3167
rect 2022 3164 2023 3168
rect 2027 3164 2028 3168
rect 2022 3163 2028 3164
rect 2238 3168 2244 3169
rect 2238 3164 2239 3168
rect 2243 3164 2244 3168
rect 2238 3163 2244 3164
rect 2462 3168 2468 3169
rect 2462 3164 2463 3168
rect 2467 3164 2468 3168
rect 2462 3163 2468 3164
rect 2678 3168 2684 3169
rect 2678 3164 2679 3168
rect 2683 3164 2684 3168
rect 2678 3163 2684 3164
rect 2878 3168 2884 3169
rect 2878 3164 2879 3168
rect 2883 3164 2884 3168
rect 2878 3163 2884 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3278 3168 3284 3169
rect 3278 3164 3279 3168
rect 3283 3164 3284 3168
rect 3278 3163 3284 3164
rect 3478 3168 3484 3169
rect 3478 3164 3479 3168
rect 3483 3164 3484 3168
rect 3478 3163 3484 3164
rect 3798 3167 3804 3168
rect 3798 3163 3799 3167
rect 3803 3163 3804 3167
rect 1974 3162 1980 3163
rect 3798 3162 3804 3163
rect 4538 3161 4544 3162
rect 3838 3160 3844 3161
rect 3838 3156 3839 3160
rect 3843 3156 3844 3160
rect 4538 3157 4539 3161
rect 4543 3157 4544 3161
rect 4538 3156 4544 3157
rect 4714 3161 4720 3162
rect 4714 3157 4715 3161
rect 4719 3157 4720 3161
rect 4714 3156 4720 3157
rect 4906 3161 4912 3162
rect 4906 3157 4907 3161
rect 4911 3157 4912 3161
rect 4906 3156 4912 3157
rect 5106 3161 5112 3162
rect 5106 3157 5107 3161
rect 5111 3157 5112 3161
rect 5106 3156 5112 3157
rect 5322 3161 5328 3162
rect 5322 3157 5323 3161
rect 5327 3157 5328 3161
rect 5322 3156 5328 3157
rect 5514 3161 5520 3162
rect 5514 3157 5515 3161
rect 5519 3157 5520 3161
rect 5514 3156 5520 3157
rect 5662 3160 5668 3161
rect 5662 3156 5663 3160
rect 5667 3156 5668 3160
rect 3838 3155 3844 3156
rect 5662 3155 5668 3156
rect 110 3153 116 3154
rect 1934 3153 1940 3154
rect 110 3149 111 3153
rect 115 3149 116 3153
rect 110 3148 116 3149
rect 302 3152 308 3153
rect 302 3148 303 3152
rect 307 3148 308 3152
rect 302 3147 308 3148
rect 542 3152 548 3153
rect 542 3148 543 3152
rect 547 3148 548 3152
rect 542 3147 548 3148
rect 782 3152 788 3153
rect 782 3148 783 3152
rect 787 3148 788 3152
rect 782 3147 788 3148
rect 1022 3152 1028 3153
rect 1022 3148 1023 3152
rect 1027 3148 1028 3152
rect 1022 3147 1028 3148
rect 1262 3152 1268 3153
rect 1262 3148 1263 3152
rect 1267 3148 1268 3152
rect 1262 3147 1268 3148
rect 1510 3152 1516 3153
rect 1510 3148 1511 3152
rect 1515 3148 1516 3152
rect 1934 3149 1935 3153
rect 1939 3149 1940 3153
rect 1934 3148 1940 3149
rect 1510 3147 1516 3148
rect 274 3137 280 3138
rect 110 3136 116 3137
rect 110 3132 111 3136
rect 115 3132 116 3136
rect 274 3133 275 3137
rect 279 3133 280 3137
rect 274 3132 280 3133
rect 514 3137 520 3138
rect 514 3133 515 3137
rect 519 3133 520 3137
rect 514 3132 520 3133
rect 754 3137 760 3138
rect 754 3133 755 3137
rect 759 3133 760 3137
rect 754 3132 760 3133
rect 994 3137 1000 3138
rect 994 3133 995 3137
rect 999 3133 1000 3137
rect 994 3132 1000 3133
rect 1234 3137 1240 3138
rect 1234 3133 1235 3137
rect 1239 3133 1240 3137
rect 1234 3132 1240 3133
rect 1482 3137 1488 3138
rect 1482 3133 1483 3137
rect 1487 3133 1488 3137
rect 1482 3132 1488 3133
rect 1934 3136 1940 3137
rect 1934 3132 1935 3136
rect 1939 3132 1940 3136
rect 110 3131 116 3132
rect 1934 3131 1940 3132
rect 1974 3109 1980 3110
rect 3798 3109 3804 3110
rect 1974 3105 1975 3109
rect 1979 3105 1980 3109
rect 1974 3104 1980 3105
rect 2022 3108 2028 3109
rect 2022 3104 2023 3108
rect 2027 3104 2028 3108
rect 2022 3103 2028 3104
rect 2326 3108 2332 3109
rect 2326 3104 2327 3108
rect 2331 3104 2332 3108
rect 2326 3103 2332 3104
rect 2630 3108 2636 3109
rect 2630 3104 2631 3108
rect 2635 3104 2636 3108
rect 2630 3103 2636 3104
rect 2910 3108 2916 3109
rect 2910 3104 2911 3108
rect 2915 3104 2916 3108
rect 2910 3103 2916 3104
rect 3174 3108 3180 3109
rect 3174 3104 3175 3108
rect 3179 3104 3180 3108
rect 3174 3103 3180 3104
rect 3438 3108 3444 3109
rect 3438 3104 3439 3108
rect 3443 3104 3444 3108
rect 3438 3103 3444 3104
rect 3678 3108 3684 3109
rect 3678 3104 3679 3108
rect 3683 3104 3684 3108
rect 3798 3105 3799 3109
rect 3803 3105 3804 3109
rect 3798 3104 3804 3105
rect 3678 3103 3684 3104
rect 1994 3093 2000 3094
rect 1974 3092 1980 3093
rect 1974 3088 1975 3092
rect 1979 3088 1980 3092
rect 1994 3089 1995 3093
rect 1999 3089 2000 3093
rect 1994 3088 2000 3089
rect 2298 3093 2304 3094
rect 2298 3089 2299 3093
rect 2303 3089 2304 3093
rect 2298 3088 2304 3089
rect 2602 3093 2608 3094
rect 2602 3089 2603 3093
rect 2607 3089 2608 3093
rect 2602 3088 2608 3089
rect 2882 3093 2888 3094
rect 2882 3089 2883 3093
rect 2887 3089 2888 3093
rect 2882 3088 2888 3089
rect 3146 3093 3152 3094
rect 3146 3089 3147 3093
rect 3151 3089 3152 3093
rect 3146 3088 3152 3089
rect 3410 3093 3416 3094
rect 3410 3089 3411 3093
rect 3415 3089 3416 3093
rect 3410 3088 3416 3089
rect 3650 3093 3656 3094
rect 3650 3089 3651 3093
rect 3655 3089 3656 3093
rect 3650 3088 3656 3089
rect 3798 3092 3804 3093
rect 3798 3088 3799 3092
rect 3803 3088 3804 3092
rect 1974 3087 1980 3088
rect 3798 3087 3804 3088
rect 3838 3024 3844 3025
rect 5662 3024 5668 3025
rect 3838 3020 3839 3024
rect 3843 3020 3844 3024
rect 3838 3019 3844 3020
rect 4306 3023 4312 3024
rect 4306 3019 4307 3023
rect 4311 3019 4312 3023
rect 4306 3018 4312 3019
rect 4482 3023 4488 3024
rect 4482 3019 4483 3023
rect 4487 3019 4488 3023
rect 4482 3018 4488 3019
rect 4674 3023 4680 3024
rect 4674 3019 4675 3023
rect 4679 3019 4680 3023
rect 4674 3018 4680 3019
rect 4874 3023 4880 3024
rect 4874 3019 4875 3023
rect 4879 3019 4880 3023
rect 4874 3018 4880 3019
rect 5090 3023 5096 3024
rect 5090 3019 5091 3023
rect 5095 3019 5096 3023
rect 5090 3018 5096 3019
rect 5314 3023 5320 3024
rect 5314 3019 5315 3023
rect 5319 3019 5320 3023
rect 5314 3018 5320 3019
rect 5514 3023 5520 3024
rect 5514 3019 5515 3023
rect 5519 3019 5520 3023
rect 5662 3020 5663 3024
rect 5667 3020 5668 3024
rect 5662 3019 5668 3020
rect 5514 3018 5520 3019
rect 4334 3008 4340 3009
rect 3838 3007 3844 3008
rect 110 3004 116 3005
rect 1934 3004 1940 3005
rect 110 3000 111 3004
rect 115 3000 116 3004
rect 110 2999 116 3000
rect 354 3003 360 3004
rect 354 2999 355 3003
rect 359 2999 360 3003
rect 354 2998 360 2999
rect 626 3003 632 3004
rect 626 2999 627 3003
rect 631 2999 632 3003
rect 626 2998 632 2999
rect 882 3003 888 3004
rect 882 2999 883 3003
rect 887 2999 888 3003
rect 882 2998 888 2999
rect 1122 3003 1128 3004
rect 1122 2999 1123 3003
rect 1127 2999 1128 3003
rect 1122 2998 1128 2999
rect 1354 3003 1360 3004
rect 1354 2999 1355 3003
rect 1359 2999 1360 3003
rect 1354 2998 1360 2999
rect 1578 3003 1584 3004
rect 1578 2999 1579 3003
rect 1583 2999 1584 3003
rect 1578 2998 1584 2999
rect 1786 3003 1792 3004
rect 1786 2999 1787 3003
rect 1791 2999 1792 3003
rect 1934 3000 1935 3004
rect 1939 3000 1940 3004
rect 3838 3003 3839 3007
rect 3843 3003 3844 3007
rect 4334 3004 4335 3008
rect 4339 3004 4340 3008
rect 4334 3003 4340 3004
rect 4510 3008 4516 3009
rect 4510 3004 4511 3008
rect 4515 3004 4516 3008
rect 4510 3003 4516 3004
rect 4702 3008 4708 3009
rect 4702 3004 4703 3008
rect 4707 3004 4708 3008
rect 4702 3003 4708 3004
rect 4902 3008 4908 3009
rect 4902 3004 4903 3008
rect 4907 3004 4908 3008
rect 4902 3003 4908 3004
rect 5118 3008 5124 3009
rect 5118 3004 5119 3008
rect 5123 3004 5124 3008
rect 5118 3003 5124 3004
rect 5342 3008 5348 3009
rect 5342 3004 5343 3008
rect 5347 3004 5348 3008
rect 5342 3003 5348 3004
rect 5542 3008 5548 3009
rect 5542 3004 5543 3008
rect 5547 3004 5548 3008
rect 5542 3003 5548 3004
rect 5662 3007 5668 3008
rect 5662 3003 5663 3007
rect 5667 3003 5668 3007
rect 3838 3002 3844 3003
rect 5662 3002 5668 3003
rect 1934 2999 1940 3000
rect 1786 2998 1792 2999
rect 382 2988 388 2989
rect 110 2987 116 2988
rect 110 2983 111 2987
rect 115 2983 116 2987
rect 382 2984 383 2988
rect 387 2984 388 2988
rect 382 2983 388 2984
rect 654 2988 660 2989
rect 654 2984 655 2988
rect 659 2984 660 2988
rect 654 2983 660 2984
rect 910 2988 916 2989
rect 910 2984 911 2988
rect 915 2984 916 2988
rect 910 2983 916 2984
rect 1150 2988 1156 2989
rect 1150 2984 1151 2988
rect 1155 2984 1156 2988
rect 1150 2983 1156 2984
rect 1382 2988 1388 2989
rect 1382 2984 1383 2988
rect 1387 2984 1388 2988
rect 1382 2983 1388 2984
rect 1606 2988 1612 2989
rect 1606 2984 1607 2988
rect 1611 2984 1612 2988
rect 1606 2983 1612 2984
rect 1814 2988 1820 2989
rect 1814 2984 1815 2988
rect 1819 2984 1820 2988
rect 1814 2983 1820 2984
rect 1934 2987 1940 2988
rect 1934 2983 1935 2987
rect 1939 2983 1940 2987
rect 110 2982 116 2983
rect 1934 2982 1940 2983
rect 1974 2952 1980 2953
rect 3798 2952 3804 2953
rect 1974 2948 1975 2952
rect 1979 2948 1980 2952
rect 1974 2947 1980 2948
rect 3106 2951 3112 2952
rect 3106 2947 3107 2951
rect 3111 2947 3112 2951
rect 3106 2946 3112 2947
rect 3242 2951 3248 2952
rect 3242 2947 3243 2951
rect 3247 2947 3248 2951
rect 3242 2946 3248 2947
rect 3378 2951 3384 2952
rect 3378 2947 3379 2951
rect 3383 2947 3384 2951
rect 3378 2946 3384 2947
rect 3514 2951 3520 2952
rect 3514 2947 3515 2951
rect 3519 2947 3520 2951
rect 3514 2946 3520 2947
rect 3650 2951 3656 2952
rect 3650 2947 3651 2951
rect 3655 2947 3656 2951
rect 3798 2948 3799 2952
rect 3803 2948 3804 2952
rect 3798 2947 3804 2948
rect 3650 2946 3656 2947
rect 3838 2945 3844 2946
rect 5662 2945 5668 2946
rect 3838 2941 3839 2945
rect 3843 2941 3844 2945
rect 3838 2940 3844 2941
rect 3886 2944 3892 2945
rect 3886 2940 3887 2944
rect 3891 2940 3892 2944
rect 3886 2939 3892 2940
rect 4022 2944 4028 2945
rect 4022 2940 4023 2944
rect 4027 2940 4028 2944
rect 4022 2939 4028 2940
rect 4174 2944 4180 2945
rect 4174 2940 4175 2944
rect 4179 2940 4180 2944
rect 4174 2939 4180 2940
rect 4390 2944 4396 2945
rect 4390 2940 4391 2944
rect 4395 2940 4396 2944
rect 4390 2939 4396 2940
rect 4638 2944 4644 2945
rect 4638 2940 4639 2944
rect 4643 2940 4644 2944
rect 4638 2939 4644 2940
rect 4918 2944 4924 2945
rect 4918 2940 4919 2944
rect 4923 2940 4924 2944
rect 4918 2939 4924 2940
rect 5222 2944 5228 2945
rect 5222 2940 5223 2944
rect 5227 2940 5228 2944
rect 5222 2939 5228 2940
rect 5526 2944 5532 2945
rect 5526 2940 5527 2944
rect 5531 2940 5532 2944
rect 5662 2941 5663 2945
rect 5667 2941 5668 2945
rect 5662 2940 5668 2941
rect 5526 2939 5532 2940
rect 3134 2936 3140 2937
rect 1974 2935 1980 2936
rect 1974 2931 1975 2935
rect 1979 2931 1980 2935
rect 3134 2932 3135 2936
rect 3139 2932 3140 2936
rect 3134 2931 3140 2932
rect 3270 2936 3276 2937
rect 3270 2932 3271 2936
rect 3275 2932 3276 2936
rect 3270 2931 3276 2932
rect 3406 2936 3412 2937
rect 3406 2932 3407 2936
rect 3411 2932 3412 2936
rect 3406 2931 3412 2932
rect 3542 2936 3548 2937
rect 3542 2932 3543 2936
rect 3547 2932 3548 2936
rect 3542 2931 3548 2932
rect 3678 2936 3684 2937
rect 3678 2932 3679 2936
rect 3683 2932 3684 2936
rect 3678 2931 3684 2932
rect 3798 2935 3804 2936
rect 3798 2931 3799 2935
rect 3803 2931 3804 2935
rect 1974 2930 1980 2931
rect 3798 2930 3804 2931
rect 110 2929 116 2930
rect 1934 2929 1940 2930
rect 3858 2929 3864 2930
rect 110 2925 111 2929
rect 115 2925 116 2929
rect 110 2924 116 2925
rect 342 2928 348 2929
rect 342 2924 343 2928
rect 347 2924 348 2928
rect 342 2923 348 2924
rect 550 2928 556 2929
rect 550 2924 551 2928
rect 555 2924 556 2928
rect 550 2923 556 2924
rect 758 2928 764 2929
rect 758 2924 759 2928
rect 763 2924 764 2928
rect 758 2923 764 2924
rect 950 2928 956 2929
rect 950 2924 951 2928
rect 955 2924 956 2928
rect 950 2923 956 2924
rect 1134 2928 1140 2929
rect 1134 2924 1135 2928
rect 1139 2924 1140 2928
rect 1134 2923 1140 2924
rect 1310 2928 1316 2929
rect 1310 2924 1311 2928
rect 1315 2924 1316 2928
rect 1310 2923 1316 2924
rect 1486 2928 1492 2929
rect 1486 2924 1487 2928
rect 1491 2924 1492 2928
rect 1486 2923 1492 2924
rect 1662 2928 1668 2929
rect 1662 2924 1663 2928
rect 1667 2924 1668 2928
rect 1662 2923 1668 2924
rect 1814 2928 1820 2929
rect 1814 2924 1815 2928
rect 1819 2924 1820 2928
rect 1934 2925 1935 2929
rect 1939 2925 1940 2929
rect 1934 2924 1940 2925
rect 3838 2928 3844 2929
rect 3838 2924 3839 2928
rect 3843 2924 3844 2928
rect 3858 2925 3859 2929
rect 3863 2925 3864 2929
rect 3858 2924 3864 2925
rect 3994 2929 4000 2930
rect 3994 2925 3995 2929
rect 3999 2925 4000 2929
rect 3994 2924 4000 2925
rect 4146 2929 4152 2930
rect 4146 2925 4147 2929
rect 4151 2925 4152 2929
rect 4146 2924 4152 2925
rect 4362 2929 4368 2930
rect 4362 2925 4363 2929
rect 4367 2925 4368 2929
rect 4362 2924 4368 2925
rect 4610 2929 4616 2930
rect 4610 2925 4611 2929
rect 4615 2925 4616 2929
rect 4610 2924 4616 2925
rect 4890 2929 4896 2930
rect 4890 2925 4891 2929
rect 4895 2925 4896 2929
rect 4890 2924 4896 2925
rect 5194 2929 5200 2930
rect 5194 2925 5195 2929
rect 5199 2925 5200 2929
rect 5194 2924 5200 2925
rect 5498 2929 5504 2930
rect 5498 2925 5499 2929
rect 5503 2925 5504 2929
rect 5498 2924 5504 2925
rect 5662 2928 5668 2929
rect 5662 2924 5663 2928
rect 5667 2924 5668 2928
rect 1814 2923 1820 2924
rect 3838 2923 3844 2924
rect 5662 2923 5668 2924
rect 314 2913 320 2914
rect 110 2912 116 2913
rect 110 2908 111 2912
rect 115 2908 116 2912
rect 314 2909 315 2913
rect 319 2909 320 2913
rect 314 2908 320 2909
rect 522 2913 528 2914
rect 522 2909 523 2913
rect 527 2909 528 2913
rect 522 2908 528 2909
rect 730 2913 736 2914
rect 730 2909 731 2913
rect 735 2909 736 2913
rect 730 2908 736 2909
rect 922 2913 928 2914
rect 922 2909 923 2913
rect 927 2909 928 2913
rect 922 2908 928 2909
rect 1106 2913 1112 2914
rect 1106 2909 1107 2913
rect 1111 2909 1112 2913
rect 1106 2908 1112 2909
rect 1282 2913 1288 2914
rect 1282 2909 1283 2913
rect 1287 2909 1288 2913
rect 1282 2908 1288 2909
rect 1458 2913 1464 2914
rect 1458 2909 1459 2913
rect 1463 2909 1464 2913
rect 1458 2908 1464 2909
rect 1634 2913 1640 2914
rect 1634 2909 1635 2913
rect 1639 2909 1640 2913
rect 1634 2908 1640 2909
rect 1786 2913 1792 2914
rect 1786 2909 1787 2913
rect 1791 2909 1792 2913
rect 1786 2908 1792 2909
rect 1934 2912 1940 2913
rect 1934 2908 1935 2912
rect 1939 2908 1940 2912
rect 110 2907 116 2908
rect 1934 2907 1940 2908
rect 3838 2796 3844 2797
rect 5662 2796 5668 2797
rect 3838 2792 3839 2796
rect 3843 2792 3844 2796
rect 3838 2791 3844 2792
rect 3858 2795 3864 2796
rect 3858 2791 3859 2795
rect 3863 2791 3864 2795
rect 3858 2790 3864 2791
rect 3994 2795 4000 2796
rect 3994 2791 3995 2795
rect 3999 2791 4000 2795
rect 3994 2790 4000 2791
rect 4130 2795 4136 2796
rect 4130 2791 4131 2795
rect 4135 2791 4136 2795
rect 4130 2790 4136 2791
rect 4266 2795 4272 2796
rect 4266 2791 4267 2795
rect 4271 2791 4272 2795
rect 4266 2790 4272 2791
rect 4402 2795 4408 2796
rect 4402 2791 4403 2795
rect 4407 2791 4408 2795
rect 4402 2790 4408 2791
rect 4538 2795 4544 2796
rect 4538 2791 4539 2795
rect 4543 2791 4544 2795
rect 4538 2790 4544 2791
rect 4674 2795 4680 2796
rect 4674 2791 4675 2795
rect 4679 2791 4680 2795
rect 4674 2790 4680 2791
rect 4810 2795 4816 2796
rect 4810 2791 4811 2795
rect 4815 2791 4816 2795
rect 5662 2792 5663 2796
rect 5667 2792 5668 2796
rect 5662 2791 5668 2792
rect 4810 2790 4816 2791
rect 3886 2780 3892 2781
rect 3838 2779 3844 2780
rect 3838 2775 3839 2779
rect 3843 2775 3844 2779
rect 3886 2776 3887 2780
rect 3891 2776 3892 2780
rect 3886 2775 3892 2776
rect 4022 2780 4028 2781
rect 4022 2776 4023 2780
rect 4027 2776 4028 2780
rect 4022 2775 4028 2776
rect 4158 2780 4164 2781
rect 4158 2776 4159 2780
rect 4163 2776 4164 2780
rect 4158 2775 4164 2776
rect 4294 2780 4300 2781
rect 4294 2776 4295 2780
rect 4299 2776 4300 2780
rect 4294 2775 4300 2776
rect 4430 2780 4436 2781
rect 4430 2776 4431 2780
rect 4435 2776 4436 2780
rect 4430 2775 4436 2776
rect 4566 2780 4572 2781
rect 4566 2776 4567 2780
rect 4571 2776 4572 2780
rect 4566 2775 4572 2776
rect 4702 2780 4708 2781
rect 4702 2776 4703 2780
rect 4707 2776 4708 2780
rect 4702 2775 4708 2776
rect 4838 2780 4844 2781
rect 4838 2776 4839 2780
rect 4843 2776 4844 2780
rect 4838 2775 4844 2776
rect 5662 2779 5668 2780
rect 5662 2775 5663 2779
rect 5667 2775 5668 2779
rect 3838 2774 3844 2775
rect 5662 2774 5668 2775
rect 110 2768 116 2769
rect 1934 2768 1940 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 362 2767 368 2768
rect 362 2763 363 2767
rect 367 2763 368 2767
rect 362 2762 368 2763
rect 562 2767 568 2768
rect 562 2763 563 2767
rect 567 2763 568 2767
rect 562 2762 568 2763
rect 754 2767 760 2768
rect 754 2763 755 2767
rect 759 2763 760 2767
rect 754 2762 760 2763
rect 938 2767 944 2768
rect 938 2763 939 2767
rect 943 2763 944 2767
rect 938 2762 944 2763
rect 1114 2767 1120 2768
rect 1114 2763 1115 2767
rect 1119 2763 1120 2767
rect 1114 2762 1120 2763
rect 1282 2767 1288 2768
rect 1282 2763 1283 2767
rect 1287 2763 1288 2767
rect 1282 2762 1288 2763
rect 1450 2767 1456 2768
rect 1450 2763 1451 2767
rect 1455 2763 1456 2767
rect 1450 2762 1456 2763
rect 1618 2767 1624 2768
rect 1618 2763 1619 2767
rect 1623 2763 1624 2767
rect 1618 2762 1624 2763
rect 1786 2767 1792 2768
rect 1786 2763 1787 2767
rect 1791 2763 1792 2767
rect 1934 2764 1935 2768
rect 1939 2764 1940 2768
rect 1934 2763 1940 2764
rect 1786 2762 1792 2763
rect 390 2752 396 2753
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 590 2752 596 2753
rect 590 2748 591 2752
rect 595 2748 596 2752
rect 590 2747 596 2748
rect 782 2752 788 2753
rect 782 2748 783 2752
rect 787 2748 788 2752
rect 782 2747 788 2748
rect 966 2752 972 2753
rect 966 2748 967 2752
rect 971 2748 972 2752
rect 966 2747 972 2748
rect 1142 2752 1148 2753
rect 1142 2748 1143 2752
rect 1147 2748 1148 2752
rect 1142 2747 1148 2748
rect 1310 2752 1316 2753
rect 1310 2748 1311 2752
rect 1315 2748 1316 2752
rect 1310 2747 1316 2748
rect 1478 2752 1484 2753
rect 1478 2748 1479 2752
rect 1483 2748 1484 2752
rect 1478 2747 1484 2748
rect 1646 2752 1652 2753
rect 1646 2748 1647 2752
rect 1651 2748 1652 2752
rect 1646 2747 1652 2748
rect 1814 2752 1820 2753
rect 1814 2748 1815 2752
rect 1819 2748 1820 2752
rect 1814 2747 1820 2748
rect 1934 2751 1940 2752
rect 1934 2747 1935 2751
rect 1939 2747 1940 2751
rect 110 2746 116 2747
rect 1934 2746 1940 2747
rect 3838 2705 3844 2706
rect 5662 2705 5668 2706
rect 3838 2701 3839 2705
rect 3843 2701 3844 2705
rect 3838 2700 3844 2701
rect 3886 2704 3892 2705
rect 3886 2700 3887 2704
rect 3891 2700 3892 2704
rect 3886 2699 3892 2700
rect 4022 2704 4028 2705
rect 4022 2700 4023 2704
rect 4027 2700 4028 2704
rect 4022 2699 4028 2700
rect 4158 2704 4164 2705
rect 4158 2700 4159 2704
rect 4163 2700 4164 2704
rect 4158 2699 4164 2700
rect 4294 2704 4300 2705
rect 4294 2700 4295 2704
rect 4299 2700 4300 2704
rect 4294 2699 4300 2700
rect 4430 2704 4436 2705
rect 4430 2700 4431 2704
rect 4435 2700 4436 2704
rect 4430 2699 4436 2700
rect 4566 2704 4572 2705
rect 4566 2700 4567 2704
rect 4571 2700 4572 2704
rect 4566 2699 4572 2700
rect 4710 2704 4716 2705
rect 4710 2700 4711 2704
rect 4715 2700 4716 2704
rect 4710 2699 4716 2700
rect 4878 2704 4884 2705
rect 4878 2700 4879 2704
rect 4883 2700 4884 2704
rect 4878 2699 4884 2700
rect 5062 2704 5068 2705
rect 5062 2700 5063 2704
rect 5067 2700 5068 2704
rect 5062 2699 5068 2700
rect 5254 2704 5260 2705
rect 5254 2700 5255 2704
rect 5259 2700 5260 2704
rect 5254 2699 5260 2700
rect 5446 2704 5452 2705
rect 5446 2700 5447 2704
rect 5451 2700 5452 2704
rect 5662 2701 5663 2705
rect 5667 2701 5668 2705
rect 5662 2700 5668 2701
rect 5446 2699 5452 2700
rect 110 2689 116 2690
rect 1934 2689 1940 2690
rect 3858 2689 3864 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 110 2684 116 2685
rect 446 2688 452 2689
rect 446 2684 447 2688
rect 451 2684 452 2688
rect 446 2683 452 2684
rect 614 2688 620 2689
rect 614 2684 615 2688
rect 619 2684 620 2688
rect 614 2683 620 2684
rect 774 2688 780 2689
rect 774 2684 775 2688
rect 779 2684 780 2688
rect 774 2683 780 2684
rect 934 2688 940 2689
rect 934 2684 935 2688
rect 939 2684 940 2688
rect 934 2683 940 2684
rect 1086 2688 1092 2689
rect 1086 2684 1087 2688
rect 1091 2684 1092 2688
rect 1086 2683 1092 2684
rect 1238 2688 1244 2689
rect 1238 2684 1239 2688
rect 1243 2684 1244 2688
rect 1238 2683 1244 2684
rect 1382 2688 1388 2689
rect 1382 2684 1383 2688
rect 1387 2684 1388 2688
rect 1382 2683 1388 2684
rect 1534 2688 1540 2689
rect 1534 2684 1535 2688
rect 1539 2684 1540 2688
rect 1534 2683 1540 2684
rect 1678 2688 1684 2689
rect 1678 2684 1679 2688
rect 1683 2684 1684 2688
rect 1678 2683 1684 2684
rect 1814 2688 1820 2689
rect 1814 2684 1815 2688
rect 1819 2684 1820 2688
rect 1934 2685 1935 2689
rect 1939 2685 1940 2689
rect 1934 2684 1940 2685
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3858 2685 3859 2689
rect 3863 2685 3864 2689
rect 3858 2684 3864 2685
rect 3994 2689 4000 2690
rect 3994 2685 3995 2689
rect 3999 2685 4000 2689
rect 3994 2684 4000 2685
rect 4130 2689 4136 2690
rect 4130 2685 4131 2689
rect 4135 2685 4136 2689
rect 4130 2684 4136 2685
rect 4266 2689 4272 2690
rect 4266 2685 4267 2689
rect 4271 2685 4272 2689
rect 4266 2684 4272 2685
rect 4402 2689 4408 2690
rect 4402 2685 4403 2689
rect 4407 2685 4408 2689
rect 4402 2684 4408 2685
rect 4538 2689 4544 2690
rect 4538 2685 4539 2689
rect 4543 2685 4544 2689
rect 4538 2684 4544 2685
rect 4682 2689 4688 2690
rect 4682 2685 4683 2689
rect 4687 2685 4688 2689
rect 4682 2684 4688 2685
rect 4850 2689 4856 2690
rect 4850 2685 4851 2689
rect 4855 2685 4856 2689
rect 4850 2684 4856 2685
rect 5034 2689 5040 2690
rect 5034 2685 5035 2689
rect 5039 2685 5040 2689
rect 5034 2684 5040 2685
rect 5226 2689 5232 2690
rect 5226 2685 5227 2689
rect 5231 2685 5232 2689
rect 5226 2684 5232 2685
rect 5418 2689 5424 2690
rect 5418 2685 5419 2689
rect 5423 2685 5424 2689
rect 5418 2684 5424 2685
rect 5662 2688 5668 2689
rect 5662 2684 5663 2688
rect 5667 2684 5668 2688
rect 1814 2683 1820 2684
rect 3838 2683 3844 2684
rect 5662 2683 5668 2684
rect 418 2673 424 2674
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 418 2669 419 2673
rect 423 2669 424 2673
rect 418 2668 424 2669
rect 586 2673 592 2674
rect 586 2669 587 2673
rect 591 2669 592 2673
rect 586 2668 592 2669
rect 746 2673 752 2674
rect 746 2669 747 2673
rect 751 2669 752 2673
rect 746 2668 752 2669
rect 906 2673 912 2674
rect 906 2669 907 2673
rect 911 2669 912 2673
rect 906 2668 912 2669
rect 1058 2673 1064 2674
rect 1058 2669 1059 2673
rect 1063 2669 1064 2673
rect 1058 2668 1064 2669
rect 1210 2673 1216 2674
rect 1210 2669 1211 2673
rect 1215 2669 1216 2673
rect 1210 2668 1216 2669
rect 1354 2673 1360 2674
rect 1354 2669 1355 2673
rect 1359 2669 1360 2673
rect 1354 2668 1360 2669
rect 1506 2673 1512 2674
rect 1506 2669 1507 2673
rect 1511 2669 1512 2673
rect 1506 2668 1512 2669
rect 1650 2673 1656 2674
rect 1650 2669 1651 2673
rect 1655 2669 1656 2673
rect 1650 2668 1656 2669
rect 1786 2673 1792 2674
rect 1786 2669 1787 2673
rect 1791 2669 1792 2673
rect 1786 2668 1792 2669
rect 1934 2672 1940 2673
rect 1934 2668 1935 2672
rect 1939 2668 1940 2672
rect 110 2667 116 2668
rect 1934 2667 1940 2668
rect 1974 2609 1980 2610
rect 3798 2609 3804 2610
rect 1974 2605 1975 2609
rect 1979 2605 1980 2609
rect 1974 2604 1980 2605
rect 3270 2608 3276 2609
rect 3270 2604 3271 2608
rect 3275 2604 3276 2608
rect 3270 2603 3276 2604
rect 3406 2608 3412 2609
rect 3406 2604 3407 2608
rect 3411 2604 3412 2608
rect 3406 2603 3412 2604
rect 3542 2608 3548 2609
rect 3542 2604 3543 2608
rect 3547 2604 3548 2608
rect 3542 2603 3548 2604
rect 3678 2608 3684 2609
rect 3678 2604 3679 2608
rect 3683 2604 3684 2608
rect 3798 2605 3799 2609
rect 3803 2605 3804 2609
rect 3798 2604 3804 2605
rect 3678 2603 3684 2604
rect 3242 2593 3248 2594
rect 1974 2592 1980 2593
rect 1974 2588 1975 2592
rect 1979 2588 1980 2592
rect 3242 2589 3243 2593
rect 3247 2589 3248 2593
rect 3242 2588 3248 2589
rect 3378 2593 3384 2594
rect 3378 2589 3379 2593
rect 3383 2589 3384 2593
rect 3378 2588 3384 2589
rect 3514 2593 3520 2594
rect 3514 2589 3515 2593
rect 3519 2589 3520 2593
rect 3514 2588 3520 2589
rect 3650 2593 3656 2594
rect 3650 2589 3651 2593
rect 3655 2589 3656 2593
rect 3650 2588 3656 2589
rect 3798 2592 3804 2593
rect 3798 2588 3799 2592
rect 3803 2588 3804 2592
rect 1974 2587 1980 2588
rect 3798 2587 3804 2588
rect 3838 2540 3844 2541
rect 5662 2540 5668 2541
rect 110 2536 116 2537
rect 1934 2536 1940 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 110 2531 116 2532
rect 234 2535 240 2536
rect 234 2531 235 2535
rect 239 2531 240 2535
rect 234 2530 240 2531
rect 434 2535 440 2536
rect 434 2531 435 2535
rect 439 2531 440 2535
rect 434 2530 440 2531
rect 626 2535 632 2536
rect 626 2531 627 2535
rect 631 2531 632 2535
rect 626 2530 632 2531
rect 810 2535 816 2536
rect 810 2531 811 2535
rect 815 2531 816 2535
rect 810 2530 816 2531
rect 986 2535 992 2536
rect 986 2531 987 2535
rect 991 2531 992 2535
rect 986 2530 992 2531
rect 1154 2535 1160 2536
rect 1154 2531 1155 2535
rect 1159 2531 1160 2535
rect 1154 2530 1160 2531
rect 1322 2535 1328 2536
rect 1322 2531 1323 2535
rect 1327 2531 1328 2535
rect 1322 2530 1328 2531
rect 1482 2535 1488 2536
rect 1482 2531 1483 2535
rect 1487 2531 1488 2535
rect 1482 2530 1488 2531
rect 1642 2535 1648 2536
rect 1642 2531 1643 2535
rect 1647 2531 1648 2535
rect 1642 2530 1648 2531
rect 1786 2535 1792 2536
rect 1786 2531 1787 2535
rect 1791 2531 1792 2535
rect 1934 2532 1935 2536
rect 1939 2532 1940 2536
rect 3838 2536 3839 2540
rect 3843 2536 3844 2540
rect 3838 2535 3844 2536
rect 4178 2539 4184 2540
rect 4178 2535 4179 2539
rect 4183 2535 4184 2539
rect 4178 2534 4184 2535
rect 4394 2539 4400 2540
rect 4394 2535 4395 2539
rect 4399 2535 4400 2539
rect 4394 2534 4400 2535
rect 4642 2539 4648 2540
rect 4642 2535 4643 2539
rect 4647 2535 4648 2539
rect 4642 2534 4648 2535
rect 4906 2539 4912 2540
rect 4906 2535 4907 2539
rect 4911 2535 4912 2539
rect 4906 2534 4912 2535
rect 5186 2539 5192 2540
rect 5186 2535 5187 2539
rect 5191 2535 5192 2539
rect 5186 2534 5192 2535
rect 5466 2539 5472 2540
rect 5466 2535 5467 2539
rect 5471 2535 5472 2539
rect 5662 2536 5663 2540
rect 5667 2536 5668 2540
rect 5662 2535 5668 2536
rect 5466 2534 5472 2535
rect 1934 2531 1940 2532
rect 1786 2530 1792 2531
rect 4206 2524 4212 2525
rect 3838 2523 3844 2524
rect 262 2520 268 2521
rect 110 2519 116 2520
rect 110 2515 111 2519
rect 115 2515 116 2519
rect 262 2516 263 2520
rect 267 2516 268 2520
rect 262 2515 268 2516
rect 462 2520 468 2521
rect 462 2516 463 2520
rect 467 2516 468 2520
rect 462 2515 468 2516
rect 654 2520 660 2521
rect 654 2516 655 2520
rect 659 2516 660 2520
rect 654 2515 660 2516
rect 838 2520 844 2521
rect 838 2516 839 2520
rect 843 2516 844 2520
rect 838 2515 844 2516
rect 1014 2520 1020 2521
rect 1014 2516 1015 2520
rect 1019 2516 1020 2520
rect 1014 2515 1020 2516
rect 1182 2520 1188 2521
rect 1182 2516 1183 2520
rect 1187 2516 1188 2520
rect 1182 2515 1188 2516
rect 1350 2520 1356 2521
rect 1350 2516 1351 2520
rect 1355 2516 1356 2520
rect 1350 2515 1356 2516
rect 1510 2520 1516 2521
rect 1510 2516 1511 2520
rect 1515 2516 1516 2520
rect 1510 2515 1516 2516
rect 1670 2520 1676 2521
rect 1670 2516 1671 2520
rect 1675 2516 1676 2520
rect 1670 2515 1676 2516
rect 1814 2520 1820 2521
rect 1814 2516 1815 2520
rect 1819 2516 1820 2520
rect 1814 2515 1820 2516
rect 1934 2519 1940 2520
rect 1934 2515 1935 2519
rect 1939 2515 1940 2519
rect 3838 2519 3839 2523
rect 3843 2519 3844 2523
rect 4206 2520 4207 2524
rect 4211 2520 4212 2524
rect 4206 2519 4212 2520
rect 4422 2524 4428 2525
rect 4422 2520 4423 2524
rect 4427 2520 4428 2524
rect 4422 2519 4428 2520
rect 4670 2524 4676 2525
rect 4670 2520 4671 2524
rect 4675 2520 4676 2524
rect 4670 2519 4676 2520
rect 4934 2524 4940 2525
rect 4934 2520 4935 2524
rect 4939 2520 4940 2524
rect 4934 2519 4940 2520
rect 5214 2524 5220 2525
rect 5214 2520 5215 2524
rect 5219 2520 5220 2524
rect 5214 2519 5220 2520
rect 5494 2524 5500 2525
rect 5494 2520 5495 2524
rect 5499 2520 5500 2524
rect 5494 2519 5500 2520
rect 5662 2523 5668 2524
rect 5662 2519 5663 2523
rect 5667 2519 5668 2523
rect 3838 2518 3844 2519
rect 5662 2518 5668 2519
rect 110 2514 116 2515
rect 1934 2514 1940 2515
rect 3838 2465 3844 2466
rect 5662 2465 5668 2466
rect 3838 2461 3839 2465
rect 3843 2461 3844 2465
rect 1974 2460 1980 2461
rect 3798 2460 3804 2461
rect 3838 2460 3844 2461
rect 4534 2464 4540 2465
rect 4534 2460 4535 2464
rect 4539 2460 4540 2464
rect 1974 2456 1975 2460
rect 1979 2456 1980 2460
rect 1974 2455 1980 2456
rect 1994 2459 2000 2460
rect 1994 2455 1995 2459
rect 1999 2455 2000 2459
rect 1994 2454 2000 2455
rect 2250 2459 2256 2460
rect 2250 2455 2251 2459
rect 2255 2455 2256 2459
rect 2250 2454 2256 2455
rect 2522 2459 2528 2460
rect 2522 2455 2523 2459
rect 2527 2455 2528 2459
rect 2522 2454 2528 2455
rect 2770 2459 2776 2460
rect 2770 2455 2771 2459
rect 2775 2455 2776 2459
rect 2770 2454 2776 2455
rect 3002 2459 3008 2460
rect 3002 2455 3003 2459
rect 3007 2455 3008 2459
rect 3002 2454 3008 2455
rect 3226 2459 3232 2460
rect 3226 2455 3227 2459
rect 3231 2455 3232 2459
rect 3226 2454 3232 2455
rect 3450 2459 3456 2460
rect 3450 2455 3451 2459
rect 3455 2455 3456 2459
rect 3450 2454 3456 2455
rect 3650 2459 3656 2460
rect 3650 2455 3651 2459
rect 3655 2455 3656 2459
rect 3798 2456 3799 2460
rect 3803 2456 3804 2460
rect 4534 2459 4540 2460
rect 4758 2464 4764 2465
rect 4758 2460 4759 2464
rect 4763 2460 4764 2464
rect 4758 2459 4764 2460
rect 4982 2464 4988 2465
rect 4982 2460 4983 2464
rect 4987 2460 4988 2464
rect 4982 2459 4988 2460
rect 5214 2464 5220 2465
rect 5214 2460 5215 2464
rect 5219 2460 5220 2464
rect 5214 2459 5220 2460
rect 5446 2464 5452 2465
rect 5446 2460 5447 2464
rect 5451 2460 5452 2464
rect 5662 2461 5663 2465
rect 5667 2461 5668 2465
rect 5662 2460 5668 2461
rect 5446 2459 5452 2460
rect 3798 2455 3804 2456
rect 3650 2454 3656 2455
rect 110 2453 116 2454
rect 1934 2453 1940 2454
rect 110 2449 111 2453
rect 115 2449 116 2453
rect 110 2448 116 2449
rect 222 2452 228 2453
rect 222 2448 223 2452
rect 227 2448 228 2452
rect 222 2447 228 2448
rect 422 2452 428 2453
rect 422 2448 423 2452
rect 427 2448 428 2452
rect 422 2447 428 2448
rect 622 2452 628 2453
rect 622 2448 623 2452
rect 627 2448 628 2452
rect 622 2447 628 2448
rect 814 2452 820 2453
rect 814 2448 815 2452
rect 819 2448 820 2452
rect 814 2447 820 2448
rect 1014 2452 1020 2453
rect 1014 2448 1015 2452
rect 1019 2448 1020 2452
rect 1014 2447 1020 2448
rect 1214 2452 1220 2453
rect 1214 2448 1215 2452
rect 1219 2448 1220 2452
rect 1934 2449 1935 2453
rect 1939 2449 1940 2453
rect 4506 2449 4512 2450
rect 1934 2448 1940 2449
rect 3838 2448 3844 2449
rect 1214 2447 1220 2448
rect 2022 2444 2028 2445
rect 1974 2443 1980 2444
rect 1974 2439 1975 2443
rect 1979 2439 1980 2443
rect 2022 2440 2023 2444
rect 2027 2440 2028 2444
rect 2022 2439 2028 2440
rect 2278 2444 2284 2445
rect 2278 2440 2279 2444
rect 2283 2440 2284 2444
rect 2278 2439 2284 2440
rect 2550 2444 2556 2445
rect 2550 2440 2551 2444
rect 2555 2440 2556 2444
rect 2550 2439 2556 2440
rect 2798 2444 2804 2445
rect 2798 2440 2799 2444
rect 2803 2440 2804 2444
rect 2798 2439 2804 2440
rect 3030 2444 3036 2445
rect 3030 2440 3031 2444
rect 3035 2440 3036 2444
rect 3030 2439 3036 2440
rect 3254 2444 3260 2445
rect 3254 2440 3255 2444
rect 3259 2440 3260 2444
rect 3254 2439 3260 2440
rect 3478 2444 3484 2445
rect 3478 2440 3479 2444
rect 3483 2440 3484 2444
rect 3478 2439 3484 2440
rect 3678 2444 3684 2445
rect 3838 2444 3839 2448
rect 3843 2444 3844 2448
rect 4506 2445 4507 2449
rect 4511 2445 4512 2449
rect 4506 2444 4512 2445
rect 4730 2449 4736 2450
rect 4730 2445 4731 2449
rect 4735 2445 4736 2449
rect 4730 2444 4736 2445
rect 4954 2449 4960 2450
rect 4954 2445 4955 2449
rect 4959 2445 4960 2449
rect 4954 2444 4960 2445
rect 5186 2449 5192 2450
rect 5186 2445 5187 2449
rect 5191 2445 5192 2449
rect 5186 2444 5192 2445
rect 5418 2449 5424 2450
rect 5418 2445 5419 2449
rect 5423 2445 5424 2449
rect 5418 2444 5424 2445
rect 5662 2448 5668 2449
rect 5662 2444 5663 2448
rect 5667 2444 5668 2448
rect 3678 2440 3679 2444
rect 3683 2440 3684 2444
rect 3678 2439 3684 2440
rect 3798 2443 3804 2444
rect 3838 2443 3844 2444
rect 5662 2443 5668 2444
rect 3798 2439 3799 2443
rect 3803 2439 3804 2443
rect 1974 2438 1980 2439
rect 3798 2438 3804 2439
rect 194 2437 200 2438
rect 110 2436 116 2437
rect 110 2432 111 2436
rect 115 2432 116 2436
rect 194 2433 195 2437
rect 199 2433 200 2437
rect 194 2432 200 2433
rect 394 2437 400 2438
rect 394 2433 395 2437
rect 399 2433 400 2437
rect 394 2432 400 2433
rect 594 2437 600 2438
rect 594 2433 595 2437
rect 599 2433 600 2437
rect 594 2432 600 2433
rect 786 2437 792 2438
rect 786 2433 787 2437
rect 791 2433 792 2437
rect 786 2432 792 2433
rect 986 2437 992 2438
rect 986 2433 987 2437
rect 991 2433 992 2437
rect 986 2432 992 2433
rect 1186 2437 1192 2438
rect 1186 2433 1187 2437
rect 1191 2433 1192 2437
rect 1186 2432 1192 2433
rect 1934 2436 1940 2437
rect 1934 2432 1935 2436
rect 1939 2432 1940 2436
rect 110 2431 116 2432
rect 1934 2431 1940 2432
rect 1974 2385 1980 2386
rect 3798 2385 3804 2386
rect 1974 2381 1975 2385
rect 1979 2381 1980 2385
rect 1974 2380 1980 2381
rect 2054 2384 2060 2385
rect 2054 2380 2055 2384
rect 2059 2380 2060 2384
rect 2054 2379 2060 2380
rect 2214 2384 2220 2385
rect 2214 2380 2215 2384
rect 2219 2380 2220 2384
rect 2214 2379 2220 2380
rect 2374 2384 2380 2385
rect 2374 2380 2375 2384
rect 2379 2380 2380 2384
rect 2374 2379 2380 2380
rect 2542 2384 2548 2385
rect 2542 2380 2543 2384
rect 2547 2380 2548 2384
rect 2542 2379 2548 2380
rect 2710 2384 2716 2385
rect 2710 2380 2711 2384
rect 2715 2380 2716 2384
rect 2710 2379 2716 2380
rect 2870 2384 2876 2385
rect 2870 2380 2871 2384
rect 2875 2380 2876 2384
rect 2870 2379 2876 2380
rect 3030 2384 3036 2385
rect 3030 2380 3031 2384
rect 3035 2380 3036 2384
rect 3030 2379 3036 2380
rect 3190 2384 3196 2385
rect 3190 2380 3191 2384
rect 3195 2380 3196 2384
rect 3190 2379 3196 2380
rect 3358 2384 3364 2385
rect 3358 2380 3359 2384
rect 3363 2380 3364 2384
rect 3358 2379 3364 2380
rect 3526 2384 3532 2385
rect 3526 2380 3527 2384
rect 3531 2380 3532 2384
rect 3798 2381 3799 2385
rect 3803 2381 3804 2385
rect 3798 2380 3804 2381
rect 3526 2379 3532 2380
rect 2026 2369 2032 2370
rect 1974 2368 1980 2369
rect 1974 2364 1975 2368
rect 1979 2364 1980 2368
rect 2026 2365 2027 2369
rect 2031 2365 2032 2369
rect 2026 2364 2032 2365
rect 2186 2369 2192 2370
rect 2186 2365 2187 2369
rect 2191 2365 2192 2369
rect 2186 2364 2192 2365
rect 2346 2369 2352 2370
rect 2346 2365 2347 2369
rect 2351 2365 2352 2369
rect 2346 2364 2352 2365
rect 2514 2369 2520 2370
rect 2514 2365 2515 2369
rect 2519 2365 2520 2369
rect 2514 2364 2520 2365
rect 2682 2369 2688 2370
rect 2682 2365 2683 2369
rect 2687 2365 2688 2369
rect 2682 2364 2688 2365
rect 2842 2369 2848 2370
rect 2842 2365 2843 2369
rect 2847 2365 2848 2369
rect 2842 2364 2848 2365
rect 3002 2369 3008 2370
rect 3002 2365 3003 2369
rect 3007 2365 3008 2369
rect 3002 2364 3008 2365
rect 3162 2369 3168 2370
rect 3162 2365 3163 2369
rect 3167 2365 3168 2369
rect 3162 2364 3168 2365
rect 3330 2369 3336 2370
rect 3330 2365 3331 2369
rect 3335 2365 3336 2369
rect 3330 2364 3336 2365
rect 3498 2369 3504 2370
rect 3498 2365 3499 2369
rect 3503 2365 3504 2369
rect 3498 2364 3504 2365
rect 3798 2368 3804 2369
rect 3798 2364 3799 2368
rect 3803 2364 3804 2368
rect 1974 2363 1980 2364
rect 3798 2363 3804 2364
rect 3838 2316 3844 2317
rect 5662 2316 5668 2317
rect 3838 2312 3839 2316
rect 3843 2312 3844 2316
rect 3838 2311 3844 2312
rect 4706 2315 4712 2316
rect 4706 2311 4707 2315
rect 4711 2311 4712 2315
rect 4706 2310 4712 2311
rect 4866 2315 4872 2316
rect 4866 2311 4867 2315
rect 4871 2311 4872 2315
rect 4866 2310 4872 2311
rect 5026 2315 5032 2316
rect 5026 2311 5027 2315
rect 5031 2311 5032 2315
rect 5026 2310 5032 2311
rect 5186 2315 5192 2316
rect 5186 2311 5187 2315
rect 5191 2311 5192 2315
rect 5186 2310 5192 2311
rect 5346 2315 5352 2316
rect 5346 2311 5347 2315
rect 5351 2311 5352 2315
rect 5346 2310 5352 2311
rect 5514 2315 5520 2316
rect 5514 2311 5515 2315
rect 5519 2311 5520 2315
rect 5662 2312 5663 2316
rect 5667 2312 5668 2316
rect 5662 2311 5668 2312
rect 5514 2310 5520 2311
rect 4734 2300 4740 2301
rect 3838 2299 3844 2300
rect 3838 2295 3839 2299
rect 3843 2295 3844 2299
rect 4734 2296 4735 2300
rect 4739 2296 4740 2300
rect 4734 2295 4740 2296
rect 4894 2300 4900 2301
rect 4894 2296 4895 2300
rect 4899 2296 4900 2300
rect 4894 2295 4900 2296
rect 5054 2300 5060 2301
rect 5054 2296 5055 2300
rect 5059 2296 5060 2300
rect 5054 2295 5060 2296
rect 5214 2300 5220 2301
rect 5214 2296 5215 2300
rect 5219 2296 5220 2300
rect 5214 2295 5220 2296
rect 5374 2300 5380 2301
rect 5374 2296 5375 2300
rect 5379 2296 5380 2300
rect 5374 2295 5380 2296
rect 5542 2300 5548 2301
rect 5542 2296 5543 2300
rect 5547 2296 5548 2300
rect 5542 2295 5548 2296
rect 5662 2299 5668 2300
rect 5662 2295 5663 2299
rect 5667 2295 5668 2299
rect 3838 2294 3844 2295
rect 5662 2294 5668 2295
rect 110 2292 116 2293
rect 1934 2292 1940 2293
rect 110 2288 111 2292
rect 115 2288 116 2292
rect 110 2287 116 2288
rect 130 2291 136 2292
rect 130 2287 131 2291
rect 135 2287 136 2291
rect 130 2286 136 2287
rect 290 2291 296 2292
rect 290 2287 291 2291
rect 295 2287 296 2291
rect 290 2286 296 2287
rect 482 2291 488 2292
rect 482 2287 483 2291
rect 487 2287 488 2291
rect 482 2286 488 2287
rect 674 2291 680 2292
rect 674 2287 675 2291
rect 679 2287 680 2291
rect 674 2286 680 2287
rect 866 2291 872 2292
rect 866 2287 867 2291
rect 871 2287 872 2291
rect 1934 2288 1935 2292
rect 1939 2288 1940 2292
rect 1934 2287 1940 2288
rect 866 2286 872 2287
rect 158 2276 164 2277
rect 110 2275 116 2276
rect 110 2271 111 2275
rect 115 2271 116 2275
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 510 2276 516 2277
rect 510 2272 511 2276
rect 515 2272 516 2276
rect 510 2271 516 2272
rect 702 2276 708 2277
rect 702 2272 703 2276
rect 707 2272 708 2276
rect 702 2271 708 2272
rect 894 2276 900 2277
rect 894 2272 895 2276
rect 899 2272 900 2276
rect 894 2271 900 2272
rect 1934 2275 1940 2276
rect 1934 2271 1935 2275
rect 1939 2271 1940 2275
rect 110 2270 116 2271
rect 1934 2270 1940 2271
rect 3838 2229 3844 2230
rect 5662 2229 5668 2230
rect 1974 2228 1980 2229
rect 3798 2228 3804 2229
rect 1974 2224 1975 2228
rect 1979 2224 1980 2228
rect 1974 2223 1980 2224
rect 2138 2227 2144 2228
rect 2138 2223 2139 2227
rect 2143 2223 2144 2227
rect 2138 2222 2144 2223
rect 2274 2227 2280 2228
rect 2274 2223 2275 2227
rect 2279 2223 2280 2227
rect 2274 2222 2280 2223
rect 2410 2227 2416 2228
rect 2410 2223 2411 2227
rect 2415 2223 2416 2227
rect 2410 2222 2416 2223
rect 2546 2227 2552 2228
rect 2546 2223 2547 2227
rect 2551 2223 2552 2227
rect 2546 2222 2552 2223
rect 2682 2227 2688 2228
rect 2682 2223 2683 2227
rect 2687 2223 2688 2227
rect 2682 2222 2688 2223
rect 2818 2227 2824 2228
rect 2818 2223 2819 2227
rect 2823 2223 2824 2227
rect 2818 2222 2824 2223
rect 2954 2227 2960 2228
rect 2954 2223 2955 2227
rect 2959 2223 2960 2227
rect 2954 2222 2960 2223
rect 3090 2227 3096 2228
rect 3090 2223 3091 2227
rect 3095 2223 3096 2227
rect 3090 2222 3096 2223
rect 3226 2227 3232 2228
rect 3226 2223 3227 2227
rect 3231 2223 3232 2227
rect 3226 2222 3232 2223
rect 3362 2227 3368 2228
rect 3362 2223 3363 2227
rect 3367 2223 3368 2227
rect 3798 2224 3799 2228
rect 3803 2224 3804 2228
rect 3838 2225 3839 2229
rect 3843 2225 3844 2229
rect 3838 2224 3844 2225
rect 4734 2228 4740 2229
rect 4734 2224 4735 2228
rect 4739 2224 4740 2228
rect 3798 2223 3804 2224
rect 4734 2223 4740 2224
rect 4886 2228 4892 2229
rect 4886 2224 4887 2228
rect 4891 2224 4892 2228
rect 4886 2223 4892 2224
rect 5046 2228 5052 2229
rect 5046 2224 5047 2228
rect 5051 2224 5052 2228
rect 5046 2223 5052 2224
rect 5214 2228 5220 2229
rect 5214 2224 5215 2228
rect 5219 2224 5220 2228
rect 5214 2223 5220 2224
rect 5390 2228 5396 2229
rect 5390 2224 5391 2228
rect 5395 2224 5396 2228
rect 5390 2223 5396 2224
rect 5542 2228 5548 2229
rect 5542 2224 5543 2228
rect 5547 2224 5548 2228
rect 5662 2225 5663 2229
rect 5667 2225 5668 2229
rect 5662 2224 5668 2225
rect 5542 2223 5548 2224
rect 3362 2222 3368 2223
rect 110 2217 116 2218
rect 1934 2217 1940 2218
rect 110 2213 111 2217
rect 115 2213 116 2217
rect 110 2212 116 2213
rect 158 2216 164 2217
rect 158 2212 159 2216
rect 163 2212 164 2216
rect 158 2211 164 2212
rect 294 2216 300 2217
rect 294 2212 295 2216
rect 299 2212 300 2216
rect 294 2211 300 2212
rect 438 2216 444 2217
rect 438 2212 439 2216
rect 443 2212 444 2216
rect 438 2211 444 2212
rect 590 2216 596 2217
rect 590 2212 591 2216
rect 595 2212 596 2216
rect 590 2211 596 2212
rect 742 2216 748 2217
rect 742 2212 743 2216
rect 747 2212 748 2216
rect 1934 2213 1935 2217
rect 1939 2213 1940 2217
rect 4706 2213 4712 2214
rect 1934 2212 1940 2213
rect 2166 2212 2172 2213
rect 742 2211 748 2212
rect 1974 2211 1980 2212
rect 1974 2207 1975 2211
rect 1979 2207 1980 2211
rect 2166 2208 2167 2212
rect 2171 2208 2172 2212
rect 2166 2207 2172 2208
rect 2302 2212 2308 2213
rect 2302 2208 2303 2212
rect 2307 2208 2308 2212
rect 2302 2207 2308 2208
rect 2438 2212 2444 2213
rect 2438 2208 2439 2212
rect 2443 2208 2444 2212
rect 2438 2207 2444 2208
rect 2574 2212 2580 2213
rect 2574 2208 2575 2212
rect 2579 2208 2580 2212
rect 2574 2207 2580 2208
rect 2710 2212 2716 2213
rect 2710 2208 2711 2212
rect 2715 2208 2716 2212
rect 2710 2207 2716 2208
rect 2846 2212 2852 2213
rect 2846 2208 2847 2212
rect 2851 2208 2852 2212
rect 2846 2207 2852 2208
rect 2982 2212 2988 2213
rect 2982 2208 2983 2212
rect 2987 2208 2988 2212
rect 2982 2207 2988 2208
rect 3118 2212 3124 2213
rect 3118 2208 3119 2212
rect 3123 2208 3124 2212
rect 3118 2207 3124 2208
rect 3254 2212 3260 2213
rect 3254 2208 3255 2212
rect 3259 2208 3260 2212
rect 3254 2207 3260 2208
rect 3390 2212 3396 2213
rect 3838 2212 3844 2213
rect 3390 2208 3391 2212
rect 3395 2208 3396 2212
rect 3390 2207 3396 2208
rect 3798 2211 3804 2212
rect 3798 2207 3799 2211
rect 3803 2207 3804 2211
rect 3838 2208 3839 2212
rect 3843 2208 3844 2212
rect 4706 2209 4707 2213
rect 4711 2209 4712 2213
rect 4706 2208 4712 2209
rect 4858 2213 4864 2214
rect 4858 2209 4859 2213
rect 4863 2209 4864 2213
rect 4858 2208 4864 2209
rect 5018 2213 5024 2214
rect 5018 2209 5019 2213
rect 5023 2209 5024 2213
rect 5018 2208 5024 2209
rect 5186 2213 5192 2214
rect 5186 2209 5187 2213
rect 5191 2209 5192 2213
rect 5186 2208 5192 2209
rect 5362 2213 5368 2214
rect 5362 2209 5363 2213
rect 5367 2209 5368 2213
rect 5362 2208 5368 2209
rect 5514 2213 5520 2214
rect 5514 2209 5515 2213
rect 5519 2209 5520 2213
rect 5514 2208 5520 2209
rect 5662 2212 5668 2213
rect 5662 2208 5663 2212
rect 5667 2208 5668 2212
rect 3838 2207 3844 2208
rect 5662 2207 5668 2208
rect 1974 2206 1980 2207
rect 3798 2206 3804 2207
rect 130 2201 136 2202
rect 110 2200 116 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 130 2197 131 2201
rect 135 2197 136 2201
rect 130 2196 136 2197
rect 266 2201 272 2202
rect 266 2197 267 2201
rect 271 2197 272 2201
rect 266 2196 272 2197
rect 410 2201 416 2202
rect 410 2197 411 2201
rect 415 2197 416 2201
rect 410 2196 416 2197
rect 562 2201 568 2202
rect 562 2197 563 2201
rect 567 2197 568 2201
rect 562 2196 568 2197
rect 714 2201 720 2202
rect 714 2197 715 2201
rect 719 2197 720 2201
rect 714 2196 720 2197
rect 1934 2200 1940 2201
rect 1934 2196 1935 2200
rect 1939 2196 1940 2200
rect 110 2195 116 2196
rect 1934 2195 1940 2196
rect 1974 2149 1980 2150
rect 3798 2149 3804 2150
rect 1974 2145 1975 2149
rect 1979 2145 1980 2149
rect 1974 2144 1980 2145
rect 2022 2148 2028 2149
rect 2022 2144 2023 2148
rect 2027 2144 2028 2148
rect 2022 2143 2028 2144
rect 2158 2148 2164 2149
rect 2158 2144 2159 2148
rect 2163 2144 2164 2148
rect 2158 2143 2164 2144
rect 2294 2148 2300 2149
rect 2294 2144 2295 2148
rect 2299 2144 2300 2148
rect 2294 2143 2300 2144
rect 2430 2148 2436 2149
rect 2430 2144 2431 2148
rect 2435 2144 2436 2148
rect 2430 2143 2436 2144
rect 2566 2148 2572 2149
rect 2566 2144 2567 2148
rect 2571 2144 2572 2148
rect 2566 2143 2572 2144
rect 2702 2148 2708 2149
rect 2702 2144 2703 2148
rect 2707 2144 2708 2148
rect 2702 2143 2708 2144
rect 2838 2148 2844 2149
rect 2838 2144 2839 2148
rect 2843 2144 2844 2148
rect 2838 2143 2844 2144
rect 2974 2148 2980 2149
rect 2974 2144 2975 2148
rect 2979 2144 2980 2148
rect 2974 2143 2980 2144
rect 3110 2148 3116 2149
rect 3110 2144 3111 2148
rect 3115 2144 3116 2148
rect 3110 2143 3116 2144
rect 3246 2148 3252 2149
rect 3246 2144 3247 2148
rect 3251 2144 3252 2148
rect 3798 2145 3799 2149
rect 3803 2145 3804 2149
rect 3798 2144 3804 2145
rect 3246 2143 3252 2144
rect 1994 2133 2000 2134
rect 1974 2132 1980 2133
rect 1974 2128 1975 2132
rect 1979 2128 1980 2132
rect 1994 2129 1995 2133
rect 1999 2129 2000 2133
rect 1994 2128 2000 2129
rect 2130 2133 2136 2134
rect 2130 2129 2131 2133
rect 2135 2129 2136 2133
rect 2130 2128 2136 2129
rect 2266 2133 2272 2134
rect 2266 2129 2267 2133
rect 2271 2129 2272 2133
rect 2266 2128 2272 2129
rect 2402 2133 2408 2134
rect 2402 2129 2403 2133
rect 2407 2129 2408 2133
rect 2402 2128 2408 2129
rect 2538 2133 2544 2134
rect 2538 2129 2539 2133
rect 2543 2129 2544 2133
rect 2538 2128 2544 2129
rect 2674 2133 2680 2134
rect 2674 2129 2675 2133
rect 2679 2129 2680 2133
rect 2674 2128 2680 2129
rect 2810 2133 2816 2134
rect 2810 2129 2811 2133
rect 2815 2129 2816 2133
rect 2810 2128 2816 2129
rect 2946 2133 2952 2134
rect 2946 2129 2947 2133
rect 2951 2129 2952 2133
rect 2946 2128 2952 2129
rect 3082 2133 3088 2134
rect 3082 2129 3083 2133
rect 3087 2129 3088 2133
rect 3082 2128 3088 2129
rect 3218 2133 3224 2134
rect 3218 2129 3219 2133
rect 3223 2129 3224 2133
rect 3218 2128 3224 2129
rect 3798 2132 3804 2133
rect 3798 2128 3799 2132
rect 3803 2128 3804 2132
rect 1974 2127 1980 2128
rect 3798 2127 3804 2128
rect 3838 2072 3844 2073
rect 5662 2072 5668 2073
rect 110 2068 116 2069
rect 1934 2068 1940 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 130 2067 136 2068
rect 130 2063 131 2067
rect 135 2063 136 2067
rect 130 2062 136 2063
rect 330 2067 336 2068
rect 330 2063 331 2067
rect 335 2063 336 2067
rect 330 2062 336 2063
rect 554 2067 560 2068
rect 554 2063 555 2067
rect 559 2063 560 2067
rect 554 2062 560 2063
rect 778 2067 784 2068
rect 778 2063 779 2067
rect 783 2063 784 2067
rect 778 2062 784 2063
rect 1010 2067 1016 2068
rect 1010 2063 1011 2067
rect 1015 2063 1016 2067
rect 1934 2064 1935 2068
rect 1939 2064 1940 2068
rect 3838 2068 3839 2072
rect 3843 2068 3844 2072
rect 3838 2067 3844 2068
rect 4786 2071 4792 2072
rect 4786 2067 4787 2071
rect 4791 2067 4792 2071
rect 4786 2066 4792 2067
rect 4922 2071 4928 2072
rect 4922 2067 4923 2071
rect 4927 2067 4928 2071
rect 4922 2066 4928 2067
rect 5066 2071 5072 2072
rect 5066 2067 5067 2071
rect 5071 2067 5072 2071
rect 5066 2066 5072 2067
rect 5218 2071 5224 2072
rect 5218 2067 5219 2071
rect 5223 2067 5224 2071
rect 5218 2066 5224 2067
rect 5378 2071 5384 2072
rect 5378 2067 5379 2071
rect 5383 2067 5384 2071
rect 5378 2066 5384 2067
rect 5514 2071 5520 2072
rect 5514 2067 5515 2071
rect 5519 2067 5520 2071
rect 5662 2068 5663 2072
rect 5667 2068 5668 2072
rect 5662 2067 5668 2068
rect 5514 2066 5520 2067
rect 1934 2063 1940 2064
rect 1010 2062 1016 2063
rect 4814 2056 4820 2057
rect 3838 2055 3844 2056
rect 158 2052 164 2053
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 158 2048 159 2052
rect 163 2048 164 2052
rect 158 2047 164 2048
rect 358 2052 364 2053
rect 358 2048 359 2052
rect 363 2048 364 2052
rect 358 2047 364 2048
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 806 2052 812 2053
rect 806 2048 807 2052
rect 811 2048 812 2052
rect 806 2047 812 2048
rect 1038 2052 1044 2053
rect 1038 2048 1039 2052
rect 1043 2048 1044 2052
rect 1038 2047 1044 2048
rect 1934 2051 1940 2052
rect 1934 2047 1935 2051
rect 1939 2047 1940 2051
rect 3838 2051 3839 2055
rect 3843 2051 3844 2055
rect 4814 2052 4815 2056
rect 4819 2052 4820 2056
rect 4814 2051 4820 2052
rect 4950 2056 4956 2057
rect 4950 2052 4951 2056
rect 4955 2052 4956 2056
rect 4950 2051 4956 2052
rect 5094 2056 5100 2057
rect 5094 2052 5095 2056
rect 5099 2052 5100 2056
rect 5094 2051 5100 2052
rect 5246 2056 5252 2057
rect 5246 2052 5247 2056
rect 5251 2052 5252 2056
rect 5246 2051 5252 2052
rect 5406 2056 5412 2057
rect 5406 2052 5407 2056
rect 5411 2052 5412 2056
rect 5406 2051 5412 2052
rect 5542 2056 5548 2057
rect 5542 2052 5543 2056
rect 5547 2052 5548 2056
rect 5542 2051 5548 2052
rect 5662 2055 5668 2056
rect 5662 2051 5663 2055
rect 5667 2051 5668 2055
rect 3838 2050 3844 2051
rect 5662 2050 5668 2051
rect 110 2046 116 2047
rect 1934 2046 1940 2047
rect 3838 1993 3844 1994
rect 5662 1993 5668 1994
rect 1974 1992 1980 1993
rect 3798 1992 3804 1993
rect 110 1989 116 1990
rect 1934 1989 1940 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 110 1984 116 1985
rect 158 1988 164 1989
rect 158 1984 159 1988
rect 163 1984 164 1988
rect 158 1983 164 1984
rect 462 1988 468 1989
rect 462 1984 463 1988
rect 467 1984 468 1988
rect 462 1983 468 1984
rect 798 1988 804 1989
rect 798 1984 799 1988
rect 803 1984 804 1988
rect 798 1983 804 1984
rect 1142 1988 1148 1989
rect 1142 1984 1143 1988
rect 1147 1984 1148 1988
rect 1142 1983 1148 1984
rect 1486 1988 1492 1989
rect 1486 1984 1487 1988
rect 1491 1984 1492 1988
rect 1486 1983 1492 1984
rect 1814 1988 1820 1989
rect 1814 1984 1815 1988
rect 1819 1984 1820 1988
rect 1934 1985 1935 1989
rect 1939 1985 1940 1989
rect 1974 1988 1975 1992
rect 1979 1988 1980 1992
rect 1974 1987 1980 1988
rect 1994 1991 2000 1992
rect 1994 1987 1995 1991
rect 1999 1987 2000 1991
rect 1994 1986 2000 1987
rect 2130 1991 2136 1992
rect 2130 1987 2131 1991
rect 2135 1987 2136 1991
rect 2130 1986 2136 1987
rect 2266 1991 2272 1992
rect 2266 1987 2267 1991
rect 2271 1987 2272 1991
rect 2266 1986 2272 1987
rect 2402 1991 2408 1992
rect 2402 1987 2403 1991
rect 2407 1987 2408 1991
rect 2402 1986 2408 1987
rect 2538 1991 2544 1992
rect 2538 1987 2539 1991
rect 2543 1987 2544 1991
rect 2538 1986 2544 1987
rect 2674 1991 2680 1992
rect 2674 1987 2675 1991
rect 2679 1987 2680 1991
rect 2674 1986 2680 1987
rect 2810 1991 2816 1992
rect 2810 1987 2811 1991
rect 2815 1987 2816 1991
rect 2810 1986 2816 1987
rect 2946 1991 2952 1992
rect 2946 1987 2947 1991
rect 2951 1987 2952 1991
rect 2946 1986 2952 1987
rect 3090 1991 3096 1992
rect 3090 1987 3091 1991
rect 3095 1987 3096 1991
rect 3090 1986 3096 1987
rect 3242 1991 3248 1992
rect 3242 1987 3243 1991
rect 3247 1987 3248 1991
rect 3242 1986 3248 1987
rect 3394 1991 3400 1992
rect 3394 1987 3395 1991
rect 3399 1987 3400 1991
rect 3798 1988 3799 1992
rect 3803 1988 3804 1992
rect 3838 1989 3839 1993
rect 3843 1989 3844 1993
rect 3838 1988 3844 1989
rect 4862 1992 4868 1993
rect 4862 1988 4863 1992
rect 4867 1988 4868 1992
rect 3798 1987 3804 1988
rect 4862 1987 4868 1988
rect 4998 1992 5004 1993
rect 4998 1988 4999 1992
rect 5003 1988 5004 1992
rect 4998 1987 5004 1988
rect 5134 1992 5140 1993
rect 5134 1988 5135 1992
rect 5139 1988 5140 1992
rect 5134 1987 5140 1988
rect 5270 1992 5276 1993
rect 5270 1988 5271 1992
rect 5275 1988 5276 1992
rect 5270 1987 5276 1988
rect 5406 1992 5412 1993
rect 5406 1988 5407 1992
rect 5411 1988 5412 1992
rect 5406 1987 5412 1988
rect 5542 1992 5548 1993
rect 5542 1988 5543 1992
rect 5547 1988 5548 1992
rect 5662 1989 5663 1993
rect 5667 1989 5668 1993
rect 5662 1988 5668 1989
rect 5542 1987 5548 1988
rect 3394 1986 3400 1987
rect 1934 1984 1940 1985
rect 1814 1983 1820 1984
rect 4834 1977 4840 1978
rect 2022 1976 2028 1977
rect 1974 1975 1980 1976
rect 130 1973 136 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 130 1969 131 1973
rect 135 1969 136 1973
rect 130 1968 136 1969
rect 434 1973 440 1974
rect 434 1969 435 1973
rect 439 1969 440 1973
rect 434 1968 440 1969
rect 770 1973 776 1974
rect 770 1969 771 1973
rect 775 1969 776 1973
rect 770 1968 776 1969
rect 1114 1973 1120 1974
rect 1114 1969 1115 1973
rect 1119 1969 1120 1973
rect 1114 1968 1120 1969
rect 1458 1973 1464 1974
rect 1458 1969 1459 1973
rect 1463 1969 1464 1973
rect 1458 1968 1464 1969
rect 1786 1973 1792 1974
rect 1786 1969 1787 1973
rect 1791 1969 1792 1973
rect 1786 1968 1792 1969
rect 1934 1972 1940 1973
rect 1934 1968 1935 1972
rect 1939 1968 1940 1972
rect 1974 1971 1975 1975
rect 1979 1971 1980 1975
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2158 1976 2164 1977
rect 2158 1972 2159 1976
rect 2163 1972 2164 1976
rect 2158 1971 2164 1972
rect 2294 1976 2300 1977
rect 2294 1972 2295 1976
rect 2299 1972 2300 1976
rect 2294 1971 2300 1972
rect 2430 1976 2436 1977
rect 2430 1972 2431 1976
rect 2435 1972 2436 1976
rect 2430 1971 2436 1972
rect 2566 1976 2572 1977
rect 2566 1972 2567 1976
rect 2571 1972 2572 1976
rect 2566 1971 2572 1972
rect 2702 1976 2708 1977
rect 2702 1972 2703 1976
rect 2707 1972 2708 1976
rect 2702 1971 2708 1972
rect 2838 1976 2844 1977
rect 2838 1972 2839 1976
rect 2843 1972 2844 1976
rect 2838 1971 2844 1972
rect 2974 1976 2980 1977
rect 2974 1972 2975 1976
rect 2979 1972 2980 1976
rect 2974 1971 2980 1972
rect 3118 1976 3124 1977
rect 3118 1972 3119 1976
rect 3123 1972 3124 1976
rect 3118 1971 3124 1972
rect 3270 1976 3276 1977
rect 3270 1972 3271 1976
rect 3275 1972 3276 1976
rect 3270 1971 3276 1972
rect 3422 1976 3428 1977
rect 3838 1976 3844 1977
rect 3422 1972 3423 1976
rect 3427 1972 3428 1976
rect 3422 1971 3428 1972
rect 3798 1975 3804 1976
rect 3798 1971 3799 1975
rect 3803 1971 3804 1975
rect 3838 1972 3839 1976
rect 3843 1972 3844 1976
rect 4834 1973 4835 1977
rect 4839 1973 4840 1977
rect 4834 1972 4840 1973
rect 4970 1977 4976 1978
rect 4970 1973 4971 1977
rect 4975 1973 4976 1977
rect 4970 1972 4976 1973
rect 5106 1977 5112 1978
rect 5106 1973 5107 1977
rect 5111 1973 5112 1977
rect 5106 1972 5112 1973
rect 5242 1977 5248 1978
rect 5242 1973 5243 1977
rect 5247 1973 5248 1977
rect 5242 1972 5248 1973
rect 5378 1977 5384 1978
rect 5378 1973 5379 1977
rect 5383 1973 5384 1977
rect 5378 1972 5384 1973
rect 5514 1977 5520 1978
rect 5514 1973 5515 1977
rect 5519 1973 5520 1977
rect 5514 1972 5520 1973
rect 5662 1976 5668 1977
rect 5662 1972 5663 1976
rect 5667 1972 5668 1976
rect 3838 1971 3844 1972
rect 5662 1971 5668 1972
rect 1974 1970 1980 1971
rect 3798 1970 3804 1971
rect 110 1967 116 1968
rect 1934 1967 1940 1968
rect 1974 1909 1980 1910
rect 3798 1909 3804 1910
rect 1974 1905 1975 1909
rect 1979 1905 1980 1909
rect 1974 1904 1980 1905
rect 2526 1908 2532 1909
rect 2526 1904 2527 1908
rect 2531 1904 2532 1908
rect 2526 1903 2532 1904
rect 2662 1908 2668 1909
rect 2662 1904 2663 1908
rect 2667 1904 2668 1908
rect 2662 1903 2668 1904
rect 2798 1908 2804 1909
rect 2798 1904 2799 1908
rect 2803 1904 2804 1908
rect 2798 1903 2804 1904
rect 2934 1908 2940 1909
rect 2934 1904 2935 1908
rect 2939 1904 2940 1908
rect 2934 1903 2940 1904
rect 3070 1908 3076 1909
rect 3070 1904 3071 1908
rect 3075 1904 3076 1908
rect 3070 1903 3076 1904
rect 3206 1908 3212 1909
rect 3206 1904 3207 1908
rect 3211 1904 3212 1908
rect 3206 1903 3212 1904
rect 3350 1908 3356 1909
rect 3350 1904 3351 1908
rect 3355 1904 3356 1908
rect 3798 1905 3799 1909
rect 3803 1905 3804 1909
rect 3798 1904 3804 1905
rect 3350 1903 3356 1904
rect 2498 1893 2504 1894
rect 1974 1892 1980 1893
rect 1974 1888 1975 1892
rect 1979 1888 1980 1892
rect 2498 1889 2499 1893
rect 2503 1889 2504 1893
rect 2498 1888 2504 1889
rect 2634 1893 2640 1894
rect 2634 1889 2635 1893
rect 2639 1889 2640 1893
rect 2634 1888 2640 1889
rect 2770 1893 2776 1894
rect 2770 1889 2771 1893
rect 2775 1889 2776 1893
rect 2770 1888 2776 1889
rect 2906 1893 2912 1894
rect 2906 1889 2907 1893
rect 2911 1889 2912 1893
rect 2906 1888 2912 1889
rect 3042 1893 3048 1894
rect 3042 1889 3043 1893
rect 3047 1889 3048 1893
rect 3042 1888 3048 1889
rect 3178 1893 3184 1894
rect 3178 1889 3179 1893
rect 3183 1889 3184 1893
rect 3178 1888 3184 1889
rect 3322 1893 3328 1894
rect 3322 1889 3323 1893
rect 3327 1889 3328 1893
rect 3322 1888 3328 1889
rect 3798 1892 3804 1893
rect 3798 1888 3799 1892
rect 3803 1888 3804 1892
rect 1974 1887 1980 1888
rect 3798 1887 3804 1888
rect 110 1840 116 1841
rect 1934 1840 1940 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 110 1835 116 1836
rect 194 1839 200 1840
rect 194 1835 195 1839
rect 199 1835 200 1839
rect 194 1834 200 1835
rect 450 1839 456 1840
rect 450 1835 451 1839
rect 455 1835 456 1839
rect 450 1834 456 1835
rect 698 1839 704 1840
rect 698 1835 699 1839
rect 703 1835 704 1839
rect 698 1834 704 1835
rect 930 1839 936 1840
rect 930 1835 931 1839
rect 935 1835 936 1839
rect 930 1834 936 1835
rect 1154 1839 1160 1840
rect 1154 1835 1155 1839
rect 1159 1835 1160 1839
rect 1154 1834 1160 1835
rect 1370 1839 1376 1840
rect 1370 1835 1371 1839
rect 1375 1835 1376 1839
rect 1370 1834 1376 1835
rect 1586 1839 1592 1840
rect 1586 1835 1587 1839
rect 1591 1835 1592 1839
rect 1586 1834 1592 1835
rect 1786 1839 1792 1840
rect 1786 1835 1787 1839
rect 1791 1835 1792 1839
rect 1934 1836 1935 1840
rect 1939 1836 1940 1840
rect 1934 1835 1940 1836
rect 3838 1840 3844 1841
rect 5662 1840 5668 1841
rect 3838 1836 3839 1840
rect 3843 1836 3844 1840
rect 3838 1835 3844 1836
rect 4682 1839 4688 1840
rect 4682 1835 4683 1839
rect 4687 1835 4688 1839
rect 1786 1834 1792 1835
rect 4682 1834 4688 1835
rect 4842 1839 4848 1840
rect 4842 1835 4843 1839
rect 4847 1835 4848 1839
rect 4842 1834 4848 1835
rect 5010 1839 5016 1840
rect 5010 1835 5011 1839
rect 5015 1835 5016 1839
rect 5010 1834 5016 1835
rect 5178 1839 5184 1840
rect 5178 1835 5179 1839
rect 5183 1835 5184 1839
rect 5178 1834 5184 1835
rect 5354 1839 5360 1840
rect 5354 1835 5355 1839
rect 5359 1835 5360 1839
rect 5354 1834 5360 1835
rect 5514 1839 5520 1840
rect 5514 1835 5515 1839
rect 5519 1835 5520 1839
rect 5662 1836 5663 1840
rect 5667 1836 5668 1840
rect 5662 1835 5668 1836
rect 5514 1834 5520 1835
rect 222 1824 228 1825
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 222 1820 223 1824
rect 227 1820 228 1824
rect 222 1819 228 1820
rect 478 1824 484 1825
rect 478 1820 479 1824
rect 483 1820 484 1824
rect 478 1819 484 1820
rect 726 1824 732 1825
rect 726 1820 727 1824
rect 731 1820 732 1824
rect 726 1819 732 1820
rect 958 1824 964 1825
rect 958 1820 959 1824
rect 963 1820 964 1824
rect 958 1819 964 1820
rect 1182 1824 1188 1825
rect 1182 1820 1183 1824
rect 1187 1820 1188 1824
rect 1182 1819 1188 1820
rect 1398 1824 1404 1825
rect 1398 1820 1399 1824
rect 1403 1820 1404 1824
rect 1398 1819 1404 1820
rect 1614 1824 1620 1825
rect 1614 1820 1615 1824
rect 1619 1820 1620 1824
rect 1614 1819 1620 1820
rect 1814 1824 1820 1825
rect 4710 1824 4716 1825
rect 1814 1820 1815 1824
rect 1819 1820 1820 1824
rect 1814 1819 1820 1820
rect 1934 1823 1940 1824
rect 1934 1819 1935 1823
rect 1939 1819 1940 1823
rect 110 1818 116 1819
rect 1934 1818 1940 1819
rect 3838 1823 3844 1824
rect 3838 1819 3839 1823
rect 3843 1819 3844 1823
rect 4710 1820 4711 1824
rect 4715 1820 4716 1824
rect 4710 1819 4716 1820
rect 4870 1824 4876 1825
rect 4870 1820 4871 1824
rect 4875 1820 4876 1824
rect 4870 1819 4876 1820
rect 5038 1824 5044 1825
rect 5038 1820 5039 1824
rect 5043 1820 5044 1824
rect 5038 1819 5044 1820
rect 5206 1824 5212 1825
rect 5206 1820 5207 1824
rect 5211 1820 5212 1824
rect 5206 1819 5212 1820
rect 5382 1824 5388 1825
rect 5382 1820 5383 1824
rect 5387 1820 5388 1824
rect 5382 1819 5388 1820
rect 5542 1824 5548 1825
rect 5542 1820 5543 1824
rect 5547 1820 5548 1824
rect 5542 1819 5548 1820
rect 5662 1823 5668 1824
rect 5662 1819 5663 1823
rect 5667 1819 5668 1823
rect 3838 1818 3844 1819
rect 5662 1818 5668 1819
rect 110 1761 116 1762
rect 1934 1761 1940 1762
rect 3838 1761 3844 1762
rect 5662 1761 5668 1762
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 110 1756 116 1757
rect 230 1760 236 1761
rect 230 1756 231 1760
rect 235 1756 236 1760
rect 230 1755 236 1756
rect 446 1760 452 1761
rect 446 1756 447 1760
rect 451 1756 452 1760
rect 446 1755 452 1756
rect 670 1760 676 1761
rect 670 1756 671 1760
rect 675 1756 676 1760
rect 670 1755 676 1756
rect 894 1760 900 1761
rect 894 1756 895 1760
rect 899 1756 900 1760
rect 894 1755 900 1756
rect 1118 1760 1124 1761
rect 1118 1756 1119 1760
rect 1123 1756 1124 1760
rect 1118 1755 1124 1756
rect 1342 1760 1348 1761
rect 1342 1756 1343 1760
rect 1347 1756 1348 1760
rect 1342 1755 1348 1756
rect 1566 1760 1572 1761
rect 1566 1756 1567 1760
rect 1571 1756 1572 1760
rect 1566 1755 1572 1756
rect 1798 1760 1804 1761
rect 1798 1756 1799 1760
rect 1803 1756 1804 1760
rect 1934 1757 1935 1761
rect 1939 1757 1940 1761
rect 1934 1756 1940 1757
rect 1974 1760 1980 1761
rect 3798 1760 3804 1761
rect 1974 1756 1975 1760
rect 1979 1756 1980 1760
rect 1798 1755 1804 1756
rect 1974 1755 1980 1756
rect 2442 1759 2448 1760
rect 2442 1755 2443 1759
rect 2447 1755 2448 1759
rect 2442 1754 2448 1755
rect 2586 1759 2592 1760
rect 2586 1755 2587 1759
rect 2591 1755 2592 1759
rect 2586 1754 2592 1755
rect 2738 1759 2744 1760
rect 2738 1755 2739 1759
rect 2743 1755 2744 1759
rect 2738 1754 2744 1755
rect 2890 1759 2896 1760
rect 2890 1755 2891 1759
rect 2895 1755 2896 1759
rect 2890 1754 2896 1755
rect 3042 1759 3048 1760
rect 3042 1755 3043 1759
rect 3047 1755 3048 1759
rect 3042 1754 3048 1755
rect 3194 1759 3200 1760
rect 3194 1755 3195 1759
rect 3199 1755 3200 1759
rect 3798 1756 3799 1760
rect 3803 1756 3804 1760
rect 3838 1757 3839 1761
rect 3843 1757 3844 1761
rect 3838 1756 3844 1757
rect 3886 1760 3892 1761
rect 3886 1756 3887 1760
rect 3891 1756 3892 1760
rect 3798 1755 3804 1756
rect 3886 1755 3892 1756
rect 4022 1760 4028 1761
rect 4022 1756 4023 1760
rect 4027 1756 4028 1760
rect 4022 1755 4028 1756
rect 4190 1760 4196 1761
rect 4190 1756 4191 1760
rect 4195 1756 4196 1760
rect 4190 1755 4196 1756
rect 4366 1760 4372 1761
rect 4366 1756 4367 1760
rect 4371 1756 4372 1760
rect 4366 1755 4372 1756
rect 4558 1760 4564 1761
rect 4558 1756 4559 1760
rect 4563 1756 4564 1760
rect 4558 1755 4564 1756
rect 4766 1760 4772 1761
rect 4766 1756 4767 1760
rect 4771 1756 4772 1760
rect 4766 1755 4772 1756
rect 4982 1760 4988 1761
rect 4982 1756 4983 1760
rect 4987 1756 4988 1760
rect 4982 1755 4988 1756
rect 5214 1760 5220 1761
rect 5214 1756 5215 1760
rect 5219 1756 5220 1760
rect 5214 1755 5220 1756
rect 5446 1760 5452 1761
rect 5446 1756 5447 1760
rect 5451 1756 5452 1760
rect 5662 1757 5663 1761
rect 5667 1757 5668 1761
rect 5662 1756 5668 1757
rect 5446 1755 5452 1756
rect 3194 1754 3200 1755
rect 202 1745 208 1746
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 202 1741 203 1745
rect 207 1741 208 1745
rect 202 1740 208 1741
rect 418 1745 424 1746
rect 418 1741 419 1745
rect 423 1741 424 1745
rect 418 1740 424 1741
rect 642 1745 648 1746
rect 642 1741 643 1745
rect 647 1741 648 1745
rect 642 1740 648 1741
rect 866 1745 872 1746
rect 866 1741 867 1745
rect 871 1741 872 1745
rect 866 1740 872 1741
rect 1090 1745 1096 1746
rect 1090 1741 1091 1745
rect 1095 1741 1096 1745
rect 1090 1740 1096 1741
rect 1314 1745 1320 1746
rect 1314 1741 1315 1745
rect 1319 1741 1320 1745
rect 1314 1740 1320 1741
rect 1538 1745 1544 1746
rect 1538 1741 1539 1745
rect 1543 1741 1544 1745
rect 1538 1740 1544 1741
rect 1770 1745 1776 1746
rect 3858 1745 3864 1746
rect 1770 1741 1771 1745
rect 1775 1741 1776 1745
rect 1770 1740 1776 1741
rect 1934 1744 1940 1745
rect 2470 1744 2476 1745
rect 1934 1740 1935 1744
rect 1939 1740 1940 1744
rect 110 1739 116 1740
rect 1934 1739 1940 1740
rect 1974 1743 1980 1744
rect 1974 1739 1975 1743
rect 1979 1739 1980 1743
rect 2470 1740 2471 1744
rect 2475 1740 2476 1744
rect 2470 1739 2476 1740
rect 2614 1744 2620 1745
rect 2614 1740 2615 1744
rect 2619 1740 2620 1744
rect 2614 1739 2620 1740
rect 2766 1744 2772 1745
rect 2766 1740 2767 1744
rect 2771 1740 2772 1744
rect 2766 1739 2772 1740
rect 2918 1744 2924 1745
rect 2918 1740 2919 1744
rect 2923 1740 2924 1744
rect 2918 1739 2924 1740
rect 3070 1744 3076 1745
rect 3070 1740 3071 1744
rect 3075 1740 3076 1744
rect 3070 1739 3076 1740
rect 3222 1744 3228 1745
rect 3838 1744 3844 1745
rect 3222 1740 3223 1744
rect 3227 1740 3228 1744
rect 3222 1739 3228 1740
rect 3798 1743 3804 1744
rect 3798 1739 3799 1743
rect 3803 1739 3804 1743
rect 3838 1740 3839 1744
rect 3843 1740 3844 1744
rect 3858 1741 3859 1745
rect 3863 1741 3864 1745
rect 3858 1740 3864 1741
rect 3994 1745 4000 1746
rect 3994 1741 3995 1745
rect 3999 1741 4000 1745
rect 3994 1740 4000 1741
rect 4162 1745 4168 1746
rect 4162 1741 4163 1745
rect 4167 1741 4168 1745
rect 4162 1740 4168 1741
rect 4338 1745 4344 1746
rect 4338 1741 4339 1745
rect 4343 1741 4344 1745
rect 4338 1740 4344 1741
rect 4530 1745 4536 1746
rect 4530 1741 4531 1745
rect 4535 1741 4536 1745
rect 4530 1740 4536 1741
rect 4738 1745 4744 1746
rect 4738 1741 4739 1745
rect 4743 1741 4744 1745
rect 4738 1740 4744 1741
rect 4954 1745 4960 1746
rect 4954 1741 4955 1745
rect 4959 1741 4960 1745
rect 4954 1740 4960 1741
rect 5186 1745 5192 1746
rect 5186 1741 5187 1745
rect 5191 1741 5192 1745
rect 5186 1740 5192 1741
rect 5418 1745 5424 1746
rect 5418 1741 5419 1745
rect 5423 1741 5424 1745
rect 5418 1740 5424 1741
rect 5662 1744 5668 1745
rect 5662 1740 5663 1744
rect 5667 1740 5668 1744
rect 3838 1739 3844 1740
rect 5662 1739 5668 1740
rect 1974 1738 1980 1739
rect 3798 1738 3804 1739
rect 1974 1641 1980 1642
rect 3798 1641 3804 1642
rect 1974 1637 1975 1641
rect 1979 1637 1980 1641
rect 1974 1636 1980 1637
rect 2230 1640 2236 1641
rect 2230 1636 2231 1640
rect 2235 1636 2236 1640
rect 2230 1635 2236 1636
rect 2598 1640 2604 1641
rect 2598 1636 2599 1640
rect 2603 1636 2604 1640
rect 2598 1635 2604 1636
rect 2966 1640 2972 1641
rect 2966 1636 2967 1640
rect 2971 1636 2972 1640
rect 2966 1635 2972 1636
rect 3334 1640 3340 1641
rect 3334 1636 3335 1640
rect 3339 1636 3340 1640
rect 3334 1635 3340 1636
rect 3678 1640 3684 1641
rect 3678 1636 3679 1640
rect 3683 1636 3684 1640
rect 3798 1637 3799 1641
rect 3803 1637 3804 1641
rect 3798 1636 3804 1637
rect 3678 1635 3684 1636
rect 2202 1625 2208 1626
rect 1974 1624 1980 1625
rect 1974 1620 1975 1624
rect 1979 1620 1980 1624
rect 2202 1621 2203 1625
rect 2207 1621 2208 1625
rect 2202 1620 2208 1621
rect 2570 1625 2576 1626
rect 2570 1621 2571 1625
rect 2575 1621 2576 1625
rect 2570 1620 2576 1621
rect 2938 1625 2944 1626
rect 2938 1621 2939 1625
rect 2943 1621 2944 1625
rect 2938 1620 2944 1621
rect 3306 1625 3312 1626
rect 3306 1621 3307 1625
rect 3311 1621 3312 1625
rect 3306 1620 3312 1621
rect 3650 1625 3656 1626
rect 3650 1621 3651 1625
rect 3655 1621 3656 1625
rect 3650 1620 3656 1621
rect 3798 1624 3804 1625
rect 3798 1620 3799 1624
rect 3803 1620 3804 1624
rect 1974 1619 1980 1620
rect 3798 1619 3804 1620
rect 110 1612 116 1613
rect 1934 1612 1940 1613
rect 110 1608 111 1612
rect 115 1608 116 1612
rect 110 1607 116 1608
rect 274 1611 280 1612
rect 274 1607 275 1611
rect 279 1607 280 1611
rect 274 1606 280 1607
rect 458 1611 464 1612
rect 458 1607 459 1611
rect 463 1607 464 1611
rect 458 1606 464 1607
rect 666 1611 672 1612
rect 666 1607 667 1611
rect 671 1607 672 1611
rect 666 1606 672 1607
rect 882 1611 888 1612
rect 882 1607 883 1611
rect 887 1607 888 1611
rect 882 1606 888 1607
rect 1114 1611 1120 1612
rect 1114 1607 1115 1611
rect 1119 1607 1120 1611
rect 1114 1606 1120 1607
rect 1354 1611 1360 1612
rect 1354 1607 1355 1611
rect 1359 1607 1360 1611
rect 1354 1606 1360 1607
rect 1594 1611 1600 1612
rect 1594 1607 1595 1611
rect 1599 1607 1600 1611
rect 1934 1608 1935 1612
rect 1939 1608 1940 1612
rect 1934 1607 1940 1608
rect 3838 1612 3844 1613
rect 5662 1612 5668 1613
rect 3838 1608 3839 1612
rect 3843 1608 3844 1612
rect 3838 1607 3844 1608
rect 3858 1611 3864 1612
rect 3858 1607 3859 1611
rect 3863 1607 3864 1611
rect 1594 1606 1600 1607
rect 3858 1606 3864 1607
rect 3994 1611 4000 1612
rect 3994 1607 3995 1611
rect 3999 1607 4000 1611
rect 3994 1606 4000 1607
rect 4130 1611 4136 1612
rect 4130 1607 4131 1611
rect 4135 1607 4136 1611
rect 4130 1606 4136 1607
rect 4282 1611 4288 1612
rect 4282 1607 4283 1611
rect 4287 1607 4288 1611
rect 4282 1606 4288 1607
rect 4482 1611 4488 1612
rect 4482 1607 4483 1611
rect 4487 1607 4488 1611
rect 4482 1606 4488 1607
rect 4714 1611 4720 1612
rect 4714 1607 4715 1611
rect 4719 1607 4720 1611
rect 4714 1606 4720 1607
rect 4978 1611 4984 1612
rect 4978 1607 4979 1611
rect 4983 1607 4984 1611
rect 4978 1606 4984 1607
rect 5258 1611 5264 1612
rect 5258 1607 5259 1611
rect 5263 1607 5264 1611
rect 5258 1606 5264 1607
rect 5514 1611 5520 1612
rect 5514 1607 5515 1611
rect 5519 1607 5520 1611
rect 5662 1608 5663 1612
rect 5667 1608 5668 1612
rect 5662 1607 5668 1608
rect 5514 1606 5520 1607
rect 302 1596 308 1597
rect 110 1595 116 1596
rect 110 1591 111 1595
rect 115 1591 116 1595
rect 302 1592 303 1596
rect 307 1592 308 1596
rect 302 1591 308 1592
rect 486 1596 492 1597
rect 486 1592 487 1596
rect 491 1592 492 1596
rect 486 1591 492 1592
rect 694 1596 700 1597
rect 694 1592 695 1596
rect 699 1592 700 1596
rect 694 1591 700 1592
rect 910 1596 916 1597
rect 910 1592 911 1596
rect 915 1592 916 1596
rect 910 1591 916 1592
rect 1142 1596 1148 1597
rect 1142 1592 1143 1596
rect 1147 1592 1148 1596
rect 1142 1591 1148 1592
rect 1382 1596 1388 1597
rect 1382 1592 1383 1596
rect 1387 1592 1388 1596
rect 1382 1591 1388 1592
rect 1622 1596 1628 1597
rect 3886 1596 3892 1597
rect 1622 1592 1623 1596
rect 1627 1592 1628 1596
rect 1622 1591 1628 1592
rect 1934 1595 1940 1596
rect 1934 1591 1935 1595
rect 1939 1591 1940 1595
rect 110 1590 116 1591
rect 1934 1590 1940 1591
rect 3838 1595 3844 1596
rect 3838 1591 3839 1595
rect 3843 1591 3844 1595
rect 3886 1592 3887 1596
rect 3891 1592 3892 1596
rect 3886 1591 3892 1592
rect 4022 1596 4028 1597
rect 4022 1592 4023 1596
rect 4027 1592 4028 1596
rect 4022 1591 4028 1592
rect 4158 1596 4164 1597
rect 4158 1592 4159 1596
rect 4163 1592 4164 1596
rect 4158 1591 4164 1592
rect 4310 1596 4316 1597
rect 4310 1592 4311 1596
rect 4315 1592 4316 1596
rect 4310 1591 4316 1592
rect 4510 1596 4516 1597
rect 4510 1592 4511 1596
rect 4515 1592 4516 1596
rect 4510 1591 4516 1592
rect 4742 1596 4748 1597
rect 4742 1592 4743 1596
rect 4747 1592 4748 1596
rect 4742 1591 4748 1592
rect 5006 1596 5012 1597
rect 5006 1592 5007 1596
rect 5011 1592 5012 1596
rect 5006 1591 5012 1592
rect 5286 1596 5292 1597
rect 5286 1592 5287 1596
rect 5291 1592 5292 1596
rect 5286 1591 5292 1592
rect 5542 1596 5548 1597
rect 5542 1592 5543 1596
rect 5547 1592 5548 1596
rect 5542 1591 5548 1592
rect 5662 1595 5668 1596
rect 5662 1591 5663 1595
rect 5667 1591 5668 1595
rect 3838 1590 3844 1591
rect 5662 1590 5668 1591
rect 110 1537 116 1538
rect 1934 1537 1940 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 382 1536 388 1537
rect 382 1532 383 1536
rect 387 1532 388 1536
rect 382 1531 388 1532
rect 574 1536 580 1537
rect 574 1532 575 1536
rect 579 1532 580 1536
rect 574 1531 580 1532
rect 766 1536 772 1537
rect 766 1532 767 1536
rect 771 1532 772 1536
rect 766 1531 772 1532
rect 950 1536 956 1537
rect 950 1532 951 1536
rect 955 1532 956 1536
rect 950 1531 956 1532
rect 1126 1536 1132 1537
rect 1126 1532 1127 1536
rect 1131 1532 1132 1536
rect 1126 1531 1132 1532
rect 1302 1536 1308 1537
rect 1302 1532 1303 1536
rect 1307 1532 1308 1536
rect 1302 1531 1308 1532
rect 1478 1536 1484 1537
rect 1478 1532 1479 1536
rect 1483 1532 1484 1536
rect 1478 1531 1484 1532
rect 1662 1536 1668 1537
rect 1662 1532 1663 1536
rect 1667 1532 1668 1536
rect 1934 1533 1935 1537
rect 1939 1533 1940 1537
rect 1934 1532 1940 1533
rect 3838 1537 3844 1538
rect 5662 1537 5668 1538
rect 3838 1533 3839 1537
rect 3843 1533 3844 1537
rect 3838 1532 3844 1533
rect 3886 1536 3892 1537
rect 3886 1532 3887 1536
rect 3891 1532 3892 1536
rect 1662 1531 1668 1532
rect 3886 1531 3892 1532
rect 4046 1536 4052 1537
rect 4046 1532 4047 1536
rect 4051 1532 4052 1536
rect 4046 1531 4052 1532
rect 4270 1536 4276 1537
rect 4270 1532 4271 1536
rect 4275 1532 4276 1536
rect 4270 1531 4276 1532
rect 4542 1536 4548 1537
rect 4542 1532 4543 1536
rect 4547 1532 4548 1536
rect 4542 1531 4548 1532
rect 4854 1536 4860 1537
rect 4854 1532 4855 1536
rect 4859 1532 4860 1536
rect 4854 1531 4860 1532
rect 5190 1536 5196 1537
rect 5190 1532 5191 1536
rect 5195 1532 5196 1536
rect 5190 1531 5196 1532
rect 5526 1536 5532 1537
rect 5526 1532 5527 1536
rect 5531 1532 5532 1536
rect 5662 1533 5663 1537
rect 5667 1533 5668 1537
rect 5662 1532 5668 1533
rect 5526 1531 5532 1532
rect 354 1521 360 1522
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 354 1517 355 1521
rect 359 1517 360 1521
rect 354 1516 360 1517
rect 546 1521 552 1522
rect 546 1517 547 1521
rect 551 1517 552 1521
rect 546 1516 552 1517
rect 738 1521 744 1522
rect 738 1517 739 1521
rect 743 1517 744 1521
rect 738 1516 744 1517
rect 922 1521 928 1522
rect 922 1517 923 1521
rect 927 1517 928 1521
rect 922 1516 928 1517
rect 1098 1521 1104 1522
rect 1098 1517 1099 1521
rect 1103 1517 1104 1521
rect 1098 1516 1104 1517
rect 1274 1521 1280 1522
rect 1274 1517 1275 1521
rect 1279 1517 1280 1521
rect 1274 1516 1280 1517
rect 1450 1521 1456 1522
rect 1450 1517 1451 1521
rect 1455 1517 1456 1521
rect 1450 1516 1456 1517
rect 1634 1521 1640 1522
rect 3858 1521 3864 1522
rect 1634 1517 1635 1521
rect 1639 1517 1640 1521
rect 1634 1516 1640 1517
rect 1934 1520 1940 1521
rect 1934 1516 1935 1520
rect 1939 1516 1940 1520
rect 110 1515 116 1516
rect 1934 1515 1940 1516
rect 3838 1520 3844 1521
rect 3838 1516 3839 1520
rect 3843 1516 3844 1520
rect 3858 1517 3859 1521
rect 3863 1517 3864 1521
rect 3858 1516 3864 1517
rect 4018 1521 4024 1522
rect 4018 1517 4019 1521
rect 4023 1517 4024 1521
rect 4018 1516 4024 1517
rect 4242 1521 4248 1522
rect 4242 1517 4243 1521
rect 4247 1517 4248 1521
rect 4242 1516 4248 1517
rect 4514 1521 4520 1522
rect 4514 1517 4515 1521
rect 4519 1517 4520 1521
rect 4514 1516 4520 1517
rect 4826 1521 4832 1522
rect 4826 1517 4827 1521
rect 4831 1517 4832 1521
rect 4826 1516 4832 1517
rect 5162 1521 5168 1522
rect 5162 1517 5163 1521
rect 5167 1517 5168 1521
rect 5162 1516 5168 1517
rect 5498 1521 5504 1522
rect 5498 1517 5499 1521
rect 5503 1517 5504 1521
rect 5498 1516 5504 1517
rect 5662 1520 5668 1521
rect 5662 1516 5663 1520
rect 5667 1516 5668 1520
rect 3838 1515 3844 1516
rect 5662 1515 5668 1516
rect 1974 1480 1980 1481
rect 3798 1480 3804 1481
rect 1974 1476 1975 1480
rect 1979 1476 1980 1480
rect 1974 1475 1980 1476
rect 1994 1479 2000 1480
rect 1994 1475 1995 1479
rect 1999 1475 2000 1479
rect 1994 1474 2000 1475
rect 2274 1479 2280 1480
rect 2274 1475 2275 1479
rect 2279 1475 2280 1479
rect 2274 1474 2280 1475
rect 2538 1479 2544 1480
rect 2538 1475 2539 1479
rect 2543 1475 2544 1479
rect 2538 1474 2544 1475
rect 2778 1479 2784 1480
rect 2778 1475 2779 1479
rect 2783 1475 2784 1479
rect 2778 1474 2784 1475
rect 3010 1479 3016 1480
rect 3010 1475 3011 1479
rect 3015 1475 3016 1479
rect 3010 1474 3016 1475
rect 3234 1479 3240 1480
rect 3234 1475 3235 1479
rect 3239 1475 3240 1479
rect 3234 1474 3240 1475
rect 3450 1479 3456 1480
rect 3450 1475 3451 1479
rect 3455 1475 3456 1479
rect 3450 1474 3456 1475
rect 3650 1479 3656 1480
rect 3650 1475 3651 1479
rect 3655 1475 3656 1479
rect 3798 1476 3799 1480
rect 3803 1476 3804 1480
rect 3798 1475 3804 1476
rect 3650 1474 3656 1475
rect 2022 1464 2028 1465
rect 1974 1463 1980 1464
rect 1974 1459 1975 1463
rect 1979 1459 1980 1463
rect 2022 1460 2023 1464
rect 2027 1460 2028 1464
rect 2022 1459 2028 1460
rect 2302 1464 2308 1465
rect 2302 1460 2303 1464
rect 2307 1460 2308 1464
rect 2302 1459 2308 1460
rect 2566 1464 2572 1465
rect 2566 1460 2567 1464
rect 2571 1460 2572 1464
rect 2566 1459 2572 1460
rect 2806 1464 2812 1465
rect 2806 1460 2807 1464
rect 2811 1460 2812 1464
rect 2806 1459 2812 1460
rect 3038 1464 3044 1465
rect 3038 1460 3039 1464
rect 3043 1460 3044 1464
rect 3038 1459 3044 1460
rect 3262 1464 3268 1465
rect 3262 1460 3263 1464
rect 3267 1460 3268 1464
rect 3262 1459 3268 1460
rect 3478 1464 3484 1465
rect 3478 1460 3479 1464
rect 3483 1460 3484 1464
rect 3478 1459 3484 1460
rect 3678 1464 3684 1465
rect 3678 1460 3679 1464
rect 3683 1460 3684 1464
rect 3678 1459 3684 1460
rect 3798 1463 3804 1464
rect 3798 1459 3799 1463
rect 3803 1459 3804 1463
rect 1974 1458 1980 1459
rect 3798 1458 3804 1459
rect 1974 1405 1980 1406
rect 3798 1405 3804 1406
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2022 1404 2028 1405
rect 2022 1400 2023 1404
rect 2027 1400 2028 1404
rect 2022 1399 2028 1400
rect 2190 1404 2196 1405
rect 2190 1400 2191 1404
rect 2195 1400 2196 1404
rect 2190 1399 2196 1400
rect 2398 1404 2404 1405
rect 2398 1400 2399 1404
rect 2403 1400 2404 1404
rect 2398 1399 2404 1400
rect 2614 1404 2620 1405
rect 2614 1400 2615 1404
rect 2619 1400 2620 1404
rect 2614 1399 2620 1400
rect 2830 1404 2836 1405
rect 2830 1400 2831 1404
rect 2835 1400 2836 1404
rect 2830 1399 2836 1400
rect 3054 1404 3060 1405
rect 3054 1400 3055 1404
rect 3059 1400 3060 1404
rect 3054 1399 3060 1400
rect 3286 1404 3292 1405
rect 3286 1400 3287 1404
rect 3291 1400 3292 1404
rect 3286 1399 3292 1400
rect 3526 1404 3532 1405
rect 3526 1400 3527 1404
rect 3531 1400 3532 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3798 1400 3804 1401
rect 3526 1399 3532 1400
rect 1994 1389 2000 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 1994 1385 1995 1389
rect 1999 1385 2000 1389
rect 1994 1384 2000 1385
rect 2162 1389 2168 1390
rect 2162 1385 2163 1389
rect 2167 1385 2168 1389
rect 2162 1384 2168 1385
rect 2370 1389 2376 1390
rect 2370 1385 2371 1389
rect 2375 1385 2376 1389
rect 2370 1384 2376 1385
rect 2586 1389 2592 1390
rect 2586 1385 2587 1389
rect 2591 1385 2592 1389
rect 2586 1384 2592 1385
rect 2802 1389 2808 1390
rect 2802 1385 2803 1389
rect 2807 1385 2808 1389
rect 2802 1384 2808 1385
rect 3026 1389 3032 1390
rect 3026 1385 3027 1389
rect 3031 1385 3032 1389
rect 3026 1384 3032 1385
rect 3258 1389 3264 1390
rect 3258 1385 3259 1389
rect 3263 1385 3264 1389
rect 3258 1384 3264 1385
rect 3498 1389 3504 1390
rect 3498 1385 3499 1389
rect 3503 1385 3504 1389
rect 3498 1384 3504 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 1974 1383 1980 1384
rect 3798 1383 3804 1384
rect 3838 1372 3844 1373
rect 5662 1372 5668 1373
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 330 1367 336 1368
rect 330 1363 331 1367
rect 335 1363 336 1367
rect 330 1362 336 1363
rect 586 1367 592 1368
rect 586 1363 587 1367
rect 591 1363 592 1367
rect 586 1362 592 1363
rect 842 1367 848 1368
rect 842 1363 843 1367
rect 847 1363 848 1367
rect 842 1362 848 1363
rect 1098 1367 1104 1368
rect 1098 1363 1099 1367
rect 1103 1363 1104 1367
rect 1098 1362 1104 1363
rect 1362 1367 1368 1368
rect 1362 1363 1363 1367
rect 1367 1363 1368 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 3838 1368 3839 1372
rect 3843 1368 3844 1372
rect 3838 1367 3844 1368
rect 3858 1371 3864 1372
rect 3858 1367 3859 1371
rect 3863 1367 3864 1371
rect 3858 1366 3864 1367
rect 3994 1371 4000 1372
rect 3994 1367 3995 1371
rect 3999 1367 4000 1371
rect 3994 1366 4000 1367
rect 4146 1371 4152 1372
rect 4146 1367 4147 1371
rect 4151 1367 4152 1371
rect 4146 1366 4152 1367
rect 4354 1371 4360 1372
rect 4354 1367 4355 1371
rect 4359 1367 4360 1371
rect 4354 1366 4360 1367
rect 4594 1371 4600 1372
rect 4594 1367 4595 1371
rect 4599 1367 4600 1371
rect 4594 1366 4600 1367
rect 4866 1371 4872 1372
rect 4866 1367 4867 1371
rect 4871 1367 4872 1371
rect 4866 1366 4872 1367
rect 5162 1371 5168 1372
rect 5162 1367 5163 1371
rect 5167 1367 5168 1371
rect 5162 1366 5168 1367
rect 5458 1371 5464 1372
rect 5458 1367 5459 1371
rect 5463 1367 5464 1371
rect 5662 1368 5663 1372
rect 5667 1368 5668 1372
rect 5662 1367 5668 1368
rect 5458 1366 5464 1367
rect 1934 1363 1940 1364
rect 1362 1362 1368 1363
rect 3886 1356 3892 1357
rect 3838 1355 3844 1356
rect 358 1352 364 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 358 1348 359 1352
rect 363 1348 364 1352
rect 358 1347 364 1348
rect 614 1352 620 1353
rect 614 1348 615 1352
rect 619 1348 620 1352
rect 614 1347 620 1348
rect 870 1352 876 1353
rect 870 1348 871 1352
rect 875 1348 876 1352
rect 870 1347 876 1348
rect 1126 1352 1132 1353
rect 1126 1348 1127 1352
rect 1131 1348 1132 1352
rect 1126 1347 1132 1348
rect 1390 1352 1396 1353
rect 1390 1348 1391 1352
rect 1395 1348 1396 1352
rect 1390 1347 1396 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 3838 1351 3839 1355
rect 3843 1351 3844 1355
rect 3886 1352 3887 1356
rect 3891 1352 3892 1356
rect 3886 1351 3892 1352
rect 4022 1356 4028 1357
rect 4022 1352 4023 1356
rect 4027 1352 4028 1356
rect 4022 1351 4028 1352
rect 4174 1356 4180 1357
rect 4174 1352 4175 1356
rect 4179 1352 4180 1356
rect 4174 1351 4180 1352
rect 4382 1356 4388 1357
rect 4382 1352 4383 1356
rect 4387 1352 4388 1356
rect 4382 1351 4388 1352
rect 4622 1356 4628 1357
rect 4622 1352 4623 1356
rect 4627 1352 4628 1356
rect 4622 1351 4628 1352
rect 4894 1356 4900 1357
rect 4894 1352 4895 1356
rect 4899 1352 4900 1356
rect 4894 1351 4900 1352
rect 5190 1356 5196 1357
rect 5190 1352 5191 1356
rect 5195 1352 5196 1356
rect 5190 1351 5196 1352
rect 5486 1356 5492 1357
rect 5486 1352 5487 1356
rect 5491 1352 5492 1356
rect 5486 1351 5492 1352
rect 5662 1355 5668 1356
rect 5662 1351 5663 1355
rect 5667 1351 5668 1355
rect 3838 1350 3844 1351
rect 5662 1350 5668 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 366 1292 372 1293
rect 366 1288 367 1292
rect 371 1288 372 1292
rect 366 1287 372 1288
rect 550 1292 556 1293
rect 550 1288 551 1292
rect 555 1288 556 1292
rect 550 1287 556 1288
rect 726 1292 732 1293
rect 726 1288 727 1292
rect 731 1288 732 1292
rect 726 1287 732 1288
rect 894 1292 900 1293
rect 894 1288 895 1292
rect 899 1288 900 1292
rect 894 1287 900 1288
rect 1062 1292 1068 1293
rect 1062 1288 1063 1292
rect 1067 1288 1068 1292
rect 1062 1287 1068 1288
rect 1222 1292 1228 1293
rect 1222 1288 1223 1292
rect 1227 1288 1228 1292
rect 1222 1287 1228 1288
rect 1374 1292 1380 1293
rect 1374 1288 1375 1292
rect 1379 1288 1380 1292
rect 1374 1287 1380 1288
rect 1526 1292 1532 1293
rect 1526 1288 1527 1292
rect 1531 1288 1532 1292
rect 1526 1287 1532 1288
rect 1678 1292 1684 1293
rect 1678 1288 1679 1292
rect 1683 1288 1684 1292
rect 1678 1287 1684 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 3838 1293 3844 1294
rect 5662 1293 5668 1294
rect 3838 1289 3839 1293
rect 3843 1289 3844 1293
rect 3838 1288 3844 1289
rect 3886 1292 3892 1293
rect 3886 1288 3887 1292
rect 3891 1288 3892 1292
rect 1814 1287 1820 1288
rect 3886 1287 3892 1288
rect 4046 1292 4052 1293
rect 4046 1288 4047 1292
rect 4051 1288 4052 1292
rect 4046 1287 4052 1288
rect 4238 1292 4244 1293
rect 4238 1288 4239 1292
rect 4243 1288 4244 1292
rect 4238 1287 4244 1288
rect 4454 1292 4460 1293
rect 4454 1288 4455 1292
rect 4459 1288 4460 1292
rect 4454 1287 4460 1288
rect 4694 1292 4700 1293
rect 4694 1288 4695 1292
rect 4699 1288 4700 1292
rect 4694 1287 4700 1288
rect 4950 1292 4956 1293
rect 4950 1288 4951 1292
rect 4955 1288 4956 1292
rect 4950 1287 4956 1288
rect 5222 1292 5228 1293
rect 5222 1288 5223 1292
rect 5227 1288 5228 1292
rect 5222 1287 5228 1288
rect 5494 1292 5500 1293
rect 5494 1288 5495 1292
rect 5499 1288 5500 1292
rect 5662 1289 5663 1293
rect 5667 1289 5668 1293
rect 5662 1288 5668 1289
rect 5494 1287 5500 1288
rect 338 1277 344 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 338 1273 339 1277
rect 343 1273 344 1277
rect 338 1272 344 1273
rect 522 1277 528 1278
rect 522 1273 523 1277
rect 527 1273 528 1277
rect 522 1272 528 1273
rect 698 1277 704 1278
rect 698 1273 699 1277
rect 703 1273 704 1277
rect 698 1272 704 1273
rect 866 1277 872 1278
rect 866 1273 867 1277
rect 871 1273 872 1277
rect 866 1272 872 1273
rect 1034 1277 1040 1278
rect 1034 1273 1035 1277
rect 1039 1273 1040 1277
rect 1034 1272 1040 1273
rect 1194 1277 1200 1278
rect 1194 1273 1195 1277
rect 1199 1273 1200 1277
rect 1194 1272 1200 1273
rect 1346 1277 1352 1278
rect 1346 1273 1347 1277
rect 1351 1273 1352 1277
rect 1346 1272 1352 1273
rect 1498 1277 1504 1278
rect 1498 1273 1499 1277
rect 1503 1273 1504 1277
rect 1498 1272 1504 1273
rect 1650 1277 1656 1278
rect 1650 1273 1651 1277
rect 1655 1273 1656 1277
rect 1650 1272 1656 1273
rect 1786 1277 1792 1278
rect 3858 1277 3864 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 3838 1276 3844 1277
rect 3838 1272 3839 1276
rect 3843 1272 3844 1276
rect 3858 1273 3859 1277
rect 3863 1273 3864 1277
rect 3858 1272 3864 1273
rect 4018 1277 4024 1278
rect 4018 1273 4019 1277
rect 4023 1273 4024 1277
rect 4018 1272 4024 1273
rect 4210 1277 4216 1278
rect 4210 1273 4211 1277
rect 4215 1273 4216 1277
rect 4210 1272 4216 1273
rect 4426 1277 4432 1278
rect 4426 1273 4427 1277
rect 4431 1273 4432 1277
rect 4426 1272 4432 1273
rect 4666 1277 4672 1278
rect 4666 1273 4667 1277
rect 4671 1273 4672 1277
rect 4666 1272 4672 1273
rect 4922 1277 4928 1278
rect 4922 1273 4923 1277
rect 4927 1273 4928 1277
rect 4922 1272 4928 1273
rect 5194 1277 5200 1278
rect 5194 1273 5195 1277
rect 5199 1273 5200 1277
rect 5194 1272 5200 1273
rect 5466 1277 5472 1278
rect 5466 1273 5467 1277
rect 5471 1273 5472 1277
rect 5466 1272 5472 1273
rect 5662 1276 5668 1277
rect 5662 1272 5663 1276
rect 5667 1272 5668 1276
rect 3838 1271 3844 1272
rect 5662 1271 5668 1272
rect 1974 1236 1980 1237
rect 3798 1236 3804 1237
rect 1974 1232 1975 1236
rect 1979 1232 1980 1236
rect 1974 1231 1980 1232
rect 3090 1235 3096 1236
rect 3090 1231 3091 1235
rect 3095 1231 3096 1235
rect 3090 1230 3096 1231
rect 3226 1235 3232 1236
rect 3226 1231 3227 1235
rect 3231 1231 3232 1235
rect 3226 1230 3232 1231
rect 3362 1235 3368 1236
rect 3362 1231 3363 1235
rect 3367 1231 3368 1235
rect 3798 1232 3799 1236
rect 3803 1232 3804 1236
rect 3798 1231 3804 1232
rect 3362 1230 3368 1231
rect 3118 1220 3124 1221
rect 1974 1219 1980 1220
rect 1974 1215 1975 1219
rect 1979 1215 1980 1219
rect 3118 1216 3119 1220
rect 3123 1216 3124 1220
rect 3118 1215 3124 1216
rect 3254 1220 3260 1221
rect 3254 1216 3255 1220
rect 3259 1216 3260 1220
rect 3254 1215 3260 1216
rect 3390 1220 3396 1221
rect 3390 1216 3391 1220
rect 3395 1216 3396 1220
rect 3390 1215 3396 1216
rect 3798 1219 3804 1220
rect 3798 1215 3799 1219
rect 3803 1215 3804 1219
rect 1974 1214 1980 1215
rect 3798 1214 3804 1215
rect 1974 1161 1980 1162
rect 3798 1161 3804 1162
rect 1974 1157 1975 1161
rect 1979 1157 1980 1161
rect 1974 1156 1980 1157
rect 2982 1160 2988 1161
rect 2982 1156 2983 1160
rect 2987 1156 2988 1160
rect 2982 1155 2988 1156
rect 3118 1160 3124 1161
rect 3118 1156 3119 1160
rect 3123 1156 3124 1160
rect 3118 1155 3124 1156
rect 3254 1160 3260 1161
rect 3254 1156 3255 1160
rect 3259 1156 3260 1160
rect 3798 1157 3799 1161
rect 3803 1157 3804 1161
rect 3798 1156 3804 1157
rect 3254 1155 3260 1156
rect 2954 1145 2960 1146
rect 1974 1144 1980 1145
rect 1974 1140 1975 1144
rect 1979 1140 1980 1144
rect 2954 1141 2955 1145
rect 2959 1141 2960 1145
rect 2954 1140 2960 1141
rect 3090 1145 3096 1146
rect 3090 1141 3091 1145
rect 3095 1141 3096 1145
rect 3090 1140 3096 1141
rect 3226 1145 3232 1146
rect 3226 1141 3227 1145
rect 3231 1141 3232 1145
rect 3226 1140 3232 1141
rect 3798 1144 3804 1145
rect 3798 1140 3799 1144
rect 3803 1140 3804 1144
rect 1974 1139 1980 1140
rect 3798 1139 3804 1140
rect 3838 1136 3844 1137
rect 5662 1136 5668 1137
rect 110 1132 116 1133
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 234 1131 240 1132
rect 234 1127 235 1131
rect 239 1127 240 1131
rect 234 1126 240 1127
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1127 384 1131
rect 378 1126 384 1127
rect 522 1131 528 1132
rect 522 1127 523 1131
rect 527 1127 528 1131
rect 522 1126 528 1127
rect 666 1131 672 1132
rect 666 1127 667 1131
rect 671 1127 672 1131
rect 666 1126 672 1127
rect 810 1131 816 1132
rect 810 1127 811 1131
rect 815 1127 816 1131
rect 810 1126 816 1127
rect 946 1131 952 1132
rect 946 1127 947 1131
rect 951 1127 952 1131
rect 946 1126 952 1127
rect 1090 1131 1096 1132
rect 1090 1127 1091 1131
rect 1095 1127 1096 1131
rect 1090 1126 1096 1127
rect 1234 1131 1240 1132
rect 1234 1127 1235 1131
rect 1239 1127 1240 1131
rect 1234 1126 1240 1127
rect 1378 1131 1384 1132
rect 1378 1127 1379 1131
rect 1383 1127 1384 1131
rect 1378 1126 1384 1127
rect 1514 1131 1520 1132
rect 1514 1127 1515 1131
rect 1519 1127 1520 1131
rect 1514 1126 1520 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 3838 1132 3839 1136
rect 3843 1132 3844 1136
rect 3838 1131 3844 1132
rect 3858 1135 3864 1136
rect 3858 1131 3859 1135
rect 3863 1131 3864 1135
rect 3858 1130 3864 1131
rect 4090 1135 4096 1136
rect 4090 1131 4091 1135
rect 4095 1131 4096 1135
rect 4090 1130 4096 1131
rect 4338 1135 4344 1136
rect 4338 1131 4339 1135
rect 4343 1131 4344 1135
rect 4338 1130 4344 1131
rect 4578 1135 4584 1136
rect 4578 1131 4579 1135
rect 4583 1131 4584 1135
rect 4578 1130 4584 1131
rect 4810 1135 4816 1136
rect 4810 1131 4811 1135
rect 4815 1131 4816 1135
rect 4810 1130 4816 1131
rect 5042 1135 5048 1136
rect 5042 1131 5043 1135
rect 5047 1131 5048 1135
rect 5042 1130 5048 1131
rect 5274 1135 5280 1136
rect 5274 1131 5275 1135
rect 5279 1131 5280 1135
rect 5274 1130 5280 1131
rect 5514 1135 5520 1136
rect 5514 1131 5515 1135
rect 5519 1131 5520 1135
rect 5662 1132 5663 1136
rect 5667 1132 5668 1136
rect 5662 1131 5668 1132
rect 5514 1130 5520 1131
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 3886 1120 3892 1121
rect 3838 1119 3844 1120
rect 262 1116 268 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 262 1112 263 1116
rect 267 1112 268 1116
rect 262 1111 268 1112
rect 406 1116 412 1117
rect 406 1112 407 1116
rect 411 1112 412 1116
rect 406 1111 412 1112
rect 550 1116 556 1117
rect 550 1112 551 1116
rect 555 1112 556 1116
rect 550 1111 556 1112
rect 694 1116 700 1117
rect 694 1112 695 1116
rect 699 1112 700 1116
rect 694 1111 700 1112
rect 838 1116 844 1117
rect 838 1112 839 1116
rect 843 1112 844 1116
rect 838 1111 844 1112
rect 974 1116 980 1117
rect 974 1112 975 1116
rect 979 1112 980 1116
rect 974 1111 980 1112
rect 1118 1116 1124 1117
rect 1118 1112 1119 1116
rect 1123 1112 1124 1116
rect 1118 1111 1124 1112
rect 1262 1116 1268 1117
rect 1262 1112 1263 1116
rect 1267 1112 1268 1116
rect 1262 1111 1268 1112
rect 1406 1116 1412 1117
rect 1406 1112 1407 1116
rect 1411 1112 1412 1116
rect 1406 1111 1412 1112
rect 1542 1116 1548 1117
rect 1542 1112 1543 1116
rect 1547 1112 1548 1116
rect 1542 1111 1548 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 3838 1115 3839 1119
rect 3843 1115 3844 1119
rect 3886 1116 3887 1120
rect 3891 1116 3892 1120
rect 3886 1115 3892 1116
rect 4118 1120 4124 1121
rect 4118 1116 4119 1120
rect 4123 1116 4124 1120
rect 4118 1115 4124 1116
rect 4366 1120 4372 1121
rect 4366 1116 4367 1120
rect 4371 1116 4372 1120
rect 4366 1115 4372 1116
rect 4606 1120 4612 1121
rect 4606 1116 4607 1120
rect 4611 1116 4612 1120
rect 4606 1115 4612 1116
rect 4838 1120 4844 1121
rect 4838 1116 4839 1120
rect 4843 1116 4844 1120
rect 4838 1115 4844 1116
rect 5070 1120 5076 1121
rect 5070 1116 5071 1120
rect 5075 1116 5076 1120
rect 5070 1115 5076 1116
rect 5302 1120 5308 1121
rect 5302 1116 5303 1120
rect 5307 1116 5308 1120
rect 5302 1115 5308 1116
rect 5542 1120 5548 1121
rect 5542 1116 5543 1120
rect 5547 1116 5548 1120
rect 5542 1115 5548 1116
rect 5662 1119 5668 1120
rect 5662 1115 5663 1119
rect 5667 1115 5668 1119
rect 3838 1114 3844 1115
rect 5662 1114 5668 1115
rect 110 1110 116 1111
rect 1934 1110 1940 1111
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 462 1044 468 1045
rect 462 1040 463 1044
rect 467 1040 468 1044
rect 462 1039 468 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 870 1044 876 1045
rect 870 1040 871 1044
rect 875 1040 876 1044
rect 870 1039 876 1040
rect 1078 1044 1084 1045
rect 1078 1040 1079 1044
rect 1083 1040 1084 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 3838 1041 3844 1042
rect 5662 1041 5668 1042
rect 1078 1039 1084 1040
rect 3838 1037 3839 1041
rect 3843 1037 3844 1041
rect 3838 1036 3844 1037
rect 4862 1040 4868 1041
rect 4862 1036 4863 1040
rect 4867 1036 4868 1040
rect 4862 1035 4868 1036
rect 4998 1040 5004 1041
rect 4998 1036 4999 1040
rect 5003 1036 5004 1040
rect 4998 1035 5004 1036
rect 5134 1040 5140 1041
rect 5134 1036 5135 1040
rect 5139 1036 5140 1040
rect 5134 1035 5140 1036
rect 5270 1040 5276 1041
rect 5270 1036 5271 1040
rect 5275 1036 5276 1040
rect 5270 1035 5276 1036
rect 5406 1040 5412 1041
rect 5406 1036 5407 1040
rect 5411 1036 5412 1040
rect 5406 1035 5412 1036
rect 5542 1040 5548 1041
rect 5542 1036 5543 1040
rect 5547 1036 5548 1040
rect 5662 1037 5663 1041
rect 5667 1037 5668 1041
rect 5662 1036 5668 1037
rect 5542 1035 5548 1036
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 434 1029 440 1030
rect 434 1025 435 1029
rect 439 1025 440 1029
rect 434 1024 440 1025
rect 634 1029 640 1030
rect 634 1025 635 1029
rect 639 1025 640 1029
rect 634 1024 640 1025
rect 842 1029 848 1030
rect 842 1025 843 1029
rect 847 1025 848 1029
rect 842 1024 848 1025
rect 1050 1029 1056 1030
rect 1050 1025 1051 1029
rect 1055 1025 1056 1029
rect 1050 1024 1056 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 4834 1025 4840 1026
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 3838 1024 3844 1025
rect 3838 1020 3839 1024
rect 3843 1020 3844 1024
rect 4834 1021 4835 1025
rect 4839 1021 4840 1025
rect 4834 1020 4840 1021
rect 4970 1025 4976 1026
rect 4970 1021 4971 1025
rect 4975 1021 4976 1025
rect 4970 1020 4976 1021
rect 5106 1025 5112 1026
rect 5106 1021 5107 1025
rect 5111 1021 5112 1025
rect 5106 1020 5112 1021
rect 5242 1025 5248 1026
rect 5242 1021 5243 1025
rect 5247 1021 5248 1025
rect 5242 1020 5248 1021
rect 5378 1025 5384 1026
rect 5378 1021 5379 1025
rect 5383 1021 5384 1025
rect 5378 1020 5384 1021
rect 5514 1025 5520 1026
rect 5514 1021 5515 1025
rect 5519 1021 5520 1025
rect 5514 1020 5520 1021
rect 5662 1024 5668 1025
rect 5662 1020 5663 1024
rect 5667 1020 5668 1024
rect 3838 1019 3844 1020
rect 5662 1019 5668 1020
rect 1974 1012 1980 1013
rect 3798 1012 3804 1013
rect 1974 1008 1975 1012
rect 1979 1008 1980 1012
rect 1974 1007 1980 1008
rect 1994 1011 2000 1012
rect 1994 1007 1995 1011
rect 1999 1007 2000 1011
rect 1994 1006 2000 1007
rect 2130 1011 2136 1012
rect 2130 1007 2131 1011
rect 2135 1007 2136 1011
rect 2130 1006 2136 1007
rect 2274 1011 2280 1012
rect 2274 1007 2275 1011
rect 2279 1007 2280 1011
rect 2274 1006 2280 1007
rect 2442 1011 2448 1012
rect 2442 1007 2443 1011
rect 2447 1007 2448 1011
rect 2442 1006 2448 1007
rect 2626 1011 2632 1012
rect 2626 1007 2627 1011
rect 2631 1007 2632 1011
rect 2626 1006 2632 1007
rect 2818 1011 2824 1012
rect 2818 1007 2819 1011
rect 2823 1007 2824 1011
rect 2818 1006 2824 1007
rect 3026 1011 3032 1012
rect 3026 1007 3027 1011
rect 3031 1007 3032 1011
rect 3026 1006 3032 1007
rect 3234 1011 3240 1012
rect 3234 1007 3235 1011
rect 3239 1007 3240 1011
rect 3234 1006 3240 1007
rect 3450 1011 3456 1012
rect 3450 1007 3451 1011
rect 3455 1007 3456 1011
rect 3450 1006 3456 1007
rect 3650 1011 3656 1012
rect 3650 1007 3651 1011
rect 3655 1007 3656 1011
rect 3798 1008 3799 1012
rect 3803 1008 3804 1012
rect 3798 1007 3804 1008
rect 3650 1006 3656 1007
rect 2022 996 2028 997
rect 1974 995 1980 996
rect 1974 991 1975 995
rect 1979 991 1980 995
rect 2022 992 2023 996
rect 2027 992 2028 996
rect 2022 991 2028 992
rect 2158 996 2164 997
rect 2158 992 2159 996
rect 2163 992 2164 996
rect 2158 991 2164 992
rect 2302 996 2308 997
rect 2302 992 2303 996
rect 2307 992 2308 996
rect 2302 991 2308 992
rect 2470 996 2476 997
rect 2470 992 2471 996
rect 2475 992 2476 996
rect 2470 991 2476 992
rect 2654 996 2660 997
rect 2654 992 2655 996
rect 2659 992 2660 996
rect 2654 991 2660 992
rect 2846 996 2852 997
rect 2846 992 2847 996
rect 2851 992 2852 996
rect 2846 991 2852 992
rect 3054 996 3060 997
rect 3054 992 3055 996
rect 3059 992 3060 996
rect 3054 991 3060 992
rect 3262 996 3268 997
rect 3262 992 3263 996
rect 3267 992 3268 996
rect 3262 991 3268 992
rect 3478 996 3484 997
rect 3478 992 3479 996
rect 3483 992 3484 996
rect 3478 991 3484 992
rect 3678 996 3684 997
rect 3678 992 3679 996
rect 3683 992 3684 996
rect 3678 991 3684 992
rect 3798 995 3804 996
rect 3798 991 3799 995
rect 3803 991 3804 995
rect 1974 990 1980 991
rect 3798 990 3804 991
rect 1974 937 1980 938
rect 3798 937 3804 938
rect 1974 933 1975 937
rect 1979 933 1980 937
rect 1974 932 1980 933
rect 2094 936 2100 937
rect 2094 932 2095 936
rect 2099 932 2100 936
rect 2094 931 2100 932
rect 2230 936 2236 937
rect 2230 932 2231 936
rect 2235 932 2236 936
rect 2230 931 2236 932
rect 2366 936 2372 937
rect 2366 932 2367 936
rect 2371 932 2372 936
rect 2366 931 2372 932
rect 2502 936 2508 937
rect 2502 932 2503 936
rect 2507 932 2508 936
rect 2502 931 2508 932
rect 2654 936 2660 937
rect 2654 932 2655 936
rect 2659 932 2660 936
rect 2654 931 2660 932
rect 2830 936 2836 937
rect 2830 932 2831 936
rect 2835 932 2836 936
rect 2830 931 2836 932
rect 3022 936 3028 937
rect 3022 932 3023 936
rect 3027 932 3028 936
rect 3022 931 3028 932
rect 3230 936 3236 937
rect 3230 932 3231 936
rect 3235 932 3236 936
rect 3230 931 3236 932
rect 3454 936 3460 937
rect 3454 932 3455 936
rect 3459 932 3460 936
rect 3454 931 3460 932
rect 3678 936 3684 937
rect 3678 932 3679 936
rect 3683 932 3684 936
rect 3798 933 3799 937
rect 3803 933 3804 937
rect 3798 932 3804 933
rect 3678 931 3684 932
rect 2066 921 2072 922
rect 1974 920 1980 921
rect 1974 916 1975 920
rect 1979 916 1980 920
rect 2066 917 2067 921
rect 2071 917 2072 921
rect 2066 916 2072 917
rect 2202 921 2208 922
rect 2202 917 2203 921
rect 2207 917 2208 921
rect 2202 916 2208 917
rect 2338 921 2344 922
rect 2338 917 2339 921
rect 2343 917 2344 921
rect 2338 916 2344 917
rect 2474 921 2480 922
rect 2474 917 2475 921
rect 2479 917 2480 921
rect 2474 916 2480 917
rect 2626 921 2632 922
rect 2626 917 2627 921
rect 2631 917 2632 921
rect 2626 916 2632 917
rect 2802 921 2808 922
rect 2802 917 2803 921
rect 2807 917 2808 921
rect 2802 916 2808 917
rect 2994 921 3000 922
rect 2994 917 2995 921
rect 2999 917 3000 921
rect 2994 916 3000 917
rect 3202 921 3208 922
rect 3202 917 3203 921
rect 3207 917 3208 921
rect 3202 916 3208 917
rect 3426 921 3432 922
rect 3426 917 3427 921
rect 3431 917 3432 921
rect 3426 916 3432 917
rect 3650 921 3656 922
rect 3650 917 3651 921
rect 3655 917 3656 921
rect 3650 916 3656 917
rect 3798 920 3804 921
rect 3798 916 3799 920
rect 3803 916 3804 920
rect 1974 915 1980 916
rect 3798 915 3804 916
rect 110 884 116 885
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 194 883 200 884
rect 194 879 195 883
rect 199 879 200 883
rect 194 878 200 879
rect 370 883 376 884
rect 370 879 371 883
rect 375 879 376 883
rect 370 878 376 879
rect 546 883 552 884
rect 546 879 547 883
rect 551 879 552 883
rect 546 878 552 879
rect 722 883 728 884
rect 722 879 723 883
rect 727 879 728 883
rect 722 878 728 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1090 883 1096 884
rect 1090 879 1091 883
rect 1095 879 1096 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 3838 880 3844 881
rect 5662 880 5668 881
rect 1090 878 1096 879
rect 3838 876 3839 880
rect 3843 876 3844 880
rect 3838 875 3844 876
rect 4586 879 4592 880
rect 4586 875 4587 879
rect 4591 875 4592 879
rect 4586 874 4592 875
rect 4754 879 4760 880
rect 4754 875 4755 879
rect 4759 875 4760 879
rect 4754 874 4760 875
rect 4938 879 4944 880
rect 4938 875 4939 879
rect 4943 875 4944 879
rect 4938 874 4944 875
rect 5130 879 5136 880
rect 5130 875 5131 879
rect 5135 875 5136 879
rect 5130 874 5136 875
rect 5330 879 5336 880
rect 5330 875 5331 879
rect 5335 875 5336 879
rect 5330 874 5336 875
rect 5514 879 5520 880
rect 5514 875 5515 879
rect 5519 875 5520 879
rect 5662 876 5663 880
rect 5667 876 5668 880
rect 5662 875 5668 876
rect 5514 874 5520 875
rect 222 868 228 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 222 864 223 868
rect 227 864 228 868
rect 222 863 228 864
rect 398 868 404 869
rect 398 864 399 868
rect 403 864 404 868
rect 398 863 404 864
rect 574 868 580 869
rect 574 864 575 868
rect 579 864 580 868
rect 574 863 580 864
rect 750 868 756 869
rect 750 864 751 868
rect 755 864 756 868
rect 750 863 756 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1118 868 1124 869
rect 1118 864 1119 868
rect 1123 864 1124 868
rect 1118 863 1124 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 4614 864 4620 865
rect 110 862 116 863
rect 1934 862 1940 863
rect 3838 863 3844 864
rect 3838 859 3839 863
rect 3843 859 3844 863
rect 4614 860 4615 864
rect 4619 860 4620 864
rect 4614 859 4620 860
rect 4782 864 4788 865
rect 4782 860 4783 864
rect 4787 860 4788 864
rect 4782 859 4788 860
rect 4966 864 4972 865
rect 4966 860 4967 864
rect 4971 860 4972 864
rect 4966 859 4972 860
rect 5158 864 5164 865
rect 5158 860 5159 864
rect 5163 860 5164 864
rect 5158 859 5164 860
rect 5358 864 5364 865
rect 5358 860 5359 864
rect 5363 860 5364 864
rect 5358 859 5364 860
rect 5542 864 5548 865
rect 5542 860 5543 864
rect 5547 860 5548 864
rect 5542 859 5548 860
rect 5662 863 5668 864
rect 5662 859 5663 863
rect 5667 859 5668 863
rect 3838 858 3844 859
rect 5662 858 5668 859
rect 3838 797 3844 798
rect 5662 797 5668 798
rect 110 793 116 794
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 158 792 164 793
rect 158 788 159 792
rect 163 788 164 792
rect 158 787 164 788
rect 350 792 356 793
rect 350 788 351 792
rect 355 788 356 792
rect 350 787 356 788
rect 582 792 588 793
rect 582 788 583 792
rect 587 788 588 792
rect 582 787 588 788
rect 838 792 844 793
rect 838 788 839 792
rect 843 788 844 792
rect 838 787 844 788
rect 1110 792 1116 793
rect 1110 788 1111 792
rect 1115 788 1116 792
rect 1110 787 1116 788
rect 1398 792 1404 793
rect 1398 788 1399 792
rect 1403 788 1404 792
rect 1398 787 1404 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3982 796 3988 797
rect 3982 792 3983 796
rect 3987 792 3988 796
rect 3982 791 3988 792
rect 4238 796 4244 797
rect 4238 792 4239 796
rect 4243 792 4244 796
rect 4238 791 4244 792
rect 4534 796 4540 797
rect 4534 792 4535 796
rect 4539 792 4540 796
rect 4534 791 4540 792
rect 4862 796 4868 797
rect 4862 792 4863 796
rect 4867 792 4868 796
rect 4862 791 4868 792
rect 5214 796 5220 797
rect 5214 792 5215 796
rect 5219 792 5220 796
rect 5214 791 5220 792
rect 5542 796 5548 797
rect 5542 792 5543 796
rect 5547 792 5548 796
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5542 791 5548 792
rect 1934 788 1940 789
rect 1974 788 1980 789
rect 3798 788 3804 789
rect 1686 787 1692 788
rect 1974 784 1975 788
rect 1979 784 1980 788
rect 1974 783 1980 784
rect 2306 787 2312 788
rect 2306 783 2307 787
rect 2311 783 2312 787
rect 2306 782 2312 783
rect 2482 787 2488 788
rect 2482 783 2483 787
rect 2487 783 2488 787
rect 2482 782 2488 783
rect 2658 787 2664 788
rect 2658 783 2659 787
rect 2663 783 2664 787
rect 2658 782 2664 783
rect 2826 787 2832 788
rect 2826 783 2827 787
rect 2831 783 2832 787
rect 2826 782 2832 783
rect 2994 787 3000 788
rect 2994 783 2995 787
rect 2999 783 3000 787
rect 2994 782 3000 783
rect 3162 787 3168 788
rect 3162 783 3163 787
rect 3167 783 3168 787
rect 3162 782 3168 783
rect 3330 787 3336 788
rect 3330 783 3331 787
rect 3335 783 3336 787
rect 3330 782 3336 783
rect 3498 787 3504 788
rect 3498 783 3499 787
rect 3503 783 3504 787
rect 3498 782 3504 783
rect 3650 787 3656 788
rect 3650 783 3651 787
rect 3655 783 3656 787
rect 3798 784 3799 788
rect 3803 784 3804 788
rect 3798 783 3804 784
rect 3650 782 3656 783
rect 3954 781 3960 782
rect 3838 780 3844 781
rect 130 777 136 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 130 773 131 777
rect 135 773 136 777
rect 130 772 136 773
rect 322 777 328 778
rect 322 773 323 777
rect 327 773 328 777
rect 322 772 328 773
rect 554 777 560 778
rect 554 773 555 777
rect 559 773 560 777
rect 554 772 560 773
rect 810 777 816 778
rect 810 773 811 777
rect 815 773 816 777
rect 810 772 816 773
rect 1082 777 1088 778
rect 1082 773 1083 777
rect 1087 773 1088 777
rect 1082 772 1088 773
rect 1370 777 1376 778
rect 1370 773 1371 777
rect 1375 773 1376 777
rect 1370 772 1376 773
rect 1658 777 1664 778
rect 1658 773 1659 777
rect 1663 773 1664 777
rect 1658 772 1664 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3954 777 3955 781
rect 3959 777 3960 781
rect 3954 776 3960 777
rect 4210 781 4216 782
rect 4210 777 4211 781
rect 4215 777 4216 781
rect 4210 776 4216 777
rect 4506 781 4512 782
rect 4506 777 4507 781
rect 4511 777 4512 781
rect 4506 776 4512 777
rect 4834 781 4840 782
rect 4834 777 4835 781
rect 4839 777 4840 781
rect 4834 776 4840 777
rect 5186 781 5192 782
rect 5186 777 5187 781
rect 5191 777 5192 781
rect 5186 776 5192 777
rect 5514 781 5520 782
rect 5514 777 5515 781
rect 5519 777 5520 781
rect 5514 776 5520 777
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 3838 775 3844 776
rect 5662 775 5668 776
rect 2334 772 2340 773
rect 110 771 116 772
rect 1934 771 1940 772
rect 1974 771 1980 772
rect 1974 767 1975 771
rect 1979 767 1980 771
rect 2334 768 2335 772
rect 2339 768 2340 772
rect 2334 767 2340 768
rect 2510 772 2516 773
rect 2510 768 2511 772
rect 2515 768 2516 772
rect 2510 767 2516 768
rect 2686 772 2692 773
rect 2686 768 2687 772
rect 2691 768 2692 772
rect 2686 767 2692 768
rect 2854 772 2860 773
rect 2854 768 2855 772
rect 2859 768 2860 772
rect 2854 767 2860 768
rect 3022 772 3028 773
rect 3022 768 3023 772
rect 3027 768 3028 772
rect 3022 767 3028 768
rect 3190 772 3196 773
rect 3190 768 3191 772
rect 3195 768 3196 772
rect 3190 767 3196 768
rect 3358 772 3364 773
rect 3358 768 3359 772
rect 3363 768 3364 772
rect 3358 767 3364 768
rect 3526 772 3532 773
rect 3526 768 3527 772
rect 3531 768 3532 772
rect 3526 767 3532 768
rect 3678 772 3684 773
rect 3678 768 3679 772
rect 3683 768 3684 772
rect 3678 767 3684 768
rect 3798 771 3804 772
rect 3798 767 3799 771
rect 3803 767 3804 771
rect 1974 766 1980 767
rect 3798 766 3804 767
rect 1974 709 1980 710
rect 3798 709 3804 710
rect 1974 705 1975 709
rect 1979 705 1980 709
rect 1974 704 1980 705
rect 3134 708 3140 709
rect 3134 704 3135 708
rect 3139 704 3140 708
rect 3134 703 3140 704
rect 3270 708 3276 709
rect 3270 704 3271 708
rect 3275 704 3276 708
rect 3270 703 3276 704
rect 3406 708 3412 709
rect 3406 704 3407 708
rect 3411 704 3412 708
rect 3406 703 3412 704
rect 3542 708 3548 709
rect 3542 704 3543 708
rect 3547 704 3548 708
rect 3542 703 3548 704
rect 3678 708 3684 709
rect 3678 704 3679 708
rect 3683 704 3684 708
rect 3798 705 3799 709
rect 3803 705 3804 709
rect 3798 704 3804 705
rect 3678 703 3684 704
rect 3106 693 3112 694
rect 1974 692 1980 693
rect 1974 688 1975 692
rect 1979 688 1980 692
rect 3106 689 3107 693
rect 3111 689 3112 693
rect 3106 688 3112 689
rect 3242 693 3248 694
rect 3242 689 3243 693
rect 3247 689 3248 693
rect 3242 688 3248 689
rect 3378 693 3384 694
rect 3378 689 3379 693
rect 3383 689 3384 693
rect 3378 688 3384 689
rect 3514 693 3520 694
rect 3514 689 3515 693
rect 3519 689 3520 693
rect 3514 688 3520 689
rect 3650 693 3656 694
rect 3650 689 3651 693
rect 3655 689 3656 693
rect 3650 688 3656 689
rect 3798 692 3804 693
rect 3798 688 3799 692
rect 3803 688 3804 692
rect 1974 687 1980 688
rect 3798 687 3804 688
rect 110 644 116 645
rect 1934 644 1940 645
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 290 643 296 644
rect 290 639 291 643
rect 295 639 296 643
rect 290 638 296 639
rect 482 643 488 644
rect 482 639 483 643
rect 487 639 488 643
rect 482 638 488 639
rect 674 643 680 644
rect 674 639 675 643
rect 679 639 680 643
rect 674 638 680 639
rect 866 643 872 644
rect 866 639 867 643
rect 871 639 872 643
rect 866 638 872 639
rect 1058 643 1064 644
rect 1058 639 1059 643
rect 1063 639 1064 643
rect 1058 638 1064 639
rect 1250 643 1256 644
rect 1250 639 1251 643
rect 1255 639 1256 643
rect 1250 638 1256 639
rect 1434 643 1440 644
rect 1434 639 1435 643
rect 1439 639 1440 643
rect 1434 638 1440 639
rect 1618 643 1624 644
rect 1618 639 1619 643
rect 1623 639 1624 643
rect 1618 638 1624 639
rect 1786 643 1792 644
rect 1786 639 1787 643
rect 1791 639 1792 643
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 1786 638 1792 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 318 628 324 629
rect 318 624 319 628
rect 323 624 324 628
rect 318 623 324 624
rect 510 628 516 629
rect 510 624 511 628
rect 515 624 516 628
rect 510 623 516 624
rect 702 628 708 629
rect 702 624 703 628
rect 707 624 708 628
rect 702 623 708 624
rect 894 628 900 629
rect 894 624 895 628
rect 899 624 900 628
rect 894 623 900 624
rect 1086 628 1092 629
rect 1086 624 1087 628
rect 1091 624 1092 628
rect 1086 623 1092 624
rect 1278 628 1284 629
rect 1278 624 1279 628
rect 1283 624 1284 628
rect 1278 623 1284 624
rect 1462 628 1468 629
rect 1462 624 1463 628
rect 1467 624 1468 628
rect 1462 623 1468 624
rect 1646 628 1652 629
rect 1646 624 1647 628
rect 1651 624 1652 628
rect 1646 623 1652 624
rect 1814 628 1820 629
rect 1814 624 1815 628
rect 1819 624 1820 628
rect 1814 623 1820 624
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 110 622 116 623
rect 1934 622 1940 623
rect 3838 624 3844 625
rect 5662 624 5668 625
rect 3838 620 3839 624
rect 3843 620 3844 624
rect 3838 619 3844 620
rect 3858 623 3864 624
rect 3858 619 3859 623
rect 3863 619 3864 623
rect 3858 618 3864 619
rect 3994 623 4000 624
rect 3994 619 3995 623
rect 3999 619 4000 623
rect 3994 618 4000 619
rect 4138 623 4144 624
rect 4138 619 4139 623
rect 4143 619 4144 623
rect 4138 618 4144 619
rect 4322 623 4328 624
rect 4322 619 4323 623
rect 4327 619 4328 623
rect 4322 618 4328 619
rect 4530 623 4536 624
rect 4530 619 4531 623
rect 4535 619 4536 623
rect 4530 618 4536 619
rect 4754 623 4760 624
rect 4754 619 4755 623
rect 4759 619 4760 623
rect 4754 618 4760 619
rect 4994 623 5000 624
rect 4994 619 4995 623
rect 4999 619 5000 623
rect 4994 618 5000 619
rect 5242 623 5248 624
rect 5242 619 5243 623
rect 5247 619 5248 623
rect 5242 618 5248 619
rect 5498 623 5504 624
rect 5498 619 5499 623
rect 5503 619 5504 623
rect 5662 620 5663 624
rect 5667 620 5668 624
rect 5662 619 5668 620
rect 5498 618 5504 619
rect 3886 608 3892 609
rect 3838 607 3844 608
rect 3838 603 3839 607
rect 3843 603 3844 607
rect 3886 604 3887 608
rect 3891 604 3892 608
rect 3886 603 3892 604
rect 4022 608 4028 609
rect 4022 604 4023 608
rect 4027 604 4028 608
rect 4022 603 4028 604
rect 4166 608 4172 609
rect 4166 604 4167 608
rect 4171 604 4172 608
rect 4166 603 4172 604
rect 4350 608 4356 609
rect 4350 604 4351 608
rect 4355 604 4356 608
rect 4350 603 4356 604
rect 4558 608 4564 609
rect 4558 604 4559 608
rect 4563 604 4564 608
rect 4558 603 4564 604
rect 4782 608 4788 609
rect 4782 604 4783 608
rect 4787 604 4788 608
rect 4782 603 4788 604
rect 5022 608 5028 609
rect 5022 604 5023 608
rect 5027 604 5028 608
rect 5022 603 5028 604
rect 5270 608 5276 609
rect 5270 604 5271 608
rect 5275 604 5276 608
rect 5270 603 5276 604
rect 5526 608 5532 609
rect 5526 604 5527 608
rect 5531 604 5532 608
rect 5526 603 5532 604
rect 5662 607 5668 608
rect 5662 603 5663 607
rect 5667 603 5668 607
rect 3838 602 3844 603
rect 5662 602 5668 603
rect 110 569 116 570
rect 1934 569 1940 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 326 568 332 569
rect 326 564 327 568
rect 331 564 332 568
rect 326 563 332 564
rect 518 568 524 569
rect 518 564 519 568
rect 523 564 524 568
rect 518 563 524 564
rect 710 568 716 569
rect 710 564 711 568
rect 715 564 716 568
rect 710 563 716 564
rect 902 568 908 569
rect 902 564 903 568
rect 907 564 908 568
rect 902 563 908 564
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 1094 563 1100 564
rect 1278 568 1284 569
rect 1278 564 1279 568
rect 1283 564 1284 568
rect 1278 563 1284 564
rect 1462 568 1468 569
rect 1462 564 1463 568
rect 1467 564 1468 568
rect 1462 563 1468 564
rect 1646 568 1652 569
rect 1646 564 1647 568
rect 1651 564 1652 568
rect 1646 563 1652 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 1814 563 1820 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 298 553 304 554
rect 298 549 299 553
rect 303 549 304 553
rect 298 548 304 549
rect 490 553 496 554
rect 490 549 491 553
rect 495 549 496 553
rect 490 548 496 549
rect 682 553 688 554
rect 682 549 683 553
rect 687 549 688 553
rect 682 548 688 549
rect 874 553 880 554
rect 874 549 875 553
rect 879 549 880 553
rect 874 548 880 549
rect 1066 553 1072 554
rect 1066 549 1067 553
rect 1071 549 1072 553
rect 1066 548 1072 549
rect 1250 553 1256 554
rect 1250 549 1251 553
rect 1255 549 1256 553
rect 1250 548 1256 549
rect 1434 553 1440 554
rect 1434 549 1435 553
rect 1439 549 1440 553
rect 1434 548 1440 549
rect 1618 553 1624 554
rect 1618 549 1619 553
rect 1623 549 1624 553
rect 1618 548 1624 549
rect 1786 553 1792 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 110 547 116 548
rect 1934 547 1940 548
rect 3838 549 3844 550
rect 5662 549 5668 550
rect 3838 545 3839 549
rect 3843 545 3844 549
rect 3838 544 3844 545
rect 3886 548 3892 549
rect 3886 544 3887 548
rect 3891 544 3892 548
rect 3886 543 3892 544
rect 4022 548 4028 549
rect 4022 544 4023 548
rect 4027 544 4028 548
rect 4022 543 4028 544
rect 4158 548 4164 549
rect 4158 544 4159 548
rect 4163 544 4164 548
rect 4158 543 4164 544
rect 4294 548 4300 549
rect 4294 544 4295 548
rect 4299 544 4300 548
rect 4294 543 4300 544
rect 4430 548 4436 549
rect 4430 544 4431 548
rect 4435 544 4436 548
rect 4430 543 4436 544
rect 4574 548 4580 549
rect 4574 544 4575 548
rect 4579 544 4580 548
rect 4574 543 4580 544
rect 4742 548 4748 549
rect 4742 544 4743 548
rect 4747 544 4748 548
rect 4742 543 4748 544
rect 4926 548 4932 549
rect 4926 544 4927 548
rect 4931 544 4932 548
rect 4926 543 4932 544
rect 5118 548 5124 549
rect 5118 544 5119 548
rect 5123 544 5124 548
rect 5118 543 5124 544
rect 5318 548 5324 549
rect 5318 544 5319 548
rect 5323 544 5324 548
rect 5318 543 5324 544
rect 5526 548 5532 549
rect 5526 544 5527 548
rect 5531 544 5532 548
rect 5662 545 5663 549
rect 5667 545 5668 549
rect 5662 544 5668 545
rect 5526 543 5532 544
rect 3858 533 3864 534
rect 3838 532 3844 533
rect 3838 528 3839 532
rect 3843 528 3844 532
rect 3858 529 3859 533
rect 3863 529 3864 533
rect 3858 528 3864 529
rect 3994 533 4000 534
rect 3994 529 3995 533
rect 3999 529 4000 533
rect 3994 528 4000 529
rect 4130 533 4136 534
rect 4130 529 4131 533
rect 4135 529 4136 533
rect 4130 528 4136 529
rect 4266 533 4272 534
rect 4266 529 4267 533
rect 4271 529 4272 533
rect 4266 528 4272 529
rect 4402 533 4408 534
rect 4402 529 4403 533
rect 4407 529 4408 533
rect 4402 528 4408 529
rect 4546 533 4552 534
rect 4546 529 4547 533
rect 4551 529 4552 533
rect 4546 528 4552 529
rect 4714 533 4720 534
rect 4714 529 4715 533
rect 4719 529 4720 533
rect 4714 528 4720 529
rect 4898 533 4904 534
rect 4898 529 4899 533
rect 4903 529 4904 533
rect 4898 528 4904 529
rect 5090 533 5096 534
rect 5090 529 5091 533
rect 5095 529 5096 533
rect 5090 528 5096 529
rect 5290 533 5296 534
rect 5290 529 5291 533
rect 5295 529 5296 533
rect 5290 528 5296 529
rect 5498 533 5504 534
rect 5498 529 5499 533
rect 5503 529 5504 533
rect 5498 528 5504 529
rect 5662 532 5668 533
rect 5662 528 5663 532
rect 5667 528 5668 532
rect 3838 527 3844 528
rect 5662 527 5668 528
rect 110 420 116 421
rect 1934 420 1940 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 394 419 400 420
rect 394 415 395 419
rect 399 415 400 419
rect 394 414 400 415
rect 586 419 592 420
rect 586 415 587 419
rect 591 415 592 419
rect 586 414 592 415
rect 786 419 792 420
rect 786 415 787 419
rect 791 415 792 419
rect 786 414 792 415
rect 986 419 992 420
rect 986 415 987 419
rect 991 415 992 419
rect 986 414 992 415
rect 1194 419 1200 420
rect 1194 415 1195 419
rect 1199 415 1200 419
rect 1194 414 1200 415
rect 1410 419 1416 420
rect 1410 415 1411 419
rect 1415 415 1416 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 1410 414 1416 415
rect 422 404 428 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 422 400 423 404
rect 427 400 428 404
rect 422 399 428 400
rect 614 404 620 405
rect 614 400 615 404
rect 619 400 620 404
rect 614 399 620 400
rect 814 404 820 405
rect 814 400 815 404
rect 819 400 820 404
rect 814 399 820 400
rect 1014 404 1020 405
rect 1014 400 1015 404
rect 1019 400 1020 404
rect 1014 399 1020 400
rect 1222 404 1228 405
rect 1222 400 1223 404
rect 1227 400 1228 404
rect 1222 399 1228 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1934 403 1940 404
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 110 398 116 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 3798 400 3804 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2866 399 2872 400
rect 2866 395 2867 399
rect 2871 395 2872 399
rect 2866 394 2872 395
rect 3074 399 3080 400
rect 3074 395 3075 399
rect 3079 395 3080 399
rect 3074 394 3080 395
rect 3274 399 3280 400
rect 3274 395 3275 399
rect 3279 395 3280 399
rect 3274 394 3280 395
rect 3474 399 3480 400
rect 3474 395 3475 399
rect 3479 395 3480 399
rect 3474 394 3480 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3838 400 3844 401
rect 5662 400 5668 401
rect 3838 396 3839 400
rect 3843 396 3844 400
rect 3838 395 3844 396
rect 4378 399 4384 400
rect 4378 395 4379 399
rect 4383 395 4384 399
rect 3650 394 3656 395
rect 4378 394 4384 395
rect 4594 399 4600 400
rect 4594 395 4595 399
rect 4599 395 4600 399
rect 4594 394 4600 395
rect 4818 399 4824 400
rect 4818 395 4819 399
rect 4823 395 4824 399
rect 4818 394 4824 395
rect 5050 399 5056 400
rect 5050 395 5051 399
rect 5055 395 5056 399
rect 5050 394 5056 395
rect 5282 399 5288 400
rect 5282 395 5283 399
rect 5287 395 5288 399
rect 5662 396 5663 400
rect 5667 396 5668 400
rect 5662 395 5668 396
rect 5282 394 5288 395
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 2894 384 2900 385
rect 2894 380 2895 384
rect 2899 380 2900 384
rect 2894 379 2900 380
rect 3102 384 3108 385
rect 3102 380 3103 384
rect 3107 380 3108 384
rect 3102 379 3108 380
rect 3302 384 3308 385
rect 3302 380 3303 384
rect 3307 380 3308 384
rect 3302 379 3308 380
rect 3502 384 3508 385
rect 3502 380 3503 384
rect 3507 380 3508 384
rect 3502 379 3508 380
rect 3678 384 3684 385
rect 4406 384 4412 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 3798 378 3804 379
rect 3838 383 3844 384
rect 3838 379 3839 383
rect 3843 379 3844 383
rect 4406 380 4407 384
rect 4411 380 4412 384
rect 4406 379 4412 380
rect 4622 384 4628 385
rect 4622 380 4623 384
rect 4627 380 4628 384
rect 4622 379 4628 380
rect 4846 384 4852 385
rect 4846 380 4847 384
rect 4851 380 4852 384
rect 4846 379 4852 380
rect 5078 384 5084 385
rect 5078 380 5079 384
rect 5083 380 5084 384
rect 5078 379 5084 380
rect 5310 384 5316 385
rect 5310 380 5311 384
rect 5315 380 5316 384
rect 5310 379 5316 380
rect 5662 383 5668 384
rect 5662 379 5663 383
rect 5667 379 5668 383
rect 3838 378 3844 379
rect 5662 378 5668 379
rect 110 333 116 334
rect 1934 333 1940 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 646 332 652 333
rect 646 328 647 332
rect 651 328 652 332
rect 646 327 652 328
rect 814 332 820 333
rect 814 328 815 332
rect 819 328 820 332
rect 814 327 820 328
rect 990 332 996 333
rect 990 328 991 332
rect 995 328 996 332
rect 990 327 996 328
rect 1166 332 1172 333
rect 1166 328 1167 332
rect 1171 328 1172 332
rect 1166 327 1172 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 1342 327 1348 328
rect 3838 325 3844 326
rect 5662 325 5668 326
rect 3838 321 3839 325
rect 3843 321 3844 325
rect 3838 320 3844 321
rect 4638 324 4644 325
rect 4638 320 4639 324
rect 4643 320 4644 324
rect 4638 319 4644 320
rect 4806 324 4812 325
rect 4806 320 4807 324
rect 4811 320 4812 324
rect 4806 319 4812 320
rect 4982 324 4988 325
rect 4982 320 4983 324
rect 4987 320 4988 324
rect 4982 319 4988 320
rect 5166 324 5172 325
rect 5166 320 5167 324
rect 5171 320 5172 324
rect 5166 319 5172 320
rect 5358 324 5364 325
rect 5358 320 5359 324
rect 5363 320 5364 324
rect 5358 319 5364 320
rect 5542 324 5548 325
rect 5542 320 5543 324
rect 5547 320 5548 324
rect 5662 321 5663 325
rect 5667 321 5668 325
rect 5662 320 5668 321
rect 5542 319 5548 320
rect 618 317 624 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 618 313 619 317
rect 623 313 624 317
rect 618 312 624 313
rect 786 317 792 318
rect 786 313 787 317
rect 791 313 792 317
rect 786 312 792 313
rect 962 317 968 318
rect 962 313 963 317
rect 967 313 968 317
rect 962 312 968 313
rect 1138 317 1144 318
rect 1138 313 1139 317
rect 1143 313 1144 317
rect 1138 312 1144 313
rect 1314 317 1320 318
rect 1314 313 1315 317
rect 1319 313 1320 317
rect 1314 312 1320 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 110 311 116 312
rect 1934 311 1940 312
rect 1974 309 1980 310
rect 3798 309 3804 310
rect 4610 309 4616 310
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3798 304 3804 305
rect 3838 308 3844 309
rect 3838 304 3839 308
rect 3843 304 3844 308
rect 4610 305 4611 309
rect 4615 305 4616 309
rect 4610 304 4616 305
rect 4778 309 4784 310
rect 4778 305 4779 309
rect 4783 305 4784 309
rect 4778 304 4784 305
rect 4954 309 4960 310
rect 4954 305 4955 309
rect 4959 305 4960 309
rect 4954 304 4960 305
rect 5138 309 5144 310
rect 5138 305 5139 309
rect 5143 305 5144 309
rect 5138 304 5144 305
rect 5330 309 5336 310
rect 5330 305 5331 309
rect 5335 305 5336 309
rect 5330 304 5336 305
rect 5514 309 5520 310
rect 5514 305 5515 309
rect 5519 305 5520 309
rect 5514 304 5520 305
rect 5662 308 5668 309
rect 5662 304 5663 308
rect 5667 304 5668 308
rect 3654 303 3660 304
rect 3838 303 3844 304
rect 5662 303 5668 304
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 1974 287 1980 288
rect 3798 287 3804 288
rect 3838 148 3844 149
rect 5662 148 5668 149
rect 110 144 116 145
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1082 138 1088 139
rect 1218 143 1224 144
rect 1218 139 1219 143
rect 1223 139 1224 143
rect 1218 138 1224 139
rect 1354 143 1360 144
rect 1354 139 1355 143
rect 1359 139 1360 143
rect 1354 138 1360 139
rect 1490 143 1496 144
rect 1490 139 1491 143
rect 1495 139 1496 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 3838 144 3839 148
rect 3843 144 3844 148
rect 3838 143 3844 144
rect 4290 147 4296 148
rect 4290 143 4291 147
rect 4295 143 4296 147
rect 4290 142 4296 143
rect 4426 147 4432 148
rect 4426 143 4427 147
rect 4431 143 4432 147
rect 4426 142 4432 143
rect 4562 147 4568 148
rect 4562 143 4563 147
rect 4567 143 4568 147
rect 4562 142 4568 143
rect 4698 147 4704 148
rect 4698 143 4699 147
rect 4703 143 4704 147
rect 4698 142 4704 143
rect 4834 147 4840 148
rect 4834 143 4835 147
rect 4839 143 4840 147
rect 4834 142 4840 143
rect 4970 147 4976 148
rect 4970 143 4971 147
rect 4975 143 4976 147
rect 4970 142 4976 143
rect 5106 147 5112 148
rect 5106 143 5107 147
rect 5111 143 5112 147
rect 5106 142 5112 143
rect 5242 147 5248 148
rect 5242 143 5243 147
rect 5247 143 5248 147
rect 5242 142 5248 143
rect 5378 147 5384 148
rect 5378 143 5379 147
rect 5383 143 5384 147
rect 5378 142 5384 143
rect 5514 147 5520 148
rect 5514 143 5515 147
rect 5519 143 5520 147
rect 5662 144 5663 148
rect 5667 144 5668 148
rect 5662 143 5668 144
rect 5514 142 5520 143
rect 1934 139 1940 140
rect 1490 138 1496 139
rect 4318 132 4324 133
rect 3838 131 3844 132
rect 566 128 572 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1246 128 1252 129
rect 1246 124 1247 128
rect 1251 124 1252 128
rect 1246 123 1252 124
rect 1382 128 1388 129
rect 1382 124 1383 128
rect 1387 124 1388 128
rect 1382 123 1388 124
rect 1518 128 1524 129
rect 1518 124 1519 128
rect 1523 124 1524 128
rect 1518 123 1524 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 3838 127 3839 131
rect 3843 127 3844 131
rect 4318 128 4319 132
rect 4323 128 4324 132
rect 4318 127 4324 128
rect 4454 132 4460 133
rect 4454 128 4455 132
rect 4459 128 4460 132
rect 4454 127 4460 128
rect 4590 132 4596 133
rect 4590 128 4591 132
rect 4595 128 4596 132
rect 4590 127 4596 128
rect 4726 132 4732 133
rect 4726 128 4727 132
rect 4731 128 4732 132
rect 4726 127 4732 128
rect 4862 132 4868 133
rect 4862 128 4863 132
rect 4867 128 4868 132
rect 4862 127 4868 128
rect 4998 132 5004 133
rect 4998 128 4999 132
rect 5003 128 5004 132
rect 4998 127 5004 128
rect 5134 132 5140 133
rect 5134 128 5135 132
rect 5139 128 5140 132
rect 5134 127 5140 128
rect 5270 132 5276 133
rect 5270 128 5271 132
rect 5275 128 5276 132
rect 5270 127 5276 128
rect 5406 132 5412 133
rect 5406 128 5407 132
rect 5411 128 5412 132
rect 5406 127 5412 128
rect 5542 132 5548 133
rect 5542 128 5543 132
rect 5547 128 5548 132
rect 5542 127 5548 128
rect 5662 131 5668 132
rect 5662 127 5663 131
rect 5667 127 5668 131
rect 3838 126 3844 127
rect 5662 126 5668 127
rect 110 122 116 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 3798 124 3804 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3626 118 3632 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 3798 102 3804 103
<< m3c >>
rect 111 5689 115 5693
rect 159 5688 163 5692
rect 303 5688 307 5692
rect 503 5688 507 5692
rect 727 5688 731 5692
rect 983 5688 987 5692
rect 1255 5688 1259 5692
rect 1543 5688 1547 5692
rect 1815 5688 1819 5692
rect 1935 5689 1939 5693
rect 111 5672 115 5676
rect 131 5673 135 5677
rect 275 5673 279 5677
rect 475 5673 479 5677
rect 699 5673 703 5677
rect 955 5673 959 5677
rect 1227 5673 1231 5677
rect 1515 5673 1519 5677
rect 1787 5673 1791 5677
rect 1935 5672 1939 5676
rect 1975 5624 1979 5628
rect 1995 5623 1999 5627
rect 2179 5623 2183 5627
rect 2387 5623 2391 5627
rect 2587 5623 2591 5627
rect 2779 5623 2783 5627
rect 2963 5623 2967 5627
rect 3147 5623 3151 5627
rect 3323 5623 3327 5627
rect 3499 5623 3503 5627
rect 3651 5623 3655 5627
rect 3799 5624 3803 5628
rect 1975 5607 1979 5611
rect 2023 5608 2027 5612
rect 2207 5608 2211 5612
rect 2415 5608 2419 5612
rect 2615 5608 2619 5612
rect 2807 5608 2811 5612
rect 2991 5608 2995 5612
rect 3175 5608 3179 5612
rect 3351 5608 3355 5612
rect 3527 5608 3531 5612
rect 3679 5608 3683 5612
rect 3799 5607 3803 5611
rect 3839 5580 3843 5584
rect 4291 5579 4295 5583
rect 4427 5579 4431 5583
rect 4563 5579 4567 5583
rect 4699 5579 4703 5583
rect 4835 5579 4839 5583
rect 4971 5579 4975 5583
rect 5107 5579 5111 5583
rect 5663 5580 5667 5584
rect 3839 5563 3843 5567
rect 4319 5564 4323 5568
rect 4455 5564 4459 5568
rect 4591 5564 4595 5568
rect 4727 5564 4731 5568
rect 4863 5564 4867 5568
rect 4999 5564 5003 5568
rect 5135 5564 5139 5568
rect 5663 5563 5667 5567
rect 1975 5549 1979 5553
rect 2263 5548 2267 5552
rect 2503 5548 2507 5552
rect 2743 5548 2747 5552
rect 2983 5548 2987 5552
rect 3223 5548 3227 5552
rect 3463 5548 3467 5552
rect 3679 5548 3683 5552
rect 3799 5549 3803 5553
rect 111 5536 115 5540
rect 563 5535 567 5539
rect 723 5535 727 5539
rect 883 5535 887 5539
rect 1051 5535 1055 5539
rect 1227 5535 1231 5539
rect 1403 5535 1407 5539
rect 1579 5535 1583 5539
rect 1763 5535 1767 5539
rect 1935 5536 1939 5540
rect 1975 5532 1979 5536
rect 2235 5533 2239 5537
rect 2475 5533 2479 5537
rect 2715 5533 2719 5537
rect 2955 5533 2959 5537
rect 3195 5533 3199 5537
rect 3435 5533 3439 5537
rect 3651 5533 3655 5537
rect 3799 5532 3803 5536
rect 111 5519 115 5523
rect 591 5520 595 5524
rect 751 5520 755 5524
rect 911 5520 915 5524
rect 1079 5520 1083 5524
rect 1255 5520 1259 5524
rect 1431 5520 1435 5524
rect 1607 5520 1611 5524
rect 1791 5520 1795 5524
rect 1935 5519 1939 5523
rect 3839 5505 3843 5509
rect 3887 5504 3891 5508
rect 4127 5504 4131 5508
rect 4375 5504 4379 5508
rect 4615 5504 4619 5508
rect 4847 5504 4851 5508
rect 5079 5504 5083 5508
rect 5311 5504 5315 5508
rect 5663 5505 5667 5509
rect 3839 5488 3843 5492
rect 3859 5489 3863 5493
rect 4099 5489 4103 5493
rect 4347 5489 4351 5493
rect 4587 5489 4591 5493
rect 4819 5489 4823 5493
rect 5051 5489 5055 5493
rect 5283 5489 5287 5493
rect 5663 5488 5667 5492
rect 111 5449 115 5453
rect 591 5448 595 5452
rect 727 5448 731 5452
rect 863 5448 867 5452
rect 999 5448 1003 5452
rect 1135 5448 1139 5452
rect 1271 5448 1275 5452
rect 1407 5448 1411 5452
rect 1543 5448 1547 5452
rect 1679 5448 1683 5452
rect 1815 5448 1819 5452
rect 1935 5449 1939 5453
rect 111 5432 115 5436
rect 563 5433 567 5437
rect 699 5433 703 5437
rect 835 5433 839 5437
rect 971 5433 975 5437
rect 1107 5433 1111 5437
rect 1243 5433 1247 5437
rect 1379 5433 1383 5437
rect 1515 5433 1519 5437
rect 1651 5433 1655 5437
rect 1787 5433 1791 5437
rect 1935 5432 1939 5436
rect 1975 5392 1979 5396
rect 2427 5391 2431 5395
rect 2643 5391 2647 5395
rect 2859 5391 2863 5395
rect 3075 5391 3079 5395
rect 3291 5391 3295 5395
rect 3799 5392 3803 5396
rect 1975 5375 1979 5379
rect 2455 5376 2459 5380
rect 2671 5376 2675 5380
rect 2887 5376 2891 5380
rect 3103 5376 3107 5380
rect 3319 5376 3323 5380
rect 3799 5375 3803 5379
rect 3839 5352 3843 5356
rect 3859 5351 3863 5355
rect 4075 5351 4079 5355
rect 4307 5351 4311 5355
rect 4531 5351 4535 5355
rect 4739 5351 4743 5355
rect 4939 5351 4943 5355
rect 5139 5351 5143 5355
rect 5339 5351 5343 5355
rect 5515 5351 5519 5355
rect 5663 5352 5667 5356
rect 3839 5335 3843 5339
rect 3887 5336 3891 5340
rect 4103 5336 4107 5340
rect 4335 5336 4339 5340
rect 4559 5336 4563 5340
rect 4767 5336 4771 5340
rect 4967 5336 4971 5340
rect 5167 5336 5171 5340
rect 5367 5336 5371 5340
rect 5543 5336 5547 5340
rect 5663 5335 5667 5339
rect 1975 5317 1979 5321
rect 2447 5316 2451 5320
rect 2583 5316 2587 5320
rect 2719 5316 2723 5320
rect 2855 5316 2859 5320
rect 2991 5316 2995 5320
rect 3135 5316 3139 5320
rect 3287 5316 3291 5320
rect 3799 5317 3803 5321
rect 1975 5300 1979 5304
rect 2419 5301 2423 5305
rect 2555 5301 2559 5305
rect 2691 5301 2695 5305
rect 2827 5301 2831 5305
rect 2963 5301 2967 5305
rect 3107 5301 3111 5305
rect 3259 5301 3263 5305
rect 3799 5300 3803 5304
rect 3839 5261 3843 5265
rect 3887 5260 3891 5264
rect 4095 5260 4099 5264
rect 4343 5260 4347 5264
rect 4615 5260 4619 5264
rect 4911 5260 4915 5264
rect 5215 5260 5219 5264
rect 5527 5260 5531 5264
rect 5663 5261 5667 5265
rect 3839 5244 3843 5248
rect 3859 5245 3863 5249
rect 4067 5245 4071 5249
rect 4315 5245 4319 5249
rect 4587 5245 4591 5249
rect 4883 5245 4887 5249
rect 5187 5245 5191 5249
rect 5499 5245 5503 5249
rect 5663 5244 5667 5248
rect 111 5196 115 5200
rect 459 5195 463 5199
rect 595 5195 599 5199
rect 731 5195 735 5199
rect 867 5195 871 5199
rect 1003 5195 1007 5199
rect 1139 5195 1143 5199
rect 1275 5195 1279 5199
rect 1411 5195 1415 5199
rect 1547 5195 1551 5199
rect 1935 5196 1939 5200
rect 111 5179 115 5183
rect 487 5180 491 5184
rect 623 5180 627 5184
rect 759 5180 763 5184
rect 895 5180 899 5184
rect 1031 5180 1035 5184
rect 1167 5180 1171 5184
rect 1303 5180 1307 5184
rect 1439 5180 1443 5184
rect 1575 5180 1579 5184
rect 1935 5179 1939 5183
rect 1975 5168 1979 5172
rect 2099 5167 2103 5171
rect 2235 5167 2239 5171
rect 2379 5167 2383 5171
rect 2531 5167 2535 5171
rect 2699 5167 2703 5171
rect 2883 5167 2887 5171
rect 3067 5167 3071 5171
rect 3259 5167 3263 5171
rect 3799 5168 3803 5172
rect 1975 5151 1979 5155
rect 2127 5152 2131 5156
rect 2263 5152 2267 5156
rect 2407 5152 2411 5156
rect 2559 5152 2563 5156
rect 2727 5152 2731 5156
rect 2911 5152 2915 5156
rect 3095 5152 3099 5156
rect 3287 5152 3291 5156
rect 3799 5151 3803 5155
rect 111 5105 115 5109
rect 319 5104 323 5108
rect 503 5104 507 5108
rect 703 5104 707 5108
rect 919 5104 923 5108
rect 1151 5104 1155 5108
rect 1391 5104 1395 5108
rect 1631 5104 1635 5108
rect 1935 5105 1939 5109
rect 3839 5104 3843 5108
rect 3859 5103 3863 5107
rect 3995 5103 3999 5107
rect 4155 5103 4159 5107
rect 4363 5103 4367 5107
rect 4611 5103 4615 5107
rect 4883 5103 4887 5107
rect 5171 5103 5175 5107
rect 5467 5103 5471 5107
rect 5663 5104 5667 5108
rect 111 5088 115 5092
rect 291 5089 295 5093
rect 475 5089 479 5093
rect 675 5089 679 5093
rect 891 5089 895 5093
rect 1123 5089 1127 5093
rect 1363 5089 1367 5093
rect 1603 5089 1607 5093
rect 1935 5088 1939 5092
rect 3839 5087 3843 5091
rect 3887 5088 3891 5092
rect 4023 5088 4027 5092
rect 4183 5088 4187 5092
rect 4391 5088 4395 5092
rect 4639 5088 4643 5092
rect 4911 5088 4915 5092
rect 5199 5088 5203 5092
rect 5495 5088 5499 5092
rect 5663 5087 5667 5091
rect 1975 5069 1979 5073
rect 2079 5068 2083 5072
rect 2359 5068 2363 5072
rect 2639 5068 2643 5072
rect 2911 5068 2915 5072
rect 3175 5068 3179 5072
rect 3439 5068 3443 5072
rect 3679 5068 3683 5072
rect 3799 5069 3803 5073
rect 1975 5052 1979 5056
rect 2051 5053 2055 5057
rect 2331 5053 2335 5057
rect 2611 5053 2615 5057
rect 2883 5053 2887 5057
rect 3147 5053 3151 5057
rect 3411 5053 3415 5057
rect 3651 5053 3655 5057
rect 3799 5052 3803 5056
rect 3839 5013 3843 5017
rect 4447 5012 4451 5016
rect 4631 5012 4635 5016
rect 4831 5012 4835 5016
rect 5047 5012 5051 5016
rect 5279 5012 5283 5016
rect 5511 5012 5515 5016
rect 5663 5013 5667 5017
rect 3839 4996 3843 5000
rect 4419 4997 4423 5001
rect 4603 4997 4607 5001
rect 4803 4997 4807 5001
rect 5019 4997 5023 5001
rect 5251 4997 5255 5001
rect 5483 4997 5487 5001
rect 5663 4996 5667 5000
rect 111 4956 115 4960
rect 139 4955 143 4959
rect 411 4955 415 4959
rect 683 4955 687 4959
rect 963 4955 967 4959
rect 1243 4955 1247 4959
rect 1523 4955 1527 4959
rect 1787 4955 1791 4959
rect 1935 4956 1939 4960
rect 111 4939 115 4943
rect 167 4940 171 4944
rect 439 4940 443 4944
rect 711 4940 715 4944
rect 991 4940 995 4944
rect 1271 4940 1275 4944
rect 1551 4940 1555 4944
rect 1815 4940 1819 4944
rect 1935 4939 1939 4943
rect 1975 4900 1979 4904
rect 1995 4899 1999 4903
rect 2131 4899 2135 4903
rect 2299 4899 2303 4903
rect 2467 4899 2471 4903
rect 2643 4899 2647 4903
rect 2819 4899 2823 4903
rect 2987 4899 2991 4903
rect 3155 4899 3159 4903
rect 3323 4899 3327 4903
rect 3499 4899 3503 4903
rect 3651 4899 3655 4903
rect 3799 4900 3803 4904
rect 111 4881 115 4885
rect 159 4880 163 4884
rect 415 4880 419 4884
rect 735 4880 739 4884
rect 1087 4880 1091 4884
rect 1463 4880 1467 4884
rect 1815 4880 1819 4884
rect 1935 4881 1939 4885
rect 1975 4883 1979 4887
rect 2023 4884 2027 4888
rect 2159 4884 2163 4888
rect 2327 4884 2331 4888
rect 2495 4884 2499 4888
rect 2671 4884 2675 4888
rect 2847 4884 2851 4888
rect 3015 4884 3019 4888
rect 3183 4884 3187 4888
rect 3351 4884 3355 4888
rect 3527 4884 3531 4888
rect 3679 4884 3683 4888
rect 3799 4883 3803 4887
rect 111 4864 115 4868
rect 131 4865 135 4869
rect 387 4865 391 4869
rect 707 4865 711 4869
rect 1059 4865 1063 4869
rect 1435 4865 1439 4869
rect 1787 4865 1791 4869
rect 1935 4864 1939 4868
rect 3839 4848 3843 4852
rect 4675 4847 4679 4851
rect 4827 4847 4831 4851
rect 4987 4847 4991 4851
rect 5155 4847 5159 4851
rect 5323 4847 5327 4851
rect 5499 4847 5503 4851
rect 5663 4848 5667 4852
rect 3839 4831 3843 4835
rect 4703 4832 4707 4836
rect 4855 4832 4859 4836
rect 5015 4832 5019 4836
rect 5183 4832 5187 4836
rect 5351 4832 5355 4836
rect 5527 4832 5531 4836
rect 5663 4831 5667 4835
rect 1975 4797 1979 4801
rect 2391 4796 2395 4800
rect 2527 4796 2531 4800
rect 2663 4796 2667 4800
rect 2807 4796 2811 4800
rect 2951 4796 2955 4800
rect 3095 4796 3099 4800
rect 3239 4796 3243 4800
rect 3383 4796 3387 4800
rect 3527 4796 3531 4800
rect 3799 4797 3803 4801
rect 1975 4780 1979 4784
rect 2363 4781 2367 4785
rect 2499 4781 2503 4785
rect 2635 4781 2639 4785
rect 2779 4781 2783 4785
rect 2923 4781 2927 4785
rect 3067 4781 3071 4785
rect 3211 4781 3215 4785
rect 3355 4781 3359 4785
rect 3499 4781 3503 4785
rect 3799 4780 3803 4784
rect 3839 4753 3843 4757
rect 4855 4752 4859 4756
rect 4991 4752 4995 4756
rect 5127 4752 5131 4756
rect 5263 4752 5267 4756
rect 5399 4752 5403 4756
rect 5535 4752 5539 4756
rect 5663 4753 5667 4757
rect 3839 4736 3843 4740
rect 4827 4737 4831 4741
rect 4963 4737 4967 4741
rect 5099 4737 5103 4741
rect 5235 4737 5239 4741
rect 5371 4737 5375 4741
rect 5507 4737 5511 4741
rect 5663 4736 5667 4740
rect 111 4720 115 4724
rect 131 4719 135 4723
rect 267 4719 271 4723
rect 403 4719 407 4723
rect 539 4719 543 4723
rect 675 4719 679 4723
rect 1935 4720 1939 4724
rect 111 4703 115 4707
rect 159 4704 163 4708
rect 295 4704 299 4708
rect 431 4704 435 4708
rect 567 4704 571 4708
rect 703 4704 707 4708
rect 1935 4703 1939 4707
rect 111 4641 115 4645
rect 159 4640 163 4644
rect 295 4640 299 4644
rect 431 4640 435 4644
rect 567 4640 571 4644
rect 703 4640 707 4644
rect 1935 4641 1939 4645
rect 1975 4640 1979 4644
rect 1995 4639 1999 4643
rect 2131 4639 2135 4643
rect 2267 4639 2271 4643
rect 2427 4639 2431 4643
rect 2587 4639 2591 4643
rect 2747 4639 2751 4643
rect 2907 4639 2911 4643
rect 3067 4639 3071 4643
rect 3235 4639 3239 4643
rect 3799 4640 3803 4644
rect 111 4624 115 4628
rect 131 4625 135 4629
rect 267 4625 271 4629
rect 403 4625 407 4629
rect 539 4625 543 4629
rect 675 4625 679 4629
rect 1935 4624 1939 4628
rect 1975 4623 1979 4627
rect 2023 4624 2027 4628
rect 2159 4624 2163 4628
rect 2295 4624 2299 4628
rect 2455 4624 2459 4628
rect 2615 4624 2619 4628
rect 2775 4624 2779 4628
rect 2935 4624 2939 4628
rect 3095 4624 3099 4628
rect 3263 4624 3267 4628
rect 3799 4623 3803 4627
rect 3839 4584 3843 4588
rect 4715 4583 4719 4587
rect 4859 4583 4863 4587
rect 5011 4583 5015 4587
rect 5171 4583 5175 4587
rect 5339 4583 5343 4587
rect 5515 4583 5519 4587
rect 5663 4584 5667 4588
rect 1975 4565 1979 4569
rect 2023 4564 2027 4568
rect 2175 4564 2179 4568
rect 2351 4564 2355 4568
rect 2527 4564 2531 4568
rect 2695 4564 2699 4568
rect 2871 4564 2875 4568
rect 3047 4564 3051 4568
rect 3799 4565 3803 4569
rect 3839 4567 3843 4571
rect 4743 4568 4747 4572
rect 4887 4568 4891 4572
rect 5039 4568 5043 4572
rect 5199 4568 5203 4572
rect 5367 4568 5371 4572
rect 5543 4568 5547 4572
rect 5663 4567 5667 4571
rect 1975 4548 1979 4552
rect 1995 4549 1999 4553
rect 2147 4549 2151 4553
rect 2323 4549 2327 4553
rect 2499 4549 2503 4553
rect 2667 4549 2671 4553
rect 2843 4549 2847 4553
rect 3019 4549 3023 4553
rect 3799 4548 3803 4552
rect 3839 4485 3843 4489
rect 3887 4484 3891 4488
rect 111 4480 115 4484
rect 299 4479 303 4483
rect 491 4479 495 4483
rect 691 4479 695 4483
rect 907 4479 911 4483
rect 1123 4479 1127 4483
rect 1347 4479 1351 4483
rect 1579 4479 1583 4483
rect 1787 4479 1791 4483
rect 1935 4480 1939 4484
rect 4063 4484 4067 4488
rect 4279 4484 4283 4488
rect 4503 4484 4507 4488
rect 4751 4484 4755 4488
rect 5007 4484 5011 4488
rect 5271 4484 5275 4488
rect 5543 4484 5547 4488
rect 5663 4485 5667 4489
rect 111 4463 115 4467
rect 327 4464 331 4468
rect 519 4464 523 4468
rect 719 4464 723 4468
rect 935 4464 939 4468
rect 1151 4464 1155 4468
rect 1375 4464 1379 4468
rect 1607 4464 1611 4468
rect 3839 4468 3843 4472
rect 3859 4469 3863 4473
rect 4035 4469 4039 4473
rect 4251 4469 4255 4473
rect 4475 4469 4479 4473
rect 4723 4469 4727 4473
rect 4979 4469 4983 4473
rect 5243 4469 5247 4473
rect 5515 4469 5519 4473
rect 5663 4468 5667 4472
rect 1815 4464 1819 4468
rect 1935 4463 1939 4467
rect 111 4405 115 4409
rect 559 4404 563 4408
rect 719 4404 723 4408
rect 887 4404 891 4408
rect 1063 4404 1067 4408
rect 1247 4404 1251 4408
rect 1439 4404 1443 4408
rect 1631 4404 1635 4408
rect 1815 4404 1819 4408
rect 1935 4405 1939 4409
rect 111 4388 115 4392
rect 531 4389 535 4393
rect 691 4389 695 4393
rect 859 4389 863 4393
rect 1035 4389 1039 4393
rect 1219 4389 1223 4393
rect 1411 4389 1415 4393
rect 1603 4389 1607 4393
rect 1787 4389 1791 4393
rect 1935 4388 1939 4392
rect 1975 4376 1979 4380
rect 2571 4375 2575 4379
rect 3123 4375 3127 4379
rect 3651 4375 3655 4379
rect 3799 4376 3803 4380
rect 1975 4359 1979 4363
rect 2599 4360 2603 4364
rect 3151 4360 3155 4364
rect 3679 4360 3683 4364
rect 3799 4359 3803 4363
rect 3839 4336 3843 4340
rect 3859 4335 3863 4339
rect 3995 4335 3999 4339
rect 4131 4335 4135 4339
rect 4267 4335 4271 4339
rect 4403 4335 4407 4339
rect 4587 4335 4591 4339
rect 4795 4335 4799 4339
rect 5027 4335 5031 4339
rect 5275 4335 5279 4339
rect 5515 4335 5519 4339
rect 5663 4336 5667 4340
rect 3839 4319 3843 4323
rect 3887 4320 3891 4324
rect 4023 4320 4027 4324
rect 4159 4320 4163 4324
rect 4295 4320 4299 4324
rect 4431 4320 4435 4324
rect 4615 4320 4619 4324
rect 4823 4320 4827 4324
rect 5055 4320 5059 4324
rect 5303 4320 5307 4324
rect 5543 4320 5547 4324
rect 5663 4319 5667 4323
rect 1975 4297 1979 4301
rect 2399 4296 2403 4300
rect 2599 4296 2603 4300
rect 2791 4296 2795 4300
rect 2983 4296 2987 4300
rect 3167 4296 3171 4300
rect 3343 4296 3347 4300
rect 3519 4296 3523 4300
rect 3679 4296 3683 4300
rect 3799 4297 3803 4301
rect 1975 4280 1979 4284
rect 2371 4281 2375 4285
rect 2571 4281 2575 4285
rect 2763 4281 2767 4285
rect 2955 4281 2959 4285
rect 3139 4281 3143 4285
rect 3315 4281 3319 4285
rect 3491 4281 3495 4285
rect 3651 4281 3655 4285
rect 3799 4280 3803 4284
rect 3839 4261 3843 4265
rect 4047 4260 4051 4264
rect 4223 4260 4227 4264
rect 4431 4260 4435 4264
rect 4679 4260 4683 4264
rect 4959 4260 4963 4264
rect 5255 4260 5259 4264
rect 5543 4260 5547 4264
rect 5663 4261 5667 4265
rect 111 4248 115 4252
rect 747 4247 751 4251
rect 883 4247 887 4251
rect 1019 4247 1023 4251
rect 1155 4247 1159 4251
rect 1291 4247 1295 4251
rect 1427 4247 1431 4251
rect 1563 4247 1567 4251
rect 1699 4247 1703 4251
rect 1935 4248 1939 4252
rect 3839 4244 3843 4248
rect 4019 4245 4023 4249
rect 4195 4245 4199 4249
rect 4403 4245 4407 4249
rect 4651 4245 4655 4249
rect 4931 4245 4935 4249
rect 5227 4245 5231 4249
rect 5515 4245 5519 4249
rect 5663 4244 5667 4248
rect 111 4231 115 4235
rect 775 4232 779 4236
rect 911 4232 915 4236
rect 1047 4232 1051 4236
rect 1183 4232 1187 4236
rect 1319 4232 1323 4236
rect 1455 4232 1459 4236
rect 1591 4232 1595 4236
rect 1727 4232 1731 4236
rect 1935 4231 1939 4235
rect 111 4161 115 4165
rect 727 4160 731 4164
rect 863 4160 867 4164
rect 999 4160 1003 4164
rect 1135 4160 1139 4164
rect 1271 4160 1275 4164
rect 1407 4160 1411 4164
rect 1543 4160 1547 4164
rect 1679 4160 1683 4164
rect 1815 4160 1819 4164
rect 1935 4161 1939 4165
rect 111 4144 115 4148
rect 699 4145 703 4149
rect 835 4145 839 4149
rect 971 4145 975 4149
rect 1107 4145 1111 4149
rect 1243 4145 1247 4149
rect 1379 4145 1383 4149
rect 1515 4145 1519 4149
rect 1651 4145 1655 4149
rect 1787 4145 1791 4149
rect 1935 4144 1939 4148
rect 1975 4136 1979 4140
rect 2371 4135 2375 4139
rect 2611 4135 2615 4139
rect 2835 4135 2839 4139
rect 3051 4135 3055 4139
rect 3259 4135 3263 4139
rect 3467 4135 3471 4139
rect 3651 4135 3655 4139
rect 3799 4136 3803 4140
rect 1975 4119 1979 4123
rect 2399 4120 2403 4124
rect 2639 4120 2643 4124
rect 2863 4120 2867 4124
rect 3079 4120 3083 4124
rect 3287 4120 3291 4124
rect 3495 4120 3499 4124
rect 3679 4120 3683 4124
rect 3799 4119 3803 4123
rect 1975 4057 1979 4061
rect 2375 4056 2379 4060
rect 2623 4056 2627 4060
rect 2855 4056 2859 4060
rect 3071 4056 3075 4060
rect 3279 4056 3283 4060
rect 3487 4056 3491 4060
rect 3679 4056 3683 4060
rect 3799 4057 3803 4061
rect 1975 4040 1979 4044
rect 2347 4041 2351 4045
rect 2595 4041 2599 4045
rect 2827 4041 2831 4045
rect 3043 4041 3047 4045
rect 3251 4041 3255 4045
rect 3459 4041 3463 4045
rect 3651 4041 3655 4045
rect 3799 4040 3803 4044
rect 3839 4028 3843 4032
rect 5515 4027 5519 4031
rect 5663 4028 5667 4032
rect 3839 4011 3843 4015
rect 5543 4012 5547 4016
rect 5663 4011 5667 4015
rect 111 4000 115 4004
rect 627 3999 631 4003
rect 763 3999 767 4003
rect 899 3999 903 4003
rect 1035 3999 1039 4003
rect 1171 3999 1175 4003
rect 1307 3999 1311 4003
rect 1443 3999 1447 4003
rect 1579 3999 1583 4003
rect 1715 3999 1719 4003
rect 1935 4000 1939 4004
rect 111 3983 115 3987
rect 655 3984 659 3988
rect 791 3984 795 3988
rect 927 3984 931 3988
rect 1063 3984 1067 3988
rect 1199 3984 1203 3988
rect 1335 3984 1339 3988
rect 1471 3984 1475 3988
rect 1607 3984 1611 3988
rect 1743 3984 1747 3988
rect 1935 3983 1939 3987
rect 3839 3945 3843 3949
rect 4183 3944 4187 3948
rect 4319 3944 4323 3948
rect 4455 3944 4459 3948
rect 4591 3944 4595 3948
rect 4727 3944 4731 3948
rect 4863 3944 4867 3948
rect 4999 3944 5003 3948
rect 5135 3944 5139 3948
rect 5271 3944 5275 3948
rect 5407 3944 5411 3948
rect 5543 3944 5547 3948
rect 5663 3945 5667 3949
rect 3839 3928 3843 3932
rect 4155 3929 4159 3933
rect 4291 3929 4295 3933
rect 4427 3929 4431 3933
rect 4563 3929 4567 3933
rect 4699 3929 4703 3933
rect 4835 3929 4839 3933
rect 4971 3929 4975 3933
rect 5107 3929 5111 3933
rect 5243 3929 5247 3933
rect 5379 3929 5383 3933
rect 5515 3929 5519 3933
rect 5663 3928 5667 3932
rect 111 3913 115 3917
rect 599 3912 603 3916
rect 743 3912 747 3916
rect 895 3912 899 3916
rect 1047 3912 1051 3916
rect 1199 3912 1203 3916
rect 1359 3912 1363 3916
rect 1519 3912 1523 3916
rect 1679 3912 1683 3916
rect 1935 3913 1939 3917
rect 1975 3908 1979 3912
rect 2323 3907 2327 3911
rect 2571 3907 2575 3911
rect 2803 3907 2807 3911
rect 3027 3907 3031 3911
rect 3243 3907 3247 3911
rect 3459 3907 3463 3911
rect 3651 3907 3655 3911
rect 3799 3908 3803 3912
rect 111 3896 115 3900
rect 571 3897 575 3901
rect 715 3897 719 3901
rect 867 3897 871 3901
rect 1019 3897 1023 3901
rect 1171 3897 1175 3901
rect 1331 3897 1335 3901
rect 1491 3897 1495 3901
rect 1651 3897 1655 3901
rect 1935 3896 1939 3900
rect 1975 3891 1979 3895
rect 2351 3892 2355 3896
rect 2599 3892 2603 3896
rect 2831 3892 2835 3896
rect 3055 3892 3059 3896
rect 3271 3892 3275 3896
rect 3487 3892 3491 3896
rect 3679 3892 3683 3896
rect 3799 3891 3803 3895
rect 1975 3829 1979 3833
rect 2239 3828 2243 3832
rect 2479 3828 2483 3832
rect 2703 3828 2707 3832
rect 2919 3828 2923 3832
rect 3119 3828 3123 3832
rect 3311 3828 3315 3832
rect 3503 3828 3507 3832
rect 3679 3828 3683 3832
rect 3799 3829 3803 3833
rect 1975 3812 1979 3816
rect 2211 3813 2215 3817
rect 2451 3813 2455 3817
rect 2675 3813 2679 3817
rect 2891 3813 2895 3817
rect 3091 3813 3095 3817
rect 3283 3813 3287 3817
rect 3475 3813 3479 3817
rect 3651 3813 3655 3817
rect 3799 3812 3803 3816
rect 3839 3764 3843 3768
rect 4139 3763 4143 3767
rect 4323 3763 4327 3767
rect 4531 3763 4535 3767
rect 4763 3763 4767 3767
rect 5011 3763 5015 3767
rect 5275 3763 5279 3767
rect 5515 3763 5519 3767
rect 5663 3764 5667 3768
rect 111 3756 115 3760
rect 427 3755 431 3759
rect 587 3755 591 3759
rect 755 3755 759 3759
rect 923 3755 927 3759
rect 1099 3755 1103 3759
rect 1275 3755 1279 3759
rect 1459 3755 1463 3759
rect 1643 3755 1647 3759
rect 1935 3756 1939 3760
rect 3839 3747 3843 3751
rect 4167 3748 4171 3752
rect 4351 3748 4355 3752
rect 4559 3748 4563 3752
rect 4791 3748 4795 3752
rect 5039 3748 5043 3752
rect 5303 3748 5307 3752
rect 5543 3748 5547 3752
rect 5663 3747 5667 3751
rect 111 3739 115 3743
rect 455 3740 459 3744
rect 615 3740 619 3744
rect 783 3740 787 3744
rect 951 3740 955 3744
rect 1127 3740 1131 3744
rect 1303 3740 1307 3744
rect 1487 3740 1491 3744
rect 1671 3740 1675 3744
rect 1935 3739 1939 3743
rect 111 3669 115 3673
rect 327 3668 331 3672
rect 495 3668 499 3672
rect 679 3668 683 3672
rect 863 3668 867 3672
rect 1055 3668 1059 3672
rect 1255 3668 1259 3672
rect 1455 3668 1459 3672
rect 1655 3668 1659 3672
rect 1935 3669 1939 3673
rect 1975 3672 1979 3676
rect 2227 3671 2231 3675
rect 2451 3671 2455 3675
rect 2667 3671 2671 3675
rect 2875 3671 2879 3675
rect 3075 3671 3079 3675
rect 3275 3671 3279 3675
rect 3475 3671 3479 3675
rect 3799 3672 3803 3676
rect 3839 3669 3843 3673
rect 4303 3668 4307 3672
rect 4479 3668 4483 3672
rect 4671 3668 4675 3672
rect 4879 3668 4883 3672
rect 5103 3668 5107 3672
rect 5335 3668 5339 3672
rect 5543 3668 5547 3672
rect 5663 3669 5667 3673
rect 111 3652 115 3656
rect 299 3653 303 3657
rect 467 3653 471 3657
rect 651 3653 655 3657
rect 835 3653 839 3657
rect 1027 3653 1031 3657
rect 1227 3653 1231 3657
rect 1427 3653 1431 3657
rect 1627 3653 1631 3657
rect 1935 3652 1939 3656
rect 1975 3655 1979 3659
rect 2255 3656 2259 3660
rect 2479 3656 2483 3660
rect 2695 3656 2699 3660
rect 2903 3656 2907 3660
rect 3103 3656 3107 3660
rect 3303 3656 3307 3660
rect 3503 3656 3507 3660
rect 3799 3655 3803 3659
rect 3839 3652 3843 3656
rect 4275 3653 4279 3657
rect 4451 3653 4455 3657
rect 4643 3653 4647 3657
rect 4851 3653 4855 3657
rect 5075 3653 5079 3657
rect 5307 3653 5311 3657
rect 5515 3653 5519 3657
rect 5663 3652 5667 3656
rect 1975 3593 1979 3597
rect 2135 3592 2139 3596
rect 2311 3592 2315 3596
rect 2479 3592 2483 3596
rect 2647 3592 2651 3596
rect 2807 3592 2811 3596
rect 2967 3592 2971 3596
rect 3135 3592 3139 3596
rect 3303 3592 3307 3596
rect 3799 3593 3803 3597
rect 1975 3576 1979 3580
rect 2107 3577 2111 3581
rect 2283 3577 2287 3581
rect 2451 3577 2455 3581
rect 2619 3577 2623 3581
rect 2779 3577 2783 3581
rect 2939 3577 2943 3581
rect 3107 3577 3111 3581
rect 3275 3577 3279 3581
rect 3799 3576 3803 3580
rect 111 3500 115 3504
rect 203 3499 207 3503
rect 379 3499 383 3503
rect 563 3499 567 3503
rect 755 3499 759 3503
rect 955 3499 959 3503
rect 1163 3499 1167 3503
rect 1379 3499 1383 3503
rect 1595 3499 1599 3503
rect 1935 3500 1939 3504
rect 3839 3492 3843 3496
rect 4555 3491 4559 3495
rect 4699 3491 4703 3495
rect 4851 3491 4855 3495
rect 5011 3491 5015 3495
rect 5179 3491 5183 3495
rect 5355 3491 5359 3495
rect 5515 3491 5519 3495
rect 5663 3492 5667 3496
rect 111 3483 115 3487
rect 231 3484 235 3488
rect 407 3484 411 3488
rect 591 3484 595 3488
rect 783 3484 787 3488
rect 983 3484 987 3488
rect 1191 3484 1195 3488
rect 1407 3484 1411 3488
rect 1623 3484 1627 3488
rect 1935 3483 1939 3487
rect 3839 3475 3843 3479
rect 4583 3476 4587 3480
rect 4727 3476 4731 3480
rect 4879 3476 4883 3480
rect 5039 3476 5043 3480
rect 5207 3476 5211 3480
rect 5383 3476 5387 3480
rect 5543 3476 5547 3480
rect 5663 3475 5667 3479
rect 1975 3420 1979 3424
rect 2035 3419 2039 3423
rect 2187 3419 2191 3423
rect 2339 3419 2343 3423
rect 2491 3419 2495 3423
rect 2643 3419 2647 3423
rect 2795 3419 2799 3423
rect 2947 3419 2951 3423
rect 3099 3419 3103 3423
rect 3799 3420 3803 3424
rect 111 3405 115 3409
rect 255 3404 259 3408
rect 471 3404 475 3408
rect 695 3404 699 3408
rect 919 3404 923 3408
rect 1143 3404 1147 3408
rect 1367 3404 1371 3408
rect 1591 3404 1595 3408
rect 1935 3405 1939 3409
rect 1975 3403 1979 3407
rect 2063 3404 2067 3408
rect 2215 3404 2219 3408
rect 2367 3404 2371 3408
rect 2519 3404 2523 3408
rect 2671 3404 2675 3408
rect 2823 3404 2827 3408
rect 2975 3404 2979 3408
rect 3127 3404 3131 3408
rect 3799 3403 3803 3407
rect 3839 3405 3843 3409
rect 4903 3404 4907 3408
rect 5039 3404 5043 3408
rect 5175 3404 5179 3408
rect 5311 3404 5315 3408
rect 5447 3404 5451 3408
rect 5663 3405 5667 3409
rect 111 3388 115 3392
rect 227 3389 231 3393
rect 443 3389 447 3393
rect 667 3389 671 3393
rect 891 3389 895 3393
rect 1115 3389 1119 3393
rect 1339 3389 1343 3393
rect 1563 3389 1567 3393
rect 1935 3388 1939 3392
rect 3839 3388 3843 3392
rect 4875 3389 4879 3393
rect 5011 3389 5015 3393
rect 5147 3389 5151 3393
rect 5283 3389 5287 3393
rect 5419 3389 5423 3393
rect 5663 3388 5667 3392
rect 1975 3333 1979 3337
rect 2023 3332 2027 3336
rect 2191 3332 2195 3336
rect 2375 3332 2379 3336
rect 2551 3332 2555 3336
rect 2727 3332 2731 3336
rect 2895 3332 2899 3336
rect 3071 3332 3075 3336
rect 3247 3332 3251 3336
rect 3799 3333 3803 3337
rect 1975 3316 1979 3320
rect 1995 3317 1999 3321
rect 2163 3317 2167 3321
rect 2347 3317 2351 3321
rect 2523 3317 2527 3321
rect 2699 3317 2703 3321
rect 2867 3317 2871 3321
rect 3043 3317 3047 3321
rect 3219 3317 3223 3321
rect 3799 3316 3803 3320
rect 3839 3256 3843 3260
rect 4699 3255 4703 3259
rect 4835 3255 4839 3259
rect 4971 3255 4975 3259
rect 5107 3255 5111 3259
rect 5243 3255 5247 3259
rect 5379 3255 5383 3259
rect 5515 3255 5519 3259
rect 5663 3256 5667 3260
rect 111 3240 115 3244
rect 211 3239 215 3243
rect 419 3239 423 3243
rect 635 3239 639 3243
rect 851 3239 855 3243
rect 1075 3239 1079 3243
rect 1299 3239 1303 3243
rect 1523 3239 1527 3243
rect 1935 3240 1939 3244
rect 3839 3239 3843 3243
rect 4727 3240 4731 3244
rect 4863 3240 4867 3244
rect 4999 3240 5003 3244
rect 5135 3240 5139 3244
rect 5271 3240 5275 3244
rect 5407 3240 5411 3244
rect 5543 3240 5547 3244
rect 5663 3239 5667 3243
rect 111 3223 115 3227
rect 239 3224 243 3228
rect 447 3224 451 3228
rect 663 3224 667 3228
rect 879 3224 883 3228
rect 1103 3224 1107 3228
rect 1327 3224 1331 3228
rect 1551 3224 1555 3228
rect 1935 3223 1939 3227
rect 1975 3180 1979 3184
rect 1995 3179 1999 3183
rect 2211 3179 2215 3183
rect 2435 3179 2439 3183
rect 2651 3179 2655 3183
rect 2851 3179 2855 3183
rect 3051 3179 3055 3183
rect 3251 3179 3255 3183
rect 3451 3179 3455 3183
rect 3799 3180 3803 3184
rect 3839 3173 3843 3177
rect 4567 3172 4571 3176
rect 4743 3172 4747 3176
rect 4935 3172 4939 3176
rect 5135 3172 5139 3176
rect 5351 3172 5355 3176
rect 5543 3172 5547 3176
rect 5663 3173 5667 3177
rect 1975 3163 1979 3167
rect 2023 3164 2027 3168
rect 2239 3164 2243 3168
rect 2463 3164 2467 3168
rect 2679 3164 2683 3168
rect 2879 3164 2883 3168
rect 3079 3164 3083 3168
rect 3279 3164 3283 3168
rect 3479 3164 3483 3168
rect 3799 3163 3803 3167
rect 3839 3156 3843 3160
rect 4539 3157 4543 3161
rect 4715 3157 4719 3161
rect 4907 3157 4911 3161
rect 5107 3157 5111 3161
rect 5323 3157 5327 3161
rect 5515 3157 5519 3161
rect 5663 3156 5667 3160
rect 111 3149 115 3153
rect 303 3148 307 3152
rect 543 3148 547 3152
rect 783 3148 787 3152
rect 1023 3148 1027 3152
rect 1263 3148 1267 3152
rect 1511 3148 1515 3152
rect 1935 3149 1939 3153
rect 111 3132 115 3136
rect 275 3133 279 3137
rect 515 3133 519 3137
rect 755 3133 759 3137
rect 995 3133 999 3137
rect 1235 3133 1239 3137
rect 1483 3133 1487 3137
rect 1935 3132 1939 3136
rect 1975 3105 1979 3109
rect 2023 3104 2027 3108
rect 2327 3104 2331 3108
rect 2631 3104 2635 3108
rect 2911 3104 2915 3108
rect 3175 3104 3179 3108
rect 3439 3104 3443 3108
rect 3679 3104 3683 3108
rect 3799 3105 3803 3109
rect 1975 3088 1979 3092
rect 1995 3089 1999 3093
rect 2299 3089 2303 3093
rect 2603 3089 2607 3093
rect 2883 3089 2887 3093
rect 3147 3089 3151 3093
rect 3411 3089 3415 3093
rect 3651 3089 3655 3093
rect 3799 3088 3803 3092
rect 3839 3020 3843 3024
rect 4307 3019 4311 3023
rect 4483 3019 4487 3023
rect 4675 3019 4679 3023
rect 4875 3019 4879 3023
rect 5091 3019 5095 3023
rect 5315 3019 5319 3023
rect 5515 3019 5519 3023
rect 5663 3020 5667 3024
rect 111 3000 115 3004
rect 355 2999 359 3003
rect 627 2999 631 3003
rect 883 2999 887 3003
rect 1123 2999 1127 3003
rect 1355 2999 1359 3003
rect 1579 2999 1583 3003
rect 1787 2999 1791 3003
rect 1935 3000 1939 3004
rect 3839 3003 3843 3007
rect 4335 3004 4339 3008
rect 4511 3004 4515 3008
rect 4703 3004 4707 3008
rect 4903 3004 4907 3008
rect 5119 3004 5123 3008
rect 5343 3004 5347 3008
rect 5543 3004 5547 3008
rect 5663 3003 5667 3007
rect 111 2983 115 2987
rect 383 2984 387 2988
rect 655 2984 659 2988
rect 911 2984 915 2988
rect 1151 2984 1155 2988
rect 1383 2984 1387 2988
rect 1607 2984 1611 2988
rect 1815 2984 1819 2988
rect 1935 2983 1939 2987
rect 1975 2948 1979 2952
rect 3107 2947 3111 2951
rect 3243 2947 3247 2951
rect 3379 2947 3383 2951
rect 3515 2947 3519 2951
rect 3651 2947 3655 2951
rect 3799 2948 3803 2952
rect 3839 2941 3843 2945
rect 3887 2940 3891 2944
rect 4023 2940 4027 2944
rect 4175 2940 4179 2944
rect 4391 2940 4395 2944
rect 4639 2940 4643 2944
rect 4919 2940 4923 2944
rect 5223 2940 5227 2944
rect 5527 2940 5531 2944
rect 5663 2941 5667 2945
rect 1975 2931 1979 2935
rect 3135 2932 3139 2936
rect 3271 2932 3275 2936
rect 3407 2932 3411 2936
rect 3543 2932 3547 2936
rect 3679 2932 3683 2936
rect 3799 2931 3803 2935
rect 111 2925 115 2929
rect 343 2924 347 2928
rect 551 2924 555 2928
rect 759 2924 763 2928
rect 951 2924 955 2928
rect 1135 2924 1139 2928
rect 1311 2924 1315 2928
rect 1487 2924 1491 2928
rect 1663 2924 1667 2928
rect 1815 2924 1819 2928
rect 1935 2925 1939 2929
rect 3839 2924 3843 2928
rect 3859 2925 3863 2929
rect 3995 2925 3999 2929
rect 4147 2925 4151 2929
rect 4363 2925 4367 2929
rect 4611 2925 4615 2929
rect 4891 2925 4895 2929
rect 5195 2925 5199 2929
rect 5499 2925 5503 2929
rect 5663 2924 5667 2928
rect 111 2908 115 2912
rect 315 2909 319 2913
rect 523 2909 527 2913
rect 731 2909 735 2913
rect 923 2909 927 2913
rect 1107 2909 1111 2913
rect 1283 2909 1287 2913
rect 1459 2909 1463 2913
rect 1635 2909 1639 2913
rect 1787 2909 1791 2913
rect 1935 2908 1939 2912
rect 3839 2792 3843 2796
rect 3859 2791 3863 2795
rect 3995 2791 3999 2795
rect 4131 2791 4135 2795
rect 4267 2791 4271 2795
rect 4403 2791 4407 2795
rect 4539 2791 4543 2795
rect 4675 2791 4679 2795
rect 4811 2791 4815 2795
rect 5663 2792 5667 2796
rect 3839 2775 3843 2779
rect 3887 2776 3891 2780
rect 4023 2776 4027 2780
rect 4159 2776 4163 2780
rect 4295 2776 4299 2780
rect 4431 2776 4435 2780
rect 4567 2776 4571 2780
rect 4703 2776 4707 2780
rect 4839 2776 4843 2780
rect 5663 2775 5667 2779
rect 111 2764 115 2768
rect 363 2763 367 2767
rect 563 2763 567 2767
rect 755 2763 759 2767
rect 939 2763 943 2767
rect 1115 2763 1119 2767
rect 1283 2763 1287 2767
rect 1451 2763 1455 2767
rect 1619 2763 1623 2767
rect 1787 2763 1791 2767
rect 1935 2764 1939 2768
rect 111 2747 115 2751
rect 391 2748 395 2752
rect 591 2748 595 2752
rect 783 2748 787 2752
rect 967 2748 971 2752
rect 1143 2748 1147 2752
rect 1311 2748 1315 2752
rect 1479 2748 1483 2752
rect 1647 2748 1651 2752
rect 1815 2748 1819 2752
rect 1935 2747 1939 2751
rect 3839 2701 3843 2705
rect 3887 2700 3891 2704
rect 4023 2700 4027 2704
rect 4159 2700 4163 2704
rect 4295 2700 4299 2704
rect 4431 2700 4435 2704
rect 4567 2700 4571 2704
rect 4711 2700 4715 2704
rect 4879 2700 4883 2704
rect 5063 2700 5067 2704
rect 5255 2700 5259 2704
rect 5447 2700 5451 2704
rect 5663 2701 5667 2705
rect 111 2685 115 2689
rect 447 2684 451 2688
rect 615 2684 619 2688
rect 775 2684 779 2688
rect 935 2684 939 2688
rect 1087 2684 1091 2688
rect 1239 2684 1243 2688
rect 1383 2684 1387 2688
rect 1535 2684 1539 2688
rect 1679 2684 1683 2688
rect 1815 2684 1819 2688
rect 1935 2685 1939 2689
rect 3839 2684 3843 2688
rect 3859 2685 3863 2689
rect 3995 2685 3999 2689
rect 4131 2685 4135 2689
rect 4267 2685 4271 2689
rect 4403 2685 4407 2689
rect 4539 2685 4543 2689
rect 4683 2685 4687 2689
rect 4851 2685 4855 2689
rect 5035 2685 5039 2689
rect 5227 2685 5231 2689
rect 5419 2685 5423 2689
rect 5663 2684 5667 2688
rect 111 2668 115 2672
rect 419 2669 423 2673
rect 587 2669 591 2673
rect 747 2669 751 2673
rect 907 2669 911 2673
rect 1059 2669 1063 2673
rect 1211 2669 1215 2673
rect 1355 2669 1359 2673
rect 1507 2669 1511 2673
rect 1651 2669 1655 2673
rect 1787 2669 1791 2673
rect 1935 2668 1939 2672
rect 1975 2605 1979 2609
rect 3271 2604 3275 2608
rect 3407 2604 3411 2608
rect 3543 2604 3547 2608
rect 3679 2604 3683 2608
rect 3799 2605 3803 2609
rect 1975 2588 1979 2592
rect 3243 2589 3247 2593
rect 3379 2589 3383 2593
rect 3515 2589 3519 2593
rect 3651 2589 3655 2593
rect 3799 2588 3803 2592
rect 111 2532 115 2536
rect 235 2531 239 2535
rect 435 2531 439 2535
rect 627 2531 631 2535
rect 811 2531 815 2535
rect 987 2531 991 2535
rect 1155 2531 1159 2535
rect 1323 2531 1327 2535
rect 1483 2531 1487 2535
rect 1643 2531 1647 2535
rect 1787 2531 1791 2535
rect 1935 2532 1939 2536
rect 3839 2536 3843 2540
rect 4179 2535 4183 2539
rect 4395 2535 4399 2539
rect 4643 2535 4647 2539
rect 4907 2535 4911 2539
rect 5187 2535 5191 2539
rect 5467 2535 5471 2539
rect 5663 2536 5667 2540
rect 111 2515 115 2519
rect 263 2516 267 2520
rect 463 2516 467 2520
rect 655 2516 659 2520
rect 839 2516 843 2520
rect 1015 2516 1019 2520
rect 1183 2516 1187 2520
rect 1351 2516 1355 2520
rect 1511 2516 1515 2520
rect 1671 2516 1675 2520
rect 1815 2516 1819 2520
rect 1935 2515 1939 2519
rect 3839 2519 3843 2523
rect 4207 2520 4211 2524
rect 4423 2520 4427 2524
rect 4671 2520 4675 2524
rect 4935 2520 4939 2524
rect 5215 2520 5219 2524
rect 5495 2520 5499 2524
rect 5663 2519 5667 2523
rect 3839 2461 3843 2465
rect 4535 2460 4539 2464
rect 1975 2456 1979 2460
rect 1995 2455 1999 2459
rect 2251 2455 2255 2459
rect 2523 2455 2527 2459
rect 2771 2455 2775 2459
rect 3003 2455 3007 2459
rect 3227 2455 3231 2459
rect 3451 2455 3455 2459
rect 3651 2455 3655 2459
rect 3799 2456 3803 2460
rect 4759 2460 4763 2464
rect 4983 2460 4987 2464
rect 5215 2460 5219 2464
rect 5447 2460 5451 2464
rect 5663 2461 5667 2465
rect 111 2449 115 2453
rect 223 2448 227 2452
rect 423 2448 427 2452
rect 623 2448 627 2452
rect 815 2448 819 2452
rect 1015 2448 1019 2452
rect 1215 2448 1219 2452
rect 1935 2449 1939 2453
rect 1975 2439 1979 2443
rect 2023 2440 2027 2444
rect 2279 2440 2283 2444
rect 2551 2440 2555 2444
rect 2799 2440 2803 2444
rect 3031 2440 3035 2444
rect 3255 2440 3259 2444
rect 3479 2440 3483 2444
rect 3839 2444 3843 2448
rect 4507 2445 4511 2449
rect 4731 2445 4735 2449
rect 4955 2445 4959 2449
rect 5187 2445 5191 2449
rect 5419 2445 5423 2449
rect 5663 2444 5667 2448
rect 3679 2440 3683 2444
rect 3799 2439 3803 2443
rect 111 2432 115 2436
rect 195 2433 199 2437
rect 395 2433 399 2437
rect 595 2433 599 2437
rect 787 2433 791 2437
rect 987 2433 991 2437
rect 1187 2433 1191 2437
rect 1935 2432 1939 2436
rect 1975 2381 1979 2385
rect 2055 2380 2059 2384
rect 2215 2380 2219 2384
rect 2375 2380 2379 2384
rect 2543 2380 2547 2384
rect 2711 2380 2715 2384
rect 2871 2380 2875 2384
rect 3031 2380 3035 2384
rect 3191 2380 3195 2384
rect 3359 2380 3363 2384
rect 3527 2380 3531 2384
rect 3799 2381 3803 2385
rect 1975 2364 1979 2368
rect 2027 2365 2031 2369
rect 2187 2365 2191 2369
rect 2347 2365 2351 2369
rect 2515 2365 2519 2369
rect 2683 2365 2687 2369
rect 2843 2365 2847 2369
rect 3003 2365 3007 2369
rect 3163 2365 3167 2369
rect 3331 2365 3335 2369
rect 3499 2365 3503 2369
rect 3799 2364 3803 2368
rect 3839 2312 3843 2316
rect 4707 2311 4711 2315
rect 4867 2311 4871 2315
rect 5027 2311 5031 2315
rect 5187 2311 5191 2315
rect 5347 2311 5351 2315
rect 5515 2311 5519 2315
rect 5663 2312 5667 2316
rect 3839 2295 3843 2299
rect 4735 2296 4739 2300
rect 4895 2296 4899 2300
rect 5055 2296 5059 2300
rect 5215 2296 5219 2300
rect 5375 2296 5379 2300
rect 5543 2296 5547 2300
rect 5663 2295 5667 2299
rect 111 2288 115 2292
rect 131 2287 135 2291
rect 291 2287 295 2291
rect 483 2287 487 2291
rect 675 2287 679 2291
rect 867 2287 871 2291
rect 1935 2288 1939 2292
rect 111 2271 115 2275
rect 159 2272 163 2276
rect 319 2272 323 2276
rect 511 2272 515 2276
rect 703 2272 707 2276
rect 895 2272 899 2276
rect 1935 2271 1939 2275
rect 1975 2224 1979 2228
rect 2139 2223 2143 2227
rect 2275 2223 2279 2227
rect 2411 2223 2415 2227
rect 2547 2223 2551 2227
rect 2683 2223 2687 2227
rect 2819 2223 2823 2227
rect 2955 2223 2959 2227
rect 3091 2223 3095 2227
rect 3227 2223 3231 2227
rect 3363 2223 3367 2227
rect 3799 2224 3803 2228
rect 3839 2225 3843 2229
rect 4735 2224 4739 2228
rect 4887 2224 4891 2228
rect 5047 2224 5051 2228
rect 5215 2224 5219 2228
rect 5391 2224 5395 2228
rect 5543 2224 5547 2228
rect 5663 2225 5667 2229
rect 111 2213 115 2217
rect 159 2212 163 2216
rect 295 2212 299 2216
rect 439 2212 443 2216
rect 591 2212 595 2216
rect 743 2212 747 2216
rect 1935 2213 1939 2217
rect 1975 2207 1979 2211
rect 2167 2208 2171 2212
rect 2303 2208 2307 2212
rect 2439 2208 2443 2212
rect 2575 2208 2579 2212
rect 2711 2208 2715 2212
rect 2847 2208 2851 2212
rect 2983 2208 2987 2212
rect 3119 2208 3123 2212
rect 3255 2208 3259 2212
rect 3391 2208 3395 2212
rect 3799 2207 3803 2211
rect 3839 2208 3843 2212
rect 4707 2209 4711 2213
rect 4859 2209 4863 2213
rect 5019 2209 5023 2213
rect 5187 2209 5191 2213
rect 5363 2209 5367 2213
rect 5515 2209 5519 2213
rect 5663 2208 5667 2212
rect 111 2196 115 2200
rect 131 2197 135 2201
rect 267 2197 271 2201
rect 411 2197 415 2201
rect 563 2197 567 2201
rect 715 2197 719 2201
rect 1935 2196 1939 2200
rect 1975 2145 1979 2149
rect 2023 2144 2027 2148
rect 2159 2144 2163 2148
rect 2295 2144 2299 2148
rect 2431 2144 2435 2148
rect 2567 2144 2571 2148
rect 2703 2144 2707 2148
rect 2839 2144 2843 2148
rect 2975 2144 2979 2148
rect 3111 2144 3115 2148
rect 3247 2144 3251 2148
rect 3799 2145 3803 2149
rect 1975 2128 1979 2132
rect 1995 2129 1999 2133
rect 2131 2129 2135 2133
rect 2267 2129 2271 2133
rect 2403 2129 2407 2133
rect 2539 2129 2543 2133
rect 2675 2129 2679 2133
rect 2811 2129 2815 2133
rect 2947 2129 2951 2133
rect 3083 2129 3087 2133
rect 3219 2129 3223 2133
rect 3799 2128 3803 2132
rect 111 2064 115 2068
rect 131 2063 135 2067
rect 331 2063 335 2067
rect 555 2063 559 2067
rect 779 2063 783 2067
rect 1011 2063 1015 2067
rect 1935 2064 1939 2068
rect 3839 2068 3843 2072
rect 4787 2067 4791 2071
rect 4923 2067 4927 2071
rect 5067 2067 5071 2071
rect 5219 2067 5223 2071
rect 5379 2067 5383 2071
rect 5515 2067 5519 2071
rect 5663 2068 5667 2072
rect 111 2047 115 2051
rect 159 2048 163 2052
rect 359 2048 363 2052
rect 583 2048 587 2052
rect 807 2048 811 2052
rect 1039 2048 1043 2052
rect 1935 2047 1939 2051
rect 3839 2051 3843 2055
rect 4815 2052 4819 2056
rect 4951 2052 4955 2056
rect 5095 2052 5099 2056
rect 5247 2052 5251 2056
rect 5407 2052 5411 2056
rect 5543 2052 5547 2056
rect 5663 2051 5667 2055
rect 111 1985 115 1989
rect 159 1984 163 1988
rect 463 1984 467 1988
rect 799 1984 803 1988
rect 1143 1984 1147 1988
rect 1487 1984 1491 1988
rect 1815 1984 1819 1988
rect 1935 1985 1939 1989
rect 1975 1988 1979 1992
rect 1995 1987 1999 1991
rect 2131 1987 2135 1991
rect 2267 1987 2271 1991
rect 2403 1987 2407 1991
rect 2539 1987 2543 1991
rect 2675 1987 2679 1991
rect 2811 1987 2815 1991
rect 2947 1987 2951 1991
rect 3091 1987 3095 1991
rect 3243 1987 3247 1991
rect 3395 1987 3399 1991
rect 3799 1988 3803 1992
rect 3839 1989 3843 1993
rect 4863 1988 4867 1992
rect 4999 1988 5003 1992
rect 5135 1988 5139 1992
rect 5271 1988 5275 1992
rect 5407 1988 5411 1992
rect 5543 1988 5547 1992
rect 5663 1989 5667 1993
rect 111 1968 115 1972
rect 131 1969 135 1973
rect 435 1969 439 1973
rect 771 1969 775 1973
rect 1115 1969 1119 1973
rect 1459 1969 1463 1973
rect 1787 1969 1791 1973
rect 1935 1968 1939 1972
rect 1975 1971 1979 1975
rect 2023 1972 2027 1976
rect 2159 1972 2163 1976
rect 2295 1972 2299 1976
rect 2431 1972 2435 1976
rect 2567 1972 2571 1976
rect 2703 1972 2707 1976
rect 2839 1972 2843 1976
rect 2975 1972 2979 1976
rect 3119 1972 3123 1976
rect 3271 1972 3275 1976
rect 3423 1972 3427 1976
rect 3799 1971 3803 1975
rect 3839 1972 3843 1976
rect 4835 1973 4839 1977
rect 4971 1973 4975 1977
rect 5107 1973 5111 1977
rect 5243 1973 5247 1977
rect 5379 1973 5383 1977
rect 5515 1973 5519 1977
rect 5663 1972 5667 1976
rect 1975 1905 1979 1909
rect 2527 1904 2531 1908
rect 2663 1904 2667 1908
rect 2799 1904 2803 1908
rect 2935 1904 2939 1908
rect 3071 1904 3075 1908
rect 3207 1904 3211 1908
rect 3351 1904 3355 1908
rect 3799 1905 3803 1909
rect 1975 1888 1979 1892
rect 2499 1889 2503 1893
rect 2635 1889 2639 1893
rect 2771 1889 2775 1893
rect 2907 1889 2911 1893
rect 3043 1889 3047 1893
rect 3179 1889 3183 1893
rect 3323 1889 3327 1893
rect 3799 1888 3803 1892
rect 111 1836 115 1840
rect 195 1835 199 1839
rect 451 1835 455 1839
rect 699 1835 703 1839
rect 931 1835 935 1839
rect 1155 1835 1159 1839
rect 1371 1835 1375 1839
rect 1587 1835 1591 1839
rect 1787 1835 1791 1839
rect 1935 1836 1939 1840
rect 3839 1836 3843 1840
rect 4683 1835 4687 1839
rect 4843 1835 4847 1839
rect 5011 1835 5015 1839
rect 5179 1835 5183 1839
rect 5355 1835 5359 1839
rect 5515 1835 5519 1839
rect 5663 1836 5667 1840
rect 111 1819 115 1823
rect 223 1820 227 1824
rect 479 1820 483 1824
rect 727 1820 731 1824
rect 959 1820 963 1824
rect 1183 1820 1187 1824
rect 1399 1820 1403 1824
rect 1615 1820 1619 1824
rect 1815 1820 1819 1824
rect 1935 1819 1939 1823
rect 3839 1819 3843 1823
rect 4711 1820 4715 1824
rect 4871 1820 4875 1824
rect 5039 1820 5043 1824
rect 5207 1820 5211 1824
rect 5383 1820 5387 1824
rect 5543 1820 5547 1824
rect 5663 1819 5667 1823
rect 111 1757 115 1761
rect 231 1756 235 1760
rect 447 1756 451 1760
rect 671 1756 675 1760
rect 895 1756 899 1760
rect 1119 1756 1123 1760
rect 1343 1756 1347 1760
rect 1567 1756 1571 1760
rect 1799 1756 1803 1760
rect 1935 1757 1939 1761
rect 1975 1756 1979 1760
rect 2443 1755 2447 1759
rect 2587 1755 2591 1759
rect 2739 1755 2743 1759
rect 2891 1755 2895 1759
rect 3043 1755 3047 1759
rect 3195 1755 3199 1759
rect 3799 1756 3803 1760
rect 3839 1757 3843 1761
rect 3887 1756 3891 1760
rect 4023 1756 4027 1760
rect 4191 1756 4195 1760
rect 4367 1756 4371 1760
rect 4559 1756 4563 1760
rect 4767 1756 4771 1760
rect 4983 1756 4987 1760
rect 5215 1756 5219 1760
rect 5447 1756 5451 1760
rect 5663 1757 5667 1761
rect 111 1740 115 1744
rect 203 1741 207 1745
rect 419 1741 423 1745
rect 643 1741 647 1745
rect 867 1741 871 1745
rect 1091 1741 1095 1745
rect 1315 1741 1319 1745
rect 1539 1741 1543 1745
rect 1771 1741 1775 1745
rect 1935 1740 1939 1744
rect 1975 1739 1979 1743
rect 2471 1740 2475 1744
rect 2615 1740 2619 1744
rect 2767 1740 2771 1744
rect 2919 1740 2923 1744
rect 3071 1740 3075 1744
rect 3223 1740 3227 1744
rect 3799 1739 3803 1743
rect 3839 1740 3843 1744
rect 3859 1741 3863 1745
rect 3995 1741 3999 1745
rect 4163 1741 4167 1745
rect 4339 1741 4343 1745
rect 4531 1741 4535 1745
rect 4739 1741 4743 1745
rect 4955 1741 4959 1745
rect 5187 1741 5191 1745
rect 5419 1741 5423 1745
rect 5663 1740 5667 1744
rect 1975 1637 1979 1641
rect 2231 1636 2235 1640
rect 2599 1636 2603 1640
rect 2967 1636 2971 1640
rect 3335 1636 3339 1640
rect 3679 1636 3683 1640
rect 3799 1637 3803 1641
rect 1975 1620 1979 1624
rect 2203 1621 2207 1625
rect 2571 1621 2575 1625
rect 2939 1621 2943 1625
rect 3307 1621 3311 1625
rect 3651 1621 3655 1625
rect 3799 1620 3803 1624
rect 111 1608 115 1612
rect 275 1607 279 1611
rect 459 1607 463 1611
rect 667 1607 671 1611
rect 883 1607 887 1611
rect 1115 1607 1119 1611
rect 1355 1607 1359 1611
rect 1595 1607 1599 1611
rect 1935 1608 1939 1612
rect 3839 1608 3843 1612
rect 3859 1607 3863 1611
rect 3995 1607 3999 1611
rect 4131 1607 4135 1611
rect 4283 1607 4287 1611
rect 4483 1607 4487 1611
rect 4715 1607 4719 1611
rect 4979 1607 4983 1611
rect 5259 1607 5263 1611
rect 5515 1607 5519 1611
rect 5663 1608 5667 1612
rect 111 1591 115 1595
rect 303 1592 307 1596
rect 487 1592 491 1596
rect 695 1592 699 1596
rect 911 1592 915 1596
rect 1143 1592 1147 1596
rect 1383 1592 1387 1596
rect 1623 1592 1627 1596
rect 1935 1591 1939 1595
rect 3839 1591 3843 1595
rect 3887 1592 3891 1596
rect 4023 1592 4027 1596
rect 4159 1592 4163 1596
rect 4311 1592 4315 1596
rect 4511 1592 4515 1596
rect 4743 1592 4747 1596
rect 5007 1592 5011 1596
rect 5287 1592 5291 1596
rect 5543 1592 5547 1596
rect 5663 1591 5667 1595
rect 111 1533 115 1537
rect 383 1532 387 1536
rect 575 1532 579 1536
rect 767 1532 771 1536
rect 951 1532 955 1536
rect 1127 1532 1131 1536
rect 1303 1532 1307 1536
rect 1479 1532 1483 1536
rect 1663 1532 1667 1536
rect 1935 1533 1939 1537
rect 3839 1533 3843 1537
rect 3887 1532 3891 1536
rect 4047 1532 4051 1536
rect 4271 1532 4275 1536
rect 4543 1532 4547 1536
rect 4855 1532 4859 1536
rect 5191 1532 5195 1536
rect 5527 1532 5531 1536
rect 5663 1533 5667 1537
rect 111 1516 115 1520
rect 355 1517 359 1521
rect 547 1517 551 1521
rect 739 1517 743 1521
rect 923 1517 927 1521
rect 1099 1517 1103 1521
rect 1275 1517 1279 1521
rect 1451 1517 1455 1521
rect 1635 1517 1639 1521
rect 1935 1516 1939 1520
rect 3839 1516 3843 1520
rect 3859 1517 3863 1521
rect 4019 1517 4023 1521
rect 4243 1517 4247 1521
rect 4515 1517 4519 1521
rect 4827 1517 4831 1521
rect 5163 1517 5167 1521
rect 5499 1517 5503 1521
rect 5663 1516 5667 1520
rect 1975 1476 1979 1480
rect 1995 1475 1999 1479
rect 2275 1475 2279 1479
rect 2539 1475 2543 1479
rect 2779 1475 2783 1479
rect 3011 1475 3015 1479
rect 3235 1475 3239 1479
rect 3451 1475 3455 1479
rect 3651 1475 3655 1479
rect 3799 1476 3803 1480
rect 1975 1459 1979 1463
rect 2023 1460 2027 1464
rect 2303 1460 2307 1464
rect 2567 1460 2571 1464
rect 2807 1460 2811 1464
rect 3039 1460 3043 1464
rect 3263 1460 3267 1464
rect 3479 1460 3483 1464
rect 3679 1460 3683 1464
rect 3799 1459 3803 1463
rect 1975 1401 1979 1405
rect 2023 1400 2027 1404
rect 2191 1400 2195 1404
rect 2399 1400 2403 1404
rect 2615 1400 2619 1404
rect 2831 1400 2835 1404
rect 3055 1400 3059 1404
rect 3287 1400 3291 1404
rect 3527 1400 3531 1404
rect 3799 1401 3803 1405
rect 1975 1384 1979 1388
rect 1995 1385 1999 1389
rect 2163 1385 2167 1389
rect 2371 1385 2375 1389
rect 2587 1385 2591 1389
rect 2803 1385 2807 1389
rect 3027 1385 3031 1389
rect 3259 1385 3263 1389
rect 3499 1385 3503 1389
rect 3799 1384 3803 1388
rect 111 1364 115 1368
rect 331 1363 335 1367
rect 587 1363 591 1367
rect 843 1363 847 1367
rect 1099 1363 1103 1367
rect 1363 1363 1367 1367
rect 1935 1364 1939 1368
rect 3839 1368 3843 1372
rect 3859 1367 3863 1371
rect 3995 1367 3999 1371
rect 4147 1367 4151 1371
rect 4355 1367 4359 1371
rect 4595 1367 4599 1371
rect 4867 1367 4871 1371
rect 5163 1367 5167 1371
rect 5459 1367 5463 1371
rect 5663 1368 5667 1372
rect 111 1347 115 1351
rect 359 1348 363 1352
rect 615 1348 619 1352
rect 871 1348 875 1352
rect 1127 1348 1131 1352
rect 1391 1348 1395 1352
rect 1935 1347 1939 1351
rect 3839 1351 3843 1355
rect 3887 1352 3891 1356
rect 4023 1352 4027 1356
rect 4175 1352 4179 1356
rect 4383 1352 4387 1356
rect 4623 1352 4627 1356
rect 4895 1352 4899 1356
rect 5191 1352 5195 1356
rect 5487 1352 5491 1356
rect 5663 1351 5667 1355
rect 111 1289 115 1293
rect 367 1288 371 1292
rect 551 1288 555 1292
rect 727 1288 731 1292
rect 895 1288 899 1292
rect 1063 1288 1067 1292
rect 1223 1288 1227 1292
rect 1375 1288 1379 1292
rect 1527 1288 1531 1292
rect 1679 1288 1683 1292
rect 1815 1288 1819 1292
rect 1935 1289 1939 1293
rect 3839 1289 3843 1293
rect 3887 1288 3891 1292
rect 4047 1288 4051 1292
rect 4239 1288 4243 1292
rect 4455 1288 4459 1292
rect 4695 1288 4699 1292
rect 4951 1288 4955 1292
rect 5223 1288 5227 1292
rect 5495 1288 5499 1292
rect 5663 1289 5667 1293
rect 111 1272 115 1276
rect 339 1273 343 1277
rect 523 1273 527 1277
rect 699 1273 703 1277
rect 867 1273 871 1277
rect 1035 1273 1039 1277
rect 1195 1273 1199 1277
rect 1347 1273 1351 1277
rect 1499 1273 1503 1277
rect 1651 1273 1655 1277
rect 1787 1273 1791 1277
rect 1935 1272 1939 1276
rect 3839 1272 3843 1276
rect 3859 1273 3863 1277
rect 4019 1273 4023 1277
rect 4211 1273 4215 1277
rect 4427 1273 4431 1277
rect 4667 1273 4671 1277
rect 4923 1273 4927 1277
rect 5195 1273 5199 1277
rect 5467 1273 5471 1277
rect 5663 1272 5667 1276
rect 1975 1232 1979 1236
rect 3091 1231 3095 1235
rect 3227 1231 3231 1235
rect 3363 1231 3367 1235
rect 3799 1232 3803 1236
rect 1975 1215 1979 1219
rect 3119 1216 3123 1220
rect 3255 1216 3259 1220
rect 3391 1216 3395 1220
rect 3799 1215 3803 1219
rect 1975 1157 1979 1161
rect 2983 1156 2987 1160
rect 3119 1156 3123 1160
rect 3255 1156 3259 1160
rect 3799 1157 3803 1161
rect 1975 1140 1979 1144
rect 2955 1141 2959 1145
rect 3091 1141 3095 1145
rect 3227 1141 3231 1145
rect 3799 1140 3803 1144
rect 111 1128 115 1132
rect 235 1127 239 1131
rect 379 1127 383 1131
rect 523 1127 527 1131
rect 667 1127 671 1131
rect 811 1127 815 1131
rect 947 1127 951 1131
rect 1091 1127 1095 1131
rect 1235 1127 1239 1131
rect 1379 1127 1383 1131
rect 1515 1127 1519 1131
rect 1651 1127 1655 1131
rect 1787 1127 1791 1131
rect 1935 1128 1939 1132
rect 3839 1132 3843 1136
rect 3859 1131 3863 1135
rect 4091 1131 4095 1135
rect 4339 1131 4343 1135
rect 4579 1131 4583 1135
rect 4811 1131 4815 1135
rect 5043 1131 5047 1135
rect 5275 1131 5279 1135
rect 5515 1131 5519 1135
rect 5663 1132 5667 1136
rect 111 1111 115 1115
rect 263 1112 267 1116
rect 407 1112 411 1116
rect 551 1112 555 1116
rect 695 1112 699 1116
rect 839 1112 843 1116
rect 975 1112 979 1116
rect 1119 1112 1123 1116
rect 1263 1112 1267 1116
rect 1407 1112 1411 1116
rect 1543 1112 1547 1116
rect 1679 1112 1683 1116
rect 1815 1112 1819 1116
rect 1935 1111 1939 1115
rect 3839 1115 3843 1119
rect 3887 1116 3891 1120
rect 4119 1116 4123 1120
rect 4367 1116 4371 1120
rect 4607 1116 4611 1120
rect 4839 1116 4843 1120
rect 5071 1116 5075 1120
rect 5303 1116 5307 1120
rect 5543 1116 5547 1120
rect 5663 1115 5667 1119
rect 111 1041 115 1045
rect 263 1040 267 1044
rect 463 1040 467 1044
rect 663 1040 667 1044
rect 871 1040 875 1044
rect 1079 1040 1083 1044
rect 1935 1041 1939 1045
rect 3839 1037 3843 1041
rect 4863 1036 4867 1040
rect 4999 1036 5003 1040
rect 5135 1036 5139 1040
rect 5271 1036 5275 1040
rect 5407 1036 5411 1040
rect 5543 1036 5547 1040
rect 5663 1037 5667 1041
rect 111 1024 115 1028
rect 235 1025 239 1029
rect 435 1025 439 1029
rect 635 1025 639 1029
rect 843 1025 847 1029
rect 1051 1025 1055 1029
rect 1935 1024 1939 1028
rect 3839 1020 3843 1024
rect 4835 1021 4839 1025
rect 4971 1021 4975 1025
rect 5107 1021 5111 1025
rect 5243 1021 5247 1025
rect 5379 1021 5383 1025
rect 5515 1021 5519 1025
rect 5663 1020 5667 1024
rect 1975 1008 1979 1012
rect 1995 1007 1999 1011
rect 2131 1007 2135 1011
rect 2275 1007 2279 1011
rect 2443 1007 2447 1011
rect 2627 1007 2631 1011
rect 2819 1007 2823 1011
rect 3027 1007 3031 1011
rect 3235 1007 3239 1011
rect 3451 1007 3455 1011
rect 3651 1007 3655 1011
rect 3799 1008 3803 1012
rect 1975 991 1979 995
rect 2023 992 2027 996
rect 2159 992 2163 996
rect 2303 992 2307 996
rect 2471 992 2475 996
rect 2655 992 2659 996
rect 2847 992 2851 996
rect 3055 992 3059 996
rect 3263 992 3267 996
rect 3479 992 3483 996
rect 3679 992 3683 996
rect 3799 991 3803 995
rect 1975 933 1979 937
rect 2095 932 2099 936
rect 2231 932 2235 936
rect 2367 932 2371 936
rect 2503 932 2507 936
rect 2655 932 2659 936
rect 2831 932 2835 936
rect 3023 932 3027 936
rect 3231 932 3235 936
rect 3455 932 3459 936
rect 3679 932 3683 936
rect 3799 933 3803 937
rect 1975 916 1979 920
rect 2067 917 2071 921
rect 2203 917 2207 921
rect 2339 917 2343 921
rect 2475 917 2479 921
rect 2627 917 2631 921
rect 2803 917 2807 921
rect 2995 917 2999 921
rect 3203 917 3207 921
rect 3427 917 3431 921
rect 3651 917 3655 921
rect 3799 916 3803 920
rect 111 880 115 884
rect 195 879 199 883
rect 371 879 375 883
rect 547 879 551 883
rect 723 879 727 883
rect 907 879 911 883
rect 1091 879 1095 883
rect 1935 880 1939 884
rect 3839 876 3843 880
rect 4587 875 4591 879
rect 4755 875 4759 879
rect 4939 875 4943 879
rect 5131 875 5135 879
rect 5331 875 5335 879
rect 5515 875 5519 879
rect 5663 876 5667 880
rect 111 863 115 867
rect 223 864 227 868
rect 399 864 403 868
rect 575 864 579 868
rect 751 864 755 868
rect 935 864 939 868
rect 1119 864 1123 868
rect 1935 863 1939 867
rect 3839 859 3843 863
rect 4615 860 4619 864
rect 4783 860 4787 864
rect 4967 860 4971 864
rect 5159 860 5163 864
rect 5359 860 5363 864
rect 5543 860 5547 864
rect 5663 859 5667 863
rect 111 789 115 793
rect 159 788 163 792
rect 351 788 355 792
rect 583 788 587 792
rect 839 788 843 792
rect 1111 788 1115 792
rect 1399 788 1403 792
rect 1687 788 1691 792
rect 1935 789 1939 793
rect 3839 793 3843 797
rect 3983 792 3987 796
rect 4239 792 4243 796
rect 4535 792 4539 796
rect 4863 792 4867 796
rect 5215 792 5219 796
rect 5543 792 5547 796
rect 5663 793 5667 797
rect 1975 784 1979 788
rect 2307 783 2311 787
rect 2483 783 2487 787
rect 2659 783 2663 787
rect 2827 783 2831 787
rect 2995 783 2999 787
rect 3163 783 3167 787
rect 3331 783 3335 787
rect 3499 783 3503 787
rect 3651 783 3655 787
rect 3799 784 3803 788
rect 111 772 115 776
rect 131 773 135 777
rect 323 773 327 777
rect 555 773 559 777
rect 811 773 815 777
rect 1083 773 1087 777
rect 1371 773 1375 777
rect 1659 773 1663 777
rect 1935 772 1939 776
rect 3839 776 3843 780
rect 3955 777 3959 781
rect 4211 777 4215 781
rect 4507 777 4511 781
rect 4835 777 4839 781
rect 5187 777 5191 781
rect 5515 777 5519 781
rect 5663 776 5667 780
rect 1975 767 1979 771
rect 2335 768 2339 772
rect 2511 768 2515 772
rect 2687 768 2691 772
rect 2855 768 2859 772
rect 3023 768 3027 772
rect 3191 768 3195 772
rect 3359 768 3363 772
rect 3527 768 3531 772
rect 3679 768 3683 772
rect 3799 767 3803 771
rect 1975 705 1979 709
rect 3135 704 3139 708
rect 3271 704 3275 708
rect 3407 704 3411 708
rect 3543 704 3547 708
rect 3679 704 3683 708
rect 3799 705 3803 709
rect 1975 688 1979 692
rect 3107 689 3111 693
rect 3243 689 3247 693
rect 3379 689 3383 693
rect 3515 689 3519 693
rect 3651 689 3655 693
rect 3799 688 3803 692
rect 111 640 115 644
rect 131 639 135 643
rect 291 639 295 643
rect 483 639 487 643
rect 675 639 679 643
rect 867 639 871 643
rect 1059 639 1063 643
rect 1251 639 1255 643
rect 1435 639 1439 643
rect 1619 639 1623 643
rect 1787 639 1791 643
rect 1935 640 1939 644
rect 111 623 115 627
rect 159 624 163 628
rect 319 624 323 628
rect 511 624 515 628
rect 703 624 707 628
rect 895 624 899 628
rect 1087 624 1091 628
rect 1279 624 1283 628
rect 1463 624 1467 628
rect 1647 624 1651 628
rect 1815 624 1819 628
rect 1935 623 1939 627
rect 3839 620 3843 624
rect 3859 619 3863 623
rect 3995 619 3999 623
rect 4139 619 4143 623
rect 4323 619 4327 623
rect 4531 619 4535 623
rect 4755 619 4759 623
rect 4995 619 4999 623
rect 5243 619 5247 623
rect 5499 619 5503 623
rect 5663 620 5667 624
rect 3839 603 3843 607
rect 3887 604 3891 608
rect 4023 604 4027 608
rect 4167 604 4171 608
rect 4351 604 4355 608
rect 4559 604 4563 608
rect 4783 604 4787 608
rect 5023 604 5027 608
rect 5271 604 5275 608
rect 5527 604 5531 608
rect 5663 603 5667 607
rect 111 565 115 569
rect 159 564 163 568
rect 327 564 331 568
rect 519 564 523 568
rect 711 564 715 568
rect 903 564 907 568
rect 1095 564 1099 568
rect 1279 564 1283 568
rect 1463 564 1467 568
rect 1647 564 1651 568
rect 1815 564 1819 568
rect 1935 565 1939 569
rect 111 548 115 552
rect 131 549 135 553
rect 299 549 303 553
rect 491 549 495 553
rect 683 549 687 553
rect 875 549 879 553
rect 1067 549 1071 553
rect 1251 549 1255 553
rect 1435 549 1439 553
rect 1619 549 1623 553
rect 1787 549 1791 553
rect 1935 548 1939 552
rect 3839 545 3843 549
rect 3887 544 3891 548
rect 4023 544 4027 548
rect 4159 544 4163 548
rect 4295 544 4299 548
rect 4431 544 4435 548
rect 4575 544 4579 548
rect 4743 544 4747 548
rect 4927 544 4931 548
rect 5119 544 5123 548
rect 5319 544 5323 548
rect 5527 544 5531 548
rect 5663 545 5667 549
rect 3839 528 3843 532
rect 3859 529 3863 533
rect 3995 529 3999 533
rect 4131 529 4135 533
rect 4267 529 4271 533
rect 4403 529 4407 533
rect 4547 529 4551 533
rect 4715 529 4719 533
rect 4899 529 4903 533
rect 5091 529 5095 533
rect 5291 529 5295 533
rect 5499 529 5503 533
rect 5663 528 5667 532
rect 111 416 115 420
rect 395 415 399 419
rect 587 415 591 419
rect 787 415 791 419
rect 987 415 991 419
rect 1195 415 1199 419
rect 1411 415 1415 419
rect 1935 416 1939 420
rect 111 399 115 403
rect 423 400 427 404
rect 615 400 619 404
rect 815 400 819 404
rect 1015 400 1019 404
rect 1223 400 1227 404
rect 1439 400 1443 404
rect 1935 399 1939 403
rect 1975 396 1979 400
rect 1995 395 1999 399
rect 2203 395 2207 399
rect 2427 395 2431 399
rect 2651 395 2655 399
rect 2867 395 2871 399
rect 3075 395 3079 399
rect 3275 395 3279 399
rect 3475 395 3479 399
rect 3651 395 3655 399
rect 3799 396 3803 400
rect 3839 396 3843 400
rect 4379 395 4383 399
rect 4595 395 4599 399
rect 4819 395 4823 399
rect 5051 395 5055 399
rect 5283 395 5287 399
rect 5663 396 5667 400
rect 1975 379 1979 383
rect 2023 380 2027 384
rect 2231 380 2235 384
rect 2455 380 2459 384
rect 2679 380 2683 384
rect 2895 380 2899 384
rect 3103 380 3107 384
rect 3303 380 3307 384
rect 3503 380 3507 384
rect 3679 380 3683 384
rect 3799 379 3803 383
rect 3839 379 3843 383
rect 4407 380 4411 384
rect 4623 380 4627 384
rect 4847 380 4851 384
rect 5079 380 5083 384
rect 5311 380 5315 384
rect 5663 379 5667 383
rect 111 329 115 333
rect 647 328 651 332
rect 815 328 819 332
rect 991 328 995 332
rect 1167 328 1171 332
rect 1343 328 1347 332
rect 1935 329 1939 333
rect 3839 321 3843 325
rect 4639 320 4643 324
rect 4807 320 4811 324
rect 4983 320 4987 324
rect 5167 320 5171 324
rect 5359 320 5363 324
rect 5543 320 5547 324
rect 5663 321 5667 325
rect 111 312 115 316
rect 619 313 623 317
rect 787 313 791 317
rect 963 313 967 317
rect 1139 313 1143 317
rect 1315 313 1319 317
rect 1935 312 1939 316
rect 1975 305 1979 309
rect 2023 304 2027 308
rect 2159 304 2163 308
rect 2295 304 2299 308
rect 2431 304 2435 308
rect 2567 304 2571 308
rect 2703 304 2707 308
rect 2839 304 2843 308
rect 2975 304 2979 308
rect 3111 304 3115 308
rect 3247 304 3251 308
rect 3383 304 3387 308
rect 3519 304 3523 308
rect 3655 304 3659 308
rect 3799 305 3803 309
rect 3839 304 3843 308
rect 4611 305 4615 309
rect 4779 305 4783 309
rect 4955 305 4959 309
rect 5139 305 5143 309
rect 5331 305 5335 309
rect 5515 305 5519 309
rect 5663 304 5667 308
rect 1975 288 1979 292
rect 1995 289 1999 293
rect 2131 289 2135 293
rect 2267 289 2271 293
rect 2403 289 2407 293
rect 2539 289 2543 293
rect 2675 289 2679 293
rect 2811 289 2815 293
rect 2947 289 2951 293
rect 3083 289 3087 293
rect 3219 289 3223 293
rect 3355 289 3359 293
rect 3491 289 3495 293
rect 3627 289 3631 293
rect 3799 288 3803 292
rect 111 140 115 144
rect 539 139 543 143
rect 675 139 679 143
rect 811 139 815 143
rect 947 139 951 143
rect 1083 139 1087 143
rect 1219 139 1223 143
rect 1355 139 1359 143
rect 1491 139 1495 143
rect 1935 140 1939 144
rect 3839 144 3843 148
rect 4291 143 4295 147
rect 4427 143 4431 147
rect 4563 143 4567 147
rect 4699 143 4703 147
rect 4835 143 4839 147
rect 4971 143 4975 147
rect 5107 143 5111 147
rect 5243 143 5247 147
rect 5379 143 5383 147
rect 5515 143 5519 147
rect 5663 144 5667 148
rect 111 123 115 127
rect 567 124 571 128
rect 703 124 707 128
rect 839 124 843 128
rect 975 124 979 128
rect 1111 124 1115 128
rect 1247 124 1251 128
rect 1383 124 1387 128
rect 1519 124 1523 128
rect 1935 123 1939 127
rect 3839 127 3843 131
rect 4319 128 4323 132
rect 4455 128 4459 132
rect 4591 128 4595 132
rect 4727 128 4731 132
rect 4863 128 4867 132
rect 4999 128 5003 132
rect 5135 128 5139 132
rect 5271 128 5275 132
rect 5407 128 5411 132
rect 5543 128 5547 132
rect 5663 127 5667 131
rect 1975 120 1979 124
rect 1995 119 1999 123
rect 2131 119 2135 123
rect 2267 119 2271 123
rect 2403 119 2407 123
rect 2539 119 2543 123
rect 2675 119 2679 123
rect 2811 119 2815 123
rect 2947 119 2951 123
rect 3083 119 3087 123
rect 3219 119 3223 123
rect 3355 119 3359 123
rect 3491 119 3495 123
rect 3627 119 3631 123
rect 3799 120 3803 124
rect 1975 103 1979 107
rect 2023 104 2027 108
rect 2159 104 2163 108
rect 2295 104 2299 108
rect 2431 104 2435 108
rect 2567 104 2571 108
rect 2703 104 2707 108
rect 2839 104 2843 108
rect 2975 104 2979 108
rect 3111 104 3115 108
rect 3247 104 3251 108
rect 3383 104 3387 108
rect 3519 104 3523 108
rect 3655 104 3659 108
rect 3799 103 3803 107
<< m3 >>
rect 111 5722 115 5723
rect 111 5717 115 5718
rect 159 5722 163 5723
rect 159 5717 163 5718
rect 303 5722 307 5723
rect 303 5717 307 5718
rect 503 5722 507 5723
rect 503 5717 507 5718
rect 727 5722 731 5723
rect 727 5717 731 5718
rect 983 5722 987 5723
rect 983 5717 987 5718
rect 1255 5722 1259 5723
rect 1255 5717 1259 5718
rect 1543 5722 1547 5723
rect 1543 5717 1547 5718
rect 1815 5722 1819 5723
rect 1815 5717 1819 5718
rect 1935 5722 1939 5723
rect 1935 5717 1939 5718
rect 112 5694 114 5717
rect 110 5693 116 5694
rect 160 5693 162 5717
rect 304 5693 306 5717
rect 504 5693 506 5717
rect 728 5693 730 5717
rect 984 5693 986 5717
rect 1256 5693 1258 5717
rect 1544 5693 1546 5717
rect 1816 5693 1818 5717
rect 1936 5694 1938 5717
rect 1975 5694 1979 5695
rect 1934 5693 1940 5694
rect 110 5689 111 5693
rect 115 5689 116 5693
rect 110 5688 116 5689
rect 158 5692 164 5693
rect 158 5688 159 5692
rect 163 5688 164 5692
rect 158 5687 164 5688
rect 302 5692 308 5693
rect 302 5688 303 5692
rect 307 5688 308 5692
rect 302 5687 308 5688
rect 502 5692 508 5693
rect 502 5688 503 5692
rect 507 5688 508 5692
rect 502 5687 508 5688
rect 726 5692 732 5693
rect 726 5688 727 5692
rect 731 5688 732 5692
rect 726 5687 732 5688
rect 982 5692 988 5693
rect 982 5688 983 5692
rect 987 5688 988 5692
rect 982 5687 988 5688
rect 1254 5692 1260 5693
rect 1254 5688 1255 5692
rect 1259 5688 1260 5692
rect 1254 5687 1260 5688
rect 1542 5692 1548 5693
rect 1542 5688 1543 5692
rect 1547 5688 1548 5692
rect 1542 5687 1548 5688
rect 1814 5692 1820 5693
rect 1814 5688 1815 5692
rect 1819 5688 1820 5692
rect 1934 5689 1935 5693
rect 1939 5689 1940 5693
rect 1975 5689 1979 5690
rect 1995 5694 1999 5695
rect 1995 5689 1999 5690
rect 2179 5694 2183 5695
rect 2179 5689 2183 5690
rect 2387 5694 2391 5695
rect 2387 5689 2391 5690
rect 2587 5694 2591 5695
rect 2587 5689 2591 5690
rect 2779 5694 2783 5695
rect 2779 5689 2783 5690
rect 2963 5694 2967 5695
rect 2963 5689 2967 5690
rect 3147 5694 3151 5695
rect 3147 5689 3151 5690
rect 3323 5694 3327 5695
rect 3323 5689 3327 5690
rect 3499 5694 3503 5695
rect 3499 5689 3503 5690
rect 3651 5694 3655 5695
rect 3651 5689 3655 5690
rect 3799 5694 3803 5695
rect 3799 5689 3803 5690
rect 1934 5688 1940 5689
rect 1814 5687 1820 5688
rect 130 5677 136 5678
rect 110 5676 116 5677
rect 110 5672 111 5676
rect 115 5672 116 5676
rect 130 5673 131 5677
rect 135 5673 136 5677
rect 130 5672 136 5673
rect 274 5677 280 5678
rect 274 5673 275 5677
rect 279 5673 280 5677
rect 274 5672 280 5673
rect 474 5677 480 5678
rect 474 5673 475 5677
rect 479 5673 480 5677
rect 474 5672 480 5673
rect 698 5677 704 5678
rect 698 5673 699 5677
rect 703 5673 704 5677
rect 698 5672 704 5673
rect 954 5677 960 5678
rect 954 5673 955 5677
rect 959 5673 960 5677
rect 954 5672 960 5673
rect 1226 5677 1232 5678
rect 1226 5673 1227 5677
rect 1231 5673 1232 5677
rect 1226 5672 1232 5673
rect 1514 5677 1520 5678
rect 1514 5673 1515 5677
rect 1519 5673 1520 5677
rect 1514 5672 1520 5673
rect 1786 5677 1792 5678
rect 1786 5673 1787 5677
rect 1791 5673 1792 5677
rect 1786 5672 1792 5673
rect 1934 5676 1940 5677
rect 1934 5672 1935 5676
rect 1939 5672 1940 5676
rect 110 5671 116 5672
rect 112 5607 114 5671
rect 132 5607 134 5672
rect 276 5607 278 5672
rect 476 5607 478 5672
rect 700 5607 702 5672
rect 956 5607 958 5672
rect 1228 5607 1230 5672
rect 1516 5607 1518 5672
rect 1788 5607 1790 5672
rect 1934 5671 1940 5672
rect 1936 5607 1938 5671
rect 1976 5629 1978 5689
rect 1974 5628 1980 5629
rect 1996 5628 1998 5689
rect 2180 5628 2182 5689
rect 2388 5628 2390 5689
rect 2588 5628 2590 5689
rect 2780 5628 2782 5689
rect 2964 5628 2966 5689
rect 3148 5628 3150 5689
rect 3324 5628 3326 5689
rect 3500 5628 3502 5689
rect 3652 5628 3654 5689
rect 3800 5629 3802 5689
rect 3839 5650 3843 5651
rect 3839 5645 3843 5646
rect 4291 5650 4295 5651
rect 4291 5645 4295 5646
rect 4427 5650 4431 5651
rect 4427 5645 4431 5646
rect 4563 5650 4567 5651
rect 4563 5645 4567 5646
rect 4699 5650 4703 5651
rect 4699 5645 4703 5646
rect 4835 5650 4839 5651
rect 4835 5645 4839 5646
rect 4971 5650 4975 5651
rect 4971 5645 4975 5646
rect 5107 5650 5111 5651
rect 5107 5645 5111 5646
rect 5663 5650 5667 5651
rect 5663 5645 5667 5646
rect 3798 5628 3804 5629
rect 1974 5624 1975 5628
rect 1979 5624 1980 5628
rect 1974 5623 1980 5624
rect 1994 5627 2000 5628
rect 1994 5623 1995 5627
rect 1999 5623 2000 5627
rect 1994 5622 2000 5623
rect 2178 5627 2184 5628
rect 2178 5623 2179 5627
rect 2183 5623 2184 5627
rect 2178 5622 2184 5623
rect 2386 5627 2392 5628
rect 2386 5623 2387 5627
rect 2391 5623 2392 5627
rect 2386 5622 2392 5623
rect 2586 5627 2592 5628
rect 2586 5623 2587 5627
rect 2591 5623 2592 5627
rect 2586 5622 2592 5623
rect 2778 5627 2784 5628
rect 2778 5623 2779 5627
rect 2783 5623 2784 5627
rect 2778 5622 2784 5623
rect 2962 5627 2968 5628
rect 2962 5623 2963 5627
rect 2967 5623 2968 5627
rect 2962 5622 2968 5623
rect 3146 5627 3152 5628
rect 3146 5623 3147 5627
rect 3151 5623 3152 5627
rect 3146 5622 3152 5623
rect 3322 5627 3328 5628
rect 3322 5623 3323 5627
rect 3327 5623 3328 5627
rect 3322 5622 3328 5623
rect 3498 5627 3504 5628
rect 3498 5623 3499 5627
rect 3503 5623 3504 5627
rect 3498 5622 3504 5623
rect 3650 5627 3656 5628
rect 3650 5623 3651 5627
rect 3655 5623 3656 5627
rect 3798 5624 3799 5628
rect 3803 5624 3804 5628
rect 3798 5623 3804 5624
rect 3650 5622 3656 5623
rect 2022 5612 2028 5613
rect 1974 5611 1980 5612
rect 1974 5607 1975 5611
rect 1979 5607 1980 5611
rect 2022 5608 2023 5612
rect 2027 5608 2028 5612
rect 2022 5607 2028 5608
rect 2206 5612 2212 5613
rect 2206 5608 2207 5612
rect 2211 5608 2212 5612
rect 2206 5607 2212 5608
rect 2414 5612 2420 5613
rect 2414 5608 2415 5612
rect 2419 5608 2420 5612
rect 2414 5607 2420 5608
rect 2614 5612 2620 5613
rect 2614 5608 2615 5612
rect 2619 5608 2620 5612
rect 2614 5607 2620 5608
rect 2806 5612 2812 5613
rect 2806 5608 2807 5612
rect 2811 5608 2812 5612
rect 2806 5607 2812 5608
rect 2990 5612 2996 5613
rect 2990 5608 2991 5612
rect 2995 5608 2996 5612
rect 2990 5607 2996 5608
rect 3174 5612 3180 5613
rect 3174 5608 3175 5612
rect 3179 5608 3180 5612
rect 3174 5607 3180 5608
rect 3350 5612 3356 5613
rect 3350 5608 3351 5612
rect 3355 5608 3356 5612
rect 3350 5607 3356 5608
rect 3526 5612 3532 5613
rect 3526 5608 3527 5612
rect 3531 5608 3532 5612
rect 3526 5607 3532 5608
rect 3678 5612 3684 5613
rect 3678 5608 3679 5612
rect 3683 5608 3684 5612
rect 3678 5607 3684 5608
rect 3798 5611 3804 5612
rect 3798 5607 3799 5611
rect 3803 5607 3804 5611
rect 111 5606 115 5607
rect 111 5601 115 5602
rect 131 5606 135 5607
rect 131 5601 135 5602
rect 275 5606 279 5607
rect 275 5601 279 5602
rect 475 5606 479 5607
rect 475 5601 479 5602
rect 563 5606 567 5607
rect 563 5601 567 5602
rect 699 5606 703 5607
rect 699 5601 703 5602
rect 723 5606 727 5607
rect 723 5601 727 5602
rect 883 5606 887 5607
rect 883 5601 887 5602
rect 955 5606 959 5607
rect 955 5601 959 5602
rect 1051 5606 1055 5607
rect 1051 5601 1055 5602
rect 1227 5606 1231 5607
rect 1227 5601 1231 5602
rect 1403 5606 1407 5607
rect 1403 5601 1407 5602
rect 1515 5606 1519 5607
rect 1515 5601 1519 5602
rect 1579 5606 1583 5607
rect 1579 5601 1583 5602
rect 1763 5606 1767 5607
rect 1763 5601 1767 5602
rect 1787 5606 1791 5607
rect 1787 5601 1791 5602
rect 1935 5606 1939 5607
rect 1974 5606 1980 5607
rect 1935 5601 1939 5602
rect 112 5541 114 5601
rect 110 5540 116 5541
rect 564 5540 566 5601
rect 724 5540 726 5601
rect 884 5540 886 5601
rect 1052 5540 1054 5601
rect 1228 5540 1230 5601
rect 1404 5540 1406 5601
rect 1580 5540 1582 5601
rect 1764 5540 1766 5601
rect 1936 5541 1938 5601
rect 1976 5583 1978 5606
rect 2024 5583 2026 5607
rect 2208 5583 2210 5607
rect 2416 5583 2418 5607
rect 2616 5583 2618 5607
rect 2808 5583 2810 5607
rect 2992 5583 2994 5607
rect 3176 5583 3178 5607
rect 3352 5583 3354 5607
rect 3528 5583 3530 5607
rect 3680 5583 3682 5607
rect 3798 5606 3804 5607
rect 3800 5583 3802 5606
rect 3840 5585 3842 5645
rect 3838 5584 3844 5585
rect 4292 5584 4294 5645
rect 4428 5584 4430 5645
rect 4564 5584 4566 5645
rect 4700 5584 4702 5645
rect 4836 5584 4838 5645
rect 4972 5584 4974 5645
rect 5108 5584 5110 5645
rect 5664 5585 5666 5645
rect 5662 5584 5668 5585
rect 1975 5582 1979 5583
rect 1975 5577 1979 5578
rect 2023 5582 2027 5583
rect 2023 5577 2027 5578
rect 2207 5582 2211 5583
rect 2207 5577 2211 5578
rect 2263 5582 2267 5583
rect 2263 5577 2267 5578
rect 2415 5582 2419 5583
rect 2415 5577 2419 5578
rect 2503 5582 2507 5583
rect 2503 5577 2507 5578
rect 2615 5582 2619 5583
rect 2615 5577 2619 5578
rect 2743 5582 2747 5583
rect 2743 5577 2747 5578
rect 2807 5582 2811 5583
rect 2807 5577 2811 5578
rect 2983 5582 2987 5583
rect 2983 5577 2987 5578
rect 2991 5582 2995 5583
rect 2991 5577 2995 5578
rect 3175 5582 3179 5583
rect 3175 5577 3179 5578
rect 3223 5582 3227 5583
rect 3223 5577 3227 5578
rect 3351 5582 3355 5583
rect 3351 5577 3355 5578
rect 3463 5582 3467 5583
rect 3463 5577 3467 5578
rect 3527 5582 3531 5583
rect 3527 5577 3531 5578
rect 3679 5582 3683 5583
rect 3679 5577 3683 5578
rect 3799 5582 3803 5583
rect 3838 5580 3839 5584
rect 3843 5580 3844 5584
rect 3838 5579 3844 5580
rect 4290 5583 4296 5584
rect 4290 5579 4291 5583
rect 4295 5579 4296 5583
rect 4290 5578 4296 5579
rect 4426 5583 4432 5584
rect 4426 5579 4427 5583
rect 4431 5579 4432 5583
rect 4426 5578 4432 5579
rect 4562 5583 4568 5584
rect 4562 5579 4563 5583
rect 4567 5579 4568 5583
rect 4562 5578 4568 5579
rect 4698 5583 4704 5584
rect 4698 5579 4699 5583
rect 4703 5579 4704 5583
rect 4698 5578 4704 5579
rect 4834 5583 4840 5584
rect 4834 5579 4835 5583
rect 4839 5579 4840 5583
rect 4834 5578 4840 5579
rect 4970 5583 4976 5584
rect 4970 5579 4971 5583
rect 4975 5579 4976 5583
rect 4970 5578 4976 5579
rect 5106 5583 5112 5584
rect 5106 5579 5107 5583
rect 5111 5579 5112 5583
rect 5662 5580 5663 5584
rect 5667 5580 5668 5584
rect 5662 5579 5668 5580
rect 5106 5578 5112 5579
rect 3799 5577 3803 5578
rect 1976 5554 1978 5577
rect 1974 5553 1980 5554
rect 2264 5553 2266 5577
rect 2504 5553 2506 5577
rect 2744 5553 2746 5577
rect 2984 5553 2986 5577
rect 3224 5553 3226 5577
rect 3464 5553 3466 5577
rect 3680 5553 3682 5577
rect 3800 5554 3802 5577
rect 4318 5568 4324 5569
rect 3838 5567 3844 5568
rect 3838 5563 3839 5567
rect 3843 5563 3844 5567
rect 4318 5564 4319 5568
rect 4323 5564 4324 5568
rect 4318 5563 4324 5564
rect 4454 5568 4460 5569
rect 4454 5564 4455 5568
rect 4459 5564 4460 5568
rect 4454 5563 4460 5564
rect 4590 5568 4596 5569
rect 4590 5564 4591 5568
rect 4595 5564 4596 5568
rect 4590 5563 4596 5564
rect 4726 5568 4732 5569
rect 4726 5564 4727 5568
rect 4731 5564 4732 5568
rect 4726 5563 4732 5564
rect 4862 5568 4868 5569
rect 4862 5564 4863 5568
rect 4867 5564 4868 5568
rect 4862 5563 4868 5564
rect 4998 5568 5004 5569
rect 4998 5564 4999 5568
rect 5003 5564 5004 5568
rect 4998 5563 5004 5564
rect 5134 5568 5140 5569
rect 5134 5564 5135 5568
rect 5139 5564 5140 5568
rect 5134 5563 5140 5564
rect 5662 5567 5668 5568
rect 5662 5563 5663 5567
rect 5667 5563 5668 5567
rect 3838 5562 3844 5563
rect 3798 5553 3804 5554
rect 1974 5549 1975 5553
rect 1979 5549 1980 5553
rect 1974 5548 1980 5549
rect 2262 5552 2268 5553
rect 2262 5548 2263 5552
rect 2267 5548 2268 5552
rect 2262 5547 2268 5548
rect 2502 5552 2508 5553
rect 2502 5548 2503 5552
rect 2507 5548 2508 5552
rect 2502 5547 2508 5548
rect 2742 5552 2748 5553
rect 2742 5548 2743 5552
rect 2747 5548 2748 5552
rect 2742 5547 2748 5548
rect 2982 5552 2988 5553
rect 2982 5548 2983 5552
rect 2987 5548 2988 5552
rect 2982 5547 2988 5548
rect 3222 5552 3228 5553
rect 3222 5548 3223 5552
rect 3227 5548 3228 5552
rect 3222 5547 3228 5548
rect 3462 5552 3468 5553
rect 3462 5548 3463 5552
rect 3467 5548 3468 5552
rect 3462 5547 3468 5548
rect 3678 5552 3684 5553
rect 3678 5548 3679 5552
rect 3683 5548 3684 5552
rect 3798 5549 3799 5553
rect 3803 5549 3804 5553
rect 3798 5548 3804 5549
rect 3678 5547 3684 5548
rect 1934 5540 1940 5541
rect 110 5536 111 5540
rect 115 5536 116 5540
rect 110 5535 116 5536
rect 562 5539 568 5540
rect 562 5535 563 5539
rect 567 5535 568 5539
rect 562 5534 568 5535
rect 722 5539 728 5540
rect 722 5535 723 5539
rect 727 5535 728 5539
rect 722 5534 728 5535
rect 882 5539 888 5540
rect 882 5535 883 5539
rect 887 5535 888 5539
rect 882 5534 888 5535
rect 1050 5539 1056 5540
rect 1050 5535 1051 5539
rect 1055 5535 1056 5539
rect 1050 5534 1056 5535
rect 1226 5539 1232 5540
rect 1226 5535 1227 5539
rect 1231 5535 1232 5539
rect 1226 5534 1232 5535
rect 1402 5539 1408 5540
rect 1402 5535 1403 5539
rect 1407 5535 1408 5539
rect 1402 5534 1408 5535
rect 1578 5539 1584 5540
rect 1578 5535 1579 5539
rect 1583 5535 1584 5539
rect 1578 5534 1584 5535
rect 1762 5539 1768 5540
rect 1762 5535 1763 5539
rect 1767 5535 1768 5539
rect 1934 5536 1935 5540
rect 1939 5536 1940 5540
rect 3840 5539 3842 5562
rect 4320 5539 4322 5563
rect 4456 5539 4458 5563
rect 4592 5539 4594 5563
rect 4728 5539 4730 5563
rect 4864 5539 4866 5563
rect 5000 5539 5002 5563
rect 5136 5539 5138 5563
rect 5662 5562 5668 5563
rect 5664 5539 5666 5562
rect 3839 5538 3843 5539
rect 2234 5537 2240 5538
rect 1934 5535 1940 5536
rect 1974 5536 1980 5537
rect 1762 5534 1768 5535
rect 1974 5532 1975 5536
rect 1979 5532 1980 5536
rect 2234 5533 2235 5537
rect 2239 5533 2240 5537
rect 2234 5532 2240 5533
rect 2474 5537 2480 5538
rect 2474 5533 2475 5537
rect 2479 5533 2480 5537
rect 2474 5532 2480 5533
rect 2714 5537 2720 5538
rect 2714 5533 2715 5537
rect 2719 5533 2720 5537
rect 2714 5532 2720 5533
rect 2954 5537 2960 5538
rect 2954 5533 2955 5537
rect 2959 5533 2960 5537
rect 2954 5532 2960 5533
rect 3194 5537 3200 5538
rect 3194 5533 3195 5537
rect 3199 5533 3200 5537
rect 3194 5532 3200 5533
rect 3434 5537 3440 5538
rect 3434 5533 3435 5537
rect 3439 5533 3440 5537
rect 3434 5532 3440 5533
rect 3650 5537 3656 5538
rect 3650 5533 3651 5537
rect 3655 5533 3656 5537
rect 3650 5532 3656 5533
rect 3798 5536 3804 5537
rect 3798 5532 3799 5536
rect 3803 5532 3804 5536
rect 3839 5533 3843 5534
rect 3887 5538 3891 5539
rect 3887 5533 3891 5534
rect 4127 5538 4131 5539
rect 4127 5533 4131 5534
rect 4319 5538 4323 5539
rect 4319 5533 4323 5534
rect 4375 5538 4379 5539
rect 4375 5533 4379 5534
rect 4455 5538 4459 5539
rect 4455 5533 4459 5534
rect 4591 5538 4595 5539
rect 4591 5533 4595 5534
rect 4615 5538 4619 5539
rect 4615 5533 4619 5534
rect 4727 5538 4731 5539
rect 4727 5533 4731 5534
rect 4847 5538 4851 5539
rect 4847 5533 4851 5534
rect 4863 5538 4867 5539
rect 4863 5533 4867 5534
rect 4999 5538 5003 5539
rect 4999 5533 5003 5534
rect 5079 5538 5083 5539
rect 5079 5533 5083 5534
rect 5135 5538 5139 5539
rect 5135 5533 5139 5534
rect 5311 5538 5315 5539
rect 5311 5533 5315 5534
rect 5663 5538 5667 5539
rect 5663 5533 5667 5534
rect 1974 5531 1980 5532
rect 590 5524 596 5525
rect 110 5523 116 5524
rect 110 5519 111 5523
rect 115 5519 116 5523
rect 590 5520 591 5524
rect 595 5520 596 5524
rect 590 5519 596 5520
rect 750 5524 756 5525
rect 750 5520 751 5524
rect 755 5520 756 5524
rect 750 5519 756 5520
rect 910 5524 916 5525
rect 910 5520 911 5524
rect 915 5520 916 5524
rect 910 5519 916 5520
rect 1078 5524 1084 5525
rect 1078 5520 1079 5524
rect 1083 5520 1084 5524
rect 1078 5519 1084 5520
rect 1254 5524 1260 5525
rect 1254 5520 1255 5524
rect 1259 5520 1260 5524
rect 1254 5519 1260 5520
rect 1430 5524 1436 5525
rect 1430 5520 1431 5524
rect 1435 5520 1436 5524
rect 1430 5519 1436 5520
rect 1606 5524 1612 5525
rect 1606 5520 1607 5524
rect 1611 5520 1612 5524
rect 1606 5519 1612 5520
rect 1790 5524 1796 5525
rect 1790 5520 1791 5524
rect 1795 5520 1796 5524
rect 1790 5519 1796 5520
rect 1934 5523 1940 5524
rect 1934 5519 1935 5523
rect 1939 5519 1940 5523
rect 110 5518 116 5519
rect 112 5483 114 5518
rect 592 5483 594 5519
rect 752 5483 754 5519
rect 912 5483 914 5519
rect 1080 5483 1082 5519
rect 1256 5483 1258 5519
rect 1432 5483 1434 5519
rect 1608 5483 1610 5519
rect 1792 5483 1794 5519
rect 1934 5518 1940 5519
rect 1936 5483 1938 5518
rect 111 5482 115 5483
rect 111 5477 115 5478
rect 591 5482 595 5483
rect 591 5477 595 5478
rect 727 5482 731 5483
rect 727 5477 731 5478
rect 751 5482 755 5483
rect 751 5477 755 5478
rect 863 5482 867 5483
rect 863 5477 867 5478
rect 911 5482 915 5483
rect 911 5477 915 5478
rect 999 5482 1003 5483
rect 999 5477 1003 5478
rect 1079 5482 1083 5483
rect 1079 5477 1083 5478
rect 1135 5482 1139 5483
rect 1135 5477 1139 5478
rect 1255 5482 1259 5483
rect 1255 5477 1259 5478
rect 1271 5482 1275 5483
rect 1271 5477 1275 5478
rect 1407 5482 1411 5483
rect 1407 5477 1411 5478
rect 1431 5482 1435 5483
rect 1431 5477 1435 5478
rect 1543 5482 1547 5483
rect 1543 5477 1547 5478
rect 1607 5482 1611 5483
rect 1607 5477 1611 5478
rect 1679 5482 1683 5483
rect 1679 5477 1683 5478
rect 1791 5482 1795 5483
rect 1791 5477 1795 5478
rect 1815 5482 1819 5483
rect 1815 5477 1819 5478
rect 1935 5482 1939 5483
rect 1935 5477 1939 5478
rect 112 5454 114 5477
rect 110 5453 116 5454
rect 592 5453 594 5477
rect 728 5453 730 5477
rect 864 5453 866 5477
rect 1000 5453 1002 5477
rect 1136 5453 1138 5477
rect 1272 5453 1274 5477
rect 1408 5453 1410 5477
rect 1544 5453 1546 5477
rect 1680 5453 1682 5477
rect 1816 5453 1818 5477
rect 1936 5454 1938 5477
rect 1976 5463 1978 5531
rect 2236 5463 2238 5532
rect 2476 5463 2478 5532
rect 2716 5463 2718 5532
rect 2956 5463 2958 5532
rect 3196 5463 3198 5532
rect 3436 5463 3438 5532
rect 3652 5463 3654 5532
rect 3798 5531 3804 5532
rect 3800 5463 3802 5531
rect 3840 5510 3842 5533
rect 3838 5509 3844 5510
rect 3888 5509 3890 5533
rect 4128 5509 4130 5533
rect 4376 5509 4378 5533
rect 4616 5509 4618 5533
rect 4848 5509 4850 5533
rect 5080 5509 5082 5533
rect 5312 5509 5314 5533
rect 5664 5510 5666 5533
rect 5662 5509 5668 5510
rect 3838 5505 3839 5509
rect 3843 5505 3844 5509
rect 3838 5504 3844 5505
rect 3886 5508 3892 5509
rect 3886 5504 3887 5508
rect 3891 5504 3892 5508
rect 3886 5503 3892 5504
rect 4126 5508 4132 5509
rect 4126 5504 4127 5508
rect 4131 5504 4132 5508
rect 4126 5503 4132 5504
rect 4374 5508 4380 5509
rect 4374 5504 4375 5508
rect 4379 5504 4380 5508
rect 4374 5503 4380 5504
rect 4614 5508 4620 5509
rect 4614 5504 4615 5508
rect 4619 5504 4620 5508
rect 4614 5503 4620 5504
rect 4846 5508 4852 5509
rect 4846 5504 4847 5508
rect 4851 5504 4852 5508
rect 4846 5503 4852 5504
rect 5078 5508 5084 5509
rect 5078 5504 5079 5508
rect 5083 5504 5084 5508
rect 5078 5503 5084 5504
rect 5310 5508 5316 5509
rect 5310 5504 5311 5508
rect 5315 5504 5316 5508
rect 5662 5505 5663 5509
rect 5667 5505 5668 5509
rect 5662 5504 5668 5505
rect 5310 5503 5316 5504
rect 3858 5493 3864 5494
rect 3838 5492 3844 5493
rect 3838 5488 3839 5492
rect 3843 5488 3844 5492
rect 3858 5489 3859 5493
rect 3863 5489 3864 5493
rect 3858 5488 3864 5489
rect 4098 5493 4104 5494
rect 4098 5489 4099 5493
rect 4103 5489 4104 5493
rect 4098 5488 4104 5489
rect 4346 5493 4352 5494
rect 4346 5489 4347 5493
rect 4351 5489 4352 5493
rect 4346 5488 4352 5489
rect 4586 5493 4592 5494
rect 4586 5489 4587 5493
rect 4591 5489 4592 5493
rect 4586 5488 4592 5489
rect 4818 5493 4824 5494
rect 4818 5489 4819 5493
rect 4823 5489 4824 5493
rect 4818 5488 4824 5489
rect 5050 5493 5056 5494
rect 5050 5489 5051 5493
rect 5055 5489 5056 5493
rect 5050 5488 5056 5489
rect 5282 5493 5288 5494
rect 5282 5489 5283 5493
rect 5287 5489 5288 5493
rect 5282 5488 5288 5489
rect 5662 5492 5668 5493
rect 5662 5488 5663 5492
rect 5667 5488 5668 5492
rect 3838 5487 3844 5488
rect 1975 5462 1979 5463
rect 1975 5457 1979 5458
rect 2235 5462 2239 5463
rect 2235 5457 2239 5458
rect 2427 5462 2431 5463
rect 2427 5457 2431 5458
rect 2475 5462 2479 5463
rect 2475 5457 2479 5458
rect 2643 5462 2647 5463
rect 2643 5457 2647 5458
rect 2715 5462 2719 5463
rect 2715 5457 2719 5458
rect 2859 5462 2863 5463
rect 2859 5457 2863 5458
rect 2955 5462 2959 5463
rect 2955 5457 2959 5458
rect 3075 5462 3079 5463
rect 3075 5457 3079 5458
rect 3195 5462 3199 5463
rect 3195 5457 3199 5458
rect 3291 5462 3295 5463
rect 3291 5457 3295 5458
rect 3435 5462 3439 5463
rect 3435 5457 3439 5458
rect 3651 5462 3655 5463
rect 3651 5457 3655 5458
rect 3799 5462 3803 5463
rect 3799 5457 3803 5458
rect 1934 5453 1940 5454
rect 110 5449 111 5453
rect 115 5449 116 5453
rect 110 5448 116 5449
rect 590 5452 596 5453
rect 590 5448 591 5452
rect 595 5448 596 5452
rect 590 5447 596 5448
rect 726 5452 732 5453
rect 726 5448 727 5452
rect 731 5448 732 5452
rect 726 5447 732 5448
rect 862 5452 868 5453
rect 862 5448 863 5452
rect 867 5448 868 5452
rect 862 5447 868 5448
rect 998 5452 1004 5453
rect 998 5448 999 5452
rect 1003 5448 1004 5452
rect 998 5447 1004 5448
rect 1134 5452 1140 5453
rect 1134 5448 1135 5452
rect 1139 5448 1140 5452
rect 1134 5447 1140 5448
rect 1270 5452 1276 5453
rect 1270 5448 1271 5452
rect 1275 5448 1276 5452
rect 1270 5447 1276 5448
rect 1406 5452 1412 5453
rect 1406 5448 1407 5452
rect 1411 5448 1412 5452
rect 1406 5447 1412 5448
rect 1542 5452 1548 5453
rect 1542 5448 1543 5452
rect 1547 5448 1548 5452
rect 1542 5447 1548 5448
rect 1678 5452 1684 5453
rect 1678 5448 1679 5452
rect 1683 5448 1684 5452
rect 1678 5447 1684 5448
rect 1814 5452 1820 5453
rect 1814 5448 1815 5452
rect 1819 5448 1820 5452
rect 1934 5449 1935 5453
rect 1939 5449 1940 5453
rect 1934 5448 1940 5449
rect 1814 5447 1820 5448
rect 562 5437 568 5438
rect 110 5436 116 5437
rect 110 5432 111 5436
rect 115 5432 116 5436
rect 562 5433 563 5437
rect 567 5433 568 5437
rect 562 5432 568 5433
rect 698 5437 704 5438
rect 698 5433 699 5437
rect 703 5433 704 5437
rect 698 5432 704 5433
rect 834 5437 840 5438
rect 834 5433 835 5437
rect 839 5433 840 5437
rect 834 5432 840 5433
rect 970 5437 976 5438
rect 970 5433 971 5437
rect 975 5433 976 5437
rect 970 5432 976 5433
rect 1106 5437 1112 5438
rect 1106 5433 1107 5437
rect 1111 5433 1112 5437
rect 1106 5432 1112 5433
rect 1242 5437 1248 5438
rect 1242 5433 1243 5437
rect 1247 5433 1248 5437
rect 1242 5432 1248 5433
rect 1378 5437 1384 5438
rect 1378 5433 1379 5437
rect 1383 5433 1384 5437
rect 1378 5432 1384 5433
rect 1514 5437 1520 5438
rect 1514 5433 1515 5437
rect 1519 5433 1520 5437
rect 1514 5432 1520 5433
rect 1650 5437 1656 5438
rect 1650 5433 1651 5437
rect 1655 5433 1656 5437
rect 1650 5432 1656 5433
rect 1786 5437 1792 5438
rect 1786 5433 1787 5437
rect 1791 5433 1792 5437
rect 1786 5432 1792 5433
rect 1934 5436 1940 5437
rect 1934 5432 1935 5436
rect 1939 5432 1940 5436
rect 110 5431 116 5432
rect 112 5267 114 5431
rect 564 5267 566 5432
rect 700 5267 702 5432
rect 836 5267 838 5432
rect 972 5267 974 5432
rect 1108 5267 1110 5432
rect 1244 5267 1246 5432
rect 1380 5267 1382 5432
rect 1516 5267 1518 5432
rect 1652 5267 1654 5432
rect 1788 5267 1790 5432
rect 1934 5431 1940 5432
rect 1936 5267 1938 5431
rect 1976 5397 1978 5457
rect 1974 5396 1980 5397
rect 2428 5396 2430 5457
rect 2644 5396 2646 5457
rect 2860 5396 2862 5457
rect 3076 5396 3078 5457
rect 3292 5396 3294 5457
rect 3800 5397 3802 5457
rect 3840 5423 3842 5487
rect 3860 5423 3862 5488
rect 4100 5423 4102 5488
rect 4348 5423 4350 5488
rect 4588 5423 4590 5488
rect 4820 5423 4822 5488
rect 5052 5423 5054 5488
rect 5284 5423 5286 5488
rect 5662 5487 5668 5488
rect 5664 5423 5666 5487
rect 3839 5422 3843 5423
rect 3839 5417 3843 5418
rect 3859 5422 3863 5423
rect 3859 5417 3863 5418
rect 4075 5422 4079 5423
rect 4075 5417 4079 5418
rect 4099 5422 4103 5423
rect 4099 5417 4103 5418
rect 4307 5422 4311 5423
rect 4307 5417 4311 5418
rect 4347 5422 4351 5423
rect 4347 5417 4351 5418
rect 4531 5422 4535 5423
rect 4531 5417 4535 5418
rect 4587 5422 4591 5423
rect 4587 5417 4591 5418
rect 4739 5422 4743 5423
rect 4739 5417 4743 5418
rect 4819 5422 4823 5423
rect 4819 5417 4823 5418
rect 4939 5422 4943 5423
rect 4939 5417 4943 5418
rect 5051 5422 5055 5423
rect 5051 5417 5055 5418
rect 5139 5422 5143 5423
rect 5139 5417 5143 5418
rect 5283 5422 5287 5423
rect 5283 5417 5287 5418
rect 5339 5422 5343 5423
rect 5339 5417 5343 5418
rect 5515 5422 5519 5423
rect 5515 5417 5519 5418
rect 5663 5422 5667 5423
rect 5663 5417 5667 5418
rect 3798 5396 3804 5397
rect 1974 5392 1975 5396
rect 1979 5392 1980 5396
rect 1974 5391 1980 5392
rect 2426 5395 2432 5396
rect 2426 5391 2427 5395
rect 2431 5391 2432 5395
rect 2426 5390 2432 5391
rect 2642 5395 2648 5396
rect 2642 5391 2643 5395
rect 2647 5391 2648 5395
rect 2642 5390 2648 5391
rect 2858 5395 2864 5396
rect 2858 5391 2859 5395
rect 2863 5391 2864 5395
rect 2858 5390 2864 5391
rect 3074 5395 3080 5396
rect 3074 5391 3075 5395
rect 3079 5391 3080 5395
rect 3074 5390 3080 5391
rect 3290 5395 3296 5396
rect 3290 5391 3291 5395
rect 3295 5391 3296 5395
rect 3798 5392 3799 5396
rect 3803 5392 3804 5396
rect 3798 5391 3804 5392
rect 3290 5390 3296 5391
rect 2454 5380 2460 5381
rect 1974 5379 1980 5380
rect 1974 5375 1975 5379
rect 1979 5375 1980 5379
rect 2454 5376 2455 5380
rect 2459 5376 2460 5380
rect 2454 5375 2460 5376
rect 2670 5380 2676 5381
rect 2670 5376 2671 5380
rect 2675 5376 2676 5380
rect 2670 5375 2676 5376
rect 2886 5380 2892 5381
rect 2886 5376 2887 5380
rect 2891 5376 2892 5380
rect 2886 5375 2892 5376
rect 3102 5380 3108 5381
rect 3102 5376 3103 5380
rect 3107 5376 3108 5380
rect 3102 5375 3108 5376
rect 3318 5380 3324 5381
rect 3318 5376 3319 5380
rect 3323 5376 3324 5380
rect 3318 5375 3324 5376
rect 3798 5379 3804 5380
rect 3798 5375 3799 5379
rect 3803 5375 3804 5379
rect 1974 5374 1980 5375
rect 1976 5351 1978 5374
rect 2456 5351 2458 5375
rect 2672 5351 2674 5375
rect 2888 5351 2890 5375
rect 3104 5351 3106 5375
rect 3320 5351 3322 5375
rect 3798 5374 3804 5375
rect 3800 5351 3802 5374
rect 3840 5357 3842 5417
rect 3838 5356 3844 5357
rect 3860 5356 3862 5417
rect 4076 5356 4078 5417
rect 4308 5356 4310 5417
rect 4532 5356 4534 5417
rect 4740 5356 4742 5417
rect 4940 5356 4942 5417
rect 5140 5356 5142 5417
rect 5340 5356 5342 5417
rect 5516 5356 5518 5417
rect 5664 5357 5666 5417
rect 5662 5356 5668 5357
rect 3838 5352 3839 5356
rect 3843 5352 3844 5356
rect 3838 5351 3844 5352
rect 3858 5355 3864 5356
rect 3858 5351 3859 5355
rect 3863 5351 3864 5355
rect 1975 5350 1979 5351
rect 1975 5345 1979 5346
rect 2447 5350 2451 5351
rect 2447 5345 2451 5346
rect 2455 5350 2459 5351
rect 2455 5345 2459 5346
rect 2583 5350 2587 5351
rect 2583 5345 2587 5346
rect 2671 5350 2675 5351
rect 2671 5345 2675 5346
rect 2719 5350 2723 5351
rect 2719 5345 2723 5346
rect 2855 5350 2859 5351
rect 2855 5345 2859 5346
rect 2887 5350 2891 5351
rect 2887 5345 2891 5346
rect 2991 5350 2995 5351
rect 2991 5345 2995 5346
rect 3103 5350 3107 5351
rect 3103 5345 3107 5346
rect 3135 5350 3139 5351
rect 3135 5345 3139 5346
rect 3287 5350 3291 5351
rect 3287 5345 3291 5346
rect 3319 5350 3323 5351
rect 3319 5345 3323 5346
rect 3799 5350 3803 5351
rect 3858 5350 3864 5351
rect 4074 5355 4080 5356
rect 4074 5351 4075 5355
rect 4079 5351 4080 5355
rect 4074 5350 4080 5351
rect 4306 5355 4312 5356
rect 4306 5351 4307 5355
rect 4311 5351 4312 5355
rect 4306 5350 4312 5351
rect 4530 5355 4536 5356
rect 4530 5351 4531 5355
rect 4535 5351 4536 5355
rect 4530 5350 4536 5351
rect 4738 5355 4744 5356
rect 4738 5351 4739 5355
rect 4743 5351 4744 5355
rect 4738 5350 4744 5351
rect 4938 5355 4944 5356
rect 4938 5351 4939 5355
rect 4943 5351 4944 5355
rect 4938 5350 4944 5351
rect 5138 5355 5144 5356
rect 5138 5351 5139 5355
rect 5143 5351 5144 5355
rect 5138 5350 5144 5351
rect 5338 5355 5344 5356
rect 5338 5351 5339 5355
rect 5343 5351 5344 5355
rect 5338 5350 5344 5351
rect 5514 5355 5520 5356
rect 5514 5351 5515 5355
rect 5519 5351 5520 5355
rect 5662 5352 5663 5356
rect 5667 5352 5668 5356
rect 5662 5351 5668 5352
rect 5514 5350 5520 5351
rect 3799 5345 3803 5346
rect 1976 5322 1978 5345
rect 1974 5321 1980 5322
rect 2448 5321 2450 5345
rect 2584 5321 2586 5345
rect 2720 5321 2722 5345
rect 2856 5321 2858 5345
rect 2992 5321 2994 5345
rect 3136 5321 3138 5345
rect 3288 5321 3290 5345
rect 3800 5322 3802 5345
rect 3886 5340 3892 5341
rect 3838 5339 3844 5340
rect 3838 5335 3839 5339
rect 3843 5335 3844 5339
rect 3886 5336 3887 5340
rect 3891 5336 3892 5340
rect 3886 5335 3892 5336
rect 4102 5340 4108 5341
rect 4102 5336 4103 5340
rect 4107 5336 4108 5340
rect 4102 5335 4108 5336
rect 4334 5340 4340 5341
rect 4334 5336 4335 5340
rect 4339 5336 4340 5340
rect 4334 5335 4340 5336
rect 4558 5340 4564 5341
rect 4558 5336 4559 5340
rect 4563 5336 4564 5340
rect 4558 5335 4564 5336
rect 4766 5340 4772 5341
rect 4766 5336 4767 5340
rect 4771 5336 4772 5340
rect 4766 5335 4772 5336
rect 4966 5340 4972 5341
rect 4966 5336 4967 5340
rect 4971 5336 4972 5340
rect 4966 5335 4972 5336
rect 5166 5340 5172 5341
rect 5166 5336 5167 5340
rect 5171 5336 5172 5340
rect 5166 5335 5172 5336
rect 5366 5340 5372 5341
rect 5366 5336 5367 5340
rect 5371 5336 5372 5340
rect 5366 5335 5372 5336
rect 5542 5340 5548 5341
rect 5542 5336 5543 5340
rect 5547 5336 5548 5340
rect 5542 5335 5548 5336
rect 5662 5339 5668 5340
rect 5662 5335 5663 5339
rect 5667 5335 5668 5339
rect 3838 5334 3844 5335
rect 3798 5321 3804 5322
rect 1974 5317 1975 5321
rect 1979 5317 1980 5321
rect 1974 5316 1980 5317
rect 2446 5320 2452 5321
rect 2446 5316 2447 5320
rect 2451 5316 2452 5320
rect 2446 5315 2452 5316
rect 2582 5320 2588 5321
rect 2582 5316 2583 5320
rect 2587 5316 2588 5320
rect 2582 5315 2588 5316
rect 2718 5320 2724 5321
rect 2718 5316 2719 5320
rect 2723 5316 2724 5320
rect 2718 5315 2724 5316
rect 2854 5320 2860 5321
rect 2854 5316 2855 5320
rect 2859 5316 2860 5320
rect 2854 5315 2860 5316
rect 2990 5320 2996 5321
rect 2990 5316 2991 5320
rect 2995 5316 2996 5320
rect 2990 5315 2996 5316
rect 3134 5320 3140 5321
rect 3134 5316 3135 5320
rect 3139 5316 3140 5320
rect 3134 5315 3140 5316
rect 3286 5320 3292 5321
rect 3286 5316 3287 5320
rect 3291 5316 3292 5320
rect 3798 5317 3799 5321
rect 3803 5317 3804 5321
rect 3798 5316 3804 5317
rect 3286 5315 3292 5316
rect 2418 5305 2424 5306
rect 1974 5304 1980 5305
rect 1974 5300 1975 5304
rect 1979 5300 1980 5304
rect 2418 5301 2419 5305
rect 2423 5301 2424 5305
rect 2418 5300 2424 5301
rect 2554 5305 2560 5306
rect 2554 5301 2555 5305
rect 2559 5301 2560 5305
rect 2554 5300 2560 5301
rect 2690 5305 2696 5306
rect 2690 5301 2691 5305
rect 2695 5301 2696 5305
rect 2690 5300 2696 5301
rect 2826 5305 2832 5306
rect 2826 5301 2827 5305
rect 2831 5301 2832 5305
rect 2826 5300 2832 5301
rect 2962 5305 2968 5306
rect 2962 5301 2963 5305
rect 2967 5301 2968 5305
rect 2962 5300 2968 5301
rect 3106 5305 3112 5306
rect 3106 5301 3107 5305
rect 3111 5301 3112 5305
rect 3106 5300 3112 5301
rect 3258 5305 3264 5306
rect 3258 5301 3259 5305
rect 3263 5301 3264 5305
rect 3258 5300 3264 5301
rect 3798 5304 3804 5305
rect 3798 5300 3799 5304
rect 3803 5300 3804 5304
rect 1974 5299 1980 5300
rect 111 5266 115 5267
rect 111 5261 115 5262
rect 459 5266 463 5267
rect 459 5261 463 5262
rect 563 5266 567 5267
rect 563 5261 567 5262
rect 595 5266 599 5267
rect 595 5261 599 5262
rect 699 5266 703 5267
rect 699 5261 703 5262
rect 731 5266 735 5267
rect 731 5261 735 5262
rect 835 5266 839 5267
rect 835 5261 839 5262
rect 867 5266 871 5267
rect 867 5261 871 5262
rect 971 5266 975 5267
rect 971 5261 975 5262
rect 1003 5266 1007 5267
rect 1003 5261 1007 5262
rect 1107 5266 1111 5267
rect 1107 5261 1111 5262
rect 1139 5266 1143 5267
rect 1139 5261 1143 5262
rect 1243 5266 1247 5267
rect 1243 5261 1247 5262
rect 1275 5266 1279 5267
rect 1275 5261 1279 5262
rect 1379 5266 1383 5267
rect 1379 5261 1383 5262
rect 1411 5266 1415 5267
rect 1411 5261 1415 5262
rect 1515 5266 1519 5267
rect 1515 5261 1519 5262
rect 1547 5266 1551 5267
rect 1547 5261 1551 5262
rect 1651 5266 1655 5267
rect 1651 5261 1655 5262
rect 1787 5266 1791 5267
rect 1787 5261 1791 5262
rect 1935 5266 1939 5267
rect 1935 5261 1939 5262
rect 112 5201 114 5261
rect 110 5200 116 5201
rect 460 5200 462 5261
rect 596 5200 598 5261
rect 732 5200 734 5261
rect 868 5200 870 5261
rect 1004 5200 1006 5261
rect 1140 5200 1142 5261
rect 1276 5200 1278 5261
rect 1412 5200 1414 5261
rect 1548 5200 1550 5261
rect 1936 5201 1938 5261
rect 1976 5239 1978 5299
rect 2420 5239 2422 5300
rect 2556 5239 2558 5300
rect 2692 5239 2694 5300
rect 2828 5239 2830 5300
rect 2964 5239 2966 5300
rect 3108 5239 3110 5300
rect 3260 5239 3262 5300
rect 3798 5299 3804 5300
rect 3800 5239 3802 5299
rect 3840 5295 3842 5334
rect 3888 5295 3890 5335
rect 4104 5295 4106 5335
rect 4336 5295 4338 5335
rect 4560 5295 4562 5335
rect 4768 5295 4770 5335
rect 4968 5295 4970 5335
rect 5168 5295 5170 5335
rect 5368 5295 5370 5335
rect 5544 5295 5546 5335
rect 5662 5334 5668 5335
rect 5664 5295 5666 5334
rect 3839 5294 3843 5295
rect 3839 5289 3843 5290
rect 3887 5294 3891 5295
rect 3887 5289 3891 5290
rect 4095 5294 4099 5295
rect 4095 5289 4099 5290
rect 4103 5294 4107 5295
rect 4103 5289 4107 5290
rect 4335 5294 4339 5295
rect 4335 5289 4339 5290
rect 4343 5294 4347 5295
rect 4343 5289 4347 5290
rect 4559 5294 4563 5295
rect 4559 5289 4563 5290
rect 4615 5294 4619 5295
rect 4615 5289 4619 5290
rect 4767 5294 4771 5295
rect 4767 5289 4771 5290
rect 4911 5294 4915 5295
rect 4911 5289 4915 5290
rect 4967 5294 4971 5295
rect 4967 5289 4971 5290
rect 5167 5294 5171 5295
rect 5167 5289 5171 5290
rect 5215 5294 5219 5295
rect 5215 5289 5219 5290
rect 5367 5294 5371 5295
rect 5367 5289 5371 5290
rect 5527 5294 5531 5295
rect 5527 5289 5531 5290
rect 5543 5294 5547 5295
rect 5543 5289 5547 5290
rect 5663 5294 5667 5295
rect 5663 5289 5667 5290
rect 3840 5266 3842 5289
rect 3838 5265 3844 5266
rect 3888 5265 3890 5289
rect 4096 5265 4098 5289
rect 4344 5265 4346 5289
rect 4616 5265 4618 5289
rect 4912 5265 4914 5289
rect 5216 5265 5218 5289
rect 5528 5265 5530 5289
rect 5664 5266 5666 5289
rect 5662 5265 5668 5266
rect 3838 5261 3839 5265
rect 3843 5261 3844 5265
rect 3838 5260 3844 5261
rect 3886 5264 3892 5265
rect 3886 5260 3887 5264
rect 3891 5260 3892 5264
rect 3886 5259 3892 5260
rect 4094 5264 4100 5265
rect 4094 5260 4095 5264
rect 4099 5260 4100 5264
rect 4094 5259 4100 5260
rect 4342 5264 4348 5265
rect 4342 5260 4343 5264
rect 4347 5260 4348 5264
rect 4342 5259 4348 5260
rect 4614 5264 4620 5265
rect 4614 5260 4615 5264
rect 4619 5260 4620 5264
rect 4614 5259 4620 5260
rect 4910 5264 4916 5265
rect 4910 5260 4911 5264
rect 4915 5260 4916 5264
rect 4910 5259 4916 5260
rect 5214 5264 5220 5265
rect 5214 5260 5215 5264
rect 5219 5260 5220 5264
rect 5214 5259 5220 5260
rect 5526 5264 5532 5265
rect 5526 5260 5527 5264
rect 5531 5260 5532 5264
rect 5662 5261 5663 5265
rect 5667 5261 5668 5265
rect 5662 5260 5668 5261
rect 5526 5259 5532 5260
rect 3858 5249 3864 5250
rect 3838 5248 3844 5249
rect 3838 5244 3839 5248
rect 3843 5244 3844 5248
rect 3858 5245 3859 5249
rect 3863 5245 3864 5249
rect 3858 5244 3864 5245
rect 4066 5249 4072 5250
rect 4066 5245 4067 5249
rect 4071 5245 4072 5249
rect 4066 5244 4072 5245
rect 4314 5249 4320 5250
rect 4314 5245 4315 5249
rect 4319 5245 4320 5249
rect 4314 5244 4320 5245
rect 4586 5249 4592 5250
rect 4586 5245 4587 5249
rect 4591 5245 4592 5249
rect 4586 5244 4592 5245
rect 4882 5249 4888 5250
rect 4882 5245 4883 5249
rect 4887 5245 4888 5249
rect 4882 5244 4888 5245
rect 5186 5249 5192 5250
rect 5186 5245 5187 5249
rect 5191 5245 5192 5249
rect 5186 5244 5192 5245
rect 5498 5249 5504 5250
rect 5498 5245 5499 5249
rect 5503 5245 5504 5249
rect 5498 5244 5504 5245
rect 5662 5248 5668 5249
rect 5662 5244 5663 5248
rect 5667 5244 5668 5248
rect 3838 5243 3844 5244
rect 1975 5238 1979 5239
rect 1975 5233 1979 5234
rect 2099 5238 2103 5239
rect 2099 5233 2103 5234
rect 2235 5238 2239 5239
rect 2235 5233 2239 5234
rect 2379 5238 2383 5239
rect 2379 5233 2383 5234
rect 2419 5238 2423 5239
rect 2419 5233 2423 5234
rect 2531 5238 2535 5239
rect 2531 5233 2535 5234
rect 2555 5238 2559 5239
rect 2555 5233 2559 5234
rect 2691 5238 2695 5239
rect 2691 5233 2695 5234
rect 2699 5238 2703 5239
rect 2699 5233 2703 5234
rect 2827 5238 2831 5239
rect 2827 5233 2831 5234
rect 2883 5238 2887 5239
rect 2883 5233 2887 5234
rect 2963 5238 2967 5239
rect 2963 5233 2967 5234
rect 3067 5238 3071 5239
rect 3067 5233 3071 5234
rect 3107 5238 3111 5239
rect 3107 5233 3111 5234
rect 3259 5238 3263 5239
rect 3259 5233 3263 5234
rect 3799 5238 3803 5239
rect 3799 5233 3803 5234
rect 1934 5200 1940 5201
rect 110 5196 111 5200
rect 115 5196 116 5200
rect 110 5195 116 5196
rect 458 5199 464 5200
rect 458 5195 459 5199
rect 463 5195 464 5199
rect 458 5194 464 5195
rect 594 5199 600 5200
rect 594 5195 595 5199
rect 599 5195 600 5199
rect 594 5194 600 5195
rect 730 5199 736 5200
rect 730 5195 731 5199
rect 735 5195 736 5199
rect 730 5194 736 5195
rect 866 5199 872 5200
rect 866 5195 867 5199
rect 871 5195 872 5199
rect 866 5194 872 5195
rect 1002 5199 1008 5200
rect 1002 5195 1003 5199
rect 1007 5195 1008 5199
rect 1002 5194 1008 5195
rect 1138 5199 1144 5200
rect 1138 5195 1139 5199
rect 1143 5195 1144 5199
rect 1138 5194 1144 5195
rect 1274 5199 1280 5200
rect 1274 5195 1275 5199
rect 1279 5195 1280 5199
rect 1274 5194 1280 5195
rect 1410 5199 1416 5200
rect 1410 5195 1411 5199
rect 1415 5195 1416 5199
rect 1410 5194 1416 5195
rect 1546 5199 1552 5200
rect 1546 5195 1547 5199
rect 1551 5195 1552 5199
rect 1934 5196 1935 5200
rect 1939 5196 1940 5200
rect 1934 5195 1940 5196
rect 1546 5194 1552 5195
rect 486 5184 492 5185
rect 110 5183 116 5184
rect 110 5179 111 5183
rect 115 5179 116 5183
rect 486 5180 487 5184
rect 491 5180 492 5184
rect 486 5179 492 5180
rect 622 5184 628 5185
rect 622 5180 623 5184
rect 627 5180 628 5184
rect 622 5179 628 5180
rect 758 5184 764 5185
rect 758 5180 759 5184
rect 763 5180 764 5184
rect 758 5179 764 5180
rect 894 5184 900 5185
rect 894 5180 895 5184
rect 899 5180 900 5184
rect 894 5179 900 5180
rect 1030 5184 1036 5185
rect 1030 5180 1031 5184
rect 1035 5180 1036 5184
rect 1030 5179 1036 5180
rect 1166 5184 1172 5185
rect 1166 5180 1167 5184
rect 1171 5180 1172 5184
rect 1166 5179 1172 5180
rect 1302 5184 1308 5185
rect 1302 5180 1303 5184
rect 1307 5180 1308 5184
rect 1302 5179 1308 5180
rect 1438 5184 1444 5185
rect 1438 5180 1439 5184
rect 1443 5180 1444 5184
rect 1438 5179 1444 5180
rect 1574 5184 1580 5185
rect 1574 5180 1575 5184
rect 1579 5180 1580 5184
rect 1574 5179 1580 5180
rect 1934 5183 1940 5184
rect 1934 5179 1935 5183
rect 1939 5179 1940 5183
rect 110 5178 116 5179
rect 112 5139 114 5178
rect 488 5139 490 5179
rect 624 5139 626 5179
rect 760 5139 762 5179
rect 896 5139 898 5179
rect 1032 5139 1034 5179
rect 1168 5139 1170 5179
rect 1304 5139 1306 5179
rect 1440 5139 1442 5179
rect 1576 5139 1578 5179
rect 1934 5178 1940 5179
rect 1936 5139 1938 5178
rect 1976 5173 1978 5233
rect 1974 5172 1980 5173
rect 2100 5172 2102 5233
rect 2236 5172 2238 5233
rect 2380 5172 2382 5233
rect 2532 5172 2534 5233
rect 2700 5172 2702 5233
rect 2884 5172 2886 5233
rect 3068 5172 3070 5233
rect 3260 5172 3262 5233
rect 3800 5173 3802 5233
rect 3840 5175 3842 5243
rect 3860 5175 3862 5244
rect 4068 5175 4070 5244
rect 4316 5175 4318 5244
rect 4588 5175 4590 5244
rect 4884 5175 4886 5244
rect 5188 5175 5190 5244
rect 5500 5175 5502 5244
rect 5662 5243 5668 5244
rect 5664 5175 5666 5243
rect 3839 5174 3843 5175
rect 3798 5172 3804 5173
rect 1974 5168 1975 5172
rect 1979 5168 1980 5172
rect 1974 5167 1980 5168
rect 2098 5171 2104 5172
rect 2098 5167 2099 5171
rect 2103 5167 2104 5171
rect 2098 5166 2104 5167
rect 2234 5171 2240 5172
rect 2234 5167 2235 5171
rect 2239 5167 2240 5171
rect 2234 5166 2240 5167
rect 2378 5171 2384 5172
rect 2378 5167 2379 5171
rect 2383 5167 2384 5171
rect 2378 5166 2384 5167
rect 2530 5171 2536 5172
rect 2530 5167 2531 5171
rect 2535 5167 2536 5171
rect 2530 5166 2536 5167
rect 2698 5171 2704 5172
rect 2698 5167 2699 5171
rect 2703 5167 2704 5171
rect 2698 5166 2704 5167
rect 2882 5171 2888 5172
rect 2882 5167 2883 5171
rect 2887 5167 2888 5171
rect 2882 5166 2888 5167
rect 3066 5171 3072 5172
rect 3066 5167 3067 5171
rect 3071 5167 3072 5171
rect 3066 5166 3072 5167
rect 3258 5171 3264 5172
rect 3258 5167 3259 5171
rect 3263 5167 3264 5171
rect 3798 5168 3799 5172
rect 3803 5168 3804 5172
rect 3839 5169 3843 5170
rect 3859 5174 3863 5175
rect 3859 5169 3863 5170
rect 3995 5174 3999 5175
rect 3995 5169 3999 5170
rect 4067 5174 4071 5175
rect 4067 5169 4071 5170
rect 4155 5174 4159 5175
rect 4155 5169 4159 5170
rect 4315 5174 4319 5175
rect 4315 5169 4319 5170
rect 4363 5174 4367 5175
rect 4363 5169 4367 5170
rect 4587 5174 4591 5175
rect 4587 5169 4591 5170
rect 4611 5174 4615 5175
rect 4611 5169 4615 5170
rect 4883 5174 4887 5175
rect 4883 5169 4887 5170
rect 5171 5174 5175 5175
rect 5171 5169 5175 5170
rect 5187 5174 5191 5175
rect 5187 5169 5191 5170
rect 5467 5174 5471 5175
rect 5467 5169 5471 5170
rect 5499 5174 5503 5175
rect 5499 5169 5503 5170
rect 5663 5174 5667 5175
rect 5663 5169 5667 5170
rect 3798 5167 3804 5168
rect 3258 5166 3264 5167
rect 2126 5156 2132 5157
rect 1974 5155 1980 5156
rect 1974 5151 1975 5155
rect 1979 5151 1980 5155
rect 2126 5152 2127 5156
rect 2131 5152 2132 5156
rect 2126 5151 2132 5152
rect 2262 5156 2268 5157
rect 2262 5152 2263 5156
rect 2267 5152 2268 5156
rect 2262 5151 2268 5152
rect 2406 5156 2412 5157
rect 2406 5152 2407 5156
rect 2411 5152 2412 5156
rect 2406 5151 2412 5152
rect 2558 5156 2564 5157
rect 2558 5152 2559 5156
rect 2563 5152 2564 5156
rect 2558 5151 2564 5152
rect 2726 5156 2732 5157
rect 2726 5152 2727 5156
rect 2731 5152 2732 5156
rect 2726 5151 2732 5152
rect 2910 5156 2916 5157
rect 2910 5152 2911 5156
rect 2915 5152 2916 5156
rect 2910 5151 2916 5152
rect 3094 5156 3100 5157
rect 3094 5152 3095 5156
rect 3099 5152 3100 5156
rect 3094 5151 3100 5152
rect 3286 5156 3292 5157
rect 3286 5152 3287 5156
rect 3291 5152 3292 5156
rect 3286 5151 3292 5152
rect 3798 5155 3804 5156
rect 3798 5151 3799 5155
rect 3803 5151 3804 5155
rect 1974 5150 1980 5151
rect 111 5138 115 5139
rect 111 5133 115 5134
rect 319 5138 323 5139
rect 319 5133 323 5134
rect 487 5138 491 5139
rect 487 5133 491 5134
rect 503 5138 507 5139
rect 503 5133 507 5134
rect 623 5138 627 5139
rect 623 5133 627 5134
rect 703 5138 707 5139
rect 703 5133 707 5134
rect 759 5138 763 5139
rect 759 5133 763 5134
rect 895 5138 899 5139
rect 895 5133 899 5134
rect 919 5138 923 5139
rect 919 5133 923 5134
rect 1031 5138 1035 5139
rect 1031 5133 1035 5134
rect 1151 5138 1155 5139
rect 1151 5133 1155 5134
rect 1167 5138 1171 5139
rect 1167 5133 1171 5134
rect 1303 5138 1307 5139
rect 1303 5133 1307 5134
rect 1391 5138 1395 5139
rect 1391 5133 1395 5134
rect 1439 5138 1443 5139
rect 1439 5133 1443 5134
rect 1575 5138 1579 5139
rect 1575 5133 1579 5134
rect 1631 5138 1635 5139
rect 1631 5133 1635 5134
rect 1935 5138 1939 5139
rect 1935 5133 1939 5134
rect 112 5110 114 5133
rect 110 5109 116 5110
rect 320 5109 322 5133
rect 504 5109 506 5133
rect 704 5109 706 5133
rect 920 5109 922 5133
rect 1152 5109 1154 5133
rect 1392 5109 1394 5133
rect 1632 5109 1634 5133
rect 1936 5110 1938 5133
rect 1934 5109 1940 5110
rect 110 5105 111 5109
rect 115 5105 116 5109
rect 110 5104 116 5105
rect 318 5108 324 5109
rect 318 5104 319 5108
rect 323 5104 324 5108
rect 318 5103 324 5104
rect 502 5108 508 5109
rect 502 5104 503 5108
rect 507 5104 508 5108
rect 502 5103 508 5104
rect 702 5108 708 5109
rect 702 5104 703 5108
rect 707 5104 708 5108
rect 702 5103 708 5104
rect 918 5108 924 5109
rect 918 5104 919 5108
rect 923 5104 924 5108
rect 918 5103 924 5104
rect 1150 5108 1156 5109
rect 1150 5104 1151 5108
rect 1155 5104 1156 5108
rect 1150 5103 1156 5104
rect 1390 5108 1396 5109
rect 1390 5104 1391 5108
rect 1395 5104 1396 5108
rect 1390 5103 1396 5104
rect 1630 5108 1636 5109
rect 1630 5104 1631 5108
rect 1635 5104 1636 5108
rect 1934 5105 1935 5109
rect 1939 5105 1940 5109
rect 1934 5104 1940 5105
rect 1630 5103 1636 5104
rect 1976 5103 1978 5150
rect 2128 5103 2130 5151
rect 2264 5103 2266 5151
rect 2408 5103 2410 5151
rect 2560 5103 2562 5151
rect 2728 5103 2730 5151
rect 2912 5103 2914 5151
rect 3096 5103 3098 5151
rect 3288 5103 3290 5151
rect 3798 5150 3804 5151
rect 3800 5103 3802 5150
rect 3840 5109 3842 5169
rect 3838 5108 3844 5109
rect 3860 5108 3862 5169
rect 3996 5108 3998 5169
rect 4156 5108 4158 5169
rect 4364 5108 4366 5169
rect 4612 5108 4614 5169
rect 4884 5108 4886 5169
rect 5172 5108 5174 5169
rect 5468 5108 5470 5169
rect 5664 5109 5666 5169
rect 5662 5108 5668 5109
rect 3838 5104 3839 5108
rect 3843 5104 3844 5108
rect 3838 5103 3844 5104
rect 3858 5107 3864 5108
rect 3858 5103 3859 5107
rect 3863 5103 3864 5107
rect 1975 5102 1979 5103
rect 1975 5097 1979 5098
rect 2079 5102 2083 5103
rect 2079 5097 2083 5098
rect 2127 5102 2131 5103
rect 2127 5097 2131 5098
rect 2263 5102 2267 5103
rect 2263 5097 2267 5098
rect 2359 5102 2363 5103
rect 2359 5097 2363 5098
rect 2407 5102 2411 5103
rect 2407 5097 2411 5098
rect 2559 5102 2563 5103
rect 2559 5097 2563 5098
rect 2639 5102 2643 5103
rect 2639 5097 2643 5098
rect 2727 5102 2731 5103
rect 2727 5097 2731 5098
rect 2911 5102 2915 5103
rect 2911 5097 2915 5098
rect 3095 5102 3099 5103
rect 3095 5097 3099 5098
rect 3175 5102 3179 5103
rect 3175 5097 3179 5098
rect 3287 5102 3291 5103
rect 3287 5097 3291 5098
rect 3439 5102 3443 5103
rect 3439 5097 3443 5098
rect 3679 5102 3683 5103
rect 3679 5097 3683 5098
rect 3799 5102 3803 5103
rect 3858 5102 3864 5103
rect 3994 5107 4000 5108
rect 3994 5103 3995 5107
rect 3999 5103 4000 5107
rect 3994 5102 4000 5103
rect 4154 5107 4160 5108
rect 4154 5103 4155 5107
rect 4159 5103 4160 5107
rect 4154 5102 4160 5103
rect 4362 5107 4368 5108
rect 4362 5103 4363 5107
rect 4367 5103 4368 5107
rect 4362 5102 4368 5103
rect 4610 5107 4616 5108
rect 4610 5103 4611 5107
rect 4615 5103 4616 5107
rect 4610 5102 4616 5103
rect 4882 5107 4888 5108
rect 4882 5103 4883 5107
rect 4887 5103 4888 5107
rect 4882 5102 4888 5103
rect 5170 5107 5176 5108
rect 5170 5103 5171 5107
rect 5175 5103 5176 5107
rect 5170 5102 5176 5103
rect 5466 5107 5472 5108
rect 5466 5103 5467 5107
rect 5471 5103 5472 5107
rect 5662 5104 5663 5108
rect 5667 5104 5668 5108
rect 5662 5103 5668 5104
rect 5466 5102 5472 5103
rect 3799 5097 3803 5098
rect 290 5093 296 5094
rect 110 5092 116 5093
rect 110 5088 111 5092
rect 115 5088 116 5092
rect 290 5089 291 5093
rect 295 5089 296 5093
rect 290 5088 296 5089
rect 474 5093 480 5094
rect 474 5089 475 5093
rect 479 5089 480 5093
rect 474 5088 480 5089
rect 674 5093 680 5094
rect 674 5089 675 5093
rect 679 5089 680 5093
rect 674 5088 680 5089
rect 890 5093 896 5094
rect 890 5089 891 5093
rect 895 5089 896 5093
rect 890 5088 896 5089
rect 1122 5093 1128 5094
rect 1122 5089 1123 5093
rect 1127 5089 1128 5093
rect 1122 5088 1128 5089
rect 1362 5093 1368 5094
rect 1362 5089 1363 5093
rect 1367 5089 1368 5093
rect 1362 5088 1368 5089
rect 1602 5093 1608 5094
rect 1602 5089 1603 5093
rect 1607 5089 1608 5093
rect 1602 5088 1608 5089
rect 1934 5092 1940 5093
rect 1934 5088 1935 5092
rect 1939 5088 1940 5092
rect 110 5087 116 5088
rect 112 5027 114 5087
rect 292 5027 294 5088
rect 476 5027 478 5088
rect 676 5027 678 5088
rect 892 5027 894 5088
rect 1124 5027 1126 5088
rect 1364 5027 1366 5088
rect 1604 5027 1606 5088
rect 1934 5087 1940 5088
rect 1936 5027 1938 5087
rect 1976 5074 1978 5097
rect 1974 5073 1980 5074
rect 2080 5073 2082 5097
rect 2360 5073 2362 5097
rect 2640 5073 2642 5097
rect 2912 5073 2914 5097
rect 3176 5073 3178 5097
rect 3440 5073 3442 5097
rect 3680 5073 3682 5097
rect 3800 5074 3802 5097
rect 3886 5092 3892 5093
rect 3838 5091 3844 5092
rect 3838 5087 3839 5091
rect 3843 5087 3844 5091
rect 3886 5088 3887 5092
rect 3891 5088 3892 5092
rect 3886 5087 3892 5088
rect 4022 5092 4028 5093
rect 4022 5088 4023 5092
rect 4027 5088 4028 5092
rect 4022 5087 4028 5088
rect 4182 5092 4188 5093
rect 4182 5088 4183 5092
rect 4187 5088 4188 5092
rect 4182 5087 4188 5088
rect 4390 5092 4396 5093
rect 4390 5088 4391 5092
rect 4395 5088 4396 5092
rect 4390 5087 4396 5088
rect 4638 5092 4644 5093
rect 4638 5088 4639 5092
rect 4643 5088 4644 5092
rect 4638 5087 4644 5088
rect 4910 5092 4916 5093
rect 4910 5088 4911 5092
rect 4915 5088 4916 5092
rect 4910 5087 4916 5088
rect 5198 5092 5204 5093
rect 5198 5088 5199 5092
rect 5203 5088 5204 5092
rect 5198 5087 5204 5088
rect 5494 5092 5500 5093
rect 5494 5088 5495 5092
rect 5499 5088 5500 5092
rect 5494 5087 5500 5088
rect 5662 5091 5668 5092
rect 5662 5087 5663 5091
rect 5667 5087 5668 5091
rect 3838 5086 3844 5087
rect 3798 5073 3804 5074
rect 1974 5069 1975 5073
rect 1979 5069 1980 5073
rect 1974 5068 1980 5069
rect 2078 5072 2084 5073
rect 2078 5068 2079 5072
rect 2083 5068 2084 5072
rect 2078 5067 2084 5068
rect 2358 5072 2364 5073
rect 2358 5068 2359 5072
rect 2363 5068 2364 5072
rect 2358 5067 2364 5068
rect 2638 5072 2644 5073
rect 2638 5068 2639 5072
rect 2643 5068 2644 5072
rect 2638 5067 2644 5068
rect 2910 5072 2916 5073
rect 2910 5068 2911 5072
rect 2915 5068 2916 5072
rect 2910 5067 2916 5068
rect 3174 5072 3180 5073
rect 3174 5068 3175 5072
rect 3179 5068 3180 5072
rect 3174 5067 3180 5068
rect 3438 5072 3444 5073
rect 3438 5068 3439 5072
rect 3443 5068 3444 5072
rect 3438 5067 3444 5068
rect 3678 5072 3684 5073
rect 3678 5068 3679 5072
rect 3683 5068 3684 5072
rect 3798 5069 3799 5073
rect 3803 5069 3804 5073
rect 3798 5068 3804 5069
rect 3678 5067 3684 5068
rect 2050 5057 2056 5058
rect 1974 5056 1980 5057
rect 1974 5052 1975 5056
rect 1979 5052 1980 5056
rect 2050 5053 2051 5057
rect 2055 5053 2056 5057
rect 2050 5052 2056 5053
rect 2330 5057 2336 5058
rect 2330 5053 2331 5057
rect 2335 5053 2336 5057
rect 2330 5052 2336 5053
rect 2610 5057 2616 5058
rect 2610 5053 2611 5057
rect 2615 5053 2616 5057
rect 2610 5052 2616 5053
rect 2882 5057 2888 5058
rect 2882 5053 2883 5057
rect 2887 5053 2888 5057
rect 2882 5052 2888 5053
rect 3146 5057 3152 5058
rect 3146 5053 3147 5057
rect 3151 5053 3152 5057
rect 3146 5052 3152 5053
rect 3410 5057 3416 5058
rect 3410 5053 3411 5057
rect 3415 5053 3416 5057
rect 3410 5052 3416 5053
rect 3650 5057 3656 5058
rect 3650 5053 3651 5057
rect 3655 5053 3656 5057
rect 3650 5052 3656 5053
rect 3798 5056 3804 5057
rect 3798 5052 3799 5056
rect 3803 5052 3804 5056
rect 1974 5051 1980 5052
rect 111 5026 115 5027
rect 111 5021 115 5022
rect 139 5026 143 5027
rect 139 5021 143 5022
rect 291 5026 295 5027
rect 291 5021 295 5022
rect 411 5026 415 5027
rect 411 5021 415 5022
rect 475 5026 479 5027
rect 475 5021 479 5022
rect 675 5026 679 5027
rect 675 5021 679 5022
rect 683 5026 687 5027
rect 683 5021 687 5022
rect 891 5026 895 5027
rect 891 5021 895 5022
rect 963 5026 967 5027
rect 963 5021 967 5022
rect 1123 5026 1127 5027
rect 1123 5021 1127 5022
rect 1243 5026 1247 5027
rect 1243 5021 1247 5022
rect 1363 5026 1367 5027
rect 1363 5021 1367 5022
rect 1523 5026 1527 5027
rect 1523 5021 1527 5022
rect 1603 5026 1607 5027
rect 1603 5021 1607 5022
rect 1787 5026 1791 5027
rect 1787 5021 1791 5022
rect 1935 5026 1939 5027
rect 1935 5021 1939 5022
rect 112 4961 114 5021
rect 110 4960 116 4961
rect 140 4960 142 5021
rect 412 4960 414 5021
rect 684 4960 686 5021
rect 964 4960 966 5021
rect 1244 4960 1246 5021
rect 1524 4960 1526 5021
rect 1788 4960 1790 5021
rect 1936 4961 1938 5021
rect 1976 4971 1978 5051
rect 2052 4971 2054 5052
rect 2332 4971 2334 5052
rect 2612 4971 2614 5052
rect 2884 4971 2886 5052
rect 3148 4971 3150 5052
rect 3412 4971 3414 5052
rect 3652 4971 3654 5052
rect 3798 5051 3804 5052
rect 3800 4971 3802 5051
rect 3840 5047 3842 5086
rect 3888 5047 3890 5087
rect 4024 5047 4026 5087
rect 4184 5047 4186 5087
rect 4392 5047 4394 5087
rect 4640 5047 4642 5087
rect 4912 5047 4914 5087
rect 5200 5047 5202 5087
rect 5496 5047 5498 5087
rect 5662 5086 5668 5087
rect 5664 5047 5666 5086
rect 3839 5046 3843 5047
rect 3839 5041 3843 5042
rect 3887 5046 3891 5047
rect 3887 5041 3891 5042
rect 4023 5046 4027 5047
rect 4023 5041 4027 5042
rect 4183 5046 4187 5047
rect 4183 5041 4187 5042
rect 4391 5046 4395 5047
rect 4391 5041 4395 5042
rect 4447 5046 4451 5047
rect 4447 5041 4451 5042
rect 4631 5046 4635 5047
rect 4631 5041 4635 5042
rect 4639 5046 4643 5047
rect 4639 5041 4643 5042
rect 4831 5046 4835 5047
rect 4831 5041 4835 5042
rect 4911 5046 4915 5047
rect 4911 5041 4915 5042
rect 5047 5046 5051 5047
rect 5047 5041 5051 5042
rect 5199 5046 5203 5047
rect 5199 5041 5203 5042
rect 5279 5046 5283 5047
rect 5279 5041 5283 5042
rect 5495 5046 5499 5047
rect 5495 5041 5499 5042
rect 5511 5046 5515 5047
rect 5511 5041 5515 5042
rect 5663 5046 5667 5047
rect 5663 5041 5667 5042
rect 3840 5018 3842 5041
rect 3838 5017 3844 5018
rect 4448 5017 4450 5041
rect 4632 5017 4634 5041
rect 4832 5017 4834 5041
rect 5048 5017 5050 5041
rect 5280 5017 5282 5041
rect 5512 5017 5514 5041
rect 5664 5018 5666 5041
rect 5662 5017 5668 5018
rect 3838 5013 3839 5017
rect 3843 5013 3844 5017
rect 3838 5012 3844 5013
rect 4446 5016 4452 5017
rect 4446 5012 4447 5016
rect 4451 5012 4452 5016
rect 4446 5011 4452 5012
rect 4630 5016 4636 5017
rect 4630 5012 4631 5016
rect 4635 5012 4636 5016
rect 4630 5011 4636 5012
rect 4830 5016 4836 5017
rect 4830 5012 4831 5016
rect 4835 5012 4836 5016
rect 4830 5011 4836 5012
rect 5046 5016 5052 5017
rect 5046 5012 5047 5016
rect 5051 5012 5052 5016
rect 5046 5011 5052 5012
rect 5278 5016 5284 5017
rect 5278 5012 5279 5016
rect 5283 5012 5284 5016
rect 5278 5011 5284 5012
rect 5510 5016 5516 5017
rect 5510 5012 5511 5016
rect 5515 5012 5516 5016
rect 5662 5013 5663 5017
rect 5667 5013 5668 5017
rect 5662 5012 5668 5013
rect 5510 5011 5516 5012
rect 4418 5001 4424 5002
rect 3838 5000 3844 5001
rect 3838 4996 3839 5000
rect 3843 4996 3844 5000
rect 4418 4997 4419 5001
rect 4423 4997 4424 5001
rect 4418 4996 4424 4997
rect 4602 5001 4608 5002
rect 4602 4997 4603 5001
rect 4607 4997 4608 5001
rect 4602 4996 4608 4997
rect 4802 5001 4808 5002
rect 4802 4997 4803 5001
rect 4807 4997 4808 5001
rect 4802 4996 4808 4997
rect 5018 5001 5024 5002
rect 5018 4997 5019 5001
rect 5023 4997 5024 5001
rect 5018 4996 5024 4997
rect 5250 5001 5256 5002
rect 5250 4997 5251 5001
rect 5255 4997 5256 5001
rect 5250 4996 5256 4997
rect 5482 5001 5488 5002
rect 5482 4997 5483 5001
rect 5487 4997 5488 5001
rect 5482 4996 5488 4997
rect 5662 5000 5668 5001
rect 5662 4996 5663 5000
rect 5667 4996 5668 5000
rect 3838 4995 3844 4996
rect 1975 4970 1979 4971
rect 1975 4965 1979 4966
rect 1995 4970 1999 4971
rect 1995 4965 1999 4966
rect 2051 4970 2055 4971
rect 2051 4965 2055 4966
rect 2131 4970 2135 4971
rect 2131 4965 2135 4966
rect 2299 4970 2303 4971
rect 2299 4965 2303 4966
rect 2331 4970 2335 4971
rect 2331 4965 2335 4966
rect 2467 4970 2471 4971
rect 2467 4965 2471 4966
rect 2611 4970 2615 4971
rect 2611 4965 2615 4966
rect 2643 4970 2647 4971
rect 2643 4965 2647 4966
rect 2819 4970 2823 4971
rect 2819 4965 2823 4966
rect 2883 4970 2887 4971
rect 2883 4965 2887 4966
rect 2987 4970 2991 4971
rect 2987 4965 2991 4966
rect 3147 4970 3151 4971
rect 3147 4965 3151 4966
rect 3155 4970 3159 4971
rect 3155 4965 3159 4966
rect 3323 4970 3327 4971
rect 3323 4965 3327 4966
rect 3411 4970 3415 4971
rect 3411 4965 3415 4966
rect 3499 4970 3503 4971
rect 3499 4965 3503 4966
rect 3651 4970 3655 4971
rect 3651 4965 3655 4966
rect 3799 4970 3803 4971
rect 3799 4965 3803 4966
rect 1934 4960 1940 4961
rect 110 4956 111 4960
rect 115 4956 116 4960
rect 110 4955 116 4956
rect 138 4959 144 4960
rect 138 4955 139 4959
rect 143 4955 144 4959
rect 138 4954 144 4955
rect 410 4959 416 4960
rect 410 4955 411 4959
rect 415 4955 416 4959
rect 410 4954 416 4955
rect 682 4959 688 4960
rect 682 4955 683 4959
rect 687 4955 688 4959
rect 682 4954 688 4955
rect 962 4959 968 4960
rect 962 4955 963 4959
rect 967 4955 968 4959
rect 962 4954 968 4955
rect 1242 4959 1248 4960
rect 1242 4955 1243 4959
rect 1247 4955 1248 4959
rect 1242 4954 1248 4955
rect 1522 4959 1528 4960
rect 1522 4955 1523 4959
rect 1527 4955 1528 4959
rect 1522 4954 1528 4955
rect 1786 4959 1792 4960
rect 1786 4955 1787 4959
rect 1791 4955 1792 4959
rect 1934 4956 1935 4960
rect 1939 4956 1940 4960
rect 1934 4955 1940 4956
rect 1786 4954 1792 4955
rect 166 4944 172 4945
rect 110 4943 116 4944
rect 110 4939 111 4943
rect 115 4939 116 4943
rect 166 4940 167 4944
rect 171 4940 172 4944
rect 166 4939 172 4940
rect 438 4944 444 4945
rect 438 4940 439 4944
rect 443 4940 444 4944
rect 438 4939 444 4940
rect 710 4944 716 4945
rect 710 4940 711 4944
rect 715 4940 716 4944
rect 710 4939 716 4940
rect 990 4944 996 4945
rect 990 4940 991 4944
rect 995 4940 996 4944
rect 990 4939 996 4940
rect 1270 4944 1276 4945
rect 1270 4940 1271 4944
rect 1275 4940 1276 4944
rect 1270 4939 1276 4940
rect 1550 4944 1556 4945
rect 1550 4940 1551 4944
rect 1555 4940 1556 4944
rect 1550 4939 1556 4940
rect 1814 4944 1820 4945
rect 1814 4940 1815 4944
rect 1819 4940 1820 4944
rect 1814 4939 1820 4940
rect 1934 4943 1940 4944
rect 1934 4939 1935 4943
rect 1939 4939 1940 4943
rect 110 4938 116 4939
rect 112 4915 114 4938
rect 168 4915 170 4939
rect 440 4915 442 4939
rect 712 4915 714 4939
rect 992 4915 994 4939
rect 1272 4915 1274 4939
rect 1552 4915 1554 4939
rect 1816 4915 1818 4939
rect 1934 4938 1940 4939
rect 1936 4915 1938 4938
rect 111 4914 115 4915
rect 111 4909 115 4910
rect 159 4914 163 4915
rect 159 4909 163 4910
rect 167 4914 171 4915
rect 167 4909 171 4910
rect 415 4914 419 4915
rect 415 4909 419 4910
rect 439 4914 443 4915
rect 439 4909 443 4910
rect 711 4914 715 4915
rect 711 4909 715 4910
rect 735 4914 739 4915
rect 735 4909 739 4910
rect 991 4914 995 4915
rect 991 4909 995 4910
rect 1087 4914 1091 4915
rect 1087 4909 1091 4910
rect 1271 4914 1275 4915
rect 1271 4909 1275 4910
rect 1463 4914 1467 4915
rect 1463 4909 1467 4910
rect 1551 4914 1555 4915
rect 1551 4909 1555 4910
rect 1815 4914 1819 4915
rect 1815 4909 1819 4910
rect 1935 4914 1939 4915
rect 1935 4909 1939 4910
rect 112 4886 114 4909
rect 110 4885 116 4886
rect 160 4885 162 4909
rect 416 4885 418 4909
rect 736 4885 738 4909
rect 1088 4885 1090 4909
rect 1464 4885 1466 4909
rect 1816 4885 1818 4909
rect 1936 4886 1938 4909
rect 1976 4905 1978 4965
rect 1974 4904 1980 4905
rect 1996 4904 1998 4965
rect 2132 4904 2134 4965
rect 2300 4904 2302 4965
rect 2468 4904 2470 4965
rect 2644 4904 2646 4965
rect 2820 4904 2822 4965
rect 2988 4904 2990 4965
rect 3156 4904 3158 4965
rect 3324 4904 3326 4965
rect 3500 4904 3502 4965
rect 3652 4904 3654 4965
rect 3800 4905 3802 4965
rect 3840 4919 3842 4995
rect 4420 4919 4422 4996
rect 4604 4919 4606 4996
rect 4804 4919 4806 4996
rect 5020 4919 5022 4996
rect 5252 4919 5254 4996
rect 5484 4919 5486 4996
rect 5662 4995 5668 4996
rect 5664 4919 5666 4995
rect 3839 4918 3843 4919
rect 3839 4913 3843 4914
rect 4419 4918 4423 4919
rect 4419 4913 4423 4914
rect 4603 4918 4607 4919
rect 4603 4913 4607 4914
rect 4675 4918 4679 4919
rect 4675 4913 4679 4914
rect 4803 4918 4807 4919
rect 4803 4913 4807 4914
rect 4827 4918 4831 4919
rect 4827 4913 4831 4914
rect 4987 4918 4991 4919
rect 4987 4913 4991 4914
rect 5019 4918 5023 4919
rect 5019 4913 5023 4914
rect 5155 4918 5159 4919
rect 5155 4913 5159 4914
rect 5251 4918 5255 4919
rect 5251 4913 5255 4914
rect 5323 4918 5327 4919
rect 5323 4913 5327 4914
rect 5483 4918 5487 4919
rect 5483 4913 5487 4914
rect 5499 4918 5503 4919
rect 5499 4913 5503 4914
rect 5663 4918 5667 4919
rect 5663 4913 5667 4914
rect 3798 4904 3804 4905
rect 1974 4900 1975 4904
rect 1979 4900 1980 4904
rect 1974 4899 1980 4900
rect 1994 4903 2000 4904
rect 1994 4899 1995 4903
rect 1999 4899 2000 4903
rect 1994 4898 2000 4899
rect 2130 4903 2136 4904
rect 2130 4899 2131 4903
rect 2135 4899 2136 4903
rect 2130 4898 2136 4899
rect 2298 4903 2304 4904
rect 2298 4899 2299 4903
rect 2303 4899 2304 4903
rect 2298 4898 2304 4899
rect 2466 4903 2472 4904
rect 2466 4899 2467 4903
rect 2471 4899 2472 4903
rect 2466 4898 2472 4899
rect 2642 4903 2648 4904
rect 2642 4899 2643 4903
rect 2647 4899 2648 4903
rect 2642 4898 2648 4899
rect 2818 4903 2824 4904
rect 2818 4899 2819 4903
rect 2823 4899 2824 4903
rect 2818 4898 2824 4899
rect 2986 4903 2992 4904
rect 2986 4899 2987 4903
rect 2991 4899 2992 4903
rect 2986 4898 2992 4899
rect 3154 4903 3160 4904
rect 3154 4899 3155 4903
rect 3159 4899 3160 4903
rect 3154 4898 3160 4899
rect 3322 4903 3328 4904
rect 3322 4899 3323 4903
rect 3327 4899 3328 4903
rect 3322 4898 3328 4899
rect 3498 4903 3504 4904
rect 3498 4899 3499 4903
rect 3503 4899 3504 4903
rect 3498 4898 3504 4899
rect 3650 4903 3656 4904
rect 3650 4899 3651 4903
rect 3655 4899 3656 4903
rect 3798 4900 3799 4904
rect 3803 4900 3804 4904
rect 3798 4899 3804 4900
rect 3650 4898 3656 4899
rect 2022 4888 2028 4889
rect 1974 4887 1980 4888
rect 1934 4885 1940 4886
rect 110 4881 111 4885
rect 115 4881 116 4885
rect 110 4880 116 4881
rect 158 4884 164 4885
rect 158 4880 159 4884
rect 163 4880 164 4884
rect 158 4879 164 4880
rect 414 4884 420 4885
rect 414 4880 415 4884
rect 419 4880 420 4884
rect 414 4879 420 4880
rect 734 4884 740 4885
rect 734 4880 735 4884
rect 739 4880 740 4884
rect 734 4879 740 4880
rect 1086 4884 1092 4885
rect 1086 4880 1087 4884
rect 1091 4880 1092 4884
rect 1086 4879 1092 4880
rect 1462 4884 1468 4885
rect 1462 4880 1463 4884
rect 1467 4880 1468 4884
rect 1462 4879 1468 4880
rect 1814 4884 1820 4885
rect 1814 4880 1815 4884
rect 1819 4880 1820 4884
rect 1934 4881 1935 4885
rect 1939 4881 1940 4885
rect 1974 4883 1975 4887
rect 1979 4883 1980 4887
rect 2022 4884 2023 4888
rect 2027 4884 2028 4888
rect 2022 4883 2028 4884
rect 2158 4888 2164 4889
rect 2158 4884 2159 4888
rect 2163 4884 2164 4888
rect 2158 4883 2164 4884
rect 2326 4888 2332 4889
rect 2326 4884 2327 4888
rect 2331 4884 2332 4888
rect 2326 4883 2332 4884
rect 2494 4888 2500 4889
rect 2494 4884 2495 4888
rect 2499 4884 2500 4888
rect 2494 4883 2500 4884
rect 2670 4888 2676 4889
rect 2670 4884 2671 4888
rect 2675 4884 2676 4888
rect 2670 4883 2676 4884
rect 2846 4888 2852 4889
rect 2846 4884 2847 4888
rect 2851 4884 2852 4888
rect 2846 4883 2852 4884
rect 3014 4888 3020 4889
rect 3014 4884 3015 4888
rect 3019 4884 3020 4888
rect 3014 4883 3020 4884
rect 3182 4888 3188 4889
rect 3182 4884 3183 4888
rect 3187 4884 3188 4888
rect 3182 4883 3188 4884
rect 3350 4888 3356 4889
rect 3350 4884 3351 4888
rect 3355 4884 3356 4888
rect 3350 4883 3356 4884
rect 3526 4888 3532 4889
rect 3526 4884 3527 4888
rect 3531 4884 3532 4888
rect 3526 4883 3532 4884
rect 3678 4888 3684 4889
rect 3678 4884 3679 4888
rect 3683 4884 3684 4888
rect 3678 4883 3684 4884
rect 3798 4887 3804 4888
rect 3798 4883 3799 4887
rect 3803 4883 3804 4887
rect 1974 4882 1980 4883
rect 1934 4880 1940 4881
rect 1814 4879 1820 4880
rect 130 4869 136 4870
rect 110 4868 116 4869
rect 110 4864 111 4868
rect 115 4864 116 4868
rect 130 4865 131 4869
rect 135 4865 136 4869
rect 130 4864 136 4865
rect 386 4869 392 4870
rect 386 4865 387 4869
rect 391 4865 392 4869
rect 386 4864 392 4865
rect 706 4869 712 4870
rect 706 4865 707 4869
rect 711 4865 712 4869
rect 706 4864 712 4865
rect 1058 4869 1064 4870
rect 1058 4865 1059 4869
rect 1063 4865 1064 4869
rect 1058 4864 1064 4865
rect 1434 4869 1440 4870
rect 1434 4865 1435 4869
rect 1439 4865 1440 4869
rect 1434 4864 1440 4865
rect 1786 4869 1792 4870
rect 1786 4865 1787 4869
rect 1791 4865 1792 4869
rect 1786 4864 1792 4865
rect 1934 4868 1940 4869
rect 1934 4864 1935 4868
rect 1939 4864 1940 4868
rect 110 4863 116 4864
rect 112 4791 114 4863
rect 132 4791 134 4864
rect 388 4791 390 4864
rect 708 4791 710 4864
rect 1060 4791 1062 4864
rect 1436 4791 1438 4864
rect 1788 4791 1790 4864
rect 1934 4863 1940 4864
rect 1936 4791 1938 4863
rect 1976 4831 1978 4882
rect 2024 4831 2026 4883
rect 2160 4831 2162 4883
rect 2328 4831 2330 4883
rect 2496 4831 2498 4883
rect 2672 4831 2674 4883
rect 2848 4831 2850 4883
rect 3016 4831 3018 4883
rect 3184 4831 3186 4883
rect 3352 4831 3354 4883
rect 3528 4831 3530 4883
rect 3680 4831 3682 4883
rect 3798 4882 3804 4883
rect 3800 4831 3802 4882
rect 3840 4853 3842 4913
rect 3838 4852 3844 4853
rect 4676 4852 4678 4913
rect 4828 4852 4830 4913
rect 4988 4852 4990 4913
rect 5156 4852 5158 4913
rect 5324 4852 5326 4913
rect 5500 4852 5502 4913
rect 5664 4853 5666 4913
rect 5662 4852 5668 4853
rect 3838 4848 3839 4852
rect 3843 4848 3844 4852
rect 3838 4847 3844 4848
rect 4674 4851 4680 4852
rect 4674 4847 4675 4851
rect 4679 4847 4680 4851
rect 4674 4846 4680 4847
rect 4826 4851 4832 4852
rect 4826 4847 4827 4851
rect 4831 4847 4832 4851
rect 4826 4846 4832 4847
rect 4986 4851 4992 4852
rect 4986 4847 4987 4851
rect 4991 4847 4992 4851
rect 4986 4846 4992 4847
rect 5154 4851 5160 4852
rect 5154 4847 5155 4851
rect 5159 4847 5160 4851
rect 5154 4846 5160 4847
rect 5322 4851 5328 4852
rect 5322 4847 5323 4851
rect 5327 4847 5328 4851
rect 5322 4846 5328 4847
rect 5498 4851 5504 4852
rect 5498 4847 5499 4851
rect 5503 4847 5504 4851
rect 5662 4848 5663 4852
rect 5667 4848 5668 4852
rect 5662 4847 5668 4848
rect 5498 4846 5504 4847
rect 4702 4836 4708 4837
rect 3838 4835 3844 4836
rect 3838 4831 3839 4835
rect 3843 4831 3844 4835
rect 4702 4832 4703 4836
rect 4707 4832 4708 4836
rect 4702 4831 4708 4832
rect 4854 4836 4860 4837
rect 4854 4832 4855 4836
rect 4859 4832 4860 4836
rect 4854 4831 4860 4832
rect 5014 4836 5020 4837
rect 5014 4832 5015 4836
rect 5019 4832 5020 4836
rect 5014 4831 5020 4832
rect 5182 4836 5188 4837
rect 5182 4832 5183 4836
rect 5187 4832 5188 4836
rect 5182 4831 5188 4832
rect 5350 4836 5356 4837
rect 5350 4832 5351 4836
rect 5355 4832 5356 4836
rect 5350 4831 5356 4832
rect 5526 4836 5532 4837
rect 5526 4832 5527 4836
rect 5531 4832 5532 4836
rect 5526 4831 5532 4832
rect 5662 4835 5668 4836
rect 5662 4831 5663 4835
rect 5667 4831 5668 4835
rect 1975 4830 1979 4831
rect 1975 4825 1979 4826
rect 2023 4830 2027 4831
rect 2023 4825 2027 4826
rect 2159 4830 2163 4831
rect 2159 4825 2163 4826
rect 2327 4830 2331 4831
rect 2327 4825 2331 4826
rect 2391 4830 2395 4831
rect 2391 4825 2395 4826
rect 2495 4830 2499 4831
rect 2495 4825 2499 4826
rect 2527 4830 2531 4831
rect 2527 4825 2531 4826
rect 2663 4830 2667 4831
rect 2663 4825 2667 4826
rect 2671 4830 2675 4831
rect 2671 4825 2675 4826
rect 2807 4830 2811 4831
rect 2807 4825 2811 4826
rect 2847 4830 2851 4831
rect 2847 4825 2851 4826
rect 2951 4830 2955 4831
rect 2951 4825 2955 4826
rect 3015 4830 3019 4831
rect 3015 4825 3019 4826
rect 3095 4830 3099 4831
rect 3095 4825 3099 4826
rect 3183 4830 3187 4831
rect 3183 4825 3187 4826
rect 3239 4830 3243 4831
rect 3239 4825 3243 4826
rect 3351 4830 3355 4831
rect 3351 4825 3355 4826
rect 3383 4830 3387 4831
rect 3383 4825 3387 4826
rect 3527 4830 3531 4831
rect 3527 4825 3531 4826
rect 3679 4830 3683 4831
rect 3679 4825 3683 4826
rect 3799 4830 3803 4831
rect 3838 4830 3844 4831
rect 3799 4825 3803 4826
rect 1976 4802 1978 4825
rect 1974 4801 1980 4802
rect 2392 4801 2394 4825
rect 2528 4801 2530 4825
rect 2664 4801 2666 4825
rect 2808 4801 2810 4825
rect 2952 4801 2954 4825
rect 3096 4801 3098 4825
rect 3240 4801 3242 4825
rect 3384 4801 3386 4825
rect 3528 4801 3530 4825
rect 3800 4802 3802 4825
rect 3798 4801 3804 4802
rect 1974 4797 1975 4801
rect 1979 4797 1980 4801
rect 1974 4796 1980 4797
rect 2390 4800 2396 4801
rect 2390 4796 2391 4800
rect 2395 4796 2396 4800
rect 2390 4795 2396 4796
rect 2526 4800 2532 4801
rect 2526 4796 2527 4800
rect 2531 4796 2532 4800
rect 2526 4795 2532 4796
rect 2662 4800 2668 4801
rect 2662 4796 2663 4800
rect 2667 4796 2668 4800
rect 2662 4795 2668 4796
rect 2806 4800 2812 4801
rect 2806 4796 2807 4800
rect 2811 4796 2812 4800
rect 2806 4795 2812 4796
rect 2950 4800 2956 4801
rect 2950 4796 2951 4800
rect 2955 4796 2956 4800
rect 2950 4795 2956 4796
rect 3094 4800 3100 4801
rect 3094 4796 3095 4800
rect 3099 4796 3100 4800
rect 3094 4795 3100 4796
rect 3238 4800 3244 4801
rect 3238 4796 3239 4800
rect 3243 4796 3244 4800
rect 3238 4795 3244 4796
rect 3382 4800 3388 4801
rect 3382 4796 3383 4800
rect 3387 4796 3388 4800
rect 3382 4795 3388 4796
rect 3526 4800 3532 4801
rect 3526 4796 3527 4800
rect 3531 4796 3532 4800
rect 3798 4797 3799 4801
rect 3803 4797 3804 4801
rect 3798 4796 3804 4797
rect 3526 4795 3532 4796
rect 111 4790 115 4791
rect 111 4785 115 4786
rect 131 4790 135 4791
rect 131 4785 135 4786
rect 267 4790 271 4791
rect 267 4785 271 4786
rect 387 4790 391 4791
rect 387 4785 391 4786
rect 403 4790 407 4791
rect 403 4785 407 4786
rect 539 4790 543 4791
rect 539 4785 543 4786
rect 675 4790 679 4791
rect 675 4785 679 4786
rect 707 4790 711 4791
rect 707 4785 711 4786
rect 1059 4790 1063 4791
rect 1059 4785 1063 4786
rect 1435 4790 1439 4791
rect 1435 4785 1439 4786
rect 1787 4790 1791 4791
rect 1787 4785 1791 4786
rect 1935 4790 1939 4791
rect 3840 4787 3842 4830
rect 4704 4787 4706 4831
rect 4856 4787 4858 4831
rect 5016 4787 5018 4831
rect 5184 4787 5186 4831
rect 5352 4787 5354 4831
rect 5528 4787 5530 4831
rect 5662 4830 5668 4831
rect 5664 4787 5666 4830
rect 3839 4786 3843 4787
rect 1935 4785 1939 4786
rect 2362 4785 2368 4786
rect 112 4725 114 4785
rect 110 4724 116 4725
rect 132 4724 134 4785
rect 268 4724 270 4785
rect 404 4724 406 4785
rect 540 4724 542 4785
rect 676 4724 678 4785
rect 1936 4725 1938 4785
rect 1974 4784 1980 4785
rect 1974 4780 1975 4784
rect 1979 4780 1980 4784
rect 2362 4781 2363 4785
rect 2367 4781 2368 4785
rect 2362 4780 2368 4781
rect 2498 4785 2504 4786
rect 2498 4781 2499 4785
rect 2503 4781 2504 4785
rect 2498 4780 2504 4781
rect 2634 4785 2640 4786
rect 2634 4781 2635 4785
rect 2639 4781 2640 4785
rect 2634 4780 2640 4781
rect 2778 4785 2784 4786
rect 2778 4781 2779 4785
rect 2783 4781 2784 4785
rect 2778 4780 2784 4781
rect 2922 4785 2928 4786
rect 2922 4781 2923 4785
rect 2927 4781 2928 4785
rect 2922 4780 2928 4781
rect 3066 4785 3072 4786
rect 3066 4781 3067 4785
rect 3071 4781 3072 4785
rect 3066 4780 3072 4781
rect 3210 4785 3216 4786
rect 3210 4781 3211 4785
rect 3215 4781 3216 4785
rect 3210 4780 3216 4781
rect 3354 4785 3360 4786
rect 3354 4781 3355 4785
rect 3359 4781 3360 4785
rect 3354 4780 3360 4781
rect 3498 4785 3504 4786
rect 3498 4781 3499 4785
rect 3503 4781 3504 4785
rect 3498 4780 3504 4781
rect 3798 4784 3804 4785
rect 3798 4780 3799 4784
rect 3803 4780 3804 4784
rect 3839 4781 3843 4782
rect 4703 4786 4707 4787
rect 4703 4781 4707 4782
rect 4855 4786 4859 4787
rect 4855 4781 4859 4782
rect 4991 4786 4995 4787
rect 4991 4781 4995 4782
rect 5015 4786 5019 4787
rect 5015 4781 5019 4782
rect 5127 4786 5131 4787
rect 5127 4781 5131 4782
rect 5183 4786 5187 4787
rect 5183 4781 5187 4782
rect 5263 4786 5267 4787
rect 5263 4781 5267 4782
rect 5351 4786 5355 4787
rect 5351 4781 5355 4782
rect 5399 4786 5403 4787
rect 5399 4781 5403 4782
rect 5527 4786 5531 4787
rect 5527 4781 5531 4782
rect 5535 4786 5539 4787
rect 5535 4781 5539 4782
rect 5663 4786 5667 4787
rect 5663 4781 5667 4782
rect 1974 4779 1980 4780
rect 1934 4724 1940 4725
rect 110 4720 111 4724
rect 115 4720 116 4724
rect 110 4719 116 4720
rect 130 4723 136 4724
rect 130 4719 131 4723
rect 135 4719 136 4723
rect 130 4718 136 4719
rect 266 4723 272 4724
rect 266 4719 267 4723
rect 271 4719 272 4723
rect 266 4718 272 4719
rect 402 4723 408 4724
rect 402 4719 403 4723
rect 407 4719 408 4723
rect 402 4718 408 4719
rect 538 4723 544 4724
rect 538 4719 539 4723
rect 543 4719 544 4723
rect 538 4718 544 4719
rect 674 4723 680 4724
rect 674 4719 675 4723
rect 679 4719 680 4723
rect 1934 4720 1935 4724
rect 1939 4720 1940 4724
rect 1934 4719 1940 4720
rect 674 4718 680 4719
rect 1976 4711 1978 4779
rect 2364 4711 2366 4780
rect 2500 4711 2502 4780
rect 2636 4711 2638 4780
rect 2780 4711 2782 4780
rect 2924 4711 2926 4780
rect 3068 4711 3070 4780
rect 3212 4711 3214 4780
rect 3356 4711 3358 4780
rect 3500 4711 3502 4780
rect 3798 4779 3804 4780
rect 3800 4711 3802 4779
rect 3840 4758 3842 4781
rect 3838 4757 3844 4758
rect 4856 4757 4858 4781
rect 4992 4757 4994 4781
rect 5128 4757 5130 4781
rect 5264 4757 5266 4781
rect 5400 4757 5402 4781
rect 5536 4757 5538 4781
rect 5664 4758 5666 4781
rect 5662 4757 5668 4758
rect 3838 4753 3839 4757
rect 3843 4753 3844 4757
rect 3838 4752 3844 4753
rect 4854 4756 4860 4757
rect 4854 4752 4855 4756
rect 4859 4752 4860 4756
rect 4854 4751 4860 4752
rect 4990 4756 4996 4757
rect 4990 4752 4991 4756
rect 4995 4752 4996 4756
rect 4990 4751 4996 4752
rect 5126 4756 5132 4757
rect 5126 4752 5127 4756
rect 5131 4752 5132 4756
rect 5126 4751 5132 4752
rect 5262 4756 5268 4757
rect 5262 4752 5263 4756
rect 5267 4752 5268 4756
rect 5262 4751 5268 4752
rect 5398 4756 5404 4757
rect 5398 4752 5399 4756
rect 5403 4752 5404 4756
rect 5398 4751 5404 4752
rect 5534 4756 5540 4757
rect 5534 4752 5535 4756
rect 5539 4752 5540 4756
rect 5662 4753 5663 4757
rect 5667 4753 5668 4757
rect 5662 4752 5668 4753
rect 5534 4751 5540 4752
rect 4826 4741 4832 4742
rect 3838 4740 3844 4741
rect 3838 4736 3839 4740
rect 3843 4736 3844 4740
rect 4826 4737 4827 4741
rect 4831 4737 4832 4741
rect 4826 4736 4832 4737
rect 4962 4741 4968 4742
rect 4962 4737 4963 4741
rect 4967 4737 4968 4741
rect 4962 4736 4968 4737
rect 5098 4741 5104 4742
rect 5098 4737 5099 4741
rect 5103 4737 5104 4741
rect 5098 4736 5104 4737
rect 5234 4741 5240 4742
rect 5234 4737 5235 4741
rect 5239 4737 5240 4741
rect 5234 4736 5240 4737
rect 5370 4741 5376 4742
rect 5370 4737 5371 4741
rect 5375 4737 5376 4741
rect 5370 4736 5376 4737
rect 5506 4741 5512 4742
rect 5506 4737 5507 4741
rect 5511 4737 5512 4741
rect 5506 4736 5512 4737
rect 5662 4740 5668 4741
rect 5662 4736 5663 4740
rect 5667 4736 5668 4740
rect 3838 4735 3844 4736
rect 1975 4710 1979 4711
rect 158 4708 164 4709
rect 110 4707 116 4708
rect 110 4703 111 4707
rect 115 4703 116 4707
rect 158 4704 159 4708
rect 163 4704 164 4708
rect 158 4703 164 4704
rect 294 4708 300 4709
rect 294 4704 295 4708
rect 299 4704 300 4708
rect 294 4703 300 4704
rect 430 4708 436 4709
rect 430 4704 431 4708
rect 435 4704 436 4708
rect 430 4703 436 4704
rect 566 4708 572 4709
rect 566 4704 567 4708
rect 571 4704 572 4708
rect 566 4703 572 4704
rect 702 4708 708 4709
rect 702 4704 703 4708
rect 707 4704 708 4708
rect 702 4703 708 4704
rect 1934 4707 1940 4708
rect 1934 4703 1935 4707
rect 1939 4703 1940 4707
rect 1975 4705 1979 4706
rect 1995 4710 1999 4711
rect 1995 4705 1999 4706
rect 2131 4710 2135 4711
rect 2131 4705 2135 4706
rect 2267 4710 2271 4711
rect 2267 4705 2271 4706
rect 2363 4710 2367 4711
rect 2363 4705 2367 4706
rect 2427 4710 2431 4711
rect 2427 4705 2431 4706
rect 2499 4710 2503 4711
rect 2499 4705 2503 4706
rect 2587 4710 2591 4711
rect 2587 4705 2591 4706
rect 2635 4710 2639 4711
rect 2635 4705 2639 4706
rect 2747 4710 2751 4711
rect 2747 4705 2751 4706
rect 2779 4710 2783 4711
rect 2779 4705 2783 4706
rect 2907 4710 2911 4711
rect 2907 4705 2911 4706
rect 2923 4710 2927 4711
rect 2923 4705 2927 4706
rect 3067 4710 3071 4711
rect 3067 4705 3071 4706
rect 3211 4710 3215 4711
rect 3211 4705 3215 4706
rect 3235 4710 3239 4711
rect 3235 4705 3239 4706
rect 3355 4710 3359 4711
rect 3355 4705 3359 4706
rect 3499 4710 3503 4711
rect 3499 4705 3503 4706
rect 3799 4710 3803 4711
rect 3799 4705 3803 4706
rect 110 4702 116 4703
rect 112 4675 114 4702
rect 160 4675 162 4703
rect 296 4675 298 4703
rect 432 4675 434 4703
rect 568 4675 570 4703
rect 704 4675 706 4703
rect 1934 4702 1940 4703
rect 1936 4675 1938 4702
rect 111 4674 115 4675
rect 111 4669 115 4670
rect 159 4674 163 4675
rect 159 4669 163 4670
rect 295 4674 299 4675
rect 295 4669 299 4670
rect 431 4674 435 4675
rect 431 4669 435 4670
rect 567 4674 571 4675
rect 567 4669 571 4670
rect 703 4674 707 4675
rect 703 4669 707 4670
rect 1935 4674 1939 4675
rect 1935 4669 1939 4670
rect 112 4646 114 4669
rect 110 4645 116 4646
rect 160 4645 162 4669
rect 296 4645 298 4669
rect 432 4645 434 4669
rect 568 4645 570 4669
rect 704 4645 706 4669
rect 1936 4646 1938 4669
rect 1934 4645 1940 4646
rect 1976 4645 1978 4705
rect 110 4641 111 4645
rect 115 4641 116 4645
rect 110 4640 116 4641
rect 158 4644 164 4645
rect 158 4640 159 4644
rect 163 4640 164 4644
rect 158 4639 164 4640
rect 294 4644 300 4645
rect 294 4640 295 4644
rect 299 4640 300 4644
rect 294 4639 300 4640
rect 430 4644 436 4645
rect 430 4640 431 4644
rect 435 4640 436 4644
rect 430 4639 436 4640
rect 566 4644 572 4645
rect 566 4640 567 4644
rect 571 4640 572 4644
rect 566 4639 572 4640
rect 702 4644 708 4645
rect 702 4640 703 4644
rect 707 4640 708 4644
rect 1934 4641 1935 4645
rect 1939 4641 1940 4645
rect 1934 4640 1940 4641
rect 1974 4644 1980 4645
rect 1996 4644 1998 4705
rect 2132 4644 2134 4705
rect 2268 4644 2270 4705
rect 2428 4644 2430 4705
rect 2588 4644 2590 4705
rect 2748 4644 2750 4705
rect 2908 4644 2910 4705
rect 3068 4644 3070 4705
rect 3236 4644 3238 4705
rect 3800 4645 3802 4705
rect 3840 4655 3842 4735
rect 4828 4655 4830 4736
rect 4964 4655 4966 4736
rect 5100 4655 5102 4736
rect 5236 4655 5238 4736
rect 5372 4655 5374 4736
rect 5508 4655 5510 4736
rect 5662 4735 5668 4736
rect 5664 4655 5666 4735
rect 3839 4654 3843 4655
rect 3839 4649 3843 4650
rect 4715 4654 4719 4655
rect 4715 4649 4719 4650
rect 4827 4654 4831 4655
rect 4827 4649 4831 4650
rect 4859 4654 4863 4655
rect 4859 4649 4863 4650
rect 4963 4654 4967 4655
rect 4963 4649 4967 4650
rect 5011 4654 5015 4655
rect 5011 4649 5015 4650
rect 5099 4654 5103 4655
rect 5099 4649 5103 4650
rect 5171 4654 5175 4655
rect 5171 4649 5175 4650
rect 5235 4654 5239 4655
rect 5235 4649 5239 4650
rect 5339 4654 5343 4655
rect 5339 4649 5343 4650
rect 5371 4654 5375 4655
rect 5371 4649 5375 4650
rect 5507 4654 5511 4655
rect 5507 4649 5511 4650
rect 5515 4654 5519 4655
rect 5515 4649 5519 4650
rect 5663 4654 5667 4655
rect 5663 4649 5667 4650
rect 3798 4644 3804 4645
rect 1974 4640 1975 4644
rect 1979 4640 1980 4644
rect 702 4639 708 4640
rect 1974 4639 1980 4640
rect 1994 4643 2000 4644
rect 1994 4639 1995 4643
rect 1999 4639 2000 4643
rect 1994 4638 2000 4639
rect 2130 4643 2136 4644
rect 2130 4639 2131 4643
rect 2135 4639 2136 4643
rect 2130 4638 2136 4639
rect 2266 4643 2272 4644
rect 2266 4639 2267 4643
rect 2271 4639 2272 4643
rect 2266 4638 2272 4639
rect 2426 4643 2432 4644
rect 2426 4639 2427 4643
rect 2431 4639 2432 4643
rect 2426 4638 2432 4639
rect 2586 4643 2592 4644
rect 2586 4639 2587 4643
rect 2591 4639 2592 4643
rect 2586 4638 2592 4639
rect 2746 4643 2752 4644
rect 2746 4639 2747 4643
rect 2751 4639 2752 4643
rect 2746 4638 2752 4639
rect 2906 4643 2912 4644
rect 2906 4639 2907 4643
rect 2911 4639 2912 4643
rect 2906 4638 2912 4639
rect 3066 4643 3072 4644
rect 3066 4639 3067 4643
rect 3071 4639 3072 4643
rect 3066 4638 3072 4639
rect 3234 4643 3240 4644
rect 3234 4639 3235 4643
rect 3239 4639 3240 4643
rect 3798 4640 3799 4644
rect 3803 4640 3804 4644
rect 3798 4639 3804 4640
rect 3234 4638 3240 4639
rect 130 4629 136 4630
rect 110 4628 116 4629
rect 110 4624 111 4628
rect 115 4624 116 4628
rect 130 4625 131 4629
rect 135 4625 136 4629
rect 130 4624 136 4625
rect 266 4629 272 4630
rect 266 4625 267 4629
rect 271 4625 272 4629
rect 266 4624 272 4625
rect 402 4629 408 4630
rect 402 4625 403 4629
rect 407 4625 408 4629
rect 402 4624 408 4625
rect 538 4629 544 4630
rect 538 4625 539 4629
rect 543 4625 544 4629
rect 538 4624 544 4625
rect 674 4629 680 4630
rect 674 4625 675 4629
rect 679 4625 680 4629
rect 674 4624 680 4625
rect 1934 4628 1940 4629
rect 2022 4628 2028 4629
rect 1934 4624 1935 4628
rect 1939 4624 1940 4628
rect 110 4623 116 4624
rect 112 4551 114 4623
rect 132 4551 134 4624
rect 268 4551 270 4624
rect 404 4551 406 4624
rect 540 4551 542 4624
rect 676 4551 678 4624
rect 1934 4623 1940 4624
rect 1974 4627 1980 4628
rect 1974 4623 1975 4627
rect 1979 4623 1980 4627
rect 2022 4624 2023 4628
rect 2027 4624 2028 4628
rect 2022 4623 2028 4624
rect 2158 4628 2164 4629
rect 2158 4624 2159 4628
rect 2163 4624 2164 4628
rect 2158 4623 2164 4624
rect 2294 4628 2300 4629
rect 2294 4624 2295 4628
rect 2299 4624 2300 4628
rect 2294 4623 2300 4624
rect 2454 4628 2460 4629
rect 2454 4624 2455 4628
rect 2459 4624 2460 4628
rect 2454 4623 2460 4624
rect 2614 4628 2620 4629
rect 2614 4624 2615 4628
rect 2619 4624 2620 4628
rect 2614 4623 2620 4624
rect 2774 4628 2780 4629
rect 2774 4624 2775 4628
rect 2779 4624 2780 4628
rect 2774 4623 2780 4624
rect 2934 4628 2940 4629
rect 2934 4624 2935 4628
rect 2939 4624 2940 4628
rect 2934 4623 2940 4624
rect 3094 4628 3100 4629
rect 3094 4624 3095 4628
rect 3099 4624 3100 4628
rect 3094 4623 3100 4624
rect 3262 4628 3268 4629
rect 3262 4624 3263 4628
rect 3267 4624 3268 4628
rect 3262 4623 3268 4624
rect 3798 4627 3804 4628
rect 3798 4623 3799 4627
rect 3803 4623 3804 4627
rect 1936 4551 1938 4623
rect 1974 4622 1980 4623
rect 1976 4599 1978 4622
rect 2024 4599 2026 4623
rect 2160 4599 2162 4623
rect 2296 4599 2298 4623
rect 2456 4599 2458 4623
rect 2616 4599 2618 4623
rect 2776 4599 2778 4623
rect 2936 4599 2938 4623
rect 3096 4599 3098 4623
rect 3264 4599 3266 4623
rect 3798 4622 3804 4623
rect 3800 4599 3802 4622
rect 1975 4598 1979 4599
rect 1975 4593 1979 4594
rect 2023 4598 2027 4599
rect 2023 4593 2027 4594
rect 2159 4598 2163 4599
rect 2159 4593 2163 4594
rect 2175 4598 2179 4599
rect 2175 4593 2179 4594
rect 2295 4598 2299 4599
rect 2295 4593 2299 4594
rect 2351 4598 2355 4599
rect 2351 4593 2355 4594
rect 2455 4598 2459 4599
rect 2455 4593 2459 4594
rect 2527 4598 2531 4599
rect 2527 4593 2531 4594
rect 2615 4598 2619 4599
rect 2615 4593 2619 4594
rect 2695 4598 2699 4599
rect 2695 4593 2699 4594
rect 2775 4598 2779 4599
rect 2775 4593 2779 4594
rect 2871 4598 2875 4599
rect 2871 4593 2875 4594
rect 2935 4598 2939 4599
rect 2935 4593 2939 4594
rect 3047 4598 3051 4599
rect 3047 4593 3051 4594
rect 3095 4598 3099 4599
rect 3095 4593 3099 4594
rect 3263 4598 3267 4599
rect 3263 4593 3267 4594
rect 3799 4598 3803 4599
rect 3799 4593 3803 4594
rect 1976 4570 1978 4593
rect 1974 4569 1980 4570
rect 2024 4569 2026 4593
rect 2176 4569 2178 4593
rect 2352 4569 2354 4593
rect 2528 4569 2530 4593
rect 2696 4569 2698 4593
rect 2872 4569 2874 4593
rect 3048 4569 3050 4593
rect 3800 4570 3802 4593
rect 3840 4589 3842 4649
rect 3838 4588 3844 4589
rect 4716 4588 4718 4649
rect 4860 4588 4862 4649
rect 5012 4588 5014 4649
rect 5172 4588 5174 4649
rect 5340 4588 5342 4649
rect 5516 4588 5518 4649
rect 5664 4589 5666 4649
rect 5662 4588 5668 4589
rect 3838 4584 3839 4588
rect 3843 4584 3844 4588
rect 3838 4583 3844 4584
rect 4714 4587 4720 4588
rect 4714 4583 4715 4587
rect 4719 4583 4720 4587
rect 4714 4582 4720 4583
rect 4858 4587 4864 4588
rect 4858 4583 4859 4587
rect 4863 4583 4864 4587
rect 4858 4582 4864 4583
rect 5010 4587 5016 4588
rect 5010 4583 5011 4587
rect 5015 4583 5016 4587
rect 5010 4582 5016 4583
rect 5170 4587 5176 4588
rect 5170 4583 5171 4587
rect 5175 4583 5176 4587
rect 5170 4582 5176 4583
rect 5338 4587 5344 4588
rect 5338 4583 5339 4587
rect 5343 4583 5344 4587
rect 5338 4582 5344 4583
rect 5514 4587 5520 4588
rect 5514 4583 5515 4587
rect 5519 4583 5520 4587
rect 5662 4584 5663 4588
rect 5667 4584 5668 4588
rect 5662 4583 5668 4584
rect 5514 4582 5520 4583
rect 4742 4572 4748 4573
rect 3838 4571 3844 4572
rect 3798 4569 3804 4570
rect 1974 4565 1975 4569
rect 1979 4565 1980 4569
rect 1974 4564 1980 4565
rect 2022 4568 2028 4569
rect 2022 4564 2023 4568
rect 2027 4564 2028 4568
rect 2022 4563 2028 4564
rect 2174 4568 2180 4569
rect 2174 4564 2175 4568
rect 2179 4564 2180 4568
rect 2174 4563 2180 4564
rect 2350 4568 2356 4569
rect 2350 4564 2351 4568
rect 2355 4564 2356 4568
rect 2350 4563 2356 4564
rect 2526 4568 2532 4569
rect 2526 4564 2527 4568
rect 2531 4564 2532 4568
rect 2526 4563 2532 4564
rect 2694 4568 2700 4569
rect 2694 4564 2695 4568
rect 2699 4564 2700 4568
rect 2694 4563 2700 4564
rect 2870 4568 2876 4569
rect 2870 4564 2871 4568
rect 2875 4564 2876 4568
rect 2870 4563 2876 4564
rect 3046 4568 3052 4569
rect 3046 4564 3047 4568
rect 3051 4564 3052 4568
rect 3798 4565 3799 4569
rect 3803 4565 3804 4569
rect 3838 4567 3839 4571
rect 3843 4567 3844 4571
rect 4742 4568 4743 4572
rect 4747 4568 4748 4572
rect 4742 4567 4748 4568
rect 4886 4572 4892 4573
rect 4886 4568 4887 4572
rect 4891 4568 4892 4572
rect 4886 4567 4892 4568
rect 5038 4572 5044 4573
rect 5038 4568 5039 4572
rect 5043 4568 5044 4572
rect 5038 4567 5044 4568
rect 5198 4572 5204 4573
rect 5198 4568 5199 4572
rect 5203 4568 5204 4572
rect 5198 4567 5204 4568
rect 5366 4572 5372 4573
rect 5366 4568 5367 4572
rect 5371 4568 5372 4572
rect 5366 4567 5372 4568
rect 5542 4572 5548 4573
rect 5542 4568 5543 4572
rect 5547 4568 5548 4572
rect 5542 4567 5548 4568
rect 5662 4571 5668 4572
rect 5662 4567 5663 4571
rect 5667 4567 5668 4571
rect 3838 4566 3844 4567
rect 3798 4564 3804 4565
rect 3046 4563 3052 4564
rect 1994 4553 2000 4554
rect 1974 4552 1980 4553
rect 111 4550 115 4551
rect 111 4545 115 4546
rect 131 4550 135 4551
rect 131 4545 135 4546
rect 267 4550 271 4551
rect 267 4545 271 4546
rect 299 4550 303 4551
rect 299 4545 303 4546
rect 403 4550 407 4551
rect 403 4545 407 4546
rect 491 4550 495 4551
rect 491 4545 495 4546
rect 539 4550 543 4551
rect 539 4545 543 4546
rect 675 4550 679 4551
rect 675 4545 679 4546
rect 691 4550 695 4551
rect 691 4545 695 4546
rect 907 4550 911 4551
rect 907 4545 911 4546
rect 1123 4550 1127 4551
rect 1123 4545 1127 4546
rect 1347 4550 1351 4551
rect 1347 4545 1351 4546
rect 1579 4550 1583 4551
rect 1579 4545 1583 4546
rect 1787 4550 1791 4551
rect 1787 4545 1791 4546
rect 1935 4550 1939 4551
rect 1974 4548 1975 4552
rect 1979 4548 1980 4552
rect 1994 4549 1995 4553
rect 1999 4549 2000 4553
rect 1994 4548 2000 4549
rect 2146 4553 2152 4554
rect 2146 4549 2147 4553
rect 2151 4549 2152 4553
rect 2146 4548 2152 4549
rect 2322 4553 2328 4554
rect 2322 4549 2323 4553
rect 2327 4549 2328 4553
rect 2322 4548 2328 4549
rect 2498 4553 2504 4554
rect 2498 4549 2499 4553
rect 2503 4549 2504 4553
rect 2498 4548 2504 4549
rect 2666 4553 2672 4554
rect 2666 4549 2667 4553
rect 2671 4549 2672 4553
rect 2666 4548 2672 4549
rect 2842 4553 2848 4554
rect 2842 4549 2843 4553
rect 2847 4549 2848 4553
rect 2842 4548 2848 4549
rect 3018 4553 3024 4554
rect 3018 4549 3019 4553
rect 3023 4549 3024 4553
rect 3018 4548 3024 4549
rect 3798 4552 3804 4553
rect 3798 4548 3799 4552
rect 3803 4548 3804 4552
rect 1974 4547 1980 4548
rect 1935 4545 1939 4546
rect 112 4485 114 4545
rect 110 4484 116 4485
rect 300 4484 302 4545
rect 492 4484 494 4545
rect 692 4484 694 4545
rect 908 4484 910 4545
rect 1124 4484 1126 4545
rect 1348 4484 1350 4545
rect 1580 4484 1582 4545
rect 1788 4484 1790 4545
rect 1936 4485 1938 4545
rect 1934 4484 1940 4485
rect 110 4480 111 4484
rect 115 4480 116 4484
rect 110 4479 116 4480
rect 298 4483 304 4484
rect 298 4479 299 4483
rect 303 4479 304 4483
rect 298 4478 304 4479
rect 490 4483 496 4484
rect 490 4479 491 4483
rect 495 4479 496 4483
rect 490 4478 496 4479
rect 690 4483 696 4484
rect 690 4479 691 4483
rect 695 4479 696 4483
rect 690 4478 696 4479
rect 906 4483 912 4484
rect 906 4479 907 4483
rect 911 4479 912 4483
rect 906 4478 912 4479
rect 1122 4483 1128 4484
rect 1122 4479 1123 4483
rect 1127 4479 1128 4483
rect 1122 4478 1128 4479
rect 1346 4483 1352 4484
rect 1346 4479 1347 4483
rect 1351 4479 1352 4483
rect 1346 4478 1352 4479
rect 1578 4483 1584 4484
rect 1578 4479 1579 4483
rect 1583 4479 1584 4483
rect 1578 4478 1584 4479
rect 1786 4483 1792 4484
rect 1786 4479 1787 4483
rect 1791 4479 1792 4483
rect 1934 4480 1935 4484
rect 1939 4480 1940 4484
rect 1934 4479 1940 4480
rect 1786 4478 1792 4479
rect 326 4468 332 4469
rect 110 4467 116 4468
rect 110 4463 111 4467
rect 115 4463 116 4467
rect 326 4464 327 4468
rect 331 4464 332 4468
rect 326 4463 332 4464
rect 518 4468 524 4469
rect 518 4464 519 4468
rect 523 4464 524 4468
rect 518 4463 524 4464
rect 718 4468 724 4469
rect 718 4464 719 4468
rect 723 4464 724 4468
rect 718 4463 724 4464
rect 934 4468 940 4469
rect 934 4464 935 4468
rect 939 4464 940 4468
rect 934 4463 940 4464
rect 1150 4468 1156 4469
rect 1150 4464 1151 4468
rect 1155 4464 1156 4468
rect 1150 4463 1156 4464
rect 1374 4468 1380 4469
rect 1374 4464 1375 4468
rect 1379 4464 1380 4468
rect 1374 4463 1380 4464
rect 1606 4468 1612 4469
rect 1606 4464 1607 4468
rect 1611 4464 1612 4468
rect 1606 4463 1612 4464
rect 1814 4468 1820 4469
rect 1814 4464 1815 4468
rect 1819 4464 1820 4468
rect 1814 4463 1820 4464
rect 1934 4467 1940 4468
rect 1934 4463 1935 4467
rect 1939 4463 1940 4467
rect 110 4462 116 4463
rect 112 4439 114 4462
rect 328 4439 330 4463
rect 520 4439 522 4463
rect 720 4439 722 4463
rect 936 4439 938 4463
rect 1152 4439 1154 4463
rect 1376 4439 1378 4463
rect 1608 4439 1610 4463
rect 1816 4439 1818 4463
rect 1934 4462 1940 4463
rect 1936 4439 1938 4462
rect 1976 4447 1978 4547
rect 1996 4447 1998 4548
rect 2148 4447 2150 4548
rect 2324 4447 2326 4548
rect 2500 4447 2502 4548
rect 2668 4447 2670 4548
rect 2844 4447 2846 4548
rect 3020 4447 3022 4548
rect 3798 4547 3804 4548
rect 3800 4447 3802 4547
rect 3840 4519 3842 4566
rect 4744 4519 4746 4567
rect 4888 4519 4890 4567
rect 5040 4519 5042 4567
rect 5200 4519 5202 4567
rect 5368 4519 5370 4567
rect 5544 4519 5546 4567
rect 5662 4566 5668 4567
rect 5664 4519 5666 4566
rect 3839 4518 3843 4519
rect 3839 4513 3843 4514
rect 3887 4518 3891 4519
rect 3887 4513 3891 4514
rect 4063 4518 4067 4519
rect 4063 4513 4067 4514
rect 4279 4518 4283 4519
rect 4279 4513 4283 4514
rect 4503 4518 4507 4519
rect 4503 4513 4507 4514
rect 4743 4518 4747 4519
rect 4743 4513 4747 4514
rect 4751 4518 4755 4519
rect 4751 4513 4755 4514
rect 4887 4518 4891 4519
rect 4887 4513 4891 4514
rect 5007 4518 5011 4519
rect 5007 4513 5011 4514
rect 5039 4518 5043 4519
rect 5039 4513 5043 4514
rect 5199 4518 5203 4519
rect 5199 4513 5203 4514
rect 5271 4518 5275 4519
rect 5271 4513 5275 4514
rect 5367 4518 5371 4519
rect 5367 4513 5371 4514
rect 5543 4518 5547 4519
rect 5543 4513 5547 4514
rect 5663 4518 5667 4519
rect 5663 4513 5667 4514
rect 3840 4490 3842 4513
rect 3838 4489 3844 4490
rect 3888 4489 3890 4513
rect 4064 4489 4066 4513
rect 4280 4489 4282 4513
rect 4504 4489 4506 4513
rect 4752 4489 4754 4513
rect 5008 4489 5010 4513
rect 5272 4489 5274 4513
rect 5544 4489 5546 4513
rect 5664 4490 5666 4513
rect 5662 4489 5668 4490
rect 3838 4485 3839 4489
rect 3843 4485 3844 4489
rect 3838 4484 3844 4485
rect 3886 4488 3892 4489
rect 3886 4484 3887 4488
rect 3891 4484 3892 4488
rect 3886 4483 3892 4484
rect 4062 4488 4068 4489
rect 4062 4484 4063 4488
rect 4067 4484 4068 4488
rect 4062 4483 4068 4484
rect 4278 4488 4284 4489
rect 4278 4484 4279 4488
rect 4283 4484 4284 4488
rect 4278 4483 4284 4484
rect 4502 4488 4508 4489
rect 4502 4484 4503 4488
rect 4507 4484 4508 4488
rect 4502 4483 4508 4484
rect 4750 4488 4756 4489
rect 4750 4484 4751 4488
rect 4755 4484 4756 4488
rect 4750 4483 4756 4484
rect 5006 4488 5012 4489
rect 5006 4484 5007 4488
rect 5011 4484 5012 4488
rect 5006 4483 5012 4484
rect 5270 4488 5276 4489
rect 5270 4484 5271 4488
rect 5275 4484 5276 4488
rect 5270 4483 5276 4484
rect 5542 4488 5548 4489
rect 5542 4484 5543 4488
rect 5547 4484 5548 4488
rect 5662 4485 5663 4489
rect 5667 4485 5668 4489
rect 5662 4484 5668 4485
rect 5542 4483 5548 4484
rect 3858 4473 3864 4474
rect 3838 4472 3844 4473
rect 3838 4468 3839 4472
rect 3843 4468 3844 4472
rect 3858 4469 3859 4473
rect 3863 4469 3864 4473
rect 3858 4468 3864 4469
rect 4034 4473 4040 4474
rect 4034 4469 4035 4473
rect 4039 4469 4040 4473
rect 4034 4468 4040 4469
rect 4250 4473 4256 4474
rect 4250 4469 4251 4473
rect 4255 4469 4256 4473
rect 4250 4468 4256 4469
rect 4474 4473 4480 4474
rect 4474 4469 4475 4473
rect 4479 4469 4480 4473
rect 4474 4468 4480 4469
rect 4722 4473 4728 4474
rect 4722 4469 4723 4473
rect 4727 4469 4728 4473
rect 4722 4468 4728 4469
rect 4978 4473 4984 4474
rect 4978 4469 4979 4473
rect 4983 4469 4984 4473
rect 4978 4468 4984 4469
rect 5242 4473 5248 4474
rect 5242 4469 5243 4473
rect 5247 4469 5248 4473
rect 5242 4468 5248 4469
rect 5514 4473 5520 4474
rect 5514 4469 5515 4473
rect 5519 4469 5520 4473
rect 5514 4468 5520 4469
rect 5662 4472 5668 4473
rect 5662 4468 5663 4472
rect 5667 4468 5668 4472
rect 3838 4467 3844 4468
rect 1975 4446 1979 4447
rect 1975 4441 1979 4442
rect 1995 4446 1999 4447
rect 1995 4441 1999 4442
rect 2147 4446 2151 4447
rect 2147 4441 2151 4442
rect 2323 4446 2327 4447
rect 2323 4441 2327 4442
rect 2499 4446 2503 4447
rect 2499 4441 2503 4442
rect 2571 4446 2575 4447
rect 2571 4441 2575 4442
rect 2667 4446 2671 4447
rect 2667 4441 2671 4442
rect 2843 4446 2847 4447
rect 2843 4441 2847 4442
rect 3019 4446 3023 4447
rect 3019 4441 3023 4442
rect 3123 4446 3127 4447
rect 3123 4441 3127 4442
rect 3651 4446 3655 4447
rect 3651 4441 3655 4442
rect 3799 4446 3803 4447
rect 3799 4441 3803 4442
rect 111 4438 115 4439
rect 111 4433 115 4434
rect 327 4438 331 4439
rect 327 4433 331 4434
rect 519 4438 523 4439
rect 519 4433 523 4434
rect 559 4438 563 4439
rect 559 4433 563 4434
rect 719 4438 723 4439
rect 719 4433 723 4434
rect 887 4438 891 4439
rect 887 4433 891 4434
rect 935 4438 939 4439
rect 935 4433 939 4434
rect 1063 4438 1067 4439
rect 1063 4433 1067 4434
rect 1151 4438 1155 4439
rect 1151 4433 1155 4434
rect 1247 4438 1251 4439
rect 1247 4433 1251 4434
rect 1375 4438 1379 4439
rect 1375 4433 1379 4434
rect 1439 4438 1443 4439
rect 1439 4433 1443 4434
rect 1607 4438 1611 4439
rect 1607 4433 1611 4434
rect 1631 4438 1635 4439
rect 1631 4433 1635 4434
rect 1815 4438 1819 4439
rect 1815 4433 1819 4434
rect 1935 4438 1939 4439
rect 1935 4433 1939 4434
rect 112 4410 114 4433
rect 110 4409 116 4410
rect 560 4409 562 4433
rect 720 4409 722 4433
rect 888 4409 890 4433
rect 1064 4409 1066 4433
rect 1248 4409 1250 4433
rect 1440 4409 1442 4433
rect 1632 4409 1634 4433
rect 1816 4409 1818 4433
rect 1936 4410 1938 4433
rect 1934 4409 1940 4410
rect 110 4405 111 4409
rect 115 4405 116 4409
rect 110 4404 116 4405
rect 558 4408 564 4409
rect 558 4404 559 4408
rect 563 4404 564 4408
rect 558 4403 564 4404
rect 718 4408 724 4409
rect 718 4404 719 4408
rect 723 4404 724 4408
rect 718 4403 724 4404
rect 886 4408 892 4409
rect 886 4404 887 4408
rect 891 4404 892 4408
rect 886 4403 892 4404
rect 1062 4408 1068 4409
rect 1062 4404 1063 4408
rect 1067 4404 1068 4408
rect 1062 4403 1068 4404
rect 1246 4408 1252 4409
rect 1246 4404 1247 4408
rect 1251 4404 1252 4408
rect 1246 4403 1252 4404
rect 1438 4408 1444 4409
rect 1438 4404 1439 4408
rect 1443 4404 1444 4408
rect 1438 4403 1444 4404
rect 1630 4408 1636 4409
rect 1630 4404 1631 4408
rect 1635 4404 1636 4408
rect 1630 4403 1636 4404
rect 1814 4408 1820 4409
rect 1814 4404 1815 4408
rect 1819 4404 1820 4408
rect 1934 4405 1935 4409
rect 1939 4405 1940 4409
rect 1934 4404 1940 4405
rect 1814 4403 1820 4404
rect 530 4393 536 4394
rect 110 4392 116 4393
rect 110 4388 111 4392
rect 115 4388 116 4392
rect 530 4389 531 4393
rect 535 4389 536 4393
rect 530 4388 536 4389
rect 690 4393 696 4394
rect 690 4389 691 4393
rect 695 4389 696 4393
rect 690 4388 696 4389
rect 858 4393 864 4394
rect 858 4389 859 4393
rect 863 4389 864 4393
rect 858 4388 864 4389
rect 1034 4393 1040 4394
rect 1034 4389 1035 4393
rect 1039 4389 1040 4393
rect 1034 4388 1040 4389
rect 1218 4393 1224 4394
rect 1218 4389 1219 4393
rect 1223 4389 1224 4393
rect 1218 4388 1224 4389
rect 1410 4393 1416 4394
rect 1410 4389 1411 4393
rect 1415 4389 1416 4393
rect 1410 4388 1416 4389
rect 1602 4393 1608 4394
rect 1602 4389 1603 4393
rect 1607 4389 1608 4393
rect 1602 4388 1608 4389
rect 1786 4393 1792 4394
rect 1786 4389 1787 4393
rect 1791 4389 1792 4393
rect 1786 4388 1792 4389
rect 1934 4392 1940 4393
rect 1934 4388 1935 4392
rect 1939 4388 1940 4392
rect 110 4387 116 4388
rect 112 4319 114 4387
rect 532 4319 534 4388
rect 692 4319 694 4388
rect 860 4319 862 4388
rect 1036 4319 1038 4388
rect 1220 4319 1222 4388
rect 1412 4319 1414 4388
rect 1604 4319 1606 4388
rect 1788 4319 1790 4388
rect 1934 4387 1940 4388
rect 1936 4319 1938 4387
rect 1976 4381 1978 4441
rect 1974 4380 1980 4381
rect 2572 4380 2574 4441
rect 3124 4380 3126 4441
rect 3652 4380 3654 4441
rect 3800 4381 3802 4441
rect 3840 4407 3842 4467
rect 3860 4407 3862 4468
rect 4036 4407 4038 4468
rect 4252 4407 4254 4468
rect 4476 4407 4478 4468
rect 4724 4407 4726 4468
rect 4980 4407 4982 4468
rect 5244 4407 5246 4468
rect 5516 4407 5518 4468
rect 5662 4467 5668 4468
rect 5664 4407 5666 4467
rect 3839 4406 3843 4407
rect 3839 4401 3843 4402
rect 3859 4406 3863 4407
rect 3859 4401 3863 4402
rect 3995 4406 3999 4407
rect 3995 4401 3999 4402
rect 4035 4406 4039 4407
rect 4035 4401 4039 4402
rect 4131 4406 4135 4407
rect 4131 4401 4135 4402
rect 4251 4406 4255 4407
rect 4251 4401 4255 4402
rect 4267 4406 4271 4407
rect 4267 4401 4271 4402
rect 4403 4406 4407 4407
rect 4403 4401 4407 4402
rect 4475 4406 4479 4407
rect 4475 4401 4479 4402
rect 4587 4406 4591 4407
rect 4587 4401 4591 4402
rect 4723 4406 4727 4407
rect 4723 4401 4727 4402
rect 4795 4406 4799 4407
rect 4795 4401 4799 4402
rect 4979 4406 4983 4407
rect 4979 4401 4983 4402
rect 5027 4406 5031 4407
rect 5027 4401 5031 4402
rect 5243 4406 5247 4407
rect 5243 4401 5247 4402
rect 5275 4406 5279 4407
rect 5275 4401 5279 4402
rect 5515 4406 5519 4407
rect 5515 4401 5519 4402
rect 5663 4406 5667 4407
rect 5663 4401 5667 4402
rect 3798 4380 3804 4381
rect 1974 4376 1975 4380
rect 1979 4376 1980 4380
rect 1974 4375 1980 4376
rect 2570 4379 2576 4380
rect 2570 4375 2571 4379
rect 2575 4375 2576 4379
rect 2570 4374 2576 4375
rect 3122 4379 3128 4380
rect 3122 4375 3123 4379
rect 3127 4375 3128 4379
rect 3122 4374 3128 4375
rect 3650 4379 3656 4380
rect 3650 4375 3651 4379
rect 3655 4375 3656 4379
rect 3798 4376 3799 4380
rect 3803 4376 3804 4380
rect 3798 4375 3804 4376
rect 3650 4374 3656 4375
rect 2598 4364 2604 4365
rect 1974 4363 1980 4364
rect 1974 4359 1975 4363
rect 1979 4359 1980 4363
rect 2598 4360 2599 4364
rect 2603 4360 2604 4364
rect 2598 4359 2604 4360
rect 3150 4364 3156 4365
rect 3150 4360 3151 4364
rect 3155 4360 3156 4364
rect 3150 4359 3156 4360
rect 3678 4364 3684 4365
rect 3678 4360 3679 4364
rect 3683 4360 3684 4364
rect 3678 4359 3684 4360
rect 3798 4363 3804 4364
rect 3798 4359 3799 4363
rect 3803 4359 3804 4363
rect 1974 4358 1980 4359
rect 1976 4331 1978 4358
rect 2600 4331 2602 4359
rect 3152 4331 3154 4359
rect 3680 4331 3682 4359
rect 3798 4358 3804 4359
rect 3800 4331 3802 4358
rect 3840 4341 3842 4401
rect 3838 4340 3844 4341
rect 3860 4340 3862 4401
rect 3996 4340 3998 4401
rect 4132 4340 4134 4401
rect 4268 4340 4270 4401
rect 4404 4340 4406 4401
rect 4588 4340 4590 4401
rect 4796 4340 4798 4401
rect 5028 4340 5030 4401
rect 5276 4340 5278 4401
rect 5516 4340 5518 4401
rect 5664 4341 5666 4401
rect 5662 4340 5668 4341
rect 3838 4336 3839 4340
rect 3843 4336 3844 4340
rect 3838 4335 3844 4336
rect 3858 4339 3864 4340
rect 3858 4335 3859 4339
rect 3863 4335 3864 4339
rect 3858 4334 3864 4335
rect 3994 4339 4000 4340
rect 3994 4335 3995 4339
rect 3999 4335 4000 4339
rect 3994 4334 4000 4335
rect 4130 4339 4136 4340
rect 4130 4335 4131 4339
rect 4135 4335 4136 4339
rect 4130 4334 4136 4335
rect 4266 4339 4272 4340
rect 4266 4335 4267 4339
rect 4271 4335 4272 4339
rect 4266 4334 4272 4335
rect 4402 4339 4408 4340
rect 4402 4335 4403 4339
rect 4407 4335 4408 4339
rect 4402 4334 4408 4335
rect 4586 4339 4592 4340
rect 4586 4335 4587 4339
rect 4591 4335 4592 4339
rect 4586 4334 4592 4335
rect 4794 4339 4800 4340
rect 4794 4335 4795 4339
rect 4799 4335 4800 4339
rect 4794 4334 4800 4335
rect 5026 4339 5032 4340
rect 5026 4335 5027 4339
rect 5031 4335 5032 4339
rect 5026 4334 5032 4335
rect 5274 4339 5280 4340
rect 5274 4335 5275 4339
rect 5279 4335 5280 4339
rect 5274 4334 5280 4335
rect 5514 4339 5520 4340
rect 5514 4335 5515 4339
rect 5519 4335 5520 4339
rect 5662 4336 5663 4340
rect 5667 4336 5668 4340
rect 5662 4335 5668 4336
rect 5514 4334 5520 4335
rect 1975 4330 1979 4331
rect 1975 4325 1979 4326
rect 2399 4330 2403 4331
rect 2399 4325 2403 4326
rect 2599 4330 2603 4331
rect 2599 4325 2603 4326
rect 2791 4330 2795 4331
rect 2791 4325 2795 4326
rect 2983 4330 2987 4331
rect 2983 4325 2987 4326
rect 3151 4330 3155 4331
rect 3151 4325 3155 4326
rect 3167 4330 3171 4331
rect 3167 4325 3171 4326
rect 3343 4330 3347 4331
rect 3343 4325 3347 4326
rect 3519 4330 3523 4331
rect 3519 4325 3523 4326
rect 3679 4330 3683 4331
rect 3679 4325 3683 4326
rect 3799 4330 3803 4331
rect 3799 4325 3803 4326
rect 111 4318 115 4319
rect 111 4313 115 4314
rect 531 4318 535 4319
rect 531 4313 535 4314
rect 691 4318 695 4319
rect 691 4313 695 4314
rect 747 4318 751 4319
rect 747 4313 751 4314
rect 859 4318 863 4319
rect 859 4313 863 4314
rect 883 4318 887 4319
rect 883 4313 887 4314
rect 1019 4318 1023 4319
rect 1019 4313 1023 4314
rect 1035 4318 1039 4319
rect 1035 4313 1039 4314
rect 1155 4318 1159 4319
rect 1155 4313 1159 4314
rect 1219 4318 1223 4319
rect 1219 4313 1223 4314
rect 1291 4318 1295 4319
rect 1291 4313 1295 4314
rect 1411 4318 1415 4319
rect 1411 4313 1415 4314
rect 1427 4318 1431 4319
rect 1427 4313 1431 4314
rect 1563 4318 1567 4319
rect 1563 4313 1567 4314
rect 1603 4318 1607 4319
rect 1603 4313 1607 4314
rect 1699 4318 1703 4319
rect 1699 4313 1703 4314
rect 1787 4318 1791 4319
rect 1787 4313 1791 4314
rect 1935 4318 1939 4319
rect 1935 4313 1939 4314
rect 112 4253 114 4313
rect 110 4252 116 4253
rect 748 4252 750 4313
rect 884 4252 886 4313
rect 1020 4252 1022 4313
rect 1156 4252 1158 4313
rect 1292 4252 1294 4313
rect 1428 4252 1430 4313
rect 1564 4252 1566 4313
rect 1700 4252 1702 4313
rect 1936 4253 1938 4313
rect 1976 4302 1978 4325
rect 1974 4301 1980 4302
rect 2400 4301 2402 4325
rect 2600 4301 2602 4325
rect 2792 4301 2794 4325
rect 2984 4301 2986 4325
rect 3168 4301 3170 4325
rect 3344 4301 3346 4325
rect 3520 4301 3522 4325
rect 3680 4301 3682 4325
rect 3800 4302 3802 4325
rect 3886 4324 3892 4325
rect 3838 4323 3844 4324
rect 3838 4319 3839 4323
rect 3843 4319 3844 4323
rect 3886 4320 3887 4324
rect 3891 4320 3892 4324
rect 3886 4319 3892 4320
rect 4022 4324 4028 4325
rect 4022 4320 4023 4324
rect 4027 4320 4028 4324
rect 4022 4319 4028 4320
rect 4158 4324 4164 4325
rect 4158 4320 4159 4324
rect 4163 4320 4164 4324
rect 4158 4319 4164 4320
rect 4294 4324 4300 4325
rect 4294 4320 4295 4324
rect 4299 4320 4300 4324
rect 4294 4319 4300 4320
rect 4430 4324 4436 4325
rect 4430 4320 4431 4324
rect 4435 4320 4436 4324
rect 4430 4319 4436 4320
rect 4614 4324 4620 4325
rect 4614 4320 4615 4324
rect 4619 4320 4620 4324
rect 4614 4319 4620 4320
rect 4822 4324 4828 4325
rect 4822 4320 4823 4324
rect 4827 4320 4828 4324
rect 4822 4319 4828 4320
rect 5054 4324 5060 4325
rect 5054 4320 5055 4324
rect 5059 4320 5060 4324
rect 5054 4319 5060 4320
rect 5302 4324 5308 4325
rect 5302 4320 5303 4324
rect 5307 4320 5308 4324
rect 5302 4319 5308 4320
rect 5542 4324 5548 4325
rect 5542 4320 5543 4324
rect 5547 4320 5548 4324
rect 5542 4319 5548 4320
rect 5662 4323 5668 4324
rect 5662 4319 5663 4323
rect 5667 4319 5668 4323
rect 3838 4318 3844 4319
rect 3798 4301 3804 4302
rect 1974 4297 1975 4301
rect 1979 4297 1980 4301
rect 1974 4296 1980 4297
rect 2398 4300 2404 4301
rect 2398 4296 2399 4300
rect 2403 4296 2404 4300
rect 2398 4295 2404 4296
rect 2598 4300 2604 4301
rect 2598 4296 2599 4300
rect 2603 4296 2604 4300
rect 2598 4295 2604 4296
rect 2790 4300 2796 4301
rect 2790 4296 2791 4300
rect 2795 4296 2796 4300
rect 2790 4295 2796 4296
rect 2982 4300 2988 4301
rect 2982 4296 2983 4300
rect 2987 4296 2988 4300
rect 2982 4295 2988 4296
rect 3166 4300 3172 4301
rect 3166 4296 3167 4300
rect 3171 4296 3172 4300
rect 3166 4295 3172 4296
rect 3342 4300 3348 4301
rect 3342 4296 3343 4300
rect 3347 4296 3348 4300
rect 3342 4295 3348 4296
rect 3518 4300 3524 4301
rect 3518 4296 3519 4300
rect 3523 4296 3524 4300
rect 3518 4295 3524 4296
rect 3678 4300 3684 4301
rect 3678 4296 3679 4300
rect 3683 4296 3684 4300
rect 3798 4297 3799 4301
rect 3803 4297 3804 4301
rect 3798 4296 3804 4297
rect 3678 4295 3684 4296
rect 3840 4295 3842 4318
rect 3888 4295 3890 4319
rect 4024 4295 4026 4319
rect 4160 4295 4162 4319
rect 4296 4295 4298 4319
rect 4432 4295 4434 4319
rect 4616 4295 4618 4319
rect 4824 4295 4826 4319
rect 5056 4295 5058 4319
rect 5304 4295 5306 4319
rect 5544 4295 5546 4319
rect 5662 4318 5668 4319
rect 5664 4295 5666 4318
rect 3839 4294 3843 4295
rect 3839 4289 3843 4290
rect 3887 4294 3891 4295
rect 3887 4289 3891 4290
rect 4023 4294 4027 4295
rect 4023 4289 4027 4290
rect 4047 4294 4051 4295
rect 4047 4289 4051 4290
rect 4159 4294 4163 4295
rect 4159 4289 4163 4290
rect 4223 4294 4227 4295
rect 4223 4289 4227 4290
rect 4295 4294 4299 4295
rect 4295 4289 4299 4290
rect 4431 4294 4435 4295
rect 4431 4289 4435 4290
rect 4615 4294 4619 4295
rect 4615 4289 4619 4290
rect 4679 4294 4683 4295
rect 4679 4289 4683 4290
rect 4823 4294 4827 4295
rect 4823 4289 4827 4290
rect 4959 4294 4963 4295
rect 4959 4289 4963 4290
rect 5055 4294 5059 4295
rect 5055 4289 5059 4290
rect 5255 4294 5259 4295
rect 5255 4289 5259 4290
rect 5303 4294 5307 4295
rect 5303 4289 5307 4290
rect 5543 4294 5547 4295
rect 5543 4289 5547 4290
rect 5663 4294 5667 4295
rect 5663 4289 5667 4290
rect 2370 4285 2376 4286
rect 1974 4284 1980 4285
rect 1974 4280 1975 4284
rect 1979 4280 1980 4284
rect 2370 4281 2371 4285
rect 2375 4281 2376 4285
rect 2370 4280 2376 4281
rect 2570 4285 2576 4286
rect 2570 4281 2571 4285
rect 2575 4281 2576 4285
rect 2570 4280 2576 4281
rect 2762 4285 2768 4286
rect 2762 4281 2763 4285
rect 2767 4281 2768 4285
rect 2762 4280 2768 4281
rect 2954 4285 2960 4286
rect 2954 4281 2955 4285
rect 2959 4281 2960 4285
rect 2954 4280 2960 4281
rect 3138 4285 3144 4286
rect 3138 4281 3139 4285
rect 3143 4281 3144 4285
rect 3138 4280 3144 4281
rect 3314 4285 3320 4286
rect 3314 4281 3315 4285
rect 3319 4281 3320 4285
rect 3314 4280 3320 4281
rect 3490 4285 3496 4286
rect 3490 4281 3491 4285
rect 3495 4281 3496 4285
rect 3490 4280 3496 4281
rect 3650 4285 3656 4286
rect 3650 4281 3651 4285
rect 3655 4281 3656 4285
rect 3650 4280 3656 4281
rect 3798 4284 3804 4285
rect 3798 4280 3799 4284
rect 3803 4280 3804 4284
rect 1974 4279 1980 4280
rect 1934 4252 1940 4253
rect 110 4248 111 4252
rect 115 4248 116 4252
rect 110 4247 116 4248
rect 746 4251 752 4252
rect 746 4247 747 4251
rect 751 4247 752 4251
rect 746 4246 752 4247
rect 882 4251 888 4252
rect 882 4247 883 4251
rect 887 4247 888 4251
rect 882 4246 888 4247
rect 1018 4251 1024 4252
rect 1018 4247 1019 4251
rect 1023 4247 1024 4251
rect 1018 4246 1024 4247
rect 1154 4251 1160 4252
rect 1154 4247 1155 4251
rect 1159 4247 1160 4251
rect 1154 4246 1160 4247
rect 1290 4251 1296 4252
rect 1290 4247 1291 4251
rect 1295 4247 1296 4251
rect 1290 4246 1296 4247
rect 1426 4251 1432 4252
rect 1426 4247 1427 4251
rect 1431 4247 1432 4251
rect 1426 4246 1432 4247
rect 1562 4251 1568 4252
rect 1562 4247 1563 4251
rect 1567 4247 1568 4251
rect 1562 4246 1568 4247
rect 1698 4251 1704 4252
rect 1698 4247 1699 4251
rect 1703 4247 1704 4251
rect 1934 4248 1935 4252
rect 1939 4248 1940 4252
rect 1934 4247 1940 4248
rect 1698 4246 1704 4247
rect 774 4236 780 4237
rect 110 4235 116 4236
rect 110 4231 111 4235
rect 115 4231 116 4235
rect 774 4232 775 4236
rect 779 4232 780 4236
rect 774 4231 780 4232
rect 910 4236 916 4237
rect 910 4232 911 4236
rect 915 4232 916 4236
rect 910 4231 916 4232
rect 1046 4236 1052 4237
rect 1046 4232 1047 4236
rect 1051 4232 1052 4236
rect 1046 4231 1052 4232
rect 1182 4236 1188 4237
rect 1182 4232 1183 4236
rect 1187 4232 1188 4236
rect 1182 4231 1188 4232
rect 1318 4236 1324 4237
rect 1318 4232 1319 4236
rect 1323 4232 1324 4236
rect 1318 4231 1324 4232
rect 1454 4236 1460 4237
rect 1454 4232 1455 4236
rect 1459 4232 1460 4236
rect 1454 4231 1460 4232
rect 1590 4236 1596 4237
rect 1590 4232 1591 4236
rect 1595 4232 1596 4236
rect 1590 4231 1596 4232
rect 1726 4236 1732 4237
rect 1726 4232 1727 4236
rect 1731 4232 1732 4236
rect 1726 4231 1732 4232
rect 1934 4235 1940 4236
rect 1934 4231 1935 4235
rect 1939 4231 1940 4235
rect 110 4230 116 4231
rect 112 4195 114 4230
rect 776 4195 778 4231
rect 912 4195 914 4231
rect 1048 4195 1050 4231
rect 1184 4195 1186 4231
rect 1320 4195 1322 4231
rect 1456 4195 1458 4231
rect 1592 4195 1594 4231
rect 1728 4195 1730 4231
rect 1934 4230 1940 4231
rect 1936 4195 1938 4230
rect 1976 4207 1978 4279
rect 2372 4207 2374 4280
rect 2572 4207 2574 4280
rect 2764 4207 2766 4280
rect 2956 4207 2958 4280
rect 3140 4207 3142 4280
rect 3316 4207 3318 4280
rect 3492 4207 3494 4280
rect 3652 4207 3654 4280
rect 3798 4279 3804 4280
rect 3800 4207 3802 4279
rect 3840 4266 3842 4289
rect 3838 4265 3844 4266
rect 4048 4265 4050 4289
rect 4224 4265 4226 4289
rect 4432 4265 4434 4289
rect 4680 4265 4682 4289
rect 4960 4265 4962 4289
rect 5256 4265 5258 4289
rect 5544 4265 5546 4289
rect 5664 4266 5666 4289
rect 5662 4265 5668 4266
rect 3838 4261 3839 4265
rect 3843 4261 3844 4265
rect 3838 4260 3844 4261
rect 4046 4264 4052 4265
rect 4046 4260 4047 4264
rect 4051 4260 4052 4264
rect 4046 4259 4052 4260
rect 4222 4264 4228 4265
rect 4222 4260 4223 4264
rect 4227 4260 4228 4264
rect 4222 4259 4228 4260
rect 4430 4264 4436 4265
rect 4430 4260 4431 4264
rect 4435 4260 4436 4264
rect 4430 4259 4436 4260
rect 4678 4264 4684 4265
rect 4678 4260 4679 4264
rect 4683 4260 4684 4264
rect 4678 4259 4684 4260
rect 4958 4264 4964 4265
rect 4958 4260 4959 4264
rect 4963 4260 4964 4264
rect 4958 4259 4964 4260
rect 5254 4264 5260 4265
rect 5254 4260 5255 4264
rect 5259 4260 5260 4264
rect 5254 4259 5260 4260
rect 5542 4264 5548 4265
rect 5542 4260 5543 4264
rect 5547 4260 5548 4264
rect 5662 4261 5663 4265
rect 5667 4261 5668 4265
rect 5662 4260 5668 4261
rect 5542 4259 5548 4260
rect 4018 4249 4024 4250
rect 3838 4248 3844 4249
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 4018 4245 4019 4249
rect 4023 4245 4024 4249
rect 4018 4244 4024 4245
rect 4194 4249 4200 4250
rect 4194 4245 4195 4249
rect 4199 4245 4200 4249
rect 4194 4244 4200 4245
rect 4402 4249 4408 4250
rect 4402 4245 4403 4249
rect 4407 4245 4408 4249
rect 4402 4244 4408 4245
rect 4650 4249 4656 4250
rect 4650 4245 4651 4249
rect 4655 4245 4656 4249
rect 4650 4244 4656 4245
rect 4930 4249 4936 4250
rect 4930 4245 4931 4249
rect 4935 4245 4936 4249
rect 4930 4244 4936 4245
rect 5226 4249 5232 4250
rect 5226 4245 5227 4249
rect 5231 4245 5232 4249
rect 5226 4244 5232 4245
rect 5514 4249 5520 4250
rect 5514 4245 5515 4249
rect 5519 4245 5520 4249
rect 5514 4244 5520 4245
rect 5662 4248 5668 4249
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 3838 4243 3844 4244
rect 1975 4206 1979 4207
rect 1975 4201 1979 4202
rect 2371 4206 2375 4207
rect 2371 4201 2375 4202
rect 2571 4206 2575 4207
rect 2571 4201 2575 4202
rect 2611 4206 2615 4207
rect 2611 4201 2615 4202
rect 2763 4206 2767 4207
rect 2763 4201 2767 4202
rect 2835 4206 2839 4207
rect 2835 4201 2839 4202
rect 2955 4206 2959 4207
rect 2955 4201 2959 4202
rect 3051 4206 3055 4207
rect 3051 4201 3055 4202
rect 3139 4206 3143 4207
rect 3139 4201 3143 4202
rect 3259 4206 3263 4207
rect 3259 4201 3263 4202
rect 3315 4206 3319 4207
rect 3315 4201 3319 4202
rect 3467 4206 3471 4207
rect 3467 4201 3471 4202
rect 3491 4206 3495 4207
rect 3491 4201 3495 4202
rect 3651 4206 3655 4207
rect 3651 4201 3655 4202
rect 3799 4206 3803 4207
rect 3799 4201 3803 4202
rect 111 4194 115 4195
rect 111 4189 115 4190
rect 727 4194 731 4195
rect 727 4189 731 4190
rect 775 4194 779 4195
rect 775 4189 779 4190
rect 863 4194 867 4195
rect 863 4189 867 4190
rect 911 4194 915 4195
rect 911 4189 915 4190
rect 999 4194 1003 4195
rect 999 4189 1003 4190
rect 1047 4194 1051 4195
rect 1047 4189 1051 4190
rect 1135 4194 1139 4195
rect 1135 4189 1139 4190
rect 1183 4194 1187 4195
rect 1183 4189 1187 4190
rect 1271 4194 1275 4195
rect 1271 4189 1275 4190
rect 1319 4194 1323 4195
rect 1319 4189 1323 4190
rect 1407 4194 1411 4195
rect 1407 4189 1411 4190
rect 1455 4194 1459 4195
rect 1455 4189 1459 4190
rect 1543 4194 1547 4195
rect 1543 4189 1547 4190
rect 1591 4194 1595 4195
rect 1591 4189 1595 4190
rect 1679 4194 1683 4195
rect 1679 4189 1683 4190
rect 1727 4194 1731 4195
rect 1727 4189 1731 4190
rect 1815 4194 1819 4195
rect 1815 4189 1819 4190
rect 1935 4194 1939 4195
rect 1935 4189 1939 4190
rect 112 4166 114 4189
rect 110 4165 116 4166
rect 728 4165 730 4189
rect 864 4165 866 4189
rect 1000 4165 1002 4189
rect 1136 4165 1138 4189
rect 1272 4165 1274 4189
rect 1408 4165 1410 4189
rect 1544 4165 1546 4189
rect 1680 4165 1682 4189
rect 1816 4165 1818 4189
rect 1936 4166 1938 4189
rect 1934 4165 1940 4166
rect 110 4161 111 4165
rect 115 4161 116 4165
rect 110 4160 116 4161
rect 726 4164 732 4165
rect 726 4160 727 4164
rect 731 4160 732 4164
rect 726 4159 732 4160
rect 862 4164 868 4165
rect 862 4160 863 4164
rect 867 4160 868 4164
rect 862 4159 868 4160
rect 998 4164 1004 4165
rect 998 4160 999 4164
rect 1003 4160 1004 4164
rect 998 4159 1004 4160
rect 1134 4164 1140 4165
rect 1134 4160 1135 4164
rect 1139 4160 1140 4164
rect 1134 4159 1140 4160
rect 1270 4164 1276 4165
rect 1270 4160 1271 4164
rect 1275 4160 1276 4164
rect 1270 4159 1276 4160
rect 1406 4164 1412 4165
rect 1406 4160 1407 4164
rect 1411 4160 1412 4164
rect 1406 4159 1412 4160
rect 1542 4164 1548 4165
rect 1542 4160 1543 4164
rect 1547 4160 1548 4164
rect 1542 4159 1548 4160
rect 1678 4164 1684 4165
rect 1678 4160 1679 4164
rect 1683 4160 1684 4164
rect 1678 4159 1684 4160
rect 1814 4164 1820 4165
rect 1814 4160 1815 4164
rect 1819 4160 1820 4164
rect 1934 4161 1935 4165
rect 1939 4161 1940 4165
rect 1934 4160 1940 4161
rect 1814 4159 1820 4160
rect 698 4149 704 4150
rect 110 4148 116 4149
rect 110 4144 111 4148
rect 115 4144 116 4148
rect 698 4145 699 4149
rect 703 4145 704 4149
rect 698 4144 704 4145
rect 834 4149 840 4150
rect 834 4145 835 4149
rect 839 4145 840 4149
rect 834 4144 840 4145
rect 970 4149 976 4150
rect 970 4145 971 4149
rect 975 4145 976 4149
rect 970 4144 976 4145
rect 1106 4149 1112 4150
rect 1106 4145 1107 4149
rect 1111 4145 1112 4149
rect 1106 4144 1112 4145
rect 1242 4149 1248 4150
rect 1242 4145 1243 4149
rect 1247 4145 1248 4149
rect 1242 4144 1248 4145
rect 1378 4149 1384 4150
rect 1378 4145 1379 4149
rect 1383 4145 1384 4149
rect 1378 4144 1384 4145
rect 1514 4149 1520 4150
rect 1514 4145 1515 4149
rect 1519 4145 1520 4149
rect 1514 4144 1520 4145
rect 1650 4149 1656 4150
rect 1650 4145 1651 4149
rect 1655 4145 1656 4149
rect 1650 4144 1656 4145
rect 1786 4149 1792 4150
rect 1786 4145 1787 4149
rect 1791 4145 1792 4149
rect 1786 4144 1792 4145
rect 1934 4148 1940 4149
rect 1934 4144 1935 4148
rect 1939 4144 1940 4148
rect 110 4143 116 4144
rect 112 4071 114 4143
rect 700 4071 702 4144
rect 836 4071 838 4144
rect 972 4071 974 4144
rect 1108 4071 1110 4144
rect 1244 4071 1246 4144
rect 1380 4071 1382 4144
rect 1516 4071 1518 4144
rect 1652 4071 1654 4144
rect 1788 4071 1790 4144
rect 1934 4143 1940 4144
rect 1936 4071 1938 4143
rect 1976 4141 1978 4201
rect 1974 4140 1980 4141
rect 2372 4140 2374 4201
rect 2612 4140 2614 4201
rect 2836 4140 2838 4201
rect 3052 4140 3054 4201
rect 3260 4140 3262 4201
rect 3468 4140 3470 4201
rect 3652 4140 3654 4201
rect 3800 4141 3802 4201
rect 3798 4140 3804 4141
rect 1974 4136 1975 4140
rect 1979 4136 1980 4140
rect 1974 4135 1980 4136
rect 2370 4139 2376 4140
rect 2370 4135 2371 4139
rect 2375 4135 2376 4139
rect 2370 4134 2376 4135
rect 2610 4139 2616 4140
rect 2610 4135 2611 4139
rect 2615 4135 2616 4139
rect 2610 4134 2616 4135
rect 2834 4139 2840 4140
rect 2834 4135 2835 4139
rect 2839 4135 2840 4139
rect 2834 4134 2840 4135
rect 3050 4139 3056 4140
rect 3050 4135 3051 4139
rect 3055 4135 3056 4139
rect 3050 4134 3056 4135
rect 3258 4139 3264 4140
rect 3258 4135 3259 4139
rect 3263 4135 3264 4139
rect 3258 4134 3264 4135
rect 3466 4139 3472 4140
rect 3466 4135 3467 4139
rect 3471 4135 3472 4139
rect 3466 4134 3472 4135
rect 3650 4139 3656 4140
rect 3650 4135 3651 4139
rect 3655 4135 3656 4139
rect 3798 4136 3799 4140
rect 3803 4136 3804 4140
rect 3798 4135 3804 4136
rect 3650 4134 3656 4135
rect 2398 4124 2404 4125
rect 1974 4123 1980 4124
rect 1974 4119 1975 4123
rect 1979 4119 1980 4123
rect 2398 4120 2399 4124
rect 2403 4120 2404 4124
rect 2398 4119 2404 4120
rect 2638 4124 2644 4125
rect 2638 4120 2639 4124
rect 2643 4120 2644 4124
rect 2638 4119 2644 4120
rect 2862 4124 2868 4125
rect 2862 4120 2863 4124
rect 2867 4120 2868 4124
rect 2862 4119 2868 4120
rect 3078 4124 3084 4125
rect 3078 4120 3079 4124
rect 3083 4120 3084 4124
rect 3078 4119 3084 4120
rect 3286 4124 3292 4125
rect 3286 4120 3287 4124
rect 3291 4120 3292 4124
rect 3286 4119 3292 4120
rect 3494 4124 3500 4125
rect 3494 4120 3495 4124
rect 3499 4120 3500 4124
rect 3494 4119 3500 4120
rect 3678 4124 3684 4125
rect 3678 4120 3679 4124
rect 3683 4120 3684 4124
rect 3678 4119 3684 4120
rect 3798 4123 3804 4124
rect 3798 4119 3799 4123
rect 3803 4119 3804 4123
rect 1974 4118 1980 4119
rect 1976 4091 1978 4118
rect 2400 4091 2402 4119
rect 2640 4091 2642 4119
rect 2864 4091 2866 4119
rect 3080 4091 3082 4119
rect 3288 4091 3290 4119
rect 3496 4091 3498 4119
rect 3680 4091 3682 4119
rect 3798 4118 3804 4119
rect 3800 4091 3802 4118
rect 3840 4099 3842 4243
rect 4020 4099 4022 4244
rect 4196 4099 4198 4244
rect 4404 4099 4406 4244
rect 4652 4099 4654 4244
rect 4932 4099 4934 4244
rect 5228 4099 5230 4244
rect 5516 4099 5518 4244
rect 5662 4243 5668 4244
rect 5664 4099 5666 4243
rect 3839 4098 3843 4099
rect 3839 4093 3843 4094
rect 4019 4098 4023 4099
rect 4019 4093 4023 4094
rect 4195 4098 4199 4099
rect 4195 4093 4199 4094
rect 4403 4098 4407 4099
rect 4403 4093 4407 4094
rect 4651 4098 4655 4099
rect 4651 4093 4655 4094
rect 4931 4098 4935 4099
rect 4931 4093 4935 4094
rect 5227 4098 5231 4099
rect 5227 4093 5231 4094
rect 5515 4098 5519 4099
rect 5515 4093 5519 4094
rect 5663 4098 5667 4099
rect 5663 4093 5667 4094
rect 1975 4090 1979 4091
rect 1975 4085 1979 4086
rect 2375 4090 2379 4091
rect 2375 4085 2379 4086
rect 2399 4090 2403 4091
rect 2399 4085 2403 4086
rect 2623 4090 2627 4091
rect 2623 4085 2627 4086
rect 2639 4090 2643 4091
rect 2639 4085 2643 4086
rect 2855 4090 2859 4091
rect 2855 4085 2859 4086
rect 2863 4090 2867 4091
rect 2863 4085 2867 4086
rect 3071 4090 3075 4091
rect 3071 4085 3075 4086
rect 3079 4090 3083 4091
rect 3079 4085 3083 4086
rect 3279 4090 3283 4091
rect 3279 4085 3283 4086
rect 3287 4090 3291 4091
rect 3287 4085 3291 4086
rect 3487 4090 3491 4091
rect 3487 4085 3491 4086
rect 3495 4090 3499 4091
rect 3495 4085 3499 4086
rect 3679 4090 3683 4091
rect 3679 4085 3683 4086
rect 3799 4090 3803 4091
rect 3799 4085 3803 4086
rect 111 4070 115 4071
rect 111 4065 115 4066
rect 627 4070 631 4071
rect 627 4065 631 4066
rect 699 4070 703 4071
rect 699 4065 703 4066
rect 763 4070 767 4071
rect 763 4065 767 4066
rect 835 4070 839 4071
rect 835 4065 839 4066
rect 899 4070 903 4071
rect 899 4065 903 4066
rect 971 4070 975 4071
rect 971 4065 975 4066
rect 1035 4070 1039 4071
rect 1035 4065 1039 4066
rect 1107 4070 1111 4071
rect 1107 4065 1111 4066
rect 1171 4070 1175 4071
rect 1171 4065 1175 4066
rect 1243 4070 1247 4071
rect 1243 4065 1247 4066
rect 1307 4070 1311 4071
rect 1307 4065 1311 4066
rect 1379 4070 1383 4071
rect 1379 4065 1383 4066
rect 1443 4070 1447 4071
rect 1443 4065 1447 4066
rect 1515 4070 1519 4071
rect 1515 4065 1519 4066
rect 1579 4070 1583 4071
rect 1579 4065 1583 4066
rect 1651 4070 1655 4071
rect 1651 4065 1655 4066
rect 1715 4070 1719 4071
rect 1715 4065 1719 4066
rect 1787 4070 1791 4071
rect 1787 4065 1791 4066
rect 1935 4070 1939 4071
rect 1935 4065 1939 4066
rect 112 4005 114 4065
rect 110 4004 116 4005
rect 628 4004 630 4065
rect 764 4004 766 4065
rect 900 4004 902 4065
rect 1036 4004 1038 4065
rect 1172 4004 1174 4065
rect 1308 4004 1310 4065
rect 1444 4004 1446 4065
rect 1580 4004 1582 4065
rect 1716 4004 1718 4065
rect 1936 4005 1938 4065
rect 1976 4062 1978 4085
rect 1974 4061 1980 4062
rect 2376 4061 2378 4085
rect 2624 4061 2626 4085
rect 2856 4061 2858 4085
rect 3072 4061 3074 4085
rect 3280 4061 3282 4085
rect 3488 4061 3490 4085
rect 3680 4061 3682 4085
rect 3800 4062 3802 4085
rect 3798 4061 3804 4062
rect 1974 4057 1975 4061
rect 1979 4057 1980 4061
rect 1974 4056 1980 4057
rect 2374 4060 2380 4061
rect 2374 4056 2375 4060
rect 2379 4056 2380 4060
rect 2374 4055 2380 4056
rect 2622 4060 2628 4061
rect 2622 4056 2623 4060
rect 2627 4056 2628 4060
rect 2622 4055 2628 4056
rect 2854 4060 2860 4061
rect 2854 4056 2855 4060
rect 2859 4056 2860 4060
rect 2854 4055 2860 4056
rect 3070 4060 3076 4061
rect 3070 4056 3071 4060
rect 3075 4056 3076 4060
rect 3070 4055 3076 4056
rect 3278 4060 3284 4061
rect 3278 4056 3279 4060
rect 3283 4056 3284 4060
rect 3278 4055 3284 4056
rect 3486 4060 3492 4061
rect 3486 4056 3487 4060
rect 3491 4056 3492 4060
rect 3486 4055 3492 4056
rect 3678 4060 3684 4061
rect 3678 4056 3679 4060
rect 3683 4056 3684 4060
rect 3798 4057 3799 4061
rect 3803 4057 3804 4061
rect 3798 4056 3804 4057
rect 3678 4055 3684 4056
rect 2346 4045 2352 4046
rect 1974 4044 1980 4045
rect 1974 4040 1975 4044
rect 1979 4040 1980 4044
rect 2346 4041 2347 4045
rect 2351 4041 2352 4045
rect 2346 4040 2352 4041
rect 2594 4045 2600 4046
rect 2594 4041 2595 4045
rect 2599 4041 2600 4045
rect 2594 4040 2600 4041
rect 2826 4045 2832 4046
rect 2826 4041 2827 4045
rect 2831 4041 2832 4045
rect 2826 4040 2832 4041
rect 3042 4045 3048 4046
rect 3042 4041 3043 4045
rect 3047 4041 3048 4045
rect 3042 4040 3048 4041
rect 3250 4045 3256 4046
rect 3250 4041 3251 4045
rect 3255 4041 3256 4045
rect 3250 4040 3256 4041
rect 3458 4045 3464 4046
rect 3458 4041 3459 4045
rect 3463 4041 3464 4045
rect 3458 4040 3464 4041
rect 3650 4045 3656 4046
rect 3650 4041 3651 4045
rect 3655 4041 3656 4045
rect 3650 4040 3656 4041
rect 3798 4044 3804 4045
rect 3798 4040 3799 4044
rect 3803 4040 3804 4044
rect 1974 4039 1980 4040
rect 1934 4004 1940 4005
rect 110 4000 111 4004
rect 115 4000 116 4004
rect 110 3999 116 4000
rect 626 4003 632 4004
rect 626 3999 627 4003
rect 631 3999 632 4003
rect 626 3998 632 3999
rect 762 4003 768 4004
rect 762 3999 763 4003
rect 767 3999 768 4003
rect 762 3998 768 3999
rect 898 4003 904 4004
rect 898 3999 899 4003
rect 903 3999 904 4003
rect 898 3998 904 3999
rect 1034 4003 1040 4004
rect 1034 3999 1035 4003
rect 1039 3999 1040 4003
rect 1034 3998 1040 3999
rect 1170 4003 1176 4004
rect 1170 3999 1171 4003
rect 1175 3999 1176 4003
rect 1170 3998 1176 3999
rect 1306 4003 1312 4004
rect 1306 3999 1307 4003
rect 1311 3999 1312 4003
rect 1306 3998 1312 3999
rect 1442 4003 1448 4004
rect 1442 3999 1443 4003
rect 1447 3999 1448 4003
rect 1442 3998 1448 3999
rect 1578 4003 1584 4004
rect 1578 3999 1579 4003
rect 1583 3999 1584 4003
rect 1578 3998 1584 3999
rect 1714 4003 1720 4004
rect 1714 3999 1715 4003
rect 1719 3999 1720 4003
rect 1934 4000 1935 4004
rect 1939 4000 1940 4004
rect 1934 3999 1940 4000
rect 1714 3998 1720 3999
rect 654 3988 660 3989
rect 110 3987 116 3988
rect 110 3983 111 3987
rect 115 3983 116 3987
rect 654 3984 655 3988
rect 659 3984 660 3988
rect 654 3983 660 3984
rect 790 3988 796 3989
rect 790 3984 791 3988
rect 795 3984 796 3988
rect 790 3983 796 3984
rect 926 3988 932 3989
rect 926 3984 927 3988
rect 931 3984 932 3988
rect 926 3983 932 3984
rect 1062 3988 1068 3989
rect 1062 3984 1063 3988
rect 1067 3984 1068 3988
rect 1062 3983 1068 3984
rect 1198 3988 1204 3989
rect 1198 3984 1199 3988
rect 1203 3984 1204 3988
rect 1198 3983 1204 3984
rect 1334 3988 1340 3989
rect 1334 3984 1335 3988
rect 1339 3984 1340 3988
rect 1334 3983 1340 3984
rect 1470 3988 1476 3989
rect 1470 3984 1471 3988
rect 1475 3984 1476 3988
rect 1470 3983 1476 3984
rect 1606 3988 1612 3989
rect 1606 3984 1607 3988
rect 1611 3984 1612 3988
rect 1606 3983 1612 3984
rect 1742 3988 1748 3989
rect 1742 3984 1743 3988
rect 1747 3984 1748 3988
rect 1742 3983 1748 3984
rect 1934 3987 1940 3988
rect 1934 3983 1935 3987
rect 1939 3983 1940 3987
rect 110 3982 116 3983
rect 112 3947 114 3982
rect 656 3947 658 3983
rect 792 3947 794 3983
rect 928 3947 930 3983
rect 1064 3947 1066 3983
rect 1200 3947 1202 3983
rect 1336 3947 1338 3983
rect 1472 3947 1474 3983
rect 1608 3947 1610 3983
rect 1744 3947 1746 3983
rect 1934 3982 1940 3983
rect 1936 3947 1938 3982
rect 1976 3979 1978 4039
rect 2348 3979 2350 4040
rect 2596 3979 2598 4040
rect 2828 3979 2830 4040
rect 3044 3979 3046 4040
rect 3252 3979 3254 4040
rect 3460 3979 3462 4040
rect 3652 3979 3654 4040
rect 3798 4039 3804 4040
rect 3800 3979 3802 4039
rect 3840 4033 3842 4093
rect 3838 4032 3844 4033
rect 5516 4032 5518 4093
rect 5664 4033 5666 4093
rect 5662 4032 5668 4033
rect 3838 4028 3839 4032
rect 3843 4028 3844 4032
rect 3838 4027 3844 4028
rect 5514 4031 5520 4032
rect 5514 4027 5515 4031
rect 5519 4027 5520 4031
rect 5662 4028 5663 4032
rect 5667 4028 5668 4032
rect 5662 4027 5668 4028
rect 5514 4026 5520 4027
rect 5542 4016 5548 4017
rect 3838 4015 3844 4016
rect 3838 4011 3839 4015
rect 3843 4011 3844 4015
rect 5542 4012 5543 4016
rect 5547 4012 5548 4016
rect 5542 4011 5548 4012
rect 5662 4015 5668 4016
rect 5662 4011 5663 4015
rect 5667 4011 5668 4015
rect 3838 4010 3844 4011
rect 3840 3979 3842 4010
rect 5544 3979 5546 4011
rect 5662 4010 5668 4011
rect 5664 3979 5666 4010
rect 1975 3978 1979 3979
rect 1975 3973 1979 3974
rect 2323 3978 2327 3979
rect 2323 3973 2327 3974
rect 2347 3978 2351 3979
rect 2347 3973 2351 3974
rect 2571 3978 2575 3979
rect 2571 3973 2575 3974
rect 2595 3978 2599 3979
rect 2595 3973 2599 3974
rect 2803 3978 2807 3979
rect 2803 3973 2807 3974
rect 2827 3978 2831 3979
rect 2827 3973 2831 3974
rect 3027 3978 3031 3979
rect 3027 3973 3031 3974
rect 3043 3978 3047 3979
rect 3043 3973 3047 3974
rect 3243 3978 3247 3979
rect 3243 3973 3247 3974
rect 3251 3978 3255 3979
rect 3251 3973 3255 3974
rect 3459 3978 3463 3979
rect 3459 3973 3463 3974
rect 3651 3978 3655 3979
rect 3651 3973 3655 3974
rect 3799 3978 3803 3979
rect 3799 3973 3803 3974
rect 3839 3978 3843 3979
rect 3839 3973 3843 3974
rect 4183 3978 4187 3979
rect 4183 3973 4187 3974
rect 4319 3978 4323 3979
rect 4319 3973 4323 3974
rect 4455 3978 4459 3979
rect 4455 3973 4459 3974
rect 4591 3978 4595 3979
rect 4591 3973 4595 3974
rect 4727 3978 4731 3979
rect 4727 3973 4731 3974
rect 4863 3978 4867 3979
rect 4863 3973 4867 3974
rect 4999 3978 5003 3979
rect 4999 3973 5003 3974
rect 5135 3978 5139 3979
rect 5135 3973 5139 3974
rect 5271 3978 5275 3979
rect 5271 3973 5275 3974
rect 5407 3978 5411 3979
rect 5407 3973 5411 3974
rect 5543 3978 5547 3979
rect 5543 3973 5547 3974
rect 5663 3978 5667 3979
rect 5663 3973 5667 3974
rect 111 3946 115 3947
rect 111 3941 115 3942
rect 599 3946 603 3947
rect 599 3941 603 3942
rect 655 3946 659 3947
rect 655 3941 659 3942
rect 743 3946 747 3947
rect 743 3941 747 3942
rect 791 3946 795 3947
rect 791 3941 795 3942
rect 895 3946 899 3947
rect 895 3941 899 3942
rect 927 3946 931 3947
rect 927 3941 931 3942
rect 1047 3946 1051 3947
rect 1047 3941 1051 3942
rect 1063 3946 1067 3947
rect 1063 3941 1067 3942
rect 1199 3946 1203 3947
rect 1199 3941 1203 3942
rect 1335 3946 1339 3947
rect 1335 3941 1339 3942
rect 1359 3946 1363 3947
rect 1359 3941 1363 3942
rect 1471 3946 1475 3947
rect 1471 3941 1475 3942
rect 1519 3946 1523 3947
rect 1519 3941 1523 3942
rect 1607 3946 1611 3947
rect 1607 3941 1611 3942
rect 1679 3946 1683 3947
rect 1679 3941 1683 3942
rect 1743 3946 1747 3947
rect 1743 3941 1747 3942
rect 1935 3946 1939 3947
rect 1935 3941 1939 3942
rect 112 3918 114 3941
rect 110 3917 116 3918
rect 600 3917 602 3941
rect 744 3917 746 3941
rect 896 3917 898 3941
rect 1048 3917 1050 3941
rect 1200 3917 1202 3941
rect 1360 3917 1362 3941
rect 1520 3917 1522 3941
rect 1680 3917 1682 3941
rect 1936 3918 1938 3941
rect 1934 3917 1940 3918
rect 110 3913 111 3917
rect 115 3913 116 3917
rect 110 3912 116 3913
rect 598 3916 604 3917
rect 598 3912 599 3916
rect 603 3912 604 3916
rect 598 3911 604 3912
rect 742 3916 748 3917
rect 742 3912 743 3916
rect 747 3912 748 3916
rect 742 3911 748 3912
rect 894 3916 900 3917
rect 894 3912 895 3916
rect 899 3912 900 3916
rect 894 3911 900 3912
rect 1046 3916 1052 3917
rect 1046 3912 1047 3916
rect 1051 3912 1052 3916
rect 1046 3911 1052 3912
rect 1198 3916 1204 3917
rect 1198 3912 1199 3916
rect 1203 3912 1204 3916
rect 1198 3911 1204 3912
rect 1358 3916 1364 3917
rect 1358 3912 1359 3916
rect 1363 3912 1364 3916
rect 1358 3911 1364 3912
rect 1518 3916 1524 3917
rect 1518 3912 1519 3916
rect 1523 3912 1524 3916
rect 1518 3911 1524 3912
rect 1678 3916 1684 3917
rect 1678 3912 1679 3916
rect 1683 3912 1684 3916
rect 1934 3913 1935 3917
rect 1939 3913 1940 3917
rect 1976 3913 1978 3973
rect 1934 3912 1940 3913
rect 1974 3912 1980 3913
rect 2324 3912 2326 3973
rect 2572 3912 2574 3973
rect 2804 3912 2806 3973
rect 3028 3912 3030 3973
rect 3244 3912 3246 3973
rect 3460 3912 3462 3973
rect 3652 3912 3654 3973
rect 3800 3913 3802 3973
rect 3840 3950 3842 3973
rect 3838 3949 3844 3950
rect 4184 3949 4186 3973
rect 4320 3949 4322 3973
rect 4456 3949 4458 3973
rect 4592 3949 4594 3973
rect 4728 3949 4730 3973
rect 4864 3949 4866 3973
rect 5000 3949 5002 3973
rect 5136 3949 5138 3973
rect 5272 3949 5274 3973
rect 5408 3949 5410 3973
rect 5544 3949 5546 3973
rect 5664 3950 5666 3973
rect 5662 3949 5668 3950
rect 3838 3945 3839 3949
rect 3843 3945 3844 3949
rect 3838 3944 3844 3945
rect 4182 3948 4188 3949
rect 4182 3944 4183 3948
rect 4187 3944 4188 3948
rect 4182 3943 4188 3944
rect 4318 3948 4324 3949
rect 4318 3944 4319 3948
rect 4323 3944 4324 3948
rect 4318 3943 4324 3944
rect 4454 3948 4460 3949
rect 4454 3944 4455 3948
rect 4459 3944 4460 3948
rect 4454 3943 4460 3944
rect 4590 3948 4596 3949
rect 4590 3944 4591 3948
rect 4595 3944 4596 3948
rect 4590 3943 4596 3944
rect 4726 3948 4732 3949
rect 4726 3944 4727 3948
rect 4731 3944 4732 3948
rect 4726 3943 4732 3944
rect 4862 3948 4868 3949
rect 4862 3944 4863 3948
rect 4867 3944 4868 3948
rect 4862 3943 4868 3944
rect 4998 3948 5004 3949
rect 4998 3944 4999 3948
rect 5003 3944 5004 3948
rect 4998 3943 5004 3944
rect 5134 3948 5140 3949
rect 5134 3944 5135 3948
rect 5139 3944 5140 3948
rect 5134 3943 5140 3944
rect 5270 3948 5276 3949
rect 5270 3944 5271 3948
rect 5275 3944 5276 3948
rect 5270 3943 5276 3944
rect 5406 3948 5412 3949
rect 5406 3944 5407 3948
rect 5411 3944 5412 3948
rect 5406 3943 5412 3944
rect 5542 3948 5548 3949
rect 5542 3944 5543 3948
rect 5547 3944 5548 3948
rect 5662 3945 5663 3949
rect 5667 3945 5668 3949
rect 5662 3944 5668 3945
rect 5542 3943 5548 3944
rect 4154 3933 4160 3934
rect 3838 3932 3844 3933
rect 3838 3928 3839 3932
rect 3843 3928 3844 3932
rect 4154 3929 4155 3933
rect 4159 3929 4160 3933
rect 4154 3928 4160 3929
rect 4290 3933 4296 3934
rect 4290 3929 4291 3933
rect 4295 3929 4296 3933
rect 4290 3928 4296 3929
rect 4426 3933 4432 3934
rect 4426 3929 4427 3933
rect 4431 3929 4432 3933
rect 4426 3928 4432 3929
rect 4562 3933 4568 3934
rect 4562 3929 4563 3933
rect 4567 3929 4568 3933
rect 4562 3928 4568 3929
rect 4698 3933 4704 3934
rect 4698 3929 4699 3933
rect 4703 3929 4704 3933
rect 4698 3928 4704 3929
rect 4834 3933 4840 3934
rect 4834 3929 4835 3933
rect 4839 3929 4840 3933
rect 4834 3928 4840 3929
rect 4970 3933 4976 3934
rect 4970 3929 4971 3933
rect 4975 3929 4976 3933
rect 4970 3928 4976 3929
rect 5106 3933 5112 3934
rect 5106 3929 5107 3933
rect 5111 3929 5112 3933
rect 5106 3928 5112 3929
rect 5242 3933 5248 3934
rect 5242 3929 5243 3933
rect 5247 3929 5248 3933
rect 5242 3928 5248 3929
rect 5378 3933 5384 3934
rect 5378 3929 5379 3933
rect 5383 3929 5384 3933
rect 5378 3928 5384 3929
rect 5514 3933 5520 3934
rect 5514 3929 5515 3933
rect 5519 3929 5520 3933
rect 5514 3928 5520 3929
rect 5662 3932 5668 3933
rect 5662 3928 5663 3932
rect 5667 3928 5668 3932
rect 3838 3927 3844 3928
rect 3798 3912 3804 3913
rect 1678 3911 1684 3912
rect 1974 3908 1975 3912
rect 1979 3908 1980 3912
rect 1974 3907 1980 3908
rect 2322 3911 2328 3912
rect 2322 3907 2323 3911
rect 2327 3907 2328 3911
rect 2322 3906 2328 3907
rect 2570 3911 2576 3912
rect 2570 3907 2571 3911
rect 2575 3907 2576 3911
rect 2570 3906 2576 3907
rect 2802 3911 2808 3912
rect 2802 3907 2803 3911
rect 2807 3907 2808 3911
rect 2802 3906 2808 3907
rect 3026 3911 3032 3912
rect 3026 3907 3027 3911
rect 3031 3907 3032 3911
rect 3026 3906 3032 3907
rect 3242 3911 3248 3912
rect 3242 3907 3243 3911
rect 3247 3907 3248 3911
rect 3242 3906 3248 3907
rect 3458 3911 3464 3912
rect 3458 3907 3459 3911
rect 3463 3907 3464 3911
rect 3458 3906 3464 3907
rect 3650 3911 3656 3912
rect 3650 3907 3651 3911
rect 3655 3907 3656 3911
rect 3798 3908 3799 3912
rect 3803 3908 3804 3912
rect 3798 3907 3804 3908
rect 3650 3906 3656 3907
rect 570 3901 576 3902
rect 110 3900 116 3901
rect 110 3896 111 3900
rect 115 3896 116 3900
rect 570 3897 571 3901
rect 575 3897 576 3901
rect 570 3896 576 3897
rect 714 3901 720 3902
rect 714 3897 715 3901
rect 719 3897 720 3901
rect 714 3896 720 3897
rect 866 3901 872 3902
rect 866 3897 867 3901
rect 871 3897 872 3901
rect 866 3896 872 3897
rect 1018 3901 1024 3902
rect 1018 3897 1019 3901
rect 1023 3897 1024 3901
rect 1018 3896 1024 3897
rect 1170 3901 1176 3902
rect 1170 3897 1171 3901
rect 1175 3897 1176 3901
rect 1170 3896 1176 3897
rect 1330 3901 1336 3902
rect 1330 3897 1331 3901
rect 1335 3897 1336 3901
rect 1330 3896 1336 3897
rect 1490 3901 1496 3902
rect 1490 3897 1491 3901
rect 1495 3897 1496 3901
rect 1490 3896 1496 3897
rect 1650 3901 1656 3902
rect 1650 3897 1651 3901
rect 1655 3897 1656 3901
rect 1650 3896 1656 3897
rect 1934 3900 1940 3901
rect 1934 3896 1935 3900
rect 1939 3896 1940 3900
rect 2350 3896 2356 3897
rect 110 3895 116 3896
rect 112 3827 114 3895
rect 572 3827 574 3896
rect 716 3827 718 3896
rect 868 3827 870 3896
rect 1020 3827 1022 3896
rect 1172 3827 1174 3896
rect 1332 3827 1334 3896
rect 1492 3827 1494 3896
rect 1652 3827 1654 3896
rect 1934 3895 1940 3896
rect 1974 3895 1980 3896
rect 1936 3827 1938 3895
rect 1974 3891 1975 3895
rect 1979 3891 1980 3895
rect 2350 3892 2351 3896
rect 2355 3892 2356 3896
rect 2350 3891 2356 3892
rect 2598 3896 2604 3897
rect 2598 3892 2599 3896
rect 2603 3892 2604 3896
rect 2598 3891 2604 3892
rect 2830 3896 2836 3897
rect 2830 3892 2831 3896
rect 2835 3892 2836 3896
rect 2830 3891 2836 3892
rect 3054 3896 3060 3897
rect 3054 3892 3055 3896
rect 3059 3892 3060 3896
rect 3054 3891 3060 3892
rect 3270 3896 3276 3897
rect 3270 3892 3271 3896
rect 3275 3892 3276 3896
rect 3270 3891 3276 3892
rect 3486 3896 3492 3897
rect 3486 3892 3487 3896
rect 3491 3892 3492 3896
rect 3486 3891 3492 3892
rect 3678 3896 3684 3897
rect 3678 3892 3679 3896
rect 3683 3892 3684 3896
rect 3678 3891 3684 3892
rect 3798 3895 3804 3896
rect 3798 3891 3799 3895
rect 3803 3891 3804 3895
rect 1974 3890 1980 3891
rect 1976 3863 1978 3890
rect 2352 3863 2354 3891
rect 2600 3863 2602 3891
rect 2832 3863 2834 3891
rect 3056 3863 3058 3891
rect 3272 3863 3274 3891
rect 3488 3863 3490 3891
rect 3680 3863 3682 3891
rect 3798 3890 3804 3891
rect 3800 3863 3802 3890
rect 1975 3862 1979 3863
rect 1975 3857 1979 3858
rect 2239 3862 2243 3863
rect 2239 3857 2243 3858
rect 2351 3862 2355 3863
rect 2351 3857 2355 3858
rect 2479 3862 2483 3863
rect 2479 3857 2483 3858
rect 2599 3862 2603 3863
rect 2599 3857 2603 3858
rect 2703 3862 2707 3863
rect 2703 3857 2707 3858
rect 2831 3862 2835 3863
rect 2831 3857 2835 3858
rect 2919 3862 2923 3863
rect 2919 3857 2923 3858
rect 3055 3862 3059 3863
rect 3055 3857 3059 3858
rect 3119 3862 3123 3863
rect 3119 3857 3123 3858
rect 3271 3862 3275 3863
rect 3271 3857 3275 3858
rect 3311 3862 3315 3863
rect 3311 3857 3315 3858
rect 3487 3862 3491 3863
rect 3487 3857 3491 3858
rect 3503 3862 3507 3863
rect 3503 3857 3507 3858
rect 3679 3862 3683 3863
rect 3679 3857 3683 3858
rect 3799 3862 3803 3863
rect 3799 3857 3803 3858
rect 1976 3834 1978 3857
rect 1974 3833 1980 3834
rect 2240 3833 2242 3857
rect 2480 3833 2482 3857
rect 2704 3833 2706 3857
rect 2920 3833 2922 3857
rect 3120 3833 3122 3857
rect 3312 3833 3314 3857
rect 3504 3833 3506 3857
rect 3680 3833 3682 3857
rect 3800 3834 3802 3857
rect 3840 3835 3842 3927
rect 4156 3835 4158 3928
rect 4292 3835 4294 3928
rect 4428 3835 4430 3928
rect 4564 3835 4566 3928
rect 4700 3835 4702 3928
rect 4836 3835 4838 3928
rect 4972 3835 4974 3928
rect 5108 3835 5110 3928
rect 5244 3835 5246 3928
rect 5380 3835 5382 3928
rect 5516 3835 5518 3928
rect 5662 3927 5668 3928
rect 5664 3835 5666 3927
rect 3839 3834 3843 3835
rect 3798 3833 3804 3834
rect 1974 3829 1975 3833
rect 1979 3829 1980 3833
rect 1974 3828 1980 3829
rect 2238 3832 2244 3833
rect 2238 3828 2239 3832
rect 2243 3828 2244 3832
rect 2238 3827 2244 3828
rect 2478 3832 2484 3833
rect 2478 3828 2479 3832
rect 2483 3828 2484 3832
rect 2478 3827 2484 3828
rect 2702 3832 2708 3833
rect 2702 3828 2703 3832
rect 2707 3828 2708 3832
rect 2702 3827 2708 3828
rect 2918 3832 2924 3833
rect 2918 3828 2919 3832
rect 2923 3828 2924 3832
rect 2918 3827 2924 3828
rect 3118 3832 3124 3833
rect 3118 3828 3119 3832
rect 3123 3828 3124 3832
rect 3118 3827 3124 3828
rect 3310 3832 3316 3833
rect 3310 3828 3311 3832
rect 3315 3828 3316 3832
rect 3310 3827 3316 3828
rect 3502 3832 3508 3833
rect 3502 3828 3503 3832
rect 3507 3828 3508 3832
rect 3502 3827 3508 3828
rect 3678 3832 3684 3833
rect 3678 3828 3679 3832
rect 3683 3828 3684 3832
rect 3798 3829 3799 3833
rect 3803 3829 3804 3833
rect 3839 3829 3843 3830
rect 4139 3834 4143 3835
rect 4139 3829 4143 3830
rect 4155 3834 4159 3835
rect 4155 3829 4159 3830
rect 4291 3834 4295 3835
rect 4291 3829 4295 3830
rect 4323 3834 4327 3835
rect 4323 3829 4327 3830
rect 4427 3834 4431 3835
rect 4427 3829 4431 3830
rect 4531 3834 4535 3835
rect 4531 3829 4535 3830
rect 4563 3834 4567 3835
rect 4563 3829 4567 3830
rect 4699 3834 4703 3835
rect 4699 3829 4703 3830
rect 4763 3834 4767 3835
rect 4763 3829 4767 3830
rect 4835 3834 4839 3835
rect 4835 3829 4839 3830
rect 4971 3834 4975 3835
rect 4971 3829 4975 3830
rect 5011 3834 5015 3835
rect 5011 3829 5015 3830
rect 5107 3834 5111 3835
rect 5107 3829 5111 3830
rect 5243 3834 5247 3835
rect 5243 3829 5247 3830
rect 5275 3834 5279 3835
rect 5275 3829 5279 3830
rect 5379 3834 5383 3835
rect 5379 3829 5383 3830
rect 5515 3834 5519 3835
rect 5515 3829 5519 3830
rect 5663 3834 5667 3835
rect 5663 3829 5667 3830
rect 3798 3828 3804 3829
rect 3678 3827 3684 3828
rect 111 3826 115 3827
rect 111 3821 115 3822
rect 427 3826 431 3827
rect 427 3821 431 3822
rect 571 3826 575 3827
rect 571 3821 575 3822
rect 587 3826 591 3827
rect 587 3821 591 3822
rect 715 3826 719 3827
rect 715 3821 719 3822
rect 755 3826 759 3827
rect 755 3821 759 3822
rect 867 3826 871 3827
rect 867 3821 871 3822
rect 923 3826 927 3827
rect 923 3821 927 3822
rect 1019 3826 1023 3827
rect 1019 3821 1023 3822
rect 1099 3826 1103 3827
rect 1099 3821 1103 3822
rect 1171 3826 1175 3827
rect 1171 3821 1175 3822
rect 1275 3826 1279 3827
rect 1275 3821 1279 3822
rect 1331 3826 1335 3827
rect 1331 3821 1335 3822
rect 1459 3826 1463 3827
rect 1459 3821 1463 3822
rect 1491 3826 1495 3827
rect 1491 3821 1495 3822
rect 1643 3826 1647 3827
rect 1643 3821 1647 3822
rect 1651 3826 1655 3827
rect 1651 3821 1655 3822
rect 1935 3826 1939 3827
rect 1935 3821 1939 3822
rect 112 3761 114 3821
rect 110 3760 116 3761
rect 428 3760 430 3821
rect 588 3760 590 3821
rect 756 3760 758 3821
rect 924 3760 926 3821
rect 1100 3760 1102 3821
rect 1276 3760 1278 3821
rect 1460 3760 1462 3821
rect 1644 3760 1646 3821
rect 1936 3761 1938 3821
rect 2210 3817 2216 3818
rect 1974 3816 1980 3817
rect 1974 3812 1975 3816
rect 1979 3812 1980 3816
rect 2210 3813 2211 3817
rect 2215 3813 2216 3817
rect 2210 3812 2216 3813
rect 2450 3817 2456 3818
rect 2450 3813 2451 3817
rect 2455 3813 2456 3817
rect 2450 3812 2456 3813
rect 2674 3817 2680 3818
rect 2674 3813 2675 3817
rect 2679 3813 2680 3817
rect 2674 3812 2680 3813
rect 2890 3817 2896 3818
rect 2890 3813 2891 3817
rect 2895 3813 2896 3817
rect 2890 3812 2896 3813
rect 3090 3817 3096 3818
rect 3090 3813 3091 3817
rect 3095 3813 3096 3817
rect 3090 3812 3096 3813
rect 3282 3817 3288 3818
rect 3282 3813 3283 3817
rect 3287 3813 3288 3817
rect 3282 3812 3288 3813
rect 3474 3817 3480 3818
rect 3474 3813 3475 3817
rect 3479 3813 3480 3817
rect 3474 3812 3480 3813
rect 3650 3817 3656 3818
rect 3650 3813 3651 3817
rect 3655 3813 3656 3817
rect 3650 3812 3656 3813
rect 3798 3816 3804 3817
rect 3798 3812 3799 3816
rect 3803 3812 3804 3816
rect 1974 3811 1980 3812
rect 1934 3760 1940 3761
rect 110 3756 111 3760
rect 115 3756 116 3760
rect 110 3755 116 3756
rect 426 3759 432 3760
rect 426 3755 427 3759
rect 431 3755 432 3759
rect 426 3754 432 3755
rect 586 3759 592 3760
rect 586 3755 587 3759
rect 591 3755 592 3759
rect 586 3754 592 3755
rect 754 3759 760 3760
rect 754 3755 755 3759
rect 759 3755 760 3759
rect 754 3754 760 3755
rect 922 3759 928 3760
rect 922 3755 923 3759
rect 927 3755 928 3759
rect 922 3754 928 3755
rect 1098 3759 1104 3760
rect 1098 3755 1099 3759
rect 1103 3755 1104 3759
rect 1098 3754 1104 3755
rect 1274 3759 1280 3760
rect 1274 3755 1275 3759
rect 1279 3755 1280 3759
rect 1274 3754 1280 3755
rect 1458 3759 1464 3760
rect 1458 3755 1459 3759
rect 1463 3755 1464 3759
rect 1458 3754 1464 3755
rect 1642 3759 1648 3760
rect 1642 3755 1643 3759
rect 1647 3755 1648 3759
rect 1934 3756 1935 3760
rect 1939 3756 1940 3760
rect 1934 3755 1940 3756
rect 1642 3754 1648 3755
rect 454 3744 460 3745
rect 110 3743 116 3744
rect 110 3739 111 3743
rect 115 3739 116 3743
rect 454 3740 455 3744
rect 459 3740 460 3744
rect 454 3739 460 3740
rect 614 3744 620 3745
rect 614 3740 615 3744
rect 619 3740 620 3744
rect 614 3739 620 3740
rect 782 3744 788 3745
rect 782 3740 783 3744
rect 787 3740 788 3744
rect 782 3739 788 3740
rect 950 3744 956 3745
rect 950 3740 951 3744
rect 955 3740 956 3744
rect 950 3739 956 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1302 3744 1308 3745
rect 1302 3740 1303 3744
rect 1307 3740 1308 3744
rect 1302 3739 1308 3740
rect 1486 3744 1492 3745
rect 1486 3740 1487 3744
rect 1491 3740 1492 3744
rect 1486 3739 1492 3740
rect 1670 3744 1676 3745
rect 1670 3740 1671 3744
rect 1675 3740 1676 3744
rect 1670 3739 1676 3740
rect 1934 3743 1940 3744
rect 1976 3743 1978 3811
rect 2212 3743 2214 3812
rect 2452 3743 2454 3812
rect 2676 3743 2678 3812
rect 2892 3743 2894 3812
rect 3092 3743 3094 3812
rect 3284 3743 3286 3812
rect 3476 3743 3478 3812
rect 3652 3743 3654 3812
rect 3798 3811 3804 3812
rect 3800 3743 3802 3811
rect 3840 3769 3842 3829
rect 3838 3768 3844 3769
rect 4140 3768 4142 3829
rect 4324 3768 4326 3829
rect 4532 3768 4534 3829
rect 4764 3768 4766 3829
rect 5012 3768 5014 3829
rect 5276 3768 5278 3829
rect 5516 3768 5518 3829
rect 5664 3769 5666 3829
rect 5662 3768 5668 3769
rect 3838 3764 3839 3768
rect 3843 3764 3844 3768
rect 3838 3763 3844 3764
rect 4138 3767 4144 3768
rect 4138 3763 4139 3767
rect 4143 3763 4144 3767
rect 4138 3762 4144 3763
rect 4322 3767 4328 3768
rect 4322 3763 4323 3767
rect 4327 3763 4328 3767
rect 4322 3762 4328 3763
rect 4530 3767 4536 3768
rect 4530 3763 4531 3767
rect 4535 3763 4536 3767
rect 4530 3762 4536 3763
rect 4762 3767 4768 3768
rect 4762 3763 4763 3767
rect 4767 3763 4768 3767
rect 4762 3762 4768 3763
rect 5010 3767 5016 3768
rect 5010 3763 5011 3767
rect 5015 3763 5016 3767
rect 5010 3762 5016 3763
rect 5274 3767 5280 3768
rect 5274 3763 5275 3767
rect 5279 3763 5280 3767
rect 5274 3762 5280 3763
rect 5514 3767 5520 3768
rect 5514 3763 5515 3767
rect 5519 3763 5520 3767
rect 5662 3764 5663 3768
rect 5667 3764 5668 3768
rect 5662 3763 5668 3764
rect 5514 3762 5520 3763
rect 4166 3752 4172 3753
rect 3838 3751 3844 3752
rect 3838 3747 3839 3751
rect 3843 3747 3844 3751
rect 4166 3748 4167 3752
rect 4171 3748 4172 3752
rect 4166 3747 4172 3748
rect 4350 3752 4356 3753
rect 4350 3748 4351 3752
rect 4355 3748 4356 3752
rect 4350 3747 4356 3748
rect 4558 3752 4564 3753
rect 4558 3748 4559 3752
rect 4563 3748 4564 3752
rect 4558 3747 4564 3748
rect 4790 3752 4796 3753
rect 4790 3748 4791 3752
rect 4795 3748 4796 3752
rect 4790 3747 4796 3748
rect 5038 3752 5044 3753
rect 5038 3748 5039 3752
rect 5043 3748 5044 3752
rect 5038 3747 5044 3748
rect 5302 3752 5308 3753
rect 5302 3748 5303 3752
rect 5307 3748 5308 3752
rect 5302 3747 5308 3748
rect 5542 3752 5548 3753
rect 5542 3748 5543 3752
rect 5547 3748 5548 3752
rect 5542 3747 5548 3748
rect 5662 3751 5668 3752
rect 5662 3747 5663 3751
rect 5667 3747 5668 3751
rect 3838 3746 3844 3747
rect 1934 3739 1935 3743
rect 1939 3739 1940 3743
rect 110 3738 116 3739
rect 112 3703 114 3738
rect 456 3703 458 3739
rect 616 3703 618 3739
rect 784 3703 786 3739
rect 952 3703 954 3739
rect 1128 3703 1130 3739
rect 1304 3703 1306 3739
rect 1488 3703 1490 3739
rect 1672 3703 1674 3739
rect 1934 3738 1940 3739
rect 1975 3742 1979 3743
rect 1936 3703 1938 3738
rect 1975 3737 1979 3738
rect 2211 3742 2215 3743
rect 2211 3737 2215 3738
rect 2227 3742 2231 3743
rect 2227 3737 2231 3738
rect 2451 3742 2455 3743
rect 2451 3737 2455 3738
rect 2667 3742 2671 3743
rect 2667 3737 2671 3738
rect 2675 3742 2679 3743
rect 2675 3737 2679 3738
rect 2875 3742 2879 3743
rect 2875 3737 2879 3738
rect 2891 3742 2895 3743
rect 2891 3737 2895 3738
rect 3075 3742 3079 3743
rect 3075 3737 3079 3738
rect 3091 3742 3095 3743
rect 3091 3737 3095 3738
rect 3275 3742 3279 3743
rect 3275 3737 3279 3738
rect 3283 3742 3287 3743
rect 3283 3737 3287 3738
rect 3475 3742 3479 3743
rect 3475 3737 3479 3738
rect 3651 3742 3655 3743
rect 3651 3737 3655 3738
rect 3799 3742 3803 3743
rect 3799 3737 3803 3738
rect 111 3702 115 3703
rect 111 3697 115 3698
rect 327 3702 331 3703
rect 327 3697 331 3698
rect 455 3702 459 3703
rect 455 3697 459 3698
rect 495 3702 499 3703
rect 495 3697 499 3698
rect 615 3702 619 3703
rect 615 3697 619 3698
rect 679 3702 683 3703
rect 679 3697 683 3698
rect 783 3702 787 3703
rect 783 3697 787 3698
rect 863 3702 867 3703
rect 863 3697 867 3698
rect 951 3702 955 3703
rect 951 3697 955 3698
rect 1055 3702 1059 3703
rect 1055 3697 1059 3698
rect 1127 3702 1131 3703
rect 1127 3697 1131 3698
rect 1255 3702 1259 3703
rect 1255 3697 1259 3698
rect 1303 3702 1307 3703
rect 1303 3697 1307 3698
rect 1455 3702 1459 3703
rect 1455 3697 1459 3698
rect 1487 3702 1491 3703
rect 1487 3697 1491 3698
rect 1655 3702 1659 3703
rect 1655 3697 1659 3698
rect 1671 3702 1675 3703
rect 1671 3697 1675 3698
rect 1935 3702 1939 3703
rect 1935 3697 1939 3698
rect 112 3674 114 3697
rect 110 3673 116 3674
rect 328 3673 330 3697
rect 496 3673 498 3697
rect 680 3673 682 3697
rect 864 3673 866 3697
rect 1056 3673 1058 3697
rect 1256 3673 1258 3697
rect 1456 3673 1458 3697
rect 1656 3673 1658 3697
rect 1936 3674 1938 3697
rect 1976 3677 1978 3737
rect 1974 3676 1980 3677
rect 2228 3676 2230 3737
rect 2452 3676 2454 3737
rect 2668 3676 2670 3737
rect 2876 3676 2878 3737
rect 3076 3676 3078 3737
rect 3276 3676 3278 3737
rect 3476 3676 3478 3737
rect 3800 3677 3802 3737
rect 3840 3703 3842 3746
rect 4168 3703 4170 3747
rect 4352 3703 4354 3747
rect 4560 3703 4562 3747
rect 4792 3703 4794 3747
rect 5040 3703 5042 3747
rect 5304 3703 5306 3747
rect 5544 3703 5546 3747
rect 5662 3746 5668 3747
rect 5664 3703 5666 3746
rect 3839 3702 3843 3703
rect 3839 3697 3843 3698
rect 4167 3702 4171 3703
rect 4167 3697 4171 3698
rect 4303 3702 4307 3703
rect 4303 3697 4307 3698
rect 4351 3702 4355 3703
rect 4351 3697 4355 3698
rect 4479 3702 4483 3703
rect 4479 3697 4483 3698
rect 4559 3702 4563 3703
rect 4559 3697 4563 3698
rect 4671 3702 4675 3703
rect 4671 3697 4675 3698
rect 4791 3702 4795 3703
rect 4791 3697 4795 3698
rect 4879 3702 4883 3703
rect 4879 3697 4883 3698
rect 5039 3702 5043 3703
rect 5039 3697 5043 3698
rect 5103 3702 5107 3703
rect 5103 3697 5107 3698
rect 5303 3702 5307 3703
rect 5303 3697 5307 3698
rect 5335 3702 5339 3703
rect 5335 3697 5339 3698
rect 5543 3702 5547 3703
rect 5543 3697 5547 3698
rect 5663 3702 5667 3703
rect 5663 3697 5667 3698
rect 3798 3676 3804 3677
rect 1934 3673 1940 3674
rect 110 3669 111 3673
rect 115 3669 116 3673
rect 110 3668 116 3669
rect 326 3672 332 3673
rect 326 3668 327 3672
rect 331 3668 332 3672
rect 326 3667 332 3668
rect 494 3672 500 3673
rect 494 3668 495 3672
rect 499 3668 500 3672
rect 494 3667 500 3668
rect 678 3672 684 3673
rect 678 3668 679 3672
rect 683 3668 684 3672
rect 678 3667 684 3668
rect 862 3672 868 3673
rect 862 3668 863 3672
rect 867 3668 868 3672
rect 862 3667 868 3668
rect 1054 3672 1060 3673
rect 1054 3668 1055 3672
rect 1059 3668 1060 3672
rect 1054 3667 1060 3668
rect 1254 3672 1260 3673
rect 1254 3668 1255 3672
rect 1259 3668 1260 3672
rect 1254 3667 1260 3668
rect 1454 3672 1460 3673
rect 1454 3668 1455 3672
rect 1459 3668 1460 3672
rect 1454 3667 1460 3668
rect 1654 3672 1660 3673
rect 1654 3668 1655 3672
rect 1659 3668 1660 3672
rect 1934 3669 1935 3673
rect 1939 3669 1940 3673
rect 1974 3672 1975 3676
rect 1979 3672 1980 3676
rect 1974 3671 1980 3672
rect 2226 3675 2232 3676
rect 2226 3671 2227 3675
rect 2231 3671 2232 3675
rect 2226 3670 2232 3671
rect 2450 3675 2456 3676
rect 2450 3671 2451 3675
rect 2455 3671 2456 3675
rect 2450 3670 2456 3671
rect 2666 3675 2672 3676
rect 2666 3671 2667 3675
rect 2671 3671 2672 3675
rect 2666 3670 2672 3671
rect 2874 3675 2880 3676
rect 2874 3671 2875 3675
rect 2879 3671 2880 3675
rect 2874 3670 2880 3671
rect 3074 3675 3080 3676
rect 3074 3671 3075 3675
rect 3079 3671 3080 3675
rect 3074 3670 3080 3671
rect 3274 3675 3280 3676
rect 3274 3671 3275 3675
rect 3279 3671 3280 3675
rect 3274 3670 3280 3671
rect 3474 3675 3480 3676
rect 3474 3671 3475 3675
rect 3479 3671 3480 3675
rect 3798 3672 3799 3676
rect 3803 3672 3804 3676
rect 3840 3674 3842 3697
rect 3798 3671 3804 3672
rect 3838 3673 3844 3674
rect 4304 3673 4306 3697
rect 4480 3673 4482 3697
rect 4672 3673 4674 3697
rect 4880 3673 4882 3697
rect 5104 3673 5106 3697
rect 5336 3673 5338 3697
rect 5544 3673 5546 3697
rect 5664 3674 5666 3697
rect 5662 3673 5668 3674
rect 3474 3670 3480 3671
rect 1934 3668 1940 3669
rect 3838 3669 3839 3673
rect 3843 3669 3844 3673
rect 3838 3668 3844 3669
rect 4302 3672 4308 3673
rect 4302 3668 4303 3672
rect 4307 3668 4308 3672
rect 1654 3667 1660 3668
rect 4302 3667 4308 3668
rect 4478 3672 4484 3673
rect 4478 3668 4479 3672
rect 4483 3668 4484 3672
rect 4478 3667 4484 3668
rect 4670 3672 4676 3673
rect 4670 3668 4671 3672
rect 4675 3668 4676 3672
rect 4670 3667 4676 3668
rect 4878 3672 4884 3673
rect 4878 3668 4879 3672
rect 4883 3668 4884 3672
rect 4878 3667 4884 3668
rect 5102 3672 5108 3673
rect 5102 3668 5103 3672
rect 5107 3668 5108 3672
rect 5102 3667 5108 3668
rect 5334 3672 5340 3673
rect 5334 3668 5335 3672
rect 5339 3668 5340 3672
rect 5334 3667 5340 3668
rect 5542 3672 5548 3673
rect 5542 3668 5543 3672
rect 5547 3668 5548 3672
rect 5662 3669 5663 3673
rect 5667 3669 5668 3673
rect 5662 3668 5668 3669
rect 5542 3667 5548 3668
rect 2254 3660 2260 3661
rect 1974 3659 1980 3660
rect 298 3657 304 3658
rect 110 3656 116 3657
rect 110 3652 111 3656
rect 115 3652 116 3656
rect 298 3653 299 3657
rect 303 3653 304 3657
rect 298 3652 304 3653
rect 466 3657 472 3658
rect 466 3653 467 3657
rect 471 3653 472 3657
rect 466 3652 472 3653
rect 650 3657 656 3658
rect 650 3653 651 3657
rect 655 3653 656 3657
rect 650 3652 656 3653
rect 834 3657 840 3658
rect 834 3653 835 3657
rect 839 3653 840 3657
rect 834 3652 840 3653
rect 1026 3657 1032 3658
rect 1026 3653 1027 3657
rect 1031 3653 1032 3657
rect 1026 3652 1032 3653
rect 1226 3657 1232 3658
rect 1226 3653 1227 3657
rect 1231 3653 1232 3657
rect 1226 3652 1232 3653
rect 1426 3657 1432 3658
rect 1426 3653 1427 3657
rect 1431 3653 1432 3657
rect 1426 3652 1432 3653
rect 1626 3657 1632 3658
rect 1626 3653 1627 3657
rect 1631 3653 1632 3657
rect 1626 3652 1632 3653
rect 1934 3656 1940 3657
rect 1934 3652 1935 3656
rect 1939 3652 1940 3656
rect 1974 3655 1975 3659
rect 1979 3655 1980 3659
rect 2254 3656 2255 3660
rect 2259 3656 2260 3660
rect 2254 3655 2260 3656
rect 2478 3660 2484 3661
rect 2478 3656 2479 3660
rect 2483 3656 2484 3660
rect 2478 3655 2484 3656
rect 2694 3660 2700 3661
rect 2694 3656 2695 3660
rect 2699 3656 2700 3660
rect 2694 3655 2700 3656
rect 2902 3660 2908 3661
rect 2902 3656 2903 3660
rect 2907 3656 2908 3660
rect 2902 3655 2908 3656
rect 3102 3660 3108 3661
rect 3102 3656 3103 3660
rect 3107 3656 3108 3660
rect 3102 3655 3108 3656
rect 3302 3660 3308 3661
rect 3302 3656 3303 3660
rect 3307 3656 3308 3660
rect 3302 3655 3308 3656
rect 3502 3660 3508 3661
rect 3502 3656 3503 3660
rect 3507 3656 3508 3660
rect 3502 3655 3508 3656
rect 3798 3659 3804 3660
rect 3798 3655 3799 3659
rect 3803 3655 3804 3659
rect 4274 3657 4280 3658
rect 1974 3654 1980 3655
rect 110 3651 116 3652
rect 112 3571 114 3651
rect 300 3571 302 3652
rect 468 3571 470 3652
rect 652 3571 654 3652
rect 836 3571 838 3652
rect 1028 3571 1030 3652
rect 1228 3571 1230 3652
rect 1428 3571 1430 3652
rect 1628 3571 1630 3652
rect 1934 3651 1940 3652
rect 1936 3571 1938 3651
rect 1976 3627 1978 3654
rect 2256 3627 2258 3655
rect 2480 3627 2482 3655
rect 2696 3627 2698 3655
rect 2904 3627 2906 3655
rect 3104 3627 3106 3655
rect 3304 3627 3306 3655
rect 3504 3627 3506 3655
rect 3798 3654 3804 3655
rect 3838 3656 3844 3657
rect 3800 3627 3802 3654
rect 3838 3652 3839 3656
rect 3843 3652 3844 3656
rect 4274 3653 4275 3657
rect 4279 3653 4280 3657
rect 4274 3652 4280 3653
rect 4450 3657 4456 3658
rect 4450 3653 4451 3657
rect 4455 3653 4456 3657
rect 4450 3652 4456 3653
rect 4642 3657 4648 3658
rect 4642 3653 4643 3657
rect 4647 3653 4648 3657
rect 4642 3652 4648 3653
rect 4850 3657 4856 3658
rect 4850 3653 4851 3657
rect 4855 3653 4856 3657
rect 4850 3652 4856 3653
rect 5074 3657 5080 3658
rect 5074 3653 5075 3657
rect 5079 3653 5080 3657
rect 5074 3652 5080 3653
rect 5306 3657 5312 3658
rect 5306 3653 5307 3657
rect 5311 3653 5312 3657
rect 5306 3652 5312 3653
rect 5514 3657 5520 3658
rect 5514 3653 5515 3657
rect 5519 3653 5520 3657
rect 5514 3652 5520 3653
rect 5662 3656 5668 3657
rect 5662 3652 5663 3656
rect 5667 3652 5668 3656
rect 3838 3651 3844 3652
rect 1975 3626 1979 3627
rect 1975 3621 1979 3622
rect 2135 3626 2139 3627
rect 2135 3621 2139 3622
rect 2255 3626 2259 3627
rect 2255 3621 2259 3622
rect 2311 3626 2315 3627
rect 2311 3621 2315 3622
rect 2479 3626 2483 3627
rect 2479 3621 2483 3622
rect 2647 3626 2651 3627
rect 2647 3621 2651 3622
rect 2695 3626 2699 3627
rect 2695 3621 2699 3622
rect 2807 3626 2811 3627
rect 2807 3621 2811 3622
rect 2903 3626 2907 3627
rect 2903 3621 2907 3622
rect 2967 3626 2971 3627
rect 2967 3621 2971 3622
rect 3103 3626 3107 3627
rect 3103 3621 3107 3622
rect 3135 3626 3139 3627
rect 3135 3621 3139 3622
rect 3303 3626 3307 3627
rect 3303 3621 3307 3622
rect 3503 3626 3507 3627
rect 3503 3621 3507 3622
rect 3799 3626 3803 3627
rect 3799 3621 3803 3622
rect 1976 3598 1978 3621
rect 1974 3597 1980 3598
rect 2136 3597 2138 3621
rect 2312 3597 2314 3621
rect 2480 3597 2482 3621
rect 2648 3597 2650 3621
rect 2808 3597 2810 3621
rect 2968 3597 2970 3621
rect 3136 3597 3138 3621
rect 3304 3597 3306 3621
rect 3800 3598 3802 3621
rect 3798 3597 3804 3598
rect 1974 3593 1975 3597
rect 1979 3593 1980 3597
rect 1974 3592 1980 3593
rect 2134 3596 2140 3597
rect 2134 3592 2135 3596
rect 2139 3592 2140 3596
rect 2134 3591 2140 3592
rect 2310 3596 2316 3597
rect 2310 3592 2311 3596
rect 2315 3592 2316 3596
rect 2310 3591 2316 3592
rect 2478 3596 2484 3597
rect 2478 3592 2479 3596
rect 2483 3592 2484 3596
rect 2478 3591 2484 3592
rect 2646 3596 2652 3597
rect 2646 3592 2647 3596
rect 2651 3592 2652 3596
rect 2646 3591 2652 3592
rect 2806 3596 2812 3597
rect 2806 3592 2807 3596
rect 2811 3592 2812 3596
rect 2806 3591 2812 3592
rect 2966 3596 2972 3597
rect 2966 3592 2967 3596
rect 2971 3592 2972 3596
rect 2966 3591 2972 3592
rect 3134 3596 3140 3597
rect 3134 3592 3135 3596
rect 3139 3592 3140 3596
rect 3134 3591 3140 3592
rect 3302 3596 3308 3597
rect 3302 3592 3303 3596
rect 3307 3592 3308 3596
rect 3798 3593 3799 3597
rect 3803 3593 3804 3597
rect 3798 3592 3804 3593
rect 3302 3591 3308 3592
rect 2106 3581 2112 3582
rect 1974 3580 1980 3581
rect 1974 3576 1975 3580
rect 1979 3576 1980 3580
rect 2106 3577 2107 3581
rect 2111 3577 2112 3581
rect 2106 3576 2112 3577
rect 2282 3581 2288 3582
rect 2282 3577 2283 3581
rect 2287 3577 2288 3581
rect 2282 3576 2288 3577
rect 2450 3581 2456 3582
rect 2450 3577 2451 3581
rect 2455 3577 2456 3581
rect 2450 3576 2456 3577
rect 2618 3581 2624 3582
rect 2618 3577 2619 3581
rect 2623 3577 2624 3581
rect 2618 3576 2624 3577
rect 2778 3581 2784 3582
rect 2778 3577 2779 3581
rect 2783 3577 2784 3581
rect 2778 3576 2784 3577
rect 2938 3581 2944 3582
rect 2938 3577 2939 3581
rect 2943 3577 2944 3581
rect 2938 3576 2944 3577
rect 3106 3581 3112 3582
rect 3106 3577 3107 3581
rect 3111 3577 3112 3581
rect 3106 3576 3112 3577
rect 3274 3581 3280 3582
rect 3274 3577 3275 3581
rect 3279 3577 3280 3581
rect 3274 3576 3280 3577
rect 3798 3580 3804 3581
rect 3798 3576 3799 3580
rect 3803 3576 3804 3580
rect 1974 3575 1980 3576
rect 111 3570 115 3571
rect 111 3565 115 3566
rect 203 3570 207 3571
rect 203 3565 207 3566
rect 299 3570 303 3571
rect 299 3565 303 3566
rect 379 3570 383 3571
rect 379 3565 383 3566
rect 467 3570 471 3571
rect 467 3565 471 3566
rect 563 3570 567 3571
rect 563 3565 567 3566
rect 651 3570 655 3571
rect 651 3565 655 3566
rect 755 3570 759 3571
rect 755 3565 759 3566
rect 835 3570 839 3571
rect 835 3565 839 3566
rect 955 3570 959 3571
rect 955 3565 959 3566
rect 1027 3570 1031 3571
rect 1027 3565 1031 3566
rect 1163 3570 1167 3571
rect 1163 3565 1167 3566
rect 1227 3570 1231 3571
rect 1227 3565 1231 3566
rect 1379 3570 1383 3571
rect 1379 3565 1383 3566
rect 1427 3570 1431 3571
rect 1427 3565 1431 3566
rect 1595 3570 1599 3571
rect 1595 3565 1599 3566
rect 1627 3570 1631 3571
rect 1627 3565 1631 3566
rect 1935 3570 1939 3571
rect 1935 3565 1939 3566
rect 112 3505 114 3565
rect 110 3504 116 3505
rect 204 3504 206 3565
rect 380 3504 382 3565
rect 564 3504 566 3565
rect 756 3504 758 3565
rect 956 3504 958 3565
rect 1164 3504 1166 3565
rect 1380 3504 1382 3565
rect 1596 3504 1598 3565
rect 1936 3505 1938 3565
rect 1934 3504 1940 3505
rect 110 3500 111 3504
rect 115 3500 116 3504
rect 110 3499 116 3500
rect 202 3503 208 3504
rect 202 3499 203 3503
rect 207 3499 208 3503
rect 202 3498 208 3499
rect 378 3503 384 3504
rect 378 3499 379 3503
rect 383 3499 384 3503
rect 378 3498 384 3499
rect 562 3503 568 3504
rect 562 3499 563 3503
rect 567 3499 568 3503
rect 562 3498 568 3499
rect 754 3503 760 3504
rect 754 3499 755 3503
rect 759 3499 760 3503
rect 754 3498 760 3499
rect 954 3503 960 3504
rect 954 3499 955 3503
rect 959 3499 960 3503
rect 954 3498 960 3499
rect 1162 3503 1168 3504
rect 1162 3499 1163 3503
rect 1167 3499 1168 3503
rect 1162 3498 1168 3499
rect 1378 3503 1384 3504
rect 1378 3499 1379 3503
rect 1383 3499 1384 3503
rect 1378 3498 1384 3499
rect 1594 3503 1600 3504
rect 1594 3499 1595 3503
rect 1599 3499 1600 3503
rect 1934 3500 1935 3504
rect 1939 3500 1940 3504
rect 1934 3499 1940 3500
rect 1594 3498 1600 3499
rect 1976 3491 1978 3575
rect 2108 3491 2110 3576
rect 2284 3491 2286 3576
rect 2452 3491 2454 3576
rect 2620 3491 2622 3576
rect 2780 3491 2782 3576
rect 2940 3491 2942 3576
rect 3108 3491 3110 3576
rect 3276 3491 3278 3576
rect 3798 3575 3804 3576
rect 3800 3491 3802 3575
rect 3840 3563 3842 3651
rect 4276 3563 4278 3652
rect 4452 3563 4454 3652
rect 4644 3563 4646 3652
rect 4852 3563 4854 3652
rect 5076 3563 5078 3652
rect 5308 3563 5310 3652
rect 5516 3563 5518 3652
rect 5662 3651 5668 3652
rect 5664 3563 5666 3651
rect 3839 3562 3843 3563
rect 3839 3557 3843 3558
rect 4275 3562 4279 3563
rect 4275 3557 4279 3558
rect 4451 3562 4455 3563
rect 4451 3557 4455 3558
rect 4555 3562 4559 3563
rect 4555 3557 4559 3558
rect 4643 3562 4647 3563
rect 4643 3557 4647 3558
rect 4699 3562 4703 3563
rect 4699 3557 4703 3558
rect 4851 3562 4855 3563
rect 4851 3557 4855 3558
rect 5011 3562 5015 3563
rect 5011 3557 5015 3558
rect 5075 3562 5079 3563
rect 5075 3557 5079 3558
rect 5179 3562 5183 3563
rect 5179 3557 5183 3558
rect 5307 3562 5311 3563
rect 5307 3557 5311 3558
rect 5355 3562 5359 3563
rect 5355 3557 5359 3558
rect 5515 3562 5519 3563
rect 5515 3557 5519 3558
rect 5663 3562 5667 3563
rect 5663 3557 5667 3558
rect 3840 3497 3842 3557
rect 3838 3496 3844 3497
rect 4556 3496 4558 3557
rect 4700 3496 4702 3557
rect 4852 3496 4854 3557
rect 5012 3496 5014 3557
rect 5180 3496 5182 3557
rect 5356 3496 5358 3557
rect 5516 3496 5518 3557
rect 5664 3497 5666 3557
rect 5662 3496 5668 3497
rect 3838 3492 3839 3496
rect 3843 3492 3844 3496
rect 3838 3491 3844 3492
rect 4554 3495 4560 3496
rect 4554 3491 4555 3495
rect 4559 3491 4560 3495
rect 1975 3490 1979 3491
rect 230 3488 236 3489
rect 110 3487 116 3488
rect 110 3483 111 3487
rect 115 3483 116 3487
rect 230 3484 231 3488
rect 235 3484 236 3488
rect 230 3483 236 3484
rect 406 3488 412 3489
rect 406 3484 407 3488
rect 411 3484 412 3488
rect 406 3483 412 3484
rect 590 3488 596 3489
rect 590 3484 591 3488
rect 595 3484 596 3488
rect 590 3483 596 3484
rect 782 3488 788 3489
rect 782 3484 783 3488
rect 787 3484 788 3488
rect 782 3483 788 3484
rect 982 3488 988 3489
rect 982 3484 983 3488
rect 987 3484 988 3488
rect 982 3483 988 3484
rect 1190 3488 1196 3489
rect 1190 3484 1191 3488
rect 1195 3484 1196 3488
rect 1190 3483 1196 3484
rect 1406 3488 1412 3489
rect 1406 3484 1407 3488
rect 1411 3484 1412 3488
rect 1406 3483 1412 3484
rect 1622 3488 1628 3489
rect 1622 3484 1623 3488
rect 1627 3484 1628 3488
rect 1622 3483 1628 3484
rect 1934 3487 1940 3488
rect 1934 3483 1935 3487
rect 1939 3483 1940 3487
rect 1975 3485 1979 3486
rect 2035 3490 2039 3491
rect 2035 3485 2039 3486
rect 2107 3490 2111 3491
rect 2107 3485 2111 3486
rect 2187 3490 2191 3491
rect 2187 3485 2191 3486
rect 2283 3490 2287 3491
rect 2283 3485 2287 3486
rect 2339 3490 2343 3491
rect 2339 3485 2343 3486
rect 2451 3490 2455 3491
rect 2451 3485 2455 3486
rect 2491 3490 2495 3491
rect 2491 3485 2495 3486
rect 2619 3490 2623 3491
rect 2619 3485 2623 3486
rect 2643 3490 2647 3491
rect 2643 3485 2647 3486
rect 2779 3490 2783 3491
rect 2779 3485 2783 3486
rect 2795 3490 2799 3491
rect 2795 3485 2799 3486
rect 2939 3490 2943 3491
rect 2939 3485 2943 3486
rect 2947 3490 2951 3491
rect 2947 3485 2951 3486
rect 3099 3490 3103 3491
rect 3099 3485 3103 3486
rect 3107 3490 3111 3491
rect 3107 3485 3111 3486
rect 3275 3490 3279 3491
rect 3275 3485 3279 3486
rect 3799 3490 3803 3491
rect 4554 3490 4560 3491
rect 4698 3495 4704 3496
rect 4698 3491 4699 3495
rect 4703 3491 4704 3495
rect 4698 3490 4704 3491
rect 4850 3495 4856 3496
rect 4850 3491 4851 3495
rect 4855 3491 4856 3495
rect 4850 3490 4856 3491
rect 5010 3495 5016 3496
rect 5010 3491 5011 3495
rect 5015 3491 5016 3495
rect 5010 3490 5016 3491
rect 5178 3495 5184 3496
rect 5178 3491 5179 3495
rect 5183 3491 5184 3495
rect 5178 3490 5184 3491
rect 5354 3495 5360 3496
rect 5354 3491 5355 3495
rect 5359 3491 5360 3495
rect 5354 3490 5360 3491
rect 5514 3495 5520 3496
rect 5514 3491 5515 3495
rect 5519 3491 5520 3495
rect 5662 3492 5663 3496
rect 5667 3492 5668 3496
rect 5662 3491 5668 3492
rect 5514 3490 5520 3491
rect 3799 3485 3803 3486
rect 110 3482 116 3483
rect 112 3439 114 3482
rect 232 3439 234 3483
rect 408 3439 410 3483
rect 592 3439 594 3483
rect 784 3439 786 3483
rect 984 3439 986 3483
rect 1192 3439 1194 3483
rect 1408 3439 1410 3483
rect 1624 3439 1626 3483
rect 1934 3482 1940 3483
rect 1936 3439 1938 3482
rect 111 3438 115 3439
rect 111 3433 115 3434
rect 231 3438 235 3439
rect 231 3433 235 3434
rect 255 3438 259 3439
rect 255 3433 259 3434
rect 407 3438 411 3439
rect 407 3433 411 3434
rect 471 3438 475 3439
rect 471 3433 475 3434
rect 591 3438 595 3439
rect 591 3433 595 3434
rect 695 3438 699 3439
rect 695 3433 699 3434
rect 783 3438 787 3439
rect 783 3433 787 3434
rect 919 3438 923 3439
rect 919 3433 923 3434
rect 983 3438 987 3439
rect 983 3433 987 3434
rect 1143 3438 1147 3439
rect 1143 3433 1147 3434
rect 1191 3438 1195 3439
rect 1191 3433 1195 3434
rect 1367 3438 1371 3439
rect 1367 3433 1371 3434
rect 1407 3438 1411 3439
rect 1407 3433 1411 3434
rect 1591 3438 1595 3439
rect 1591 3433 1595 3434
rect 1623 3438 1627 3439
rect 1623 3433 1627 3434
rect 1935 3438 1939 3439
rect 1935 3433 1939 3434
rect 112 3410 114 3433
rect 110 3409 116 3410
rect 256 3409 258 3433
rect 472 3409 474 3433
rect 696 3409 698 3433
rect 920 3409 922 3433
rect 1144 3409 1146 3433
rect 1368 3409 1370 3433
rect 1592 3409 1594 3433
rect 1936 3410 1938 3433
rect 1976 3425 1978 3485
rect 1974 3424 1980 3425
rect 2036 3424 2038 3485
rect 2188 3424 2190 3485
rect 2340 3424 2342 3485
rect 2492 3424 2494 3485
rect 2644 3424 2646 3485
rect 2796 3424 2798 3485
rect 2948 3424 2950 3485
rect 3100 3424 3102 3485
rect 3800 3425 3802 3485
rect 4582 3480 4588 3481
rect 3838 3479 3844 3480
rect 3838 3475 3839 3479
rect 3843 3475 3844 3479
rect 4582 3476 4583 3480
rect 4587 3476 4588 3480
rect 4582 3475 4588 3476
rect 4726 3480 4732 3481
rect 4726 3476 4727 3480
rect 4731 3476 4732 3480
rect 4726 3475 4732 3476
rect 4878 3480 4884 3481
rect 4878 3476 4879 3480
rect 4883 3476 4884 3480
rect 4878 3475 4884 3476
rect 5038 3480 5044 3481
rect 5038 3476 5039 3480
rect 5043 3476 5044 3480
rect 5038 3475 5044 3476
rect 5206 3480 5212 3481
rect 5206 3476 5207 3480
rect 5211 3476 5212 3480
rect 5206 3475 5212 3476
rect 5382 3480 5388 3481
rect 5382 3476 5383 3480
rect 5387 3476 5388 3480
rect 5382 3475 5388 3476
rect 5542 3480 5548 3481
rect 5542 3476 5543 3480
rect 5547 3476 5548 3480
rect 5542 3475 5548 3476
rect 5662 3479 5668 3480
rect 5662 3475 5663 3479
rect 5667 3475 5668 3479
rect 3838 3474 3844 3475
rect 3840 3439 3842 3474
rect 4584 3439 4586 3475
rect 4728 3439 4730 3475
rect 4880 3439 4882 3475
rect 5040 3439 5042 3475
rect 5208 3439 5210 3475
rect 5384 3439 5386 3475
rect 5544 3439 5546 3475
rect 5662 3474 5668 3475
rect 5664 3439 5666 3474
rect 3839 3438 3843 3439
rect 3839 3433 3843 3434
rect 4583 3438 4587 3439
rect 4583 3433 4587 3434
rect 4727 3438 4731 3439
rect 4727 3433 4731 3434
rect 4879 3438 4883 3439
rect 4879 3433 4883 3434
rect 4903 3438 4907 3439
rect 4903 3433 4907 3434
rect 5039 3438 5043 3439
rect 5039 3433 5043 3434
rect 5175 3438 5179 3439
rect 5175 3433 5179 3434
rect 5207 3438 5211 3439
rect 5207 3433 5211 3434
rect 5311 3438 5315 3439
rect 5311 3433 5315 3434
rect 5383 3438 5387 3439
rect 5383 3433 5387 3434
rect 5447 3438 5451 3439
rect 5447 3433 5451 3434
rect 5543 3438 5547 3439
rect 5543 3433 5547 3434
rect 5663 3438 5667 3439
rect 5663 3433 5667 3434
rect 3798 3424 3804 3425
rect 1974 3420 1975 3424
rect 1979 3420 1980 3424
rect 1974 3419 1980 3420
rect 2034 3423 2040 3424
rect 2034 3419 2035 3423
rect 2039 3419 2040 3423
rect 2034 3418 2040 3419
rect 2186 3423 2192 3424
rect 2186 3419 2187 3423
rect 2191 3419 2192 3423
rect 2186 3418 2192 3419
rect 2338 3423 2344 3424
rect 2338 3419 2339 3423
rect 2343 3419 2344 3423
rect 2338 3418 2344 3419
rect 2490 3423 2496 3424
rect 2490 3419 2491 3423
rect 2495 3419 2496 3423
rect 2490 3418 2496 3419
rect 2642 3423 2648 3424
rect 2642 3419 2643 3423
rect 2647 3419 2648 3423
rect 2642 3418 2648 3419
rect 2794 3423 2800 3424
rect 2794 3419 2795 3423
rect 2799 3419 2800 3423
rect 2794 3418 2800 3419
rect 2946 3423 2952 3424
rect 2946 3419 2947 3423
rect 2951 3419 2952 3423
rect 2946 3418 2952 3419
rect 3098 3423 3104 3424
rect 3098 3419 3099 3423
rect 3103 3419 3104 3423
rect 3798 3420 3799 3424
rect 3803 3420 3804 3424
rect 3798 3419 3804 3420
rect 3098 3418 3104 3419
rect 3840 3410 3842 3433
rect 1934 3409 1940 3410
rect 3838 3409 3844 3410
rect 4904 3409 4906 3433
rect 5040 3409 5042 3433
rect 5176 3409 5178 3433
rect 5312 3409 5314 3433
rect 5448 3409 5450 3433
rect 5664 3410 5666 3433
rect 5662 3409 5668 3410
rect 110 3405 111 3409
rect 115 3405 116 3409
rect 110 3404 116 3405
rect 254 3408 260 3409
rect 254 3404 255 3408
rect 259 3404 260 3408
rect 254 3403 260 3404
rect 470 3408 476 3409
rect 470 3404 471 3408
rect 475 3404 476 3408
rect 470 3403 476 3404
rect 694 3408 700 3409
rect 694 3404 695 3408
rect 699 3404 700 3408
rect 694 3403 700 3404
rect 918 3408 924 3409
rect 918 3404 919 3408
rect 923 3404 924 3408
rect 918 3403 924 3404
rect 1142 3408 1148 3409
rect 1142 3404 1143 3408
rect 1147 3404 1148 3408
rect 1142 3403 1148 3404
rect 1366 3408 1372 3409
rect 1366 3404 1367 3408
rect 1371 3404 1372 3408
rect 1366 3403 1372 3404
rect 1590 3408 1596 3409
rect 1590 3404 1591 3408
rect 1595 3404 1596 3408
rect 1934 3405 1935 3409
rect 1939 3405 1940 3409
rect 2062 3408 2068 3409
rect 1934 3404 1940 3405
rect 1974 3407 1980 3408
rect 1590 3403 1596 3404
rect 1974 3403 1975 3407
rect 1979 3403 1980 3407
rect 2062 3404 2063 3408
rect 2067 3404 2068 3408
rect 2062 3403 2068 3404
rect 2214 3408 2220 3409
rect 2214 3404 2215 3408
rect 2219 3404 2220 3408
rect 2214 3403 2220 3404
rect 2366 3408 2372 3409
rect 2366 3404 2367 3408
rect 2371 3404 2372 3408
rect 2366 3403 2372 3404
rect 2518 3408 2524 3409
rect 2518 3404 2519 3408
rect 2523 3404 2524 3408
rect 2518 3403 2524 3404
rect 2670 3408 2676 3409
rect 2670 3404 2671 3408
rect 2675 3404 2676 3408
rect 2670 3403 2676 3404
rect 2822 3408 2828 3409
rect 2822 3404 2823 3408
rect 2827 3404 2828 3408
rect 2822 3403 2828 3404
rect 2974 3408 2980 3409
rect 2974 3404 2975 3408
rect 2979 3404 2980 3408
rect 2974 3403 2980 3404
rect 3126 3408 3132 3409
rect 3126 3404 3127 3408
rect 3131 3404 3132 3408
rect 3126 3403 3132 3404
rect 3798 3407 3804 3408
rect 3798 3403 3799 3407
rect 3803 3403 3804 3407
rect 3838 3405 3839 3409
rect 3843 3405 3844 3409
rect 3838 3404 3844 3405
rect 4902 3408 4908 3409
rect 4902 3404 4903 3408
rect 4907 3404 4908 3408
rect 4902 3403 4908 3404
rect 5038 3408 5044 3409
rect 5038 3404 5039 3408
rect 5043 3404 5044 3408
rect 5038 3403 5044 3404
rect 5174 3408 5180 3409
rect 5174 3404 5175 3408
rect 5179 3404 5180 3408
rect 5174 3403 5180 3404
rect 5310 3408 5316 3409
rect 5310 3404 5311 3408
rect 5315 3404 5316 3408
rect 5310 3403 5316 3404
rect 5446 3408 5452 3409
rect 5446 3404 5447 3408
rect 5451 3404 5452 3408
rect 5662 3405 5663 3409
rect 5667 3405 5668 3409
rect 5662 3404 5668 3405
rect 5446 3403 5452 3404
rect 1974 3402 1980 3403
rect 226 3393 232 3394
rect 110 3392 116 3393
rect 110 3388 111 3392
rect 115 3388 116 3392
rect 226 3389 227 3393
rect 231 3389 232 3393
rect 226 3388 232 3389
rect 442 3393 448 3394
rect 442 3389 443 3393
rect 447 3389 448 3393
rect 442 3388 448 3389
rect 666 3393 672 3394
rect 666 3389 667 3393
rect 671 3389 672 3393
rect 666 3388 672 3389
rect 890 3393 896 3394
rect 890 3389 891 3393
rect 895 3389 896 3393
rect 890 3388 896 3389
rect 1114 3393 1120 3394
rect 1114 3389 1115 3393
rect 1119 3389 1120 3393
rect 1114 3388 1120 3389
rect 1338 3393 1344 3394
rect 1338 3389 1339 3393
rect 1343 3389 1344 3393
rect 1338 3388 1344 3389
rect 1562 3393 1568 3394
rect 1562 3389 1563 3393
rect 1567 3389 1568 3393
rect 1562 3388 1568 3389
rect 1934 3392 1940 3393
rect 1934 3388 1935 3392
rect 1939 3388 1940 3392
rect 110 3387 116 3388
rect 112 3311 114 3387
rect 228 3311 230 3388
rect 444 3311 446 3388
rect 668 3311 670 3388
rect 892 3311 894 3388
rect 1116 3311 1118 3388
rect 1340 3311 1342 3388
rect 1564 3311 1566 3388
rect 1934 3387 1940 3388
rect 1936 3311 1938 3387
rect 1976 3367 1978 3402
rect 2064 3367 2066 3403
rect 2216 3367 2218 3403
rect 2368 3367 2370 3403
rect 2520 3367 2522 3403
rect 2672 3367 2674 3403
rect 2824 3367 2826 3403
rect 2976 3367 2978 3403
rect 3128 3367 3130 3403
rect 3798 3402 3804 3403
rect 3800 3367 3802 3402
rect 4874 3393 4880 3394
rect 3838 3392 3844 3393
rect 3838 3388 3839 3392
rect 3843 3388 3844 3392
rect 4874 3389 4875 3393
rect 4879 3389 4880 3393
rect 4874 3388 4880 3389
rect 5010 3393 5016 3394
rect 5010 3389 5011 3393
rect 5015 3389 5016 3393
rect 5010 3388 5016 3389
rect 5146 3393 5152 3394
rect 5146 3389 5147 3393
rect 5151 3389 5152 3393
rect 5146 3388 5152 3389
rect 5282 3393 5288 3394
rect 5282 3389 5283 3393
rect 5287 3389 5288 3393
rect 5282 3388 5288 3389
rect 5418 3393 5424 3394
rect 5418 3389 5419 3393
rect 5423 3389 5424 3393
rect 5418 3388 5424 3389
rect 5662 3392 5668 3393
rect 5662 3388 5663 3392
rect 5667 3388 5668 3392
rect 3838 3387 3844 3388
rect 1975 3366 1979 3367
rect 1975 3361 1979 3362
rect 2023 3366 2027 3367
rect 2023 3361 2027 3362
rect 2063 3366 2067 3367
rect 2063 3361 2067 3362
rect 2191 3366 2195 3367
rect 2191 3361 2195 3362
rect 2215 3366 2219 3367
rect 2215 3361 2219 3362
rect 2367 3366 2371 3367
rect 2367 3361 2371 3362
rect 2375 3366 2379 3367
rect 2375 3361 2379 3362
rect 2519 3366 2523 3367
rect 2519 3361 2523 3362
rect 2551 3366 2555 3367
rect 2551 3361 2555 3362
rect 2671 3366 2675 3367
rect 2671 3361 2675 3362
rect 2727 3366 2731 3367
rect 2727 3361 2731 3362
rect 2823 3366 2827 3367
rect 2823 3361 2827 3362
rect 2895 3366 2899 3367
rect 2895 3361 2899 3362
rect 2975 3366 2979 3367
rect 2975 3361 2979 3362
rect 3071 3366 3075 3367
rect 3071 3361 3075 3362
rect 3127 3366 3131 3367
rect 3127 3361 3131 3362
rect 3247 3366 3251 3367
rect 3247 3361 3251 3362
rect 3799 3366 3803 3367
rect 3799 3361 3803 3362
rect 1976 3338 1978 3361
rect 1974 3337 1980 3338
rect 2024 3337 2026 3361
rect 2192 3337 2194 3361
rect 2376 3337 2378 3361
rect 2552 3337 2554 3361
rect 2728 3337 2730 3361
rect 2896 3337 2898 3361
rect 3072 3337 3074 3361
rect 3248 3337 3250 3361
rect 3800 3338 3802 3361
rect 3798 3337 3804 3338
rect 1974 3333 1975 3337
rect 1979 3333 1980 3337
rect 1974 3332 1980 3333
rect 2022 3336 2028 3337
rect 2022 3332 2023 3336
rect 2027 3332 2028 3336
rect 2022 3331 2028 3332
rect 2190 3336 2196 3337
rect 2190 3332 2191 3336
rect 2195 3332 2196 3336
rect 2190 3331 2196 3332
rect 2374 3336 2380 3337
rect 2374 3332 2375 3336
rect 2379 3332 2380 3336
rect 2374 3331 2380 3332
rect 2550 3336 2556 3337
rect 2550 3332 2551 3336
rect 2555 3332 2556 3336
rect 2550 3331 2556 3332
rect 2726 3336 2732 3337
rect 2726 3332 2727 3336
rect 2731 3332 2732 3336
rect 2726 3331 2732 3332
rect 2894 3336 2900 3337
rect 2894 3332 2895 3336
rect 2899 3332 2900 3336
rect 2894 3331 2900 3332
rect 3070 3336 3076 3337
rect 3070 3332 3071 3336
rect 3075 3332 3076 3336
rect 3070 3331 3076 3332
rect 3246 3336 3252 3337
rect 3246 3332 3247 3336
rect 3251 3332 3252 3336
rect 3798 3333 3799 3337
rect 3803 3333 3804 3337
rect 3798 3332 3804 3333
rect 3246 3331 3252 3332
rect 3840 3327 3842 3387
rect 4876 3327 4878 3388
rect 5012 3327 5014 3388
rect 5148 3327 5150 3388
rect 5284 3327 5286 3388
rect 5420 3327 5422 3388
rect 5662 3387 5668 3388
rect 5664 3327 5666 3387
rect 3839 3326 3843 3327
rect 1994 3321 2000 3322
rect 1974 3320 1980 3321
rect 1974 3316 1975 3320
rect 1979 3316 1980 3320
rect 1994 3317 1995 3321
rect 1999 3317 2000 3321
rect 1994 3316 2000 3317
rect 2162 3321 2168 3322
rect 2162 3317 2163 3321
rect 2167 3317 2168 3321
rect 2162 3316 2168 3317
rect 2346 3321 2352 3322
rect 2346 3317 2347 3321
rect 2351 3317 2352 3321
rect 2346 3316 2352 3317
rect 2522 3321 2528 3322
rect 2522 3317 2523 3321
rect 2527 3317 2528 3321
rect 2522 3316 2528 3317
rect 2698 3321 2704 3322
rect 2698 3317 2699 3321
rect 2703 3317 2704 3321
rect 2698 3316 2704 3317
rect 2866 3321 2872 3322
rect 2866 3317 2867 3321
rect 2871 3317 2872 3321
rect 2866 3316 2872 3317
rect 3042 3321 3048 3322
rect 3042 3317 3043 3321
rect 3047 3317 3048 3321
rect 3042 3316 3048 3317
rect 3218 3321 3224 3322
rect 3839 3321 3843 3322
rect 4699 3326 4703 3327
rect 4699 3321 4703 3322
rect 4835 3326 4839 3327
rect 4835 3321 4839 3322
rect 4875 3326 4879 3327
rect 4875 3321 4879 3322
rect 4971 3326 4975 3327
rect 4971 3321 4975 3322
rect 5011 3326 5015 3327
rect 5011 3321 5015 3322
rect 5107 3326 5111 3327
rect 5107 3321 5111 3322
rect 5147 3326 5151 3327
rect 5147 3321 5151 3322
rect 5243 3326 5247 3327
rect 5243 3321 5247 3322
rect 5283 3326 5287 3327
rect 5283 3321 5287 3322
rect 5379 3326 5383 3327
rect 5379 3321 5383 3322
rect 5419 3326 5423 3327
rect 5419 3321 5423 3322
rect 5515 3326 5519 3327
rect 5515 3321 5519 3322
rect 5663 3326 5667 3327
rect 5663 3321 5667 3322
rect 3218 3317 3219 3321
rect 3223 3317 3224 3321
rect 3218 3316 3224 3317
rect 3798 3320 3804 3321
rect 3798 3316 3799 3320
rect 3803 3316 3804 3320
rect 1974 3315 1980 3316
rect 111 3310 115 3311
rect 111 3305 115 3306
rect 211 3310 215 3311
rect 211 3305 215 3306
rect 227 3310 231 3311
rect 227 3305 231 3306
rect 419 3310 423 3311
rect 419 3305 423 3306
rect 443 3310 447 3311
rect 443 3305 447 3306
rect 635 3310 639 3311
rect 635 3305 639 3306
rect 667 3310 671 3311
rect 667 3305 671 3306
rect 851 3310 855 3311
rect 851 3305 855 3306
rect 891 3310 895 3311
rect 891 3305 895 3306
rect 1075 3310 1079 3311
rect 1075 3305 1079 3306
rect 1115 3310 1119 3311
rect 1115 3305 1119 3306
rect 1299 3310 1303 3311
rect 1299 3305 1303 3306
rect 1339 3310 1343 3311
rect 1339 3305 1343 3306
rect 1523 3310 1527 3311
rect 1523 3305 1527 3306
rect 1563 3310 1567 3311
rect 1563 3305 1567 3306
rect 1935 3310 1939 3311
rect 1935 3305 1939 3306
rect 112 3245 114 3305
rect 110 3244 116 3245
rect 212 3244 214 3305
rect 420 3244 422 3305
rect 636 3244 638 3305
rect 852 3244 854 3305
rect 1076 3244 1078 3305
rect 1300 3244 1302 3305
rect 1524 3244 1526 3305
rect 1936 3245 1938 3305
rect 1976 3251 1978 3315
rect 1996 3251 1998 3316
rect 2164 3251 2166 3316
rect 2348 3251 2350 3316
rect 2524 3251 2526 3316
rect 2700 3251 2702 3316
rect 2868 3251 2870 3316
rect 3044 3251 3046 3316
rect 3220 3251 3222 3316
rect 3798 3315 3804 3316
rect 3800 3251 3802 3315
rect 3840 3261 3842 3321
rect 3838 3260 3844 3261
rect 4700 3260 4702 3321
rect 4836 3260 4838 3321
rect 4972 3260 4974 3321
rect 5108 3260 5110 3321
rect 5244 3260 5246 3321
rect 5380 3260 5382 3321
rect 5516 3260 5518 3321
rect 5664 3261 5666 3321
rect 5662 3260 5668 3261
rect 3838 3256 3839 3260
rect 3843 3256 3844 3260
rect 3838 3255 3844 3256
rect 4698 3259 4704 3260
rect 4698 3255 4699 3259
rect 4703 3255 4704 3259
rect 4698 3254 4704 3255
rect 4834 3259 4840 3260
rect 4834 3255 4835 3259
rect 4839 3255 4840 3259
rect 4834 3254 4840 3255
rect 4970 3259 4976 3260
rect 4970 3255 4971 3259
rect 4975 3255 4976 3259
rect 4970 3254 4976 3255
rect 5106 3259 5112 3260
rect 5106 3255 5107 3259
rect 5111 3255 5112 3259
rect 5106 3254 5112 3255
rect 5242 3259 5248 3260
rect 5242 3255 5243 3259
rect 5247 3255 5248 3259
rect 5242 3254 5248 3255
rect 5378 3259 5384 3260
rect 5378 3255 5379 3259
rect 5383 3255 5384 3259
rect 5378 3254 5384 3255
rect 5514 3259 5520 3260
rect 5514 3255 5515 3259
rect 5519 3255 5520 3259
rect 5662 3256 5663 3260
rect 5667 3256 5668 3260
rect 5662 3255 5668 3256
rect 5514 3254 5520 3255
rect 1975 3250 1979 3251
rect 1975 3245 1979 3246
rect 1995 3250 1999 3251
rect 1995 3245 1999 3246
rect 2163 3250 2167 3251
rect 2163 3245 2167 3246
rect 2211 3250 2215 3251
rect 2211 3245 2215 3246
rect 2347 3250 2351 3251
rect 2347 3245 2351 3246
rect 2435 3250 2439 3251
rect 2435 3245 2439 3246
rect 2523 3250 2527 3251
rect 2523 3245 2527 3246
rect 2651 3250 2655 3251
rect 2651 3245 2655 3246
rect 2699 3250 2703 3251
rect 2699 3245 2703 3246
rect 2851 3250 2855 3251
rect 2851 3245 2855 3246
rect 2867 3250 2871 3251
rect 2867 3245 2871 3246
rect 3043 3250 3047 3251
rect 3043 3245 3047 3246
rect 3051 3250 3055 3251
rect 3051 3245 3055 3246
rect 3219 3250 3223 3251
rect 3219 3245 3223 3246
rect 3251 3250 3255 3251
rect 3251 3245 3255 3246
rect 3451 3250 3455 3251
rect 3451 3245 3455 3246
rect 3799 3250 3803 3251
rect 3799 3245 3803 3246
rect 1934 3244 1940 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 110 3239 116 3240
rect 210 3243 216 3244
rect 210 3239 211 3243
rect 215 3239 216 3243
rect 210 3238 216 3239
rect 418 3243 424 3244
rect 418 3239 419 3243
rect 423 3239 424 3243
rect 418 3238 424 3239
rect 634 3243 640 3244
rect 634 3239 635 3243
rect 639 3239 640 3243
rect 634 3238 640 3239
rect 850 3243 856 3244
rect 850 3239 851 3243
rect 855 3239 856 3243
rect 850 3238 856 3239
rect 1074 3243 1080 3244
rect 1074 3239 1075 3243
rect 1079 3239 1080 3243
rect 1074 3238 1080 3239
rect 1298 3243 1304 3244
rect 1298 3239 1299 3243
rect 1303 3239 1304 3243
rect 1298 3238 1304 3239
rect 1522 3243 1528 3244
rect 1522 3239 1523 3243
rect 1527 3239 1528 3243
rect 1934 3240 1935 3244
rect 1939 3240 1940 3244
rect 1934 3239 1940 3240
rect 1522 3238 1528 3239
rect 238 3228 244 3229
rect 110 3227 116 3228
rect 110 3223 111 3227
rect 115 3223 116 3227
rect 238 3224 239 3228
rect 243 3224 244 3228
rect 238 3223 244 3224
rect 446 3228 452 3229
rect 446 3224 447 3228
rect 451 3224 452 3228
rect 446 3223 452 3224
rect 662 3228 668 3229
rect 662 3224 663 3228
rect 667 3224 668 3228
rect 662 3223 668 3224
rect 878 3228 884 3229
rect 878 3224 879 3228
rect 883 3224 884 3228
rect 878 3223 884 3224
rect 1102 3228 1108 3229
rect 1102 3224 1103 3228
rect 1107 3224 1108 3228
rect 1102 3223 1108 3224
rect 1326 3228 1332 3229
rect 1326 3224 1327 3228
rect 1331 3224 1332 3228
rect 1326 3223 1332 3224
rect 1550 3228 1556 3229
rect 1550 3224 1551 3228
rect 1555 3224 1556 3228
rect 1550 3223 1556 3224
rect 1934 3227 1940 3228
rect 1934 3223 1935 3227
rect 1939 3223 1940 3227
rect 110 3222 116 3223
rect 112 3183 114 3222
rect 240 3183 242 3223
rect 448 3183 450 3223
rect 664 3183 666 3223
rect 880 3183 882 3223
rect 1104 3183 1106 3223
rect 1328 3183 1330 3223
rect 1552 3183 1554 3223
rect 1934 3222 1940 3223
rect 1936 3183 1938 3222
rect 1976 3185 1978 3245
rect 1974 3184 1980 3185
rect 1996 3184 1998 3245
rect 2212 3184 2214 3245
rect 2436 3184 2438 3245
rect 2652 3184 2654 3245
rect 2852 3184 2854 3245
rect 3052 3184 3054 3245
rect 3252 3184 3254 3245
rect 3452 3184 3454 3245
rect 3800 3185 3802 3245
rect 4726 3244 4732 3245
rect 3838 3243 3844 3244
rect 3838 3239 3839 3243
rect 3843 3239 3844 3243
rect 4726 3240 4727 3244
rect 4731 3240 4732 3244
rect 4726 3239 4732 3240
rect 4862 3244 4868 3245
rect 4862 3240 4863 3244
rect 4867 3240 4868 3244
rect 4862 3239 4868 3240
rect 4998 3244 5004 3245
rect 4998 3240 4999 3244
rect 5003 3240 5004 3244
rect 4998 3239 5004 3240
rect 5134 3244 5140 3245
rect 5134 3240 5135 3244
rect 5139 3240 5140 3244
rect 5134 3239 5140 3240
rect 5270 3244 5276 3245
rect 5270 3240 5271 3244
rect 5275 3240 5276 3244
rect 5270 3239 5276 3240
rect 5406 3244 5412 3245
rect 5406 3240 5407 3244
rect 5411 3240 5412 3244
rect 5406 3239 5412 3240
rect 5542 3244 5548 3245
rect 5542 3240 5543 3244
rect 5547 3240 5548 3244
rect 5542 3239 5548 3240
rect 5662 3243 5668 3244
rect 5662 3239 5663 3243
rect 5667 3239 5668 3243
rect 3838 3238 3844 3239
rect 3840 3207 3842 3238
rect 4728 3207 4730 3239
rect 4864 3207 4866 3239
rect 5000 3207 5002 3239
rect 5136 3207 5138 3239
rect 5272 3207 5274 3239
rect 5408 3207 5410 3239
rect 5544 3207 5546 3239
rect 5662 3238 5668 3239
rect 5664 3207 5666 3238
rect 3839 3206 3843 3207
rect 3839 3201 3843 3202
rect 4567 3206 4571 3207
rect 4567 3201 4571 3202
rect 4727 3206 4731 3207
rect 4727 3201 4731 3202
rect 4743 3206 4747 3207
rect 4743 3201 4747 3202
rect 4863 3206 4867 3207
rect 4863 3201 4867 3202
rect 4935 3206 4939 3207
rect 4935 3201 4939 3202
rect 4999 3206 5003 3207
rect 4999 3201 5003 3202
rect 5135 3206 5139 3207
rect 5135 3201 5139 3202
rect 5271 3206 5275 3207
rect 5271 3201 5275 3202
rect 5351 3206 5355 3207
rect 5351 3201 5355 3202
rect 5407 3206 5411 3207
rect 5407 3201 5411 3202
rect 5543 3206 5547 3207
rect 5543 3201 5547 3202
rect 5663 3206 5667 3207
rect 5663 3201 5667 3202
rect 3798 3184 3804 3185
rect 111 3182 115 3183
rect 111 3177 115 3178
rect 239 3182 243 3183
rect 239 3177 243 3178
rect 303 3182 307 3183
rect 303 3177 307 3178
rect 447 3182 451 3183
rect 447 3177 451 3178
rect 543 3182 547 3183
rect 543 3177 547 3178
rect 663 3182 667 3183
rect 663 3177 667 3178
rect 783 3182 787 3183
rect 783 3177 787 3178
rect 879 3182 883 3183
rect 879 3177 883 3178
rect 1023 3182 1027 3183
rect 1023 3177 1027 3178
rect 1103 3182 1107 3183
rect 1103 3177 1107 3178
rect 1263 3182 1267 3183
rect 1263 3177 1267 3178
rect 1327 3182 1331 3183
rect 1327 3177 1331 3178
rect 1511 3182 1515 3183
rect 1511 3177 1515 3178
rect 1551 3182 1555 3183
rect 1551 3177 1555 3178
rect 1935 3182 1939 3183
rect 1974 3180 1975 3184
rect 1979 3180 1980 3184
rect 1974 3179 1980 3180
rect 1994 3183 2000 3184
rect 1994 3179 1995 3183
rect 1999 3179 2000 3183
rect 1994 3178 2000 3179
rect 2210 3183 2216 3184
rect 2210 3179 2211 3183
rect 2215 3179 2216 3183
rect 2210 3178 2216 3179
rect 2434 3183 2440 3184
rect 2434 3179 2435 3183
rect 2439 3179 2440 3183
rect 2434 3178 2440 3179
rect 2650 3183 2656 3184
rect 2650 3179 2651 3183
rect 2655 3179 2656 3183
rect 2650 3178 2656 3179
rect 2850 3183 2856 3184
rect 2850 3179 2851 3183
rect 2855 3179 2856 3183
rect 2850 3178 2856 3179
rect 3050 3183 3056 3184
rect 3050 3179 3051 3183
rect 3055 3179 3056 3183
rect 3050 3178 3056 3179
rect 3250 3183 3256 3184
rect 3250 3179 3251 3183
rect 3255 3179 3256 3183
rect 3250 3178 3256 3179
rect 3450 3183 3456 3184
rect 3450 3179 3451 3183
rect 3455 3179 3456 3183
rect 3798 3180 3799 3184
rect 3803 3180 3804 3184
rect 3798 3179 3804 3180
rect 3450 3178 3456 3179
rect 3840 3178 3842 3201
rect 1935 3177 1939 3178
rect 3838 3177 3844 3178
rect 4568 3177 4570 3201
rect 4744 3177 4746 3201
rect 4936 3177 4938 3201
rect 5136 3177 5138 3201
rect 5352 3177 5354 3201
rect 5544 3177 5546 3201
rect 5664 3178 5666 3201
rect 5662 3177 5668 3178
rect 112 3154 114 3177
rect 110 3153 116 3154
rect 304 3153 306 3177
rect 544 3153 546 3177
rect 784 3153 786 3177
rect 1024 3153 1026 3177
rect 1264 3153 1266 3177
rect 1512 3153 1514 3177
rect 1936 3154 1938 3177
rect 3838 3173 3839 3177
rect 3843 3173 3844 3177
rect 3838 3172 3844 3173
rect 4566 3176 4572 3177
rect 4566 3172 4567 3176
rect 4571 3172 4572 3176
rect 4566 3171 4572 3172
rect 4742 3176 4748 3177
rect 4742 3172 4743 3176
rect 4747 3172 4748 3176
rect 4742 3171 4748 3172
rect 4934 3176 4940 3177
rect 4934 3172 4935 3176
rect 4939 3172 4940 3176
rect 4934 3171 4940 3172
rect 5134 3176 5140 3177
rect 5134 3172 5135 3176
rect 5139 3172 5140 3176
rect 5134 3171 5140 3172
rect 5350 3176 5356 3177
rect 5350 3172 5351 3176
rect 5355 3172 5356 3176
rect 5350 3171 5356 3172
rect 5542 3176 5548 3177
rect 5542 3172 5543 3176
rect 5547 3172 5548 3176
rect 5662 3173 5663 3177
rect 5667 3173 5668 3177
rect 5662 3172 5668 3173
rect 5542 3171 5548 3172
rect 2022 3168 2028 3169
rect 1974 3167 1980 3168
rect 1974 3163 1975 3167
rect 1979 3163 1980 3167
rect 2022 3164 2023 3168
rect 2027 3164 2028 3168
rect 2022 3163 2028 3164
rect 2238 3168 2244 3169
rect 2238 3164 2239 3168
rect 2243 3164 2244 3168
rect 2238 3163 2244 3164
rect 2462 3168 2468 3169
rect 2462 3164 2463 3168
rect 2467 3164 2468 3168
rect 2462 3163 2468 3164
rect 2678 3168 2684 3169
rect 2678 3164 2679 3168
rect 2683 3164 2684 3168
rect 2678 3163 2684 3164
rect 2878 3168 2884 3169
rect 2878 3164 2879 3168
rect 2883 3164 2884 3168
rect 2878 3163 2884 3164
rect 3078 3168 3084 3169
rect 3078 3164 3079 3168
rect 3083 3164 3084 3168
rect 3078 3163 3084 3164
rect 3278 3168 3284 3169
rect 3278 3164 3279 3168
rect 3283 3164 3284 3168
rect 3278 3163 3284 3164
rect 3478 3168 3484 3169
rect 3478 3164 3479 3168
rect 3483 3164 3484 3168
rect 3478 3163 3484 3164
rect 3798 3167 3804 3168
rect 3798 3163 3799 3167
rect 3803 3163 3804 3167
rect 1974 3162 1980 3163
rect 1934 3153 1940 3154
rect 110 3149 111 3153
rect 115 3149 116 3153
rect 110 3148 116 3149
rect 302 3152 308 3153
rect 302 3148 303 3152
rect 307 3148 308 3152
rect 302 3147 308 3148
rect 542 3152 548 3153
rect 542 3148 543 3152
rect 547 3148 548 3152
rect 542 3147 548 3148
rect 782 3152 788 3153
rect 782 3148 783 3152
rect 787 3148 788 3152
rect 782 3147 788 3148
rect 1022 3152 1028 3153
rect 1022 3148 1023 3152
rect 1027 3148 1028 3152
rect 1022 3147 1028 3148
rect 1262 3152 1268 3153
rect 1262 3148 1263 3152
rect 1267 3148 1268 3152
rect 1262 3147 1268 3148
rect 1510 3152 1516 3153
rect 1510 3148 1511 3152
rect 1515 3148 1516 3152
rect 1934 3149 1935 3153
rect 1939 3149 1940 3153
rect 1934 3148 1940 3149
rect 1510 3147 1516 3148
rect 1976 3139 1978 3162
rect 2024 3139 2026 3163
rect 2240 3139 2242 3163
rect 2464 3139 2466 3163
rect 2680 3139 2682 3163
rect 2880 3139 2882 3163
rect 3080 3139 3082 3163
rect 3280 3139 3282 3163
rect 3480 3139 3482 3163
rect 3798 3162 3804 3163
rect 3800 3139 3802 3162
rect 4538 3161 4544 3162
rect 3838 3160 3844 3161
rect 3838 3156 3839 3160
rect 3843 3156 3844 3160
rect 4538 3157 4539 3161
rect 4543 3157 4544 3161
rect 4538 3156 4544 3157
rect 4714 3161 4720 3162
rect 4714 3157 4715 3161
rect 4719 3157 4720 3161
rect 4714 3156 4720 3157
rect 4906 3161 4912 3162
rect 4906 3157 4907 3161
rect 4911 3157 4912 3161
rect 4906 3156 4912 3157
rect 5106 3161 5112 3162
rect 5106 3157 5107 3161
rect 5111 3157 5112 3161
rect 5106 3156 5112 3157
rect 5322 3161 5328 3162
rect 5322 3157 5323 3161
rect 5327 3157 5328 3161
rect 5322 3156 5328 3157
rect 5514 3161 5520 3162
rect 5514 3157 5515 3161
rect 5519 3157 5520 3161
rect 5514 3156 5520 3157
rect 5662 3160 5668 3161
rect 5662 3156 5663 3160
rect 5667 3156 5668 3160
rect 3838 3155 3844 3156
rect 1975 3138 1979 3139
rect 274 3137 280 3138
rect 110 3136 116 3137
rect 110 3132 111 3136
rect 115 3132 116 3136
rect 274 3133 275 3137
rect 279 3133 280 3137
rect 274 3132 280 3133
rect 514 3137 520 3138
rect 514 3133 515 3137
rect 519 3133 520 3137
rect 514 3132 520 3133
rect 754 3137 760 3138
rect 754 3133 755 3137
rect 759 3133 760 3137
rect 754 3132 760 3133
rect 994 3137 1000 3138
rect 994 3133 995 3137
rect 999 3133 1000 3137
rect 994 3132 1000 3133
rect 1234 3137 1240 3138
rect 1234 3133 1235 3137
rect 1239 3133 1240 3137
rect 1234 3132 1240 3133
rect 1482 3137 1488 3138
rect 1482 3133 1483 3137
rect 1487 3133 1488 3137
rect 1482 3132 1488 3133
rect 1934 3136 1940 3137
rect 1934 3132 1935 3136
rect 1939 3132 1940 3136
rect 1975 3133 1979 3134
rect 2023 3138 2027 3139
rect 2023 3133 2027 3134
rect 2239 3138 2243 3139
rect 2239 3133 2243 3134
rect 2327 3138 2331 3139
rect 2327 3133 2331 3134
rect 2463 3138 2467 3139
rect 2463 3133 2467 3134
rect 2631 3138 2635 3139
rect 2631 3133 2635 3134
rect 2679 3138 2683 3139
rect 2679 3133 2683 3134
rect 2879 3138 2883 3139
rect 2879 3133 2883 3134
rect 2911 3138 2915 3139
rect 2911 3133 2915 3134
rect 3079 3138 3083 3139
rect 3079 3133 3083 3134
rect 3175 3138 3179 3139
rect 3175 3133 3179 3134
rect 3279 3138 3283 3139
rect 3279 3133 3283 3134
rect 3439 3138 3443 3139
rect 3439 3133 3443 3134
rect 3479 3138 3483 3139
rect 3479 3133 3483 3134
rect 3679 3138 3683 3139
rect 3679 3133 3683 3134
rect 3799 3138 3803 3139
rect 3799 3133 3803 3134
rect 110 3131 116 3132
rect 112 3071 114 3131
rect 276 3071 278 3132
rect 516 3071 518 3132
rect 756 3071 758 3132
rect 996 3071 998 3132
rect 1236 3071 1238 3132
rect 1484 3071 1486 3132
rect 1934 3131 1940 3132
rect 1936 3071 1938 3131
rect 1976 3110 1978 3133
rect 1974 3109 1980 3110
rect 2024 3109 2026 3133
rect 2328 3109 2330 3133
rect 2632 3109 2634 3133
rect 2912 3109 2914 3133
rect 3176 3109 3178 3133
rect 3440 3109 3442 3133
rect 3680 3109 3682 3133
rect 3800 3110 3802 3133
rect 3798 3109 3804 3110
rect 1974 3105 1975 3109
rect 1979 3105 1980 3109
rect 1974 3104 1980 3105
rect 2022 3108 2028 3109
rect 2022 3104 2023 3108
rect 2027 3104 2028 3108
rect 2022 3103 2028 3104
rect 2326 3108 2332 3109
rect 2326 3104 2327 3108
rect 2331 3104 2332 3108
rect 2326 3103 2332 3104
rect 2630 3108 2636 3109
rect 2630 3104 2631 3108
rect 2635 3104 2636 3108
rect 2630 3103 2636 3104
rect 2910 3108 2916 3109
rect 2910 3104 2911 3108
rect 2915 3104 2916 3108
rect 2910 3103 2916 3104
rect 3174 3108 3180 3109
rect 3174 3104 3175 3108
rect 3179 3104 3180 3108
rect 3174 3103 3180 3104
rect 3438 3108 3444 3109
rect 3438 3104 3439 3108
rect 3443 3104 3444 3108
rect 3438 3103 3444 3104
rect 3678 3108 3684 3109
rect 3678 3104 3679 3108
rect 3683 3104 3684 3108
rect 3798 3105 3799 3109
rect 3803 3105 3804 3109
rect 3798 3104 3804 3105
rect 3678 3103 3684 3104
rect 1994 3093 2000 3094
rect 1974 3092 1980 3093
rect 1974 3088 1975 3092
rect 1979 3088 1980 3092
rect 1994 3089 1995 3093
rect 1999 3089 2000 3093
rect 1994 3088 2000 3089
rect 2298 3093 2304 3094
rect 2298 3089 2299 3093
rect 2303 3089 2304 3093
rect 2298 3088 2304 3089
rect 2602 3093 2608 3094
rect 2602 3089 2603 3093
rect 2607 3089 2608 3093
rect 2602 3088 2608 3089
rect 2882 3093 2888 3094
rect 2882 3089 2883 3093
rect 2887 3089 2888 3093
rect 2882 3088 2888 3089
rect 3146 3093 3152 3094
rect 3146 3089 3147 3093
rect 3151 3089 3152 3093
rect 3146 3088 3152 3089
rect 3410 3093 3416 3094
rect 3410 3089 3411 3093
rect 3415 3089 3416 3093
rect 3410 3088 3416 3089
rect 3650 3093 3656 3094
rect 3650 3089 3651 3093
rect 3655 3089 3656 3093
rect 3650 3088 3656 3089
rect 3798 3092 3804 3093
rect 3798 3088 3799 3092
rect 3803 3088 3804 3092
rect 3840 3091 3842 3155
rect 4540 3091 4542 3156
rect 4716 3091 4718 3156
rect 4908 3091 4910 3156
rect 5108 3091 5110 3156
rect 5324 3091 5326 3156
rect 5516 3091 5518 3156
rect 5662 3155 5668 3156
rect 5664 3091 5666 3155
rect 1974 3087 1980 3088
rect 111 3070 115 3071
rect 111 3065 115 3066
rect 275 3070 279 3071
rect 275 3065 279 3066
rect 355 3070 359 3071
rect 355 3065 359 3066
rect 515 3070 519 3071
rect 515 3065 519 3066
rect 627 3070 631 3071
rect 627 3065 631 3066
rect 755 3070 759 3071
rect 755 3065 759 3066
rect 883 3070 887 3071
rect 883 3065 887 3066
rect 995 3070 999 3071
rect 995 3065 999 3066
rect 1123 3070 1127 3071
rect 1123 3065 1127 3066
rect 1235 3070 1239 3071
rect 1235 3065 1239 3066
rect 1355 3070 1359 3071
rect 1355 3065 1359 3066
rect 1483 3070 1487 3071
rect 1483 3065 1487 3066
rect 1579 3070 1583 3071
rect 1579 3065 1583 3066
rect 1787 3070 1791 3071
rect 1787 3065 1791 3066
rect 1935 3070 1939 3071
rect 1935 3065 1939 3066
rect 112 3005 114 3065
rect 110 3004 116 3005
rect 356 3004 358 3065
rect 628 3004 630 3065
rect 884 3004 886 3065
rect 1124 3004 1126 3065
rect 1356 3004 1358 3065
rect 1580 3004 1582 3065
rect 1788 3004 1790 3065
rect 1936 3005 1938 3065
rect 1976 3019 1978 3087
rect 1996 3019 1998 3088
rect 2300 3019 2302 3088
rect 2604 3019 2606 3088
rect 2884 3019 2886 3088
rect 3148 3019 3150 3088
rect 3412 3019 3414 3088
rect 3652 3019 3654 3088
rect 3798 3087 3804 3088
rect 3839 3090 3843 3091
rect 3800 3019 3802 3087
rect 3839 3085 3843 3086
rect 4307 3090 4311 3091
rect 4307 3085 4311 3086
rect 4483 3090 4487 3091
rect 4483 3085 4487 3086
rect 4539 3090 4543 3091
rect 4539 3085 4543 3086
rect 4675 3090 4679 3091
rect 4675 3085 4679 3086
rect 4715 3090 4719 3091
rect 4715 3085 4719 3086
rect 4875 3090 4879 3091
rect 4875 3085 4879 3086
rect 4907 3090 4911 3091
rect 4907 3085 4911 3086
rect 5091 3090 5095 3091
rect 5091 3085 5095 3086
rect 5107 3090 5111 3091
rect 5107 3085 5111 3086
rect 5315 3090 5319 3091
rect 5315 3085 5319 3086
rect 5323 3090 5327 3091
rect 5323 3085 5327 3086
rect 5515 3090 5519 3091
rect 5515 3085 5519 3086
rect 5663 3090 5667 3091
rect 5663 3085 5667 3086
rect 3840 3025 3842 3085
rect 3838 3024 3844 3025
rect 4308 3024 4310 3085
rect 4484 3024 4486 3085
rect 4676 3024 4678 3085
rect 4876 3024 4878 3085
rect 5092 3024 5094 3085
rect 5316 3024 5318 3085
rect 5516 3024 5518 3085
rect 5664 3025 5666 3085
rect 5662 3024 5668 3025
rect 3838 3020 3839 3024
rect 3843 3020 3844 3024
rect 3838 3019 3844 3020
rect 4306 3023 4312 3024
rect 4306 3019 4307 3023
rect 4311 3019 4312 3023
rect 1975 3018 1979 3019
rect 1975 3013 1979 3014
rect 1995 3018 1999 3019
rect 1995 3013 1999 3014
rect 2299 3018 2303 3019
rect 2299 3013 2303 3014
rect 2603 3018 2607 3019
rect 2603 3013 2607 3014
rect 2883 3018 2887 3019
rect 2883 3013 2887 3014
rect 3107 3018 3111 3019
rect 3107 3013 3111 3014
rect 3147 3018 3151 3019
rect 3147 3013 3151 3014
rect 3243 3018 3247 3019
rect 3243 3013 3247 3014
rect 3379 3018 3383 3019
rect 3379 3013 3383 3014
rect 3411 3018 3415 3019
rect 3411 3013 3415 3014
rect 3515 3018 3519 3019
rect 3515 3013 3519 3014
rect 3651 3018 3655 3019
rect 3651 3013 3655 3014
rect 3799 3018 3803 3019
rect 4306 3018 4312 3019
rect 4482 3023 4488 3024
rect 4482 3019 4483 3023
rect 4487 3019 4488 3023
rect 4482 3018 4488 3019
rect 4674 3023 4680 3024
rect 4674 3019 4675 3023
rect 4679 3019 4680 3023
rect 4674 3018 4680 3019
rect 4874 3023 4880 3024
rect 4874 3019 4875 3023
rect 4879 3019 4880 3023
rect 4874 3018 4880 3019
rect 5090 3023 5096 3024
rect 5090 3019 5091 3023
rect 5095 3019 5096 3023
rect 5090 3018 5096 3019
rect 5314 3023 5320 3024
rect 5314 3019 5315 3023
rect 5319 3019 5320 3023
rect 5314 3018 5320 3019
rect 5514 3023 5520 3024
rect 5514 3019 5515 3023
rect 5519 3019 5520 3023
rect 5662 3020 5663 3024
rect 5667 3020 5668 3024
rect 5662 3019 5668 3020
rect 5514 3018 5520 3019
rect 3799 3013 3803 3014
rect 1934 3004 1940 3005
rect 110 3000 111 3004
rect 115 3000 116 3004
rect 110 2999 116 3000
rect 354 3003 360 3004
rect 354 2999 355 3003
rect 359 2999 360 3003
rect 354 2998 360 2999
rect 626 3003 632 3004
rect 626 2999 627 3003
rect 631 2999 632 3003
rect 626 2998 632 2999
rect 882 3003 888 3004
rect 882 2999 883 3003
rect 887 2999 888 3003
rect 882 2998 888 2999
rect 1122 3003 1128 3004
rect 1122 2999 1123 3003
rect 1127 2999 1128 3003
rect 1122 2998 1128 2999
rect 1354 3003 1360 3004
rect 1354 2999 1355 3003
rect 1359 2999 1360 3003
rect 1354 2998 1360 2999
rect 1578 3003 1584 3004
rect 1578 2999 1579 3003
rect 1583 2999 1584 3003
rect 1578 2998 1584 2999
rect 1786 3003 1792 3004
rect 1786 2999 1787 3003
rect 1791 2999 1792 3003
rect 1934 3000 1935 3004
rect 1939 3000 1940 3004
rect 1934 2999 1940 3000
rect 1786 2998 1792 2999
rect 382 2988 388 2989
rect 110 2987 116 2988
rect 110 2983 111 2987
rect 115 2983 116 2987
rect 382 2984 383 2988
rect 387 2984 388 2988
rect 382 2983 388 2984
rect 654 2988 660 2989
rect 654 2984 655 2988
rect 659 2984 660 2988
rect 654 2983 660 2984
rect 910 2988 916 2989
rect 910 2984 911 2988
rect 915 2984 916 2988
rect 910 2983 916 2984
rect 1150 2988 1156 2989
rect 1150 2984 1151 2988
rect 1155 2984 1156 2988
rect 1150 2983 1156 2984
rect 1382 2988 1388 2989
rect 1382 2984 1383 2988
rect 1387 2984 1388 2988
rect 1382 2983 1388 2984
rect 1606 2988 1612 2989
rect 1606 2984 1607 2988
rect 1611 2984 1612 2988
rect 1606 2983 1612 2984
rect 1814 2988 1820 2989
rect 1814 2984 1815 2988
rect 1819 2984 1820 2988
rect 1814 2983 1820 2984
rect 1934 2987 1940 2988
rect 1934 2983 1935 2987
rect 1939 2983 1940 2987
rect 110 2982 116 2983
rect 112 2959 114 2982
rect 384 2959 386 2983
rect 656 2959 658 2983
rect 912 2959 914 2983
rect 1152 2959 1154 2983
rect 1384 2959 1386 2983
rect 1608 2959 1610 2983
rect 1816 2959 1818 2983
rect 1934 2982 1940 2983
rect 1936 2959 1938 2982
rect 111 2958 115 2959
rect 111 2953 115 2954
rect 343 2958 347 2959
rect 343 2953 347 2954
rect 383 2958 387 2959
rect 383 2953 387 2954
rect 551 2958 555 2959
rect 551 2953 555 2954
rect 655 2958 659 2959
rect 655 2953 659 2954
rect 759 2958 763 2959
rect 759 2953 763 2954
rect 911 2958 915 2959
rect 911 2953 915 2954
rect 951 2958 955 2959
rect 951 2953 955 2954
rect 1135 2958 1139 2959
rect 1135 2953 1139 2954
rect 1151 2958 1155 2959
rect 1151 2953 1155 2954
rect 1311 2958 1315 2959
rect 1311 2953 1315 2954
rect 1383 2958 1387 2959
rect 1383 2953 1387 2954
rect 1487 2958 1491 2959
rect 1487 2953 1491 2954
rect 1607 2958 1611 2959
rect 1607 2953 1611 2954
rect 1663 2958 1667 2959
rect 1663 2953 1667 2954
rect 1815 2958 1819 2959
rect 1815 2953 1819 2954
rect 1935 2958 1939 2959
rect 1935 2953 1939 2954
rect 1976 2953 1978 3013
rect 112 2930 114 2953
rect 110 2929 116 2930
rect 344 2929 346 2953
rect 552 2929 554 2953
rect 760 2929 762 2953
rect 952 2929 954 2953
rect 1136 2929 1138 2953
rect 1312 2929 1314 2953
rect 1488 2929 1490 2953
rect 1664 2929 1666 2953
rect 1816 2929 1818 2953
rect 1936 2930 1938 2953
rect 1974 2952 1980 2953
rect 3108 2952 3110 3013
rect 3244 2952 3246 3013
rect 3380 2952 3382 3013
rect 3516 2952 3518 3013
rect 3652 2952 3654 3013
rect 3800 2953 3802 3013
rect 4334 3008 4340 3009
rect 3838 3007 3844 3008
rect 3838 3003 3839 3007
rect 3843 3003 3844 3007
rect 4334 3004 4335 3008
rect 4339 3004 4340 3008
rect 4334 3003 4340 3004
rect 4510 3008 4516 3009
rect 4510 3004 4511 3008
rect 4515 3004 4516 3008
rect 4510 3003 4516 3004
rect 4702 3008 4708 3009
rect 4702 3004 4703 3008
rect 4707 3004 4708 3008
rect 4702 3003 4708 3004
rect 4902 3008 4908 3009
rect 4902 3004 4903 3008
rect 4907 3004 4908 3008
rect 4902 3003 4908 3004
rect 5118 3008 5124 3009
rect 5118 3004 5119 3008
rect 5123 3004 5124 3008
rect 5118 3003 5124 3004
rect 5342 3008 5348 3009
rect 5342 3004 5343 3008
rect 5347 3004 5348 3008
rect 5342 3003 5348 3004
rect 5542 3008 5548 3009
rect 5542 3004 5543 3008
rect 5547 3004 5548 3008
rect 5542 3003 5548 3004
rect 5662 3007 5668 3008
rect 5662 3003 5663 3007
rect 5667 3003 5668 3007
rect 3838 3002 3844 3003
rect 3840 2975 3842 3002
rect 4336 2975 4338 3003
rect 4512 2975 4514 3003
rect 4704 2975 4706 3003
rect 4904 2975 4906 3003
rect 5120 2975 5122 3003
rect 5344 2975 5346 3003
rect 5544 2975 5546 3003
rect 5662 3002 5668 3003
rect 5664 2975 5666 3002
rect 3839 2974 3843 2975
rect 3839 2969 3843 2970
rect 3887 2974 3891 2975
rect 3887 2969 3891 2970
rect 4023 2974 4027 2975
rect 4023 2969 4027 2970
rect 4175 2974 4179 2975
rect 4175 2969 4179 2970
rect 4335 2974 4339 2975
rect 4335 2969 4339 2970
rect 4391 2974 4395 2975
rect 4391 2969 4395 2970
rect 4511 2974 4515 2975
rect 4511 2969 4515 2970
rect 4639 2974 4643 2975
rect 4639 2969 4643 2970
rect 4703 2974 4707 2975
rect 4703 2969 4707 2970
rect 4903 2974 4907 2975
rect 4903 2969 4907 2970
rect 4919 2974 4923 2975
rect 4919 2969 4923 2970
rect 5119 2974 5123 2975
rect 5119 2969 5123 2970
rect 5223 2974 5227 2975
rect 5223 2969 5227 2970
rect 5343 2974 5347 2975
rect 5343 2969 5347 2970
rect 5527 2974 5531 2975
rect 5527 2969 5531 2970
rect 5543 2974 5547 2975
rect 5543 2969 5547 2970
rect 5663 2974 5667 2975
rect 5663 2969 5667 2970
rect 3798 2952 3804 2953
rect 1974 2948 1975 2952
rect 1979 2948 1980 2952
rect 1974 2947 1980 2948
rect 3106 2951 3112 2952
rect 3106 2947 3107 2951
rect 3111 2947 3112 2951
rect 3106 2946 3112 2947
rect 3242 2951 3248 2952
rect 3242 2947 3243 2951
rect 3247 2947 3248 2951
rect 3242 2946 3248 2947
rect 3378 2951 3384 2952
rect 3378 2947 3379 2951
rect 3383 2947 3384 2951
rect 3378 2946 3384 2947
rect 3514 2951 3520 2952
rect 3514 2947 3515 2951
rect 3519 2947 3520 2951
rect 3514 2946 3520 2947
rect 3650 2951 3656 2952
rect 3650 2947 3651 2951
rect 3655 2947 3656 2951
rect 3798 2948 3799 2952
rect 3803 2948 3804 2952
rect 3798 2947 3804 2948
rect 3650 2946 3656 2947
rect 3840 2946 3842 2969
rect 3838 2945 3844 2946
rect 3888 2945 3890 2969
rect 4024 2945 4026 2969
rect 4176 2945 4178 2969
rect 4392 2945 4394 2969
rect 4640 2945 4642 2969
rect 4920 2945 4922 2969
rect 5224 2945 5226 2969
rect 5528 2945 5530 2969
rect 5664 2946 5666 2969
rect 5662 2945 5668 2946
rect 3838 2941 3839 2945
rect 3843 2941 3844 2945
rect 3838 2940 3844 2941
rect 3886 2944 3892 2945
rect 3886 2940 3887 2944
rect 3891 2940 3892 2944
rect 3886 2939 3892 2940
rect 4022 2944 4028 2945
rect 4022 2940 4023 2944
rect 4027 2940 4028 2944
rect 4022 2939 4028 2940
rect 4174 2944 4180 2945
rect 4174 2940 4175 2944
rect 4179 2940 4180 2944
rect 4174 2939 4180 2940
rect 4390 2944 4396 2945
rect 4390 2940 4391 2944
rect 4395 2940 4396 2944
rect 4390 2939 4396 2940
rect 4638 2944 4644 2945
rect 4638 2940 4639 2944
rect 4643 2940 4644 2944
rect 4638 2939 4644 2940
rect 4918 2944 4924 2945
rect 4918 2940 4919 2944
rect 4923 2940 4924 2944
rect 4918 2939 4924 2940
rect 5222 2944 5228 2945
rect 5222 2940 5223 2944
rect 5227 2940 5228 2944
rect 5222 2939 5228 2940
rect 5526 2944 5532 2945
rect 5526 2940 5527 2944
rect 5531 2940 5532 2944
rect 5662 2941 5663 2945
rect 5667 2941 5668 2945
rect 5662 2940 5668 2941
rect 5526 2939 5532 2940
rect 3134 2936 3140 2937
rect 1974 2935 1980 2936
rect 1974 2931 1975 2935
rect 1979 2931 1980 2935
rect 3134 2932 3135 2936
rect 3139 2932 3140 2936
rect 3134 2931 3140 2932
rect 3270 2936 3276 2937
rect 3270 2932 3271 2936
rect 3275 2932 3276 2936
rect 3270 2931 3276 2932
rect 3406 2936 3412 2937
rect 3406 2932 3407 2936
rect 3411 2932 3412 2936
rect 3406 2931 3412 2932
rect 3542 2936 3548 2937
rect 3542 2932 3543 2936
rect 3547 2932 3548 2936
rect 3542 2931 3548 2932
rect 3678 2936 3684 2937
rect 3678 2932 3679 2936
rect 3683 2932 3684 2936
rect 3678 2931 3684 2932
rect 3798 2935 3804 2936
rect 3798 2931 3799 2935
rect 3803 2931 3804 2935
rect 1974 2930 1980 2931
rect 1934 2929 1940 2930
rect 110 2925 111 2929
rect 115 2925 116 2929
rect 110 2924 116 2925
rect 342 2928 348 2929
rect 342 2924 343 2928
rect 347 2924 348 2928
rect 342 2923 348 2924
rect 550 2928 556 2929
rect 550 2924 551 2928
rect 555 2924 556 2928
rect 550 2923 556 2924
rect 758 2928 764 2929
rect 758 2924 759 2928
rect 763 2924 764 2928
rect 758 2923 764 2924
rect 950 2928 956 2929
rect 950 2924 951 2928
rect 955 2924 956 2928
rect 950 2923 956 2924
rect 1134 2928 1140 2929
rect 1134 2924 1135 2928
rect 1139 2924 1140 2928
rect 1134 2923 1140 2924
rect 1310 2928 1316 2929
rect 1310 2924 1311 2928
rect 1315 2924 1316 2928
rect 1310 2923 1316 2924
rect 1486 2928 1492 2929
rect 1486 2924 1487 2928
rect 1491 2924 1492 2928
rect 1486 2923 1492 2924
rect 1662 2928 1668 2929
rect 1662 2924 1663 2928
rect 1667 2924 1668 2928
rect 1662 2923 1668 2924
rect 1814 2928 1820 2929
rect 1814 2924 1815 2928
rect 1819 2924 1820 2928
rect 1934 2925 1935 2929
rect 1939 2925 1940 2929
rect 1934 2924 1940 2925
rect 1814 2923 1820 2924
rect 314 2913 320 2914
rect 110 2912 116 2913
rect 110 2908 111 2912
rect 115 2908 116 2912
rect 314 2909 315 2913
rect 319 2909 320 2913
rect 314 2908 320 2909
rect 522 2913 528 2914
rect 522 2909 523 2913
rect 527 2909 528 2913
rect 522 2908 528 2909
rect 730 2913 736 2914
rect 730 2909 731 2913
rect 735 2909 736 2913
rect 730 2908 736 2909
rect 922 2913 928 2914
rect 922 2909 923 2913
rect 927 2909 928 2913
rect 922 2908 928 2909
rect 1106 2913 1112 2914
rect 1106 2909 1107 2913
rect 1111 2909 1112 2913
rect 1106 2908 1112 2909
rect 1282 2913 1288 2914
rect 1282 2909 1283 2913
rect 1287 2909 1288 2913
rect 1282 2908 1288 2909
rect 1458 2913 1464 2914
rect 1458 2909 1459 2913
rect 1463 2909 1464 2913
rect 1458 2908 1464 2909
rect 1634 2913 1640 2914
rect 1634 2909 1635 2913
rect 1639 2909 1640 2913
rect 1634 2908 1640 2909
rect 1786 2913 1792 2914
rect 1786 2909 1787 2913
rect 1791 2909 1792 2913
rect 1786 2908 1792 2909
rect 1934 2912 1940 2913
rect 1934 2908 1935 2912
rect 1939 2908 1940 2912
rect 110 2907 116 2908
rect 112 2835 114 2907
rect 316 2835 318 2908
rect 524 2835 526 2908
rect 732 2835 734 2908
rect 924 2835 926 2908
rect 1108 2835 1110 2908
rect 1284 2835 1286 2908
rect 1460 2835 1462 2908
rect 1636 2835 1638 2908
rect 1788 2835 1790 2908
rect 1934 2907 1940 2908
rect 1936 2835 1938 2907
rect 111 2834 115 2835
rect 111 2829 115 2830
rect 315 2834 319 2835
rect 315 2829 319 2830
rect 363 2834 367 2835
rect 363 2829 367 2830
rect 523 2834 527 2835
rect 523 2829 527 2830
rect 563 2834 567 2835
rect 563 2829 567 2830
rect 731 2834 735 2835
rect 731 2829 735 2830
rect 755 2834 759 2835
rect 755 2829 759 2830
rect 923 2834 927 2835
rect 923 2829 927 2830
rect 939 2834 943 2835
rect 939 2829 943 2830
rect 1107 2834 1111 2835
rect 1107 2829 1111 2830
rect 1115 2834 1119 2835
rect 1115 2829 1119 2830
rect 1283 2834 1287 2835
rect 1283 2829 1287 2830
rect 1451 2834 1455 2835
rect 1451 2829 1455 2830
rect 1459 2834 1463 2835
rect 1459 2829 1463 2830
rect 1619 2834 1623 2835
rect 1619 2829 1623 2830
rect 1635 2834 1639 2835
rect 1635 2829 1639 2830
rect 1787 2834 1791 2835
rect 1787 2829 1791 2830
rect 1935 2834 1939 2835
rect 1935 2829 1939 2830
rect 112 2769 114 2829
rect 110 2768 116 2769
rect 364 2768 366 2829
rect 564 2768 566 2829
rect 756 2768 758 2829
rect 940 2768 942 2829
rect 1116 2768 1118 2829
rect 1284 2768 1286 2829
rect 1452 2768 1454 2829
rect 1620 2768 1622 2829
rect 1788 2768 1790 2829
rect 1936 2769 1938 2829
rect 1934 2768 1940 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 362 2767 368 2768
rect 362 2763 363 2767
rect 367 2763 368 2767
rect 362 2762 368 2763
rect 562 2767 568 2768
rect 562 2763 563 2767
rect 567 2763 568 2767
rect 562 2762 568 2763
rect 754 2767 760 2768
rect 754 2763 755 2767
rect 759 2763 760 2767
rect 754 2762 760 2763
rect 938 2767 944 2768
rect 938 2763 939 2767
rect 943 2763 944 2767
rect 938 2762 944 2763
rect 1114 2767 1120 2768
rect 1114 2763 1115 2767
rect 1119 2763 1120 2767
rect 1114 2762 1120 2763
rect 1282 2767 1288 2768
rect 1282 2763 1283 2767
rect 1287 2763 1288 2767
rect 1282 2762 1288 2763
rect 1450 2767 1456 2768
rect 1450 2763 1451 2767
rect 1455 2763 1456 2767
rect 1450 2762 1456 2763
rect 1618 2767 1624 2768
rect 1618 2763 1619 2767
rect 1623 2763 1624 2767
rect 1618 2762 1624 2763
rect 1786 2767 1792 2768
rect 1786 2763 1787 2767
rect 1791 2763 1792 2767
rect 1934 2764 1935 2768
rect 1939 2764 1940 2768
rect 1934 2763 1940 2764
rect 1786 2762 1792 2763
rect 390 2752 396 2753
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 390 2748 391 2752
rect 395 2748 396 2752
rect 390 2747 396 2748
rect 590 2752 596 2753
rect 590 2748 591 2752
rect 595 2748 596 2752
rect 590 2747 596 2748
rect 782 2752 788 2753
rect 782 2748 783 2752
rect 787 2748 788 2752
rect 782 2747 788 2748
rect 966 2752 972 2753
rect 966 2748 967 2752
rect 971 2748 972 2752
rect 966 2747 972 2748
rect 1142 2752 1148 2753
rect 1142 2748 1143 2752
rect 1147 2748 1148 2752
rect 1142 2747 1148 2748
rect 1310 2752 1316 2753
rect 1310 2748 1311 2752
rect 1315 2748 1316 2752
rect 1310 2747 1316 2748
rect 1478 2752 1484 2753
rect 1478 2748 1479 2752
rect 1483 2748 1484 2752
rect 1478 2747 1484 2748
rect 1646 2752 1652 2753
rect 1646 2748 1647 2752
rect 1651 2748 1652 2752
rect 1646 2747 1652 2748
rect 1814 2752 1820 2753
rect 1814 2748 1815 2752
rect 1819 2748 1820 2752
rect 1814 2747 1820 2748
rect 1934 2751 1940 2752
rect 1934 2747 1935 2751
rect 1939 2747 1940 2751
rect 110 2746 116 2747
rect 112 2719 114 2746
rect 392 2719 394 2747
rect 592 2719 594 2747
rect 784 2719 786 2747
rect 968 2719 970 2747
rect 1144 2719 1146 2747
rect 1312 2719 1314 2747
rect 1480 2719 1482 2747
rect 1648 2719 1650 2747
rect 1816 2719 1818 2747
rect 1934 2746 1940 2747
rect 1936 2719 1938 2746
rect 111 2718 115 2719
rect 111 2713 115 2714
rect 391 2718 395 2719
rect 391 2713 395 2714
rect 447 2718 451 2719
rect 447 2713 451 2714
rect 591 2718 595 2719
rect 591 2713 595 2714
rect 615 2718 619 2719
rect 615 2713 619 2714
rect 775 2718 779 2719
rect 775 2713 779 2714
rect 783 2718 787 2719
rect 783 2713 787 2714
rect 935 2718 939 2719
rect 935 2713 939 2714
rect 967 2718 971 2719
rect 967 2713 971 2714
rect 1087 2718 1091 2719
rect 1087 2713 1091 2714
rect 1143 2718 1147 2719
rect 1143 2713 1147 2714
rect 1239 2718 1243 2719
rect 1239 2713 1243 2714
rect 1311 2718 1315 2719
rect 1311 2713 1315 2714
rect 1383 2718 1387 2719
rect 1383 2713 1387 2714
rect 1479 2718 1483 2719
rect 1479 2713 1483 2714
rect 1535 2718 1539 2719
rect 1535 2713 1539 2714
rect 1647 2718 1651 2719
rect 1647 2713 1651 2714
rect 1679 2718 1683 2719
rect 1679 2713 1683 2714
rect 1815 2718 1819 2719
rect 1815 2713 1819 2714
rect 1935 2718 1939 2719
rect 1935 2713 1939 2714
rect 112 2690 114 2713
rect 110 2689 116 2690
rect 448 2689 450 2713
rect 616 2689 618 2713
rect 776 2689 778 2713
rect 936 2689 938 2713
rect 1088 2689 1090 2713
rect 1240 2689 1242 2713
rect 1384 2689 1386 2713
rect 1536 2689 1538 2713
rect 1680 2689 1682 2713
rect 1816 2689 1818 2713
rect 1936 2690 1938 2713
rect 1934 2689 1940 2690
rect 110 2685 111 2689
rect 115 2685 116 2689
rect 110 2684 116 2685
rect 446 2688 452 2689
rect 446 2684 447 2688
rect 451 2684 452 2688
rect 446 2683 452 2684
rect 614 2688 620 2689
rect 614 2684 615 2688
rect 619 2684 620 2688
rect 614 2683 620 2684
rect 774 2688 780 2689
rect 774 2684 775 2688
rect 779 2684 780 2688
rect 774 2683 780 2684
rect 934 2688 940 2689
rect 934 2684 935 2688
rect 939 2684 940 2688
rect 934 2683 940 2684
rect 1086 2688 1092 2689
rect 1086 2684 1087 2688
rect 1091 2684 1092 2688
rect 1086 2683 1092 2684
rect 1238 2688 1244 2689
rect 1238 2684 1239 2688
rect 1243 2684 1244 2688
rect 1238 2683 1244 2684
rect 1382 2688 1388 2689
rect 1382 2684 1383 2688
rect 1387 2684 1388 2688
rect 1382 2683 1388 2684
rect 1534 2688 1540 2689
rect 1534 2684 1535 2688
rect 1539 2684 1540 2688
rect 1534 2683 1540 2684
rect 1678 2688 1684 2689
rect 1678 2684 1679 2688
rect 1683 2684 1684 2688
rect 1678 2683 1684 2684
rect 1814 2688 1820 2689
rect 1814 2684 1815 2688
rect 1819 2684 1820 2688
rect 1934 2685 1935 2689
rect 1939 2685 1940 2689
rect 1934 2684 1940 2685
rect 1814 2683 1820 2684
rect 418 2673 424 2674
rect 110 2672 116 2673
rect 110 2668 111 2672
rect 115 2668 116 2672
rect 418 2669 419 2673
rect 423 2669 424 2673
rect 418 2668 424 2669
rect 586 2673 592 2674
rect 586 2669 587 2673
rect 591 2669 592 2673
rect 586 2668 592 2669
rect 746 2673 752 2674
rect 746 2669 747 2673
rect 751 2669 752 2673
rect 746 2668 752 2669
rect 906 2673 912 2674
rect 906 2669 907 2673
rect 911 2669 912 2673
rect 906 2668 912 2669
rect 1058 2673 1064 2674
rect 1058 2669 1059 2673
rect 1063 2669 1064 2673
rect 1058 2668 1064 2669
rect 1210 2673 1216 2674
rect 1210 2669 1211 2673
rect 1215 2669 1216 2673
rect 1210 2668 1216 2669
rect 1354 2673 1360 2674
rect 1354 2669 1355 2673
rect 1359 2669 1360 2673
rect 1354 2668 1360 2669
rect 1506 2673 1512 2674
rect 1506 2669 1507 2673
rect 1511 2669 1512 2673
rect 1506 2668 1512 2669
rect 1650 2673 1656 2674
rect 1650 2669 1651 2673
rect 1655 2669 1656 2673
rect 1650 2668 1656 2669
rect 1786 2673 1792 2674
rect 1786 2669 1787 2673
rect 1791 2669 1792 2673
rect 1786 2668 1792 2669
rect 1934 2672 1940 2673
rect 1934 2668 1935 2672
rect 1939 2668 1940 2672
rect 110 2667 116 2668
rect 112 2603 114 2667
rect 420 2603 422 2668
rect 588 2603 590 2668
rect 748 2603 750 2668
rect 908 2603 910 2668
rect 1060 2603 1062 2668
rect 1212 2603 1214 2668
rect 1356 2603 1358 2668
rect 1508 2603 1510 2668
rect 1652 2603 1654 2668
rect 1788 2603 1790 2668
rect 1934 2667 1940 2668
rect 1936 2603 1938 2667
rect 1976 2639 1978 2930
rect 3136 2639 3138 2931
rect 3272 2639 3274 2931
rect 3408 2639 3410 2931
rect 3544 2639 3546 2931
rect 3680 2639 3682 2931
rect 3798 2930 3804 2931
rect 3800 2639 3802 2930
rect 3858 2929 3864 2930
rect 3838 2928 3844 2929
rect 3838 2924 3839 2928
rect 3843 2924 3844 2928
rect 3858 2925 3859 2929
rect 3863 2925 3864 2929
rect 3858 2924 3864 2925
rect 3994 2929 4000 2930
rect 3994 2925 3995 2929
rect 3999 2925 4000 2929
rect 3994 2924 4000 2925
rect 4146 2929 4152 2930
rect 4146 2925 4147 2929
rect 4151 2925 4152 2929
rect 4146 2924 4152 2925
rect 4362 2929 4368 2930
rect 4362 2925 4363 2929
rect 4367 2925 4368 2929
rect 4362 2924 4368 2925
rect 4610 2929 4616 2930
rect 4610 2925 4611 2929
rect 4615 2925 4616 2929
rect 4610 2924 4616 2925
rect 4890 2929 4896 2930
rect 4890 2925 4891 2929
rect 4895 2925 4896 2929
rect 4890 2924 4896 2925
rect 5194 2929 5200 2930
rect 5194 2925 5195 2929
rect 5199 2925 5200 2929
rect 5194 2924 5200 2925
rect 5498 2929 5504 2930
rect 5498 2925 5499 2929
rect 5503 2925 5504 2929
rect 5498 2924 5504 2925
rect 5662 2928 5668 2929
rect 5662 2924 5663 2928
rect 5667 2924 5668 2928
rect 3838 2923 3844 2924
rect 3840 2863 3842 2923
rect 3860 2863 3862 2924
rect 3996 2863 3998 2924
rect 4148 2863 4150 2924
rect 4364 2863 4366 2924
rect 4612 2863 4614 2924
rect 4892 2863 4894 2924
rect 5196 2863 5198 2924
rect 5500 2863 5502 2924
rect 5662 2923 5668 2924
rect 5664 2863 5666 2923
rect 3839 2862 3843 2863
rect 3839 2857 3843 2858
rect 3859 2862 3863 2863
rect 3859 2857 3863 2858
rect 3995 2862 3999 2863
rect 3995 2857 3999 2858
rect 4131 2862 4135 2863
rect 4131 2857 4135 2858
rect 4147 2862 4151 2863
rect 4147 2857 4151 2858
rect 4267 2862 4271 2863
rect 4267 2857 4271 2858
rect 4363 2862 4367 2863
rect 4363 2857 4367 2858
rect 4403 2862 4407 2863
rect 4403 2857 4407 2858
rect 4539 2862 4543 2863
rect 4539 2857 4543 2858
rect 4611 2862 4615 2863
rect 4611 2857 4615 2858
rect 4675 2862 4679 2863
rect 4675 2857 4679 2858
rect 4811 2862 4815 2863
rect 4811 2857 4815 2858
rect 4891 2862 4895 2863
rect 4891 2857 4895 2858
rect 5195 2862 5199 2863
rect 5195 2857 5199 2858
rect 5499 2862 5503 2863
rect 5499 2857 5503 2858
rect 5663 2862 5667 2863
rect 5663 2857 5667 2858
rect 3840 2797 3842 2857
rect 3838 2796 3844 2797
rect 3860 2796 3862 2857
rect 3996 2796 3998 2857
rect 4132 2796 4134 2857
rect 4268 2796 4270 2857
rect 4404 2796 4406 2857
rect 4540 2796 4542 2857
rect 4676 2796 4678 2857
rect 4812 2796 4814 2857
rect 5664 2797 5666 2857
rect 5662 2796 5668 2797
rect 3838 2792 3839 2796
rect 3843 2792 3844 2796
rect 3838 2791 3844 2792
rect 3858 2795 3864 2796
rect 3858 2791 3859 2795
rect 3863 2791 3864 2795
rect 3858 2790 3864 2791
rect 3994 2795 4000 2796
rect 3994 2791 3995 2795
rect 3999 2791 4000 2795
rect 3994 2790 4000 2791
rect 4130 2795 4136 2796
rect 4130 2791 4131 2795
rect 4135 2791 4136 2795
rect 4130 2790 4136 2791
rect 4266 2795 4272 2796
rect 4266 2791 4267 2795
rect 4271 2791 4272 2795
rect 4266 2790 4272 2791
rect 4402 2795 4408 2796
rect 4402 2791 4403 2795
rect 4407 2791 4408 2795
rect 4402 2790 4408 2791
rect 4538 2795 4544 2796
rect 4538 2791 4539 2795
rect 4543 2791 4544 2795
rect 4538 2790 4544 2791
rect 4674 2795 4680 2796
rect 4674 2791 4675 2795
rect 4679 2791 4680 2795
rect 4674 2790 4680 2791
rect 4810 2795 4816 2796
rect 4810 2791 4811 2795
rect 4815 2791 4816 2795
rect 5662 2792 5663 2796
rect 5667 2792 5668 2796
rect 5662 2791 5668 2792
rect 4810 2790 4816 2791
rect 3886 2780 3892 2781
rect 3838 2779 3844 2780
rect 3838 2775 3839 2779
rect 3843 2775 3844 2779
rect 3886 2776 3887 2780
rect 3891 2776 3892 2780
rect 3886 2775 3892 2776
rect 4022 2780 4028 2781
rect 4022 2776 4023 2780
rect 4027 2776 4028 2780
rect 4022 2775 4028 2776
rect 4158 2780 4164 2781
rect 4158 2776 4159 2780
rect 4163 2776 4164 2780
rect 4158 2775 4164 2776
rect 4294 2780 4300 2781
rect 4294 2776 4295 2780
rect 4299 2776 4300 2780
rect 4294 2775 4300 2776
rect 4430 2780 4436 2781
rect 4430 2776 4431 2780
rect 4435 2776 4436 2780
rect 4430 2775 4436 2776
rect 4566 2780 4572 2781
rect 4566 2776 4567 2780
rect 4571 2776 4572 2780
rect 4566 2775 4572 2776
rect 4702 2780 4708 2781
rect 4702 2776 4703 2780
rect 4707 2776 4708 2780
rect 4702 2775 4708 2776
rect 4838 2780 4844 2781
rect 4838 2776 4839 2780
rect 4843 2776 4844 2780
rect 4838 2775 4844 2776
rect 5662 2779 5668 2780
rect 5662 2775 5663 2779
rect 5667 2775 5668 2779
rect 3838 2774 3844 2775
rect 3840 2735 3842 2774
rect 3888 2735 3890 2775
rect 4024 2735 4026 2775
rect 4160 2735 4162 2775
rect 4296 2735 4298 2775
rect 4432 2735 4434 2775
rect 4568 2735 4570 2775
rect 4704 2735 4706 2775
rect 4840 2735 4842 2775
rect 5662 2774 5668 2775
rect 5664 2735 5666 2774
rect 3839 2734 3843 2735
rect 3839 2729 3843 2730
rect 3887 2734 3891 2735
rect 3887 2729 3891 2730
rect 4023 2734 4027 2735
rect 4023 2729 4027 2730
rect 4159 2734 4163 2735
rect 4159 2729 4163 2730
rect 4295 2734 4299 2735
rect 4295 2729 4299 2730
rect 4431 2734 4435 2735
rect 4431 2729 4435 2730
rect 4567 2734 4571 2735
rect 4567 2729 4571 2730
rect 4703 2734 4707 2735
rect 4703 2729 4707 2730
rect 4711 2734 4715 2735
rect 4711 2729 4715 2730
rect 4839 2734 4843 2735
rect 4839 2729 4843 2730
rect 4879 2734 4883 2735
rect 4879 2729 4883 2730
rect 5063 2734 5067 2735
rect 5063 2729 5067 2730
rect 5255 2734 5259 2735
rect 5255 2729 5259 2730
rect 5447 2734 5451 2735
rect 5447 2729 5451 2730
rect 5663 2734 5667 2735
rect 5663 2729 5667 2730
rect 3840 2706 3842 2729
rect 3838 2705 3844 2706
rect 3888 2705 3890 2729
rect 4024 2705 4026 2729
rect 4160 2705 4162 2729
rect 4296 2705 4298 2729
rect 4432 2705 4434 2729
rect 4568 2705 4570 2729
rect 4712 2705 4714 2729
rect 4880 2705 4882 2729
rect 5064 2705 5066 2729
rect 5256 2705 5258 2729
rect 5448 2705 5450 2729
rect 5664 2706 5666 2729
rect 5662 2705 5668 2706
rect 3838 2701 3839 2705
rect 3843 2701 3844 2705
rect 3838 2700 3844 2701
rect 3886 2704 3892 2705
rect 3886 2700 3887 2704
rect 3891 2700 3892 2704
rect 3886 2699 3892 2700
rect 4022 2704 4028 2705
rect 4022 2700 4023 2704
rect 4027 2700 4028 2704
rect 4022 2699 4028 2700
rect 4158 2704 4164 2705
rect 4158 2700 4159 2704
rect 4163 2700 4164 2704
rect 4158 2699 4164 2700
rect 4294 2704 4300 2705
rect 4294 2700 4295 2704
rect 4299 2700 4300 2704
rect 4294 2699 4300 2700
rect 4430 2704 4436 2705
rect 4430 2700 4431 2704
rect 4435 2700 4436 2704
rect 4430 2699 4436 2700
rect 4566 2704 4572 2705
rect 4566 2700 4567 2704
rect 4571 2700 4572 2704
rect 4566 2699 4572 2700
rect 4710 2704 4716 2705
rect 4710 2700 4711 2704
rect 4715 2700 4716 2704
rect 4710 2699 4716 2700
rect 4878 2704 4884 2705
rect 4878 2700 4879 2704
rect 4883 2700 4884 2704
rect 4878 2699 4884 2700
rect 5062 2704 5068 2705
rect 5062 2700 5063 2704
rect 5067 2700 5068 2704
rect 5062 2699 5068 2700
rect 5254 2704 5260 2705
rect 5254 2700 5255 2704
rect 5259 2700 5260 2704
rect 5254 2699 5260 2700
rect 5446 2704 5452 2705
rect 5446 2700 5447 2704
rect 5451 2700 5452 2704
rect 5662 2701 5663 2705
rect 5667 2701 5668 2705
rect 5662 2700 5668 2701
rect 5446 2699 5452 2700
rect 3858 2689 3864 2690
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3858 2685 3859 2689
rect 3863 2685 3864 2689
rect 3858 2684 3864 2685
rect 3994 2689 4000 2690
rect 3994 2685 3995 2689
rect 3999 2685 4000 2689
rect 3994 2684 4000 2685
rect 4130 2689 4136 2690
rect 4130 2685 4131 2689
rect 4135 2685 4136 2689
rect 4130 2684 4136 2685
rect 4266 2689 4272 2690
rect 4266 2685 4267 2689
rect 4271 2685 4272 2689
rect 4266 2684 4272 2685
rect 4402 2689 4408 2690
rect 4402 2685 4403 2689
rect 4407 2685 4408 2689
rect 4402 2684 4408 2685
rect 4538 2689 4544 2690
rect 4538 2685 4539 2689
rect 4543 2685 4544 2689
rect 4538 2684 4544 2685
rect 4682 2689 4688 2690
rect 4682 2685 4683 2689
rect 4687 2685 4688 2689
rect 4682 2684 4688 2685
rect 4850 2689 4856 2690
rect 4850 2685 4851 2689
rect 4855 2685 4856 2689
rect 4850 2684 4856 2685
rect 5034 2689 5040 2690
rect 5034 2685 5035 2689
rect 5039 2685 5040 2689
rect 5034 2684 5040 2685
rect 5226 2689 5232 2690
rect 5226 2685 5227 2689
rect 5231 2685 5232 2689
rect 5226 2684 5232 2685
rect 5418 2689 5424 2690
rect 5418 2685 5419 2689
rect 5423 2685 5424 2689
rect 5418 2684 5424 2685
rect 5662 2688 5668 2689
rect 5662 2684 5663 2688
rect 5667 2684 5668 2688
rect 3838 2683 3844 2684
rect 1975 2638 1979 2639
rect 1975 2633 1979 2634
rect 3135 2638 3139 2639
rect 3135 2633 3139 2634
rect 3271 2638 3275 2639
rect 3271 2633 3275 2634
rect 3407 2638 3411 2639
rect 3407 2633 3411 2634
rect 3543 2638 3547 2639
rect 3543 2633 3547 2634
rect 3679 2638 3683 2639
rect 3679 2633 3683 2634
rect 3799 2638 3803 2639
rect 3799 2633 3803 2634
rect 1976 2610 1978 2633
rect 1974 2609 1980 2610
rect 3272 2609 3274 2633
rect 3408 2609 3410 2633
rect 3544 2609 3546 2633
rect 3680 2609 3682 2633
rect 3800 2610 3802 2633
rect 3798 2609 3804 2610
rect 1974 2605 1975 2609
rect 1979 2605 1980 2609
rect 1974 2604 1980 2605
rect 3270 2608 3276 2609
rect 3270 2604 3271 2608
rect 3275 2604 3276 2608
rect 3270 2603 3276 2604
rect 3406 2608 3412 2609
rect 3406 2604 3407 2608
rect 3411 2604 3412 2608
rect 3406 2603 3412 2604
rect 3542 2608 3548 2609
rect 3542 2604 3543 2608
rect 3547 2604 3548 2608
rect 3542 2603 3548 2604
rect 3678 2608 3684 2609
rect 3678 2604 3679 2608
rect 3683 2604 3684 2608
rect 3798 2605 3799 2609
rect 3803 2605 3804 2609
rect 3840 2607 3842 2683
rect 3860 2607 3862 2684
rect 3996 2607 3998 2684
rect 4132 2607 4134 2684
rect 4268 2607 4270 2684
rect 4404 2607 4406 2684
rect 4540 2607 4542 2684
rect 4684 2607 4686 2684
rect 4852 2607 4854 2684
rect 5036 2607 5038 2684
rect 5228 2607 5230 2684
rect 5420 2607 5422 2684
rect 5662 2683 5668 2684
rect 5664 2607 5666 2683
rect 3798 2604 3804 2605
rect 3839 2606 3843 2607
rect 3678 2603 3684 2604
rect 111 2602 115 2603
rect 111 2597 115 2598
rect 235 2602 239 2603
rect 235 2597 239 2598
rect 419 2602 423 2603
rect 419 2597 423 2598
rect 435 2602 439 2603
rect 435 2597 439 2598
rect 587 2602 591 2603
rect 587 2597 591 2598
rect 627 2602 631 2603
rect 627 2597 631 2598
rect 747 2602 751 2603
rect 747 2597 751 2598
rect 811 2602 815 2603
rect 811 2597 815 2598
rect 907 2602 911 2603
rect 907 2597 911 2598
rect 987 2602 991 2603
rect 987 2597 991 2598
rect 1059 2602 1063 2603
rect 1059 2597 1063 2598
rect 1155 2602 1159 2603
rect 1155 2597 1159 2598
rect 1211 2602 1215 2603
rect 1211 2597 1215 2598
rect 1323 2602 1327 2603
rect 1323 2597 1327 2598
rect 1355 2602 1359 2603
rect 1355 2597 1359 2598
rect 1483 2602 1487 2603
rect 1483 2597 1487 2598
rect 1507 2602 1511 2603
rect 1507 2597 1511 2598
rect 1643 2602 1647 2603
rect 1643 2597 1647 2598
rect 1651 2602 1655 2603
rect 1651 2597 1655 2598
rect 1787 2602 1791 2603
rect 1787 2597 1791 2598
rect 1935 2602 1939 2603
rect 3839 2601 3843 2602
rect 3859 2606 3863 2607
rect 3859 2601 3863 2602
rect 3995 2606 3999 2607
rect 3995 2601 3999 2602
rect 4131 2606 4135 2607
rect 4131 2601 4135 2602
rect 4179 2606 4183 2607
rect 4179 2601 4183 2602
rect 4267 2606 4271 2607
rect 4267 2601 4271 2602
rect 4395 2606 4399 2607
rect 4395 2601 4399 2602
rect 4403 2606 4407 2607
rect 4403 2601 4407 2602
rect 4539 2606 4543 2607
rect 4539 2601 4543 2602
rect 4643 2606 4647 2607
rect 4643 2601 4647 2602
rect 4683 2606 4687 2607
rect 4683 2601 4687 2602
rect 4851 2606 4855 2607
rect 4851 2601 4855 2602
rect 4907 2606 4911 2607
rect 4907 2601 4911 2602
rect 5035 2606 5039 2607
rect 5035 2601 5039 2602
rect 5187 2606 5191 2607
rect 5187 2601 5191 2602
rect 5227 2606 5231 2607
rect 5227 2601 5231 2602
rect 5419 2606 5423 2607
rect 5419 2601 5423 2602
rect 5467 2606 5471 2607
rect 5467 2601 5471 2602
rect 5663 2606 5667 2607
rect 5663 2601 5667 2602
rect 1935 2597 1939 2598
rect 112 2537 114 2597
rect 110 2536 116 2537
rect 236 2536 238 2597
rect 436 2536 438 2597
rect 628 2536 630 2597
rect 812 2536 814 2597
rect 988 2536 990 2597
rect 1156 2536 1158 2597
rect 1324 2536 1326 2597
rect 1484 2536 1486 2597
rect 1644 2536 1646 2597
rect 1788 2536 1790 2597
rect 1936 2537 1938 2597
rect 3242 2593 3248 2594
rect 1974 2592 1980 2593
rect 1974 2588 1975 2592
rect 1979 2588 1980 2592
rect 3242 2589 3243 2593
rect 3247 2589 3248 2593
rect 3242 2588 3248 2589
rect 3378 2593 3384 2594
rect 3378 2589 3379 2593
rect 3383 2589 3384 2593
rect 3378 2588 3384 2589
rect 3514 2593 3520 2594
rect 3514 2589 3515 2593
rect 3519 2589 3520 2593
rect 3514 2588 3520 2589
rect 3650 2593 3656 2594
rect 3650 2589 3651 2593
rect 3655 2589 3656 2593
rect 3650 2588 3656 2589
rect 3798 2592 3804 2593
rect 3798 2588 3799 2592
rect 3803 2588 3804 2592
rect 1974 2587 1980 2588
rect 1934 2536 1940 2537
rect 110 2532 111 2536
rect 115 2532 116 2536
rect 110 2531 116 2532
rect 234 2535 240 2536
rect 234 2531 235 2535
rect 239 2531 240 2535
rect 234 2530 240 2531
rect 434 2535 440 2536
rect 434 2531 435 2535
rect 439 2531 440 2535
rect 434 2530 440 2531
rect 626 2535 632 2536
rect 626 2531 627 2535
rect 631 2531 632 2535
rect 626 2530 632 2531
rect 810 2535 816 2536
rect 810 2531 811 2535
rect 815 2531 816 2535
rect 810 2530 816 2531
rect 986 2535 992 2536
rect 986 2531 987 2535
rect 991 2531 992 2535
rect 986 2530 992 2531
rect 1154 2535 1160 2536
rect 1154 2531 1155 2535
rect 1159 2531 1160 2535
rect 1154 2530 1160 2531
rect 1322 2535 1328 2536
rect 1322 2531 1323 2535
rect 1327 2531 1328 2535
rect 1322 2530 1328 2531
rect 1482 2535 1488 2536
rect 1482 2531 1483 2535
rect 1487 2531 1488 2535
rect 1482 2530 1488 2531
rect 1642 2535 1648 2536
rect 1642 2531 1643 2535
rect 1647 2531 1648 2535
rect 1642 2530 1648 2531
rect 1786 2535 1792 2536
rect 1786 2531 1787 2535
rect 1791 2531 1792 2535
rect 1934 2532 1935 2536
rect 1939 2532 1940 2536
rect 1934 2531 1940 2532
rect 1786 2530 1792 2531
rect 1976 2527 1978 2587
rect 3244 2527 3246 2588
rect 3380 2527 3382 2588
rect 3516 2527 3518 2588
rect 3652 2527 3654 2588
rect 3798 2587 3804 2588
rect 3800 2527 3802 2587
rect 3840 2541 3842 2601
rect 3838 2540 3844 2541
rect 4180 2540 4182 2601
rect 4396 2540 4398 2601
rect 4644 2540 4646 2601
rect 4908 2540 4910 2601
rect 5188 2540 5190 2601
rect 5468 2540 5470 2601
rect 5664 2541 5666 2601
rect 5662 2540 5668 2541
rect 3838 2536 3839 2540
rect 3843 2536 3844 2540
rect 3838 2535 3844 2536
rect 4178 2539 4184 2540
rect 4178 2535 4179 2539
rect 4183 2535 4184 2539
rect 4178 2534 4184 2535
rect 4394 2539 4400 2540
rect 4394 2535 4395 2539
rect 4399 2535 4400 2539
rect 4394 2534 4400 2535
rect 4642 2539 4648 2540
rect 4642 2535 4643 2539
rect 4647 2535 4648 2539
rect 4642 2534 4648 2535
rect 4906 2539 4912 2540
rect 4906 2535 4907 2539
rect 4911 2535 4912 2539
rect 4906 2534 4912 2535
rect 5186 2539 5192 2540
rect 5186 2535 5187 2539
rect 5191 2535 5192 2539
rect 5186 2534 5192 2535
rect 5466 2539 5472 2540
rect 5466 2535 5467 2539
rect 5471 2535 5472 2539
rect 5662 2536 5663 2540
rect 5667 2536 5668 2540
rect 5662 2535 5668 2536
rect 5466 2534 5472 2535
rect 1975 2526 1979 2527
rect 1975 2521 1979 2522
rect 1995 2526 1999 2527
rect 1995 2521 1999 2522
rect 2251 2526 2255 2527
rect 2251 2521 2255 2522
rect 2523 2526 2527 2527
rect 2523 2521 2527 2522
rect 2771 2526 2775 2527
rect 2771 2521 2775 2522
rect 3003 2526 3007 2527
rect 3003 2521 3007 2522
rect 3227 2526 3231 2527
rect 3227 2521 3231 2522
rect 3243 2526 3247 2527
rect 3243 2521 3247 2522
rect 3379 2526 3383 2527
rect 3379 2521 3383 2522
rect 3451 2526 3455 2527
rect 3451 2521 3455 2522
rect 3515 2526 3519 2527
rect 3515 2521 3519 2522
rect 3651 2526 3655 2527
rect 3651 2521 3655 2522
rect 3799 2526 3803 2527
rect 4206 2524 4212 2525
rect 3799 2521 3803 2522
rect 3838 2523 3844 2524
rect 262 2520 268 2521
rect 110 2519 116 2520
rect 110 2515 111 2519
rect 115 2515 116 2519
rect 262 2516 263 2520
rect 267 2516 268 2520
rect 262 2515 268 2516
rect 462 2520 468 2521
rect 462 2516 463 2520
rect 467 2516 468 2520
rect 462 2515 468 2516
rect 654 2520 660 2521
rect 654 2516 655 2520
rect 659 2516 660 2520
rect 654 2515 660 2516
rect 838 2520 844 2521
rect 838 2516 839 2520
rect 843 2516 844 2520
rect 838 2515 844 2516
rect 1014 2520 1020 2521
rect 1014 2516 1015 2520
rect 1019 2516 1020 2520
rect 1014 2515 1020 2516
rect 1182 2520 1188 2521
rect 1182 2516 1183 2520
rect 1187 2516 1188 2520
rect 1182 2515 1188 2516
rect 1350 2520 1356 2521
rect 1350 2516 1351 2520
rect 1355 2516 1356 2520
rect 1350 2515 1356 2516
rect 1510 2520 1516 2521
rect 1510 2516 1511 2520
rect 1515 2516 1516 2520
rect 1510 2515 1516 2516
rect 1670 2520 1676 2521
rect 1670 2516 1671 2520
rect 1675 2516 1676 2520
rect 1670 2515 1676 2516
rect 1814 2520 1820 2521
rect 1814 2516 1815 2520
rect 1819 2516 1820 2520
rect 1814 2515 1820 2516
rect 1934 2519 1940 2520
rect 1934 2515 1935 2519
rect 1939 2515 1940 2519
rect 110 2514 116 2515
rect 112 2483 114 2514
rect 264 2483 266 2515
rect 464 2483 466 2515
rect 656 2483 658 2515
rect 840 2483 842 2515
rect 1016 2483 1018 2515
rect 1184 2483 1186 2515
rect 1352 2483 1354 2515
rect 1512 2483 1514 2515
rect 1672 2483 1674 2515
rect 1816 2483 1818 2515
rect 1934 2514 1940 2515
rect 1936 2483 1938 2514
rect 111 2482 115 2483
rect 111 2477 115 2478
rect 223 2482 227 2483
rect 223 2477 227 2478
rect 263 2482 267 2483
rect 263 2477 267 2478
rect 423 2482 427 2483
rect 423 2477 427 2478
rect 463 2482 467 2483
rect 463 2477 467 2478
rect 623 2482 627 2483
rect 623 2477 627 2478
rect 655 2482 659 2483
rect 655 2477 659 2478
rect 815 2482 819 2483
rect 815 2477 819 2478
rect 839 2482 843 2483
rect 839 2477 843 2478
rect 1015 2482 1019 2483
rect 1015 2477 1019 2478
rect 1183 2482 1187 2483
rect 1183 2477 1187 2478
rect 1215 2482 1219 2483
rect 1215 2477 1219 2478
rect 1351 2482 1355 2483
rect 1351 2477 1355 2478
rect 1511 2482 1515 2483
rect 1511 2477 1515 2478
rect 1671 2482 1675 2483
rect 1671 2477 1675 2478
rect 1815 2482 1819 2483
rect 1815 2477 1819 2478
rect 1935 2482 1939 2483
rect 1935 2477 1939 2478
rect 112 2454 114 2477
rect 110 2453 116 2454
rect 224 2453 226 2477
rect 424 2453 426 2477
rect 624 2453 626 2477
rect 816 2453 818 2477
rect 1016 2453 1018 2477
rect 1216 2453 1218 2477
rect 1936 2454 1938 2477
rect 1976 2461 1978 2521
rect 1974 2460 1980 2461
rect 1996 2460 1998 2521
rect 2252 2460 2254 2521
rect 2524 2460 2526 2521
rect 2772 2460 2774 2521
rect 3004 2460 3006 2521
rect 3228 2460 3230 2521
rect 3452 2460 3454 2521
rect 3652 2460 3654 2521
rect 3800 2461 3802 2521
rect 3838 2519 3839 2523
rect 3843 2519 3844 2523
rect 4206 2520 4207 2524
rect 4211 2520 4212 2524
rect 4206 2519 4212 2520
rect 4422 2524 4428 2525
rect 4422 2520 4423 2524
rect 4427 2520 4428 2524
rect 4422 2519 4428 2520
rect 4670 2524 4676 2525
rect 4670 2520 4671 2524
rect 4675 2520 4676 2524
rect 4670 2519 4676 2520
rect 4934 2524 4940 2525
rect 4934 2520 4935 2524
rect 4939 2520 4940 2524
rect 4934 2519 4940 2520
rect 5214 2524 5220 2525
rect 5214 2520 5215 2524
rect 5219 2520 5220 2524
rect 5214 2519 5220 2520
rect 5494 2524 5500 2525
rect 5494 2520 5495 2524
rect 5499 2520 5500 2524
rect 5494 2519 5500 2520
rect 5662 2523 5668 2524
rect 5662 2519 5663 2523
rect 5667 2519 5668 2523
rect 3838 2518 3844 2519
rect 3840 2495 3842 2518
rect 4208 2495 4210 2519
rect 4424 2495 4426 2519
rect 4672 2495 4674 2519
rect 4936 2495 4938 2519
rect 5216 2495 5218 2519
rect 5496 2495 5498 2519
rect 5662 2518 5668 2519
rect 5664 2495 5666 2518
rect 3839 2494 3843 2495
rect 3839 2489 3843 2490
rect 4207 2494 4211 2495
rect 4207 2489 4211 2490
rect 4423 2494 4427 2495
rect 4423 2489 4427 2490
rect 4535 2494 4539 2495
rect 4535 2489 4539 2490
rect 4671 2494 4675 2495
rect 4671 2489 4675 2490
rect 4759 2494 4763 2495
rect 4759 2489 4763 2490
rect 4935 2494 4939 2495
rect 4935 2489 4939 2490
rect 4983 2494 4987 2495
rect 4983 2489 4987 2490
rect 5215 2494 5219 2495
rect 5215 2489 5219 2490
rect 5447 2494 5451 2495
rect 5447 2489 5451 2490
rect 5495 2494 5499 2495
rect 5495 2489 5499 2490
rect 5663 2494 5667 2495
rect 5663 2489 5667 2490
rect 3840 2466 3842 2489
rect 3838 2465 3844 2466
rect 4536 2465 4538 2489
rect 4760 2465 4762 2489
rect 4984 2465 4986 2489
rect 5216 2465 5218 2489
rect 5448 2465 5450 2489
rect 5664 2466 5666 2489
rect 5662 2465 5668 2466
rect 3838 2461 3839 2465
rect 3843 2461 3844 2465
rect 3798 2460 3804 2461
rect 3838 2460 3844 2461
rect 4534 2464 4540 2465
rect 4534 2460 4535 2464
rect 4539 2460 4540 2464
rect 1974 2456 1975 2460
rect 1979 2456 1980 2460
rect 1974 2455 1980 2456
rect 1994 2459 2000 2460
rect 1994 2455 1995 2459
rect 1999 2455 2000 2459
rect 1994 2454 2000 2455
rect 2250 2459 2256 2460
rect 2250 2455 2251 2459
rect 2255 2455 2256 2459
rect 2250 2454 2256 2455
rect 2522 2459 2528 2460
rect 2522 2455 2523 2459
rect 2527 2455 2528 2459
rect 2522 2454 2528 2455
rect 2770 2459 2776 2460
rect 2770 2455 2771 2459
rect 2775 2455 2776 2459
rect 2770 2454 2776 2455
rect 3002 2459 3008 2460
rect 3002 2455 3003 2459
rect 3007 2455 3008 2459
rect 3002 2454 3008 2455
rect 3226 2459 3232 2460
rect 3226 2455 3227 2459
rect 3231 2455 3232 2459
rect 3226 2454 3232 2455
rect 3450 2459 3456 2460
rect 3450 2455 3451 2459
rect 3455 2455 3456 2459
rect 3450 2454 3456 2455
rect 3650 2459 3656 2460
rect 3650 2455 3651 2459
rect 3655 2455 3656 2459
rect 3798 2456 3799 2460
rect 3803 2456 3804 2460
rect 4534 2459 4540 2460
rect 4758 2464 4764 2465
rect 4758 2460 4759 2464
rect 4763 2460 4764 2464
rect 4758 2459 4764 2460
rect 4982 2464 4988 2465
rect 4982 2460 4983 2464
rect 4987 2460 4988 2464
rect 4982 2459 4988 2460
rect 5214 2464 5220 2465
rect 5214 2460 5215 2464
rect 5219 2460 5220 2464
rect 5214 2459 5220 2460
rect 5446 2464 5452 2465
rect 5446 2460 5447 2464
rect 5451 2460 5452 2464
rect 5662 2461 5663 2465
rect 5667 2461 5668 2465
rect 5662 2460 5668 2461
rect 5446 2459 5452 2460
rect 3798 2455 3804 2456
rect 3650 2454 3656 2455
rect 1934 2453 1940 2454
rect 110 2449 111 2453
rect 115 2449 116 2453
rect 110 2448 116 2449
rect 222 2452 228 2453
rect 222 2448 223 2452
rect 227 2448 228 2452
rect 222 2447 228 2448
rect 422 2452 428 2453
rect 422 2448 423 2452
rect 427 2448 428 2452
rect 422 2447 428 2448
rect 622 2452 628 2453
rect 622 2448 623 2452
rect 627 2448 628 2452
rect 622 2447 628 2448
rect 814 2452 820 2453
rect 814 2448 815 2452
rect 819 2448 820 2452
rect 814 2447 820 2448
rect 1014 2452 1020 2453
rect 1014 2448 1015 2452
rect 1019 2448 1020 2452
rect 1014 2447 1020 2448
rect 1214 2452 1220 2453
rect 1214 2448 1215 2452
rect 1219 2448 1220 2452
rect 1934 2449 1935 2453
rect 1939 2449 1940 2453
rect 4506 2449 4512 2450
rect 1934 2448 1940 2449
rect 3838 2448 3844 2449
rect 1214 2447 1220 2448
rect 2022 2444 2028 2445
rect 1974 2443 1980 2444
rect 1974 2439 1975 2443
rect 1979 2439 1980 2443
rect 2022 2440 2023 2444
rect 2027 2440 2028 2444
rect 2022 2439 2028 2440
rect 2278 2444 2284 2445
rect 2278 2440 2279 2444
rect 2283 2440 2284 2444
rect 2278 2439 2284 2440
rect 2550 2444 2556 2445
rect 2550 2440 2551 2444
rect 2555 2440 2556 2444
rect 2550 2439 2556 2440
rect 2798 2444 2804 2445
rect 2798 2440 2799 2444
rect 2803 2440 2804 2444
rect 2798 2439 2804 2440
rect 3030 2444 3036 2445
rect 3030 2440 3031 2444
rect 3035 2440 3036 2444
rect 3030 2439 3036 2440
rect 3254 2444 3260 2445
rect 3254 2440 3255 2444
rect 3259 2440 3260 2444
rect 3254 2439 3260 2440
rect 3478 2444 3484 2445
rect 3478 2440 3479 2444
rect 3483 2440 3484 2444
rect 3478 2439 3484 2440
rect 3678 2444 3684 2445
rect 3838 2444 3839 2448
rect 3843 2444 3844 2448
rect 4506 2445 4507 2449
rect 4511 2445 4512 2449
rect 4506 2444 4512 2445
rect 4730 2449 4736 2450
rect 4730 2445 4731 2449
rect 4735 2445 4736 2449
rect 4730 2444 4736 2445
rect 4954 2449 4960 2450
rect 4954 2445 4955 2449
rect 4959 2445 4960 2449
rect 4954 2444 4960 2445
rect 5186 2449 5192 2450
rect 5186 2445 5187 2449
rect 5191 2445 5192 2449
rect 5186 2444 5192 2445
rect 5418 2449 5424 2450
rect 5418 2445 5419 2449
rect 5423 2445 5424 2449
rect 5418 2444 5424 2445
rect 5662 2448 5668 2449
rect 5662 2444 5663 2448
rect 5667 2444 5668 2448
rect 3678 2440 3679 2444
rect 3683 2440 3684 2444
rect 3678 2439 3684 2440
rect 3798 2443 3804 2444
rect 3838 2443 3844 2444
rect 3798 2439 3799 2443
rect 3803 2439 3804 2443
rect 1974 2438 1980 2439
rect 194 2437 200 2438
rect 110 2436 116 2437
rect 110 2432 111 2436
rect 115 2432 116 2436
rect 194 2433 195 2437
rect 199 2433 200 2437
rect 194 2432 200 2433
rect 394 2437 400 2438
rect 394 2433 395 2437
rect 399 2433 400 2437
rect 394 2432 400 2433
rect 594 2437 600 2438
rect 594 2433 595 2437
rect 599 2433 600 2437
rect 594 2432 600 2433
rect 786 2437 792 2438
rect 786 2433 787 2437
rect 791 2433 792 2437
rect 786 2432 792 2433
rect 986 2437 992 2438
rect 986 2433 987 2437
rect 991 2433 992 2437
rect 986 2432 992 2433
rect 1186 2437 1192 2438
rect 1186 2433 1187 2437
rect 1191 2433 1192 2437
rect 1186 2432 1192 2433
rect 1934 2436 1940 2437
rect 1934 2432 1935 2436
rect 1939 2432 1940 2436
rect 110 2431 116 2432
rect 112 2359 114 2431
rect 196 2359 198 2432
rect 396 2359 398 2432
rect 596 2359 598 2432
rect 788 2359 790 2432
rect 988 2359 990 2432
rect 1188 2359 1190 2432
rect 1934 2431 1940 2432
rect 1936 2359 1938 2431
rect 1976 2415 1978 2438
rect 2024 2415 2026 2439
rect 2280 2415 2282 2439
rect 2552 2415 2554 2439
rect 2800 2415 2802 2439
rect 3032 2415 3034 2439
rect 3256 2415 3258 2439
rect 3480 2415 3482 2439
rect 3680 2415 3682 2439
rect 3798 2438 3804 2439
rect 3800 2415 3802 2438
rect 1975 2414 1979 2415
rect 1975 2409 1979 2410
rect 2023 2414 2027 2415
rect 2023 2409 2027 2410
rect 2055 2414 2059 2415
rect 2055 2409 2059 2410
rect 2215 2414 2219 2415
rect 2215 2409 2219 2410
rect 2279 2414 2283 2415
rect 2279 2409 2283 2410
rect 2375 2414 2379 2415
rect 2375 2409 2379 2410
rect 2543 2414 2547 2415
rect 2543 2409 2547 2410
rect 2551 2414 2555 2415
rect 2551 2409 2555 2410
rect 2711 2414 2715 2415
rect 2711 2409 2715 2410
rect 2799 2414 2803 2415
rect 2799 2409 2803 2410
rect 2871 2414 2875 2415
rect 2871 2409 2875 2410
rect 3031 2414 3035 2415
rect 3031 2409 3035 2410
rect 3191 2414 3195 2415
rect 3191 2409 3195 2410
rect 3255 2414 3259 2415
rect 3255 2409 3259 2410
rect 3359 2414 3363 2415
rect 3359 2409 3363 2410
rect 3479 2414 3483 2415
rect 3479 2409 3483 2410
rect 3527 2414 3531 2415
rect 3527 2409 3531 2410
rect 3679 2414 3683 2415
rect 3679 2409 3683 2410
rect 3799 2414 3803 2415
rect 3799 2409 3803 2410
rect 1976 2386 1978 2409
rect 1974 2385 1980 2386
rect 2056 2385 2058 2409
rect 2216 2385 2218 2409
rect 2376 2385 2378 2409
rect 2544 2385 2546 2409
rect 2712 2385 2714 2409
rect 2872 2385 2874 2409
rect 3032 2385 3034 2409
rect 3192 2385 3194 2409
rect 3360 2385 3362 2409
rect 3528 2385 3530 2409
rect 3800 2386 3802 2409
rect 3798 2385 3804 2386
rect 1974 2381 1975 2385
rect 1979 2381 1980 2385
rect 1974 2380 1980 2381
rect 2054 2384 2060 2385
rect 2054 2380 2055 2384
rect 2059 2380 2060 2384
rect 2054 2379 2060 2380
rect 2214 2384 2220 2385
rect 2214 2380 2215 2384
rect 2219 2380 2220 2384
rect 2214 2379 2220 2380
rect 2374 2384 2380 2385
rect 2374 2380 2375 2384
rect 2379 2380 2380 2384
rect 2374 2379 2380 2380
rect 2542 2384 2548 2385
rect 2542 2380 2543 2384
rect 2547 2380 2548 2384
rect 2542 2379 2548 2380
rect 2710 2384 2716 2385
rect 2710 2380 2711 2384
rect 2715 2380 2716 2384
rect 2710 2379 2716 2380
rect 2870 2384 2876 2385
rect 2870 2380 2871 2384
rect 2875 2380 2876 2384
rect 2870 2379 2876 2380
rect 3030 2384 3036 2385
rect 3030 2380 3031 2384
rect 3035 2380 3036 2384
rect 3030 2379 3036 2380
rect 3190 2384 3196 2385
rect 3190 2380 3191 2384
rect 3195 2380 3196 2384
rect 3190 2379 3196 2380
rect 3358 2384 3364 2385
rect 3358 2380 3359 2384
rect 3363 2380 3364 2384
rect 3358 2379 3364 2380
rect 3526 2384 3532 2385
rect 3526 2380 3527 2384
rect 3531 2380 3532 2384
rect 3798 2381 3799 2385
rect 3803 2381 3804 2385
rect 3840 2383 3842 2443
rect 4508 2383 4510 2444
rect 4732 2383 4734 2444
rect 4956 2383 4958 2444
rect 5188 2383 5190 2444
rect 5420 2383 5422 2444
rect 5662 2443 5668 2444
rect 5664 2383 5666 2443
rect 3798 2380 3804 2381
rect 3839 2382 3843 2383
rect 3526 2379 3532 2380
rect 3839 2377 3843 2378
rect 4507 2382 4511 2383
rect 4507 2377 4511 2378
rect 4707 2382 4711 2383
rect 4707 2377 4711 2378
rect 4731 2382 4735 2383
rect 4731 2377 4735 2378
rect 4867 2382 4871 2383
rect 4867 2377 4871 2378
rect 4955 2382 4959 2383
rect 4955 2377 4959 2378
rect 5027 2382 5031 2383
rect 5027 2377 5031 2378
rect 5187 2382 5191 2383
rect 5187 2377 5191 2378
rect 5347 2382 5351 2383
rect 5347 2377 5351 2378
rect 5419 2382 5423 2383
rect 5419 2377 5423 2378
rect 5515 2382 5519 2383
rect 5515 2377 5519 2378
rect 5663 2382 5667 2383
rect 5663 2377 5667 2378
rect 2026 2369 2032 2370
rect 1974 2368 1980 2369
rect 1974 2364 1975 2368
rect 1979 2364 1980 2368
rect 2026 2365 2027 2369
rect 2031 2365 2032 2369
rect 2026 2364 2032 2365
rect 2186 2369 2192 2370
rect 2186 2365 2187 2369
rect 2191 2365 2192 2369
rect 2186 2364 2192 2365
rect 2346 2369 2352 2370
rect 2346 2365 2347 2369
rect 2351 2365 2352 2369
rect 2346 2364 2352 2365
rect 2514 2369 2520 2370
rect 2514 2365 2515 2369
rect 2519 2365 2520 2369
rect 2514 2364 2520 2365
rect 2682 2369 2688 2370
rect 2682 2365 2683 2369
rect 2687 2365 2688 2369
rect 2682 2364 2688 2365
rect 2842 2369 2848 2370
rect 2842 2365 2843 2369
rect 2847 2365 2848 2369
rect 2842 2364 2848 2365
rect 3002 2369 3008 2370
rect 3002 2365 3003 2369
rect 3007 2365 3008 2369
rect 3002 2364 3008 2365
rect 3162 2369 3168 2370
rect 3162 2365 3163 2369
rect 3167 2365 3168 2369
rect 3162 2364 3168 2365
rect 3330 2369 3336 2370
rect 3330 2365 3331 2369
rect 3335 2365 3336 2369
rect 3330 2364 3336 2365
rect 3498 2369 3504 2370
rect 3498 2365 3499 2369
rect 3503 2365 3504 2369
rect 3498 2364 3504 2365
rect 3798 2368 3804 2369
rect 3798 2364 3799 2368
rect 3803 2364 3804 2368
rect 1974 2363 1980 2364
rect 111 2358 115 2359
rect 111 2353 115 2354
rect 131 2358 135 2359
rect 131 2353 135 2354
rect 195 2358 199 2359
rect 195 2353 199 2354
rect 291 2358 295 2359
rect 291 2353 295 2354
rect 395 2358 399 2359
rect 395 2353 399 2354
rect 483 2358 487 2359
rect 483 2353 487 2354
rect 595 2358 599 2359
rect 595 2353 599 2354
rect 675 2358 679 2359
rect 675 2353 679 2354
rect 787 2358 791 2359
rect 787 2353 791 2354
rect 867 2358 871 2359
rect 867 2353 871 2354
rect 987 2358 991 2359
rect 987 2353 991 2354
rect 1187 2358 1191 2359
rect 1187 2353 1191 2354
rect 1935 2358 1939 2359
rect 1935 2353 1939 2354
rect 112 2293 114 2353
rect 110 2292 116 2293
rect 132 2292 134 2353
rect 292 2292 294 2353
rect 484 2292 486 2353
rect 676 2292 678 2353
rect 868 2292 870 2353
rect 1936 2293 1938 2353
rect 1976 2295 1978 2363
rect 2028 2295 2030 2364
rect 2188 2295 2190 2364
rect 2348 2295 2350 2364
rect 2516 2295 2518 2364
rect 2684 2295 2686 2364
rect 2844 2295 2846 2364
rect 3004 2295 3006 2364
rect 3164 2295 3166 2364
rect 3332 2295 3334 2364
rect 3500 2295 3502 2364
rect 3798 2363 3804 2364
rect 3800 2295 3802 2363
rect 3840 2317 3842 2377
rect 3838 2316 3844 2317
rect 4708 2316 4710 2377
rect 4868 2316 4870 2377
rect 5028 2316 5030 2377
rect 5188 2316 5190 2377
rect 5348 2316 5350 2377
rect 5516 2316 5518 2377
rect 5664 2317 5666 2377
rect 5662 2316 5668 2317
rect 3838 2312 3839 2316
rect 3843 2312 3844 2316
rect 3838 2311 3844 2312
rect 4706 2315 4712 2316
rect 4706 2311 4707 2315
rect 4711 2311 4712 2315
rect 4706 2310 4712 2311
rect 4866 2315 4872 2316
rect 4866 2311 4867 2315
rect 4871 2311 4872 2315
rect 4866 2310 4872 2311
rect 5026 2315 5032 2316
rect 5026 2311 5027 2315
rect 5031 2311 5032 2315
rect 5026 2310 5032 2311
rect 5186 2315 5192 2316
rect 5186 2311 5187 2315
rect 5191 2311 5192 2315
rect 5186 2310 5192 2311
rect 5346 2315 5352 2316
rect 5346 2311 5347 2315
rect 5351 2311 5352 2315
rect 5346 2310 5352 2311
rect 5514 2315 5520 2316
rect 5514 2311 5515 2315
rect 5519 2311 5520 2315
rect 5662 2312 5663 2316
rect 5667 2312 5668 2316
rect 5662 2311 5668 2312
rect 5514 2310 5520 2311
rect 4734 2300 4740 2301
rect 3838 2299 3844 2300
rect 3838 2295 3839 2299
rect 3843 2295 3844 2299
rect 4734 2296 4735 2300
rect 4739 2296 4740 2300
rect 4734 2295 4740 2296
rect 4894 2300 4900 2301
rect 4894 2296 4895 2300
rect 4899 2296 4900 2300
rect 4894 2295 4900 2296
rect 5054 2300 5060 2301
rect 5054 2296 5055 2300
rect 5059 2296 5060 2300
rect 5054 2295 5060 2296
rect 5214 2300 5220 2301
rect 5214 2296 5215 2300
rect 5219 2296 5220 2300
rect 5214 2295 5220 2296
rect 5374 2300 5380 2301
rect 5374 2296 5375 2300
rect 5379 2296 5380 2300
rect 5374 2295 5380 2296
rect 5542 2300 5548 2301
rect 5542 2296 5543 2300
rect 5547 2296 5548 2300
rect 5542 2295 5548 2296
rect 5662 2299 5668 2300
rect 5662 2295 5663 2299
rect 5667 2295 5668 2299
rect 1975 2294 1979 2295
rect 1934 2292 1940 2293
rect 110 2288 111 2292
rect 115 2288 116 2292
rect 110 2287 116 2288
rect 130 2291 136 2292
rect 130 2287 131 2291
rect 135 2287 136 2291
rect 130 2286 136 2287
rect 290 2291 296 2292
rect 290 2287 291 2291
rect 295 2287 296 2291
rect 290 2286 296 2287
rect 482 2291 488 2292
rect 482 2287 483 2291
rect 487 2287 488 2291
rect 482 2286 488 2287
rect 674 2291 680 2292
rect 674 2287 675 2291
rect 679 2287 680 2291
rect 674 2286 680 2287
rect 866 2291 872 2292
rect 866 2287 867 2291
rect 871 2287 872 2291
rect 1934 2288 1935 2292
rect 1939 2288 1940 2292
rect 1975 2289 1979 2290
rect 2027 2294 2031 2295
rect 2027 2289 2031 2290
rect 2139 2294 2143 2295
rect 2139 2289 2143 2290
rect 2187 2294 2191 2295
rect 2187 2289 2191 2290
rect 2275 2294 2279 2295
rect 2275 2289 2279 2290
rect 2347 2294 2351 2295
rect 2347 2289 2351 2290
rect 2411 2294 2415 2295
rect 2411 2289 2415 2290
rect 2515 2294 2519 2295
rect 2515 2289 2519 2290
rect 2547 2294 2551 2295
rect 2547 2289 2551 2290
rect 2683 2294 2687 2295
rect 2683 2289 2687 2290
rect 2819 2294 2823 2295
rect 2819 2289 2823 2290
rect 2843 2294 2847 2295
rect 2843 2289 2847 2290
rect 2955 2294 2959 2295
rect 2955 2289 2959 2290
rect 3003 2294 3007 2295
rect 3003 2289 3007 2290
rect 3091 2294 3095 2295
rect 3091 2289 3095 2290
rect 3163 2294 3167 2295
rect 3163 2289 3167 2290
rect 3227 2294 3231 2295
rect 3227 2289 3231 2290
rect 3331 2294 3335 2295
rect 3331 2289 3335 2290
rect 3363 2294 3367 2295
rect 3363 2289 3367 2290
rect 3499 2294 3503 2295
rect 3499 2289 3503 2290
rect 3799 2294 3803 2295
rect 3838 2294 3844 2295
rect 3799 2289 3803 2290
rect 1934 2287 1940 2288
rect 866 2286 872 2287
rect 158 2276 164 2277
rect 110 2275 116 2276
rect 110 2271 111 2275
rect 115 2271 116 2275
rect 158 2272 159 2276
rect 163 2272 164 2276
rect 158 2271 164 2272
rect 318 2276 324 2277
rect 318 2272 319 2276
rect 323 2272 324 2276
rect 318 2271 324 2272
rect 510 2276 516 2277
rect 510 2272 511 2276
rect 515 2272 516 2276
rect 510 2271 516 2272
rect 702 2276 708 2277
rect 702 2272 703 2276
rect 707 2272 708 2276
rect 702 2271 708 2272
rect 894 2276 900 2277
rect 894 2272 895 2276
rect 899 2272 900 2276
rect 894 2271 900 2272
rect 1934 2275 1940 2276
rect 1934 2271 1935 2275
rect 1939 2271 1940 2275
rect 110 2270 116 2271
rect 112 2247 114 2270
rect 160 2247 162 2271
rect 320 2247 322 2271
rect 512 2247 514 2271
rect 704 2247 706 2271
rect 896 2247 898 2271
rect 1934 2270 1940 2271
rect 1936 2247 1938 2270
rect 111 2246 115 2247
rect 111 2241 115 2242
rect 159 2246 163 2247
rect 159 2241 163 2242
rect 295 2246 299 2247
rect 295 2241 299 2242
rect 319 2246 323 2247
rect 319 2241 323 2242
rect 439 2246 443 2247
rect 439 2241 443 2242
rect 511 2246 515 2247
rect 511 2241 515 2242
rect 591 2246 595 2247
rect 591 2241 595 2242
rect 703 2246 707 2247
rect 703 2241 707 2242
rect 743 2246 747 2247
rect 743 2241 747 2242
rect 895 2246 899 2247
rect 895 2241 899 2242
rect 1935 2246 1939 2247
rect 1935 2241 1939 2242
rect 112 2218 114 2241
rect 110 2217 116 2218
rect 160 2217 162 2241
rect 296 2217 298 2241
rect 440 2217 442 2241
rect 592 2217 594 2241
rect 744 2217 746 2241
rect 1936 2218 1938 2241
rect 1976 2229 1978 2289
rect 1974 2228 1980 2229
rect 2140 2228 2142 2289
rect 2276 2228 2278 2289
rect 2412 2228 2414 2289
rect 2548 2228 2550 2289
rect 2684 2228 2686 2289
rect 2820 2228 2822 2289
rect 2956 2228 2958 2289
rect 3092 2228 3094 2289
rect 3228 2228 3230 2289
rect 3364 2228 3366 2289
rect 3800 2229 3802 2289
rect 3840 2259 3842 2294
rect 4736 2259 4738 2295
rect 4896 2259 4898 2295
rect 5056 2259 5058 2295
rect 5216 2259 5218 2295
rect 5376 2259 5378 2295
rect 5544 2259 5546 2295
rect 5662 2294 5668 2295
rect 5664 2259 5666 2294
rect 3839 2258 3843 2259
rect 3839 2253 3843 2254
rect 4735 2258 4739 2259
rect 4735 2253 4739 2254
rect 4887 2258 4891 2259
rect 4887 2253 4891 2254
rect 4895 2258 4899 2259
rect 4895 2253 4899 2254
rect 5047 2258 5051 2259
rect 5047 2253 5051 2254
rect 5055 2258 5059 2259
rect 5055 2253 5059 2254
rect 5215 2258 5219 2259
rect 5215 2253 5219 2254
rect 5375 2258 5379 2259
rect 5375 2253 5379 2254
rect 5391 2258 5395 2259
rect 5391 2253 5395 2254
rect 5543 2258 5547 2259
rect 5543 2253 5547 2254
rect 5663 2258 5667 2259
rect 5663 2253 5667 2254
rect 3840 2230 3842 2253
rect 3838 2229 3844 2230
rect 4736 2229 4738 2253
rect 4888 2229 4890 2253
rect 5048 2229 5050 2253
rect 5216 2229 5218 2253
rect 5392 2229 5394 2253
rect 5544 2229 5546 2253
rect 5664 2230 5666 2253
rect 5662 2229 5668 2230
rect 3798 2228 3804 2229
rect 1974 2224 1975 2228
rect 1979 2224 1980 2228
rect 1974 2223 1980 2224
rect 2138 2227 2144 2228
rect 2138 2223 2139 2227
rect 2143 2223 2144 2227
rect 2138 2222 2144 2223
rect 2274 2227 2280 2228
rect 2274 2223 2275 2227
rect 2279 2223 2280 2227
rect 2274 2222 2280 2223
rect 2410 2227 2416 2228
rect 2410 2223 2411 2227
rect 2415 2223 2416 2227
rect 2410 2222 2416 2223
rect 2546 2227 2552 2228
rect 2546 2223 2547 2227
rect 2551 2223 2552 2227
rect 2546 2222 2552 2223
rect 2682 2227 2688 2228
rect 2682 2223 2683 2227
rect 2687 2223 2688 2227
rect 2682 2222 2688 2223
rect 2818 2227 2824 2228
rect 2818 2223 2819 2227
rect 2823 2223 2824 2227
rect 2818 2222 2824 2223
rect 2954 2227 2960 2228
rect 2954 2223 2955 2227
rect 2959 2223 2960 2227
rect 2954 2222 2960 2223
rect 3090 2227 3096 2228
rect 3090 2223 3091 2227
rect 3095 2223 3096 2227
rect 3090 2222 3096 2223
rect 3226 2227 3232 2228
rect 3226 2223 3227 2227
rect 3231 2223 3232 2227
rect 3226 2222 3232 2223
rect 3362 2227 3368 2228
rect 3362 2223 3363 2227
rect 3367 2223 3368 2227
rect 3798 2224 3799 2228
rect 3803 2224 3804 2228
rect 3838 2225 3839 2229
rect 3843 2225 3844 2229
rect 3838 2224 3844 2225
rect 4734 2228 4740 2229
rect 4734 2224 4735 2228
rect 4739 2224 4740 2228
rect 3798 2223 3804 2224
rect 4734 2223 4740 2224
rect 4886 2228 4892 2229
rect 4886 2224 4887 2228
rect 4891 2224 4892 2228
rect 4886 2223 4892 2224
rect 5046 2228 5052 2229
rect 5046 2224 5047 2228
rect 5051 2224 5052 2228
rect 5046 2223 5052 2224
rect 5214 2228 5220 2229
rect 5214 2224 5215 2228
rect 5219 2224 5220 2228
rect 5214 2223 5220 2224
rect 5390 2228 5396 2229
rect 5390 2224 5391 2228
rect 5395 2224 5396 2228
rect 5390 2223 5396 2224
rect 5542 2228 5548 2229
rect 5542 2224 5543 2228
rect 5547 2224 5548 2228
rect 5662 2225 5663 2229
rect 5667 2225 5668 2229
rect 5662 2224 5668 2225
rect 5542 2223 5548 2224
rect 3362 2222 3368 2223
rect 1934 2217 1940 2218
rect 110 2213 111 2217
rect 115 2213 116 2217
rect 110 2212 116 2213
rect 158 2216 164 2217
rect 158 2212 159 2216
rect 163 2212 164 2216
rect 158 2211 164 2212
rect 294 2216 300 2217
rect 294 2212 295 2216
rect 299 2212 300 2216
rect 294 2211 300 2212
rect 438 2216 444 2217
rect 438 2212 439 2216
rect 443 2212 444 2216
rect 438 2211 444 2212
rect 590 2216 596 2217
rect 590 2212 591 2216
rect 595 2212 596 2216
rect 590 2211 596 2212
rect 742 2216 748 2217
rect 742 2212 743 2216
rect 747 2212 748 2216
rect 1934 2213 1935 2217
rect 1939 2213 1940 2217
rect 4706 2213 4712 2214
rect 1934 2212 1940 2213
rect 2166 2212 2172 2213
rect 742 2211 748 2212
rect 1974 2211 1980 2212
rect 1974 2207 1975 2211
rect 1979 2207 1980 2211
rect 2166 2208 2167 2212
rect 2171 2208 2172 2212
rect 2166 2207 2172 2208
rect 2302 2212 2308 2213
rect 2302 2208 2303 2212
rect 2307 2208 2308 2212
rect 2302 2207 2308 2208
rect 2438 2212 2444 2213
rect 2438 2208 2439 2212
rect 2443 2208 2444 2212
rect 2438 2207 2444 2208
rect 2574 2212 2580 2213
rect 2574 2208 2575 2212
rect 2579 2208 2580 2212
rect 2574 2207 2580 2208
rect 2710 2212 2716 2213
rect 2710 2208 2711 2212
rect 2715 2208 2716 2212
rect 2710 2207 2716 2208
rect 2846 2212 2852 2213
rect 2846 2208 2847 2212
rect 2851 2208 2852 2212
rect 2846 2207 2852 2208
rect 2982 2212 2988 2213
rect 2982 2208 2983 2212
rect 2987 2208 2988 2212
rect 2982 2207 2988 2208
rect 3118 2212 3124 2213
rect 3118 2208 3119 2212
rect 3123 2208 3124 2212
rect 3118 2207 3124 2208
rect 3254 2212 3260 2213
rect 3254 2208 3255 2212
rect 3259 2208 3260 2212
rect 3254 2207 3260 2208
rect 3390 2212 3396 2213
rect 3838 2212 3844 2213
rect 3390 2208 3391 2212
rect 3395 2208 3396 2212
rect 3390 2207 3396 2208
rect 3798 2211 3804 2212
rect 3798 2207 3799 2211
rect 3803 2207 3804 2211
rect 3838 2208 3839 2212
rect 3843 2208 3844 2212
rect 4706 2209 4707 2213
rect 4711 2209 4712 2213
rect 4706 2208 4712 2209
rect 4858 2213 4864 2214
rect 4858 2209 4859 2213
rect 4863 2209 4864 2213
rect 4858 2208 4864 2209
rect 5018 2213 5024 2214
rect 5018 2209 5019 2213
rect 5023 2209 5024 2213
rect 5018 2208 5024 2209
rect 5186 2213 5192 2214
rect 5186 2209 5187 2213
rect 5191 2209 5192 2213
rect 5186 2208 5192 2209
rect 5362 2213 5368 2214
rect 5362 2209 5363 2213
rect 5367 2209 5368 2213
rect 5362 2208 5368 2209
rect 5514 2213 5520 2214
rect 5514 2209 5515 2213
rect 5519 2209 5520 2213
rect 5514 2208 5520 2209
rect 5662 2212 5668 2213
rect 5662 2208 5663 2212
rect 5667 2208 5668 2212
rect 3838 2207 3844 2208
rect 1974 2206 1980 2207
rect 130 2201 136 2202
rect 110 2200 116 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 130 2197 131 2201
rect 135 2197 136 2201
rect 130 2196 136 2197
rect 266 2201 272 2202
rect 266 2197 267 2201
rect 271 2197 272 2201
rect 266 2196 272 2197
rect 410 2201 416 2202
rect 410 2197 411 2201
rect 415 2197 416 2201
rect 410 2196 416 2197
rect 562 2201 568 2202
rect 562 2197 563 2201
rect 567 2197 568 2201
rect 562 2196 568 2197
rect 714 2201 720 2202
rect 714 2197 715 2201
rect 719 2197 720 2201
rect 714 2196 720 2197
rect 1934 2200 1940 2201
rect 1934 2196 1935 2200
rect 1939 2196 1940 2200
rect 110 2195 116 2196
rect 112 2135 114 2195
rect 132 2135 134 2196
rect 268 2135 270 2196
rect 412 2135 414 2196
rect 564 2135 566 2196
rect 716 2135 718 2196
rect 1934 2195 1940 2196
rect 1936 2135 1938 2195
rect 1976 2179 1978 2206
rect 2168 2179 2170 2207
rect 2304 2179 2306 2207
rect 2440 2179 2442 2207
rect 2576 2179 2578 2207
rect 2712 2179 2714 2207
rect 2848 2179 2850 2207
rect 2984 2179 2986 2207
rect 3120 2179 3122 2207
rect 3256 2179 3258 2207
rect 3392 2179 3394 2207
rect 3798 2206 3804 2207
rect 3800 2179 3802 2206
rect 1975 2178 1979 2179
rect 1975 2173 1979 2174
rect 2023 2178 2027 2179
rect 2023 2173 2027 2174
rect 2159 2178 2163 2179
rect 2159 2173 2163 2174
rect 2167 2178 2171 2179
rect 2167 2173 2171 2174
rect 2295 2178 2299 2179
rect 2295 2173 2299 2174
rect 2303 2178 2307 2179
rect 2303 2173 2307 2174
rect 2431 2178 2435 2179
rect 2431 2173 2435 2174
rect 2439 2178 2443 2179
rect 2439 2173 2443 2174
rect 2567 2178 2571 2179
rect 2567 2173 2571 2174
rect 2575 2178 2579 2179
rect 2575 2173 2579 2174
rect 2703 2178 2707 2179
rect 2703 2173 2707 2174
rect 2711 2178 2715 2179
rect 2711 2173 2715 2174
rect 2839 2178 2843 2179
rect 2839 2173 2843 2174
rect 2847 2178 2851 2179
rect 2847 2173 2851 2174
rect 2975 2178 2979 2179
rect 2975 2173 2979 2174
rect 2983 2178 2987 2179
rect 2983 2173 2987 2174
rect 3111 2178 3115 2179
rect 3111 2173 3115 2174
rect 3119 2178 3123 2179
rect 3119 2173 3123 2174
rect 3247 2178 3251 2179
rect 3247 2173 3251 2174
rect 3255 2178 3259 2179
rect 3255 2173 3259 2174
rect 3391 2178 3395 2179
rect 3391 2173 3395 2174
rect 3799 2178 3803 2179
rect 3799 2173 3803 2174
rect 1976 2150 1978 2173
rect 1974 2149 1980 2150
rect 2024 2149 2026 2173
rect 2160 2149 2162 2173
rect 2296 2149 2298 2173
rect 2432 2149 2434 2173
rect 2568 2149 2570 2173
rect 2704 2149 2706 2173
rect 2840 2149 2842 2173
rect 2976 2149 2978 2173
rect 3112 2149 3114 2173
rect 3248 2149 3250 2173
rect 3800 2150 3802 2173
rect 3798 2149 3804 2150
rect 1974 2145 1975 2149
rect 1979 2145 1980 2149
rect 1974 2144 1980 2145
rect 2022 2148 2028 2149
rect 2022 2144 2023 2148
rect 2027 2144 2028 2148
rect 2022 2143 2028 2144
rect 2158 2148 2164 2149
rect 2158 2144 2159 2148
rect 2163 2144 2164 2148
rect 2158 2143 2164 2144
rect 2294 2148 2300 2149
rect 2294 2144 2295 2148
rect 2299 2144 2300 2148
rect 2294 2143 2300 2144
rect 2430 2148 2436 2149
rect 2430 2144 2431 2148
rect 2435 2144 2436 2148
rect 2430 2143 2436 2144
rect 2566 2148 2572 2149
rect 2566 2144 2567 2148
rect 2571 2144 2572 2148
rect 2566 2143 2572 2144
rect 2702 2148 2708 2149
rect 2702 2144 2703 2148
rect 2707 2144 2708 2148
rect 2702 2143 2708 2144
rect 2838 2148 2844 2149
rect 2838 2144 2839 2148
rect 2843 2144 2844 2148
rect 2838 2143 2844 2144
rect 2974 2148 2980 2149
rect 2974 2144 2975 2148
rect 2979 2144 2980 2148
rect 2974 2143 2980 2144
rect 3110 2148 3116 2149
rect 3110 2144 3111 2148
rect 3115 2144 3116 2148
rect 3110 2143 3116 2144
rect 3246 2148 3252 2149
rect 3246 2144 3247 2148
rect 3251 2144 3252 2148
rect 3798 2145 3799 2149
rect 3803 2145 3804 2149
rect 3798 2144 3804 2145
rect 3246 2143 3252 2144
rect 3840 2139 3842 2207
rect 4708 2139 4710 2208
rect 4860 2139 4862 2208
rect 5020 2139 5022 2208
rect 5188 2139 5190 2208
rect 5364 2139 5366 2208
rect 5516 2139 5518 2208
rect 5662 2207 5668 2208
rect 5664 2139 5666 2207
rect 3839 2138 3843 2139
rect 111 2134 115 2135
rect 111 2129 115 2130
rect 131 2134 135 2135
rect 131 2129 135 2130
rect 267 2134 271 2135
rect 267 2129 271 2130
rect 331 2134 335 2135
rect 331 2129 335 2130
rect 411 2134 415 2135
rect 411 2129 415 2130
rect 555 2134 559 2135
rect 555 2129 559 2130
rect 563 2134 567 2135
rect 563 2129 567 2130
rect 715 2134 719 2135
rect 715 2129 719 2130
rect 779 2134 783 2135
rect 779 2129 783 2130
rect 1011 2134 1015 2135
rect 1011 2129 1015 2130
rect 1935 2134 1939 2135
rect 1994 2133 2000 2134
rect 1935 2129 1939 2130
rect 1974 2132 1980 2133
rect 112 2069 114 2129
rect 110 2068 116 2069
rect 132 2068 134 2129
rect 332 2068 334 2129
rect 556 2068 558 2129
rect 780 2068 782 2129
rect 1012 2068 1014 2129
rect 1936 2069 1938 2129
rect 1974 2128 1975 2132
rect 1979 2128 1980 2132
rect 1994 2129 1995 2133
rect 1999 2129 2000 2133
rect 1994 2128 2000 2129
rect 2130 2133 2136 2134
rect 2130 2129 2131 2133
rect 2135 2129 2136 2133
rect 2130 2128 2136 2129
rect 2266 2133 2272 2134
rect 2266 2129 2267 2133
rect 2271 2129 2272 2133
rect 2266 2128 2272 2129
rect 2402 2133 2408 2134
rect 2402 2129 2403 2133
rect 2407 2129 2408 2133
rect 2402 2128 2408 2129
rect 2538 2133 2544 2134
rect 2538 2129 2539 2133
rect 2543 2129 2544 2133
rect 2538 2128 2544 2129
rect 2674 2133 2680 2134
rect 2674 2129 2675 2133
rect 2679 2129 2680 2133
rect 2674 2128 2680 2129
rect 2810 2133 2816 2134
rect 2810 2129 2811 2133
rect 2815 2129 2816 2133
rect 2810 2128 2816 2129
rect 2946 2133 2952 2134
rect 2946 2129 2947 2133
rect 2951 2129 2952 2133
rect 2946 2128 2952 2129
rect 3082 2133 3088 2134
rect 3082 2129 3083 2133
rect 3087 2129 3088 2133
rect 3082 2128 3088 2129
rect 3218 2133 3224 2134
rect 3839 2133 3843 2134
rect 4707 2138 4711 2139
rect 4707 2133 4711 2134
rect 4787 2138 4791 2139
rect 4787 2133 4791 2134
rect 4859 2138 4863 2139
rect 4859 2133 4863 2134
rect 4923 2138 4927 2139
rect 4923 2133 4927 2134
rect 5019 2138 5023 2139
rect 5019 2133 5023 2134
rect 5067 2138 5071 2139
rect 5067 2133 5071 2134
rect 5187 2138 5191 2139
rect 5187 2133 5191 2134
rect 5219 2138 5223 2139
rect 5219 2133 5223 2134
rect 5363 2138 5367 2139
rect 5363 2133 5367 2134
rect 5379 2138 5383 2139
rect 5379 2133 5383 2134
rect 5515 2138 5519 2139
rect 5515 2133 5519 2134
rect 5663 2138 5667 2139
rect 5663 2133 5667 2134
rect 3218 2129 3219 2133
rect 3223 2129 3224 2133
rect 3218 2128 3224 2129
rect 3798 2132 3804 2133
rect 3798 2128 3799 2132
rect 3803 2128 3804 2132
rect 1974 2127 1980 2128
rect 1934 2068 1940 2069
rect 110 2064 111 2068
rect 115 2064 116 2068
rect 110 2063 116 2064
rect 130 2067 136 2068
rect 130 2063 131 2067
rect 135 2063 136 2067
rect 130 2062 136 2063
rect 330 2067 336 2068
rect 330 2063 331 2067
rect 335 2063 336 2067
rect 330 2062 336 2063
rect 554 2067 560 2068
rect 554 2063 555 2067
rect 559 2063 560 2067
rect 554 2062 560 2063
rect 778 2067 784 2068
rect 778 2063 779 2067
rect 783 2063 784 2067
rect 778 2062 784 2063
rect 1010 2067 1016 2068
rect 1010 2063 1011 2067
rect 1015 2063 1016 2067
rect 1934 2064 1935 2068
rect 1939 2064 1940 2068
rect 1934 2063 1940 2064
rect 1010 2062 1016 2063
rect 1976 2059 1978 2127
rect 1996 2059 1998 2128
rect 2132 2059 2134 2128
rect 2268 2059 2270 2128
rect 2404 2059 2406 2128
rect 2540 2059 2542 2128
rect 2676 2059 2678 2128
rect 2812 2059 2814 2128
rect 2948 2059 2950 2128
rect 3084 2059 3086 2128
rect 3220 2059 3222 2128
rect 3798 2127 3804 2128
rect 3800 2059 3802 2127
rect 3840 2073 3842 2133
rect 3838 2072 3844 2073
rect 4788 2072 4790 2133
rect 4924 2072 4926 2133
rect 5068 2072 5070 2133
rect 5220 2072 5222 2133
rect 5380 2072 5382 2133
rect 5516 2072 5518 2133
rect 5664 2073 5666 2133
rect 5662 2072 5668 2073
rect 3838 2068 3839 2072
rect 3843 2068 3844 2072
rect 3838 2067 3844 2068
rect 4786 2071 4792 2072
rect 4786 2067 4787 2071
rect 4791 2067 4792 2071
rect 4786 2066 4792 2067
rect 4922 2071 4928 2072
rect 4922 2067 4923 2071
rect 4927 2067 4928 2071
rect 4922 2066 4928 2067
rect 5066 2071 5072 2072
rect 5066 2067 5067 2071
rect 5071 2067 5072 2071
rect 5066 2066 5072 2067
rect 5218 2071 5224 2072
rect 5218 2067 5219 2071
rect 5223 2067 5224 2071
rect 5218 2066 5224 2067
rect 5378 2071 5384 2072
rect 5378 2067 5379 2071
rect 5383 2067 5384 2071
rect 5378 2066 5384 2067
rect 5514 2071 5520 2072
rect 5514 2067 5515 2071
rect 5519 2067 5520 2071
rect 5662 2068 5663 2072
rect 5667 2068 5668 2072
rect 5662 2067 5668 2068
rect 5514 2066 5520 2067
rect 1975 2058 1979 2059
rect 1975 2053 1979 2054
rect 1995 2058 1999 2059
rect 1995 2053 1999 2054
rect 2131 2058 2135 2059
rect 2131 2053 2135 2054
rect 2267 2058 2271 2059
rect 2267 2053 2271 2054
rect 2403 2058 2407 2059
rect 2403 2053 2407 2054
rect 2539 2058 2543 2059
rect 2539 2053 2543 2054
rect 2675 2058 2679 2059
rect 2675 2053 2679 2054
rect 2811 2058 2815 2059
rect 2811 2053 2815 2054
rect 2947 2058 2951 2059
rect 2947 2053 2951 2054
rect 3083 2058 3087 2059
rect 3083 2053 3087 2054
rect 3091 2058 3095 2059
rect 3091 2053 3095 2054
rect 3219 2058 3223 2059
rect 3219 2053 3223 2054
rect 3243 2058 3247 2059
rect 3243 2053 3247 2054
rect 3395 2058 3399 2059
rect 3395 2053 3399 2054
rect 3799 2058 3803 2059
rect 4814 2056 4820 2057
rect 3799 2053 3803 2054
rect 3838 2055 3844 2056
rect 158 2052 164 2053
rect 110 2051 116 2052
rect 110 2047 111 2051
rect 115 2047 116 2051
rect 158 2048 159 2052
rect 163 2048 164 2052
rect 158 2047 164 2048
rect 358 2052 364 2053
rect 358 2048 359 2052
rect 363 2048 364 2052
rect 358 2047 364 2048
rect 582 2052 588 2053
rect 582 2048 583 2052
rect 587 2048 588 2052
rect 582 2047 588 2048
rect 806 2052 812 2053
rect 806 2048 807 2052
rect 811 2048 812 2052
rect 806 2047 812 2048
rect 1038 2052 1044 2053
rect 1038 2048 1039 2052
rect 1043 2048 1044 2052
rect 1038 2047 1044 2048
rect 1934 2051 1940 2052
rect 1934 2047 1935 2051
rect 1939 2047 1940 2051
rect 110 2046 116 2047
rect 112 2019 114 2046
rect 160 2019 162 2047
rect 360 2019 362 2047
rect 584 2019 586 2047
rect 808 2019 810 2047
rect 1040 2019 1042 2047
rect 1934 2046 1940 2047
rect 1936 2019 1938 2046
rect 111 2018 115 2019
rect 111 2013 115 2014
rect 159 2018 163 2019
rect 159 2013 163 2014
rect 359 2018 363 2019
rect 359 2013 363 2014
rect 463 2018 467 2019
rect 463 2013 467 2014
rect 583 2018 587 2019
rect 583 2013 587 2014
rect 799 2018 803 2019
rect 799 2013 803 2014
rect 807 2018 811 2019
rect 807 2013 811 2014
rect 1039 2018 1043 2019
rect 1039 2013 1043 2014
rect 1143 2018 1147 2019
rect 1143 2013 1147 2014
rect 1487 2018 1491 2019
rect 1487 2013 1491 2014
rect 1815 2018 1819 2019
rect 1815 2013 1819 2014
rect 1935 2018 1939 2019
rect 1935 2013 1939 2014
rect 112 1990 114 2013
rect 110 1989 116 1990
rect 160 1989 162 2013
rect 464 1989 466 2013
rect 800 1989 802 2013
rect 1144 1989 1146 2013
rect 1488 1989 1490 2013
rect 1816 1989 1818 2013
rect 1936 1990 1938 2013
rect 1976 1993 1978 2053
rect 1974 1992 1980 1993
rect 1996 1992 1998 2053
rect 2132 1992 2134 2053
rect 2268 1992 2270 2053
rect 2404 1992 2406 2053
rect 2540 1992 2542 2053
rect 2676 1992 2678 2053
rect 2812 1992 2814 2053
rect 2948 1992 2950 2053
rect 3092 1992 3094 2053
rect 3244 1992 3246 2053
rect 3396 1992 3398 2053
rect 3800 1993 3802 2053
rect 3838 2051 3839 2055
rect 3843 2051 3844 2055
rect 4814 2052 4815 2056
rect 4819 2052 4820 2056
rect 4814 2051 4820 2052
rect 4950 2056 4956 2057
rect 4950 2052 4951 2056
rect 4955 2052 4956 2056
rect 4950 2051 4956 2052
rect 5094 2056 5100 2057
rect 5094 2052 5095 2056
rect 5099 2052 5100 2056
rect 5094 2051 5100 2052
rect 5246 2056 5252 2057
rect 5246 2052 5247 2056
rect 5251 2052 5252 2056
rect 5246 2051 5252 2052
rect 5406 2056 5412 2057
rect 5406 2052 5407 2056
rect 5411 2052 5412 2056
rect 5406 2051 5412 2052
rect 5542 2056 5548 2057
rect 5542 2052 5543 2056
rect 5547 2052 5548 2056
rect 5542 2051 5548 2052
rect 5662 2055 5668 2056
rect 5662 2051 5663 2055
rect 5667 2051 5668 2055
rect 3838 2050 3844 2051
rect 3840 2023 3842 2050
rect 4816 2023 4818 2051
rect 4952 2023 4954 2051
rect 5096 2023 5098 2051
rect 5248 2023 5250 2051
rect 5408 2023 5410 2051
rect 5544 2023 5546 2051
rect 5662 2050 5668 2051
rect 5664 2023 5666 2050
rect 3839 2022 3843 2023
rect 3839 2017 3843 2018
rect 4815 2022 4819 2023
rect 4815 2017 4819 2018
rect 4863 2022 4867 2023
rect 4863 2017 4867 2018
rect 4951 2022 4955 2023
rect 4951 2017 4955 2018
rect 4999 2022 5003 2023
rect 4999 2017 5003 2018
rect 5095 2022 5099 2023
rect 5095 2017 5099 2018
rect 5135 2022 5139 2023
rect 5135 2017 5139 2018
rect 5247 2022 5251 2023
rect 5247 2017 5251 2018
rect 5271 2022 5275 2023
rect 5271 2017 5275 2018
rect 5407 2022 5411 2023
rect 5407 2017 5411 2018
rect 5543 2022 5547 2023
rect 5543 2017 5547 2018
rect 5663 2022 5667 2023
rect 5663 2017 5667 2018
rect 3840 1994 3842 2017
rect 3838 1993 3844 1994
rect 4864 1993 4866 2017
rect 5000 1993 5002 2017
rect 5136 1993 5138 2017
rect 5272 1993 5274 2017
rect 5408 1993 5410 2017
rect 5544 1993 5546 2017
rect 5664 1994 5666 2017
rect 5662 1993 5668 1994
rect 3798 1992 3804 1993
rect 1934 1989 1940 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 110 1984 116 1985
rect 158 1988 164 1989
rect 158 1984 159 1988
rect 163 1984 164 1988
rect 158 1983 164 1984
rect 462 1988 468 1989
rect 462 1984 463 1988
rect 467 1984 468 1988
rect 462 1983 468 1984
rect 798 1988 804 1989
rect 798 1984 799 1988
rect 803 1984 804 1988
rect 798 1983 804 1984
rect 1142 1988 1148 1989
rect 1142 1984 1143 1988
rect 1147 1984 1148 1988
rect 1142 1983 1148 1984
rect 1486 1988 1492 1989
rect 1486 1984 1487 1988
rect 1491 1984 1492 1988
rect 1486 1983 1492 1984
rect 1814 1988 1820 1989
rect 1814 1984 1815 1988
rect 1819 1984 1820 1988
rect 1934 1985 1935 1989
rect 1939 1985 1940 1989
rect 1974 1988 1975 1992
rect 1979 1988 1980 1992
rect 1974 1987 1980 1988
rect 1994 1991 2000 1992
rect 1994 1987 1995 1991
rect 1999 1987 2000 1991
rect 1994 1986 2000 1987
rect 2130 1991 2136 1992
rect 2130 1987 2131 1991
rect 2135 1987 2136 1991
rect 2130 1986 2136 1987
rect 2266 1991 2272 1992
rect 2266 1987 2267 1991
rect 2271 1987 2272 1991
rect 2266 1986 2272 1987
rect 2402 1991 2408 1992
rect 2402 1987 2403 1991
rect 2407 1987 2408 1991
rect 2402 1986 2408 1987
rect 2538 1991 2544 1992
rect 2538 1987 2539 1991
rect 2543 1987 2544 1991
rect 2538 1986 2544 1987
rect 2674 1991 2680 1992
rect 2674 1987 2675 1991
rect 2679 1987 2680 1991
rect 2674 1986 2680 1987
rect 2810 1991 2816 1992
rect 2810 1987 2811 1991
rect 2815 1987 2816 1991
rect 2810 1986 2816 1987
rect 2946 1991 2952 1992
rect 2946 1987 2947 1991
rect 2951 1987 2952 1991
rect 2946 1986 2952 1987
rect 3090 1991 3096 1992
rect 3090 1987 3091 1991
rect 3095 1987 3096 1991
rect 3090 1986 3096 1987
rect 3242 1991 3248 1992
rect 3242 1987 3243 1991
rect 3247 1987 3248 1991
rect 3242 1986 3248 1987
rect 3394 1991 3400 1992
rect 3394 1987 3395 1991
rect 3399 1987 3400 1991
rect 3798 1988 3799 1992
rect 3803 1988 3804 1992
rect 3838 1989 3839 1993
rect 3843 1989 3844 1993
rect 3838 1988 3844 1989
rect 4862 1992 4868 1993
rect 4862 1988 4863 1992
rect 4867 1988 4868 1992
rect 3798 1987 3804 1988
rect 4862 1987 4868 1988
rect 4998 1992 5004 1993
rect 4998 1988 4999 1992
rect 5003 1988 5004 1992
rect 4998 1987 5004 1988
rect 5134 1992 5140 1993
rect 5134 1988 5135 1992
rect 5139 1988 5140 1992
rect 5134 1987 5140 1988
rect 5270 1992 5276 1993
rect 5270 1988 5271 1992
rect 5275 1988 5276 1992
rect 5270 1987 5276 1988
rect 5406 1992 5412 1993
rect 5406 1988 5407 1992
rect 5411 1988 5412 1992
rect 5406 1987 5412 1988
rect 5542 1992 5548 1993
rect 5542 1988 5543 1992
rect 5547 1988 5548 1992
rect 5662 1989 5663 1993
rect 5667 1989 5668 1993
rect 5662 1988 5668 1989
rect 5542 1987 5548 1988
rect 3394 1986 3400 1987
rect 1934 1984 1940 1985
rect 1814 1983 1820 1984
rect 4834 1977 4840 1978
rect 2022 1976 2028 1977
rect 1974 1975 1980 1976
rect 130 1973 136 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 130 1969 131 1973
rect 135 1969 136 1973
rect 130 1968 136 1969
rect 434 1973 440 1974
rect 434 1969 435 1973
rect 439 1969 440 1973
rect 434 1968 440 1969
rect 770 1973 776 1974
rect 770 1969 771 1973
rect 775 1969 776 1973
rect 770 1968 776 1969
rect 1114 1973 1120 1974
rect 1114 1969 1115 1973
rect 1119 1969 1120 1973
rect 1114 1968 1120 1969
rect 1458 1973 1464 1974
rect 1458 1969 1459 1973
rect 1463 1969 1464 1973
rect 1458 1968 1464 1969
rect 1786 1973 1792 1974
rect 1786 1969 1787 1973
rect 1791 1969 1792 1973
rect 1786 1968 1792 1969
rect 1934 1972 1940 1973
rect 1934 1968 1935 1972
rect 1939 1968 1940 1972
rect 1974 1971 1975 1975
rect 1979 1971 1980 1975
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2158 1976 2164 1977
rect 2158 1972 2159 1976
rect 2163 1972 2164 1976
rect 2158 1971 2164 1972
rect 2294 1976 2300 1977
rect 2294 1972 2295 1976
rect 2299 1972 2300 1976
rect 2294 1971 2300 1972
rect 2430 1976 2436 1977
rect 2430 1972 2431 1976
rect 2435 1972 2436 1976
rect 2430 1971 2436 1972
rect 2566 1976 2572 1977
rect 2566 1972 2567 1976
rect 2571 1972 2572 1976
rect 2566 1971 2572 1972
rect 2702 1976 2708 1977
rect 2702 1972 2703 1976
rect 2707 1972 2708 1976
rect 2702 1971 2708 1972
rect 2838 1976 2844 1977
rect 2838 1972 2839 1976
rect 2843 1972 2844 1976
rect 2838 1971 2844 1972
rect 2974 1976 2980 1977
rect 2974 1972 2975 1976
rect 2979 1972 2980 1976
rect 2974 1971 2980 1972
rect 3118 1976 3124 1977
rect 3118 1972 3119 1976
rect 3123 1972 3124 1976
rect 3118 1971 3124 1972
rect 3270 1976 3276 1977
rect 3270 1972 3271 1976
rect 3275 1972 3276 1976
rect 3270 1971 3276 1972
rect 3422 1976 3428 1977
rect 3838 1976 3844 1977
rect 3422 1972 3423 1976
rect 3427 1972 3428 1976
rect 3422 1971 3428 1972
rect 3798 1975 3804 1976
rect 3798 1971 3799 1975
rect 3803 1971 3804 1975
rect 3838 1972 3839 1976
rect 3843 1972 3844 1976
rect 4834 1973 4835 1977
rect 4839 1973 4840 1977
rect 4834 1972 4840 1973
rect 4970 1977 4976 1978
rect 4970 1973 4971 1977
rect 4975 1973 4976 1977
rect 4970 1972 4976 1973
rect 5106 1977 5112 1978
rect 5106 1973 5107 1977
rect 5111 1973 5112 1977
rect 5106 1972 5112 1973
rect 5242 1977 5248 1978
rect 5242 1973 5243 1977
rect 5247 1973 5248 1977
rect 5242 1972 5248 1973
rect 5378 1977 5384 1978
rect 5378 1973 5379 1977
rect 5383 1973 5384 1977
rect 5378 1972 5384 1973
rect 5514 1977 5520 1978
rect 5514 1973 5515 1977
rect 5519 1973 5520 1977
rect 5514 1972 5520 1973
rect 5662 1976 5668 1977
rect 5662 1972 5663 1976
rect 5667 1972 5668 1976
rect 3838 1971 3844 1972
rect 1974 1970 1980 1971
rect 110 1967 116 1968
rect 112 1907 114 1967
rect 132 1907 134 1968
rect 436 1907 438 1968
rect 772 1907 774 1968
rect 1116 1907 1118 1968
rect 1460 1907 1462 1968
rect 1788 1907 1790 1968
rect 1934 1967 1940 1968
rect 1936 1907 1938 1967
rect 1976 1939 1978 1970
rect 2024 1939 2026 1971
rect 2160 1939 2162 1971
rect 2296 1939 2298 1971
rect 2432 1939 2434 1971
rect 2568 1939 2570 1971
rect 2704 1939 2706 1971
rect 2840 1939 2842 1971
rect 2976 1939 2978 1971
rect 3120 1939 3122 1971
rect 3272 1939 3274 1971
rect 3424 1939 3426 1971
rect 3798 1970 3804 1971
rect 3800 1939 3802 1970
rect 1975 1938 1979 1939
rect 1975 1933 1979 1934
rect 2023 1938 2027 1939
rect 2023 1933 2027 1934
rect 2159 1938 2163 1939
rect 2159 1933 2163 1934
rect 2295 1938 2299 1939
rect 2295 1933 2299 1934
rect 2431 1938 2435 1939
rect 2431 1933 2435 1934
rect 2527 1938 2531 1939
rect 2527 1933 2531 1934
rect 2567 1938 2571 1939
rect 2567 1933 2571 1934
rect 2663 1938 2667 1939
rect 2663 1933 2667 1934
rect 2703 1938 2707 1939
rect 2703 1933 2707 1934
rect 2799 1938 2803 1939
rect 2799 1933 2803 1934
rect 2839 1938 2843 1939
rect 2839 1933 2843 1934
rect 2935 1938 2939 1939
rect 2935 1933 2939 1934
rect 2975 1938 2979 1939
rect 2975 1933 2979 1934
rect 3071 1938 3075 1939
rect 3071 1933 3075 1934
rect 3119 1938 3123 1939
rect 3119 1933 3123 1934
rect 3207 1938 3211 1939
rect 3207 1933 3211 1934
rect 3271 1938 3275 1939
rect 3271 1933 3275 1934
rect 3351 1938 3355 1939
rect 3351 1933 3355 1934
rect 3423 1938 3427 1939
rect 3423 1933 3427 1934
rect 3799 1938 3803 1939
rect 3799 1933 3803 1934
rect 1976 1910 1978 1933
rect 1974 1909 1980 1910
rect 2528 1909 2530 1933
rect 2664 1909 2666 1933
rect 2800 1909 2802 1933
rect 2936 1909 2938 1933
rect 3072 1909 3074 1933
rect 3208 1909 3210 1933
rect 3352 1909 3354 1933
rect 3800 1910 3802 1933
rect 3798 1909 3804 1910
rect 111 1906 115 1907
rect 111 1901 115 1902
rect 131 1906 135 1907
rect 131 1901 135 1902
rect 195 1906 199 1907
rect 195 1901 199 1902
rect 435 1906 439 1907
rect 435 1901 439 1902
rect 451 1906 455 1907
rect 451 1901 455 1902
rect 699 1906 703 1907
rect 699 1901 703 1902
rect 771 1906 775 1907
rect 771 1901 775 1902
rect 931 1906 935 1907
rect 931 1901 935 1902
rect 1115 1906 1119 1907
rect 1115 1901 1119 1902
rect 1155 1906 1159 1907
rect 1155 1901 1159 1902
rect 1371 1906 1375 1907
rect 1371 1901 1375 1902
rect 1459 1906 1463 1907
rect 1459 1901 1463 1902
rect 1587 1906 1591 1907
rect 1587 1901 1591 1902
rect 1787 1906 1791 1907
rect 1787 1901 1791 1902
rect 1935 1906 1939 1907
rect 1974 1905 1975 1909
rect 1979 1905 1980 1909
rect 1974 1904 1980 1905
rect 2526 1908 2532 1909
rect 2526 1904 2527 1908
rect 2531 1904 2532 1908
rect 2526 1903 2532 1904
rect 2662 1908 2668 1909
rect 2662 1904 2663 1908
rect 2667 1904 2668 1908
rect 2662 1903 2668 1904
rect 2798 1908 2804 1909
rect 2798 1904 2799 1908
rect 2803 1904 2804 1908
rect 2798 1903 2804 1904
rect 2934 1908 2940 1909
rect 2934 1904 2935 1908
rect 2939 1904 2940 1908
rect 2934 1903 2940 1904
rect 3070 1908 3076 1909
rect 3070 1904 3071 1908
rect 3075 1904 3076 1908
rect 3070 1903 3076 1904
rect 3206 1908 3212 1909
rect 3206 1904 3207 1908
rect 3211 1904 3212 1908
rect 3206 1903 3212 1904
rect 3350 1908 3356 1909
rect 3350 1904 3351 1908
rect 3355 1904 3356 1908
rect 3798 1905 3799 1909
rect 3803 1905 3804 1909
rect 3840 1907 3842 1971
rect 4836 1907 4838 1972
rect 4972 1907 4974 1972
rect 5108 1907 5110 1972
rect 5244 1907 5246 1972
rect 5380 1907 5382 1972
rect 5516 1907 5518 1972
rect 5662 1971 5668 1972
rect 5664 1907 5666 1971
rect 3798 1904 3804 1905
rect 3839 1906 3843 1907
rect 3350 1903 3356 1904
rect 1935 1901 1939 1902
rect 3839 1901 3843 1902
rect 4683 1906 4687 1907
rect 4683 1901 4687 1902
rect 4835 1906 4839 1907
rect 4835 1901 4839 1902
rect 4843 1906 4847 1907
rect 4843 1901 4847 1902
rect 4971 1906 4975 1907
rect 4971 1901 4975 1902
rect 5011 1906 5015 1907
rect 5011 1901 5015 1902
rect 5107 1906 5111 1907
rect 5107 1901 5111 1902
rect 5179 1906 5183 1907
rect 5179 1901 5183 1902
rect 5243 1906 5247 1907
rect 5243 1901 5247 1902
rect 5355 1906 5359 1907
rect 5355 1901 5359 1902
rect 5379 1906 5383 1907
rect 5379 1901 5383 1902
rect 5515 1906 5519 1907
rect 5515 1901 5519 1902
rect 5663 1906 5667 1907
rect 5663 1901 5667 1902
rect 112 1841 114 1901
rect 110 1840 116 1841
rect 196 1840 198 1901
rect 452 1840 454 1901
rect 700 1840 702 1901
rect 932 1840 934 1901
rect 1156 1840 1158 1901
rect 1372 1840 1374 1901
rect 1588 1840 1590 1901
rect 1788 1840 1790 1901
rect 1936 1841 1938 1901
rect 2498 1893 2504 1894
rect 1974 1892 1980 1893
rect 1974 1888 1975 1892
rect 1979 1888 1980 1892
rect 2498 1889 2499 1893
rect 2503 1889 2504 1893
rect 2498 1888 2504 1889
rect 2634 1893 2640 1894
rect 2634 1889 2635 1893
rect 2639 1889 2640 1893
rect 2634 1888 2640 1889
rect 2770 1893 2776 1894
rect 2770 1889 2771 1893
rect 2775 1889 2776 1893
rect 2770 1888 2776 1889
rect 2906 1893 2912 1894
rect 2906 1889 2907 1893
rect 2911 1889 2912 1893
rect 2906 1888 2912 1889
rect 3042 1893 3048 1894
rect 3042 1889 3043 1893
rect 3047 1889 3048 1893
rect 3042 1888 3048 1889
rect 3178 1893 3184 1894
rect 3178 1889 3179 1893
rect 3183 1889 3184 1893
rect 3178 1888 3184 1889
rect 3322 1893 3328 1894
rect 3322 1889 3323 1893
rect 3327 1889 3328 1893
rect 3322 1888 3328 1889
rect 3798 1892 3804 1893
rect 3798 1888 3799 1892
rect 3803 1888 3804 1892
rect 1974 1887 1980 1888
rect 1934 1840 1940 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 110 1835 116 1836
rect 194 1839 200 1840
rect 194 1835 195 1839
rect 199 1835 200 1839
rect 194 1834 200 1835
rect 450 1839 456 1840
rect 450 1835 451 1839
rect 455 1835 456 1839
rect 450 1834 456 1835
rect 698 1839 704 1840
rect 698 1835 699 1839
rect 703 1835 704 1839
rect 698 1834 704 1835
rect 930 1839 936 1840
rect 930 1835 931 1839
rect 935 1835 936 1839
rect 930 1834 936 1835
rect 1154 1839 1160 1840
rect 1154 1835 1155 1839
rect 1159 1835 1160 1839
rect 1154 1834 1160 1835
rect 1370 1839 1376 1840
rect 1370 1835 1371 1839
rect 1375 1835 1376 1839
rect 1370 1834 1376 1835
rect 1586 1839 1592 1840
rect 1586 1835 1587 1839
rect 1591 1835 1592 1839
rect 1586 1834 1592 1835
rect 1786 1839 1792 1840
rect 1786 1835 1787 1839
rect 1791 1835 1792 1839
rect 1934 1836 1935 1840
rect 1939 1836 1940 1840
rect 1934 1835 1940 1836
rect 1786 1834 1792 1835
rect 1976 1827 1978 1887
rect 2500 1827 2502 1888
rect 2636 1827 2638 1888
rect 2772 1827 2774 1888
rect 2908 1827 2910 1888
rect 3044 1827 3046 1888
rect 3180 1827 3182 1888
rect 3324 1827 3326 1888
rect 3798 1887 3804 1888
rect 3800 1827 3802 1887
rect 3840 1841 3842 1901
rect 3838 1840 3844 1841
rect 4684 1840 4686 1901
rect 4844 1840 4846 1901
rect 5012 1840 5014 1901
rect 5180 1840 5182 1901
rect 5356 1840 5358 1901
rect 5516 1840 5518 1901
rect 5664 1841 5666 1901
rect 5662 1840 5668 1841
rect 3838 1836 3839 1840
rect 3843 1836 3844 1840
rect 3838 1835 3844 1836
rect 4682 1839 4688 1840
rect 4682 1835 4683 1839
rect 4687 1835 4688 1839
rect 4682 1834 4688 1835
rect 4842 1839 4848 1840
rect 4842 1835 4843 1839
rect 4847 1835 4848 1839
rect 4842 1834 4848 1835
rect 5010 1839 5016 1840
rect 5010 1835 5011 1839
rect 5015 1835 5016 1839
rect 5010 1834 5016 1835
rect 5178 1839 5184 1840
rect 5178 1835 5179 1839
rect 5183 1835 5184 1839
rect 5178 1834 5184 1835
rect 5354 1839 5360 1840
rect 5354 1835 5355 1839
rect 5359 1835 5360 1839
rect 5354 1834 5360 1835
rect 5514 1839 5520 1840
rect 5514 1835 5515 1839
rect 5519 1835 5520 1839
rect 5662 1836 5663 1840
rect 5667 1836 5668 1840
rect 5662 1835 5668 1836
rect 5514 1834 5520 1835
rect 1975 1826 1979 1827
rect 222 1824 228 1825
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 222 1820 223 1824
rect 227 1820 228 1824
rect 222 1819 228 1820
rect 478 1824 484 1825
rect 478 1820 479 1824
rect 483 1820 484 1824
rect 478 1819 484 1820
rect 726 1824 732 1825
rect 726 1820 727 1824
rect 731 1820 732 1824
rect 726 1819 732 1820
rect 958 1824 964 1825
rect 958 1820 959 1824
rect 963 1820 964 1824
rect 958 1819 964 1820
rect 1182 1824 1188 1825
rect 1182 1820 1183 1824
rect 1187 1820 1188 1824
rect 1182 1819 1188 1820
rect 1398 1824 1404 1825
rect 1398 1820 1399 1824
rect 1403 1820 1404 1824
rect 1398 1819 1404 1820
rect 1614 1824 1620 1825
rect 1614 1820 1615 1824
rect 1619 1820 1620 1824
rect 1614 1819 1620 1820
rect 1814 1824 1820 1825
rect 1814 1820 1815 1824
rect 1819 1820 1820 1824
rect 1814 1819 1820 1820
rect 1934 1823 1940 1824
rect 1934 1819 1935 1823
rect 1939 1819 1940 1823
rect 1975 1821 1979 1822
rect 2443 1826 2447 1827
rect 2443 1821 2447 1822
rect 2499 1826 2503 1827
rect 2499 1821 2503 1822
rect 2587 1826 2591 1827
rect 2587 1821 2591 1822
rect 2635 1826 2639 1827
rect 2635 1821 2639 1822
rect 2739 1826 2743 1827
rect 2739 1821 2743 1822
rect 2771 1826 2775 1827
rect 2771 1821 2775 1822
rect 2891 1826 2895 1827
rect 2891 1821 2895 1822
rect 2907 1826 2911 1827
rect 2907 1821 2911 1822
rect 3043 1826 3047 1827
rect 3043 1821 3047 1822
rect 3179 1826 3183 1827
rect 3179 1821 3183 1822
rect 3195 1826 3199 1827
rect 3195 1821 3199 1822
rect 3323 1826 3327 1827
rect 3323 1821 3327 1822
rect 3799 1826 3803 1827
rect 4710 1824 4716 1825
rect 3799 1821 3803 1822
rect 3838 1823 3844 1824
rect 110 1818 116 1819
rect 112 1791 114 1818
rect 224 1791 226 1819
rect 480 1791 482 1819
rect 728 1791 730 1819
rect 960 1791 962 1819
rect 1184 1791 1186 1819
rect 1400 1791 1402 1819
rect 1616 1791 1618 1819
rect 1816 1791 1818 1819
rect 1934 1818 1940 1819
rect 1936 1791 1938 1818
rect 111 1790 115 1791
rect 111 1785 115 1786
rect 223 1790 227 1791
rect 223 1785 227 1786
rect 231 1790 235 1791
rect 231 1785 235 1786
rect 447 1790 451 1791
rect 447 1785 451 1786
rect 479 1790 483 1791
rect 479 1785 483 1786
rect 671 1790 675 1791
rect 671 1785 675 1786
rect 727 1790 731 1791
rect 727 1785 731 1786
rect 895 1790 899 1791
rect 895 1785 899 1786
rect 959 1790 963 1791
rect 959 1785 963 1786
rect 1119 1790 1123 1791
rect 1119 1785 1123 1786
rect 1183 1790 1187 1791
rect 1183 1785 1187 1786
rect 1343 1790 1347 1791
rect 1343 1785 1347 1786
rect 1399 1790 1403 1791
rect 1399 1785 1403 1786
rect 1567 1790 1571 1791
rect 1567 1785 1571 1786
rect 1615 1790 1619 1791
rect 1615 1785 1619 1786
rect 1799 1790 1803 1791
rect 1799 1785 1803 1786
rect 1815 1790 1819 1791
rect 1815 1785 1819 1786
rect 1935 1790 1939 1791
rect 1935 1785 1939 1786
rect 112 1762 114 1785
rect 110 1761 116 1762
rect 232 1761 234 1785
rect 448 1761 450 1785
rect 672 1761 674 1785
rect 896 1761 898 1785
rect 1120 1761 1122 1785
rect 1344 1761 1346 1785
rect 1568 1761 1570 1785
rect 1800 1761 1802 1785
rect 1936 1762 1938 1785
rect 1934 1761 1940 1762
rect 1976 1761 1978 1821
rect 110 1757 111 1761
rect 115 1757 116 1761
rect 110 1756 116 1757
rect 230 1760 236 1761
rect 230 1756 231 1760
rect 235 1756 236 1760
rect 230 1755 236 1756
rect 446 1760 452 1761
rect 446 1756 447 1760
rect 451 1756 452 1760
rect 446 1755 452 1756
rect 670 1760 676 1761
rect 670 1756 671 1760
rect 675 1756 676 1760
rect 670 1755 676 1756
rect 894 1760 900 1761
rect 894 1756 895 1760
rect 899 1756 900 1760
rect 894 1755 900 1756
rect 1118 1760 1124 1761
rect 1118 1756 1119 1760
rect 1123 1756 1124 1760
rect 1118 1755 1124 1756
rect 1342 1760 1348 1761
rect 1342 1756 1343 1760
rect 1347 1756 1348 1760
rect 1342 1755 1348 1756
rect 1566 1760 1572 1761
rect 1566 1756 1567 1760
rect 1571 1756 1572 1760
rect 1566 1755 1572 1756
rect 1798 1760 1804 1761
rect 1798 1756 1799 1760
rect 1803 1756 1804 1760
rect 1934 1757 1935 1761
rect 1939 1757 1940 1761
rect 1934 1756 1940 1757
rect 1974 1760 1980 1761
rect 2444 1760 2446 1821
rect 2588 1760 2590 1821
rect 2740 1760 2742 1821
rect 2892 1760 2894 1821
rect 3044 1760 3046 1821
rect 3196 1760 3198 1821
rect 3800 1761 3802 1821
rect 3838 1819 3839 1823
rect 3843 1819 3844 1823
rect 4710 1820 4711 1824
rect 4715 1820 4716 1824
rect 4710 1819 4716 1820
rect 4870 1824 4876 1825
rect 4870 1820 4871 1824
rect 4875 1820 4876 1824
rect 4870 1819 4876 1820
rect 5038 1824 5044 1825
rect 5038 1820 5039 1824
rect 5043 1820 5044 1824
rect 5038 1819 5044 1820
rect 5206 1824 5212 1825
rect 5206 1820 5207 1824
rect 5211 1820 5212 1824
rect 5206 1819 5212 1820
rect 5382 1824 5388 1825
rect 5382 1820 5383 1824
rect 5387 1820 5388 1824
rect 5382 1819 5388 1820
rect 5542 1824 5548 1825
rect 5542 1820 5543 1824
rect 5547 1820 5548 1824
rect 5542 1819 5548 1820
rect 5662 1823 5668 1824
rect 5662 1819 5663 1823
rect 5667 1819 5668 1823
rect 3838 1818 3844 1819
rect 3840 1791 3842 1818
rect 4712 1791 4714 1819
rect 4872 1791 4874 1819
rect 5040 1791 5042 1819
rect 5208 1791 5210 1819
rect 5384 1791 5386 1819
rect 5544 1791 5546 1819
rect 5662 1818 5668 1819
rect 5664 1791 5666 1818
rect 3839 1790 3843 1791
rect 3839 1785 3843 1786
rect 3887 1790 3891 1791
rect 3887 1785 3891 1786
rect 4023 1790 4027 1791
rect 4023 1785 4027 1786
rect 4191 1790 4195 1791
rect 4191 1785 4195 1786
rect 4367 1790 4371 1791
rect 4367 1785 4371 1786
rect 4559 1790 4563 1791
rect 4559 1785 4563 1786
rect 4711 1790 4715 1791
rect 4711 1785 4715 1786
rect 4767 1790 4771 1791
rect 4767 1785 4771 1786
rect 4871 1790 4875 1791
rect 4871 1785 4875 1786
rect 4983 1790 4987 1791
rect 4983 1785 4987 1786
rect 5039 1790 5043 1791
rect 5039 1785 5043 1786
rect 5207 1790 5211 1791
rect 5207 1785 5211 1786
rect 5215 1790 5219 1791
rect 5215 1785 5219 1786
rect 5383 1790 5387 1791
rect 5383 1785 5387 1786
rect 5447 1790 5451 1791
rect 5447 1785 5451 1786
rect 5543 1790 5547 1791
rect 5543 1785 5547 1786
rect 5663 1790 5667 1791
rect 5663 1785 5667 1786
rect 3840 1762 3842 1785
rect 3838 1761 3844 1762
rect 3888 1761 3890 1785
rect 4024 1761 4026 1785
rect 4192 1761 4194 1785
rect 4368 1761 4370 1785
rect 4560 1761 4562 1785
rect 4768 1761 4770 1785
rect 4984 1761 4986 1785
rect 5216 1761 5218 1785
rect 5448 1761 5450 1785
rect 5664 1762 5666 1785
rect 5662 1761 5668 1762
rect 3798 1760 3804 1761
rect 1974 1756 1975 1760
rect 1979 1756 1980 1760
rect 1798 1755 1804 1756
rect 1974 1755 1980 1756
rect 2442 1759 2448 1760
rect 2442 1755 2443 1759
rect 2447 1755 2448 1759
rect 2442 1754 2448 1755
rect 2586 1759 2592 1760
rect 2586 1755 2587 1759
rect 2591 1755 2592 1759
rect 2586 1754 2592 1755
rect 2738 1759 2744 1760
rect 2738 1755 2739 1759
rect 2743 1755 2744 1759
rect 2738 1754 2744 1755
rect 2890 1759 2896 1760
rect 2890 1755 2891 1759
rect 2895 1755 2896 1759
rect 2890 1754 2896 1755
rect 3042 1759 3048 1760
rect 3042 1755 3043 1759
rect 3047 1755 3048 1759
rect 3042 1754 3048 1755
rect 3194 1759 3200 1760
rect 3194 1755 3195 1759
rect 3199 1755 3200 1759
rect 3798 1756 3799 1760
rect 3803 1756 3804 1760
rect 3838 1757 3839 1761
rect 3843 1757 3844 1761
rect 3838 1756 3844 1757
rect 3886 1760 3892 1761
rect 3886 1756 3887 1760
rect 3891 1756 3892 1760
rect 3798 1755 3804 1756
rect 3886 1755 3892 1756
rect 4022 1760 4028 1761
rect 4022 1756 4023 1760
rect 4027 1756 4028 1760
rect 4022 1755 4028 1756
rect 4190 1760 4196 1761
rect 4190 1756 4191 1760
rect 4195 1756 4196 1760
rect 4190 1755 4196 1756
rect 4366 1760 4372 1761
rect 4366 1756 4367 1760
rect 4371 1756 4372 1760
rect 4366 1755 4372 1756
rect 4558 1760 4564 1761
rect 4558 1756 4559 1760
rect 4563 1756 4564 1760
rect 4558 1755 4564 1756
rect 4766 1760 4772 1761
rect 4766 1756 4767 1760
rect 4771 1756 4772 1760
rect 4766 1755 4772 1756
rect 4982 1760 4988 1761
rect 4982 1756 4983 1760
rect 4987 1756 4988 1760
rect 4982 1755 4988 1756
rect 5214 1760 5220 1761
rect 5214 1756 5215 1760
rect 5219 1756 5220 1760
rect 5214 1755 5220 1756
rect 5446 1760 5452 1761
rect 5446 1756 5447 1760
rect 5451 1756 5452 1760
rect 5662 1757 5663 1761
rect 5667 1757 5668 1761
rect 5662 1756 5668 1757
rect 5446 1755 5452 1756
rect 3194 1754 3200 1755
rect 202 1745 208 1746
rect 110 1744 116 1745
rect 110 1740 111 1744
rect 115 1740 116 1744
rect 202 1741 203 1745
rect 207 1741 208 1745
rect 202 1740 208 1741
rect 418 1745 424 1746
rect 418 1741 419 1745
rect 423 1741 424 1745
rect 418 1740 424 1741
rect 642 1745 648 1746
rect 642 1741 643 1745
rect 647 1741 648 1745
rect 642 1740 648 1741
rect 866 1745 872 1746
rect 866 1741 867 1745
rect 871 1741 872 1745
rect 866 1740 872 1741
rect 1090 1745 1096 1746
rect 1090 1741 1091 1745
rect 1095 1741 1096 1745
rect 1090 1740 1096 1741
rect 1314 1745 1320 1746
rect 1314 1741 1315 1745
rect 1319 1741 1320 1745
rect 1314 1740 1320 1741
rect 1538 1745 1544 1746
rect 1538 1741 1539 1745
rect 1543 1741 1544 1745
rect 1538 1740 1544 1741
rect 1770 1745 1776 1746
rect 3858 1745 3864 1746
rect 1770 1741 1771 1745
rect 1775 1741 1776 1745
rect 1770 1740 1776 1741
rect 1934 1744 1940 1745
rect 2470 1744 2476 1745
rect 1934 1740 1935 1744
rect 1939 1740 1940 1744
rect 110 1739 116 1740
rect 112 1679 114 1739
rect 204 1679 206 1740
rect 420 1679 422 1740
rect 644 1679 646 1740
rect 868 1679 870 1740
rect 1092 1679 1094 1740
rect 1316 1679 1318 1740
rect 1540 1679 1542 1740
rect 1772 1679 1774 1740
rect 1934 1739 1940 1740
rect 1974 1743 1980 1744
rect 1974 1739 1975 1743
rect 1979 1739 1980 1743
rect 2470 1740 2471 1744
rect 2475 1740 2476 1744
rect 2470 1739 2476 1740
rect 2614 1744 2620 1745
rect 2614 1740 2615 1744
rect 2619 1740 2620 1744
rect 2614 1739 2620 1740
rect 2766 1744 2772 1745
rect 2766 1740 2767 1744
rect 2771 1740 2772 1744
rect 2766 1739 2772 1740
rect 2918 1744 2924 1745
rect 2918 1740 2919 1744
rect 2923 1740 2924 1744
rect 2918 1739 2924 1740
rect 3070 1744 3076 1745
rect 3070 1740 3071 1744
rect 3075 1740 3076 1744
rect 3070 1739 3076 1740
rect 3222 1744 3228 1745
rect 3838 1744 3844 1745
rect 3222 1740 3223 1744
rect 3227 1740 3228 1744
rect 3222 1739 3228 1740
rect 3798 1743 3804 1744
rect 3798 1739 3799 1743
rect 3803 1739 3804 1743
rect 3838 1740 3839 1744
rect 3843 1740 3844 1744
rect 3858 1741 3859 1745
rect 3863 1741 3864 1745
rect 3858 1740 3864 1741
rect 3994 1745 4000 1746
rect 3994 1741 3995 1745
rect 3999 1741 4000 1745
rect 3994 1740 4000 1741
rect 4162 1745 4168 1746
rect 4162 1741 4163 1745
rect 4167 1741 4168 1745
rect 4162 1740 4168 1741
rect 4338 1745 4344 1746
rect 4338 1741 4339 1745
rect 4343 1741 4344 1745
rect 4338 1740 4344 1741
rect 4530 1745 4536 1746
rect 4530 1741 4531 1745
rect 4535 1741 4536 1745
rect 4530 1740 4536 1741
rect 4738 1745 4744 1746
rect 4738 1741 4739 1745
rect 4743 1741 4744 1745
rect 4738 1740 4744 1741
rect 4954 1745 4960 1746
rect 4954 1741 4955 1745
rect 4959 1741 4960 1745
rect 4954 1740 4960 1741
rect 5186 1745 5192 1746
rect 5186 1741 5187 1745
rect 5191 1741 5192 1745
rect 5186 1740 5192 1741
rect 5418 1745 5424 1746
rect 5418 1741 5419 1745
rect 5423 1741 5424 1745
rect 5418 1740 5424 1741
rect 5662 1744 5668 1745
rect 5662 1740 5663 1744
rect 5667 1740 5668 1744
rect 3838 1739 3844 1740
rect 1936 1679 1938 1739
rect 1974 1738 1980 1739
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 203 1678 207 1679
rect 203 1673 207 1674
rect 275 1678 279 1679
rect 275 1673 279 1674
rect 419 1678 423 1679
rect 419 1673 423 1674
rect 459 1678 463 1679
rect 459 1673 463 1674
rect 643 1678 647 1679
rect 643 1673 647 1674
rect 667 1678 671 1679
rect 667 1673 671 1674
rect 867 1678 871 1679
rect 867 1673 871 1674
rect 883 1678 887 1679
rect 883 1673 887 1674
rect 1091 1678 1095 1679
rect 1091 1673 1095 1674
rect 1115 1678 1119 1679
rect 1115 1673 1119 1674
rect 1315 1678 1319 1679
rect 1315 1673 1319 1674
rect 1355 1678 1359 1679
rect 1355 1673 1359 1674
rect 1539 1678 1543 1679
rect 1539 1673 1543 1674
rect 1595 1678 1599 1679
rect 1595 1673 1599 1674
rect 1771 1678 1775 1679
rect 1771 1673 1775 1674
rect 1935 1678 1939 1679
rect 1935 1673 1939 1674
rect 112 1613 114 1673
rect 110 1612 116 1613
rect 276 1612 278 1673
rect 460 1612 462 1673
rect 668 1612 670 1673
rect 884 1612 886 1673
rect 1116 1612 1118 1673
rect 1356 1612 1358 1673
rect 1596 1612 1598 1673
rect 1936 1613 1938 1673
rect 1976 1671 1978 1738
rect 2472 1671 2474 1739
rect 2616 1671 2618 1739
rect 2768 1671 2770 1739
rect 2920 1671 2922 1739
rect 3072 1671 3074 1739
rect 3224 1671 3226 1739
rect 3798 1738 3804 1739
rect 3800 1671 3802 1738
rect 3840 1679 3842 1739
rect 3860 1679 3862 1740
rect 3996 1679 3998 1740
rect 4164 1679 4166 1740
rect 4340 1679 4342 1740
rect 4532 1679 4534 1740
rect 4740 1679 4742 1740
rect 4956 1679 4958 1740
rect 5188 1679 5190 1740
rect 5420 1679 5422 1740
rect 5662 1739 5668 1740
rect 5664 1679 5666 1739
rect 3839 1678 3843 1679
rect 3839 1673 3843 1674
rect 3859 1678 3863 1679
rect 3859 1673 3863 1674
rect 3995 1678 3999 1679
rect 3995 1673 3999 1674
rect 4131 1678 4135 1679
rect 4131 1673 4135 1674
rect 4163 1678 4167 1679
rect 4163 1673 4167 1674
rect 4283 1678 4287 1679
rect 4283 1673 4287 1674
rect 4339 1678 4343 1679
rect 4339 1673 4343 1674
rect 4483 1678 4487 1679
rect 4483 1673 4487 1674
rect 4531 1678 4535 1679
rect 4531 1673 4535 1674
rect 4715 1678 4719 1679
rect 4715 1673 4719 1674
rect 4739 1678 4743 1679
rect 4739 1673 4743 1674
rect 4955 1678 4959 1679
rect 4955 1673 4959 1674
rect 4979 1678 4983 1679
rect 4979 1673 4983 1674
rect 5187 1678 5191 1679
rect 5187 1673 5191 1674
rect 5259 1678 5263 1679
rect 5259 1673 5263 1674
rect 5419 1678 5423 1679
rect 5419 1673 5423 1674
rect 5515 1678 5519 1679
rect 5515 1673 5519 1674
rect 5663 1678 5667 1679
rect 5663 1673 5667 1674
rect 1975 1670 1979 1671
rect 1975 1665 1979 1666
rect 2231 1670 2235 1671
rect 2231 1665 2235 1666
rect 2471 1670 2475 1671
rect 2471 1665 2475 1666
rect 2599 1670 2603 1671
rect 2599 1665 2603 1666
rect 2615 1670 2619 1671
rect 2615 1665 2619 1666
rect 2767 1670 2771 1671
rect 2767 1665 2771 1666
rect 2919 1670 2923 1671
rect 2919 1665 2923 1666
rect 2967 1670 2971 1671
rect 2967 1665 2971 1666
rect 3071 1670 3075 1671
rect 3071 1665 3075 1666
rect 3223 1670 3227 1671
rect 3223 1665 3227 1666
rect 3335 1670 3339 1671
rect 3335 1665 3339 1666
rect 3679 1670 3683 1671
rect 3679 1665 3683 1666
rect 3799 1670 3803 1671
rect 3799 1665 3803 1666
rect 1976 1642 1978 1665
rect 1974 1641 1980 1642
rect 2232 1641 2234 1665
rect 2600 1641 2602 1665
rect 2968 1641 2970 1665
rect 3336 1641 3338 1665
rect 3680 1641 3682 1665
rect 3800 1642 3802 1665
rect 3798 1641 3804 1642
rect 1974 1637 1975 1641
rect 1979 1637 1980 1641
rect 1974 1636 1980 1637
rect 2230 1640 2236 1641
rect 2230 1636 2231 1640
rect 2235 1636 2236 1640
rect 2230 1635 2236 1636
rect 2598 1640 2604 1641
rect 2598 1636 2599 1640
rect 2603 1636 2604 1640
rect 2598 1635 2604 1636
rect 2966 1640 2972 1641
rect 2966 1636 2967 1640
rect 2971 1636 2972 1640
rect 2966 1635 2972 1636
rect 3334 1640 3340 1641
rect 3334 1636 3335 1640
rect 3339 1636 3340 1640
rect 3334 1635 3340 1636
rect 3678 1640 3684 1641
rect 3678 1636 3679 1640
rect 3683 1636 3684 1640
rect 3798 1637 3799 1641
rect 3803 1637 3804 1641
rect 3798 1636 3804 1637
rect 3678 1635 3684 1636
rect 2202 1625 2208 1626
rect 1974 1624 1980 1625
rect 1974 1620 1975 1624
rect 1979 1620 1980 1624
rect 2202 1621 2203 1625
rect 2207 1621 2208 1625
rect 2202 1620 2208 1621
rect 2570 1625 2576 1626
rect 2570 1621 2571 1625
rect 2575 1621 2576 1625
rect 2570 1620 2576 1621
rect 2938 1625 2944 1626
rect 2938 1621 2939 1625
rect 2943 1621 2944 1625
rect 2938 1620 2944 1621
rect 3306 1625 3312 1626
rect 3306 1621 3307 1625
rect 3311 1621 3312 1625
rect 3306 1620 3312 1621
rect 3650 1625 3656 1626
rect 3650 1621 3651 1625
rect 3655 1621 3656 1625
rect 3650 1620 3656 1621
rect 3798 1624 3804 1625
rect 3798 1620 3799 1624
rect 3803 1620 3804 1624
rect 1974 1619 1980 1620
rect 1934 1612 1940 1613
rect 110 1608 111 1612
rect 115 1608 116 1612
rect 110 1607 116 1608
rect 274 1611 280 1612
rect 274 1607 275 1611
rect 279 1607 280 1611
rect 274 1606 280 1607
rect 458 1611 464 1612
rect 458 1607 459 1611
rect 463 1607 464 1611
rect 458 1606 464 1607
rect 666 1611 672 1612
rect 666 1607 667 1611
rect 671 1607 672 1611
rect 666 1606 672 1607
rect 882 1611 888 1612
rect 882 1607 883 1611
rect 887 1607 888 1611
rect 882 1606 888 1607
rect 1114 1611 1120 1612
rect 1114 1607 1115 1611
rect 1119 1607 1120 1611
rect 1114 1606 1120 1607
rect 1354 1611 1360 1612
rect 1354 1607 1355 1611
rect 1359 1607 1360 1611
rect 1354 1606 1360 1607
rect 1594 1611 1600 1612
rect 1594 1607 1595 1611
rect 1599 1607 1600 1611
rect 1934 1608 1935 1612
rect 1939 1608 1940 1612
rect 1934 1607 1940 1608
rect 1594 1606 1600 1607
rect 302 1596 308 1597
rect 110 1595 116 1596
rect 110 1591 111 1595
rect 115 1591 116 1595
rect 302 1592 303 1596
rect 307 1592 308 1596
rect 302 1591 308 1592
rect 486 1596 492 1597
rect 486 1592 487 1596
rect 491 1592 492 1596
rect 486 1591 492 1592
rect 694 1596 700 1597
rect 694 1592 695 1596
rect 699 1592 700 1596
rect 694 1591 700 1592
rect 910 1596 916 1597
rect 910 1592 911 1596
rect 915 1592 916 1596
rect 910 1591 916 1592
rect 1142 1596 1148 1597
rect 1142 1592 1143 1596
rect 1147 1592 1148 1596
rect 1142 1591 1148 1592
rect 1382 1596 1388 1597
rect 1382 1592 1383 1596
rect 1387 1592 1388 1596
rect 1382 1591 1388 1592
rect 1622 1596 1628 1597
rect 1622 1592 1623 1596
rect 1627 1592 1628 1596
rect 1622 1591 1628 1592
rect 1934 1595 1940 1596
rect 1934 1591 1935 1595
rect 1939 1591 1940 1595
rect 110 1590 116 1591
rect 112 1567 114 1590
rect 304 1567 306 1591
rect 488 1567 490 1591
rect 696 1567 698 1591
rect 912 1567 914 1591
rect 1144 1567 1146 1591
rect 1384 1567 1386 1591
rect 1624 1567 1626 1591
rect 1934 1590 1940 1591
rect 1936 1567 1938 1590
rect 111 1566 115 1567
rect 111 1561 115 1562
rect 303 1566 307 1567
rect 303 1561 307 1562
rect 383 1566 387 1567
rect 383 1561 387 1562
rect 487 1566 491 1567
rect 487 1561 491 1562
rect 575 1566 579 1567
rect 575 1561 579 1562
rect 695 1566 699 1567
rect 695 1561 699 1562
rect 767 1566 771 1567
rect 767 1561 771 1562
rect 911 1566 915 1567
rect 911 1561 915 1562
rect 951 1566 955 1567
rect 951 1561 955 1562
rect 1127 1566 1131 1567
rect 1127 1561 1131 1562
rect 1143 1566 1147 1567
rect 1143 1561 1147 1562
rect 1303 1566 1307 1567
rect 1303 1561 1307 1562
rect 1383 1566 1387 1567
rect 1383 1561 1387 1562
rect 1479 1566 1483 1567
rect 1479 1561 1483 1562
rect 1623 1566 1627 1567
rect 1623 1561 1627 1562
rect 1663 1566 1667 1567
rect 1663 1561 1667 1562
rect 1935 1566 1939 1567
rect 1935 1561 1939 1562
rect 112 1538 114 1561
rect 110 1537 116 1538
rect 384 1537 386 1561
rect 576 1537 578 1561
rect 768 1537 770 1561
rect 952 1537 954 1561
rect 1128 1537 1130 1561
rect 1304 1537 1306 1561
rect 1480 1537 1482 1561
rect 1664 1537 1666 1561
rect 1936 1538 1938 1561
rect 1976 1547 1978 1619
rect 2204 1547 2206 1620
rect 2572 1547 2574 1620
rect 2940 1547 2942 1620
rect 3308 1547 3310 1620
rect 3652 1547 3654 1620
rect 3798 1619 3804 1620
rect 3800 1547 3802 1619
rect 3840 1613 3842 1673
rect 3838 1612 3844 1613
rect 3860 1612 3862 1673
rect 3996 1612 3998 1673
rect 4132 1612 4134 1673
rect 4284 1612 4286 1673
rect 4484 1612 4486 1673
rect 4716 1612 4718 1673
rect 4980 1612 4982 1673
rect 5260 1612 5262 1673
rect 5516 1612 5518 1673
rect 5664 1613 5666 1673
rect 5662 1612 5668 1613
rect 3838 1608 3839 1612
rect 3843 1608 3844 1612
rect 3838 1607 3844 1608
rect 3858 1611 3864 1612
rect 3858 1607 3859 1611
rect 3863 1607 3864 1611
rect 3858 1606 3864 1607
rect 3994 1611 4000 1612
rect 3994 1607 3995 1611
rect 3999 1607 4000 1611
rect 3994 1606 4000 1607
rect 4130 1611 4136 1612
rect 4130 1607 4131 1611
rect 4135 1607 4136 1611
rect 4130 1606 4136 1607
rect 4282 1611 4288 1612
rect 4282 1607 4283 1611
rect 4287 1607 4288 1611
rect 4282 1606 4288 1607
rect 4482 1611 4488 1612
rect 4482 1607 4483 1611
rect 4487 1607 4488 1611
rect 4482 1606 4488 1607
rect 4714 1611 4720 1612
rect 4714 1607 4715 1611
rect 4719 1607 4720 1611
rect 4714 1606 4720 1607
rect 4978 1611 4984 1612
rect 4978 1607 4979 1611
rect 4983 1607 4984 1611
rect 4978 1606 4984 1607
rect 5258 1611 5264 1612
rect 5258 1607 5259 1611
rect 5263 1607 5264 1611
rect 5258 1606 5264 1607
rect 5514 1611 5520 1612
rect 5514 1607 5515 1611
rect 5519 1607 5520 1611
rect 5662 1608 5663 1612
rect 5667 1608 5668 1612
rect 5662 1607 5668 1608
rect 5514 1606 5520 1607
rect 3886 1596 3892 1597
rect 3838 1595 3844 1596
rect 3838 1591 3839 1595
rect 3843 1591 3844 1595
rect 3886 1592 3887 1596
rect 3891 1592 3892 1596
rect 3886 1591 3892 1592
rect 4022 1596 4028 1597
rect 4022 1592 4023 1596
rect 4027 1592 4028 1596
rect 4022 1591 4028 1592
rect 4158 1596 4164 1597
rect 4158 1592 4159 1596
rect 4163 1592 4164 1596
rect 4158 1591 4164 1592
rect 4310 1596 4316 1597
rect 4310 1592 4311 1596
rect 4315 1592 4316 1596
rect 4310 1591 4316 1592
rect 4510 1596 4516 1597
rect 4510 1592 4511 1596
rect 4515 1592 4516 1596
rect 4510 1591 4516 1592
rect 4742 1596 4748 1597
rect 4742 1592 4743 1596
rect 4747 1592 4748 1596
rect 4742 1591 4748 1592
rect 5006 1596 5012 1597
rect 5006 1592 5007 1596
rect 5011 1592 5012 1596
rect 5006 1591 5012 1592
rect 5286 1596 5292 1597
rect 5286 1592 5287 1596
rect 5291 1592 5292 1596
rect 5286 1591 5292 1592
rect 5542 1596 5548 1597
rect 5542 1592 5543 1596
rect 5547 1592 5548 1596
rect 5542 1591 5548 1592
rect 5662 1595 5668 1596
rect 5662 1591 5663 1595
rect 5667 1591 5668 1595
rect 3838 1590 3844 1591
rect 3840 1567 3842 1590
rect 3888 1567 3890 1591
rect 4024 1567 4026 1591
rect 4160 1567 4162 1591
rect 4312 1567 4314 1591
rect 4512 1567 4514 1591
rect 4744 1567 4746 1591
rect 5008 1567 5010 1591
rect 5288 1567 5290 1591
rect 5544 1567 5546 1591
rect 5662 1590 5668 1591
rect 5664 1567 5666 1590
rect 3839 1566 3843 1567
rect 3839 1561 3843 1562
rect 3887 1566 3891 1567
rect 3887 1561 3891 1562
rect 4023 1566 4027 1567
rect 4023 1561 4027 1562
rect 4047 1566 4051 1567
rect 4047 1561 4051 1562
rect 4159 1566 4163 1567
rect 4159 1561 4163 1562
rect 4271 1566 4275 1567
rect 4271 1561 4275 1562
rect 4311 1566 4315 1567
rect 4311 1561 4315 1562
rect 4511 1566 4515 1567
rect 4511 1561 4515 1562
rect 4543 1566 4547 1567
rect 4543 1561 4547 1562
rect 4743 1566 4747 1567
rect 4743 1561 4747 1562
rect 4855 1566 4859 1567
rect 4855 1561 4859 1562
rect 5007 1566 5011 1567
rect 5007 1561 5011 1562
rect 5191 1566 5195 1567
rect 5191 1561 5195 1562
rect 5287 1566 5291 1567
rect 5287 1561 5291 1562
rect 5527 1566 5531 1567
rect 5527 1561 5531 1562
rect 5543 1566 5547 1567
rect 5543 1561 5547 1562
rect 5663 1566 5667 1567
rect 5663 1561 5667 1562
rect 1975 1546 1979 1547
rect 1975 1541 1979 1542
rect 1995 1546 1999 1547
rect 1995 1541 1999 1542
rect 2203 1546 2207 1547
rect 2203 1541 2207 1542
rect 2275 1546 2279 1547
rect 2275 1541 2279 1542
rect 2539 1546 2543 1547
rect 2539 1541 2543 1542
rect 2571 1546 2575 1547
rect 2571 1541 2575 1542
rect 2779 1546 2783 1547
rect 2779 1541 2783 1542
rect 2939 1546 2943 1547
rect 2939 1541 2943 1542
rect 3011 1546 3015 1547
rect 3011 1541 3015 1542
rect 3235 1546 3239 1547
rect 3235 1541 3239 1542
rect 3307 1546 3311 1547
rect 3307 1541 3311 1542
rect 3451 1546 3455 1547
rect 3451 1541 3455 1542
rect 3651 1546 3655 1547
rect 3651 1541 3655 1542
rect 3799 1546 3803 1547
rect 3799 1541 3803 1542
rect 1934 1537 1940 1538
rect 110 1533 111 1537
rect 115 1533 116 1537
rect 110 1532 116 1533
rect 382 1536 388 1537
rect 382 1532 383 1536
rect 387 1532 388 1536
rect 382 1531 388 1532
rect 574 1536 580 1537
rect 574 1532 575 1536
rect 579 1532 580 1536
rect 574 1531 580 1532
rect 766 1536 772 1537
rect 766 1532 767 1536
rect 771 1532 772 1536
rect 766 1531 772 1532
rect 950 1536 956 1537
rect 950 1532 951 1536
rect 955 1532 956 1536
rect 950 1531 956 1532
rect 1126 1536 1132 1537
rect 1126 1532 1127 1536
rect 1131 1532 1132 1536
rect 1126 1531 1132 1532
rect 1302 1536 1308 1537
rect 1302 1532 1303 1536
rect 1307 1532 1308 1536
rect 1302 1531 1308 1532
rect 1478 1536 1484 1537
rect 1478 1532 1479 1536
rect 1483 1532 1484 1536
rect 1478 1531 1484 1532
rect 1662 1536 1668 1537
rect 1662 1532 1663 1536
rect 1667 1532 1668 1536
rect 1934 1533 1935 1537
rect 1939 1533 1940 1537
rect 1934 1532 1940 1533
rect 1662 1531 1668 1532
rect 354 1521 360 1522
rect 110 1520 116 1521
rect 110 1516 111 1520
rect 115 1516 116 1520
rect 354 1517 355 1521
rect 359 1517 360 1521
rect 354 1516 360 1517
rect 546 1521 552 1522
rect 546 1517 547 1521
rect 551 1517 552 1521
rect 546 1516 552 1517
rect 738 1521 744 1522
rect 738 1517 739 1521
rect 743 1517 744 1521
rect 738 1516 744 1517
rect 922 1521 928 1522
rect 922 1517 923 1521
rect 927 1517 928 1521
rect 922 1516 928 1517
rect 1098 1521 1104 1522
rect 1098 1517 1099 1521
rect 1103 1517 1104 1521
rect 1098 1516 1104 1517
rect 1274 1521 1280 1522
rect 1274 1517 1275 1521
rect 1279 1517 1280 1521
rect 1274 1516 1280 1517
rect 1450 1521 1456 1522
rect 1450 1517 1451 1521
rect 1455 1517 1456 1521
rect 1450 1516 1456 1517
rect 1634 1521 1640 1522
rect 1634 1517 1635 1521
rect 1639 1517 1640 1521
rect 1634 1516 1640 1517
rect 1934 1520 1940 1521
rect 1934 1516 1935 1520
rect 1939 1516 1940 1520
rect 110 1515 116 1516
rect 112 1435 114 1515
rect 356 1435 358 1516
rect 548 1435 550 1516
rect 740 1435 742 1516
rect 924 1435 926 1516
rect 1100 1435 1102 1516
rect 1276 1435 1278 1516
rect 1452 1435 1454 1516
rect 1636 1435 1638 1516
rect 1934 1515 1940 1516
rect 1936 1435 1938 1515
rect 1976 1481 1978 1541
rect 1974 1480 1980 1481
rect 1996 1480 1998 1541
rect 2276 1480 2278 1541
rect 2540 1480 2542 1541
rect 2780 1480 2782 1541
rect 3012 1480 3014 1541
rect 3236 1480 3238 1541
rect 3452 1480 3454 1541
rect 3652 1480 3654 1541
rect 3800 1481 3802 1541
rect 3840 1538 3842 1561
rect 3838 1537 3844 1538
rect 3888 1537 3890 1561
rect 4048 1537 4050 1561
rect 4272 1537 4274 1561
rect 4544 1537 4546 1561
rect 4856 1537 4858 1561
rect 5192 1537 5194 1561
rect 5528 1537 5530 1561
rect 5664 1538 5666 1561
rect 5662 1537 5668 1538
rect 3838 1533 3839 1537
rect 3843 1533 3844 1537
rect 3838 1532 3844 1533
rect 3886 1536 3892 1537
rect 3886 1532 3887 1536
rect 3891 1532 3892 1536
rect 3886 1531 3892 1532
rect 4046 1536 4052 1537
rect 4046 1532 4047 1536
rect 4051 1532 4052 1536
rect 4046 1531 4052 1532
rect 4270 1536 4276 1537
rect 4270 1532 4271 1536
rect 4275 1532 4276 1536
rect 4270 1531 4276 1532
rect 4542 1536 4548 1537
rect 4542 1532 4543 1536
rect 4547 1532 4548 1536
rect 4542 1531 4548 1532
rect 4854 1536 4860 1537
rect 4854 1532 4855 1536
rect 4859 1532 4860 1536
rect 4854 1531 4860 1532
rect 5190 1536 5196 1537
rect 5190 1532 5191 1536
rect 5195 1532 5196 1536
rect 5190 1531 5196 1532
rect 5526 1536 5532 1537
rect 5526 1532 5527 1536
rect 5531 1532 5532 1536
rect 5662 1533 5663 1537
rect 5667 1533 5668 1537
rect 5662 1532 5668 1533
rect 5526 1531 5532 1532
rect 3858 1521 3864 1522
rect 3838 1520 3844 1521
rect 3838 1516 3839 1520
rect 3843 1516 3844 1520
rect 3858 1517 3859 1521
rect 3863 1517 3864 1521
rect 3858 1516 3864 1517
rect 4018 1521 4024 1522
rect 4018 1517 4019 1521
rect 4023 1517 4024 1521
rect 4018 1516 4024 1517
rect 4242 1521 4248 1522
rect 4242 1517 4243 1521
rect 4247 1517 4248 1521
rect 4242 1516 4248 1517
rect 4514 1521 4520 1522
rect 4514 1517 4515 1521
rect 4519 1517 4520 1521
rect 4514 1516 4520 1517
rect 4826 1521 4832 1522
rect 4826 1517 4827 1521
rect 4831 1517 4832 1521
rect 4826 1516 4832 1517
rect 5162 1521 5168 1522
rect 5162 1517 5163 1521
rect 5167 1517 5168 1521
rect 5162 1516 5168 1517
rect 5498 1521 5504 1522
rect 5498 1517 5499 1521
rect 5503 1517 5504 1521
rect 5498 1516 5504 1517
rect 5662 1520 5668 1521
rect 5662 1516 5663 1520
rect 5667 1516 5668 1520
rect 3838 1515 3844 1516
rect 3798 1480 3804 1481
rect 1974 1476 1975 1480
rect 1979 1476 1980 1480
rect 1974 1475 1980 1476
rect 1994 1479 2000 1480
rect 1994 1475 1995 1479
rect 1999 1475 2000 1479
rect 1994 1474 2000 1475
rect 2274 1479 2280 1480
rect 2274 1475 2275 1479
rect 2279 1475 2280 1479
rect 2274 1474 2280 1475
rect 2538 1479 2544 1480
rect 2538 1475 2539 1479
rect 2543 1475 2544 1479
rect 2538 1474 2544 1475
rect 2778 1479 2784 1480
rect 2778 1475 2779 1479
rect 2783 1475 2784 1479
rect 2778 1474 2784 1475
rect 3010 1479 3016 1480
rect 3010 1475 3011 1479
rect 3015 1475 3016 1479
rect 3010 1474 3016 1475
rect 3234 1479 3240 1480
rect 3234 1475 3235 1479
rect 3239 1475 3240 1479
rect 3234 1474 3240 1475
rect 3450 1479 3456 1480
rect 3450 1475 3451 1479
rect 3455 1475 3456 1479
rect 3450 1474 3456 1475
rect 3650 1479 3656 1480
rect 3650 1475 3651 1479
rect 3655 1475 3656 1479
rect 3798 1476 3799 1480
rect 3803 1476 3804 1480
rect 3798 1475 3804 1476
rect 3650 1474 3656 1475
rect 2022 1464 2028 1465
rect 1974 1463 1980 1464
rect 1974 1459 1975 1463
rect 1979 1459 1980 1463
rect 2022 1460 2023 1464
rect 2027 1460 2028 1464
rect 2022 1459 2028 1460
rect 2302 1464 2308 1465
rect 2302 1460 2303 1464
rect 2307 1460 2308 1464
rect 2302 1459 2308 1460
rect 2566 1464 2572 1465
rect 2566 1460 2567 1464
rect 2571 1460 2572 1464
rect 2566 1459 2572 1460
rect 2806 1464 2812 1465
rect 2806 1460 2807 1464
rect 2811 1460 2812 1464
rect 2806 1459 2812 1460
rect 3038 1464 3044 1465
rect 3038 1460 3039 1464
rect 3043 1460 3044 1464
rect 3038 1459 3044 1460
rect 3262 1464 3268 1465
rect 3262 1460 3263 1464
rect 3267 1460 3268 1464
rect 3262 1459 3268 1460
rect 3478 1464 3484 1465
rect 3478 1460 3479 1464
rect 3483 1460 3484 1464
rect 3478 1459 3484 1460
rect 3678 1464 3684 1465
rect 3678 1460 3679 1464
rect 3683 1460 3684 1464
rect 3678 1459 3684 1460
rect 3798 1463 3804 1464
rect 3798 1459 3799 1463
rect 3803 1459 3804 1463
rect 1974 1458 1980 1459
rect 1976 1435 1978 1458
rect 2024 1435 2026 1459
rect 2304 1435 2306 1459
rect 2568 1435 2570 1459
rect 2808 1435 2810 1459
rect 3040 1435 3042 1459
rect 3264 1435 3266 1459
rect 3480 1435 3482 1459
rect 3680 1435 3682 1459
rect 3798 1458 3804 1459
rect 3800 1435 3802 1458
rect 3840 1439 3842 1515
rect 3860 1439 3862 1516
rect 4020 1439 4022 1516
rect 4244 1439 4246 1516
rect 4516 1439 4518 1516
rect 4828 1439 4830 1516
rect 5164 1439 5166 1516
rect 5500 1439 5502 1516
rect 5662 1515 5668 1516
rect 5664 1439 5666 1515
rect 3839 1438 3843 1439
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 331 1434 335 1435
rect 331 1429 335 1430
rect 355 1434 359 1435
rect 355 1429 359 1430
rect 547 1434 551 1435
rect 547 1429 551 1430
rect 587 1434 591 1435
rect 587 1429 591 1430
rect 739 1434 743 1435
rect 739 1429 743 1430
rect 843 1434 847 1435
rect 843 1429 847 1430
rect 923 1434 927 1435
rect 923 1429 927 1430
rect 1099 1434 1103 1435
rect 1099 1429 1103 1430
rect 1275 1434 1279 1435
rect 1275 1429 1279 1430
rect 1363 1434 1367 1435
rect 1363 1429 1367 1430
rect 1451 1434 1455 1435
rect 1451 1429 1455 1430
rect 1635 1434 1639 1435
rect 1635 1429 1639 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 1975 1434 1979 1435
rect 1975 1429 1979 1430
rect 2023 1434 2027 1435
rect 2023 1429 2027 1430
rect 2191 1434 2195 1435
rect 2191 1429 2195 1430
rect 2303 1434 2307 1435
rect 2303 1429 2307 1430
rect 2399 1434 2403 1435
rect 2399 1429 2403 1430
rect 2567 1434 2571 1435
rect 2567 1429 2571 1430
rect 2615 1434 2619 1435
rect 2615 1429 2619 1430
rect 2807 1434 2811 1435
rect 2807 1429 2811 1430
rect 2831 1434 2835 1435
rect 2831 1429 2835 1430
rect 3039 1434 3043 1435
rect 3039 1429 3043 1430
rect 3055 1434 3059 1435
rect 3055 1429 3059 1430
rect 3263 1434 3267 1435
rect 3263 1429 3267 1430
rect 3287 1434 3291 1435
rect 3287 1429 3291 1430
rect 3479 1434 3483 1435
rect 3479 1429 3483 1430
rect 3527 1434 3531 1435
rect 3527 1429 3531 1430
rect 3679 1434 3683 1435
rect 3679 1429 3683 1430
rect 3799 1434 3803 1435
rect 3839 1433 3843 1434
rect 3859 1438 3863 1439
rect 3859 1433 3863 1434
rect 3995 1438 3999 1439
rect 3995 1433 3999 1434
rect 4019 1438 4023 1439
rect 4019 1433 4023 1434
rect 4147 1438 4151 1439
rect 4147 1433 4151 1434
rect 4243 1438 4247 1439
rect 4243 1433 4247 1434
rect 4355 1438 4359 1439
rect 4355 1433 4359 1434
rect 4515 1438 4519 1439
rect 4515 1433 4519 1434
rect 4595 1438 4599 1439
rect 4595 1433 4599 1434
rect 4827 1438 4831 1439
rect 4827 1433 4831 1434
rect 4867 1438 4871 1439
rect 4867 1433 4871 1434
rect 5163 1438 5167 1439
rect 5163 1433 5167 1434
rect 5459 1438 5463 1439
rect 5459 1433 5463 1434
rect 5499 1438 5503 1439
rect 5499 1433 5503 1434
rect 5663 1438 5667 1439
rect 5663 1433 5667 1434
rect 3799 1429 3803 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 332 1368 334 1429
rect 588 1368 590 1429
rect 844 1368 846 1429
rect 1100 1368 1102 1429
rect 1364 1368 1366 1429
rect 1936 1369 1938 1429
rect 1976 1406 1978 1429
rect 1974 1405 1980 1406
rect 2024 1405 2026 1429
rect 2192 1405 2194 1429
rect 2400 1405 2402 1429
rect 2616 1405 2618 1429
rect 2832 1405 2834 1429
rect 3056 1405 3058 1429
rect 3288 1405 3290 1429
rect 3528 1405 3530 1429
rect 3800 1406 3802 1429
rect 3798 1405 3804 1406
rect 1974 1401 1975 1405
rect 1979 1401 1980 1405
rect 1974 1400 1980 1401
rect 2022 1404 2028 1405
rect 2022 1400 2023 1404
rect 2027 1400 2028 1404
rect 2022 1399 2028 1400
rect 2190 1404 2196 1405
rect 2190 1400 2191 1404
rect 2195 1400 2196 1404
rect 2190 1399 2196 1400
rect 2398 1404 2404 1405
rect 2398 1400 2399 1404
rect 2403 1400 2404 1404
rect 2398 1399 2404 1400
rect 2614 1404 2620 1405
rect 2614 1400 2615 1404
rect 2619 1400 2620 1404
rect 2614 1399 2620 1400
rect 2830 1404 2836 1405
rect 2830 1400 2831 1404
rect 2835 1400 2836 1404
rect 2830 1399 2836 1400
rect 3054 1404 3060 1405
rect 3054 1400 3055 1404
rect 3059 1400 3060 1404
rect 3054 1399 3060 1400
rect 3286 1404 3292 1405
rect 3286 1400 3287 1404
rect 3291 1400 3292 1404
rect 3286 1399 3292 1400
rect 3526 1404 3532 1405
rect 3526 1400 3527 1404
rect 3531 1400 3532 1404
rect 3798 1401 3799 1405
rect 3803 1401 3804 1405
rect 3798 1400 3804 1401
rect 3526 1399 3532 1400
rect 1994 1389 2000 1390
rect 1974 1388 1980 1389
rect 1974 1384 1975 1388
rect 1979 1384 1980 1388
rect 1994 1385 1995 1389
rect 1999 1385 2000 1389
rect 1994 1384 2000 1385
rect 2162 1389 2168 1390
rect 2162 1385 2163 1389
rect 2167 1385 2168 1389
rect 2162 1384 2168 1385
rect 2370 1389 2376 1390
rect 2370 1385 2371 1389
rect 2375 1385 2376 1389
rect 2370 1384 2376 1385
rect 2586 1389 2592 1390
rect 2586 1385 2587 1389
rect 2591 1385 2592 1389
rect 2586 1384 2592 1385
rect 2802 1389 2808 1390
rect 2802 1385 2803 1389
rect 2807 1385 2808 1389
rect 2802 1384 2808 1385
rect 3026 1389 3032 1390
rect 3026 1385 3027 1389
rect 3031 1385 3032 1389
rect 3026 1384 3032 1385
rect 3258 1389 3264 1390
rect 3258 1385 3259 1389
rect 3263 1385 3264 1389
rect 3258 1384 3264 1385
rect 3498 1389 3504 1390
rect 3498 1385 3499 1389
rect 3503 1385 3504 1389
rect 3498 1384 3504 1385
rect 3798 1388 3804 1389
rect 3798 1384 3799 1388
rect 3803 1384 3804 1388
rect 1974 1383 1980 1384
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 330 1367 336 1368
rect 330 1363 331 1367
rect 335 1363 336 1367
rect 330 1362 336 1363
rect 586 1367 592 1368
rect 586 1363 587 1367
rect 591 1363 592 1367
rect 586 1362 592 1363
rect 842 1367 848 1368
rect 842 1363 843 1367
rect 847 1363 848 1367
rect 842 1362 848 1363
rect 1098 1367 1104 1368
rect 1098 1363 1099 1367
rect 1103 1363 1104 1367
rect 1098 1362 1104 1363
rect 1362 1367 1368 1368
rect 1362 1363 1363 1367
rect 1367 1363 1368 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1362 1362 1368 1363
rect 358 1352 364 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 358 1348 359 1352
rect 363 1348 364 1352
rect 358 1347 364 1348
rect 614 1352 620 1353
rect 614 1348 615 1352
rect 619 1348 620 1352
rect 614 1347 620 1348
rect 870 1352 876 1353
rect 870 1348 871 1352
rect 875 1348 876 1352
rect 870 1347 876 1348
rect 1126 1352 1132 1353
rect 1126 1348 1127 1352
rect 1131 1348 1132 1352
rect 1126 1347 1132 1348
rect 1390 1352 1396 1353
rect 1390 1348 1391 1352
rect 1395 1348 1396 1352
rect 1390 1347 1396 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 360 1323 362 1347
rect 616 1323 618 1347
rect 872 1323 874 1347
rect 1128 1323 1130 1347
rect 1392 1323 1394 1347
rect 1934 1346 1940 1347
rect 1936 1323 1938 1346
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 359 1322 363 1323
rect 359 1317 363 1318
rect 367 1322 371 1323
rect 367 1317 371 1318
rect 551 1322 555 1323
rect 551 1317 555 1318
rect 615 1322 619 1323
rect 615 1317 619 1318
rect 727 1322 731 1323
rect 727 1317 731 1318
rect 871 1322 875 1323
rect 871 1317 875 1318
rect 895 1322 899 1323
rect 895 1317 899 1318
rect 1063 1322 1067 1323
rect 1063 1317 1067 1318
rect 1127 1322 1131 1323
rect 1127 1317 1131 1318
rect 1223 1322 1227 1323
rect 1223 1317 1227 1318
rect 1375 1322 1379 1323
rect 1375 1317 1379 1318
rect 1391 1322 1395 1323
rect 1391 1317 1395 1318
rect 1527 1322 1531 1323
rect 1527 1317 1531 1318
rect 1679 1322 1683 1323
rect 1679 1317 1683 1318
rect 1815 1322 1819 1323
rect 1815 1317 1819 1318
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 368 1293 370 1317
rect 552 1293 554 1317
rect 728 1293 730 1317
rect 896 1293 898 1317
rect 1064 1293 1066 1317
rect 1224 1293 1226 1317
rect 1376 1293 1378 1317
rect 1528 1293 1530 1317
rect 1680 1293 1682 1317
rect 1816 1293 1818 1317
rect 1936 1294 1938 1317
rect 1976 1303 1978 1383
rect 1996 1303 1998 1384
rect 2164 1303 2166 1384
rect 2372 1303 2374 1384
rect 2588 1303 2590 1384
rect 2804 1303 2806 1384
rect 3028 1303 3030 1384
rect 3260 1303 3262 1384
rect 3500 1303 3502 1384
rect 3798 1383 3804 1384
rect 3800 1303 3802 1383
rect 3840 1373 3842 1433
rect 3838 1372 3844 1373
rect 3860 1372 3862 1433
rect 3996 1372 3998 1433
rect 4148 1372 4150 1433
rect 4356 1372 4358 1433
rect 4596 1372 4598 1433
rect 4868 1372 4870 1433
rect 5164 1372 5166 1433
rect 5460 1372 5462 1433
rect 5664 1373 5666 1433
rect 5662 1372 5668 1373
rect 3838 1368 3839 1372
rect 3843 1368 3844 1372
rect 3838 1367 3844 1368
rect 3858 1371 3864 1372
rect 3858 1367 3859 1371
rect 3863 1367 3864 1371
rect 3858 1366 3864 1367
rect 3994 1371 4000 1372
rect 3994 1367 3995 1371
rect 3999 1367 4000 1371
rect 3994 1366 4000 1367
rect 4146 1371 4152 1372
rect 4146 1367 4147 1371
rect 4151 1367 4152 1371
rect 4146 1366 4152 1367
rect 4354 1371 4360 1372
rect 4354 1367 4355 1371
rect 4359 1367 4360 1371
rect 4354 1366 4360 1367
rect 4594 1371 4600 1372
rect 4594 1367 4595 1371
rect 4599 1367 4600 1371
rect 4594 1366 4600 1367
rect 4866 1371 4872 1372
rect 4866 1367 4867 1371
rect 4871 1367 4872 1371
rect 4866 1366 4872 1367
rect 5162 1371 5168 1372
rect 5162 1367 5163 1371
rect 5167 1367 5168 1371
rect 5162 1366 5168 1367
rect 5458 1371 5464 1372
rect 5458 1367 5459 1371
rect 5463 1367 5464 1371
rect 5662 1368 5663 1372
rect 5667 1368 5668 1372
rect 5662 1367 5668 1368
rect 5458 1366 5464 1367
rect 3886 1356 3892 1357
rect 3838 1355 3844 1356
rect 3838 1351 3839 1355
rect 3843 1351 3844 1355
rect 3886 1352 3887 1356
rect 3891 1352 3892 1356
rect 3886 1351 3892 1352
rect 4022 1356 4028 1357
rect 4022 1352 4023 1356
rect 4027 1352 4028 1356
rect 4022 1351 4028 1352
rect 4174 1356 4180 1357
rect 4174 1352 4175 1356
rect 4179 1352 4180 1356
rect 4174 1351 4180 1352
rect 4382 1356 4388 1357
rect 4382 1352 4383 1356
rect 4387 1352 4388 1356
rect 4382 1351 4388 1352
rect 4622 1356 4628 1357
rect 4622 1352 4623 1356
rect 4627 1352 4628 1356
rect 4622 1351 4628 1352
rect 4894 1356 4900 1357
rect 4894 1352 4895 1356
rect 4899 1352 4900 1356
rect 4894 1351 4900 1352
rect 5190 1356 5196 1357
rect 5190 1352 5191 1356
rect 5195 1352 5196 1356
rect 5190 1351 5196 1352
rect 5486 1356 5492 1357
rect 5486 1352 5487 1356
rect 5491 1352 5492 1356
rect 5486 1351 5492 1352
rect 5662 1355 5668 1356
rect 5662 1351 5663 1355
rect 5667 1351 5668 1355
rect 3838 1350 3844 1351
rect 3840 1323 3842 1350
rect 3888 1323 3890 1351
rect 4024 1323 4026 1351
rect 4176 1323 4178 1351
rect 4384 1323 4386 1351
rect 4624 1323 4626 1351
rect 4896 1323 4898 1351
rect 5192 1323 5194 1351
rect 5488 1323 5490 1351
rect 5662 1350 5668 1351
rect 5664 1323 5666 1350
rect 3839 1322 3843 1323
rect 3839 1317 3843 1318
rect 3887 1322 3891 1323
rect 3887 1317 3891 1318
rect 4023 1322 4027 1323
rect 4023 1317 4027 1318
rect 4047 1322 4051 1323
rect 4047 1317 4051 1318
rect 4175 1322 4179 1323
rect 4175 1317 4179 1318
rect 4239 1322 4243 1323
rect 4239 1317 4243 1318
rect 4383 1322 4387 1323
rect 4383 1317 4387 1318
rect 4455 1322 4459 1323
rect 4455 1317 4459 1318
rect 4623 1322 4627 1323
rect 4623 1317 4627 1318
rect 4695 1322 4699 1323
rect 4695 1317 4699 1318
rect 4895 1322 4899 1323
rect 4895 1317 4899 1318
rect 4951 1322 4955 1323
rect 4951 1317 4955 1318
rect 5191 1322 5195 1323
rect 5191 1317 5195 1318
rect 5223 1322 5227 1323
rect 5223 1317 5227 1318
rect 5487 1322 5491 1323
rect 5487 1317 5491 1318
rect 5495 1322 5499 1323
rect 5495 1317 5499 1318
rect 5663 1322 5667 1323
rect 5663 1317 5667 1318
rect 1975 1302 1979 1303
rect 1975 1297 1979 1298
rect 1995 1302 1999 1303
rect 1995 1297 1999 1298
rect 2163 1302 2167 1303
rect 2163 1297 2167 1298
rect 2371 1302 2375 1303
rect 2371 1297 2375 1298
rect 2587 1302 2591 1303
rect 2587 1297 2591 1298
rect 2803 1302 2807 1303
rect 2803 1297 2807 1298
rect 3027 1302 3031 1303
rect 3027 1297 3031 1298
rect 3091 1302 3095 1303
rect 3091 1297 3095 1298
rect 3227 1302 3231 1303
rect 3227 1297 3231 1298
rect 3259 1302 3263 1303
rect 3259 1297 3263 1298
rect 3363 1302 3367 1303
rect 3363 1297 3367 1298
rect 3499 1302 3503 1303
rect 3499 1297 3503 1298
rect 3799 1302 3803 1303
rect 3799 1297 3803 1298
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 366 1292 372 1293
rect 366 1288 367 1292
rect 371 1288 372 1292
rect 366 1287 372 1288
rect 550 1292 556 1293
rect 550 1288 551 1292
rect 555 1288 556 1292
rect 550 1287 556 1288
rect 726 1292 732 1293
rect 726 1288 727 1292
rect 731 1288 732 1292
rect 726 1287 732 1288
rect 894 1292 900 1293
rect 894 1288 895 1292
rect 899 1288 900 1292
rect 894 1287 900 1288
rect 1062 1292 1068 1293
rect 1062 1288 1063 1292
rect 1067 1288 1068 1292
rect 1062 1287 1068 1288
rect 1222 1292 1228 1293
rect 1222 1288 1223 1292
rect 1227 1288 1228 1292
rect 1222 1287 1228 1288
rect 1374 1292 1380 1293
rect 1374 1288 1375 1292
rect 1379 1288 1380 1292
rect 1374 1287 1380 1288
rect 1526 1292 1532 1293
rect 1526 1288 1527 1292
rect 1531 1288 1532 1292
rect 1526 1287 1532 1288
rect 1678 1292 1684 1293
rect 1678 1288 1679 1292
rect 1683 1288 1684 1292
rect 1678 1287 1684 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 338 1277 344 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 338 1273 339 1277
rect 343 1273 344 1277
rect 338 1272 344 1273
rect 522 1277 528 1278
rect 522 1273 523 1277
rect 527 1273 528 1277
rect 522 1272 528 1273
rect 698 1277 704 1278
rect 698 1273 699 1277
rect 703 1273 704 1277
rect 698 1272 704 1273
rect 866 1277 872 1278
rect 866 1273 867 1277
rect 871 1273 872 1277
rect 866 1272 872 1273
rect 1034 1277 1040 1278
rect 1034 1273 1035 1277
rect 1039 1273 1040 1277
rect 1034 1272 1040 1273
rect 1194 1277 1200 1278
rect 1194 1273 1195 1277
rect 1199 1273 1200 1277
rect 1194 1272 1200 1273
rect 1346 1277 1352 1278
rect 1346 1273 1347 1277
rect 1351 1273 1352 1277
rect 1346 1272 1352 1273
rect 1498 1277 1504 1278
rect 1498 1273 1499 1277
rect 1503 1273 1504 1277
rect 1498 1272 1504 1273
rect 1650 1277 1656 1278
rect 1650 1273 1651 1277
rect 1655 1273 1656 1277
rect 1650 1272 1656 1273
rect 1786 1277 1792 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 112 1199 114 1271
rect 340 1199 342 1272
rect 524 1199 526 1272
rect 700 1199 702 1272
rect 868 1199 870 1272
rect 1036 1199 1038 1272
rect 1196 1199 1198 1272
rect 1348 1199 1350 1272
rect 1500 1199 1502 1272
rect 1652 1199 1654 1272
rect 1788 1199 1790 1272
rect 1934 1271 1940 1272
rect 1936 1199 1938 1271
rect 1976 1237 1978 1297
rect 1974 1236 1980 1237
rect 3092 1236 3094 1297
rect 3228 1236 3230 1297
rect 3364 1236 3366 1297
rect 3800 1237 3802 1297
rect 3840 1294 3842 1317
rect 3838 1293 3844 1294
rect 3888 1293 3890 1317
rect 4048 1293 4050 1317
rect 4240 1293 4242 1317
rect 4456 1293 4458 1317
rect 4696 1293 4698 1317
rect 4952 1293 4954 1317
rect 5224 1293 5226 1317
rect 5496 1293 5498 1317
rect 5664 1294 5666 1317
rect 5662 1293 5668 1294
rect 3838 1289 3839 1293
rect 3843 1289 3844 1293
rect 3838 1288 3844 1289
rect 3886 1292 3892 1293
rect 3886 1288 3887 1292
rect 3891 1288 3892 1292
rect 3886 1287 3892 1288
rect 4046 1292 4052 1293
rect 4046 1288 4047 1292
rect 4051 1288 4052 1292
rect 4046 1287 4052 1288
rect 4238 1292 4244 1293
rect 4238 1288 4239 1292
rect 4243 1288 4244 1292
rect 4238 1287 4244 1288
rect 4454 1292 4460 1293
rect 4454 1288 4455 1292
rect 4459 1288 4460 1292
rect 4454 1287 4460 1288
rect 4694 1292 4700 1293
rect 4694 1288 4695 1292
rect 4699 1288 4700 1292
rect 4694 1287 4700 1288
rect 4950 1292 4956 1293
rect 4950 1288 4951 1292
rect 4955 1288 4956 1292
rect 4950 1287 4956 1288
rect 5222 1292 5228 1293
rect 5222 1288 5223 1292
rect 5227 1288 5228 1292
rect 5222 1287 5228 1288
rect 5494 1292 5500 1293
rect 5494 1288 5495 1292
rect 5499 1288 5500 1292
rect 5662 1289 5663 1293
rect 5667 1289 5668 1293
rect 5662 1288 5668 1289
rect 5494 1287 5500 1288
rect 3858 1277 3864 1278
rect 3838 1276 3844 1277
rect 3838 1272 3839 1276
rect 3843 1272 3844 1276
rect 3858 1273 3859 1277
rect 3863 1273 3864 1277
rect 3858 1272 3864 1273
rect 4018 1277 4024 1278
rect 4018 1273 4019 1277
rect 4023 1273 4024 1277
rect 4018 1272 4024 1273
rect 4210 1277 4216 1278
rect 4210 1273 4211 1277
rect 4215 1273 4216 1277
rect 4210 1272 4216 1273
rect 4426 1277 4432 1278
rect 4426 1273 4427 1277
rect 4431 1273 4432 1277
rect 4426 1272 4432 1273
rect 4666 1277 4672 1278
rect 4666 1273 4667 1277
rect 4671 1273 4672 1277
rect 4666 1272 4672 1273
rect 4922 1277 4928 1278
rect 4922 1273 4923 1277
rect 4927 1273 4928 1277
rect 4922 1272 4928 1273
rect 5194 1277 5200 1278
rect 5194 1273 5195 1277
rect 5199 1273 5200 1277
rect 5194 1272 5200 1273
rect 5466 1277 5472 1278
rect 5466 1273 5467 1277
rect 5471 1273 5472 1277
rect 5466 1272 5472 1273
rect 5662 1276 5668 1277
rect 5662 1272 5663 1276
rect 5667 1272 5668 1276
rect 3838 1271 3844 1272
rect 3798 1236 3804 1237
rect 1974 1232 1975 1236
rect 1979 1232 1980 1236
rect 1974 1231 1980 1232
rect 3090 1235 3096 1236
rect 3090 1231 3091 1235
rect 3095 1231 3096 1235
rect 3090 1230 3096 1231
rect 3226 1235 3232 1236
rect 3226 1231 3227 1235
rect 3231 1231 3232 1235
rect 3226 1230 3232 1231
rect 3362 1235 3368 1236
rect 3362 1231 3363 1235
rect 3367 1231 3368 1235
rect 3798 1232 3799 1236
rect 3803 1232 3804 1236
rect 3798 1231 3804 1232
rect 3362 1230 3368 1231
rect 3118 1220 3124 1221
rect 1974 1219 1980 1220
rect 1974 1215 1975 1219
rect 1979 1215 1980 1219
rect 3118 1216 3119 1220
rect 3123 1216 3124 1220
rect 3118 1215 3124 1216
rect 3254 1220 3260 1221
rect 3254 1216 3255 1220
rect 3259 1216 3260 1220
rect 3254 1215 3260 1216
rect 3390 1220 3396 1221
rect 3390 1216 3391 1220
rect 3395 1216 3396 1220
rect 3390 1215 3396 1216
rect 3798 1219 3804 1220
rect 3798 1215 3799 1219
rect 3803 1215 3804 1219
rect 1974 1214 1980 1215
rect 111 1198 115 1199
rect 111 1193 115 1194
rect 235 1198 239 1199
rect 235 1193 239 1194
rect 339 1198 343 1199
rect 339 1193 343 1194
rect 379 1198 383 1199
rect 379 1193 383 1194
rect 523 1198 527 1199
rect 523 1193 527 1194
rect 667 1198 671 1199
rect 667 1193 671 1194
rect 699 1198 703 1199
rect 699 1193 703 1194
rect 811 1198 815 1199
rect 811 1193 815 1194
rect 867 1198 871 1199
rect 867 1193 871 1194
rect 947 1198 951 1199
rect 947 1193 951 1194
rect 1035 1198 1039 1199
rect 1035 1193 1039 1194
rect 1091 1198 1095 1199
rect 1091 1193 1095 1194
rect 1195 1198 1199 1199
rect 1195 1193 1199 1194
rect 1235 1198 1239 1199
rect 1235 1193 1239 1194
rect 1347 1198 1351 1199
rect 1347 1193 1351 1194
rect 1379 1198 1383 1199
rect 1379 1193 1383 1194
rect 1499 1198 1503 1199
rect 1499 1193 1503 1194
rect 1515 1198 1519 1199
rect 1515 1193 1519 1194
rect 1651 1198 1655 1199
rect 1651 1193 1655 1194
rect 1787 1198 1791 1199
rect 1787 1193 1791 1194
rect 1935 1198 1939 1199
rect 1935 1193 1939 1194
rect 112 1133 114 1193
rect 110 1132 116 1133
rect 236 1132 238 1193
rect 380 1132 382 1193
rect 524 1132 526 1193
rect 668 1132 670 1193
rect 812 1132 814 1193
rect 948 1132 950 1193
rect 1092 1132 1094 1193
rect 1236 1132 1238 1193
rect 1380 1132 1382 1193
rect 1516 1132 1518 1193
rect 1652 1132 1654 1193
rect 1788 1132 1790 1193
rect 1936 1133 1938 1193
rect 1976 1191 1978 1214
rect 3120 1191 3122 1215
rect 3256 1191 3258 1215
rect 3392 1191 3394 1215
rect 3798 1214 3804 1215
rect 3800 1191 3802 1214
rect 3840 1203 3842 1271
rect 3860 1203 3862 1272
rect 4020 1203 4022 1272
rect 4212 1203 4214 1272
rect 4428 1203 4430 1272
rect 4668 1203 4670 1272
rect 4924 1203 4926 1272
rect 5196 1203 5198 1272
rect 5468 1203 5470 1272
rect 5662 1271 5668 1272
rect 5664 1203 5666 1271
rect 3839 1202 3843 1203
rect 3839 1197 3843 1198
rect 3859 1202 3863 1203
rect 3859 1197 3863 1198
rect 4019 1202 4023 1203
rect 4019 1197 4023 1198
rect 4091 1202 4095 1203
rect 4091 1197 4095 1198
rect 4211 1202 4215 1203
rect 4211 1197 4215 1198
rect 4339 1202 4343 1203
rect 4339 1197 4343 1198
rect 4427 1202 4431 1203
rect 4427 1197 4431 1198
rect 4579 1202 4583 1203
rect 4579 1197 4583 1198
rect 4667 1202 4671 1203
rect 4667 1197 4671 1198
rect 4811 1202 4815 1203
rect 4811 1197 4815 1198
rect 4923 1202 4927 1203
rect 4923 1197 4927 1198
rect 5043 1202 5047 1203
rect 5043 1197 5047 1198
rect 5195 1202 5199 1203
rect 5195 1197 5199 1198
rect 5275 1202 5279 1203
rect 5275 1197 5279 1198
rect 5467 1202 5471 1203
rect 5467 1197 5471 1198
rect 5515 1202 5519 1203
rect 5515 1197 5519 1198
rect 5663 1202 5667 1203
rect 5663 1197 5667 1198
rect 1975 1190 1979 1191
rect 1975 1185 1979 1186
rect 2983 1190 2987 1191
rect 2983 1185 2987 1186
rect 3119 1190 3123 1191
rect 3119 1185 3123 1186
rect 3255 1190 3259 1191
rect 3255 1185 3259 1186
rect 3391 1190 3395 1191
rect 3391 1185 3395 1186
rect 3799 1190 3803 1191
rect 3799 1185 3803 1186
rect 1976 1162 1978 1185
rect 1974 1161 1980 1162
rect 2984 1161 2986 1185
rect 3120 1161 3122 1185
rect 3256 1161 3258 1185
rect 3800 1162 3802 1185
rect 3798 1161 3804 1162
rect 1974 1157 1975 1161
rect 1979 1157 1980 1161
rect 1974 1156 1980 1157
rect 2982 1160 2988 1161
rect 2982 1156 2983 1160
rect 2987 1156 2988 1160
rect 2982 1155 2988 1156
rect 3118 1160 3124 1161
rect 3118 1156 3119 1160
rect 3123 1156 3124 1160
rect 3118 1155 3124 1156
rect 3254 1160 3260 1161
rect 3254 1156 3255 1160
rect 3259 1156 3260 1160
rect 3798 1157 3799 1161
rect 3803 1157 3804 1161
rect 3798 1156 3804 1157
rect 3254 1155 3260 1156
rect 2954 1145 2960 1146
rect 1974 1144 1980 1145
rect 1974 1140 1975 1144
rect 1979 1140 1980 1144
rect 2954 1141 2955 1145
rect 2959 1141 2960 1145
rect 2954 1140 2960 1141
rect 3090 1145 3096 1146
rect 3090 1141 3091 1145
rect 3095 1141 3096 1145
rect 3090 1140 3096 1141
rect 3226 1145 3232 1146
rect 3226 1141 3227 1145
rect 3231 1141 3232 1145
rect 3226 1140 3232 1141
rect 3798 1144 3804 1145
rect 3798 1140 3799 1144
rect 3803 1140 3804 1144
rect 1974 1139 1980 1140
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 234 1131 240 1132
rect 234 1127 235 1131
rect 239 1127 240 1131
rect 234 1126 240 1127
rect 378 1131 384 1132
rect 378 1127 379 1131
rect 383 1127 384 1131
rect 378 1126 384 1127
rect 522 1131 528 1132
rect 522 1127 523 1131
rect 527 1127 528 1131
rect 522 1126 528 1127
rect 666 1131 672 1132
rect 666 1127 667 1131
rect 671 1127 672 1131
rect 666 1126 672 1127
rect 810 1131 816 1132
rect 810 1127 811 1131
rect 815 1127 816 1131
rect 810 1126 816 1127
rect 946 1131 952 1132
rect 946 1127 947 1131
rect 951 1127 952 1131
rect 946 1126 952 1127
rect 1090 1131 1096 1132
rect 1090 1127 1091 1131
rect 1095 1127 1096 1131
rect 1090 1126 1096 1127
rect 1234 1131 1240 1132
rect 1234 1127 1235 1131
rect 1239 1127 1240 1131
rect 1234 1126 1240 1127
rect 1378 1131 1384 1132
rect 1378 1127 1379 1131
rect 1383 1127 1384 1131
rect 1378 1126 1384 1127
rect 1514 1131 1520 1132
rect 1514 1127 1515 1131
rect 1519 1127 1520 1131
rect 1514 1126 1520 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 262 1116 268 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 262 1112 263 1116
rect 267 1112 268 1116
rect 262 1111 268 1112
rect 406 1116 412 1117
rect 406 1112 407 1116
rect 411 1112 412 1116
rect 406 1111 412 1112
rect 550 1116 556 1117
rect 550 1112 551 1116
rect 555 1112 556 1116
rect 550 1111 556 1112
rect 694 1116 700 1117
rect 694 1112 695 1116
rect 699 1112 700 1116
rect 694 1111 700 1112
rect 838 1116 844 1117
rect 838 1112 839 1116
rect 843 1112 844 1116
rect 838 1111 844 1112
rect 974 1116 980 1117
rect 974 1112 975 1116
rect 979 1112 980 1116
rect 974 1111 980 1112
rect 1118 1116 1124 1117
rect 1118 1112 1119 1116
rect 1123 1112 1124 1116
rect 1118 1111 1124 1112
rect 1262 1116 1268 1117
rect 1262 1112 1263 1116
rect 1267 1112 1268 1116
rect 1262 1111 1268 1112
rect 1406 1116 1412 1117
rect 1406 1112 1407 1116
rect 1411 1112 1412 1116
rect 1406 1111 1412 1112
rect 1542 1116 1548 1117
rect 1542 1112 1543 1116
rect 1547 1112 1548 1116
rect 1542 1111 1548 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 110 1110 116 1111
rect 112 1075 114 1110
rect 264 1075 266 1111
rect 408 1075 410 1111
rect 552 1075 554 1111
rect 696 1075 698 1111
rect 840 1075 842 1111
rect 976 1075 978 1111
rect 1120 1075 1122 1111
rect 1264 1075 1266 1111
rect 1408 1075 1410 1111
rect 1544 1075 1546 1111
rect 1680 1075 1682 1111
rect 1816 1075 1818 1111
rect 1934 1110 1940 1111
rect 1936 1075 1938 1110
rect 1976 1079 1978 1139
rect 2956 1079 2958 1140
rect 3092 1079 3094 1140
rect 3228 1079 3230 1140
rect 3798 1139 3804 1140
rect 3800 1079 3802 1139
rect 3840 1137 3842 1197
rect 3838 1136 3844 1137
rect 3860 1136 3862 1197
rect 4092 1136 4094 1197
rect 4340 1136 4342 1197
rect 4580 1136 4582 1197
rect 4812 1136 4814 1197
rect 5044 1136 5046 1197
rect 5276 1136 5278 1197
rect 5516 1136 5518 1197
rect 5664 1137 5666 1197
rect 5662 1136 5668 1137
rect 3838 1132 3839 1136
rect 3843 1132 3844 1136
rect 3838 1131 3844 1132
rect 3858 1135 3864 1136
rect 3858 1131 3859 1135
rect 3863 1131 3864 1135
rect 3858 1130 3864 1131
rect 4090 1135 4096 1136
rect 4090 1131 4091 1135
rect 4095 1131 4096 1135
rect 4090 1130 4096 1131
rect 4338 1135 4344 1136
rect 4338 1131 4339 1135
rect 4343 1131 4344 1135
rect 4338 1130 4344 1131
rect 4578 1135 4584 1136
rect 4578 1131 4579 1135
rect 4583 1131 4584 1135
rect 4578 1130 4584 1131
rect 4810 1135 4816 1136
rect 4810 1131 4811 1135
rect 4815 1131 4816 1135
rect 4810 1130 4816 1131
rect 5042 1135 5048 1136
rect 5042 1131 5043 1135
rect 5047 1131 5048 1135
rect 5042 1130 5048 1131
rect 5274 1135 5280 1136
rect 5274 1131 5275 1135
rect 5279 1131 5280 1135
rect 5274 1130 5280 1131
rect 5514 1135 5520 1136
rect 5514 1131 5515 1135
rect 5519 1131 5520 1135
rect 5662 1132 5663 1136
rect 5667 1132 5668 1136
rect 5662 1131 5668 1132
rect 5514 1130 5520 1131
rect 3886 1120 3892 1121
rect 3838 1119 3844 1120
rect 3838 1115 3839 1119
rect 3843 1115 3844 1119
rect 3886 1116 3887 1120
rect 3891 1116 3892 1120
rect 3886 1115 3892 1116
rect 4118 1120 4124 1121
rect 4118 1116 4119 1120
rect 4123 1116 4124 1120
rect 4118 1115 4124 1116
rect 4366 1120 4372 1121
rect 4366 1116 4367 1120
rect 4371 1116 4372 1120
rect 4366 1115 4372 1116
rect 4606 1120 4612 1121
rect 4606 1116 4607 1120
rect 4611 1116 4612 1120
rect 4606 1115 4612 1116
rect 4838 1120 4844 1121
rect 4838 1116 4839 1120
rect 4843 1116 4844 1120
rect 4838 1115 4844 1116
rect 5070 1120 5076 1121
rect 5070 1116 5071 1120
rect 5075 1116 5076 1120
rect 5070 1115 5076 1116
rect 5302 1120 5308 1121
rect 5302 1116 5303 1120
rect 5307 1116 5308 1120
rect 5302 1115 5308 1116
rect 5542 1120 5548 1121
rect 5542 1116 5543 1120
rect 5547 1116 5548 1120
rect 5542 1115 5548 1116
rect 5662 1119 5668 1120
rect 5662 1115 5663 1119
rect 5667 1115 5668 1119
rect 3838 1114 3844 1115
rect 1975 1078 1979 1079
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 263 1074 267 1075
rect 263 1069 267 1070
rect 407 1074 411 1075
rect 407 1069 411 1070
rect 463 1074 467 1075
rect 463 1069 467 1070
rect 551 1074 555 1075
rect 551 1069 555 1070
rect 663 1074 667 1075
rect 663 1069 667 1070
rect 695 1074 699 1075
rect 695 1069 699 1070
rect 839 1074 843 1075
rect 839 1069 843 1070
rect 871 1074 875 1075
rect 871 1069 875 1070
rect 975 1074 979 1075
rect 975 1069 979 1070
rect 1079 1074 1083 1075
rect 1079 1069 1083 1070
rect 1119 1074 1123 1075
rect 1119 1069 1123 1070
rect 1263 1074 1267 1075
rect 1263 1069 1267 1070
rect 1407 1074 1411 1075
rect 1407 1069 1411 1070
rect 1543 1074 1547 1075
rect 1543 1069 1547 1070
rect 1679 1074 1683 1075
rect 1679 1069 1683 1070
rect 1815 1074 1819 1075
rect 1815 1069 1819 1070
rect 1935 1074 1939 1075
rect 1975 1073 1979 1074
rect 1995 1078 1999 1079
rect 1995 1073 1999 1074
rect 2131 1078 2135 1079
rect 2131 1073 2135 1074
rect 2275 1078 2279 1079
rect 2275 1073 2279 1074
rect 2443 1078 2447 1079
rect 2443 1073 2447 1074
rect 2627 1078 2631 1079
rect 2627 1073 2631 1074
rect 2819 1078 2823 1079
rect 2819 1073 2823 1074
rect 2955 1078 2959 1079
rect 2955 1073 2959 1074
rect 3027 1078 3031 1079
rect 3027 1073 3031 1074
rect 3091 1078 3095 1079
rect 3091 1073 3095 1074
rect 3227 1078 3231 1079
rect 3227 1073 3231 1074
rect 3235 1078 3239 1079
rect 3235 1073 3239 1074
rect 3451 1078 3455 1079
rect 3451 1073 3455 1074
rect 3651 1078 3655 1079
rect 3651 1073 3655 1074
rect 3799 1078 3803 1079
rect 3799 1073 3803 1074
rect 1935 1069 1939 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 264 1045 266 1069
rect 464 1045 466 1069
rect 664 1045 666 1069
rect 872 1045 874 1069
rect 1080 1045 1082 1069
rect 1936 1046 1938 1069
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 262 1044 268 1045
rect 262 1040 263 1044
rect 267 1040 268 1044
rect 262 1039 268 1040
rect 462 1044 468 1045
rect 462 1040 463 1044
rect 467 1040 468 1044
rect 462 1039 468 1040
rect 662 1044 668 1045
rect 662 1040 663 1044
rect 667 1040 668 1044
rect 662 1039 668 1040
rect 870 1044 876 1045
rect 870 1040 871 1044
rect 875 1040 876 1044
rect 870 1039 876 1040
rect 1078 1044 1084 1045
rect 1078 1040 1079 1044
rect 1083 1040 1084 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1078 1039 1084 1040
rect 234 1029 240 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 234 1025 235 1029
rect 239 1025 240 1029
rect 234 1024 240 1025
rect 434 1029 440 1030
rect 434 1025 435 1029
rect 439 1025 440 1029
rect 434 1024 440 1025
rect 634 1029 640 1030
rect 634 1025 635 1029
rect 639 1025 640 1029
rect 634 1024 640 1025
rect 842 1029 848 1030
rect 842 1025 843 1029
rect 847 1025 848 1029
rect 842 1024 848 1025
rect 1050 1029 1056 1030
rect 1050 1025 1051 1029
rect 1055 1025 1056 1029
rect 1050 1024 1056 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 112 951 114 1023
rect 236 951 238 1024
rect 436 951 438 1024
rect 636 951 638 1024
rect 844 951 846 1024
rect 1052 951 1054 1024
rect 1934 1023 1940 1024
rect 1936 951 1938 1023
rect 1976 1013 1978 1073
rect 1974 1012 1980 1013
rect 1996 1012 1998 1073
rect 2132 1012 2134 1073
rect 2276 1012 2278 1073
rect 2444 1012 2446 1073
rect 2628 1012 2630 1073
rect 2820 1012 2822 1073
rect 3028 1012 3030 1073
rect 3236 1012 3238 1073
rect 3452 1012 3454 1073
rect 3652 1012 3654 1073
rect 3800 1013 3802 1073
rect 3840 1071 3842 1114
rect 3888 1071 3890 1115
rect 4120 1071 4122 1115
rect 4368 1071 4370 1115
rect 4608 1071 4610 1115
rect 4840 1071 4842 1115
rect 5072 1071 5074 1115
rect 5304 1071 5306 1115
rect 5544 1071 5546 1115
rect 5662 1114 5668 1115
rect 5664 1071 5666 1114
rect 3839 1070 3843 1071
rect 3839 1065 3843 1066
rect 3887 1070 3891 1071
rect 3887 1065 3891 1066
rect 4119 1070 4123 1071
rect 4119 1065 4123 1066
rect 4367 1070 4371 1071
rect 4367 1065 4371 1066
rect 4607 1070 4611 1071
rect 4607 1065 4611 1066
rect 4839 1070 4843 1071
rect 4839 1065 4843 1066
rect 4863 1070 4867 1071
rect 4863 1065 4867 1066
rect 4999 1070 5003 1071
rect 4999 1065 5003 1066
rect 5071 1070 5075 1071
rect 5071 1065 5075 1066
rect 5135 1070 5139 1071
rect 5135 1065 5139 1066
rect 5271 1070 5275 1071
rect 5271 1065 5275 1066
rect 5303 1070 5307 1071
rect 5303 1065 5307 1066
rect 5407 1070 5411 1071
rect 5407 1065 5411 1066
rect 5543 1070 5547 1071
rect 5543 1065 5547 1066
rect 5663 1070 5667 1071
rect 5663 1065 5667 1066
rect 3840 1042 3842 1065
rect 3838 1041 3844 1042
rect 4864 1041 4866 1065
rect 5000 1041 5002 1065
rect 5136 1041 5138 1065
rect 5272 1041 5274 1065
rect 5408 1041 5410 1065
rect 5544 1041 5546 1065
rect 5664 1042 5666 1065
rect 5662 1041 5668 1042
rect 3838 1037 3839 1041
rect 3843 1037 3844 1041
rect 3838 1036 3844 1037
rect 4862 1040 4868 1041
rect 4862 1036 4863 1040
rect 4867 1036 4868 1040
rect 4862 1035 4868 1036
rect 4998 1040 5004 1041
rect 4998 1036 4999 1040
rect 5003 1036 5004 1040
rect 4998 1035 5004 1036
rect 5134 1040 5140 1041
rect 5134 1036 5135 1040
rect 5139 1036 5140 1040
rect 5134 1035 5140 1036
rect 5270 1040 5276 1041
rect 5270 1036 5271 1040
rect 5275 1036 5276 1040
rect 5270 1035 5276 1036
rect 5406 1040 5412 1041
rect 5406 1036 5407 1040
rect 5411 1036 5412 1040
rect 5406 1035 5412 1036
rect 5542 1040 5548 1041
rect 5542 1036 5543 1040
rect 5547 1036 5548 1040
rect 5662 1037 5663 1041
rect 5667 1037 5668 1041
rect 5662 1036 5668 1037
rect 5542 1035 5548 1036
rect 4834 1025 4840 1026
rect 3838 1024 3844 1025
rect 3838 1020 3839 1024
rect 3843 1020 3844 1024
rect 4834 1021 4835 1025
rect 4839 1021 4840 1025
rect 4834 1020 4840 1021
rect 4970 1025 4976 1026
rect 4970 1021 4971 1025
rect 4975 1021 4976 1025
rect 4970 1020 4976 1021
rect 5106 1025 5112 1026
rect 5106 1021 5107 1025
rect 5111 1021 5112 1025
rect 5106 1020 5112 1021
rect 5242 1025 5248 1026
rect 5242 1021 5243 1025
rect 5247 1021 5248 1025
rect 5242 1020 5248 1021
rect 5378 1025 5384 1026
rect 5378 1021 5379 1025
rect 5383 1021 5384 1025
rect 5378 1020 5384 1021
rect 5514 1025 5520 1026
rect 5514 1021 5515 1025
rect 5519 1021 5520 1025
rect 5514 1020 5520 1021
rect 5662 1024 5668 1025
rect 5662 1020 5663 1024
rect 5667 1020 5668 1024
rect 3838 1019 3844 1020
rect 3798 1012 3804 1013
rect 1974 1008 1975 1012
rect 1979 1008 1980 1012
rect 1974 1007 1980 1008
rect 1994 1011 2000 1012
rect 1994 1007 1995 1011
rect 1999 1007 2000 1011
rect 1994 1006 2000 1007
rect 2130 1011 2136 1012
rect 2130 1007 2131 1011
rect 2135 1007 2136 1011
rect 2130 1006 2136 1007
rect 2274 1011 2280 1012
rect 2274 1007 2275 1011
rect 2279 1007 2280 1011
rect 2274 1006 2280 1007
rect 2442 1011 2448 1012
rect 2442 1007 2443 1011
rect 2447 1007 2448 1011
rect 2442 1006 2448 1007
rect 2626 1011 2632 1012
rect 2626 1007 2627 1011
rect 2631 1007 2632 1011
rect 2626 1006 2632 1007
rect 2818 1011 2824 1012
rect 2818 1007 2819 1011
rect 2823 1007 2824 1011
rect 2818 1006 2824 1007
rect 3026 1011 3032 1012
rect 3026 1007 3027 1011
rect 3031 1007 3032 1011
rect 3026 1006 3032 1007
rect 3234 1011 3240 1012
rect 3234 1007 3235 1011
rect 3239 1007 3240 1011
rect 3234 1006 3240 1007
rect 3450 1011 3456 1012
rect 3450 1007 3451 1011
rect 3455 1007 3456 1011
rect 3450 1006 3456 1007
rect 3650 1011 3656 1012
rect 3650 1007 3651 1011
rect 3655 1007 3656 1011
rect 3798 1008 3799 1012
rect 3803 1008 3804 1012
rect 3798 1007 3804 1008
rect 3650 1006 3656 1007
rect 2022 996 2028 997
rect 1974 995 1980 996
rect 1974 991 1975 995
rect 1979 991 1980 995
rect 2022 992 2023 996
rect 2027 992 2028 996
rect 2022 991 2028 992
rect 2158 996 2164 997
rect 2158 992 2159 996
rect 2163 992 2164 996
rect 2158 991 2164 992
rect 2302 996 2308 997
rect 2302 992 2303 996
rect 2307 992 2308 996
rect 2302 991 2308 992
rect 2470 996 2476 997
rect 2470 992 2471 996
rect 2475 992 2476 996
rect 2470 991 2476 992
rect 2654 996 2660 997
rect 2654 992 2655 996
rect 2659 992 2660 996
rect 2654 991 2660 992
rect 2846 996 2852 997
rect 2846 992 2847 996
rect 2851 992 2852 996
rect 2846 991 2852 992
rect 3054 996 3060 997
rect 3054 992 3055 996
rect 3059 992 3060 996
rect 3054 991 3060 992
rect 3262 996 3268 997
rect 3262 992 3263 996
rect 3267 992 3268 996
rect 3262 991 3268 992
rect 3478 996 3484 997
rect 3478 992 3479 996
rect 3483 992 3484 996
rect 3478 991 3484 992
rect 3678 996 3684 997
rect 3678 992 3679 996
rect 3683 992 3684 996
rect 3678 991 3684 992
rect 3798 995 3804 996
rect 3798 991 3799 995
rect 3803 991 3804 995
rect 1974 990 1980 991
rect 1976 967 1978 990
rect 2024 967 2026 991
rect 2160 967 2162 991
rect 2304 967 2306 991
rect 2472 967 2474 991
rect 2656 967 2658 991
rect 2848 967 2850 991
rect 3056 967 3058 991
rect 3264 967 3266 991
rect 3480 967 3482 991
rect 3680 967 3682 991
rect 3798 990 3804 991
rect 3800 967 3802 990
rect 1975 966 1979 967
rect 1975 961 1979 962
rect 2023 966 2027 967
rect 2023 961 2027 962
rect 2095 966 2099 967
rect 2095 961 2099 962
rect 2159 966 2163 967
rect 2159 961 2163 962
rect 2231 966 2235 967
rect 2231 961 2235 962
rect 2303 966 2307 967
rect 2303 961 2307 962
rect 2367 966 2371 967
rect 2367 961 2371 962
rect 2471 966 2475 967
rect 2471 961 2475 962
rect 2503 966 2507 967
rect 2503 961 2507 962
rect 2655 966 2659 967
rect 2655 961 2659 962
rect 2831 966 2835 967
rect 2831 961 2835 962
rect 2847 966 2851 967
rect 2847 961 2851 962
rect 3023 966 3027 967
rect 3023 961 3027 962
rect 3055 966 3059 967
rect 3055 961 3059 962
rect 3231 966 3235 967
rect 3231 961 3235 962
rect 3263 966 3267 967
rect 3263 961 3267 962
rect 3455 966 3459 967
rect 3455 961 3459 962
rect 3479 966 3483 967
rect 3479 961 3483 962
rect 3679 966 3683 967
rect 3679 961 3683 962
rect 3799 966 3803 967
rect 3799 961 3803 962
rect 111 950 115 951
rect 111 945 115 946
rect 195 950 199 951
rect 195 945 199 946
rect 235 950 239 951
rect 235 945 239 946
rect 371 950 375 951
rect 371 945 375 946
rect 435 950 439 951
rect 435 945 439 946
rect 547 950 551 951
rect 547 945 551 946
rect 635 950 639 951
rect 635 945 639 946
rect 723 950 727 951
rect 723 945 727 946
rect 843 950 847 951
rect 843 945 847 946
rect 907 950 911 951
rect 907 945 911 946
rect 1051 950 1055 951
rect 1051 945 1055 946
rect 1091 950 1095 951
rect 1091 945 1095 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 112 885 114 945
rect 110 884 116 885
rect 196 884 198 945
rect 372 884 374 945
rect 548 884 550 945
rect 724 884 726 945
rect 908 884 910 945
rect 1092 884 1094 945
rect 1936 885 1938 945
rect 1976 938 1978 961
rect 1974 937 1980 938
rect 2096 937 2098 961
rect 2232 937 2234 961
rect 2368 937 2370 961
rect 2504 937 2506 961
rect 2656 937 2658 961
rect 2832 937 2834 961
rect 3024 937 3026 961
rect 3232 937 3234 961
rect 3456 937 3458 961
rect 3680 937 3682 961
rect 3800 938 3802 961
rect 3840 947 3842 1019
rect 4836 947 4838 1020
rect 4972 947 4974 1020
rect 5108 947 5110 1020
rect 5244 947 5246 1020
rect 5380 947 5382 1020
rect 5516 947 5518 1020
rect 5662 1019 5668 1020
rect 5664 947 5666 1019
rect 3839 946 3843 947
rect 3839 941 3843 942
rect 4587 946 4591 947
rect 4587 941 4591 942
rect 4755 946 4759 947
rect 4755 941 4759 942
rect 4835 946 4839 947
rect 4835 941 4839 942
rect 4939 946 4943 947
rect 4939 941 4943 942
rect 4971 946 4975 947
rect 4971 941 4975 942
rect 5107 946 5111 947
rect 5107 941 5111 942
rect 5131 946 5135 947
rect 5131 941 5135 942
rect 5243 946 5247 947
rect 5243 941 5247 942
rect 5331 946 5335 947
rect 5331 941 5335 942
rect 5379 946 5383 947
rect 5379 941 5383 942
rect 5515 946 5519 947
rect 5515 941 5519 942
rect 5663 946 5667 947
rect 5663 941 5667 942
rect 3798 937 3804 938
rect 1974 933 1975 937
rect 1979 933 1980 937
rect 1974 932 1980 933
rect 2094 936 2100 937
rect 2094 932 2095 936
rect 2099 932 2100 936
rect 2094 931 2100 932
rect 2230 936 2236 937
rect 2230 932 2231 936
rect 2235 932 2236 936
rect 2230 931 2236 932
rect 2366 936 2372 937
rect 2366 932 2367 936
rect 2371 932 2372 936
rect 2366 931 2372 932
rect 2502 936 2508 937
rect 2502 932 2503 936
rect 2507 932 2508 936
rect 2502 931 2508 932
rect 2654 936 2660 937
rect 2654 932 2655 936
rect 2659 932 2660 936
rect 2654 931 2660 932
rect 2830 936 2836 937
rect 2830 932 2831 936
rect 2835 932 2836 936
rect 2830 931 2836 932
rect 3022 936 3028 937
rect 3022 932 3023 936
rect 3027 932 3028 936
rect 3022 931 3028 932
rect 3230 936 3236 937
rect 3230 932 3231 936
rect 3235 932 3236 936
rect 3230 931 3236 932
rect 3454 936 3460 937
rect 3454 932 3455 936
rect 3459 932 3460 936
rect 3454 931 3460 932
rect 3678 936 3684 937
rect 3678 932 3679 936
rect 3683 932 3684 936
rect 3798 933 3799 937
rect 3803 933 3804 937
rect 3798 932 3804 933
rect 3678 931 3684 932
rect 2066 921 2072 922
rect 1974 920 1980 921
rect 1974 916 1975 920
rect 1979 916 1980 920
rect 2066 917 2067 921
rect 2071 917 2072 921
rect 2066 916 2072 917
rect 2202 921 2208 922
rect 2202 917 2203 921
rect 2207 917 2208 921
rect 2202 916 2208 917
rect 2338 921 2344 922
rect 2338 917 2339 921
rect 2343 917 2344 921
rect 2338 916 2344 917
rect 2474 921 2480 922
rect 2474 917 2475 921
rect 2479 917 2480 921
rect 2474 916 2480 917
rect 2626 921 2632 922
rect 2626 917 2627 921
rect 2631 917 2632 921
rect 2626 916 2632 917
rect 2802 921 2808 922
rect 2802 917 2803 921
rect 2807 917 2808 921
rect 2802 916 2808 917
rect 2994 921 3000 922
rect 2994 917 2995 921
rect 2999 917 3000 921
rect 2994 916 3000 917
rect 3202 921 3208 922
rect 3202 917 3203 921
rect 3207 917 3208 921
rect 3202 916 3208 917
rect 3426 921 3432 922
rect 3426 917 3427 921
rect 3431 917 3432 921
rect 3426 916 3432 917
rect 3650 921 3656 922
rect 3650 917 3651 921
rect 3655 917 3656 921
rect 3650 916 3656 917
rect 3798 920 3804 921
rect 3798 916 3799 920
rect 3803 916 3804 920
rect 1974 915 1980 916
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 194 883 200 884
rect 194 879 195 883
rect 199 879 200 883
rect 194 878 200 879
rect 370 883 376 884
rect 370 879 371 883
rect 375 879 376 883
rect 370 878 376 879
rect 546 883 552 884
rect 546 879 547 883
rect 551 879 552 883
rect 546 878 552 879
rect 722 883 728 884
rect 722 879 723 883
rect 727 879 728 883
rect 722 878 728 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1090 883 1096 884
rect 1090 879 1091 883
rect 1095 879 1096 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1090 878 1096 879
rect 222 868 228 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 222 864 223 868
rect 227 864 228 868
rect 222 863 228 864
rect 398 868 404 869
rect 398 864 399 868
rect 403 864 404 868
rect 398 863 404 864
rect 574 868 580 869
rect 574 864 575 868
rect 579 864 580 868
rect 574 863 580 864
rect 750 868 756 869
rect 750 864 751 868
rect 755 864 756 868
rect 750 863 756 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1118 868 1124 869
rect 1118 864 1119 868
rect 1123 864 1124 868
rect 1118 863 1124 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 110 862 116 863
rect 112 823 114 862
rect 224 823 226 863
rect 400 823 402 863
rect 576 823 578 863
rect 752 823 754 863
rect 936 823 938 863
rect 1120 823 1122 863
rect 1934 862 1940 863
rect 1936 823 1938 862
rect 1976 855 1978 915
rect 2068 855 2070 916
rect 2204 855 2206 916
rect 2340 855 2342 916
rect 2476 855 2478 916
rect 2628 855 2630 916
rect 2804 855 2806 916
rect 2996 855 2998 916
rect 3204 855 3206 916
rect 3428 855 3430 916
rect 3652 855 3654 916
rect 3798 915 3804 916
rect 3800 855 3802 915
rect 3840 881 3842 941
rect 3838 880 3844 881
rect 4588 880 4590 941
rect 4756 880 4758 941
rect 4940 880 4942 941
rect 5132 880 5134 941
rect 5332 880 5334 941
rect 5516 880 5518 941
rect 5664 881 5666 941
rect 5662 880 5668 881
rect 3838 876 3839 880
rect 3843 876 3844 880
rect 3838 875 3844 876
rect 4586 879 4592 880
rect 4586 875 4587 879
rect 4591 875 4592 879
rect 4586 874 4592 875
rect 4754 879 4760 880
rect 4754 875 4755 879
rect 4759 875 4760 879
rect 4754 874 4760 875
rect 4938 879 4944 880
rect 4938 875 4939 879
rect 4943 875 4944 879
rect 4938 874 4944 875
rect 5130 879 5136 880
rect 5130 875 5131 879
rect 5135 875 5136 879
rect 5130 874 5136 875
rect 5330 879 5336 880
rect 5330 875 5331 879
rect 5335 875 5336 879
rect 5330 874 5336 875
rect 5514 879 5520 880
rect 5514 875 5515 879
rect 5519 875 5520 879
rect 5662 876 5663 880
rect 5667 876 5668 880
rect 5662 875 5668 876
rect 5514 874 5520 875
rect 4614 864 4620 865
rect 3838 863 3844 864
rect 3838 859 3839 863
rect 3843 859 3844 863
rect 4614 860 4615 864
rect 4619 860 4620 864
rect 4614 859 4620 860
rect 4782 864 4788 865
rect 4782 860 4783 864
rect 4787 860 4788 864
rect 4782 859 4788 860
rect 4966 864 4972 865
rect 4966 860 4967 864
rect 4971 860 4972 864
rect 4966 859 4972 860
rect 5158 864 5164 865
rect 5158 860 5159 864
rect 5163 860 5164 864
rect 5158 859 5164 860
rect 5358 864 5364 865
rect 5358 860 5359 864
rect 5363 860 5364 864
rect 5358 859 5364 860
rect 5542 864 5548 865
rect 5542 860 5543 864
rect 5547 860 5548 864
rect 5542 859 5548 860
rect 5662 863 5668 864
rect 5662 859 5663 863
rect 5667 859 5668 863
rect 3838 858 3844 859
rect 1975 854 1979 855
rect 1975 849 1979 850
rect 2067 854 2071 855
rect 2067 849 2071 850
rect 2203 854 2207 855
rect 2203 849 2207 850
rect 2307 854 2311 855
rect 2307 849 2311 850
rect 2339 854 2343 855
rect 2339 849 2343 850
rect 2475 854 2479 855
rect 2475 849 2479 850
rect 2483 854 2487 855
rect 2483 849 2487 850
rect 2627 854 2631 855
rect 2627 849 2631 850
rect 2659 854 2663 855
rect 2659 849 2663 850
rect 2803 854 2807 855
rect 2803 849 2807 850
rect 2827 854 2831 855
rect 2827 849 2831 850
rect 2995 854 2999 855
rect 2995 849 2999 850
rect 3163 854 3167 855
rect 3163 849 3167 850
rect 3203 854 3207 855
rect 3203 849 3207 850
rect 3331 854 3335 855
rect 3331 849 3335 850
rect 3427 854 3431 855
rect 3427 849 3431 850
rect 3499 854 3503 855
rect 3499 849 3503 850
rect 3651 854 3655 855
rect 3651 849 3655 850
rect 3799 854 3803 855
rect 3799 849 3803 850
rect 111 822 115 823
rect 111 817 115 818
rect 159 822 163 823
rect 159 817 163 818
rect 223 822 227 823
rect 223 817 227 818
rect 351 822 355 823
rect 351 817 355 818
rect 399 822 403 823
rect 399 817 403 818
rect 575 822 579 823
rect 575 817 579 818
rect 583 822 587 823
rect 583 817 587 818
rect 751 822 755 823
rect 751 817 755 818
rect 839 822 843 823
rect 839 817 843 818
rect 935 822 939 823
rect 935 817 939 818
rect 1111 822 1115 823
rect 1111 817 1115 818
rect 1119 822 1123 823
rect 1119 817 1123 818
rect 1399 822 1403 823
rect 1399 817 1403 818
rect 1687 822 1691 823
rect 1687 817 1691 818
rect 1935 822 1939 823
rect 1935 817 1939 818
rect 112 794 114 817
rect 110 793 116 794
rect 160 793 162 817
rect 352 793 354 817
rect 584 793 586 817
rect 840 793 842 817
rect 1112 793 1114 817
rect 1400 793 1402 817
rect 1688 793 1690 817
rect 1936 794 1938 817
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 158 792 164 793
rect 158 788 159 792
rect 163 788 164 792
rect 158 787 164 788
rect 350 792 356 793
rect 350 788 351 792
rect 355 788 356 792
rect 350 787 356 788
rect 582 792 588 793
rect 582 788 583 792
rect 587 788 588 792
rect 582 787 588 788
rect 838 792 844 793
rect 838 788 839 792
rect 843 788 844 792
rect 838 787 844 788
rect 1110 792 1116 793
rect 1110 788 1111 792
rect 1115 788 1116 792
rect 1110 787 1116 788
rect 1398 792 1404 793
rect 1398 788 1399 792
rect 1403 788 1404 792
rect 1398 787 1404 788
rect 1686 792 1692 793
rect 1686 788 1687 792
rect 1691 788 1692 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 1976 789 1978 849
rect 1934 788 1940 789
rect 1974 788 1980 789
rect 2308 788 2310 849
rect 2484 788 2486 849
rect 2660 788 2662 849
rect 2828 788 2830 849
rect 2996 788 2998 849
rect 3164 788 3166 849
rect 3332 788 3334 849
rect 3500 788 3502 849
rect 3652 788 3654 849
rect 3800 789 3802 849
rect 3840 827 3842 858
rect 4616 827 4618 859
rect 4784 827 4786 859
rect 4968 827 4970 859
rect 5160 827 5162 859
rect 5360 827 5362 859
rect 5544 827 5546 859
rect 5662 858 5668 859
rect 5664 827 5666 858
rect 3839 826 3843 827
rect 3839 821 3843 822
rect 3983 826 3987 827
rect 3983 821 3987 822
rect 4239 826 4243 827
rect 4239 821 4243 822
rect 4535 826 4539 827
rect 4535 821 4539 822
rect 4615 826 4619 827
rect 4615 821 4619 822
rect 4783 826 4787 827
rect 4783 821 4787 822
rect 4863 826 4867 827
rect 4863 821 4867 822
rect 4967 826 4971 827
rect 4967 821 4971 822
rect 5159 826 5163 827
rect 5159 821 5163 822
rect 5215 826 5219 827
rect 5215 821 5219 822
rect 5359 826 5363 827
rect 5359 821 5363 822
rect 5543 826 5547 827
rect 5543 821 5547 822
rect 5663 826 5667 827
rect 5663 821 5667 822
rect 3840 798 3842 821
rect 3838 797 3844 798
rect 3984 797 3986 821
rect 4240 797 4242 821
rect 4536 797 4538 821
rect 4864 797 4866 821
rect 5216 797 5218 821
rect 5544 797 5546 821
rect 5664 798 5666 821
rect 5662 797 5668 798
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3982 796 3988 797
rect 3982 792 3983 796
rect 3987 792 3988 796
rect 3982 791 3988 792
rect 4238 796 4244 797
rect 4238 792 4239 796
rect 4243 792 4244 796
rect 4238 791 4244 792
rect 4534 796 4540 797
rect 4534 792 4535 796
rect 4539 792 4540 796
rect 4534 791 4540 792
rect 4862 796 4868 797
rect 4862 792 4863 796
rect 4867 792 4868 796
rect 4862 791 4868 792
rect 5214 796 5220 797
rect 5214 792 5215 796
rect 5219 792 5220 796
rect 5214 791 5220 792
rect 5542 796 5548 797
rect 5542 792 5543 796
rect 5547 792 5548 796
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5542 791 5548 792
rect 3798 788 3804 789
rect 1686 787 1692 788
rect 1974 784 1975 788
rect 1979 784 1980 788
rect 1974 783 1980 784
rect 2306 787 2312 788
rect 2306 783 2307 787
rect 2311 783 2312 787
rect 2306 782 2312 783
rect 2482 787 2488 788
rect 2482 783 2483 787
rect 2487 783 2488 787
rect 2482 782 2488 783
rect 2658 787 2664 788
rect 2658 783 2659 787
rect 2663 783 2664 787
rect 2658 782 2664 783
rect 2826 787 2832 788
rect 2826 783 2827 787
rect 2831 783 2832 787
rect 2826 782 2832 783
rect 2994 787 3000 788
rect 2994 783 2995 787
rect 2999 783 3000 787
rect 2994 782 3000 783
rect 3162 787 3168 788
rect 3162 783 3163 787
rect 3167 783 3168 787
rect 3162 782 3168 783
rect 3330 787 3336 788
rect 3330 783 3331 787
rect 3335 783 3336 787
rect 3330 782 3336 783
rect 3498 787 3504 788
rect 3498 783 3499 787
rect 3503 783 3504 787
rect 3498 782 3504 783
rect 3650 787 3656 788
rect 3650 783 3651 787
rect 3655 783 3656 787
rect 3798 784 3799 788
rect 3803 784 3804 788
rect 3798 783 3804 784
rect 3650 782 3656 783
rect 3954 781 3960 782
rect 3838 780 3844 781
rect 130 777 136 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 130 773 131 777
rect 135 773 136 777
rect 130 772 136 773
rect 322 777 328 778
rect 322 773 323 777
rect 327 773 328 777
rect 322 772 328 773
rect 554 777 560 778
rect 554 773 555 777
rect 559 773 560 777
rect 554 772 560 773
rect 810 777 816 778
rect 810 773 811 777
rect 815 773 816 777
rect 810 772 816 773
rect 1082 777 1088 778
rect 1082 773 1083 777
rect 1087 773 1088 777
rect 1082 772 1088 773
rect 1370 777 1376 778
rect 1370 773 1371 777
rect 1375 773 1376 777
rect 1370 772 1376 773
rect 1658 777 1664 778
rect 1658 773 1659 777
rect 1663 773 1664 777
rect 1658 772 1664 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3954 777 3955 781
rect 3959 777 3960 781
rect 3954 776 3960 777
rect 4210 781 4216 782
rect 4210 777 4211 781
rect 4215 777 4216 781
rect 4210 776 4216 777
rect 4506 781 4512 782
rect 4506 777 4507 781
rect 4511 777 4512 781
rect 4506 776 4512 777
rect 4834 781 4840 782
rect 4834 777 4835 781
rect 4839 777 4840 781
rect 4834 776 4840 777
rect 5186 781 5192 782
rect 5186 777 5187 781
rect 5191 777 5192 781
rect 5186 776 5192 777
rect 5514 781 5520 782
rect 5514 777 5515 781
rect 5519 777 5520 781
rect 5514 776 5520 777
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 3838 775 3844 776
rect 2334 772 2340 773
rect 110 771 116 772
rect 112 711 114 771
rect 132 711 134 772
rect 324 711 326 772
rect 556 711 558 772
rect 812 711 814 772
rect 1084 711 1086 772
rect 1372 711 1374 772
rect 1660 711 1662 772
rect 1934 771 1940 772
rect 1974 771 1980 772
rect 1936 711 1938 771
rect 1974 767 1975 771
rect 1979 767 1980 771
rect 2334 768 2335 772
rect 2339 768 2340 772
rect 2334 767 2340 768
rect 2510 772 2516 773
rect 2510 768 2511 772
rect 2515 768 2516 772
rect 2510 767 2516 768
rect 2686 772 2692 773
rect 2686 768 2687 772
rect 2691 768 2692 772
rect 2686 767 2692 768
rect 2854 772 2860 773
rect 2854 768 2855 772
rect 2859 768 2860 772
rect 2854 767 2860 768
rect 3022 772 3028 773
rect 3022 768 3023 772
rect 3027 768 3028 772
rect 3022 767 3028 768
rect 3190 772 3196 773
rect 3190 768 3191 772
rect 3195 768 3196 772
rect 3190 767 3196 768
rect 3358 772 3364 773
rect 3358 768 3359 772
rect 3363 768 3364 772
rect 3358 767 3364 768
rect 3526 772 3532 773
rect 3526 768 3527 772
rect 3531 768 3532 772
rect 3526 767 3532 768
rect 3678 772 3684 773
rect 3678 768 3679 772
rect 3683 768 3684 772
rect 3678 767 3684 768
rect 3798 771 3804 772
rect 3798 767 3799 771
rect 3803 767 3804 771
rect 1974 766 1980 767
rect 1976 739 1978 766
rect 2336 739 2338 767
rect 2512 739 2514 767
rect 2688 739 2690 767
rect 2856 739 2858 767
rect 3024 739 3026 767
rect 3192 739 3194 767
rect 3360 739 3362 767
rect 3528 739 3530 767
rect 3680 739 3682 767
rect 3798 766 3804 767
rect 3800 739 3802 766
rect 1975 738 1979 739
rect 1975 733 1979 734
rect 2335 738 2339 739
rect 2335 733 2339 734
rect 2511 738 2515 739
rect 2511 733 2515 734
rect 2687 738 2691 739
rect 2687 733 2691 734
rect 2855 738 2859 739
rect 2855 733 2859 734
rect 3023 738 3027 739
rect 3023 733 3027 734
rect 3135 738 3139 739
rect 3135 733 3139 734
rect 3191 738 3195 739
rect 3191 733 3195 734
rect 3271 738 3275 739
rect 3271 733 3275 734
rect 3359 738 3363 739
rect 3359 733 3363 734
rect 3407 738 3411 739
rect 3407 733 3411 734
rect 3527 738 3531 739
rect 3527 733 3531 734
rect 3543 738 3547 739
rect 3543 733 3547 734
rect 3679 738 3683 739
rect 3679 733 3683 734
rect 3799 738 3803 739
rect 3799 733 3803 734
rect 111 710 115 711
rect 111 705 115 706
rect 131 710 135 711
rect 131 705 135 706
rect 291 710 295 711
rect 291 705 295 706
rect 323 710 327 711
rect 323 705 327 706
rect 483 710 487 711
rect 483 705 487 706
rect 555 710 559 711
rect 555 705 559 706
rect 675 710 679 711
rect 675 705 679 706
rect 811 710 815 711
rect 811 705 815 706
rect 867 710 871 711
rect 867 705 871 706
rect 1059 710 1063 711
rect 1059 705 1063 706
rect 1083 710 1087 711
rect 1083 705 1087 706
rect 1251 710 1255 711
rect 1251 705 1255 706
rect 1371 710 1375 711
rect 1371 705 1375 706
rect 1435 710 1439 711
rect 1435 705 1439 706
rect 1619 710 1623 711
rect 1619 705 1623 706
rect 1659 710 1663 711
rect 1659 705 1663 706
rect 1787 710 1791 711
rect 1787 705 1791 706
rect 1935 710 1939 711
rect 1976 710 1978 733
rect 1935 705 1939 706
rect 1974 709 1980 710
rect 3136 709 3138 733
rect 3272 709 3274 733
rect 3408 709 3410 733
rect 3544 709 3546 733
rect 3680 709 3682 733
rect 3800 710 3802 733
rect 3798 709 3804 710
rect 1974 705 1975 709
rect 1979 705 1980 709
rect 112 645 114 705
rect 110 644 116 645
rect 132 644 134 705
rect 292 644 294 705
rect 484 644 486 705
rect 676 644 678 705
rect 868 644 870 705
rect 1060 644 1062 705
rect 1252 644 1254 705
rect 1436 644 1438 705
rect 1620 644 1622 705
rect 1788 644 1790 705
rect 1936 645 1938 705
rect 1974 704 1980 705
rect 3134 708 3140 709
rect 3134 704 3135 708
rect 3139 704 3140 708
rect 3134 703 3140 704
rect 3270 708 3276 709
rect 3270 704 3271 708
rect 3275 704 3276 708
rect 3270 703 3276 704
rect 3406 708 3412 709
rect 3406 704 3407 708
rect 3411 704 3412 708
rect 3406 703 3412 704
rect 3542 708 3548 709
rect 3542 704 3543 708
rect 3547 704 3548 708
rect 3542 703 3548 704
rect 3678 708 3684 709
rect 3678 704 3679 708
rect 3683 704 3684 708
rect 3798 705 3799 709
rect 3803 705 3804 709
rect 3798 704 3804 705
rect 3678 703 3684 704
rect 3106 693 3112 694
rect 1974 692 1980 693
rect 1974 688 1975 692
rect 1979 688 1980 692
rect 3106 689 3107 693
rect 3111 689 3112 693
rect 3106 688 3112 689
rect 3242 693 3248 694
rect 3242 689 3243 693
rect 3247 689 3248 693
rect 3242 688 3248 689
rect 3378 693 3384 694
rect 3378 689 3379 693
rect 3383 689 3384 693
rect 3378 688 3384 689
rect 3514 693 3520 694
rect 3514 689 3515 693
rect 3519 689 3520 693
rect 3514 688 3520 689
rect 3650 693 3656 694
rect 3650 689 3651 693
rect 3655 689 3656 693
rect 3650 688 3656 689
rect 3798 692 3804 693
rect 3798 688 3799 692
rect 3803 688 3804 692
rect 3840 691 3842 775
rect 3956 691 3958 776
rect 4212 691 4214 776
rect 4508 691 4510 776
rect 4836 691 4838 776
rect 5188 691 5190 776
rect 5516 691 5518 776
rect 5662 775 5668 776
rect 5664 691 5666 775
rect 1974 687 1980 688
rect 1934 644 1940 645
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 290 643 296 644
rect 290 639 291 643
rect 295 639 296 643
rect 290 638 296 639
rect 482 643 488 644
rect 482 639 483 643
rect 487 639 488 643
rect 482 638 488 639
rect 674 643 680 644
rect 674 639 675 643
rect 679 639 680 643
rect 674 638 680 639
rect 866 643 872 644
rect 866 639 867 643
rect 871 639 872 643
rect 866 638 872 639
rect 1058 643 1064 644
rect 1058 639 1059 643
rect 1063 639 1064 643
rect 1058 638 1064 639
rect 1250 643 1256 644
rect 1250 639 1251 643
rect 1255 639 1256 643
rect 1250 638 1256 639
rect 1434 643 1440 644
rect 1434 639 1435 643
rect 1439 639 1440 643
rect 1434 638 1440 639
rect 1618 643 1624 644
rect 1618 639 1619 643
rect 1623 639 1624 643
rect 1618 638 1624 639
rect 1786 643 1792 644
rect 1786 639 1787 643
rect 1791 639 1792 643
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 1786 638 1792 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 318 628 324 629
rect 318 624 319 628
rect 323 624 324 628
rect 318 623 324 624
rect 510 628 516 629
rect 510 624 511 628
rect 515 624 516 628
rect 510 623 516 624
rect 702 628 708 629
rect 702 624 703 628
rect 707 624 708 628
rect 702 623 708 624
rect 894 628 900 629
rect 894 624 895 628
rect 899 624 900 628
rect 894 623 900 624
rect 1086 628 1092 629
rect 1086 624 1087 628
rect 1091 624 1092 628
rect 1086 623 1092 624
rect 1278 628 1284 629
rect 1278 624 1279 628
rect 1283 624 1284 628
rect 1278 623 1284 624
rect 1462 628 1468 629
rect 1462 624 1463 628
rect 1467 624 1468 628
rect 1462 623 1468 624
rect 1646 628 1652 629
rect 1646 624 1647 628
rect 1651 624 1652 628
rect 1646 623 1652 624
rect 1814 628 1820 629
rect 1814 624 1815 628
rect 1819 624 1820 628
rect 1814 623 1820 624
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 110 622 116 623
rect 112 599 114 622
rect 160 599 162 623
rect 320 599 322 623
rect 512 599 514 623
rect 704 599 706 623
rect 896 599 898 623
rect 1088 599 1090 623
rect 1280 599 1282 623
rect 1464 599 1466 623
rect 1648 599 1650 623
rect 1816 599 1818 623
rect 1934 622 1940 623
rect 1936 599 1938 622
rect 111 598 115 599
rect 111 593 115 594
rect 159 598 163 599
rect 159 593 163 594
rect 319 598 323 599
rect 319 593 323 594
rect 327 598 331 599
rect 327 593 331 594
rect 511 598 515 599
rect 511 593 515 594
rect 519 598 523 599
rect 519 593 523 594
rect 703 598 707 599
rect 703 593 707 594
rect 711 598 715 599
rect 711 593 715 594
rect 895 598 899 599
rect 895 593 899 594
rect 903 598 907 599
rect 903 593 907 594
rect 1087 598 1091 599
rect 1087 593 1091 594
rect 1095 598 1099 599
rect 1095 593 1099 594
rect 1279 598 1283 599
rect 1279 593 1283 594
rect 1463 598 1467 599
rect 1463 593 1467 594
rect 1647 598 1651 599
rect 1647 593 1651 594
rect 1815 598 1819 599
rect 1815 593 1819 594
rect 1935 598 1939 599
rect 1935 593 1939 594
rect 112 570 114 593
rect 110 569 116 570
rect 160 569 162 593
rect 328 569 330 593
rect 520 569 522 593
rect 712 569 714 593
rect 904 569 906 593
rect 1096 569 1098 593
rect 1280 569 1282 593
rect 1464 569 1466 593
rect 1648 569 1650 593
rect 1816 569 1818 593
rect 1936 570 1938 593
rect 1934 569 1940 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 326 568 332 569
rect 326 564 327 568
rect 331 564 332 568
rect 326 563 332 564
rect 518 568 524 569
rect 518 564 519 568
rect 523 564 524 568
rect 518 563 524 564
rect 710 568 716 569
rect 710 564 711 568
rect 715 564 716 568
rect 710 563 716 564
rect 902 568 908 569
rect 902 564 903 568
rect 907 564 908 568
rect 902 563 908 564
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 1094 563 1100 564
rect 1278 568 1284 569
rect 1278 564 1279 568
rect 1283 564 1284 568
rect 1278 563 1284 564
rect 1462 568 1468 569
rect 1462 564 1463 568
rect 1467 564 1468 568
rect 1462 563 1468 564
rect 1646 568 1652 569
rect 1646 564 1647 568
rect 1651 564 1652 568
rect 1646 563 1652 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 1814 563 1820 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 298 553 304 554
rect 298 549 299 553
rect 303 549 304 553
rect 298 548 304 549
rect 490 553 496 554
rect 490 549 491 553
rect 495 549 496 553
rect 490 548 496 549
rect 682 553 688 554
rect 682 549 683 553
rect 687 549 688 553
rect 682 548 688 549
rect 874 553 880 554
rect 874 549 875 553
rect 879 549 880 553
rect 874 548 880 549
rect 1066 553 1072 554
rect 1066 549 1067 553
rect 1071 549 1072 553
rect 1066 548 1072 549
rect 1250 553 1256 554
rect 1250 549 1251 553
rect 1255 549 1256 553
rect 1250 548 1256 549
rect 1434 553 1440 554
rect 1434 549 1435 553
rect 1439 549 1440 553
rect 1434 548 1440 549
rect 1618 553 1624 554
rect 1618 549 1619 553
rect 1623 549 1624 553
rect 1618 548 1624 549
rect 1786 553 1792 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 110 547 116 548
rect 112 487 114 547
rect 132 487 134 548
rect 300 487 302 548
rect 492 487 494 548
rect 684 487 686 548
rect 876 487 878 548
rect 1068 487 1070 548
rect 1252 487 1254 548
rect 1436 487 1438 548
rect 1620 487 1622 548
rect 1788 487 1790 548
rect 1934 547 1940 548
rect 1936 487 1938 547
rect 111 486 115 487
rect 111 481 115 482
rect 131 486 135 487
rect 131 481 135 482
rect 299 486 303 487
rect 299 481 303 482
rect 395 486 399 487
rect 395 481 399 482
rect 491 486 495 487
rect 491 481 495 482
rect 587 486 591 487
rect 587 481 591 482
rect 683 486 687 487
rect 683 481 687 482
rect 787 486 791 487
rect 787 481 791 482
rect 875 486 879 487
rect 875 481 879 482
rect 987 486 991 487
rect 987 481 991 482
rect 1067 486 1071 487
rect 1067 481 1071 482
rect 1195 486 1199 487
rect 1195 481 1199 482
rect 1251 486 1255 487
rect 1251 481 1255 482
rect 1411 486 1415 487
rect 1411 481 1415 482
rect 1435 486 1439 487
rect 1435 481 1439 482
rect 1619 486 1623 487
rect 1619 481 1623 482
rect 1787 486 1791 487
rect 1787 481 1791 482
rect 1935 486 1939 487
rect 1935 481 1939 482
rect 112 421 114 481
rect 110 420 116 421
rect 396 420 398 481
rect 588 420 590 481
rect 788 420 790 481
rect 988 420 990 481
rect 1196 420 1198 481
rect 1412 420 1414 481
rect 1936 421 1938 481
rect 1976 467 1978 687
rect 3108 467 3110 688
rect 3244 467 3246 688
rect 3380 467 3382 688
rect 3516 467 3518 688
rect 3652 467 3654 688
rect 3798 687 3804 688
rect 3839 690 3843 691
rect 3800 467 3802 687
rect 3839 685 3843 686
rect 3859 690 3863 691
rect 3859 685 3863 686
rect 3955 690 3959 691
rect 3955 685 3959 686
rect 3995 690 3999 691
rect 3995 685 3999 686
rect 4139 690 4143 691
rect 4139 685 4143 686
rect 4211 690 4215 691
rect 4211 685 4215 686
rect 4323 690 4327 691
rect 4323 685 4327 686
rect 4507 690 4511 691
rect 4507 685 4511 686
rect 4531 690 4535 691
rect 4531 685 4535 686
rect 4755 690 4759 691
rect 4755 685 4759 686
rect 4835 690 4839 691
rect 4835 685 4839 686
rect 4995 690 4999 691
rect 4995 685 4999 686
rect 5187 690 5191 691
rect 5187 685 5191 686
rect 5243 690 5247 691
rect 5243 685 5247 686
rect 5499 690 5503 691
rect 5499 685 5503 686
rect 5515 690 5519 691
rect 5515 685 5519 686
rect 5663 690 5667 691
rect 5663 685 5667 686
rect 3840 625 3842 685
rect 3838 624 3844 625
rect 3860 624 3862 685
rect 3996 624 3998 685
rect 4140 624 4142 685
rect 4324 624 4326 685
rect 4532 624 4534 685
rect 4756 624 4758 685
rect 4996 624 4998 685
rect 5244 624 5246 685
rect 5500 624 5502 685
rect 5664 625 5666 685
rect 5662 624 5668 625
rect 3838 620 3839 624
rect 3843 620 3844 624
rect 3838 619 3844 620
rect 3858 623 3864 624
rect 3858 619 3859 623
rect 3863 619 3864 623
rect 3858 618 3864 619
rect 3994 623 4000 624
rect 3994 619 3995 623
rect 3999 619 4000 623
rect 3994 618 4000 619
rect 4138 623 4144 624
rect 4138 619 4139 623
rect 4143 619 4144 623
rect 4138 618 4144 619
rect 4322 623 4328 624
rect 4322 619 4323 623
rect 4327 619 4328 623
rect 4322 618 4328 619
rect 4530 623 4536 624
rect 4530 619 4531 623
rect 4535 619 4536 623
rect 4530 618 4536 619
rect 4754 623 4760 624
rect 4754 619 4755 623
rect 4759 619 4760 623
rect 4754 618 4760 619
rect 4994 623 5000 624
rect 4994 619 4995 623
rect 4999 619 5000 623
rect 4994 618 5000 619
rect 5242 623 5248 624
rect 5242 619 5243 623
rect 5247 619 5248 623
rect 5242 618 5248 619
rect 5498 623 5504 624
rect 5498 619 5499 623
rect 5503 619 5504 623
rect 5662 620 5663 624
rect 5667 620 5668 624
rect 5662 619 5668 620
rect 5498 618 5504 619
rect 3886 608 3892 609
rect 3838 607 3844 608
rect 3838 603 3839 607
rect 3843 603 3844 607
rect 3886 604 3887 608
rect 3891 604 3892 608
rect 3886 603 3892 604
rect 4022 608 4028 609
rect 4022 604 4023 608
rect 4027 604 4028 608
rect 4022 603 4028 604
rect 4166 608 4172 609
rect 4166 604 4167 608
rect 4171 604 4172 608
rect 4166 603 4172 604
rect 4350 608 4356 609
rect 4350 604 4351 608
rect 4355 604 4356 608
rect 4350 603 4356 604
rect 4558 608 4564 609
rect 4558 604 4559 608
rect 4563 604 4564 608
rect 4558 603 4564 604
rect 4782 608 4788 609
rect 4782 604 4783 608
rect 4787 604 4788 608
rect 4782 603 4788 604
rect 5022 608 5028 609
rect 5022 604 5023 608
rect 5027 604 5028 608
rect 5022 603 5028 604
rect 5270 608 5276 609
rect 5270 604 5271 608
rect 5275 604 5276 608
rect 5270 603 5276 604
rect 5526 608 5532 609
rect 5526 604 5527 608
rect 5531 604 5532 608
rect 5526 603 5532 604
rect 5662 607 5668 608
rect 5662 603 5663 607
rect 5667 603 5668 607
rect 3838 602 3844 603
rect 3840 579 3842 602
rect 3888 579 3890 603
rect 4024 579 4026 603
rect 4168 579 4170 603
rect 4352 579 4354 603
rect 4560 579 4562 603
rect 4784 579 4786 603
rect 5024 579 5026 603
rect 5272 579 5274 603
rect 5528 579 5530 603
rect 5662 602 5668 603
rect 5664 579 5666 602
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3887 578 3891 579
rect 3887 573 3891 574
rect 4023 578 4027 579
rect 4023 573 4027 574
rect 4159 578 4163 579
rect 4159 573 4163 574
rect 4167 578 4171 579
rect 4167 573 4171 574
rect 4295 578 4299 579
rect 4295 573 4299 574
rect 4351 578 4355 579
rect 4351 573 4355 574
rect 4431 578 4435 579
rect 4431 573 4435 574
rect 4559 578 4563 579
rect 4559 573 4563 574
rect 4575 578 4579 579
rect 4575 573 4579 574
rect 4743 578 4747 579
rect 4743 573 4747 574
rect 4783 578 4787 579
rect 4783 573 4787 574
rect 4927 578 4931 579
rect 4927 573 4931 574
rect 5023 578 5027 579
rect 5023 573 5027 574
rect 5119 578 5123 579
rect 5119 573 5123 574
rect 5271 578 5275 579
rect 5271 573 5275 574
rect 5319 578 5323 579
rect 5319 573 5323 574
rect 5527 578 5531 579
rect 5527 573 5531 574
rect 5663 578 5667 579
rect 5663 573 5667 574
rect 3840 550 3842 573
rect 3838 549 3844 550
rect 3888 549 3890 573
rect 4024 549 4026 573
rect 4160 549 4162 573
rect 4296 549 4298 573
rect 4432 549 4434 573
rect 4576 549 4578 573
rect 4744 549 4746 573
rect 4928 549 4930 573
rect 5120 549 5122 573
rect 5320 549 5322 573
rect 5528 549 5530 573
rect 5664 550 5666 573
rect 5662 549 5668 550
rect 3838 545 3839 549
rect 3843 545 3844 549
rect 3838 544 3844 545
rect 3886 548 3892 549
rect 3886 544 3887 548
rect 3891 544 3892 548
rect 3886 543 3892 544
rect 4022 548 4028 549
rect 4022 544 4023 548
rect 4027 544 4028 548
rect 4022 543 4028 544
rect 4158 548 4164 549
rect 4158 544 4159 548
rect 4163 544 4164 548
rect 4158 543 4164 544
rect 4294 548 4300 549
rect 4294 544 4295 548
rect 4299 544 4300 548
rect 4294 543 4300 544
rect 4430 548 4436 549
rect 4430 544 4431 548
rect 4435 544 4436 548
rect 4430 543 4436 544
rect 4574 548 4580 549
rect 4574 544 4575 548
rect 4579 544 4580 548
rect 4574 543 4580 544
rect 4742 548 4748 549
rect 4742 544 4743 548
rect 4747 544 4748 548
rect 4742 543 4748 544
rect 4926 548 4932 549
rect 4926 544 4927 548
rect 4931 544 4932 548
rect 4926 543 4932 544
rect 5118 548 5124 549
rect 5118 544 5119 548
rect 5123 544 5124 548
rect 5118 543 5124 544
rect 5318 548 5324 549
rect 5318 544 5319 548
rect 5323 544 5324 548
rect 5318 543 5324 544
rect 5526 548 5532 549
rect 5526 544 5527 548
rect 5531 544 5532 548
rect 5662 545 5663 549
rect 5667 545 5668 549
rect 5662 544 5668 545
rect 5526 543 5532 544
rect 3858 533 3864 534
rect 3838 532 3844 533
rect 3838 528 3839 532
rect 3843 528 3844 532
rect 3858 529 3859 533
rect 3863 529 3864 533
rect 3858 528 3864 529
rect 3994 533 4000 534
rect 3994 529 3995 533
rect 3999 529 4000 533
rect 3994 528 4000 529
rect 4130 533 4136 534
rect 4130 529 4131 533
rect 4135 529 4136 533
rect 4130 528 4136 529
rect 4266 533 4272 534
rect 4266 529 4267 533
rect 4271 529 4272 533
rect 4266 528 4272 529
rect 4402 533 4408 534
rect 4402 529 4403 533
rect 4407 529 4408 533
rect 4402 528 4408 529
rect 4546 533 4552 534
rect 4546 529 4547 533
rect 4551 529 4552 533
rect 4546 528 4552 529
rect 4714 533 4720 534
rect 4714 529 4715 533
rect 4719 529 4720 533
rect 4714 528 4720 529
rect 4898 533 4904 534
rect 4898 529 4899 533
rect 4903 529 4904 533
rect 4898 528 4904 529
rect 5090 533 5096 534
rect 5090 529 5091 533
rect 5095 529 5096 533
rect 5090 528 5096 529
rect 5290 533 5296 534
rect 5290 529 5291 533
rect 5295 529 5296 533
rect 5290 528 5296 529
rect 5498 533 5504 534
rect 5498 529 5499 533
rect 5503 529 5504 533
rect 5498 528 5504 529
rect 5662 532 5668 533
rect 5662 528 5663 532
rect 5667 528 5668 532
rect 3838 527 3844 528
rect 3840 467 3842 527
rect 3860 467 3862 528
rect 3996 467 3998 528
rect 4132 467 4134 528
rect 4268 467 4270 528
rect 4404 467 4406 528
rect 4548 467 4550 528
rect 4716 467 4718 528
rect 4900 467 4902 528
rect 5092 467 5094 528
rect 5292 467 5294 528
rect 5500 467 5502 528
rect 5662 527 5668 528
rect 5664 467 5666 527
rect 1975 466 1979 467
rect 1975 461 1979 462
rect 1995 466 1999 467
rect 1995 461 1999 462
rect 2203 466 2207 467
rect 2203 461 2207 462
rect 2427 466 2431 467
rect 2427 461 2431 462
rect 2651 466 2655 467
rect 2651 461 2655 462
rect 2867 466 2871 467
rect 2867 461 2871 462
rect 3075 466 3079 467
rect 3075 461 3079 462
rect 3107 466 3111 467
rect 3107 461 3111 462
rect 3243 466 3247 467
rect 3243 461 3247 462
rect 3275 466 3279 467
rect 3275 461 3279 462
rect 3379 466 3383 467
rect 3379 461 3383 462
rect 3475 466 3479 467
rect 3475 461 3479 462
rect 3515 466 3519 467
rect 3515 461 3519 462
rect 3651 466 3655 467
rect 3651 461 3655 462
rect 3799 466 3803 467
rect 3799 461 3803 462
rect 3839 466 3843 467
rect 3839 461 3843 462
rect 3859 466 3863 467
rect 3859 461 3863 462
rect 3995 466 3999 467
rect 3995 461 3999 462
rect 4131 466 4135 467
rect 4131 461 4135 462
rect 4267 466 4271 467
rect 4267 461 4271 462
rect 4379 466 4383 467
rect 4379 461 4383 462
rect 4403 466 4407 467
rect 4403 461 4407 462
rect 4547 466 4551 467
rect 4547 461 4551 462
rect 4595 466 4599 467
rect 4595 461 4599 462
rect 4715 466 4719 467
rect 4715 461 4719 462
rect 4819 466 4823 467
rect 4819 461 4823 462
rect 4899 466 4903 467
rect 4899 461 4903 462
rect 5051 466 5055 467
rect 5051 461 5055 462
rect 5091 466 5095 467
rect 5091 461 5095 462
rect 5283 466 5287 467
rect 5283 461 5287 462
rect 5291 466 5295 467
rect 5291 461 5295 462
rect 5499 466 5503 467
rect 5499 461 5503 462
rect 5663 466 5667 467
rect 5663 461 5667 462
rect 1934 420 1940 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 394 419 400 420
rect 394 415 395 419
rect 399 415 400 419
rect 394 414 400 415
rect 586 419 592 420
rect 586 415 587 419
rect 591 415 592 419
rect 586 414 592 415
rect 786 419 792 420
rect 786 415 787 419
rect 791 415 792 419
rect 786 414 792 415
rect 986 419 992 420
rect 986 415 987 419
rect 991 415 992 419
rect 986 414 992 415
rect 1194 419 1200 420
rect 1194 415 1195 419
rect 1199 415 1200 419
rect 1194 414 1200 415
rect 1410 419 1416 420
rect 1410 415 1411 419
rect 1415 415 1416 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 1410 414 1416 415
rect 422 404 428 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 422 400 423 404
rect 427 400 428 404
rect 422 399 428 400
rect 614 404 620 405
rect 614 400 615 404
rect 619 400 620 404
rect 614 399 620 400
rect 814 404 820 405
rect 814 400 815 404
rect 819 400 820 404
rect 814 399 820 400
rect 1014 404 1020 405
rect 1014 400 1015 404
rect 1019 400 1020 404
rect 1014 399 1020 400
rect 1222 404 1228 405
rect 1222 400 1223 404
rect 1227 400 1228 404
rect 1222 399 1228 400
rect 1438 404 1444 405
rect 1438 400 1439 404
rect 1443 400 1444 404
rect 1438 399 1444 400
rect 1934 403 1940 404
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 1976 401 1978 461
rect 110 398 116 399
rect 112 363 114 398
rect 424 363 426 399
rect 616 363 618 399
rect 816 363 818 399
rect 1016 363 1018 399
rect 1224 363 1226 399
rect 1440 363 1442 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 1996 400 1998 461
rect 2204 400 2206 461
rect 2428 400 2430 461
rect 2652 400 2654 461
rect 2868 400 2870 461
rect 3076 400 3078 461
rect 3276 400 3278 461
rect 3476 400 3478 461
rect 3652 400 3654 461
rect 3800 401 3802 461
rect 3840 401 3842 461
rect 3798 400 3804 401
rect 1936 363 1938 398
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2866 399 2872 400
rect 2866 395 2867 399
rect 2871 395 2872 399
rect 2866 394 2872 395
rect 3074 399 3080 400
rect 3074 395 3075 399
rect 3079 395 3080 399
rect 3074 394 3080 395
rect 3274 399 3280 400
rect 3274 395 3275 399
rect 3279 395 3280 399
rect 3274 394 3280 395
rect 3474 399 3480 400
rect 3474 395 3475 399
rect 3479 395 3480 399
rect 3474 394 3480 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3838 400 3844 401
rect 4380 400 4382 461
rect 4596 400 4598 461
rect 4820 400 4822 461
rect 5052 400 5054 461
rect 5284 400 5286 461
rect 5664 401 5666 461
rect 5662 400 5668 401
rect 3838 396 3839 400
rect 3843 396 3844 400
rect 3838 395 3844 396
rect 4378 399 4384 400
rect 4378 395 4379 399
rect 4383 395 4384 399
rect 3650 394 3656 395
rect 4378 394 4384 395
rect 4594 399 4600 400
rect 4594 395 4595 399
rect 4599 395 4600 399
rect 4594 394 4600 395
rect 4818 399 4824 400
rect 4818 395 4819 399
rect 4823 395 4824 399
rect 4818 394 4824 395
rect 5050 399 5056 400
rect 5050 395 5051 399
rect 5055 395 5056 399
rect 5050 394 5056 395
rect 5282 399 5288 400
rect 5282 395 5283 399
rect 5287 395 5288 399
rect 5662 396 5663 400
rect 5667 396 5668 400
rect 5662 395 5668 396
rect 5282 394 5288 395
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 2894 384 2900 385
rect 2894 380 2895 384
rect 2899 380 2900 384
rect 2894 379 2900 380
rect 3102 384 3108 385
rect 3102 380 3103 384
rect 3107 380 3108 384
rect 3102 379 3108 380
rect 3302 384 3308 385
rect 3302 380 3303 384
rect 3307 380 3308 384
rect 3302 379 3308 380
rect 3502 384 3508 385
rect 3502 380 3503 384
rect 3507 380 3508 384
rect 3502 379 3508 380
rect 3678 384 3684 385
rect 4406 384 4412 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 111 362 115 363
rect 111 357 115 358
rect 423 362 427 363
rect 423 357 427 358
rect 615 362 619 363
rect 615 357 619 358
rect 647 362 651 363
rect 647 357 651 358
rect 815 362 819 363
rect 815 357 819 358
rect 991 362 995 363
rect 991 357 995 358
rect 1015 362 1019 363
rect 1015 357 1019 358
rect 1167 362 1171 363
rect 1167 357 1171 358
rect 1223 362 1227 363
rect 1223 357 1227 358
rect 1343 362 1347 363
rect 1343 357 1347 358
rect 1439 362 1443 363
rect 1439 357 1443 358
rect 1935 362 1939 363
rect 1935 357 1939 358
rect 112 334 114 357
rect 110 333 116 334
rect 648 333 650 357
rect 816 333 818 357
rect 992 333 994 357
rect 1168 333 1170 357
rect 1344 333 1346 357
rect 1936 334 1938 357
rect 1976 339 1978 378
rect 2024 339 2026 379
rect 2232 339 2234 379
rect 2456 339 2458 379
rect 2680 339 2682 379
rect 2896 339 2898 379
rect 3104 339 3106 379
rect 3304 339 3306 379
rect 3504 339 3506 379
rect 3680 339 3682 379
rect 3798 378 3804 379
rect 3838 383 3844 384
rect 3838 379 3839 383
rect 3843 379 3844 383
rect 4406 380 4407 384
rect 4411 380 4412 384
rect 4406 379 4412 380
rect 4622 384 4628 385
rect 4622 380 4623 384
rect 4627 380 4628 384
rect 4622 379 4628 380
rect 4846 384 4852 385
rect 4846 380 4847 384
rect 4851 380 4852 384
rect 4846 379 4852 380
rect 5078 384 5084 385
rect 5078 380 5079 384
rect 5083 380 5084 384
rect 5078 379 5084 380
rect 5310 384 5316 385
rect 5310 380 5311 384
rect 5315 380 5316 384
rect 5310 379 5316 380
rect 5662 383 5668 384
rect 5662 379 5663 383
rect 5667 379 5668 383
rect 3838 378 3844 379
rect 3800 339 3802 378
rect 3840 355 3842 378
rect 4408 355 4410 379
rect 4624 355 4626 379
rect 4848 355 4850 379
rect 5080 355 5082 379
rect 5312 355 5314 379
rect 5662 378 5668 379
rect 5664 355 5666 378
rect 3839 354 3843 355
rect 3839 349 3843 350
rect 4407 354 4411 355
rect 4407 349 4411 350
rect 4623 354 4627 355
rect 4623 349 4627 350
rect 4639 354 4643 355
rect 4639 349 4643 350
rect 4807 354 4811 355
rect 4807 349 4811 350
rect 4847 354 4851 355
rect 4847 349 4851 350
rect 4983 354 4987 355
rect 4983 349 4987 350
rect 5079 354 5083 355
rect 5079 349 5083 350
rect 5167 354 5171 355
rect 5167 349 5171 350
rect 5311 354 5315 355
rect 5311 349 5315 350
rect 5359 354 5363 355
rect 5359 349 5363 350
rect 5543 354 5547 355
rect 5543 349 5547 350
rect 5663 354 5667 355
rect 5663 349 5667 350
rect 1975 338 1979 339
rect 1934 333 1940 334
rect 1975 333 1979 334
rect 2023 338 2027 339
rect 2023 333 2027 334
rect 2159 338 2163 339
rect 2159 333 2163 334
rect 2231 338 2235 339
rect 2231 333 2235 334
rect 2295 338 2299 339
rect 2295 333 2299 334
rect 2431 338 2435 339
rect 2431 333 2435 334
rect 2455 338 2459 339
rect 2455 333 2459 334
rect 2567 338 2571 339
rect 2567 333 2571 334
rect 2679 338 2683 339
rect 2679 333 2683 334
rect 2703 338 2707 339
rect 2703 333 2707 334
rect 2839 338 2843 339
rect 2839 333 2843 334
rect 2895 338 2899 339
rect 2895 333 2899 334
rect 2975 338 2979 339
rect 2975 333 2979 334
rect 3103 338 3107 339
rect 3103 333 3107 334
rect 3111 338 3115 339
rect 3111 333 3115 334
rect 3247 338 3251 339
rect 3247 333 3251 334
rect 3303 338 3307 339
rect 3303 333 3307 334
rect 3383 338 3387 339
rect 3383 333 3387 334
rect 3503 338 3507 339
rect 3503 333 3507 334
rect 3519 338 3523 339
rect 3519 333 3523 334
rect 3655 338 3659 339
rect 3655 333 3659 334
rect 3679 338 3683 339
rect 3679 333 3683 334
rect 3799 338 3803 339
rect 3799 333 3803 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 646 332 652 333
rect 646 328 647 332
rect 651 328 652 332
rect 646 327 652 328
rect 814 332 820 333
rect 814 328 815 332
rect 819 328 820 332
rect 814 327 820 328
rect 990 332 996 333
rect 990 328 991 332
rect 995 328 996 332
rect 990 327 996 328
rect 1166 332 1172 333
rect 1166 328 1167 332
rect 1171 328 1172 332
rect 1166 327 1172 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 1342 327 1348 328
rect 618 317 624 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 618 313 619 317
rect 623 313 624 317
rect 618 312 624 313
rect 786 317 792 318
rect 786 313 787 317
rect 791 313 792 317
rect 786 312 792 313
rect 962 317 968 318
rect 962 313 963 317
rect 967 313 968 317
rect 962 312 968 313
rect 1138 317 1144 318
rect 1138 313 1139 317
rect 1143 313 1144 317
rect 1138 312 1144 313
rect 1314 317 1320 318
rect 1314 313 1315 317
rect 1319 313 1320 317
rect 1314 312 1320 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 110 311 116 312
rect 112 211 114 311
rect 620 211 622 312
rect 788 211 790 312
rect 964 211 966 312
rect 1140 211 1142 312
rect 1316 211 1318 312
rect 1934 311 1940 312
rect 1936 211 1938 311
rect 1976 310 1978 333
rect 1974 309 1980 310
rect 2024 309 2026 333
rect 2160 309 2162 333
rect 2296 309 2298 333
rect 2432 309 2434 333
rect 2568 309 2570 333
rect 2704 309 2706 333
rect 2840 309 2842 333
rect 2976 309 2978 333
rect 3112 309 3114 333
rect 3248 309 3250 333
rect 3384 309 3386 333
rect 3520 309 3522 333
rect 3656 309 3658 333
rect 3800 310 3802 333
rect 3840 326 3842 349
rect 3838 325 3844 326
rect 4640 325 4642 349
rect 4808 325 4810 349
rect 4984 325 4986 349
rect 5168 325 5170 349
rect 5360 325 5362 349
rect 5544 325 5546 349
rect 5664 326 5666 349
rect 5662 325 5668 326
rect 3838 321 3839 325
rect 3843 321 3844 325
rect 3838 320 3844 321
rect 4638 324 4644 325
rect 4638 320 4639 324
rect 4643 320 4644 324
rect 4638 319 4644 320
rect 4806 324 4812 325
rect 4806 320 4807 324
rect 4811 320 4812 324
rect 4806 319 4812 320
rect 4982 324 4988 325
rect 4982 320 4983 324
rect 4987 320 4988 324
rect 4982 319 4988 320
rect 5166 324 5172 325
rect 5166 320 5167 324
rect 5171 320 5172 324
rect 5166 319 5172 320
rect 5358 324 5364 325
rect 5358 320 5359 324
rect 5363 320 5364 324
rect 5358 319 5364 320
rect 5542 324 5548 325
rect 5542 320 5543 324
rect 5547 320 5548 324
rect 5662 321 5663 325
rect 5667 321 5668 325
rect 5662 320 5668 321
rect 5542 319 5548 320
rect 3798 309 3804 310
rect 4610 309 4616 310
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3798 304 3804 305
rect 3838 308 3844 309
rect 3838 304 3839 308
rect 3843 304 3844 308
rect 4610 305 4611 309
rect 4615 305 4616 309
rect 4610 304 4616 305
rect 4778 309 4784 310
rect 4778 305 4779 309
rect 4783 305 4784 309
rect 4778 304 4784 305
rect 4954 309 4960 310
rect 4954 305 4955 309
rect 4959 305 4960 309
rect 4954 304 4960 305
rect 5138 309 5144 310
rect 5138 305 5139 309
rect 5143 305 5144 309
rect 5138 304 5144 305
rect 5330 309 5336 310
rect 5330 305 5331 309
rect 5335 305 5336 309
rect 5330 304 5336 305
rect 5514 309 5520 310
rect 5514 305 5515 309
rect 5519 305 5520 309
rect 5514 304 5520 305
rect 5662 308 5668 309
rect 5662 304 5663 308
rect 5667 304 5668 308
rect 3654 303 3660 304
rect 3838 303 3844 304
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 1974 287 1980 288
rect 111 210 115 211
rect 111 205 115 206
rect 539 210 543 211
rect 539 205 543 206
rect 619 210 623 211
rect 619 205 623 206
rect 675 210 679 211
rect 675 205 679 206
rect 787 210 791 211
rect 787 205 791 206
rect 811 210 815 211
rect 811 205 815 206
rect 947 210 951 211
rect 947 205 951 206
rect 963 210 967 211
rect 963 205 967 206
rect 1083 210 1087 211
rect 1083 205 1087 206
rect 1139 210 1143 211
rect 1139 205 1143 206
rect 1219 210 1223 211
rect 1219 205 1223 206
rect 1315 210 1319 211
rect 1315 205 1319 206
rect 1355 210 1359 211
rect 1355 205 1359 206
rect 1491 210 1495 211
rect 1491 205 1495 206
rect 1935 210 1939 211
rect 1935 205 1939 206
rect 112 145 114 205
rect 110 144 116 145
rect 540 144 542 205
rect 676 144 678 205
rect 812 144 814 205
rect 948 144 950 205
rect 1084 144 1086 205
rect 1220 144 1222 205
rect 1356 144 1358 205
rect 1492 144 1494 205
rect 1936 145 1938 205
rect 1976 191 1978 287
rect 1996 191 1998 288
rect 2132 191 2134 288
rect 2268 191 2270 288
rect 2404 191 2406 288
rect 2540 191 2542 288
rect 2676 191 2678 288
rect 2812 191 2814 288
rect 2948 191 2950 288
rect 3084 191 3086 288
rect 3220 191 3222 288
rect 3356 191 3358 288
rect 3492 191 3494 288
rect 3628 191 3630 288
rect 3798 287 3804 288
rect 3800 191 3802 287
rect 3840 215 3842 303
rect 4612 215 4614 304
rect 4780 215 4782 304
rect 4956 215 4958 304
rect 5140 215 5142 304
rect 5332 215 5334 304
rect 5516 215 5518 304
rect 5662 303 5668 304
rect 5664 215 5666 303
rect 3839 214 3843 215
rect 3839 209 3843 210
rect 4291 214 4295 215
rect 4291 209 4295 210
rect 4427 214 4431 215
rect 4427 209 4431 210
rect 4563 214 4567 215
rect 4563 209 4567 210
rect 4611 214 4615 215
rect 4611 209 4615 210
rect 4699 214 4703 215
rect 4699 209 4703 210
rect 4779 214 4783 215
rect 4779 209 4783 210
rect 4835 214 4839 215
rect 4835 209 4839 210
rect 4955 214 4959 215
rect 4955 209 4959 210
rect 4971 214 4975 215
rect 4971 209 4975 210
rect 5107 214 5111 215
rect 5107 209 5111 210
rect 5139 214 5143 215
rect 5139 209 5143 210
rect 5243 214 5247 215
rect 5243 209 5247 210
rect 5331 214 5335 215
rect 5331 209 5335 210
rect 5379 214 5383 215
rect 5379 209 5383 210
rect 5515 214 5519 215
rect 5515 209 5519 210
rect 5663 214 5667 215
rect 5663 209 5667 210
rect 1975 190 1979 191
rect 1975 185 1979 186
rect 1995 190 1999 191
rect 1995 185 1999 186
rect 2131 190 2135 191
rect 2131 185 2135 186
rect 2267 190 2271 191
rect 2267 185 2271 186
rect 2403 190 2407 191
rect 2403 185 2407 186
rect 2539 190 2543 191
rect 2539 185 2543 186
rect 2675 190 2679 191
rect 2675 185 2679 186
rect 2811 190 2815 191
rect 2811 185 2815 186
rect 2947 190 2951 191
rect 2947 185 2951 186
rect 3083 190 3087 191
rect 3083 185 3087 186
rect 3219 190 3223 191
rect 3219 185 3223 186
rect 3355 190 3359 191
rect 3355 185 3359 186
rect 3491 190 3495 191
rect 3491 185 3495 186
rect 3627 190 3631 191
rect 3627 185 3631 186
rect 3799 190 3803 191
rect 3799 185 3803 186
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1082 138 1088 139
rect 1218 143 1224 144
rect 1218 139 1219 143
rect 1223 139 1224 143
rect 1218 138 1224 139
rect 1354 143 1360 144
rect 1354 139 1355 143
rect 1359 139 1360 143
rect 1354 138 1360 139
rect 1490 143 1496 144
rect 1490 139 1491 143
rect 1495 139 1496 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 1490 138 1496 139
rect 566 128 572 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1246 128 1252 129
rect 1246 124 1247 128
rect 1251 124 1252 128
rect 1246 123 1252 124
rect 1382 128 1388 129
rect 1382 124 1383 128
rect 1387 124 1388 128
rect 1382 123 1388 124
rect 1518 128 1524 129
rect 1518 124 1519 128
rect 1523 124 1524 128
rect 1518 123 1524 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 1976 125 1978 185
rect 110 122 116 123
rect 112 99 114 122
rect 568 99 570 123
rect 704 99 706 123
rect 840 99 842 123
rect 976 99 978 123
rect 1112 99 1114 123
rect 1248 99 1250 123
rect 1384 99 1386 123
rect 1520 99 1522 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 1996 124 1998 185
rect 2132 124 2134 185
rect 2268 124 2270 185
rect 2404 124 2406 185
rect 2540 124 2542 185
rect 2676 124 2678 185
rect 2812 124 2814 185
rect 2948 124 2950 185
rect 3084 124 3086 185
rect 3220 124 3222 185
rect 3356 124 3358 185
rect 3492 124 3494 185
rect 3628 124 3630 185
rect 3800 125 3802 185
rect 3840 149 3842 209
rect 3838 148 3844 149
rect 4292 148 4294 209
rect 4428 148 4430 209
rect 4564 148 4566 209
rect 4700 148 4702 209
rect 4836 148 4838 209
rect 4972 148 4974 209
rect 5108 148 5110 209
rect 5244 148 5246 209
rect 5380 148 5382 209
rect 5516 148 5518 209
rect 5664 149 5666 209
rect 5662 148 5668 149
rect 3838 144 3839 148
rect 3843 144 3844 148
rect 3838 143 3844 144
rect 4290 147 4296 148
rect 4290 143 4291 147
rect 4295 143 4296 147
rect 4290 142 4296 143
rect 4426 147 4432 148
rect 4426 143 4427 147
rect 4431 143 4432 147
rect 4426 142 4432 143
rect 4562 147 4568 148
rect 4562 143 4563 147
rect 4567 143 4568 147
rect 4562 142 4568 143
rect 4698 147 4704 148
rect 4698 143 4699 147
rect 4703 143 4704 147
rect 4698 142 4704 143
rect 4834 147 4840 148
rect 4834 143 4835 147
rect 4839 143 4840 147
rect 4834 142 4840 143
rect 4970 147 4976 148
rect 4970 143 4971 147
rect 4975 143 4976 147
rect 4970 142 4976 143
rect 5106 147 5112 148
rect 5106 143 5107 147
rect 5111 143 5112 147
rect 5106 142 5112 143
rect 5242 147 5248 148
rect 5242 143 5243 147
rect 5247 143 5248 147
rect 5242 142 5248 143
rect 5378 147 5384 148
rect 5378 143 5379 147
rect 5383 143 5384 147
rect 5378 142 5384 143
rect 5514 147 5520 148
rect 5514 143 5515 147
rect 5519 143 5520 147
rect 5662 144 5663 148
rect 5667 144 5668 148
rect 5662 143 5668 144
rect 5514 142 5520 143
rect 4318 132 4324 133
rect 3838 131 3844 132
rect 3838 127 3839 131
rect 3843 127 3844 131
rect 4318 128 4319 132
rect 4323 128 4324 132
rect 4318 127 4324 128
rect 4454 132 4460 133
rect 4454 128 4455 132
rect 4459 128 4460 132
rect 4454 127 4460 128
rect 4590 132 4596 133
rect 4590 128 4591 132
rect 4595 128 4596 132
rect 4590 127 4596 128
rect 4726 132 4732 133
rect 4726 128 4727 132
rect 4731 128 4732 132
rect 4726 127 4732 128
rect 4862 132 4868 133
rect 4862 128 4863 132
rect 4867 128 4868 132
rect 4862 127 4868 128
rect 4998 132 5004 133
rect 4998 128 4999 132
rect 5003 128 5004 132
rect 4998 127 5004 128
rect 5134 132 5140 133
rect 5134 128 5135 132
rect 5139 128 5140 132
rect 5134 127 5140 128
rect 5270 132 5276 133
rect 5270 128 5271 132
rect 5275 128 5276 132
rect 5270 127 5276 128
rect 5406 132 5412 133
rect 5406 128 5407 132
rect 5411 128 5412 132
rect 5406 127 5412 128
rect 5542 132 5548 133
rect 5542 128 5543 132
rect 5547 128 5548 132
rect 5542 127 5548 128
rect 5662 131 5668 132
rect 5662 127 5663 131
rect 5667 127 5668 131
rect 3838 126 3844 127
rect 3798 124 3804 125
rect 1936 99 1938 122
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3626 118 3632 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 3840 103 3842 126
rect 4320 103 4322 127
rect 4456 103 4458 127
rect 4592 103 4594 127
rect 4728 103 4730 127
rect 4864 103 4866 127
rect 5000 103 5002 127
rect 5136 103 5138 127
rect 5272 103 5274 127
rect 5408 103 5410 127
rect 5544 103 5546 127
rect 5662 126 5668 127
rect 5664 103 5666 126
rect 1974 102 1980 103
rect 111 98 115 99
rect 111 93 115 94
rect 567 98 571 99
rect 567 93 571 94
rect 703 98 707 99
rect 703 93 707 94
rect 839 98 843 99
rect 839 93 843 94
rect 975 98 979 99
rect 975 93 979 94
rect 1111 98 1115 99
rect 1111 93 1115 94
rect 1247 98 1251 99
rect 1247 93 1251 94
rect 1383 98 1387 99
rect 1383 93 1387 94
rect 1519 98 1523 99
rect 1519 93 1523 94
rect 1935 98 1939 99
rect 1935 93 1939 94
rect 1976 79 1978 102
rect 2024 79 2026 103
rect 2160 79 2162 103
rect 2296 79 2298 103
rect 2432 79 2434 103
rect 2568 79 2570 103
rect 2704 79 2706 103
rect 2840 79 2842 103
rect 2976 79 2978 103
rect 3112 79 3114 103
rect 3248 79 3250 103
rect 3384 79 3386 103
rect 3520 79 3522 103
rect 3656 79 3658 103
rect 3798 102 3804 103
rect 3839 102 3843 103
rect 3800 79 3802 102
rect 3839 97 3843 98
rect 4319 102 4323 103
rect 4319 97 4323 98
rect 4455 102 4459 103
rect 4455 97 4459 98
rect 4591 102 4595 103
rect 4591 97 4595 98
rect 4727 102 4731 103
rect 4727 97 4731 98
rect 4863 102 4867 103
rect 4863 97 4867 98
rect 4999 102 5003 103
rect 4999 97 5003 98
rect 5135 102 5139 103
rect 5135 97 5139 98
rect 5271 102 5275 103
rect 5271 97 5275 98
rect 5407 102 5411 103
rect 5407 97 5411 98
rect 5543 102 5547 103
rect 5543 97 5547 98
rect 5663 102 5667 103
rect 5663 97 5667 98
rect 1975 78 1979 79
rect 1975 73 1979 74
rect 2023 78 2027 79
rect 2023 73 2027 74
rect 2159 78 2163 79
rect 2159 73 2163 74
rect 2295 78 2299 79
rect 2295 73 2299 74
rect 2431 78 2435 79
rect 2431 73 2435 74
rect 2567 78 2571 79
rect 2567 73 2571 74
rect 2703 78 2707 79
rect 2703 73 2707 74
rect 2839 78 2843 79
rect 2839 73 2843 74
rect 2975 78 2979 79
rect 2975 73 2979 74
rect 3111 78 3115 79
rect 3111 73 3115 74
rect 3247 78 3251 79
rect 3247 73 3251 74
rect 3383 78 3387 79
rect 3383 73 3387 74
rect 3519 78 3523 79
rect 3519 73 3523 74
rect 3655 78 3659 79
rect 3655 73 3659 74
rect 3799 78 3803 79
rect 3799 73 3803 74
<< m4c >>
rect 111 5718 115 5722
rect 159 5718 163 5722
rect 303 5718 307 5722
rect 503 5718 507 5722
rect 727 5718 731 5722
rect 983 5718 987 5722
rect 1255 5718 1259 5722
rect 1543 5718 1547 5722
rect 1815 5718 1819 5722
rect 1935 5718 1939 5722
rect 1975 5690 1979 5694
rect 1995 5690 1999 5694
rect 2179 5690 2183 5694
rect 2387 5690 2391 5694
rect 2587 5690 2591 5694
rect 2779 5690 2783 5694
rect 2963 5690 2967 5694
rect 3147 5690 3151 5694
rect 3323 5690 3327 5694
rect 3499 5690 3503 5694
rect 3651 5690 3655 5694
rect 3799 5690 3803 5694
rect 3839 5646 3843 5650
rect 4291 5646 4295 5650
rect 4427 5646 4431 5650
rect 4563 5646 4567 5650
rect 4699 5646 4703 5650
rect 4835 5646 4839 5650
rect 4971 5646 4975 5650
rect 5107 5646 5111 5650
rect 5663 5646 5667 5650
rect 111 5602 115 5606
rect 131 5602 135 5606
rect 275 5602 279 5606
rect 475 5602 479 5606
rect 563 5602 567 5606
rect 699 5602 703 5606
rect 723 5602 727 5606
rect 883 5602 887 5606
rect 955 5602 959 5606
rect 1051 5602 1055 5606
rect 1227 5602 1231 5606
rect 1403 5602 1407 5606
rect 1515 5602 1519 5606
rect 1579 5602 1583 5606
rect 1763 5602 1767 5606
rect 1787 5602 1791 5606
rect 1935 5602 1939 5606
rect 1975 5578 1979 5582
rect 2023 5578 2027 5582
rect 2207 5578 2211 5582
rect 2263 5578 2267 5582
rect 2415 5578 2419 5582
rect 2503 5578 2507 5582
rect 2615 5578 2619 5582
rect 2743 5578 2747 5582
rect 2807 5578 2811 5582
rect 2983 5578 2987 5582
rect 2991 5578 2995 5582
rect 3175 5578 3179 5582
rect 3223 5578 3227 5582
rect 3351 5578 3355 5582
rect 3463 5578 3467 5582
rect 3527 5578 3531 5582
rect 3679 5578 3683 5582
rect 3799 5578 3803 5582
rect 3839 5534 3843 5538
rect 3887 5534 3891 5538
rect 4127 5534 4131 5538
rect 4319 5534 4323 5538
rect 4375 5534 4379 5538
rect 4455 5534 4459 5538
rect 4591 5534 4595 5538
rect 4615 5534 4619 5538
rect 4727 5534 4731 5538
rect 4847 5534 4851 5538
rect 4863 5534 4867 5538
rect 4999 5534 5003 5538
rect 5079 5534 5083 5538
rect 5135 5534 5139 5538
rect 5311 5534 5315 5538
rect 5663 5534 5667 5538
rect 111 5478 115 5482
rect 591 5478 595 5482
rect 727 5478 731 5482
rect 751 5478 755 5482
rect 863 5478 867 5482
rect 911 5478 915 5482
rect 999 5478 1003 5482
rect 1079 5478 1083 5482
rect 1135 5478 1139 5482
rect 1255 5478 1259 5482
rect 1271 5478 1275 5482
rect 1407 5478 1411 5482
rect 1431 5478 1435 5482
rect 1543 5478 1547 5482
rect 1607 5478 1611 5482
rect 1679 5478 1683 5482
rect 1791 5478 1795 5482
rect 1815 5478 1819 5482
rect 1935 5478 1939 5482
rect 1975 5458 1979 5462
rect 2235 5458 2239 5462
rect 2427 5458 2431 5462
rect 2475 5458 2479 5462
rect 2643 5458 2647 5462
rect 2715 5458 2719 5462
rect 2859 5458 2863 5462
rect 2955 5458 2959 5462
rect 3075 5458 3079 5462
rect 3195 5458 3199 5462
rect 3291 5458 3295 5462
rect 3435 5458 3439 5462
rect 3651 5458 3655 5462
rect 3799 5458 3803 5462
rect 3839 5418 3843 5422
rect 3859 5418 3863 5422
rect 4075 5418 4079 5422
rect 4099 5418 4103 5422
rect 4307 5418 4311 5422
rect 4347 5418 4351 5422
rect 4531 5418 4535 5422
rect 4587 5418 4591 5422
rect 4739 5418 4743 5422
rect 4819 5418 4823 5422
rect 4939 5418 4943 5422
rect 5051 5418 5055 5422
rect 5139 5418 5143 5422
rect 5283 5418 5287 5422
rect 5339 5418 5343 5422
rect 5515 5418 5519 5422
rect 5663 5418 5667 5422
rect 1975 5346 1979 5350
rect 2447 5346 2451 5350
rect 2455 5346 2459 5350
rect 2583 5346 2587 5350
rect 2671 5346 2675 5350
rect 2719 5346 2723 5350
rect 2855 5346 2859 5350
rect 2887 5346 2891 5350
rect 2991 5346 2995 5350
rect 3103 5346 3107 5350
rect 3135 5346 3139 5350
rect 3287 5346 3291 5350
rect 3319 5346 3323 5350
rect 3799 5346 3803 5350
rect 111 5262 115 5266
rect 459 5262 463 5266
rect 563 5262 567 5266
rect 595 5262 599 5266
rect 699 5262 703 5266
rect 731 5262 735 5266
rect 835 5262 839 5266
rect 867 5262 871 5266
rect 971 5262 975 5266
rect 1003 5262 1007 5266
rect 1107 5262 1111 5266
rect 1139 5262 1143 5266
rect 1243 5262 1247 5266
rect 1275 5262 1279 5266
rect 1379 5262 1383 5266
rect 1411 5262 1415 5266
rect 1515 5262 1519 5266
rect 1547 5262 1551 5266
rect 1651 5262 1655 5266
rect 1787 5262 1791 5266
rect 1935 5262 1939 5266
rect 3839 5290 3843 5294
rect 3887 5290 3891 5294
rect 4095 5290 4099 5294
rect 4103 5290 4107 5294
rect 4335 5290 4339 5294
rect 4343 5290 4347 5294
rect 4559 5290 4563 5294
rect 4615 5290 4619 5294
rect 4767 5290 4771 5294
rect 4911 5290 4915 5294
rect 4967 5290 4971 5294
rect 5167 5290 5171 5294
rect 5215 5290 5219 5294
rect 5367 5290 5371 5294
rect 5527 5290 5531 5294
rect 5543 5290 5547 5294
rect 5663 5290 5667 5294
rect 1975 5234 1979 5238
rect 2099 5234 2103 5238
rect 2235 5234 2239 5238
rect 2379 5234 2383 5238
rect 2419 5234 2423 5238
rect 2531 5234 2535 5238
rect 2555 5234 2559 5238
rect 2691 5234 2695 5238
rect 2699 5234 2703 5238
rect 2827 5234 2831 5238
rect 2883 5234 2887 5238
rect 2963 5234 2967 5238
rect 3067 5234 3071 5238
rect 3107 5234 3111 5238
rect 3259 5234 3263 5238
rect 3799 5234 3803 5238
rect 3839 5170 3843 5174
rect 3859 5170 3863 5174
rect 3995 5170 3999 5174
rect 4067 5170 4071 5174
rect 4155 5170 4159 5174
rect 4315 5170 4319 5174
rect 4363 5170 4367 5174
rect 4587 5170 4591 5174
rect 4611 5170 4615 5174
rect 4883 5170 4887 5174
rect 5171 5170 5175 5174
rect 5187 5170 5191 5174
rect 5467 5170 5471 5174
rect 5499 5170 5503 5174
rect 5663 5170 5667 5174
rect 111 5134 115 5138
rect 319 5134 323 5138
rect 487 5134 491 5138
rect 503 5134 507 5138
rect 623 5134 627 5138
rect 703 5134 707 5138
rect 759 5134 763 5138
rect 895 5134 899 5138
rect 919 5134 923 5138
rect 1031 5134 1035 5138
rect 1151 5134 1155 5138
rect 1167 5134 1171 5138
rect 1303 5134 1307 5138
rect 1391 5134 1395 5138
rect 1439 5134 1443 5138
rect 1575 5134 1579 5138
rect 1631 5134 1635 5138
rect 1935 5134 1939 5138
rect 1975 5098 1979 5102
rect 2079 5098 2083 5102
rect 2127 5098 2131 5102
rect 2263 5098 2267 5102
rect 2359 5098 2363 5102
rect 2407 5098 2411 5102
rect 2559 5098 2563 5102
rect 2639 5098 2643 5102
rect 2727 5098 2731 5102
rect 2911 5098 2915 5102
rect 3095 5098 3099 5102
rect 3175 5098 3179 5102
rect 3287 5098 3291 5102
rect 3439 5098 3443 5102
rect 3679 5098 3683 5102
rect 3799 5098 3803 5102
rect 111 5022 115 5026
rect 139 5022 143 5026
rect 291 5022 295 5026
rect 411 5022 415 5026
rect 475 5022 479 5026
rect 675 5022 679 5026
rect 683 5022 687 5026
rect 891 5022 895 5026
rect 963 5022 967 5026
rect 1123 5022 1127 5026
rect 1243 5022 1247 5026
rect 1363 5022 1367 5026
rect 1523 5022 1527 5026
rect 1603 5022 1607 5026
rect 1787 5022 1791 5026
rect 1935 5022 1939 5026
rect 3839 5042 3843 5046
rect 3887 5042 3891 5046
rect 4023 5042 4027 5046
rect 4183 5042 4187 5046
rect 4391 5042 4395 5046
rect 4447 5042 4451 5046
rect 4631 5042 4635 5046
rect 4639 5042 4643 5046
rect 4831 5042 4835 5046
rect 4911 5042 4915 5046
rect 5047 5042 5051 5046
rect 5199 5042 5203 5046
rect 5279 5042 5283 5046
rect 5495 5042 5499 5046
rect 5511 5042 5515 5046
rect 5663 5042 5667 5046
rect 1975 4966 1979 4970
rect 1995 4966 1999 4970
rect 2051 4966 2055 4970
rect 2131 4966 2135 4970
rect 2299 4966 2303 4970
rect 2331 4966 2335 4970
rect 2467 4966 2471 4970
rect 2611 4966 2615 4970
rect 2643 4966 2647 4970
rect 2819 4966 2823 4970
rect 2883 4966 2887 4970
rect 2987 4966 2991 4970
rect 3147 4966 3151 4970
rect 3155 4966 3159 4970
rect 3323 4966 3327 4970
rect 3411 4966 3415 4970
rect 3499 4966 3503 4970
rect 3651 4966 3655 4970
rect 3799 4966 3803 4970
rect 111 4910 115 4914
rect 159 4910 163 4914
rect 167 4910 171 4914
rect 415 4910 419 4914
rect 439 4910 443 4914
rect 711 4910 715 4914
rect 735 4910 739 4914
rect 991 4910 995 4914
rect 1087 4910 1091 4914
rect 1271 4910 1275 4914
rect 1463 4910 1467 4914
rect 1551 4910 1555 4914
rect 1815 4910 1819 4914
rect 1935 4910 1939 4914
rect 3839 4914 3843 4918
rect 4419 4914 4423 4918
rect 4603 4914 4607 4918
rect 4675 4914 4679 4918
rect 4803 4914 4807 4918
rect 4827 4914 4831 4918
rect 4987 4914 4991 4918
rect 5019 4914 5023 4918
rect 5155 4914 5159 4918
rect 5251 4914 5255 4918
rect 5323 4914 5327 4918
rect 5483 4914 5487 4918
rect 5499 4914 5503 4918
rect 5663 4914 5667 4918
rect 1975 4826 1979 4830
rect 2023 4826 2027 4830
rect 2159 4826 2163 4830
rect 2327 4826 2331 4830
rect 2391 4826 2395 4830
rect 2495 4826 2499 4830
rect 2527 4826 2531 4830
rect 2663 4826 2667 4830
rect 2671 4826 2675 4830
rect 2807 4826 2811 4830
rect 2847 4826 2851 4830
rect 2951 4826 2955 4830
rect 3015 4826 3019 4830
rect 3095 4826 3099 4830
rect 3183 4826 3187 4830
rect 3239 4826 3243 4830
rect 3351 4826 3355 4830
rect 3383 4826 3387 4830
rect 3527 4826 3531 4830
rect 3679 4826 3683 4830
rect 3799 4826 3803 4830
rect 111 4786 115 4790
rect 131 4786 135 4790
rect 267 4786 271 4790
rect 387 4786 391 4790
rect 403 4786 407 4790
rect 539 4786 543 4790
rect 675 4786 679 4790
rect 707 4786 711 4790
rect 1059 4786 1063 4790
rect 1435 4786 1439 4790
rect 1787 4786 1791 4790
rect 1935 4786 1939 4790
rect 3839 4782 3843 4786
rect 4703 4782 4707 4786
rect 4855 4782 4859 4786
rect 4991 4782 4995 4786
rect 5015 4782 5019 4786
rect 5127 4782 5131 4786
rect 5183 4782 5187 4786
rect 5263 4782 5267 4786
rect 5351 4782 5355 4786
rect 5399 4782 5403 4786
rect 5527 4782 5531 4786
rect 5535 4782 5539 4786
rect 5663 4782 5667 4786
rect 1975 4706 1979 4710
rect 1995 4706 1999 4710
rect 2131 4706 2135 4710
rect 2267 4706 2271 4710
rect 2363 4706 2367 4710
rect 2427 4706 2431 4710
rect 2499 4706 2503 4710
rect 2587 4706 2591 4710
rect 2635 4706 2639 4710
rect 2747 4706 2751 4710
rect 2779 4706 2783 4710
rect 2907 4706 2911 4710
rect 2923 4706 2927 4710
rect 3067 4706 3071 4710
rect 3211 4706 3215 4710
rect 3235 4706 3239 4710
rect 3355 4706 3359 4710
rect 3499 4706 3503 4710
rect 3799 4706 3803 4710
rect 111 4670 115 4674
rect 159 4670 163 4674
rect 295 4670 299 4674
rect 431 4670 435 4674
rect 567 4670 571 4674
rect 703 4670 707 4674
rect 1935 4670 1939 4674
rect 3839 4650 3843 4654
rect 4715 4650 4719 4654
rect 4827 4650 4831 4654
rect 4859 4650 4863 4654
rect 4963 4650 4967 4654
rect 5011 4650 5015 4654
rect 5099 4650 5103 4654
rect 5171 4650 5175 4654
rect 5235 4650 5239 4654
rect 5339 4650 5343 4654
rect 5371 4650 5375 4654
rect 5507 4650 5511 4654
rect 5515 4650 5519 4654
rect 5663 4650 5667 4654
rect 1975 4594 1979 4598
rect 2023 4594 2027 4598
rect 2159 4594 2163 4598
rect 2175 4594 2179 4598
rect 2295 4594 2299 4598
rect 2351 4594 2355 4598
rect 2455 4594 2459 4598
rect 2527 4594 2531 4598
rect 2615 4594 2619 4598
rect 2695 4594 2699 4598
rect 2775 4594 2779 4598
rect 2871 4594 2875 4598
rect 2935 4594 2939 4598
rect 3047 4594 3051 4598
rect 3095 4594 3099 4598
rect 3263 4594 3267 4598
rect 3799 4594 3803 4598
rect 111 4546 115 4550
rect 131 4546 135 4550
rect 267 4546 271 4550
rect 299 4546 303 4550
rect 403 4546 407 4550
rect 491 4546 495 4550
rect 539 4546 543 4550
rect 675 4546 679 4550
rect 691 4546 695 4550
rect 907 4546 911 4550
rect 1123 4546 1127 4550
rect 1347 4546 1351 4550
rect 1579 4546 1583 4550
rect 1787 4546 1791 4550
rect 1935 4546 1939 4550
rect 3839 4514 3843 4518
rect 3887 4514 3891 4518
rect 4063 4514 4067 4518
rect 4279 4514 4283 4518
rect 4503 4514 4507 4518
rect 4743 4514 4747 4518
rect 4751 4514 4755 4518
rect 4887 4514 4891 4518
rect 5007 4514 5011 4518
rect 5039 4514 5043 4518
rect 5199 4514 5203 4518
rect 5271 4514 5275 4518
rect 5367 4514 5371 4518
rect 5543 4514 5547 4518
rect 5663 4514 5667 4518
rect 1975 4442 1979 4446
rect 1995 4442 1999 4446
rect 2147 4442 2151 4446
rect 2323 4442 2327 4446
rect 2499 4442 2503 4446
rect 2571 4442 2575 4446
rect 2667 4442 2671 4446
rect 2843 4442 2847 4446
rect 3019 4442 3023 4446
rect 3123 4442 3127 4446
rect 3651 4442 3655 4446
rect 3799 4442 3803 4446
rect 111 4434 115 4438
rect 327 4434 331 4438
rect 519 4434 523 4438
rect 559 4434 563 4438
rect 719 4434 723 4438
rect 887 4434 891 4438
rect 935 4434 939 4438
rect 1063 4434 1067 4438
rect 1151 4434 1155 4438
rect 1247 4434 1251 4438
rect 1375 4434 1379 4438
rect 1439 4434 1443 4438
rect 1607 4434 1611 4438
rect 1631 4434 1635 4438
rect 1815 4434 1819 4438
rect 1935 4434 1939 4438
rect 3839 4402 3843 4406
rect 3859 4402 3863 4406
rect 3995 4402 3999 4406
rect 4035 4402 4039 4406
rect 4131 4402 4135 4406
rect 4251 4402 4255 4406
rect 4267 4402 4271 4406
rect 4403 4402 4407 4406
rect 4475 4402 4479 4406
rect 4587 4402 4591 4406
rect 4723 4402 4727 4406
rect 4795 4402 4799 4406
rect 4979 4402 4983 4406
rect 5027 4402 5031 4406
rect 5243 4402 5247 4406
rect 5275 4402 5279 4406
rect 5515 4402 5519 4406
rect 5663 4402 5667 4406
rect 1975 4326 1979 4330
rect 2399 4326 2403 4330
rect 2599 4326 2603 4330
rect 2791 4326 2795 4330
rect 2983 4326 2987 4330
rect 3151 4326 3155 4330
rect 3167 4326 3171 4330
rect 3343 4326 3347 4330
rect 3519 4326 3523 4330
rect 3679 4326 3683 4330
rect 3799 4326 3803 4330
rect 111 4314 115 4318
rect 531 4314 535 4318
rect 691 4314 695 4318
rect 747 4314 751 4318
rect 859 4314 863 4318
rect 883 4314 887 4318
rect 1019 4314 1023 4318
rect 1035 4314 1039 4318
rect 1155 4314 1159 4318
rect 1219 4314 1223 4318
rect 1291 4314 1295 4318
rect 1411 4314 1415 4318
rect 1427 4314 1431 4318
rect 1563 4314 1567 4318
rect 1603 4314 1607 4318
rect 1699 4314 1703 4318
rect 1787 4314 1791 4318
rect 1935 4314 1939 4318
rect 3839 4290 3843 4294
rect 3887 4290 3891 4294
rect 4023 4290 4027 4294
rect 4047 4290 4051 4294
rect 4159 4290 4163 4294
rect 4223 4290 4227 4294
rect 4295 4290 4299 4294
rect 4431 4290 4435 4294
rect 4615 4290 4619 4294
rect 4679 4290 4683 4294
rect 4823 4290 4827 4294
rect 4959 4290 4963 4294
rect 5055 4290 5059 4294
rect 5255 4290 5259 4294
rect 5303 4290 5307 4294
rect 5543 4290 5547 4294
rect 5663 4290 5667 4294
rect 1975 4202 1979 4206
rect 2371 4202 2375 4206
rect 2571 4202 2575 4206
rect 2611 4202 2615 4206
rect 2763 4202 2767 4206
rect 2835 4202 2839 4206
rect 2955 4202 2959 4206
rect 3051 4202 3055 4206
rect 3139 4202 3143 4206
rect 3259 4202 3263 4206
rect 3315 4202 3319 4206
rect 3467 4202 3471 4206
rect 3491 4202 3495 4206
rect 3651 4202 3655 4206
rect 3799 4202 3803 4206
rect 111 4190 115 4194
rect 727 4190 731 4194
rect 775 4190 779 4194
rect 863 4190 867 4194
rect 911 4190 915 4194
rect 999 4190 1003 4194
rect 1047 4190 1051 4194
rect 1135 4190 1139 4194
rect 1183 4190 1187 4194
rect 1271 4190 1275 4194
rect 1319 4190 1323 4194
rect 1407 4190 1411 4194
rect 1455 4190 1459 4194
rect 1543 4190 1547 4194
rect 1591 4190 1595 4194
rect 1679 4190 1683 4194
rect 1727 4190 1731 4194
rect 1815 4190 1819 4194
rect 1935 4190 1939 4194
rect 3839 4094 3843 4098
rect 4019 4094 4023 4098
rect 4195 4094 4199 4098
rect 4403 4094 4407 4098
rect 4651 4094 4655 4098
rect 4931 4094 4935 4098
rect 5227 4094 5231 4098
rect 5515 4094 5519 4098
rect 5663 4094 5667 4098
rect 1975 4086 1979 4090
rect 2375 4086 2379 4090
rect 2399 4086 2403 4090
rect 2623 4086 2627 4090
rect 2639 4086 2643 4090
rect 2855 4086 2859 4090
rect 2863 4086 2867 4090
rect 3071 4086 3075 4090
rect 3079 4086 3083 4090
rect 3279 4086 3283 4090
rect 3287 4086 3291 4090
rect 3487 4086 3491 4090
rect 3495 4086 3499 4090
rect 3679 4086 3683 4090
rect 3799 4086 3803 4090
rect 111 4066 115 4070
rect 627 4066 631 4070
rect 699 4066 703 4070
rect 763 4066 767 4070
rect 835 4066 839 4070
rect 899 4066 903 4070
rect 971 4066 975 4070
rect 1035 4066 1039 4070
rect 1107 4066 1111 4070
rect 1171 4066 1175 4070
rect 1243 4066 1247 4070
rect 1307 4066 1311 4070
rect 1379 4066 1383 4070
rect 1443 4066 1447 4070
rect 1515 4066 1519 4070
rect 1579 4066 1583 4070
rect 1651 4066 1655 4070
rect 1715 4066 1719 4070
rect 1787 4066 1791 4070
rect 1935 4066 1939 4070
rect 1975 3974 1979 3978
rect 2323 3974 2327 3978
rect 2347 3974 2351 3978
rect 2571 3974 2575 3978
rect 2595 3974 2599 3978
rect 2803 3974 2807 3978
rect 2827 3974 2831 3978
rect 3027 3974 3031 3978
rect 3043 3974 3047 3978
rect 3243 3974 3247 3978
rect 3251 3974 3255 3978
rect 3459 3974 3463 3978
rect 3651 3974 3655 3978
rect 3799 3974 3803 3978
rect 3839 3974 3843 3978
rect 4183 3974 4187 3978
rect 4319 3974 4323 3978
rect 4455 3974 4459 3978
rect 4591 3974 4595 3978
rect 4727 3974 4731 3978
rect 4863 3974 4867 3978
rect 4999 3974 5003 3978
rect 5135 3974 5139 3978
rect 5271 3974 5275 3978
rect 5407 3974 5411 3978
rect 5543 3974 5547 3978
rect 5663 3974 5667 3978
rect 111 3942 115 3946
rect 599 3942 603 3946
rect 655 3942 659 3946
rect 743 3942 747 3946
rect 791 3942 795 3946
rect 895 3942 899 3946
rect 927 3942 931 3946
rect 1047 3942 1051 3946
rect 1063 3942 1067 3946
rect 1199 3942 1203 3946
rect 1335 3942 1339 3946
rect 1359 3942 1363 3946
rect 1471 3942 1475 3946
rect 1519 3942 1523 3946
rect 1607 3942 1611 3946
rect 1679 3942 1683 3946
rect 1743 3942 1747 3946
rect 1935 3942 1939 3946
rect 1975 3858 1979 3862
rect 2239 3858 2243 3862
rect 2351 3858 2355 3862
rect 2479 3858 2483 3862
rect 2599 3858 2603 3862
rect 2703 3858 2707 3862
rect 2831 3858 2835 3862
rect 2919 3858 2923 3862
rect 3055 3858 3059 3862
rect 3119 3858 3123 3862
rect 3271 3858 3275 3862
rect 3311 3858 3315 3862
rect 3487 3858 3491 3862
rect 3503 3858 3507 3862
rect 3679 3858 3683 3862
rect 3799 3858 3803 3862
rect 3839 3830 3843 3834
rect 4139 3830 4143 3834
rect 4155 3830 4159 3834
rect 4291 3830 4295 3834
rect 4323 3830 4327 3834
rect 4427 3830 4431 3834
rect 4531 3830 4535 3834
rect 4563 3830 4567 3834
rect 4699 3830 4703 3834
rect 4763 3830 4767 3834
rect 4835 3830 4839 3834
rect 4971 3830 4975 3834
rect 5011 3830 5015 3834
rect 5107 3830 5111 3834
rect 5243 3830 5247 3834
rect 5275 3830 5279 3834
rect 5379 3830 5383 3834
rect 5515 3830 5519 3834
rect 5663 3830 5667 3834
rect 111 3822 115 3826
rect 427 3822 431 3826
rect 571 3822 575 3826
rect 587 3822 591 3826
rect 715 3822 719 3826
rect 755 3822 759 3826
rect 867 3822 871 3826
rect 923 3822 927 3826
rect 1019 3822 1023 3826
rect 1099 3822 1103 3826
rect 1171 3822 1175 3826
rect 1275 3822 1279 3826
rect 1331 3822 1335 3826
rect 1459 3822 1463 3826
rect 1491 3822 1495 3826
rect 1643 3822 1647 3826
rect 1651 3822 1655 3826
rect 1935 3822 1939 3826
rect 1975 3738 1979 3742
rect 2211 3738 2215 3742
rect 2227 3738 2231 3742
rect 2451 3738 2455 3742
rect 2667 3738 2671 3742
rect 2675 3738 2679 3742
rect 2875 3738 2879 3742
rect 2891 3738 2895 3742
rect 3075 3738 3079 3742
rect 3091 3738 3095 3742
rect 3275 3738 3279 3742
rect 3283 3738 3287 3742
rect 3475 3738 3479 3742
rect 3651 3738 3655 3742
rect 3799 3738 3803 3742
rect 111 3698 115 3702
rect 327 3698 331 3702
rect 455 3698 459 3702
rect 495 3698 499 3702
rect 615 3698 619 3702
rect 679 3698 683 3702
rect 783 3698 787 3702
rect 863 3698 867 3702
rect 951 3698 955 3702
rect 1055 3698 1059 3702
rect 1127 3698 1131 3702
rect 1255 3698 1259 3702
rect 1303 3698 1307 3702
rect 1455 3698 1459 3702
rect 1487 3698 1491 3702
rect 1655 3698 1659 3702
rect 1671 3698 1675 3702
rect 1935 3698 1939 3702
rect 3839 3698 3843 3702
rect 4167 3698 4171 3702
rect 4303 3698 4307 3702
rect 4351 3698 4355 3702
rect 4479 3698 4483 3702
rect 4559 3698 4563 3702
rect 4671 3698 4675 3702
rect 4791 3698 4795 3702
rect 4879 3698 4883 3702
rect 5039 3698 5043 3702
rect 5103 3698 5107 3702
rect 5303 3698 5307 3702
rect 5335 3698 5339 3702
rect 5543 3698 5547 3702
rect 5663 3698 5667 3702
rect 1975 3622 1979 3626
rect 2135 3622 2139 3626
rect 2255 3622 2259 3626
rect 2311 3622 2315 3626
rect 2479 3622 2483 3626
rect 2647 3622 2651 3626
rect 2695 3622 2699 3626
rect 2807 3622 2811 3626
rect 2903 3622 2907 3626
rect 2967 3622 2971 3626
rect 3103 3622 3107 3626
rect 3135 3622 3139 3626
rect 3303 3622 3307 3626
rect 3503 3622 3507 3626
rect 3799 3622 3803 3626
rect 111 3566 115 3570
rect 203 3566 207 3570
rect 299 3566 303 3570
rect 379 3566 383 3570
rect 467 3566 471 3570
rect 563 3566 567 3570
rect 651 3566 655 3570
rect 755 3566 759 3570
rect 835 3566 839 3570
rect 955 3566 959 3570
rect 1027 3566 1031 3570
rect 1163 3566 1167 3570
rect 1227 3566 1231 3570
rect 1379 3566 1383 3570
rect 1427 3566 1431 3570
rect 1595 3566 1599 3570
rect 1627 3566 1631 3570
rect 1935 3566 1939 3570
rect 3839 3558 3843 3562
rect 4275 3558 4279 3562
rect 4451 3558 4455 3562
rect 4555 3558 4559 3562
rect 4643 3558 4647 3562
rect 4699 3558 4703 3562
rect 4851 3558 4855 3562
rect 5011 3558 5015 3562
rect 5075 3558 5079 3562
rect 5179 3558 5183 3562
rect 5307 3558 5311 3562
rect 5355 3558 5359 3562
rect 5515 3558 5519 3562
rect 5663 3558 5667 3562
rect 1975 3486 1979 3490
rect 2035 3486 2039 3490
rect 2107 3486 2111 3490
rect 2187 3486 2191 3490
rect 2283 3486 2287 3490
rect 2339 3486 2343 3490
rect 2451 3486 2455 3490
rect 2491 3486 2495 3490
rect 2619 3486 2623 3490
rect 2643 3486 2647 3490
rect 2779 3486 2783 3490
rect 2795 3486 2799 3490
rect 2939 3486 2943 3490
rect 2947 3486 2951 3490
rect 3099 3486 3103 3490
rect 3107 3486 3111 3490
rect 3275 3486 3279 3490
rect 3799 3486 3803 3490
rect 111 3434 115 3438
rect 231 3434 235 3438
rect 255 3434 259 3438
rect 407 3434 411 3438
rect 471 3434 475 3438
rect 591 3434 595 3438
rect 695 3434 699 3438
rect 783 3434 787 3438
rect 919 3434 923 3438
rect 983 3434 987 3438
rect 1143 3434 1147 3438
rect 1191 3434 1195 3438
rect 1367 3434 1371 3438
rect 1407 3434 1411 3438
rect 1591 3434 1595 3438
rect 1623 3434 1627 3438
rect 1935 3434 1939 3438
rect 3839 3434 3843 3438
rect 4583 3434 4587 3438
rect 4727 3434 4731 3438
rect 4879 3434 4883 3438
rect 4903 3434 4907 3438
rect 5039 3434 5043 3438
rect 5175 3434 5179 3438
rect 5207 3434 5211 3438
rect 5311 3434 5315 3438
rect 5383 3434 5387 3438
rect 5447 3434 5451 3438
rect 5543 3434 5547 3438
rect 5663 3434 5667 3438
rect 1975 3362 1979 3366
rect 2023 3362 2027 3366
rect 2063 3362 2067 3366
rect 2191 3362 2195 3366
rect 2215 3362 2219 3366
rect 2367 3362 2371 3366
rect 2375 3362 2379 3366
rect 2519 3362 2523 3366
rect 2551 3362 2555 3366
rect 2671 3362 2675 3366
rect 2727 3362 2731 3366
rect 2823 3362 2827 3366
rect 2895 3362 2899 3366
rect 2975 3362 2979 3366
rect 3071 3362 3075 3366
rect 3127 3362 3131 3366
rect 3247 3362 3251 3366
rect 3799 3362 3803 3366
rect 3839 3322 3843 3326
rect 4699 3322 4703 3326
rect 4835 3322 4839 3326
rect 4875 3322 4879 3326
rect 4971 3322 4975 3326
rect 5011 3322 5015 3326
rect 5107 3322 5111 3326
rect 5147 3322 5151 3326
rect 5243 3322 5247 3326
rect 5283 3322 5287 3326
rect 5379 3322 5383 3326
rect 5419 3322 5423 3326
rect 5515 3322 5519 3326
rect 5663 3322 5667 3326
rect 111 3306 115 3310
rect 211 3306 215 3310
rect 227 3306 231 3310
rect 419 3306 423 3310
rect 443 3306 447 3310
rect 635 3306 639 3310
rect 667 3306 671 3310
rect 851 3306 855 3310
rect 891 3306 895 3310
rect 1075 3306 1079 3310
rect 1115 3306 1119 3310
rect 1299 3306 1303 3310
rect 1339 3306 1343 3310
rect 1523 3306 1527 3310
rect 1563 3306 1567 3310
rect 1935 3306 1939 3310
rect 1975 3246 1979 3250
rect 1995 3246 1999 3250
rect 2163 3246 2167 3250
rect 2211 3246 2215 3250
rect 2347 3246 2351 3250
rect 2435 3246 2439 3250
rect 2523 3246 2527 3250
rect 2651 3246 2655 3250
rect 2699 3246 2703 3250
rect 2851 3246 2855 3250
rect 2867 3246 2871 3250
rect 3043 3246 3047 3250
rect 3051 3246 3055 3250
rect 3219 3246 3223 3250
rect 3251 3246 3255 3250
rect 3451 3246 3455 3250
rect 3799 3246 3803 3250
rect 3839 3202 3843 3206
rect 4567 3202 4571 3206
rect 4727 3202 4731 3206
rect 4743 3202 4747 3206
rect 4863 3202 4867 3206
rect 4935 3202 4939 3206
rect 4999 3202 5003 3206
rect 5135 3202 5139 3206
rect 5271 3202 5275 3206
rect 5351 3202 5355 3206
rect 5407 3202 5411 3206
rect 5543 3202 5547 3206
rect 5663 3202 5667 3206
rect 111 3178 115 3182
rect 239 3178 243 3182
rect 303 3178 307 3182
rect 447 3178 451 3182
rect 543 3178 547 3182
rect 663 3178 667 3182
rect 783 3178 787 3182
rect 879 3178 883 3182
rect 1023 3178 1027 3182
rect 1103 3178 1107 3182
rect 1263 3178 1267 3182
rect 1327 3178 1331 3182
rect 1511 3178 1515 3182
rect 1551 3178 1555 3182
rect 1935 3178 1939 3182
rect 1975 3134 1979 3138
rect 2023 3134 2027 3138
rect 2239 3134 2243 3138
rect 2327 3134 2331 3138
rect 2463 3134 2467 3138
rect 2631 3134 2635 3138
rect 2679 3134 2683 3138
rect 2879 3134 2883 3138
rect 2911 3134 2915 3138
rect 3079 3134 3083 3138
rect 3175 3134 3179 3138
rect 3279 3134 3283 3138
rect 3439 3134 3443 3138
rect 3479 3134 3483 3138
rect 3679 3134 3683 3138
rect 3799 3134 3803 3138
rect 111 3066 115 3070
rect 275 3066 279 3070
rect 355 3066 359 3070
rect 515 3066 519 3070
rect 627 3066 631 3070
rect 755 3066 759 3070
rect 883 3066 887 3070
rect 995 3066 999 3070
rect 1123 3066 1127 3070
rect 1235 3066 1239 3070
rect 1355 3066 1359 3070
rect 1483 3066 1487 3070
rect 1579 3066 1583 3070
rect 1787 3066 1791 3070
rect 1935 3066 1939 3070
rect 3839 3086 3843 3090
rect 4307 3086 4311 3090
rect 4483 3086 4487 3090
rect 4539 3086 4543 3090
rect 4675 3086 4679 3090
rect 4715 3086 4719 3090
rect 4875 3086 4879 3090
rect 4907 3086 4911 3090
rect 5091 3086 5095 3090
rect 5107 3086 5111 3090
rect 5315 3086 5319 3090
rect 5323 3086 5327 3090
rect 5515 3086 5519 3090
rect 5663 3086 5667 3090
rect 1975 3014 1979 3018
rect 1995 3014 1999 3018
rect 2299 3014 2303 3018
rect 2603 3014 2607 3018
rect 2883 3014 2887 3018
rect 3107 3014 3111 3018
rect 3147 3014 3151 3018
rect 3243 3014 3247 3018
rect 3379 3014 3383 3018
rect 3411 3014 3415 3018
rect 3515 3014 3519 3018
rect 3651 3014 3655 3018
rect 3799 3014 3803 3018
rect 111 2954 115 2958
rect 343 2954 347 2958
rect 383 2954 387 2958
rect 551 2954 555 2958
rect 655 2954 659 2958
rect 759 2954 763 2958
rect 911 2954 915 2958
rect 951 2954 955 2958
rect 1135 2954 1139 2958
rect 1151 2954 1155 2958
rect 1311 2954 1315 2958
rect 1383 2954 1387 2958
rect 1487 2954 1491 2958
rect 1607 2954 1611 2958
rect 1663 2954 1667 2958
rect 1815 2954 1819 2958
rect 1935 2954 1939 2958
rect 3839 2970 3843 2974
rect 3887 2970 3891 2974
rect 4023 2970 4027 2974
rect 4175 2970 4179 2974
rect 4335 2970 4339 2974
rect 4391 2970 4395 2974
rect 4511 2970 4515 2974
rect 4639 2970 4643 2974
rect 4703 2970 4707 2974
rect 4903 2970 4907 2974
rect 4919 2970 4923 2974
rect 5119 2970 5123 2974
rect 5223 2970 5227 2974
rect 5343 2970 5347 2974
rect 5527 2970 5531 2974
rect 5543 2970 5547 2974
rect 5663 2970 5667 2974
rect 111 2830 115 2834
rect 315 2830 319 2834
rect 363 2830 367 2834
rect 523 2830 527 2834
rect 563 2830 567 2834
rect 731 2830 735 2834
rect 755 2830 759 2834
rect 923 2830 927 2834
rect 939 2830 943 2834
rect 1107 2830 1111 2834
rect 1115 2830 1119 2834
rect 1283 2830 1287 2834
rect 1451 2830 1455 2834
rect 1459 2830 1463 2834
rect 1619 2830 1623 2834
rect 1635 2830 1639 2834
rect 1787 2830 1791 2834
rect 1935 2830 1939 2834
rect 111 2714 115 2718
rect 391 2714 395 2718
rect 447 2714 451 2718
rect 591 2714 595 2718
rect 615 2714 619 2718
rect 775 2714 779 2718
rect 783 2714 787 2718
rect 935 2714 939 2718
rect 967 2714 971 2718
rect 1087 2714 1091 2718
rect 1143 2714 1147 2718
rect 1239 2714 1243 2718
rect 1311 2714 1315 2718
rect 1383 2714 1387 2718
rect 1479 2714 1483 2718
rect 1535 2714 1539 2718
rect 1647 2714 1651 2718
rect 1679 2714 1683 2718
rect 1815 2714 1819 2718
rect 1935 2714 1939 2718
rect 3839 2858 3843 2862
rect 3859 2858 3863 2862
rect 3995 2858 3999 2862
rect 4131 2858 4135 2862
rect 4147 2858 4151 2862
rect 4267 2858 4271 2862
rect 4363 2858 4367 2862
rect 4403 2858 4407 2862
rect 4539 2858 4543 2862
rect 4611 2858 4615 2862
rect 4675 2858 4679 2862
rect 4811 2858 4815 2862
rect 4891 2858 4895 2862
rect 5195 2858 5199 2862
rect 5499 2858 5503 2862
rect 5663 2858 5667 2862
rect 3839 2730 3843 2734
rect 3887 2730 3891 2734
rect 4023 2730 4027 2734
rect 4159 2730 4163 2734
rect 4295 2730 4299 2734
rect 4431 2730 4435 2734
rect 4567 2730 4571 2734
rect 4703 2730 4707 2734
rect 4711 2730 4715 2734
rect 4839 2730 4843 2734
rect 4879 2730 4883 2734
rect 5063 2730 5067 2734
rect 5255 2730 5259 2734
rect 5447 2730 5451 2734
rect 5663 2730 5667 2734
rect 1975 2634 1979 2638
rect 3135 2634 3139 2638
rect 3271 2634 3275 2638
rect 3407 2634 3411 2638
rect 3543 2634 3547 2638
rect 3679 2634 3683 2638
rect 3799 2634 3803 2638
rect 111 2598 115 2602
rect 235 2598 239 2602
rect 419 2598 423 2602
rect 435 2598 439 2602
rect 587 2598 591 2602
rect 627 2598 631 2602
rect 747 2598 751 2602
rect 811 2598 815 2602
rect 907 2598 911 2602
rect 987 2598 991 2602
rect 1059 2598 1063 2602
rect 1155 2598 1159 2602
rect 1211 2598 1215 2602
rect 1323 2598 1327 2602
rect 1355 2598 1359 2602
rect 1483 2598 1487 2602
rect 1507 2598 1511 2602
rect 1643 2598 1647 2602
rect 1651 2598 1655 2602
rect 1787 2598 1791 2602
rect 1935 2598 1939 2602
rect 3839 2602 3843 2606
rect 3859 2602 3863 2606
rect 3995 2602 3999 2606
rect 4131 2602 4135 2606
rect 4179 2602 4183 2606
rect 4267 2602 4271 2606
rect 4395 2602 4399 2606
rect 4403 2602 4407 2606
rect 4539 2602 4543 2606
rect 4643 2602 4647 2606
rect 4683 2602 4687 2606
rect 4851 2602 4855 2606
rect 4907 2602 4911 2606
rect 5035 2602 5039 2606
rect 5187 2602 5191 2606
rect 5227 2602 5231 2606
rect 5419 2602 5423 2606
rect 5467 2602 5471 2606
rect 5663 2602 5667 2606
rect 1975 2522 1979 2526
rect 1995 2522 1999 2526
rect 2251 2522 2255 2526
rect 2523 2522 2527 2526
rect 2771 2522 2775 2526
rect 3003 2522 3007 2526
rect 3227 2522 3231 2526
rect 3243 2522 3247 2526
rect 3379 2522 3383 2526
rect 3451 2522 3455 2526
rect 3515 2522 3519 2526
rect 3651 2522 3655 2526
rect 3799 2522 3803 2526
rect 111 2478 115 2482
rect 223 2478 227 2482
rect 263 2478 267 2482
rect 423 2478 427 2482
rect 463 2478 467 2482
rect 623 2478 627 2482
rect 655 2478 659 2482
rect 815 2478 819 2482
rect 839 2478 843 2482
rect 1015 2478 1019 2482
rect 1183 2478 1187 2482
rect 1215 2478 1219 2482
rect 1351 2478 1355 2482
rect 1511 2478 1515 2482
rect 1671 2478 1675 2482
rect 1815 2478 1819 2482
rect 1935 2478 1939 2482
rect 3839 2490 3843 2494
rect 4207 2490 4211 2494
rect 4423 2490 4427 2494
rect 4535 2490 4539 2494
rect 4671 2490 4675 2494
rect 4759 2490 4763 2494
rect 4935 2490 4939 2494
rect 4983 2490 4987 2494
rect 5215 2490 5219 2494
rect 5447 2490 5451 2494
rect 5495 2490 5499 2494
rect 5663 2490 5667 2494
rect 1975 2410 1979 2414
rect 2023 2410 2027 2414
rect 2055 2410 2059 2414
rect 2215 2410 2219 2414
rect 2279 2410 2283 2414
rect 2375 2410 2379 2414
rect 2543 2410 2547 2414
rect 2551 2410 2555 2414
rect 2711 2410 2715 2414
rect 2799 2410 2803 2414
rect 2871 2410 2875 2414
rect 3031 2410 3035 2414
rect 3191 2410 3195 2414
rect 3255 2410 3259 2414
rect 3359 2410 3363 2414
rect 3479 2410 3483 2414
rect 3527 2410 3531 2414
rect 3679 2410 3683 2414
rect 3799 2410 3803 2414
rect 3839 2378 3843 2382
rect 4507 2378 4511 2382
rect 4707 2378 4711 2382
rect 4731 2378 4735 2382
rect 4867 2378 4871 2382
rect 4955 2378 4959 2382
rect 5027 2378 5031 2382
rect 5187 2378 5191 2382
rect 5347 2378 5351 2382
rect 5419 2378 5423 2382
rect 5515 2378 5519 2382
rect 5663 2378 5667 2382
rect 111 2354 115 2358
rect 131 2354 135 2358
rect 195 2354 199 2358
rect 291 2354 295 2358
rect 395 2354 399 2358
rect 483 2354 487 2358
rect 595 2354 599 2358
rect 675 2354 679 2358
rect 787 2354 791 2358
rect 867 2354 871 2358
rect 987 2354 991 2358
rect 1187 2354 1191 2358
rect 1935 2354 1939 2358
rect 1975 2290 1979 2294
rect 2027 2290 2031 2294
rect 2139 2290 2143 2294
rect 2187 2290 2191 2294
rect 2275 2290 2279 2294
rect 2347 2290 2351 2294
rect 2411 2290 2415 2294
rect 2515 2290 2519 2294
rect 2547 2290 2551 2294
rect 2683 2290 2687 2294
rect 2819 2290 2823 2294
rect 2843 2290 2847 2294
rect 2955 2290 2959 2294
rect 3003 2290 3007 2294
rect 3091 2290 3095 2294
rect 3163 2290 3167 2294
rect 3227 2290 3231 2294
rect 3331 2290 3335 2294
rect 3363 2290 3367 2294
rect 3499 2290 3503 2294
rect 3799 2290 3803 2294
rect 111 2242 115 2246
rect 159 2242 163 2246
rect 295 2242 299 2246
rect 319 2242 323 2246
rect 439 2242 443 2246
rect 511 2242 515 2246
rect 591 2242 595 2246
rect 703 2242 707 2246
rect 743 2242 747 2246
rect 895 2242 899 2246
rect 1935 2242 1939 2246
rect 3839 2254 3843 2258
rect 4735 2254 4739 2258
rect 4887 2254 4891 2258
rect 4895 2254 4899 2258
rect 5047 2254 5051 2258
rect 5055 2254 5059 2258
rect 5215 2254 5219 2258
rect 5375 2254 5379 2258
rect 5391 2254 5395 2258
rect 5543 2254 5547 2258
rect 5663 2254 5667 2258
rect 1975 2174 1979 2178
rect 2023 2174 2027 2178
rect 2159 2174 2163 2178
rect 2167 2174 2171 2178
rect 2295 2174 2299 2178
rect 2303 2174 2307 2178
rect 2431 2174 2435 2178
rect 2439 2174 2443 2178
rect 2567 2174 2571 2178
rect 2575 2174 2579 2178
rect 2703 2174 2707 2178
rect 2711 2174 2715 2178
rect 2839 2174 2843 2178
rect 2847 2174 2851 2178
rect 2975 2174 2979 2178
rect 2983 2174 2987 2178
rect 3111 2174 3115 2178
rect 3119 2174 3123 2178
rect 3247 2174 3251 2178
rect 3255 2174 3259 2178
rect 3391 2174 3395 2178
rect 3799 2174 3803 2178
rect 111 2130 115 2134
rect 131 2130 135 2134
rect 267 2130 271 2134
rect 331 2130 335 2134
rect 411 2130 415 2134
rect 555 2130 559 2134
rect 563 2130 567 2134
rect 715 2130 719 2134
rect 779 2130 783 2134
rect 1011 2130 1015 2134
rect 3839 2134 3843 2138
rect 1935 2130 1939 2134
rect 4707 2134 4711 2138
rect 4787 2134 4791 2138
rect 4859 2134 4863 2138
rect 4923 2134 4927 2138
rect 5019 2134 5023 2138
rect 5067 2134 5071 2138
rect 5187 2134 5191 2138
rect 5219 2134 5223 2138
rect 5363 2134 5367 2138
rect 5379 2134 5383 2138
rect 5515 2134 5519 2138
rect 5663 2134 5667 2138
rect 1975 2054 1979 2058
rect 1995 2054 1999 2058
rect 2131 2054 2135 2058
rect 2267 2054 2271 2058
rect 2403 2054 2407 2058
rect 2539 2054 2543 2058
rect 2675 2054 2679 2058
rect 2811 2054 2815 2058
rect 2947 2054 2951 2058
rect 3083 2054 3087 2058
rect 3091 2054 3095 2058
rect 3219 2054 3223 2058
rect 3243 2054 3247 2058
rect 3395 2054 3399 2058
rect 3799 2054 3803 2058
rect 111 2014 115 2018
rect 159 2014 163 2018
rect 359 2014 363 2018
rect 463 2014 467 2018
rect 583 2014 587 2018
rect 799 2014 803 2018
rect 807 2014 811 2018
rect 1039 2014 1043 2018
rect 1143 2014 1147 2018
rect 1487 2014 1491 2018
rect 1815 2014 1819 2018
rect 1935 2014 1939 2018
rect 3839 2018 3843 2022
rect 4815 2018 4819 2022
rect 4863 2018 4867 2022
rect 4951 2018 4955 2022
rect 4999 2018 5003 2022
rect 5095 2018 5099 2022
rect 5135 2018 5139 2022
rect 5247 2018 5251 2022
rect 5271 2018 5275 2022
rect 5407 2018 5411 2022
rect 5543 2018 5547 2022
rect 5663 2018 5667 2022
rect 1975 1934 1979 1938
rect 2023 1934 2027 1938
rect 2159 1934 2163 1938
rect 2295 1934 2299 1938
rect 2431 1934 2435 1938
rect 2527 1934 2531 1938
rect 2567 1934 2571 1938
rect 2663 1934 2667 1938
rect 2703 1934 2707 1938
rect 2799 1934 2803 1938
rect 2839 1934 2843 1938
rect 2935 1934 2939 1938
rect 2975 1934 2979 1938
rect 3071 1934 3075 1938
rect 3119 1934 3123 1938
rect 3207 1934 3211 1938
rect 3271 1934 3275 1938
rect 3351 1934 3355 1938
rect 3423 1934 3427 1938
rect 3799 1934 3803 1938
rect 111 1902 115 1906
rect 131 1902 135 1906
rect 195 1902 199 1906
rect 435 1902 439 1906
rect 451 1902 455 1906
rect 699 1902 703 1906
rect 771 1902 775 1906
rect 931 1902 935 1906
rect 1115 1902 1119 1906
rect 1155 1902 1159 1906
rect 1371 1902 1375 1906
rect 1459 1902 1463 1906
rect 1587 1902 1591 1906
rect 1787 1902 1791 1906
rect 1935 1902 1939 1906
rect 3839 1902 3843 1906
rect 4683 1902 4687 1906
rect 4835 1902 4839 1906
rect 4843 1902 4847 1906
rect 4971 1902 4975 1906
rect 5011 1902 5015 1906
rect 5107 1902 5111 1906
rect 5179 1902 5183 1906
rect 5243 1902 5247 1906
rect 5355 1902 5359 1906
rect 5379 1902 5383 1906
rect 5515 1902 5519 1906
rect 5663 1902 5667 1906
rect 1975 1822 1979 1826
rect 2443 1822 2447 1826
rect 2499 1822 2503 1826
rect 2587 1822 2591 1826
rect 2635 1822 2639 1826
rect 2739 1822 2743 1826
rect 2771 1822 2775 1826
rect 2891 1822 2895 1826
rect 2907 1822 2911 1826
rect 3043 1822 3047 1826
rect 3179 1822 3183 1826
rect 3195 1822 3199 1826
rect 3323 1822 3327 1826
rect 3799 1822 3803 1826
rect 111 1786 115 1790
rect 223 1786 227 1790
rect 231 1786 235 1790
rect 447 1786 451 1790
rect 479 1786 483 1790
rect 671 1786 675 1790
rect 727 1786 731 1790
rect 895 1786 899 1790
rect 959 1786 963 1790
rect 1119 1786 1123 1790
rect 1183 1786 1187 1790
rect 1343 1786 1347 1790
rect 1399 1786 1403 1790
rect 1567 1786 1571 1790
rect 1615 1786 1619 1790
rect 1799 1786 1803 1790
rect 1815 1786 1819 1790
rect 1935 1786 1939 1790
rect 3839 1786 3843 1790
rect 3887 1786 3891 1790
rect 4023 1786 4027 1790
rect 4191 1786 4195 1790
rect 4367 1786 4371 1790
rect 4559 1786 4563 1790
rect 4711 1786 4715 1790
rect 4767 1786 4771 1790
rect 4871 1786 4875 1790
rect 4983 1786 4987 1790
rect 5039 1786 5043 1790
rect 5207 1786 5211 1790
rect 5215 1786 5219 1790
rect 5383 1786 5387 1790
rect 5447 1786 5451 1790
rect 5543 1786 5547 1790
rect 5663 1786 5667 1790
rect 111 1674 115 1678
rect 203 1674 207 1678
rect 275 1674 279 1678
rect 419 1674 423 1678
rect 459 1674 463 1678
rect 643 1674 647 1678
rect 667 1674 671 1678
rect 867 1674 871 1678
rect 883 1674 887 1678
rect 1091 1674 1095 1678
rect 1115 1674 1119 1678
rect 1315 1674 1319 1678
rect 1355 1674 1359 1678
rect 1539 1674 1543 1678
rect 1595 1674 1599 1678
rect 1771 1674 1775 1678
rect 1935 1674 1939 1678
rect 3839 1674 3843 1678
rect 3859 1674 3863 1678
rect 3995 1674 3999 1678
rect 4131 1674 4135 1678
rect 4163 1674 4167 1678
rect 4283 1674 4287 1678
rect 4339 1674 4343 1678
rect 4483 1674 4487 1678
rect 4531 1674 4535 1678
rect 4715 1674 4719 1678
rect 4739 1674 4743 1678
rect 4955 1674 4959 1678
rect 4979 1674 4983 1678
rect 5187 1674 5191 1678
rect 5259 1674 5263 1678
rect 5419 1674 5423 1678
rect 5515 1674 5519 1678
rect 5663 1674 5667 1678
rect 1975 1666 1979 1670
rect 2231 1666 2235 1670
rect 2471 1666 2475 1670
rect 2599 1666 2603 1670
rect 2615 1666 2619 1670
rect 2767 1666 2771 1670
rect 2919 1666 2923 1670
rect 2967 1666 2971 1670
rect 3071 1666 3075 1670
rect 3223 1666 3227 1670
rect 3335 1666 3339 1670
rect 3679 1666 3683 1670
rect 3799 1666 3803 1670
rect 111 1562 115 1566
rect 303 1562 307 1566
rect 383 1562 387 1566
rect 487 1562 491 1566
rect 575 1562 579 1566
rect 695 1562 699 1566
rect 767 1562 771 1566
rect 911 1562 915 1566
rect 951 1562 955 1566
rect 1127 1562 1131 1566
rect 1143 1562 1147 1566
rect 1303 1562 1307 1566
rect 1383 1562 1387 1566
rect 1479 1562 1483 1566
rect 1623 1562 1627 1566
rect 1663 1562 1667 1566
rect 1935 1562 1939 1566
rect 3839 1562 3843 1566
rect 3887 1562 3891 1566
rect 4023 1562 4027 1566
rect 4047 1562 4051 1566
rect 4159 1562 4163 1566
rect 4271 1562 4275 1566
rect 4311 1562 4315 1566
rect 4511 1562 4515 1566
rect 4543 1562 4547 1566
rect 4743 1562 4747 1566
rect 4855 1562 4859 1566
rect 5007 1562 5011 1566
rect 5191 1562 5195 1566
rect 5287 1562 5291 1566
rect 5527 1562 5531 1566
rect 5543 1562 5547 1566
rect 5663 1562 5667 1566
rect 1975 1542 1979 1546
rect 1995 1542 1999 1546
rect 2203 1542 2207 1546
rect 2275 1542 2279 1546
rect 2539 1542 2543 1546
rect 2571 1542 2575 1546
rect 2779 1542 2783 1546
rect 2939 1542 2943 1546
rect 3011 1542 3015 1546
rect 3235 1542 3239 1546
rect 3307 1542 3311 1546
rect 3451 1542 3455 1546
rect 3651 1542 3655 1546
rect 3799 1542 3803 1546
rect 111 1430 115 1434
rect 331 1430 335 1434
rect 355 1430 359 1434
rect 547 1430 551 1434
rect 587 1430 591 1434
rect 739 1430 743 1434
rect 843 1430 847 1434
rect 923 1430 927 1434
rect 1099 1430 1103 1434
rect 1275 1430 1279 1434
rect 1363 1430 1367 1434
rect 1451 1430 1455 1434
rect 1635 1430 1639 1434
rect 1935 1430 1939 1434
rect 1975 1430 1979 1434
rect 2023 1430 2027 1434
rect 2191 1430 2195 1434
rect 2303 1430 2307 1434
rect 2399 1430 2403 1434
rect 2567 1430 2571 1434
rect 2615 1430 2619 1434
rect 2807 1430 2811 1434
rect 2831 1430 2835 1434
rect 3039 1430 3043 1434
rect 3055 1430 3059 1434
rect 3263 1430 3267 1434
rect 3287 1430 3291 1434
rect 3479 1430 3483 1434
rect 3527 1430 3531 1434
rect 3679 1430 3683 1434
rect 3799 1430 3803 1434
rect 3839 1434 3843 1438
rect 3859 1434 3863 1438
rect 3995 1434 3999 1438
rect 4019 1434 4023 1438
rect 4147 1434 4151 1438
rect 4243 1434 4247 1438
rect 4355 1434 4359 1438
rect 4515 1434 4519 1438
rect 4595 1434 4599 1438
rect 4827 1434 4831 1438
rect 4867 1434 4871 1438
rect 5163 1434 5167 1438
rect 5459 1434 5463 1438
rect 5499 1434 5503 1438
rect 5663 1434 5667 1438
rect 111 1318 115 1322
rect 359 1318 363 1322
rect 367 1318 371 1322
rect 551 1318 555 1322
rect 615 1318 619 1322
rect 727 1318 731 1322
rect 871 1318 875 1322
rect 895 1318 899 1322
rect 1063 1318 1067 1322
rect 1127 1318 1131 1322
rect 1223 1318 1227 1322
rect 1375 1318 1379 1322
rect 1391 1318 1395 1322
rect 1527 1318 1531 1322
rect 1679 1318 1683 1322
rect 1815 1318 1819 1322
rect 1935 1318 1939 1322
rect 3839 1318 3843 1322
rect 3887 1318 3891 1322
rect 4023 1318 4027 1322
rect 4047 1318 4051 1322
rect 4175 1318 4179 1322
rect 4239 1318 4243 1322
rect 4383 1318 4387 1322
rect 4455 1318 4459 1322
rect 4623 1318 4627 1322
rect 4695 1318 4699 1322
rect 4895 1318 4899 1322
rect 4951 1318 4955 1322
rect 5191 1318 5195 1322
rect 5223 1318 5227 1322
rect 5487 1318 5491 1322
rect 5495 1318 5499 1322
rect 5663 1318 5667 1322
rect 1975 1298 1979 1302
rect 1995 1298 1999 1302
rect 2163 1298 2167 1302
rect 2371 1298 2375 1302
rect 2587 1298 2591 1302
rect 2803 1298 2807 1302
rect 3027 1298 3031 1302
rect 3091 1298 3095 1302
rect 3227 1298 3231 1302
rect 3259 1298 3263 1302
rect 3363 1298 3367 1302
rect 3499 1298 3503 1302
rect 3799 1298 3803 1302
rect 111 1194 115 1198
rect 235 1194 239 1198
rect 339 1194 343 1198
rect 379 1194 383 1198
rect 523 1194 527 1198
rect 667 1194 671 1198
rect 699 1194 703 1198
rect 811 1194 815 1198
rect 867 1194 871 1198
rect 947 1194 951 1198
rect 1035 1194 1039 1198
rect 1091 1194 1095 1198
rect 1195 1194 1199 1198
rect 1235 1194 1239 1198
rect 1347 1194 1351 1198
rect 1379 1194 1383 1198
rect 1499 1194 1503 1198
rect 1515 1194 1519 1198
rect 1651 1194 1655 1198
rect 1787 1194 1791 1198
rect 1935 1194 1939 1198
rect 3839 1198 3843 1202
rect 3859 1198 3863 1202
rect 4019 1198 4023 1202
rect 4091 1198 4095 1202
rect 4211 1198 4215 1202
rect 4339 1198 4343 1202
rect 4427 1198 4431 1202
rect 4579 1198 4583 1202
rect 4667 1198 4671 1202
rect 4811 1198 4815 1202
rect 4923 1198 4927 1202
rect 5043 1198 5047 1202
rect 5195 1198 5199 1202
rect 5275 1198 5279 1202
rect 5467 1198 5471 1202
rect 5515 1198 5519 1202
rect 5663 1198 5667 1202
rect 1975 1186 1979 1190
rect 2983 1186 2987 1190
rect 3119 1186 3123 1190
rect 3255 1186 3259 1190
rect 3391 1186 3395 1190
rect 3799 1186 3803 1190
rect 111 1070 115 1074
rect 263 1070 267 1074
rect 407 1070 411 1074
rect 463 1070 467 1074
rect 551 1070 555 1074
rect 663 1070 667 1074
rect 695 1070 699 1074
rect 839 1070 843 1074
rect 871 1070 875 1074
rect 975 1070 979 1074
rect 1079 1070 1083 1074
rect 1119 1070 1123 1074
rect 1263 1070 1267 1074
rect 1407 1070 1411 1074
rect 1543 1070 1547 1074
rect 1679 1070 1683 1074
rect 1815 1070 1819 1074
rect 1935 1070 1939 1074
rect 1975 1074 1979 1078
rect 1995 1074 1999 1078
rect 2131 1074 2135 1078
rect 2275 1074 2279 1078
rect 2443 1074 2447 1078
rect 2627 1074 2631 1078
rect 2819 1074 2823 1078
rect 2955 1074 2959 1078
rect 3027 1074 3031 1078
rect 3091 1074 3095 1078
rect 3227 1074 3231 1078
rect 3235 1074 3239 1078
rect 3451 1074 3455 1078
rect 3651 1074 3655 1078
rect 3799 1074 3803 1078
rect 3839 1066 3843 1070
rect 3887 1066 3891 1070
rect 4119 1066 4123 1070
rect 4367 1066 4371 1070
rect 4607 1066 4611 1070
rect 4839 1066 4843 1070
rect 4863 1066 4867 1070
rect 4999 1066 5003 1070
rect 5071 1066 5075 1070
rect 5135 1066 5139 1070
rect 5271 1066 5275 1070
rect 5303 1066 5307 1070
rect 5407 1066 5411 1070
rect 5543 1066 5547 1070
rect 5663 1066 5667 1070
rect 1975 962 1979 966
rect 2023 962 2027 966
rect 2095 962 2099 966
rect 2159 962 2163 966
rect 2231 962 2235 966
rect 2303 962 2307 966
rect 2367 962 2371 966
rect 2471 962 2475 966
rect 2503 962 2507 966
rect 2655 962 2659 966
rect 2831 962 2835 966
rect 2847 962 2851 966
rect 3023 962 3027 966
rect 3055 962 3059 966
rect 3231 962 3235 966
rect 3263 962 3267 966
rect 3455 962 3459 966
rect 3479 962 3483 966
rect 3679 962 3683 966
rect 3799 962 3803 966
rect 111 946 115 950
rect 195 946 199 950
rect 235 946 239 950
rect 371 946 375 950
rect 435 946 439 950
rect 547 946 551 950
rect 635 946 639 950
rect 723 946 727 950
rect 843 946 847 950
rect 907 946 911 950
rect 1051 946 1055 950
rect 1091 946 1095 950
rect 1935 946 1939 950
rect 3839 942 3843 946
rect 4587 942 4591 946
rect 4755 942 4759 946
rect 4835 942 4839 946
rect 4939 942 4943 946
rect 4971 942 4975 946
rect 5107 942 5111 946
rect 5131 942 5135 946
rect 5243 942 5247 946
rect 5331 942 5335 946
rect 5379 942 5383 946
rect 5515 942 5519 946
rect 5663 942 5667 946
rect 1975 850 1979 854
rect 2067 850 2071 854
rect 2203 850 2207 854
rect 2307 850 2311 854
rect 2339 850 2343 854
rect 2475 850 2479 854
rect 2483 850 2487 854
rect 2627 850 2631 854
rect 2659 850 2663 854
rect 2803 850 2807 854
rect 2827 850 2831 854
rect 2995 850 2999 854
rect 3163 850 3167 854
rect 3203 850 3207 854
rect 3331 850 3335 854
rect 3427 850 3431 854
rect 3499 850 3503 854
rect 3651 850 3655 854
rect 3799 850 3803 854
rect 111 818 115 822
rect 159 818 163 822
rect 223 818 227 822
rect 351 818 355 822
rect 399 818 403 822
rect 575 818 579 822
rect 583 818 587 822
rect 751 818 755 822
rect 839 818 843 822
rect 935 818 939 822
rect 1111 818 1115 822
rect 1119 818 1123 822
rect 1399 818 1403 822
rect 1687 818 1691 822
rect 1935 818 1939 822
rect 3839 822 3843 826
rect 3983 822 3987 826
rect 4239 822 4243 826
rect 4535 822 4539 826
rect 4615 822 4619 826
rect 4783 822 4787 826
rect 4863 822 4867 826
rect 4967 822 4971 826
rect 5159 822 5163 826
rect 5215 822 5219 826
rect 5359 822 5363 826
rect 5543 822 5547 826
rect 5663 822 5667 826
rect 1975 734 1979 738
rect 2335 734 2339 738
rect 2511 734 2515 738
rect 2687 734 2691 738
rect 2855 734 2859 738
rect 3023 734 3027 738
rect 3135 734 3139 738
rect 3191 734 3195 738
rect 3271 734 3275 738
rect 3359 734 3363 738
rect 3407 734 3411 738
rect 3527 734 3531 738
rect 3543 734 3547 738
rect 3679 734 3683 738
rect 3799 734 3803 738
rect 111 706 115 710
rect 131 706 135 710
rect 291 706 295 710
rect 323 706 327 710
rect 483 706 487 710
rect 555 706 559 710
rect 675 706 679 710
rect 811 706 815 710
rect 867 706 871 710
rect 1059 706 1063 710
rect 1083 706 1087 710
rect 1251 706 1255 710
rect 1371 706 1375 710
rect 1435 706 1439 710
rect 1619 706 1623 710
rect 1659 706 1663 710
rect 1787 706 1791 710
rect 1935 706 1939 710
rect 111 594 115 598
rect 159 594 163 598
rect 319 594 323 598
rect 327 594 331 598
rect 511 594 515 598
rect 519 594 523 598
rect 703 594 707 598
rect 711 594 715 598
rect 895 594 899 598
rect 903 594 907 598
rect 1087 594 1091 598
rect 1095 594 1099 598
rect 1279 594 1283 598
rect 1463 594 1467 598
rect 1647 594 1651 598
rect 1815 594 1819 598
rect 1935 594 1939 598
rect 111 482 115 486
rect 131 482 135 486
rect 299 482 303 486
rect 395 482 399 486
rect 491 482 495 486
rect 587 482 591 486
rect 683 482 687 486
rect 787 482 791 486
rect 875 482 879 486
rect 987 482 991 486
rect 1067 482 1071 486
rect 1195 482 1199 486
rect 1251 482 1255 486
rect 1411 482 1415 486
rect 1435 482 1439 486
rect 1619 482 1623 486
rect 1787 482 1791 486
rect 1935 482 1939 486
rect 3839 686 3843 690
rect 3859 686 3863 690
rect 3955 686 3959 690
rect 3995 686 3999 690
rect 4139 686 4143 690
rect 4211 686 4215 690
rect 4323 686 4327 690
rect 4507 686 4511 690
rect 4531 686 4535 690
rect 4755 686 4759 690
rect 4835 686 4839 690
rect 4995 686 4999 690
rect 5187 686 5191 690
rect 5243 686 5247 690
rect 5499 686 5503 690
rect 5515 686 5519 690
rect 5663 686 5667 690
rect 3839 574 3843 578
rect 3887 574 3891 578
rect 4023 574 4027 578
rect 4159 574 4163 578
rect 4167 574 4171 578
rect 4295 574 4299 578
rect 4351 574 4355 578
rect 4431 574 4435 578
rect 4559 574 4563 578
rect 4575 574 4579 578
rect 4743 574 4747 578
rect 4783 574 4787 578
rect 4927 574 4931 578
rect 5023 574 5027 578
rect 5119 574 5123 578
rect 5271 574 5275 578
rect 5319 574 5323 578
rect 5527 574 5531 578
rect 5663 574 5667 578
rect 1975 462 1979 466
rect 1995 462 1999 466
rect 2203 462 2207 466
rect 2427 462 2431 466
rect 2651 462 2655 466
rect 2867 462 2871 466
rect 3075 462 3079 466
rect 3107 462 3111 466
rect 3243 462 3247 466
rect 3275 462 3279 466
rect 3379 462 3383 466
rect 3475 462 3479 466
rect 3515 462 3519 466
rect 3651 462 3655 466
rect 3799 462 3803 466
rect 3839 462 3843 466
rect 3859 462 3863 466
rect 3995 462 3999 466
rect 4131 462 4135 466
rect 4267 462 4271 466
rect 4379 462 4383 466
rect 4403 462 4407 466
rect 4547 462 4551 466
rect 4595 462 4599 466
rect 4715 462 4719 466
rect 4819 462 4823 466
rect 4899 462 4903 466
rect 5051 462 5055 466
rect 5091 462 5095 466
rect 5283 462 5287 466
rect 5291 462 5295 466
rect 5499 462 5503 466
rect 5663 462 5667 466
rect 111 358 115 362
rect 423 358 427 362
rect 615 358 619 362
rect 647 358 651 362
rect 815 358 819 362
rect 991 358 995 362
rect 1015 358 1019 362
rect 1167 358 1171 362
rect 1223 358 1227 362
rect 1343 358 1347 362
rect 1439 358 1443 362
rect 1935 358 1939 362
rect 3839 350 3843 354
rect 4407 350 4411 354
rect 4623 350 4627 354
rect 4639 350 4643 354
rect 4807 350 4811 354
rect 4847 350 4851 354
rect 4983 350 4987 354
rect 5079 350 5083 354
rect 5167 350 5171 354
rect 5311 350 5315 354
rect 5359 350 5363 354
rect 5543 350 5547 354
rect 5663 350 5667 354
rect 1975 334 1979 338
rect 2023 334 2027 338
rect 2159 334 2163 338
rect 2231 334 2235 338
rect 2295 334 2299 338
rect 2431 334 2435 338
rect 2455 334 2459 338
rect 2567 334 2571 338
rect 2679 334 2683 338
rect 2703 334 2707 338
rect 2839 334 2843 338
rect 2895 334 2899 338
rect 2975 334 2979 338
rect 3103 334 3107 338
rect 3111 334 3115 338
rect 3247 334 3251 338
rect 3303 334 3307 338
rect 3383 334 3387 338
rect 3503 334 3507 338
rect 3519 334 3523 338
rect 3655 334 3659 338
rect 3679 334 3683 338
rect 3799 334 3803 338
rect 111 206 115 210
rect 539 206 543 210
rect 619 206 623 210
rect 675 206 679 210
rect 787 206 791 210
rect 811 206 815 210
rect 947 206 951 210
rect 963 206 967 210
rect 1083 206 1087 210
rect 1139 206 1143 210
rect 1219 206 1223 210
rect 1315 206 1319 210
rect 1355 206 1359 210
rect 1491 206 1495 210
rect 1935 206 1939 210
rect 3839 210 3843 214
rect 4291 210 4295 214
rect 4427 210 4431 214
rect 4563 210 4567 214
rect 4611 210 4615 214
rect 4699 210 4703 214
rect 4779 210 4783 214
rect 4835 210 4839 214
rect 4955 210 4959 214
rect 4971 210 4975 214
rect 5107 210 5111 214
rect 5139 210 5143 214
rect 5243 210 5247 214
rect 5331 210 5335 214
rect 5379 210 5383 214
rect 5515 210 5519 214
rect 5663 210 5667 214
rect 1975 186 1979 190
rect 1995 186 1999 190
rect 2131 186 2135 190
rect 2267 186 2271 190
rect 2403 186 2407 190
rect 2539 186 2543 190
rect 2675 186 2679 190
rect 2811 186 2815 190
rect 2947 186 2951 190
rect 3083 186 3087 190
rect 3219 186 3223 190
rect 3355 186 3359 190
rect 3491 186 3495 190
rect 3627 186 3631 190
rect 3799 186 3803 190
rect 111 94 115 98
rect 567 94 571 98
rect 703 94 707 98
rect 839 94 843 98
rect 975 94 979 98
rect 1111 94 1115 98
rect 1247 94 1251 98
rect 1383 94 1387 98
rect 1519 94 1523 98
rect 1935 94 1939 98
rect 3839 98 3843 102
rect 4319 98 4323 102
rect 4455 98 4459 102
rect 4591 98 4595 102
rect 4727 98 4731 102
rect 4863 98 4867 102
rect 4999 98 5003 102
rect 5135 98 5139 102
rect 5271 98 5275 102
rect 5407 98 5411 102
rect 5543 98 5547 102
rect 5663 98 5667 102
rect 1975 74 1979 78
rect 2023 74 2027 78
rect 2159 74 2163 78
rect 2295 74 2299 78
rect 2431 74 2435 78
rect 2567 74 2571 78
rect 2703 74 2707 78
rect 2839 74 2843 78
rect 2975 74 2979 78
rect 3111 74 3115 78
rect 3247 74 3251 78
rect 3383 74 3387 78
rect 3519 74 3523 78
rect 3655 74 3659 78
rect 3799 74 3803 78
<< m4 >>
rect 84 5717 85 5723
rect 91 5722 1947 5723
rect 91 5718 111 5722
rect 115 5718 159 5722
rect 163 5718 303 5722
rect 307 5718 503 5722
rect 507 5718 727 5722
rect 731 5718 983 5722
rect 987 5718 1255 5722
rect 1259 5718 1543 5722
rect 1547 5718 1815 5722
rect 1819 5718 1935 5722
rect 1939 5718 1947 5722
rect 91 5717 1947 5718
rect 1953 5717 1954 5723
rect 1958 5689 1959 5695
rect 1965 5694 3823 5695
rect 1965 5690 1975 5694
rect 1979 5690 1995 5694
rect 1999 5690 2179 5694
rect 2183 5690 2387 5694
rect 2391 5690 2587 5694
rect 2591 5690 2779 5694
rect 2783 5690 2963 5694
rect 2967 5690 3147 5694
rect 3151 5690 3323 5694
rect 3327 5690 3499 5694
rect 3503 5690 3651 5694
rect 3655 5690 3799 5694
rect 3803 5690 3823 5694
rect 1965 5689 3823 5690
rect 3829 5689 3830 5695
rect 3822 5645 3823 5651
rect 3829 5650 5707 5651
rect 3829 5646 3839 5650
rect 3843 5646 4291 5650
rect 4295 5646 4427 5650
rect 4431 5646 4563 5650
rect 4567 5646 4699 5650
rect 4703 5646 4835 5650
rect 4839 5646 4971 5650
rect 4975 5646 5107 5650
rect 5111 5646 5663 5650
rect 5667 5646 5707 5650
rect 3829 5645 5707 5646
rect 5713 5645 5714 5651
rect 96 5601 97 5607
rect 103 5606 1959 5607
rect 103 5602 111 5606
rect 115 5602 131 5606
rect 135 5602 275 5606
rect 279 5602 475 5606
rect 479 5602 563 5606
rect 567 5602 699 5606
rect 703 5602 723 5606
rect 727 5602 883 5606
rect 887 5602 955 5606
rect 959 5602 1051 5606
rect 1055 5602 1227 5606
rect 1231 5602 1403 5606
rect 1407 5602 1515 5606
rect 1519 5602 1579 5606
rect 1583 5602 1763 5606
rect 1767 5602 1787 5606
rect 1791 5602 1935 5606
rect 1939 5602 1959 5606
rect 103 5601 1959 5602
rect 1965 5601 1966 5607
rect 1946 5577 1947 5583
rect 1953 5582 3811 5583
rect 1953 5578 1975 5582
rect 1979 5578 2023 5582
rect 2027 5578 2207 5582
rect 2211 5578 2263 5582
rect 2267 5578 2415 5582
rect 2419 5578 2503 5582
rect 2507 5578 2615 5582
rect 2619 5578 2743 5582
rect 2747 5578 2807 5582
rect 2811 5578 2983 5582
rect 2987 5578 2991 5582
rect 2995 5578 3175 5582
rect 3179 5578 3223 5582
rect 3227 5578 3351 5582
rect 3355 5578 3463 5582
rect 3467 5578 3527 5582
rect 3531 5578 3679 5582
rect 3683 5578 3799 5582
rect 3803 5578 3811 5582
rect 1953 5577 3811 5578
rect 3817 5577 3818 5583
rect 3810 5533 3811 5539
rect 3817 5538 5695 5539
rect 3817 5534 3839 5538
rect 3843 5534 3887 5538
rect 3891 5534 4127 5538
rect 4131 5534 4319 5538
rect 4323 5534 4375 5538
rect 4379 5534 4455 5538
rect 4459 5534 4591 5538
rect 4595 5534 4615 5538
rect 4619 5534 4727 5538
rect 4731 5534 4847 5538
rect 4851 5534 4863 5538
rect 4867 5534 4999 5538
rect 5003 5534 5079 5538
rect 5083 5534 5135 5538
rect 5139 5534 5311 5538
rect 5315 5534 5663 5538
rect 5667 5534 5695 5538
rect 3817 5533 5695 5534
rect 5701 5533 5702 5539
rect 84 5477 85 5483
rect 91 5482 1947 5483
rect 91 5478 111 5482
rect 115 5478 591 5482
rect 595 5478 727 5482
rect 731 5478 751 5482
rect 755 5478 863 5482
rect 867 5478 911 5482
rect 915 5478 999 5482
rect 1003 5478 1079 5482
rect 1083 5478 1135 5482
rect 1139 5478 1255 5482
rect 1259 5478 1271 5482
rect 1275 5478 1407 5482
rect 1411 5478 1431 5482
rect 1435 5478 1543 5482
rect 1547 5478 1607 5482
rect 1611 5478 1679 5482
rect 1683 5478 1791 5482
rect 1795 5478 1815 5482
rect 1819 5478 1935 5482
rect 1939 5478 1947 5482
rect 91 5477 1947 5478
rect 1953 5477 1954 5483
rect 1958 5457 1959 5463
rect 1965 5462 3823 5463
rect 1965 5458 1975 5462
rect 1979 5458 2235 5462
rect 2239 5458 2427 5462
rect 2431 5458 2475 5462
rect 2479 5458 2643 5462
rect 2647 5458 2715 5462
rect 2719 5458 2859 5462
rect 2863 5458 2955 5462
rect 2959 5458 3075 5462
rect 3079 5458 3195 5462
rect 3199 5458 3291 5462
rect 3295 5458 3435 5462
rect 3439 5458 3651 5462
rect 3655 5458 3799 5462
rect 3803 5458 3823 5462
rect 1965 5457 3823 5458
rect 3829 5457 3830 5463
rect 3822 5417 3823 5423
rect 3829 5422 5707 5423
rect 3829 5418 3839 5422
rect 3843 5418 3859 5422
rect 3863 5418 4075 5422
rect 4079 5418 4099 5422
rect 4103 5418 4307 5422
rect 4311 5418 4347 5422
rect 4351 5418 4531 5422
rect 4535 5418 4587 5422
rect 4591 5418 4739 5422
rect 4743 5418 4819 5422
rect 4823 5418 4939 5422
rect 4943 5418 5051 5422
rect 5055 5418 5139 5422
rect 5143 5418 5283 5422
rect 5287 5418 5339 5422
rect 5343 5418 5515 5422
rect 5519 5418 5663 5422
rect 5667 5418 5707 5422
rect 3829 5417 5707 5418
rect 5713 5417 5714 5423
rect 1946 5345 1947 5351
rect 1953 5350 3811 5351
rect 1953 5346 1975 5350
rect 1979 5346 2447 5350
rect 2451 5346 2455 5350
rect 2459 5346 2583 5350
rect 2587 5346 2671 5350
rect 2675 5346 2719 5350
rect 2723 5346 2855 5350
rect 2859 5346 2887 5350
rect 2891 5346 2991 5350
rect 2995 5346 3103 5350
rect 3107 5346 3135 5350
rect 3139 5346 3287 5350
rect 3291 5346 3319 5350
rect 3323 5346 3799 5350
rect 3803 5346 3811 5350
rect 1953 5345 3811 5346
rect 3817 5345 3818 5351
rect 3810 5289 3811 5295
rect 3817 5294 5695 5295
rect 3817 5290 3839 5294
rect 3843 5290 3887 5294
rect 3891 5290 4095 5294
rect 4099 5290 4103 5294
rect 4107 5290 4335 5294
rect 4339 5290 4343 5294
rect 4347 5290 4559 5294
rect 4563 5290 4615 5294
rect 4619 5290 4767 5294
rect 4771 5290 4911 5294
rect 4915 5290 4967 5294
rect 4971 5290 5167 5294
rect 5171 5290 5215 5294
rect 5219 5290 5367 5294
rect 5371 5290 5527 5294
rect 5531 5290 5543 5294
rect 5547 5290 5663 5294
rect 5667 5290 5695 5294
rect 3817 5289 5695 5290
rect 5701 5289 5702 5295
rect 96 5261 97 5267
rect 103 5266 1959 5267
rect 103 5262 111 5266
rect 115 5262 459 5266
rect 463 5262 563 5266
rect 567 5262 595 5266
rect 599 5262 699 5266
rect 703 5262 731 5266
rect 735 5262 835 5266
rect 839 5262 867 5266
rect 871 5262 971 5266
rect 975 5262 1003 5266
rect 1007 5262 1107 5266
rect 1111 5262 1139 5266
rect 1143 5262 1243 5266
rect 1247 5262 1275 5266
rect 1279 5262 1379 5266
rect 1383 5262 1411 5266
rect 1415 5262 1515 5266
rect 1519 5262 1547 5266
rect 1551 5262 1651 5266
rect 1655 5262 1787 5266
rect 1791 5262 1935 5266
rect 1939 5262 1959 5266
rect 103 5261 1959 5262
rect 1965 5261 1966 5267
rect 1958 5233 1959 5239
rect 1965 5238 3823 5239
rect 1965 5234 1975 5238
rect 1979 5234 2099 5238
rect 2103 5234 2235 5238
rect 2239 5234 2379 5238
rect 2383 5234 2419 5238
rect 2423 5234 2531 5238
rect 2535 5234 2555 5238
rect 2559 5234 2691 5238
rect 2695 5234 2699 5238
rect 2703 5234 2827 5238
rect 2831 5234 2883 5238
rect 2887 5234 2963 5238
rect 2967 5234 3067 5238
rect 3071 5234 3107 5238
rect 3111 5234 3259 5238
rect 3263 5234 3799 5238
rect 3803 5234 3823 5238
rect 1965 5233 3823 5234
rect 3829 5233 3830 5239
rect 3822 5169 3823 5175
rect 3829 5174 5707 5175
rect 3829 5170 3839 5174
rect 3843 5170 3859 5174
rect 3863 5170 3995 5174
rect 3999 5170 4067 5174
rect 4071 5170 4155 5174
rect 4159 5170 4315 5174
rect 4319 5170 4363 5174
rect 4367 5170 4587 5174
rect 4591 5170 4611 5174
rect 4615 5170 4883 5174
rect 4887 5170 5171 5174
rect 5175 5170 5187 5174
rect 5191 5170 5467 5174
rect 5471 5170 5499 5174
rect 5503 5170 5663 5174
rect 5667 5170 5707 5174
rect 3829 5169 5707 5170
rect 5713 5169 5714 5175
rect 84 5133 85 5139
rect 91 5138 1947 5139
rect 91 5134 111 5138
rect 115 5134 319 5138
rect 323 5134 487 5138
rect 491 5134 503 5138
rect 507 5134 623 5138
rect 627 5134 703 5138
rect 707 5134 759 5138
rect 763 5134 895 5138
rect 899 5134 919 5138
rect 923 5134 1031 5138
rect 1035 5134 1151 5138
rect 1155 5134 1167 5138
rect 1171 5134 1303 5138
rect 1307 5134 1391 5138
rect 1395 5134 1439 5138
rect 1443 5134 1575 5138
rect 1579 5134 1631 5138
rect 1635 5134 1935 5138
rect 1939 5134 1947 5138
rect 91 5133 1947 5134
rect 1953 5133 1954 5139
rect 1946 5097 1947 5103
rect 1953 5102 3811 5103
rect 1953 5098 1975 5102
rect 1979 5098 2079 5102
rect 2083 5098 2127 5102
rect 2131 5098 2263 5102
rect 2267 5098 2359 5102
rect 2363 5098 2407 5102
rect 2411 5098 2559 5102
rect 2563 5098 2639 5102
rect 2643 5098 2727 5102
rect 2731 5098 2911 5102
rect 2915 5098 3095 5102
rect 3099 5098 3175 5102
rect 3179 5098 3287 5102
rect 3291 5098 3439 5102
rect 3443 5098 3679 5102
rect 3683 5098 3799 5102
rect 3803 5098 3811 5102
rect 1953 5097 3811 5098
rect 3817 5097 3818 5103
rect 3810 5041 3811 5047
rect 3817 5046 5695 5047
rect 3817 5042 3839 5046
rect 3843 5042 3887 5046
rect 3891 5042 4023 5046
rect 4027 5042 4183 5046
rect 4187 5042 4391 5046
rect 4395 5042 4447 5046
rect 4451 5042 4631 5046
rect 4635 5042 4639 5046
rect 4643 5042 4831 5046
rect 4835 5042 4911 5046
rect 4915 5042 5047 5046
rect 5051 5042 5199 5046
rect 5203 5042 5279 5046
rect 5283 5042 5495 5046
rect 5499 5042 5511 5046
rect 5515 5042 5663 5046
rect 5667 5042 5695 5046
rect 3817 5041 5695 5042
rect 5701 5041 5702 5047
rect 96 5021 97 5027
rect 103 5026 1959 5027
rect 103 5022 111 5026
rect 115 5022 139 5026
rect 143 5022 291 5026
rect 295 5022 411 5026
rect 415 5022 475 5026
rect 479 5022 675 5026
rect 679 5022 683 5026
rect 687 5022 891 5026
rect 895 5022 963 5026
rect 967 5022 1123 5026
rect 1127 5022 1243 5026
rect 1247 5022 1363 5026
rect 1367 5022 1523 5026
rect 1527 5022 1603 5026
rect 1607 5022 1787 5026
rect 1791 5022 1935 5026
rect 1939 5022 1959 5026
rect 103 5021 1959 5022
rect 1965 5021 1966 5027
rect 1958 4965 1959 4971
rect 1965 4970 3823 4971
rect 1965 4966 1975 4970
rect 1979 4966 1995 4970
rect 1999 4966 2051 4970
rect 2055 4966 2131 4970
rect 2135 4966 2299 4970
rect 2303 4966 2331 4970
rect 2335 4966 2467 4970
rect 2471 4966 2611 4970
rect 2615 4966 2643 4970
rect 2647 4966 2819 4970
rect 2823 4966 2883 4970
rect 2887 4966 2987 4970
rect 2991 4966 3147 4970
rect 3151 4966 3155 4970
rect 3159 4966 3323 4970
rect 3327 4966 3411 4970
rect 3415 4966 3499 4970
rect 3503 4966 3651 4970
rect 3655 4966 3799 4970
rect 3803 4966 3823 4970
rect 1965 4965 3823 4966
rect 3829 4965 3830 4971
rect 84 4909 85 4915
rect 91 4914 1947 4915
rect 91 4910 111 4914
rect 115 4910 159 4914
rect 163 4910 167 4914
rect 171 4910 415 4914
rect 419 4910 439 4914
rect 443 4910 711 4914
rect 715 4910 735 4914
rect 739 4910 991 4914
rect 995 4910 1087 4914
rect 1091 4910 1271 4914
rect 1275 4910 1463 4914
rect 1467 4910 1551 4914
rect 1555 4910 1815 4914
rect 1819 4910 1935 4914
rect 1939 4910 1947 4914
rect 91 4909 1947 4910
rect 1953 4909 1954 4915
rect 3822 4913 3823 4919
rect 3829 4918 5707 4919
rect 3829 4914 3839 4918
rect 3843 4914 4419 4918
rect 4423 4914 4603 4918
rect 4607 4914 4675 4918
rect 4679 4914 4803 4918
rect 4807 4914 4827 4918
rect 4831 4914 4987 4918
rect 4991 4914 5019 4918
rect 5023 4914 5155 4918
rect 5159 4914 5251 4918
rect 5255 4914 5323 4918
rect 5327 4914 5483 4918
rect 5487 4914 5499 4918
rect 5503 4914 5663 4918
rect 5667 4914 5707 4918
rect 3829 4913 5707 4914
rect 5713 4913 5714 4919
rect 1946 4825 1947 4831
rect 1953 4830 3811 4831
rect 1953 4826 1975 4830
rect 1979 4826 2023 4830
rect 2027 4826 2159 4830
rect 2163 4826 2327 4830
rect 2331 4826 2391 4830
rect 2395 4826 2495 4830
rect 2499 4826 2527 4830
rect 2531 4826 2663 4830
rect 2667 4826 2671 4830
rect 2675 4826 2807 4830
rect 2811 4826 2847 4830
rect 2851 4826 2951 4830
rect 2955 4826 3015 4830
rect 3019 4826 3095 4830
rect 3099 4826 3183 4830
rect 3187 4826 3239 4830
rect 3243 4826 3351 4830
rect 3355 4826 3383 4830
rect 3387 4826 3527 4830
rect 3531 4826 3679 4830
rect 3683 4826 3799 4830
rect 3803 4826 3811 4830
rect 1953 4825 3811 4826
rect 3817 4825 3818 4831
rect 96 4785 97 4791
rect 103 4790 1959 4791
rect 103 4786 111 4790
rect 115 4786 131 4790
rect 135 4786 267 4790
rect 271 4786 387 4790
rect 391 4786 403 4790
rect 407 4786 539 4790
rect 543 4786 675 4790
rect 679 4786 707 4790
rect 711 4786 1059 4790
rect 1063 4786 1435 4790
rect 1439 4786 1787 4790
rect 1791 4786 1935 4790
rect 1939 4786 1959 4790
rect 103 4785 1959 4786
rect 1965 4785 1966 4791
rect 3810 4781 3811 4787
rect 3817 4786 5695 4787
rect 3817 4782 3839 4786
rect 3843 4782 4703 4786
rect 4707 4782 4855 4786
rect 4859 4782 4991 4786
rect 4995 4782 5015 4786
rect 5019 4782 5127 4786
rect 5131 4782 5183 4786
rect 5187 4782 5263 4786
rect 5267 4782 5351 4786
rect 5355 4782 5399 4786
rect 5403 4782 5527 4786
rect 5531 4782 5535 4786
rect 5539 4782 5663 4786
rect 5667 4782 5695 4786
rect 3817 4781 5695 4782
rect 5701 4781 5702 4787
rect 1958 4705 1959 4711
rect 1965 4710 3823 4711
rect 1965 4706 1975 4710
rect 1979 4706 1995 4710
rect 1999 4706 2131 4710
rect 2135 4706 2267 4710
rect 2271 4706 2363 4710
rect 2367 4706 2427 4710
rect 2431 4706 2499 4710
rect 2503 4706 2587 4710
rect 2591 4706 2635 4710
rect 2639 4706 2747 4710
rect 2751 4706 2779 4710
rect 2783 4706 2907 4710
rect 2911 4706 2923 4710
rect 2927 4706 3067 4710
rect 3071 4706 3211 4710
rect 3215 4706 3235 4710
rect 3239 4706 3355 4710
rect 3359 4706 3499 4710
rect 3503 4706 3799 4710
rect 3803 4706 3823 4710
rect 1965 4705 3823 4706
rect 3829 4705 3830 4711
rect 84 4669 85 4675
rect 91 4674 1947 4675
rect 91 4670 111 4674
rect 115 4670 159 4674
rect 163 4670 295 4674
rect 299 4670 431 4674
rect 435 4670 567 4674
rect 571 4670 703 4674
rect 707 4670 1935 4674
rect 1939 4670 1947 4674
rect 91 4669 1947 4670
rect 1953 4669 1954 4675
rect 3822 4649 3823 4655
rect 3829 4654 5707 4655
rect 3829 4650 3839 4654
rect 3843 4650 4715 4654
rect 4719 4650 4827 4654
rect 4831 4650 4859 4654
rect 4863 4650 4963 4654
rect 4967 4650 5011 4654
rect 5015 4650 5099 4654
rect 5103 4650 5171 4654
rect 5175 4650 5235 4654
rect 5239 4650 5339 4654
rect 5343 4650 5371 4654
rect 5375 4650 5507 4654
rect 5511 4650 5515 4654
rect 5519 4650 5663 4654
rect 5667 4650 5707 4654
rect 3829 4649 5707 4650
rect 5713 4649 5714 4655
rect 1946 4593 1947 4599
rect 1953 4598 3811 4599
rect 1953 4594 1975 4598
rect 1979 4594 2023 4598
rect 2027 4594 2159 4598
rect 2163 4594 2175 4598
rect 2179 4594 2295 4598
rect 2299 4594 2351 4598
rect 2355 4594 2455 4598
rect 2459 4594 2527 4598
rect 2531 4594 2615 4598
rect 2619 4594 2695 4598
rect 2699 4594 2775 4598
rect 2779 4594 2871 4598
rect 2875 4594 2935 4598
rect 2939 4594 3047 4598
rect 3051 4594 3095 4598
rect 3099 4594 3263 4598
rect 3267 4594 3799 4598
rect 3803 4594 3811 4598
rect 1953 4593 3811 4594
rect 3817 4593 3818 4599
rect 96 4545 97 4551
rect 103 4550 1959 4551
rect 103 4546 111 4550
rect 115 4546 131 4550
rect 135 4546 267 4550
rect 271 4546 299 4550
rect 303 4546 403 4550
rect 407 4546 491 4550
rect 495 4546 539 4550
rect 543 4546 675 4550
rect 679 4546 691 4550
rect 695 4546 907 4550
rect 911 4546 1123 4550
rect 1127 4546 1347 4550
rect 1351 4546 1579 4550
rect 1583 4546 1787 4550
rect 1791 4546 1935 4550
rect 1939 4546 1959 4550
rect 103 4545 1959 4546
rect 1965 4545 1966 4551
rect 3810 4513 3811 4519
rect 3817 4518 5695 4519
rect 3817 4514 3839 4518
rect 3843 4514 3887 4518
rect 3891 4514 4063 4518
rect 4067 4514 4279 4518
rect 4283 4514 4503 4518
rect 4507 4514 4743 4518
rect 4747 4514 4751 4518
rect 4755 4514 4887 4518
rect 4891 4514 5007 4518
rect 5011 4514 5039 4518
rect 5043 4514 5199 4518
rect 5203 4514 5271 4518
rect 5275 4514 5367 4518
rect 5371 4514 5543 4518
rect 5547 4514 5663 4518
rect 5667 4514 5695 4518
rect 3817 4513 5695 4514
rect 5701 4513 5702 4519
rect 1958 4441 1959 4447
rect 1965 4446 3823 4447
rect 1965 4442 1975 4446
rect 1979 4442 1995 4446
rect 1999 4442 2147 4446
rect 2151 4442 2323 4446
rect 2327 4442 2499 4446
rect 2503 4442 2571 4446
rect 2575 4442 2667 4446
rect 2671 4442 2843 4446
rect 2847 4442 3019 4446
rect 3023 4442 3123 4446
rect 3127 4442 3651 4446
rect 3655 4442 3799 4446
rect 3803 4442 3823 4446
rect 1965 4441 3823 4442
rect 3829 4441 3830 4447
rect 84 4433 85 4439
rect 91 4438 1947 4439
rect 91 4434 111 4438
rect 115 4434 327 4438
rect 331 4434 519 4438
rect 523 4434 559 4438
rect 563 4434 719 4438
rect 723 4434 887 4438
rect 891 4434 935 4438
rect 939 4434 1063 4438
rect 1067 4434 1151 4438
rect 1155 4434 1247 4438
rect 1251 4434 1375 4438
rect 1379 4434 1439 4438
rect 1443 4434 1607 4438
rect 1611 4434 1631 4438
rect 1635 4434 1815 4438
rect 1819 4434 1935 4438
rect 1939 4434 1947 4438
rect 91 4433 1947 4434
rect 1953 4433 1954 4439
rect 3822 4401 3823 4407
rect 3829 4406 5707 4407
rect 3829 4402 3839 4406
rect 3843 4402 3859 4406
rect 3863 4402 3995 4406
rect 3999 4402 4035 4406
rect 4039 4402 4131 4406
rect 4135 4402 4251 4406
rect 4255 4402 4267 4406
rect 4271 4402 4403 4406
rect 4407 4402 4475 4406
rect 4479 4402 4587 4406
rect 4591 4402 4723 4406
rect 4727 4402 4795 4406
rect 4799 4402 4979 4406
rect 4983 4402 5027 4406
rect 5031 4402 5243 4406
rect 5247 4402 5275 4406
rect 5279 4402 5515 4406
rect 5519 4402 5663 4406
rect 5667 4402 5707 4406
rect 3829 4401 5707 4402
rect 5713 4401 5714 4407
rect 1946 4325 1947 4331
rect 1953 4330 3811 4331
rect 1953 4326 1975 4330
rect 1979 4326 2399 4330
rect 2403 4326 2599 4330
rect 2603 4326 2791 4330
rect 2795 4326 2983 4330
rect 2987 4326 3151 4330
rect 3155 4326 3167 4330
rect 3171 4326 3343 4330
rect 3347 4326 3519 4330
rect 3523 4326 3679 4330
rect 3683 4326 3799 4330
rect 3803 4326 3811 4330
rect 1953 4325 3811 4326
rect 3817 4325 3818 4331
rect 96 4313 97 4319
rect 103 4318 1959 4319
rect 103 4314 111 4318
rect 115 4314 531 4318
rect 535 4314 691 4318
rect 695 4314 747 4318
rect 751 4314 859 4318
rect 863 4314 883 4318
rect 887 4314 1019 4318
rect 1023 4314 1035 4318
rect 1039 4314 1155 4318
rect 1159 4314 1219 4318
rect 1223 4314 1291 4318
rect 1295 4314 1411 4318
rect 1415 4314 1427 4318
rect 1431 4314 1563 4318
rect 1567 4314 1603 4318
rect 1607 4314 1699 4318
rect 1703 4314 1787 4318
rect 1791 4314 1935 4318
rect 1939 4314 1959 4318
rect 103 4313 1959 4314
rect 1965 4313 1966 4319
rect 3810 4289 3811 4295
rect 3817 4294 5695 4295
rect 3817 4290 3839 4294
rect 3843 4290 3887 4294
rect 3891 4290 4023 4294
rect 4027 4290 4047 4294
rect 4051 4290 4159 4294
rect 4163 4290 4223 4294
rect 4227 4290 4295 4294
rect 4299 4290 4431 4294
rect 4435 4290 4615 4294
rect 4619 4290 4679 4294
rect 4683 4290 4823 4294
rect 4827 4290 4959 4294
rect 4963 4290 5055 4294
rect 5059 4290 5255 4294
rect 5259 4290 5303 4294
rect 5307 4290 5543 4294
rect 5547 4290 5663 4294
rect 5667 4290 5695 4294
rect 3817 4289 5695 4290
rect 5701 4289 5702 4295
rect 1958 4201 1959 4207
rect 1965 4206 3823 4207
rect 1965 4202 1975 4206
rect 1979 4202 2371 4206
rect 2375 4202 2571 4206
rect 2575 4202 2611 4206
rect 2615 4202 2763 4206
rect 2767 4202 2835 4206
rect 2839 4202 2955 4206
rect 2959 4202 3051 4206
rect 3055 4202 3139 4206
rect 3143 4202 3259 4206
rect 3263 4202 3315 4206
rect 3319 4202 3467 4206
rect 3471 4202 3491 4206
rect 3495 4202 3651 4206
rect 3655 4202 3799 4206
rect 3803 4202 3823 4206
rect 1965 4201 3823 4202
rect 3829 4201 3830 4207
rect 84 4189 85 4195
rect 91 4194 1947 4195
rect 91 4190 111 4194
rect 115 4190 727 4194
rect 731 4190 775 4194
rect 779 4190 863 4194
rect 867 4190 911 4194
rect 915 4190 999 4194
rect 1003 4190 1047 4194
rect 1051 4190 1135 4194
rect 1139 4190 1183 4194
rect 1187 4190 1271 4194
rect 1275 4190 1319 4194
rect 1323 4190 1407 4194
rect 1411 4190 1455 4194
rect 1459 4190 1543 4194
rect 1547 4190 1591 4194
rect 1595 4190 1679 4194
rect 1683 4190 1727 4194
rect 1731 4190 1815 4194
rect 1819 4190 1935 4194
rect 1939 4190 1947 4194
rect 91 4189 1947 4190
rect 1953 4189 1954 4195
rect 3822 4093 3823 4099
rect 3829 4098 5707 4099
rect 3829 4094 3839 4098
rect 3843 4094 4019 4098
rect 4023 4094 4195 4098
rect 4199 4094 4403 4098
rect 4407 4094 4651 4098
rect 4655 4094 4931 4098
rect 4935 4094 5227 4098
rect 5231 4094 5515 4098
rect 5519 4094 5663 4098
rect 5667 4094 5707 4098
rect 3829 4093 5707 4094
rect 5713 4093 5714 4099
rect 1946 4085 1947 4091
rect 1953 4090 3811 4091
rect 1953 4086 1975 4090
rect 1979 4086 2375 4090
rect 2379 4086 2399 4090
rect 2403 4086 2623 4090
rect 2627 4086 2639 4090
rect 2643 4086 2855 4090
rect 2859 4086 2863 4090
rect 2867 4086 3071 4090
rect 3075 4086 3079 4090
rect 3083 4086 3279 4090
rect 3283 4086 3287 4090
rect 3291 4086 3487 4090
rect 3491 4086 3495 4090
rect 3499 4086 3679 4090
rect 3683 4086 3799 4090
rect 3803 4086 3811 4090
rect 1953 4085 3811 4086
rect 3817 4085 3818 4091
rect 96 4065 97 4071
rect 103 4070 1959 4071
rect 103 4066 111 4070
rect 115 4066 627 4070
rect 631 4066 699 4070
rect 703 4066 763 4070
rect 767 4066 835 4070
rect 839 4066 899 4070
rect 903 4066 971 4070
rect 975 4066 1035 4070
rect 1039 4066 1107 4070
rect 1111 4066 1171 4070
rect 1175 4066 1243 4070
rect 1247 4066 1307 4070
rect 1311 4066 1379 4070
rect 1383 4066 1443 4070
rect 1447 4066 1515 4070
rect 1519 4066 1579 4070
rect 1583 4066 1651 4070
rect 1655 4066 1715 4070
rect 1719 4066 1787 4070
rect 1791 4066 1935 4070
rect 1939 4066 1959 4070
rect 103 4065 1959 4066
rect 1965 4065 1966 4071
rect 3810 3983 3811 3989
rect 3817 3983 3842 3989
rect 3836 3979 3842 3983
rect 1958 3973 1959 3979
rect 1965 3978 3823 3979
rect 1965 3974 1975 3978
rect 1979 3974 2323 3978
rect 2327 3974 2347 3978
rect 2351 3974 2571 3978
rect 2575 3974 2595 3978
rect 2599 3974 2803 3978
rect 2807 3974 2827 3978
rect 2831 3974 3027 3978
rect 3031 3974 3043 3978
rect 3047 3974 3243 3978
rect 3247 3974 3251 3978
rect 3255 3974 3459 3978
rect 3463 3974 3651 3978
rect 3655 3974 3799 3978
rect 3803 3974 3823 3978
rect 1965 3973 3823 3974
rect 3829 3973 3830 3979
rect 3836 3978 5695 3979
rect 3836 3974 3839 3978
rect 3843 3974 4183 3978
rect 4187 3974 4319 3978
rect 4323 3974 4455 3978
rect 4459 3974 4591 3978
rect 4595 3974 4727 3978
rect 4731 3974 4863 3978
rect 4867 3974 4999 3978
rect 5003 3974 5135 3978
rect 5139 3974 5271 3978
rect 5275 3974 5407 3978
rect 5411 3974 5543 3978
rect 5547 3974 5663 3978
rect 5667 3974 5695 3978
rect 3836 3973 5695 3974
rect 5701 3973 5702 3979
rect 84 3941 85 3947
rect 91 3946 1947 3947
rect 91 3942 111 3946
rect 115 3942 599 3946
rect 603 3942 655 3946
rect 659 3942 743 3946
rect 747 3942 791 3946
rect 795 3942 895 3946
rect 899 3942 927 3946
rect 931 3942 1047 3946
rect 1051 3942 1063 3946
rect 1067 3942 1199 3946
rect 1203 3942 1335 3946
rect 1339 3942 1359 3946
rect 1363 3942 1471 3946
rect 1475 3942 1519 3946
rect 1523 3942 1607 3946
rect 1611 3942 1679 3946
rect 1683 3942 1743 3946
rect 1747 3942 1935 3946
rect 1939 3942 1947 3946
rect 91 3941 1947 3942
rect 1953 3941 1954 3947
rect 1946 3857 1947 3863
rect 1953 3862 3811 3863
rect 1953 3858 1975 3862
rect 1979 3858 2239 3862
rect 2243 3858 2351 3862
rect 2355 3858 2479 3862
rect 2483 3858 2599 3862
rect 2603 3858 2703 3862
rect 2707 3858 2831 3862
rect 2835 3858 2919 3862
rect 2923 3858 3055 3862
rect 3059 3858 3119 3862
rect 3123 3858 3271 3862
rect 3275 3858 3311 3862
rect 3315 3858 3487 3862
rect 3491 3858 3503 3862
rect 3507 3858 3679 3862
rect 3683 3858 3799 3862
rect 3803 3858 3811 3862
rect 1953 3857 3811 3858
rect 3817 3857 3818 3863
rect 3822 3829 3823 3835
rect 3829 3834 5707 3835
rect 3829 3830 3839 3834
rect 3843 3830 4139 3834
rect 4143 3830 4155 3834
rect 4159 3830 4291 3834
rect 4295 3830 4323 3834
rect 4327 3830 4427 3834
rect 4431 3830 4531 3834
rect 4535 3830 4563 3834
rect 4567 3830 4699 3834
rect 4703 3830 4763 3834
rect 4767 3830 4835 3834
rect 4839 3830 4971 3834
rect 4975 3830 5011 3834
rect 5015 3830 5107 3834
rect 5111 3830 5243 3834
rect 5247 3830 5275 3834
rect 5279 3830 5379 3834
rect 5383 3830 5515 3834
rect 5519 3830 5663 3834
rect 5667 3830 5707 3834
rect 3829 3829 5707 3830
rect 5713 3829 5714 3835
rect 96 3821 97 3827
rect 103 3826 1959 3827
rect 103 3822 111 3826
rect 115 3822 427 3826
rect 431 3822 571 3826
rect 575 3822 587 3826
rect 591 3822 715 3826
rect 719 3822 755 3826
rect 759 3822 867 3826
rect 871 3822 923 3826
rect 927 3822 1019 3826
rect 1023 3822 1099 3826
rect 1103 3822 1171 3826
rect 1175 3822 1275 3826
rect 1279 3822 1331 3826
rect 1335 3822 1459 3826
rect 1463 3822 1491 3826
rect 1495 3822 1643 3826
rect 1647 3822 1651 3826
rect 1655 3822 1935 3826
rect 1939 3822 1959 3826
rect 103 3821 1959 3822
rect 1965 3821 1966 3827
rect 1958 3737 1959 3743
rect 1965 3742 3823 3743
rect 1965 3738 1975 3742
rect 1979 3738 2211 3742
rect 2215 3738 2227 3742
rect 2231 3738 2451 3742
rect 2455 3738 2667 3742
rect 2671 3738 2675 3742
rect 2679 3738 2875 3742
rect 2879 3738 2891 3742
rect 2895 3738 3075 3742
rect 3079 3738 3091 3742
rect 3095 3738 3275 3742
rect 3279 3738 3283 3742
rect 3287 3738 3475 3742
rect 3479 3738 3651 3742
rect 3655 3738 3799 3742
rect 3803 3738 3823 3742
rect 1965 3737 3823 3738
rect 3829 3737 3830 3743
rect 84 3697 85 3703
rect 91 3702 1947 3703
rect 91 3698 111 3702
rect 115 3698 327 3702
rect 331 3698 455 3702
rect 459 3698 495 3702
rect 499 3698 615 3702
rect 619 3698 679 3702
rect 683 3698 783 3702
rect 787 3698 863 3702
rect 867 3698 951 3702
rect 955 3698 1055 3702
rect 1059 3698 1127 3702
rect 1131 3698 1255 3702
rect 1259 3698 1303 3702
rect 1307 3698 1455 3702
rect 1459 3698 1487 3702
rect 1491 3698 1655 3702
rect 1659 3698 1671 3702
rect 1675 3698 1935 3702
rect 1939 3698 1947 3702
rect 91 3697 1947 3698
rect 1953 3697 1954 3703
rect 3810 3697 3811 3703
rect 3817 3702 5695 3703
rect 3817 3698 3839 3702
rect 3843 3698 4167 3702
rect 4171 3698 4303 3702
rect 4307 3698 4351 3702
rect 4355 3698 4479 3702
rect 4483 3698 4559 3702
rect 4563 3698 4671 3702
rect 4675 3698 4791 3702
rect 4795 3698 4879 3702
rect 4883 3698 5039 3702
rect 5043 3698 5103 3702
rect 5107 3698 5303 3702
rect 5307 3698 5335 3702
rect 5339 3698 5543 3702
rect 5547 3698 5663 3702
rect 5667 3698 5695 3702
rect 3817 3697 5695 3698
rect 5701 3697 5702 3703
rect 1946 3621 1947 3627
rect 1953 3626 3811 3627
rect 1953 3622 1975 3626
rect 1979 3622 2135 3626
rect 2139 3622 2255 3626
rect 2259 3622 2311 3626
rect 2315 3622 2479 3626
rect 2483 3622 2647 3626
rect 2651 3622 2695 3626
rect 2699 3622 2807 3626
rect 2811 3622 2903 3626
rect 2907 3622 2967 3626
rect 2971 3622 3103 3626
rect 3107 3622 3135 3626
rect 3139 3622 3303 3626
rect 3307 3622 3503 3626
rect 3507 3622 3799 3626
rect 3803 3622 3811 3626
rect 1953 3621 3811 3622
rect 3817 3621 3818 3627
rect 96 3565 97 3571
rect 103 3570 1959 3571
rect 103 3566 111 3570
rect 115 3566 203 3570
rect 207 3566 299 3570
rect 303 3566 379 3570
rect 383 3566 467 3570
rect 471 3566 563 3570
rect 567 3566 651 3570
rect 655 3566 755 3570
rect 759 3566 835 3570
rect 839 3566 955 3570
rect 959 3566 1027 3570
rect 1031 3566 1163 3570
rect 1167 3566 1227 3570
rect 1231 3566 1379 3570
rect 1383 3566 1427 3570
rect 1431 3566 1595 3570
rect 1599 3566 1627 3570
rect 1631 3566 1935 3570
rect 1939 3566 1959 3570
rect 103 3565 1959 3566
rect 1965 3565 1966 3571
rect 3822 3557 3823 3563
rect 3829 3562 5707 3563
rect 3829 3558 3839 3562
rect 3843 3558 4275 3562
rect 4279 3558 4451 3562
rect 4455 3558 4555 3562
rect 4559 3558 4643 3562
rect 4647 3558 4699 3562
rect 4703 3558 4851 3562
rect 4855 3558 5011 3562
rect 5015 3558 5075 3562
rect 5079 3558 5179 3562
rect 5183 3558 5307 3562
rect 5311 3558 5355 3562
rect 5359 3558 5515 3562
rect 5519 3558 5663 3562
rect 5667 3558 5707 3562
rect 3829 3557 5707 3558
rect 5713 3557 5714 3563
rect 1958 3485 1959 3491
rect 1965 3490 3823 3491
rect 1965 3486 1975 3490
rect 1979 3486 2035 3490
rect 2039 3486 2107 3490
rect 2111 3486 2187 3490
rect 2191 3486 2283 3490
rect 2287 3486 2339 3490
rect 2343 3486 2451 3490
rect 2455 3486 2491 3490
rect 2495 3486 2619 3490
rect 2623 3486 2643 3490
rect 2647 3486 2779 3490
rect 2783 3486 2795 3490
rect 2799 3486 2939 3490
rect 2943 3486 2947 3490
rect 2951 3486 3099 3490
rect 3103 3486 3107 3490
rect 3111 3486 3275 3490
rect 3279 3486 3799 3490
rect 3803 3486 3823 3490
rect 1965 3485 3823 3486
rect 3829 3485 3830 3491
rect 84 3433 85 3439
rect 91 3438 1947 3439
rect 91 3434 111 3438
rect 115 3434 231 3438
rect 235 3434 255 3438
rect 259 3434 407 3438
rect 411 3434 471 3438
rect 475 3434 591 3438
rect 595 3434 695 3438
rect 699 3434 783 3438
rect 787 3434 919 3438
rect 923 3434 983 3438
rect 987 3434 1143 3438
rect 1147 3434 1191 3438
rect 1195 3434 1367 3438
rect 1371 3434 1407 3438
rect 1411 3434 1591 3438
rect 1595 3434 1623 3438
rect 1627 3434 1935 3438
rect 1939 3434 1947 3438
rect 91 3433 1947 3434
rect 1953 3433 1954 3439
rect 3810 3433 3811 3439
rect 3817 3438 5695 3439
rect 3817 3434 3839 3438
rect 3843 3434 4583 3438
rect 4587 3434 4727 3438
rect 4731 3434 4879 3438
rect 4883 3434 4903 3438
rect 4907 3434 5039 3438
rect 5043 3434 5175 3438
rect 5179 3434 5207 3438
rect 5211 3434 5311 3438
rect 5315 3434 5383 3438
rect 5387 3434 5447 3438
rect 5451 3434 5543 3438
rect 5547 3434 5663 3438
rect 5667 3434 5695 3438
rect 3817 3433 5695 3434
rect 5701 3433 5702 3439
rect 1946 3361 1947 3367
rect 1953 3366 3811 3367
rect 1953 3362 1975 3366
rect 1979 3362 2023 3366
rect 2027 3362 2063 3366
rect 2067 3362 2191 3366
rect 2195 3362 2215 3366
rect 2219 3362 2367 3366
rect 2371 3362 2375 3366
rect 2379 3362 2519 3366
rect 2523 3362 2551 3366
rect 2555 3362 2671 3366
rect 2675 3362 2727 3366
rect 2731 3362 2823 3366
rect 2827 3362 2895 3366
rect 2899 3362 2975 3366
rect 2979 3362 3071 3366
rect 3075 3362 3127 3366
rect 3131 3362 3247 3366
rect 3251 3362 3799 3366
rect 3803 3362 3811 3366
rect 1953 3361 3811 3362
rect 3817 3361 3818 3367
rect 3822 3321 3823 3327
rect 3829 3326 5707 3327
rect 3829 3322 3839 3326
rect 3843 3322 4699 3326
rect 4703 3322 4835 3326
rect 4839 3322 4875 3326
rect 4879 3322 4971 3326
rect 4975 3322 5011 3326
rect 5015 3322 5107 3326
rect 5111 3322 5147 3326
rect 5151 3322 5243 3326
rect 5247 3322 5283 3326
rect 5287 3322 5379 3326
rect 5383 3322 5419 3326
rect 5423 3322 5515 3326
rect 5519 3322 5663 3326
rect 5667 3322 5707 3326
rect 3829 3321 5707 3322
rect 5713 3321 5714 3327
rect 96 3305 97 3311
rect 103 3310 1959 3311
rect 103 3306 111 3310
rect 115 3306 211 3310
rect 215 3306 227 3310
rect 231 3306 419 3310
rect 423 3306 443 3310
rect 447 3306 635 3310
rect 639 3306 667 3310
rect 671 3306 851 3310
rect 855 3306 891 3310
rect 895 3306 1075 3310
rect 1079 3306 1115 3310
rect 1119 3306 1299 3310
rect 1303 3306 1339 3310
rect 1343 3306 1523 3310
rect 1527 3306 1563 3310
rect 1567 3306 1935 3310
rect 1939 3306 1959 3310
rect 103 3305 1959 3306
rect 1965 3305 1966 3311
rect 1958 3245 1959 3251
rect 1965 3250 3823 3251
rect 1965 3246 1975 3250
rect 1979 3246 1995 3250
rect 1999 3246 2163 3250
rect 2167 3246 2211 3250
rect 2215 3246 2347 3250
rect 2351 3246 2435 3250
rect 2439 3246 2523 3250
rect 2527 3246 2651 3250
rect 2655 3246 2699 3250
rect 2703 3246 2851 3250
rect 2855 3246 2867 3250
rect 2871 3246 3043 3250
rect 3047 3246 3051 3250
rect 3055 3246 3219 3250
rect 3223 3246 3251 3250
rect 3255 3246 3451 3250
rect 3455 3246 3799 3250
rect 3803 3246 3823 3250
rect 1965 3245 3823 3246
rect 3829 3245 3830 3251
rect 3810 3201 3811 3207
rect 3817 3206 5695 3207
rect 3817 3202 3839 3206
rect 3843 3202 4567 3206
rect 4571 3202 4727 3206
rect 4731 3202 4743 3206
rect 4747 3202 4863 3206
rect 4867 3202 4935 3206
rect 4939 3202 4999 3206
rect 5003 3202 5135 3206
rect 5139 3202 5271 3206
rect 5275 3202 5351 3206
rect 5355 3202 5407 3206
rect 5411 3202 5543 3206
rect 5547 3202 5663 3206
rect 5667 3202 5695 3206
rect 3817 3201 5695 3202
rect 5701 3201 5702 3207
rect 84 3177 85 3183
rect 91 3182 1947 3183
rect 91 3178 111 3182
rect 115 3178 239 3182
rect 243 3178 303 3182
rect 307 3178 447 3182
rect 451 3178 543 3182
rect 547 3178 663 3182
rect 667 3178 783 3182
rect 787 3178 879 3182
rect 883 3178 1023 3182
rect 1027 3178 1103 3182
rect 1107 3178 1263 3182
rect 1267 3178 1327 3182
rect 1331 3178 1511 3182
rect 1515 3178 1551 3182
rect 1555 3178 1935 3182
rect 1939 3178 1947 3182
rect 91 3177 1947 3178
rect 1953 3177 1954 3183
rect 1946 3133 1947 3139
rect 1953 3138 3811 3139
rect 1953 3134 1975 3138
rect 1979 3134 2023 3138
rect 2027 3134 2239 3138
rect 2243 3134 2327 3138
rect 2331 3134 2463 3138
rect 2467 3134 2631 3138
rect 2635 3134 2679 3138
rect 2683 3134 2879 3138
rect 2883 3134 2911 3138
rect 2915 3134 3079 3138
rect 3083 3134 3175 3138
rect 3179 3134 3279 3138
rect 3283 3134 3439 3138
rect 3443 3134 3479 3138
rect 3483 3134 3679 3138
rect 3683 3134 3799 3138
rect 3803 3134 3811 3138
rect 1953 3133 3811 3134
rect 3817 3133 3818 3139
rect 3822 3085 3823 3091
rect 3829 3090 5707 3091
rect 3829 3086 3839 3090
rect 3843 3086 4307 3090
rect 4311 3086 4483 3090
rect 4487 3086 4539 3090
rect 4543 3086 4675 3090
rect 4679 3086 4715 3090
rect 4719 3086 4875 3090
rect 4879 3086 4907 3090
rect 4911 3086 5091 3090
rect 5095 3086 5107 3090
rect 5111 3086 5315 3090
rect 5319 3086 5323 3090
rect 5327 3086 5515 3090
rect 5519 3086 5663 3090
rect 5667 3086 5707 3090
rect 3829 3085 5707 3086
rect 5713 3085 5714 3091
rect 96 3065 97 3071
rect 103 3070 1959 3071
rect 103 3066 111 3070
rect 115 3066 275 3070
rect 279 3066 355 3070
rect 359 3066 515 3070
rect 519 3066 627 3070
rect 631 3066 755 3070
rect 759 3066 883 3070
rect 887 3066 995 3070
rect 999 3066 1123 3070
rect 1127 3066 1235 3070
rect 1239 3066 1355 3070
rect 1359 3066 1483 3070
rect 1487 3066 1579 3070
rect 1583 3066 1787 3070
rect 1791 3066 1935 3070
rect 1939 3066 1959 3070
rect 103 3065 1959 3066
rect 1965 3065 1966 3071
rect 1958 3013 1959 3019
rect 1965 3018 3823 3019
rect 1965 3014 1975 3018
rect 1979 3014 1995 3018
rect 1999 3014 2299 3018
rect 2303 3014 2603 3018
rect 2607 3014 2883 3018
rect 2887 3014 3107 3018
rect 3111 3014 3147 3018
rect 3151 3014 3243 3018
rect 3247 3014 3379 3018
rect 3383 3014 3411 3018
rect 3415 3014 3515 3018
rect 3519 3014 3651 3018
rect 3655 3014 3799 3018
rect 3803 3014 3823 3018
rect 1965 3013 3823 3014
rect 3829 3013 3830 3019
rect 3810 2969 3811 2975
rect 3817 2974 5695 2975
rect 3817 2970 3839 2974
rect 3843 2970 3887 2974
rect 3891 2970 4023 2974
rect 4027 2970 4175 2974
rect 4179 2970 4335 2974
rect 4339 2970 4391 2974
rect 4395 2970 4511 2974
rect 4515 2970 4639 2974
rect 4643 2970 4703 2974
rect 4707 2970 4903 2974
rect 4907 2970 4919 2974
rect 4923 2970 5119 2974
rect 5123 2970 5223 2974
rect 5227 2970 5343 2974
rect 5347 2970 5527 2974
rect 5531 2970 5543 2974
rect 5547 2970 5663 2974
rect 5667 2970 5695 2974
rect 3817 2969 5695 2970
rect 5701 2969 5702 2975
rect 84 2953 85 2959
rect 91 2958 1947 2959
rect 91 2954 111 2958
rect 115 2954 343 2958
rect 347 2954 383 2958
rect 387 2954 551 2958
rect 555 2954 655 2958
rect 659 2954 759 2958
rect 763 2954 911 2958
rect 915 2954 951 2958
rect 955 2954 1135 2958
rect 1139 2954 1151 2958
rect 1155 2954 1311 2958
rect 1315 2954 1383 2958
rect 1387 2954 1487 2958
rect 1491 2954 1607 2958
rect 1611 2954 1663 2958
rect 1667 2954 1815 2958
rect 1819 2954 1935 2958
rect 1939 2954 1947 2958
rect 91 2953 1947 2954
rect 1953 2953 1954 2959
rect 3822 2857 3823 2863
rect 3829 2862 5707 2863
rect 3829 2858 3839 2862
rect 3843 2858 3859 2862
rect 3863 2858 3995 2862
rect 3999 2858 4131 2862
rect 4135 2858 4147 2862
rect 4151 2858 4267 2862
rect 4271 2858 4363 2862
rect 4367 2858 4403 2862
rect 4407 2858 4539 2862
rect 4543 2858 4611 2862
rect 4615 2858 4675 2862
rect 4679 2858 4811 2862
rect 4815 2858 4891 2862
rect 4895 2858 5195 2862
rect 5199 2858 5499 2862
rect 5503 2858 5663 2862
rect 5667 2858 5707 2862
rect 3829 2857 5707 2858
rect 5713 2857 5714 2863
rect 96 2829 97 2835
rect 103 2834 1959 2835
rect 103 2830 111 2834
rect 115 2830 315 2834
rect 319 2830 363 2834
rect 367 2830 523 2834
rect 527 2830 563 2834
rect 567 2830 731 2834
rect 735 2830 755 2834
rect 759 2830 923 2834
rect 927 2830 939 2834
rect 943 2830 1107 2834
rect 1111 2830 1115 2834
rect 1119 2830 1283 2834
rect 1287 2830 1451 2834
rect 1455 2830 1459 2834
rect 1463 2830 1619 2834
rect 1623 2830 1635 2834
rect 1639 2830 1787 2834
rect 1791 2830 1935 2834
rect 1939 2830 1959 2834
rect 103 2829 1959 2830
rect 1965 2829 1966 2835
rect 3810 2729 3811 2735
rect 3817 2734 5695 2735
rect 3817 2730 3839 2734
rect 3843 2730 3887 2734
rect 3891 2730 4023 2734
rect 4027 2730 4159 2734
rect 4163 2730 4295 2734
rect 4299 2730 4431 2734
rect 4435 2730 4567 2734
rect 4571 2730 4703 2734
rect 4707 2730 4711 2734
rect 4715 2730 4839 2734
rect 4843 2730 4879 2734
rect 4883 2730 5063 2734
rect 5067 2730 5255 2734
rect 5259 2730 5447 2734
rect 5451 2730 5663 2734
rect 5667 2730 5695 2734
rect 3817 2729 5695 2730
rect 5701 2729 5702 2735
rect 84 2713 85 2719
rect 91 2718 1947 2719
rect 91 2714 111 2718
rect 115 2714 391 2718
rect 395 2714 447 2718
rect 451 2714 591 2718
rect 595 2714 615 2718
rect 619 2714 775 2718
rect 779 2714 783 2718
rect 787 2714 935 2718
rect 939 2714 967 2718
rect 971 2714 1087 2718
rect 1091 2714 1143 2718
rect 1147 2714 1239 2718
rect 1243 2714 1311 2718
rect 1315 2714 1383 2718
rect 1387 2714 1479 2718
rect 1483 2714 1535 2718
rect 1539 2714 1647 2718
rect 1651 2714 1679 2718
rect 1683 2714 1815 2718
rect 1819 2714 1935 2718
rect 1939 2714 1947 2718
rect 91 2713 1947 2714
rect 1953 2713 1954 2719
rect 1946 2633 1947 2639
rect 1953 2638 3811 2639
rect 1953 2634 1975 2638
rect 1979 2634 3135 2638
rect 3139 2634 3271 2638
rect 3275 2634 3407 2638
rect 3411 2634 3543 2638
rect 3547 2634 3679 2638
rect 3683 2634 3799 2638
rect 3803 2634 3811 2638
rect 1953 2633 3811 2634
rect 3817 2633 3818 2639
rect 96 2597 97 2603
rect 103 2602 1959 2603
rect 103 2598 111 2602
rect 115 2598 235 2602
rect 239 2598 419 2602
rect 423 2598 435 2602
rect 439 2598 587 2602
rect 591 2598 627 2602
rect 631 2598 747 2602
rect 751 2598 811 2602
rect 815 2598 907 2602
rect 911 2598 987 2602
rect 991 2598 1059 2602
rect 1063 2598 1155 2602
rect 1159 2598 1211 2602
rect 1215 2598 1323 2602
rect 1327 2598 1355 2602
rect 1359 2598 1483 2602
rect 1487 2598 1507 2602
rect 1511 2598 1643 2602
rect 1647 2598 1651 2602
rect 1655 2598 1787 2602
rect 1791 2598 1935 2602
rect 1939 2598 1959 2602
rect 103 2597 1959 2598
rect 1965 2597 1966 2603
rect 3822 2601 3823 2607
rect 3829 2606 5707 2607
rect 3829 2602 3839 2606
rect 3843 2602 3859 2606
rect 3863 2602 3995 2606
rect 3999 2602 4131 2606
rect 4135 2602 4179 2606
rect 4183 2602 4267 2606
rect 4271 2602 4395 2606
rect 4399 2602 4403 2606
rect 4407 2602 4539 2606
rect 4543 2602 4643 2606
rect 4647 2602 4683 2606
rect 4687 2602 4851 2606
rect 4855 2602 4907 2606
rect 4911 2602 5035 2606
rect 5039 2602 5187 2606
rect 5191 2602 5227 2606
rect 5231 2602 5419 2606
rect 5423 2602 5467 2606
rect 5471 2602 5663 2606
rect 5667 2602 5707 2606
rect 3829 2601 5707 2602
rect 5713 2601 5714 2607
rect 1958 2521 1959 2527
rect 1965 2526 3823 2527
rect 1965 2522 1975 2526
rect 1979 2522 1995 2526
rect 1999 2522 2251 2526
rect 2255 2522 2523 2526
rect 2527 2522 2771 2526
rect 2775 2522 3003 2526
rect 3007 2522 3227 2526
rect 3231 2522 3243 2526
rect 3247 2522 3379 2526
rect 3383 2522 3451 2526
rect 3455 2522 3515 2526
rect 3519 2522 3651 2526
rect 3655 2522 3799 2526
rect 3803 2522 3823 2526
rect 1965 2521 3823 2522
rect 3829 2521 3830 2527
rect 3810 2489 3811 2495
rect 3817 2494 5695 2495
rect 3817 2490 3839 2494
rect 3843 2490 4207 2494
rect 4211 2490 4423 2494
rect 4427 2490 4535 2494
rect 4539 2490 4671 2494
rect 4675 2490 4759 2494
rect 4763 2490 4935 2494
rect 4939 2490 4983 2494
rect 4987 2490 5215 2494
rect 5219 2490 5447 2494
rect 5451 2490 5495 2494
rect 5499 2490 5663 2494
rect 5667 2490 5695 2494
rect 3817 2489 5695 2490
rect 5701 2489 5702 2495
rect 84 2477 85 2483
rect 91 2482 1947 2483
rect 91 2478 111 2482
rect 115 2478 223 2482
rect 227 2478 263 2482
rect 267 2478 423 2482
rect 427 2478 463 2482
rect 467 2478 623 2482
rect 627 2478 655 2482
rect 659 2478 815 2482
rect 819 2478 839 2482
rect 843 2478 1015 2482
rect 1019 2478 1183 2482
rect 1187 2478 1215 2482
rect 1219 2478 1351 2482
rect 1355 2478 1511 2482
rect 1515 2478 1671 2482
rect 1675 2478 1815 2482
rect 1819 2478 1935 2482
rect 1939 2478 1947 2482
rect 91 2477 1947 2478
rect 1953 2477 1954 2483
rect 1946 2409 1947 2415
rect 1953 2414 3811 2415
rect 1953 2410 1975 2414
rect 1979 2410 2023 2414
rect 2027 2410 2055 2414
rect 2059 2410 2215 2414
rect 2219 2410 2279 2414
rect 2283 2410 2375 2414
rect 2379 2410 2543 2414
rect 2547 2410 2551 2414
rect 2555 2410 2711 2414
rect 2715 2410 2799 2414
rect 2803 2410 2871 2414
rect 2875 2410 3031 2414
rect 3035 2410 3191 2414
rect 3195 2410 3255 2414
rect 3259 2410 3359 2414
rect 3363 2410 3479 2414
rect 3483 2410 3527 2414
rect 3531 2410 3679 2414
rect 3683 2410 3799 2414
rect 3803 2410 3811 2414
rect 1953 2409 3811 2410
rect 3817 2409 3818 2415
rect 3822 2377 3823 2383
rect 3829 2382 5707 2383
rect 3829 2378 3839 2382
rect 3843 2378 4507 2382
rect 4511 2378 4707 2382
rect 4711 2378 4731 2382
rect 4735 2378 4867 2382
rect 4871 2378 4955 2382
rect 4959 2378 5027 2382
rect 5031 2378 5187 2382
rect 5191 2378 5347 2382
rect 5351 2378 5419 2382
rect 5423 2378 5515 2382
rect 5519 2378 5663 2382
rect 5667 2378 5707 2382
rect 3829 2377 5707 2378
rect 5713 2377 5714 2383
rect 96 2353 97 2359
rect 103 2358 1959 2359
rect 103 2354 111 2358
rect 115 2354 131 2358
rect 135 2354 195 2358
rect 199 2354 291 2358
rect 295 2354 395 2358
rect 399 2354 483 2358
rect 487 2354 595 2358
rect 599 2354 675 2358
rect 679 2354 787 2358
rect 791 2354 867 2358
rect 871 2354 987 2358
rect 991 2354 1187 2358
rect 1191 2354 1935 2358
rect 1939 2354 1959 2358
rect 103 2353 1959 2354
rect 1965 2353 1966 2359
rect 1958 2289 1959 2295
rect 1965 2294 3823 2295
rect 1965 2290 1975 2294
rect 1979 2290 2027 2294
rect 2031 2290 2139 2294
rect 2143 2290 2187 2294
rect 2191 2290 2275 2294
rect 2279 2290 2347 2294
rect 2351 2290 2411 2294
rect 2415 2290 2515 2294
rect 2519 2290 2547 2294
rect 2551 2290 2683 2294
rect 2687 2290 2819 2294
rect 2823 2290 2843 2294
rect 2847 2290 2955 2294
rect 2959 2290 3003 2294
rect 3007 2290 3091 2294
rect 3095 2290 3163 2294
rect 3167 2290 3227 2294
rect 3231 2290 3331 2294
rect 3335 2290 3363 2294
rect 3367 2290 3499 2294
rect 3503 2290 3799 2294
rect 3803 2290 3823 2294
rect 1965 2289 3823 2290
rect 3829 2289 3830 2295
rect 3810 2253 3811 2259
rect 3817 2258 5695 2259
rect 3817 2254 3839 2258
rect 3843 2254 4735 2258
rect 4739 2254 4887 2258
rect 4891 2254 4895 2258
rect 4899 2254 5047 2258
rect 5051 2254 5055 2258
rect 5059 2254 5215 2258
rect 5219 2254 5375 2258
rect 5379 2254 5391 2258
rect 5395 2254 5543 2258
rect 5547 2254 5663 2258
rect 5667 2254 5695 2258
rect 3817 2253 5695 2254
rect 5701 2253 5702 2259
rect 84 2241 85 2247
rect 91 2246 1947 2247
rect 91 2242 111 2246
rect 115 2242 159 2246
rect 163 2242 295 2246
rect 299 2242 319 2246
rect 323 2242 439 2246
rect 443 2242 511 2246
rect 515 2242 591 2246
rect 595 2242 703 2246
rect 707 2242 743 2246
rect 747 2242 895 2246
rect 899 2242 1935 2246
rect 1939 2242 1947 2246
rect 91 2241 1947 2242
rect 1953 2241 1954 2247
rect 1946 2173 1947 2179
rect 1953 2178 3811 2179
rect 1953 2174 1975 2178
rect 1979 2174 2023 2178
rect 2027 2174 2159 2178
rect 2163 2174 2167 2178
rect 2171 2174 2295 2178
rect 2299 2174 2303 2178
rect 2307 2174 2431 2178
rect 2435 2174 2439 2178
rect 2443 2174 2567 2178
rect 2571 2174 2575 2178
rect 2579 2174 2703 2178
rect 2707 2174 2711 2178
rect 2715 2174 2839 2178
rect 2843 2174 2847 2178
rect 2851 2174 2975 2178
rect 2979 2174 2983 2178
rect 2987 2174 3111 2178
rect 3115 2174 3119 2178
rect 3123 2174 3247 2178
rect 3251 2174 3255 2178
rect 3259 2174 3391 2178
rect 3395 2174 3799 2178
rect 3803 2174 3811 2178
rect 1953 2173 3811 2174
rect 3817 2173 3818 2179
rect 96 2129 97 2135
rect 103 2134 1959 2135
rect 103 2130 111 2134
rect 115 2130 131 2134
rect 135 2130 267 2134
rect 271 2130 331 2134
rect 335 2130 411 2134
rect 415 2130 555 2134
rect 559 2130 563 2134
rect 567 2130 715 2134
rect 719 2130 779 2134
rect 783 2130 1011 2134
rect 1015 2130 1935 2134
rect 1939 2130 1959 2134
rect 103 2129 1959 2130
rect 1965 2129 1966 2135
rect 3822 2133 3823 2139
rect 3829 2138 5707 2139
rect 3829 2134 3839 2138
rect 3843 2134 4707 2138
rect 4711 2134 4787 2138
rect 4791 2134 4859 2138
rect 4863 2134 4923 2138
rect 4927 2134 5019 2138
rect 5023 2134 5067 2138
rect 5071 2134 5187 2138
rect 5191 2134 5219 2138
rect 5223 2134 5363 2138
rect 5367 2134 5379 2138
rect 5383 2134 5515 2138
rect 5519 2134 5663 2138
rect 5667 2134 5707 2138
rect 3829 2133 5707 2134
rect 5713 2133 5714 2139
rect 1958 2053 1959 2059
rect 1965 2058 3823 2059
rect 1965 2054 1975 2058
rect 1979 2054 1995 2058
rect 1999 2054 2131 2058
rect 2135 2054 2267 2058
rect 2271 2054 2403 2058
rect 2407 2054 2539 2058
rect 2543 2054 2675 2058
rect 2679 2054 2811 2058
rect 2815 2054 2947 2058
rect 2951 2054 3083 2058
rect 3087 2054 3091 2058
rect 3095 2054 3219 2058
rect 3223 2054 3243 2058
rect 3247 2054 3395 2058
rect 3399 2054 3799 2058
rect 3803 2054 3823 2058
rect 1965 2053 3823 2054
rect 3829 2053 3830 2059
rect 84 2013 85 2019
rect 91 2018 1947 2019
rect 91 2014 111 2018
rect 115 2014 159 2018
rect 163 2014 359 2018
rect 363 2014 463 2018
rect 467 2014 583 2018
rect 587 2014 799 2018
rect 803 2014 807 2018
rect 811 2014 1039 2018
rect 1043 2014 1143 2018
rect 1147 2014 1487 2018
rect 1491 2014 1815 2018
rect 1819 2014 1935 2018
rect 1939 2014 1947 2018
rect 91 2013 1947 2014
rect 1953 2013 1954 2019
rect 3810 2017 3811 2023
rect 3817 2022 5695 2023
rect 3817 2018 3839 2022
rect 3843 2018 4815 2022
rect 4819 2018 4863 2022
rect 4867 2018 4951 2022
rect 4955 2018 4999 2022
rect 5003 2018 5095 2022
rect 5099 2018 5135 2022
rect 5139 2018 5247 2022
rect 5251 2018 5271 2022
rect 5275 2018 5407 2022
rect 5411 2018 5543 2022
rect 5547 2018 5663 2022
rect 5667 2018 5695 2022
rect 3817 2017 5695 2018
rect 5701 2017 5702 2023
rect 1946 1933 1947 1939
rect 1953 1938 3811 1939
rect 1953 1934 1975 1938
rect 1979 1934 2023 1938
rect 2027 1934 2159 1938
rect 2163 1934 2295 1938
rect 2299 1934 2431 1938
rect 2435 1934 2527 1938
rect 2531 1934 2567 1938
rect 2571 1934 2663 1938
rect 2667 1934 2703 1938
rect 2707 1934 2799 1938
rect 2803 1934 2839 1938
rect 2843 1934 2935 1938
rect 2939 1934 2975 1938
rect 2979 1934 3071 1938
rect 3075 1934 3119 1938
rect 3123 1934 3207 1938
rect 3211 1934 3271 1938
rect 3275 1934 3351 1938
rect 3355 1934 3423 1938
rect 3427 1934 3799 1938
rect 3803 1934 3811 1938
rect 1953 1933 3811 1934
rect 3817 1933 3818 1939
rect 96 1901 97 1907
rect 103 1906 1959 1907
rect 103 1902 111 1906
rect 115 1902 131 1906
rect 135 1902 195 1906
rect 199 1902 435 1906
rect 439 1902 451 1906
rect 455 1902 699 1906
rect 703 1902 771 1906
rect 775 1902 931 1906
rect 935 1902 1115 1906
rect 1119 1902 1155 1906
rect 1159 1902 1371 1906
rect 1375 1902 1459 1906
rect 1463 1902 1587 1906
rect 1591 1902 1787 1906
rect 1791 1902 1935 1906
rect 1939 1902 1959 1906
rect 103 1901 1959 1902
rect 1965 1901 1966 1907
rect 3822 1901 3823 1907
rect 3829 1906 5707 1907
rect 3829 1902 3839 1906
rect 3843 1902 4683 1906
rect 4687 1902 4835 1906
rect 4839 1902 4843 1906
rect 4847 1902 4971 1906
rect 4975 1902 5011 1906
rect 5015 1902 5107 1906
rect 5111 1902 5179 1906
rect 5183 1902 5243 1906
rect 5247 1902 5355 1906
rect 5359 1902 5379 1906
rect 5383 1902 5515 1906
rect 5519 1902 5663 1906
rect 5667 1902 5707 1906
rect 3829 1901 5707 1902
rect 5713 1901 5714 1907
rect 1958 1821 1959 1827
rect 1965 1826 3823 1827
rect 1965 1822 1975 1826
rect 1979 1822 2443 1826
rect 2447 1822 2499 1826
rect 2503 1822 2587 1826
rect 2591 1822 2635 1826
rect 2639 1822 2739 1826
rect 2743 1822 2771 1826
rect 2775 1822 2891 1826
rect 2895 1822 2907 1826
rect 2911 1822 3043 1826
rect 3047 1822 3179 1826
rect 3183 1822 3195 1826
rect 3199 1822 3323 1826
rect 3327 1822 3799 1826
rect 3803 1822 3823 1826
rect 1965 1821 3823 1822
rect 3829 1821 3830 1827
rect 84 1785 85 1791
rect 91 1790 1947 1791
rect 91 1786 111 1790
rect 115 1786 223 1790
rect 227 1786 231 1790
rect 235 1786 447 1790
rect 451 1786 479 1790
rect 483 1786 671 1790
rect 675 1786 727 1790
rect 731 1786 895 1790
rect 899 1786 959 1790
rect 963 1786 1119 1790
rect 1123 1786 1183 1790
rect 1187 1786 1343 1790
rect 1347 1786 1399 1790
rect 1403 1786 1567 1790
rect 1571 1786 1615 1790
rect 1619 1786 1799 1790
rect 1803 1786 1815 1790
rect 1819 1786 1935 1790
rect 1939 1786 1947 1790
rect 91 1785 1947 1786
rect 1953 1785 1954 1791
rect 3810 1785 3811 1791
rect 3817 1790 5695 1791
rect 3817 1786 3839 1790
rect 3843 1786 3887 1790
rect 3891 1786 4023 1790
rect 4027 1786 4191 1790
rect 4195 1786 4367 1790
rect 4371 1786 4559 1790
rect 4563 1786 4711 1790
rect 4715 1786 4767 1790
rect 4771 1786 4871 1790
rect 4875 1786 4983 1790
rect 4987 1786 5039 1790
rect 5043 1786 5207 1790
rect 5211 1786 5215 1790
rect 5219 1786 5383 1790
rect 5387 1786 5447 1790
rect 5451 1786 5543 1790
rect 5547 1786 5663 1790
rect 5667 1786 5695 1790
rect 3817 1785 5695 1786
rect 5701 1785 5702 1791
rect 1946 1683 1947 1689
rect 1953 1683 1978 1689
rect 96 1673 97 1679
rect 103 1678 1959 1679
rect 103 1674 111 1678
rect 115 1674 203 1678
rect 207 1674 275 1678
rect 279 1674 419 1678
rect 423 1674 459 1678
rect 463 1674 643 1678
rect 647 1674 667 1678
rect 671 1674 867 1678
rect 871 1674 883 1678
rect 887 1674 1091 1678
rect 1095 1674 1115 1678
rect 1119 1674 1315 1678
rect 1319 1674 1355 1678
rect 1359 1674 1539 1678
rect 1543 1674 1595 1678
rect 1599 1674 1771 1678
rect 1775 1674 1935 1678
rect 1939 1674 1959 1678
rect 103 1673 1959 1674
rect 1965 1673 1966 1679
rect 1972 1671 1978 1683
rect 3822 1673 3823 1679
rect 3829 1678 5707 1679
rect 3829 1674 3839 1678
rect 3843 1674 3859 1678
rect 3863 1674 3995 1678
rect 3999 1674 4131 1678
rect 4135 1674 4163 1678
rect 4167 1674 4283 1678
rect 4287 1674 4339 1678
rect 4343 1674 4483 1678
rect 4487 1674 4531 1678
rect 4535 1674 4715 1678
rect 4719 1674 4739 1678
rect 4743 1674 4955 1678
rect 4959 1674 4979 1678
rect 4983 1674 5187 1678
rect 5191 1674 5259 1678
rect 5263 1674 5419 1678
rect 5423 1674 5515 1678
rect 5519 1674 5663 1678
rect 5667 1674 5707 1678
rect 3829 1673 5707 1674
rect 5713 1673 5714 1679
rect 1972 1670 3811 1671
rect 1972 1666 1975 1670
rect 1979 1666 2231 1670
rect 2235 1666 2471 1670
rect 2475 1666 2599 1670
rect 2603 1666 2615 1670
rect 2619 1666 2767 1670
rect 2771 1666 2919 1670
rect 2923 1666 2967 1670
rect 2971 1666 3071 1670
rect 3075 1666 3223 1670
rect 3227 1666 3335 1670
rect 3339 1666 3679 1670
rect 3683 1666 3799 1670
rect 3803 1666 3811 1670
rect 1972 1665 3811 1666
rect 3817 1665 3818 1671
rect 84 1561 85 1567
rect 91 1566 1947 1567
rect 91 1562 111 1566
rect 115 1562 303 1566
rect 307 1562 383 1566
rect 387 1562 487 1566
rect 491 1562 575 1566
rect 579 1562 695 1566
rect 699 1562 767 1566
rect 771 1562 911 1566
rect 915 1562 951 1566
rect 955 1562 1127 1566
rect 1131 1562 1143 1566
rect 1147 1562 1303 1566
rect 1307 1562 1383 1566
rect 1387 1562 1479 1566
rect 1483 1562 1623 1566
rect 1627 1562 1663 1566
rect 1667 1562 1935 1566
rect 1939 1562 1947 1566
rect 91 1561 1947 1562
rect 1953 1561 1954 1567
rect 3810 1561 3811 1567
rect 3817 1566 5695 1567
rect 3817 1562 3839 1566
rect 3843 1562 3887 1566
rect 3891 1562 4023 1566
rect 4027 1562 4047 1566
rect 4051 1562 4159 1566
rect 4163 1562 4271 1566
rect 4275 1562 4311 1566
rect 4315 1562 4511 1566
rect 4515 1562 4543 1566
rect 4547 1562 4743 1566
rect 4747 1562 4855 1566
rect 4859 1562 5007 1566
rect 5011 1562 5191 1566
rect 5195 1562 5287 1566
rect 5291 1562 5527 1566
rect 5531 1562 5543 1566
rect 5547 1562 5663 1566
rect 5667 1562 5695 1566
rect 3817 1561 5695 1562
rect 5701 1561 5702 1567
rect 1958 1541 1959 1547
rect 1965 1546 3823 1547
rect 1965 1542 1975 1546
rect 1979 1542 1995 1546
rect 1999 1542 2203 1546
rect 2207 1542 2275 1546
rect 2279 1542 2539 1546
rect 2543 1542 2571 1546
rect 2575 1542 2779 1546
rect 2783 1542 2939 1546
rect 2943 1542 3011 1546
rect 3015 1542 3235 1546
rect 3239 1542 3307 1546
rect 3311 1542 3451 1546
rect 3455 1542 3651 1546
rect 3655 1542 3799 1546
rect 3803 1542 3823 1546
rect 1965 1541 3823 1542
rect 3829 1541 3830 1547
rect 1946 1439 1947 1445
rect 1953 1439 1978 1445
rect 1972 1435 1978 1439
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 331 1434
rect 335 1430 355 1434
rect 359 1430 547 1434
rect 551 1430 587 1434
rect 591 1430 739 1434
rect 743 1430 843 1434
rect 847 1430 923 1434
rect 927 1430 1099 1434
rect 1103 1430 1275 1434
rect 1279 1430 1363 1434
rect 1367 1430 1451 1434
rect 1455 1430 1635 1434
rect 1639 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 1972 1434 3811 1435
rect 1972 1430 1975 1434
rect 1979 1430 2023 1434
rect 2027 1430 2191 1434
rect 2195 1430 2303 1434
rect 2307 1430 2399 1434
rect 2403 1430 2567 1434
rect 2571 1430 2615 1434
rect 2619 1430 2807 1434
rect 2811 1430 2831 1434
rect 2835 1430 3039 1434
rect 3043 1430 3055 1434
rect 3059 1430 3263 1434
rect 3267 1430 3287 1434
rect 3291 1430 3479 1434
rect 3483 1430 3527 1434
rect 3531 1430 3679 1434
rect 3683 1430 3799 1434
rect 3803 1430 3811 1434
rect 1972 1429 3811 1430
rect 3817 1429 3818 1435
rect 3822 1433 3823 1439
rect 3829 1438 5707 1439
rect 3829 1434 3839 1438
rect 3843 1434 3859 1438
rect 3863 1434 3995 1438
rect 3999 1434 4019 1438
rect 4023 1434 4147 1438
rect 4151 1434 4243 1438
rect 4247 1434 4355 1438
rect 4359 1434 4515 1438
rect 4519 1434 4595 1438
rect 4599 1434 4827 1438
rect 4831 1434 4867 1438
rect 4871 1434 5163 1438
rect 5167 1434 5459 1438
rect 5463 1434 5499 1438
rect 5503 1434 5663 1438
rect 5667 1434 5707 1438
rect 3829 1433 5707 1434
rect 5713 1433 5714 1439
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 359 1322
rect 363 1318 367 1322
rect 371 1318 551 1322
rect 555 1318 615 1322
rect 619 1318 727 1322
rect 731 1318 871 1322
rect 875 1318 895 1322
rect 899 1318 1063 1322
rect 1067 1318 1127 1322
rect 1131 1318 1223 1322
rect 1227 1318 1375 1322
rect 1379 1318 1391 1322
rect 1395 1318 1527 1322
rect 1531 1318 1679 1322
rect 1683 1318 1815 1322
rect 1819 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 3810 1317 3811 1323
rect 3817 1322 5695 1323
rect 3817 1318 3839 1322
rect 3843 1318 3887 1322
rect 3891 1318 4023 1322
rect 4027 1318 4047 1322
rect 4051 1318 4175 1322
rect 4179 1318 4239 1322
rect 4243 1318 4383 1322
rect 4387 1318 4455 1322
rect 4459 1318 4623 1322
rect 4627 1318 4695 1322
rect 4699 1318 4895 1322
rect 4899 1318 4951 1322
rect 4955 1318 5191 1322
rect 5195 1318 5223 1322
rect 5227 1318 5487 1322
rect 5491 1318 5495 1322
rect 5499 1318 5663 1322
rect 5667 1318 5695 1322
rect 3817 1317 5695 1318
rect 5701 1317 5702 1323
rect 1958 1297 1959 1303
rect 1965 1302 3823 1303
rect 1965 1298 1975 1302
rect 1979 1298 1995 1302
rect 1999 1298 2163 1302
rect 2167 1298 2371 1302
rect 2375 1298 2587 1302
rect 2591 1298 2803 1302
rect 2807 1298 3027 1302
rect 3031 1298 3091 1302
rect 3095 1298 3227 1302
rect 3231 1298 3259 1302
rect 3263 1298 3363 1302
rect 3367 1298 3499 1302
rect 3503 1298 3799 1302
rect 3803 1298 3823 1302
rect 1965 1297 3823 1298
rect 3829 1297 3830 1303
rect 1946 1203 1947 1209
rect 1953 1203 1978 1209
rect 96 1193 97 1199
rect 103 1198 1959 1199
rect 103 1194 111 1198
rect 115 1194 235 1198
rect 239 1194 339 1198
rect 343 1194 379 1198
rect 383 1194 523 1198
rect 527 1194 667 1198
rect 671 1194 699 1198
rect 703 1194 811 1198
rect 815 1194 867 1198
rect 871 1194 947 1198
rect 951 1194 1035 1198
rect 1039 1194 1091 1198
rect 1095 1194 1195 1198
rect 1199 1194 1235 1198
rect 1239 1194 1347 1198
rect 1351 1194 1379 1198
rect 1383 1194 1499 1198
rect 1503 1194 1515 1198
rect 1519 1194 1651 1198
rect 1655 1194 1787 1198
rect 1791 1194 1935 1198
rect 1939 1194 1959 1198
rect 103 1193 1959 1194
rect 1965 1193 1966 1199
rect 1972 1191 1978 1203
rect 3822 1197 3823 1203
rect 3829 1202 5707 1203
rect 3829 1198 3839 1202
rect 3843 1198 3859 1202
rect 3863 1198 4019 1202
rect 4023 1198 4091 1202
rect 4095 1198 4211 1202
rect 4215 1198 4339 1202
rect 4343 1198 4427 1202
rect 4431 1198 4579 1202
rect 4583 1198 4667 1202
rect 4671 1198 4811 1202
rect 4815 1198 4923 1202
rect 4927 1198 5043 1202
rect 5047 1198 5195 1202
rect 5199 1198 5275 1202
rect 5279 1198 5467 1202
rect 5471 1198 5515 1202
rect 5519 1198 5663 1202
rect 5667 1198 5707 1202
rect 3829 1197 5707 1198
rect 5713 1197 5714 1203
rect 1972 1190 3811 1191
rect 1972 1186 1975 1190
rect 1979 1186 2983 1190
rect 2987 1186 3119 1190
rect 3123 1186 3255 1190
rect 3259 1186 3391 1190
rect 3395 1186 3799 1190
rect 3803 1186 3811 1190
rect 1972 1185 3811 1186
rect 3817 1185 3818 1191
rect 3810 1083 3811 1089
rect 3817 1083 3842 1089
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 263 1074
rect 267 1070 407 1074
rect 411 1070 463 1074
rect 467 1070 551 1074
rect 555 1070 663 1074
rect 667 1070 695 1074
rect 699 1070 839 1074
rect 843 1070 871 1074
rect 875 1070 975 1074
rect 979 1070 1079 1074
rect 1083 1070 1119 1074
rect 1123 1070 1263 1074
rect 1267 1070 1407 1074
rect 1411 1070 1543 1074
rect 1547 1070 1679 1074
rect 1683 1070 1815 1074
rect 1819 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1069 1954 1075
rect 1958 1073 1959 1079
rect 1965 1078 3823 1079
rect 1965 1074 1975 1078
rect 1979 1074 1995 1078
rect 1999 1074 2131 1078
rect 2135 1074 2275 1078
rect 2279 1074 2443 1078
rect 2447 1074 2627 1078
rect 2631 1074 2819 1078
rect 2823 1074 2955 1078
rect 2959 1074 3027 1078
rect 3031 1074 3091 1078
rect 3095 1074 3227 1078
rect 3231 1074 3235 1078
rect 3239 1074 3451 1078
rect 3455 1074 3651 1078
rect 3655 1074 3799 1078
rect 3803 1074 3823 1078
rect 1965 1073 3823 1074
rect 3829 1073 3830 1079
rect 3836 1071 3842 1083
rect 3836 1070 5695 1071
rect 3836 1066 3839 1070
rect 3843 1066 3887 1070
rect 3891 1066 4119 1070
rect 4123 1066 4367 1070
rect 4371 1066 4607 1070
rect 4611 1066 4839 1070
rect 4843 1066 4863 1070
rect 4867 1066 4999 1070
rect 5003 1066 5071 1070
rect 5075 1066 5135 1070
rect 5139 1066 5271 1070
rect 5275 1066 5303 1070
rect 5307 1066 5407 1070
rect 5411 1066 5543 1070
rect 5547 1066 5663 1070
rect 5667 1066 5695 1070
rect 3836 1065 5695 1066
rect 5701 1065 5702 1071
rect 1946 961 1947 967
rect 1953 966 3811 967
rect 1953 962 1975 966
rect 1979 962 2023 966
rect 2027 962 2095 966
rect 2099 962 2159 966
rect 2163 962 2231 966
rect 2235 962 2303 966
rect 2307 962 2367 966
rect 2371 962 2471 966
rect 2475 962 2503 966
rect 2507 962 2655 966
rect 2659 962 2831 966
rect 2835 962 2847 966
rect 2851 962 3023 966
rect 3027 962 3055 966
rect 3059 962 3231 966
rect 3235 962 3263 966
rect 3267 962 3455 966
rect 3459 962 3479 966
rect 3483 962 3679 966
rect 3683 962 3799 966
rect 3803 962 3811 966
rect 1953 961 3811 962
rect 3817 961 3818 967
rect 96 945 97 951
rect 103 950 1959 951
rect 103 946 111 950
rect 115 946 195 950
rect 199 946 235 950
rect 239 946 371 950
rect 375 946 435 950
rect 439 946 547 950
rect 551 946 635 950
rect 639 946 723 950
rect 727 946 843 950
rect 847 946 907 950
rect 911 946 1051 950
rect 1055 946 1091 950
rect 1095 946 1935 950
rect 1939 946 1959 950
rect 103 945 1959 946
rect 1965 945 1966 951
rect 3822 941 3823 947
rect 3829 946 5707 947
rect 3829 942 3839 946
rect 3843 942 4587 946
rect 4591 942 4755 946
rect 4759 942 4835 946
rect 4839 942 4939 946
rect 4943 942 4971 946
rect 4975 942 5107 946
rect 5111 942 5131 946
rect 5135 942 5243 946
rect 5247 942 5331 946
rect 5335 942 5379 946
rect 5383 942 5515 946
rect 5519 942 5663 946
rect 5667 942 5707 946
rect 3829 941 5707 942
rect 5713 941 5714 947
rect 1958 849 1959 855
rect 1965 854 3823 855
rect 1965 850 1975 854
rect 1979 850 2067 854
rect 2071 850 2203 854
rect 2207 850 2307 854
rect 2311 850 2339 854
rect 2343 850 2475 854
rect 2479 850 2483 854
rect 2487 850 2627 854
rect 2631 850 2659 854
rect 2663 850 2803 854
rect 2807 850 2827 854
rect 2831 850 2995 854
rect 2999 850 3163 854
rect 3167 850 3203 854
rect 3207 850 3331 854
rect 3335 850 3427 854
rect 3431 850 3499 854
rect 3503 850 3651 854
rect 3655 850 3799 854
rect 3803 850 3823 854
rect 1965 849 3823 850
rect 3829 849 3830 855
rect 84 817 85 823
rect 91 822 1947 823
rect 91 818 111 822
rect 115 818 159 822
rect 163 818 223 822
rect 227 818 351 822
rect 355 818 399 822
rect 403 818 575 822
rect 579 818 583 822
rect 587 818 751 822
rect 755 818 839 822
rect 843 818 935 822
rect 939 818 1111 822
rect 1115 818 1119 822
rect 1123 818 1399 822
rect 1403 818 1687 822
rect 1691 818 1935 822
rect 1939 818 1947 822
rect 91 817 1947 818
rect 1953 817 1954 823
rect 3810 821 3811 827
rect 3817 826 5695 827
rect 3817 822 3839 826
rect 3843 822 3983 826
rect 3987 822 4239 826
rect 4243 822 4535 826
rect 4539 822 4615 826
rect 4619 822 4783 826
rect 4787 822 4863 826
rect 4867 822 4967 826
rect 4971 822 5159 826
rect 5163 822 5215 826
rect 5219 822 5359 826
rect 5363 822 5543 826
rect 5547 822 5663 826
rect 5667 822 5695 826
rect 3817 821 5695 822
rect 5701 821 5702 827
rect 1946 733 1947 739
rect 1953 738 3811 739
rect 1953 734 1975 738
rect 1979 734 2335 738
rect 2339 734 2511 738
rect 2515 734 2687 738
rect 2691 734 2855 738
rect 2859 734 3023 738
rect 3027 734 3135 738
rect 3139 734 3191 738
rect 3195 734 3271 738
rect 3275 734 3359 738
rect 3363 734 3407 738
rect 3411 734 3527 738
rect 3531 734 3543 738
rect 3547 734 3679 738
rect 3683 734 3799 738
rect 3803 734 3811 738
rect 1953 733 3811 734
rect 3817 733 3818 739
rect 96 705 97 711
rect 103 710 1959 711
rect 103 706 111 710
rect 115 706 131 710
rect 135 706 291 710
rect 295 706 323 710
rect 327 706 483 710
rect 487 706 555 710
rect 559 706 675 710
rect 679 706 811 710
rect 815 706 867 710
rect 871 706 1059 710
rect 1063 706 1083 710
rect 1087 706 1251 710
rect 1255 706 1371 710
rect 1375 706 1435 710
rect 1439 706 1619 710
rect 1623 706 1659 710
rect 1663 706 1787 710
rect 1791 706 1935 710
rect 1939 706 1959 710
rect 103 705 1959 706
rect 1965 705 1966 711
rect 3822 685 3823 691
rect 3829 690 5707 691
rect 3829 686 3839 690
rect 3843 686 3859 690
rect 3863 686 3955 690
rect 3959 686 3995 690
rect 3999 686 4139 690
rect 4143 686 4211 690
rect 4215 686 4323 690
rect 4327 686 4507 690
rect 4511 686 4531 690
rect 4535 686 4755 690
rect 4759 686 4835 690
rect 4839 686 4995 690
rect 4999 686 5187 690
rect 5191 686 5243 690
rect 5247 686 5499 690
rect 5503 686 5515 690
rect 5519 686 5663 690
rect 5667 686 5707 690
rect 3829 685 5707 686
rect 5713 685 5714 691
rect 84 593 85 599
rect 91 598 1947 599
rect 91 594 111 598
rect 115 594 159 598
rect 163 594 319 598
rect 323 594 327 598
rect 331 594 511 598
rect 515 594 519 598
rect 523 594 703 598
rect 707 594 711 598
rect 715 594 895 598
rect 899 594 903 598
rect 907 594 1087 598
rect 1091 594 1095 598
rect 1099 594 1279 598
rect 1283 594 1463 598
rect 1467 594 1647 598
rect 1651 594 1815 598
rect 1819 594 1935 598
rect 1939 594 1947 598
rect 91 593 1947 594
rect 1953 593 1954 599
rect 3810 573 3811 579
rect 3817 578 5695 579
rect 3817 574 3839 578
rect 3843 574 3887 578
rect 3891 574 4023 578
rect 4027 574 4159 578
rect 4163 574 4167 578
rect 4171 574 4295 578
rect 4299 574 4351 578
rect 4355 574 4431 578
rect 4435 574 4559 578
rect 4563 574 4575 578
rect 4579 574 4743 578
rect 4747 574 4783 578
rect 4787 574 4927 578
rect 4931 574 5023 578
rect 5027 574 5119 578
rect 5123 574 5271 578
rect 5275 574 5319 578
rect 5323 574 5527 578
rect 5531 574 5663 578
rect 5667 574 5695 578
rect 3817 573 5695 574
rect 5701 573 5702 579
rect 96 481 97 487
rect 103 486 1959 487
rect 103 482 111 486
rect 115 482 131 486
rect 135 482 299 486
rect 303 482 395 486
rect 399 482 491 486
rect 495 482 587 486
rect 591 482 683 486
rect 687 482 787 486
rect 791 482 875 486
rect 879 482 987 486
rect 991 482 1067 486
rect 1071 482 1195 486
rect 1199 482 1251 486
rect 1255 482 1411 486
rect 1415 482 1435 486
rect 1439 482 1619 486
rect 1623 482 1787 486
rect 1791 482 1935 486
rect 1939 482 1959 486
rect 103 481 1959 482
rect 1965 481 1966 487
rect 1958 461 1959 467
rect 1965 466 3823 467
rect 1965 462 1975 466
rect 1979 462 1995 466
rect 1999 462 2203 466
rect 2207 462 2427 466
rect 2431 462 2651 466
rect 2655 462 2867 466
rect 2871 462 3075 466
rect 3079 462 3107 466
rect 3111 462 3243 466
rect 3247 462 3275 466
rect 3279 462 3379 466
rect 3383 462 3475 466
rect 3479 462 3515 466
rect 3519 462 3651 466
rect 3655 462 3799 466
rect 3803 462 3823 466
rect 1965 461 3823 462
rect 3829 466 5714 467
rect 3829 462 3839 466
rect 3843 462 3859 466
rect 3863 462 3995 466
rect 3999 462 4131 466
rect 4135 462 4267 466
rect 4271 462 4379 466
rect 4383 462 4403 466
rect 4407 462 4547 466
rect 4551 462 4595 466
rect 4599 462 4715 466
rect 4719 462 4819 466
rect 4823 462 4899 466
rect 4903 462 5051 466
rect 5055 462 5091 466
rect 5095 462 5283 466
rect 5287 462 5291 466
rect 5295 462 5499 466
rect 5503 462 5663 466
rect 5667 462 5714 466
rect 3829 461 5714 462
rect 84 357 85 363
rect 91 362 1947 363
rect 91 358 111 362
rect 115 358 423 362
rect 427 358 615 362
rect 619 358 647 362
rect 651 358 815 362
rect 819 358 991 362
rect 995 358 1015 362
rect 1019 358 1167 362
rect 1171 358 1223 362
rect 1227 358 1343 362
rect 1347 358 1439 362
rect 1443 358 1935 362
rect 1939 358 1947 362
rect 91 357 1947 358
rect 1953 357 1954 363
rect 3810 349 3811 355
rect 3817 354 5695 355
rect 3817 350 3839 354
rect 3843 350 4407 354
rect 4411 350 4623 354
rect 4627 350 4639 354
rect 4643 350 4807 354
rect 4811 350 4847 354
rect 4851 350 4983 354
rect 4987 350 5079 354
rect 5083 350 5167 354
rect 5171 350 5311 354
rect 5315 350 5359 354
rect 5363 350 5543 354
rect 5547 350 5663 354
rect 5667 350 5695 354
rect 3817 349 5695 350
rect 5701 349 5702 355
rect 1946 333 1947 339
rect 1953 338 3811 339
rect 1953 334 1975 338
rect 1979 334 2023 338
rect 2027 334 2159 338
rect 2163 334 2231 338
rect 2235 334 2295 338
rect 2299 334 2431 338
rect 2435 334 2455 338
rect 2459 334 2567 338
rect 2571 334 2679 338
rect 2683 334 2703 338
rect 2707 334 2839 338
rect 2843 334 2895 338
rect 2899 334 2975 338
rect 2979 334 3103 338
rect 3107 334 3111 338
rect 3115 334 3247 338
rect 3251 334 3303 338
rect 3307 334 3383 338
rect 3387 334 3503 338
rect 3507 334 3519 338
rect 3523 334 3655 338
rect 3659 334 3679 338
rect 3683 334 3799 338
rect 3803 334 3811 338
rect 1953 333 3811 334
rect 3817 333 3818 339
rect 96 205 97 211
rect 103 210 1959 211
rect 103 206 111 210
rect 115 206 539 210
rect 543 206 619 210
rect 623 206 675 210
rect 679 206 787 210
rect 791 206 811 210
rect 815 206 947 210
rect 951 206 963 210
rect 967 206 1083 210
rect 1087 206 1139 210
rect 1143 206 1219 210
rect 1223 206 1315 210
rect 1319 206 1355 210
rect 1359 206 1491 210
rect 1495 206 1935 210
rect 1939 206 1959 210
rect 103 205 1959 206
rect 1965 205 1966 211
rect 3822 209 3823 215
rect 3829 214 5707 215
rect 3829 210 3839 214
rect 3843 210 4291 214
rect 4295 210 4427 214
rect 4431 210 4563 214
rect 4567 210 4611 214
rect 4615 210 4699 214
rect 4703 210 4779 214
rect 4783 210 4835 214
rect 4839 210 4955 214
rect 4959 210 4971 214
rect 4975 210 5107 214
rect 5111 210 5139 214
rect 5143 210 5243 214
rect 5247 210 5331 214
rect 5335 210 5379 214
rect 5383 210 5515 214
rect 5519 210 5663 214
rect 5667 210 5707 214
rect 3829 209 5707 210
rect 5713 209 5714 215
rect 1958 185 1959 191
rect 1965 190 3823 191
rect 1965 186 1975 190
rect 1979 186 1995 190
rect 1999 186 2131 190
rect 2135 186 2267 190
rect 2271 186 2403 190
rect 2407 186 2539 190
rect 2543 186 2675 190
rect 2679 186 2811 190
rect 2815 186 2947 190
rect 2951 186 3083 190
rect 3087 186 3219 190
rect 3223 186 3355 190
rect 3359 186 3491 190
rect 3495 186 3627 190
rect 3631 186 3799 190
rect 3803 186 3823 190
rect 1965 185 3823 186
rect 3829 185 3830 191
rect 84 93 85 99
rect 91 98 1947 99
rect 91 94 111 98
rect 115 94 567 98
rect 571 94 703 98
rect 707 94 839 98
rect 843 94 975 98
rect 979 94 1111 98
rect 1115 94 1247 98
rect 1251 94 1383 98
rect 1387 94 1519 98
rect 1523 94 1935 98
rect 1939 94 1947 98
rect 91 93 1947 94
rect 1953 93 1954 99
rect 3810 97 3811 103
rect 3817 102 5695 103
rect 3817 98 3839 102
rect 3843 98 4319 102
rect 4323 98 4455 102
rect 4459 98 4591 102
rect 4595 98 4727 102
rect 4731 98 4863 102
rect 4867 98 4999 102
rect 5003 98 5135 102
rect 5139 98 5271 102
rect 5275 98 5407 102
rect 5411 98 5543 102
rect 5547 98 5663 102
rect 5667 98 5695 102
rect 3817 97 5695 98
rect 5701 97 5702 103
rect 1946 73 1947 79
rect 1953 78 3811 79
rect 1953 74 1975 78
rect 1979 74 2023 78
rect 2027 74 2159 78
rect 2163 74 2295 78
rect 2299 74 2431 78
rect 2435 74 2567 78
rect 2571 74 2703 78
rect 2707 74 2839 78
rect 2843 74 2975 78
rect 2979 74 3111 78
rect 3115 74 3247 78
rect 3251 74 3383 78
rect 3387 74 3519 78
rect 3523 74 3655 78
rect 3659 74 3799 78
rect 3803 74 3811 78
rect 1953 73 3811 74
rect 3817 73 3818 79
<< m5c >>
rect 85 5717 91 5723
rect 1947 5717 1953 5723
rect 1959 5689 1965 5695
rect 3823 5689 3829 5695
rect 3823 5645 3829 5651
rect 5707 5645 5713 5651
rect 97 5601 103 5607
rect 1959 5601 1965 5607
rect 1947 5577 1953 5583
rect 3811 5577 3817 5583
rect 3811 5533 3817 5539
rect 5695 5533 5701 5539
rect 85 5477 91 5483
rect 1947 5477 1953 5483
rect 1959 5457 1965 5463
rect 3823 5457 3829 5463
rect 3823 5417 3829 5423
rect 5707 5417 5713 5423
rect 1947 5345 1953 5351
rect 3811 5345 3817 5351
rect 3811 5289 3817 5295
rect 5695 5289 5701 5295
rect 97 5261 103 5267
rect 1959 5261 1965 5267
rect 1959 5233 1965 5239
rect 3823 5233 3829 5239
rect 3823 5169 3829 5175
rect 5707 5169 5713 5175
rect 85 5133 91 5139
rect 1947 5133 1953 5139
rect 1947 5097 1953 5103
rect 3811 5097 3817 5103
rect 3811 5041 3817 5047
rect 5695 5041 5701 5047
rect 97 5021 103 5027
rect 1959 5021 1965 5027
rect 1959 4965 1965 4971
rect 3823 4965 3829 4971
rect 85 4909 91 4915
rect 1947 4909 1953 4915
rect 3823 4913 3829 4919
rect 5707 4913 5713 4919
rect 1947 4825 1953 4831
rect 3811 4825 3817 4831
rect 97 4785 103 4791
rect 1959 4785 1965 4791
rect 3811 4781 3817 4787
rect 5695 4781 5701 4787
rect 1959 4705 1965 4711
rect 3823 4705 3829 4711
rect 85 4669 91 4675
rect 1947 4669 1953 4675
rect 3823 4649 3829 4655
rect 5707 4649 5713 4655
rect 1947 4593 1953 4599
rect 3811 4593 3817 4599
rect 97 4545 103 4551
rect 1959 4545 1965 4551
rect 3811 4513 3817 4519
rect 5695 4513 5701 4519
rect 1959 4441 1965 4447
rect 3823 4441 3829 4447
rect 85 4433 91 4439
rect 1947 4433 1953 4439
rect 3823 4401 3829 4407
rect 5707 4401 5713 4407
rect 1947 4325 1953 4331
rect 3811 4325 3817 4331
rect 97 4313 103 4319
rect 1959 4313 1965 4319
rect 3811 4289 3817 4295
rect 5695 4289 5701 4295
rect 1959 4201 1965 4207
rect 3823 4201 3829 4207
rect 85 4189 91 4195
rect 1947 4189 1953 4195
rect 3823 4093 3829 4099
rect 5707 4093 5713 4099
rect 1947 4085 1953 4091
rect 3811 4085 3817 4091
rect 97 4065 103 4071
rect 1959 4065 1965 4071
rect 3811 3983 3817 3989
rect 1959 3973 1965 3979
rect 3823 3973 3829 3979
rect 5695 3973 5701 3979
rect 85 3941 91 3947
rect 1947 3941 1953 3947
rect 1947 3857 1953 3863
rect 3811 3857 3817 3863
rect 3823 3829 3829 3835
rect 5707 3829 5713 3835
rect 97 3821 103 3827
rect 1959 3821 1965 3827
rect 1959 3737 1965 3743
rect 3823 3737 3829 3743
rect 85 3697 91 3703
rect 1947 3697 1953 3703
rect 3811 3697 3817 3703
rect 5695 3697 5701 3703
rect 1947 3621 1953 3627
rect 3811 3621 3817 3627
rect 97 3565 103 3571
rect 1959 3565 1965 3571
rect 3823 3557 3829 3563
rect 5707 3557 5713 3563
rect 1959 3485 1965 3491
rect 3823 3485 3829 3491
rect 85 3433 91 3439
rect 1947 3433 1953 3439
rect 3811 3433 3817 3439
rect 5695 3433 5701 3439
rect 1947 3361 1953 3367
rect 3811 3361 3817 3367
rect 3823 3321 3829 3327
rect 5707 3321 5713 3327
rect 97 3305 103 3311
rect 1959 3305 1965 3311
rect 1959 3245 1965 3251
rect 3823 3245 3829 3251
rect 3811 3201 3817 3207
rect 5695 3201 5701 3207
rect 85 3177 91 3183
rect 1947 3177 1953 3183
rect 1947 3133 1953 3139
rect 3811 3133 3817 3139
rect 3823 3085 3829 3091
rect 5707 3085 5713 3091
rect 97 3065 103 3071
rect 1959 3065 1965 3071
rect 1959 3013 1965 3019
rect 3823 3013 3829 3019
rect 3811 2969 3817 2975
rect 5695 2969 5701 2975
rect 85 2953 91 2959
rect 1947 2953 1953 2959
rect 3823 2857 3829 2863
rect 5707 2857 5713 2863
rect 97 2829 103 2835
rect 1959 2829 1965 2835
rect 3811 2729 3817 2735
rect 5695 2729 5701 2735
rect 85 2713 91 2719
rect 1947 2713 1953 2719
rect 1947 2633 1953 2639
rect 3811 2633 3817 2639
rect 97 2597 103 2603
rect 1959 2597 1965 2603
rect 3823 2601 3829 2607
rect 5707 2601 5713 2607
rect 1959 2521 1965 2527
rect 3823 2521 3829 2527
rect 3811 2489 3817 2495
rect 5695 2489 5701 2495
rect 85 2477 91 2483
rect 1947 2477 1953 2483
rect 1947 2409 1953 2415
rect 3811 2409 3817 2415
rect 3823 2377 3829 2383
rect 5707 2377 5713 2383
rect 97 2353 103 2359
rect 1959 2353 1965 2359
rect 1959 2289 1965 2295
rect 3823 2289 3829 2295
rect 3811 2253 3817 2259
rect 5695 2253 5701 2259
rect 85 2241 91 2247
rect 1947 2241 1953 2247
rect 1947 2173 1953 2179
rect 3811 2173 3817 2179
rect 97 2129 103 2135
rect 1959 2129 1965 2135
rect 3823 2133 3829 2139
rect 5707 2133 5713 2139
rect 1959 2053 1965 2059
rect 3823 2053 3829 2059
rect 85 2013 91 2019
rect 1947 2013 1953 2019
rect 3811 2017 3817 2023
rect 5695 2017 5701 2023
rect 1947 1933 1953 1939
rect 3811 1933 3817 1939
rect 97 1901 103 1907
rect 1959 1901 1965 1907
rect 3823 1901 3829 1907
rect 5707 1901 5713 1907
rect 1959 1821 1965 1827
rect 3823 1821 3829 1827
rect 85 1785 91 1791
rect 1947 1785 1953 1791
rect 3811 1785 3817 1791
rect 5695 1785 5701 1791
rect 1947 1683 1953 1689
rect 97 1673 103 1679
rect 1959 1673 1965 1679
rect 3823 1673 3829 1679
rect 5707 1673 5713 1679
rect 3811 1665 3817 1671
rect 85 1561 91 1567
rect 1947 1561 1953 1567
rect 3811 1561 3817 1567
rect 5695 1561 5701 1567
rect 1959 1541 1965 1547
rect 3823 1541 3829 1547
rect 1947 1439 1953 1445
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3811 1429 3817 1435
rect 3823 1433 3829 1439
rect 5707 1433 5713 1439
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 3811 1317 3817 1323
rect 5695 1317 5701 1323
rect 1959 1297 1965 1303
rect 3823 1297 3829 1303
rect 1947 1203 1953 1209
rect 97 1193 103 1199
rect 1959 1193 1965 1199
rect 3823 1197 3829 1203
rect 5707 1197 5713 1203
rect 3811 1185 3817 1191
rect 3811 1083 3817 1089
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 1959 1073 1965 1079
rect 3823 1073 3829 1079
rect 5695 1065 5701 1071
rect 1947 961 1953 967
rect 3811 961 3817 967
rect 97 945 103 951
rect 1959 945 1965 951
rect 3823 941 3829 947
rect 5707 941 5713 947
rect 1959 849 1965 855
rect 3823 849 3829 855
rect 85 817 91 823
rect 1947 817 1953 823
rect 3811 821 3817 827
rect 5695 821 5701 827
rect 1947 733 1953 739
rect 3811 733 3817 739
rect 97 705 103 711
rect 1959 705 1965 711
rect 3823 685 3829 691
rect 5707 685 5713 691
rect 85 593 91 599
rect 1947 593 1953 599
rect 3811 573 3817 579
rect 5695 573 5701 579
rect 97 481 103 487
rect 1959 481 1965 487
rect 1959 461 1965 467
rect 3823 461 3829 467
rect 85 357 91 363
rect 1947 357 1953 363
rect 3811 349 3817 355
rect 5695 349 5701 355
rect 1947 333 1953 339
rect 3811 333 3817 339
rect 97 205 103 211
rect 1959 205 1965 211
rect 3823 209 3829 215
rect 5707 209 5713 215
rect 1959 185 1965 191
rect 3823 185 3829 191
rect 85 93 91 99
rect 1947 93 1953 99
rect 3811 97 3817 103
rect 5695 97 5701 103
rect 1947 73 1953 79
rect 3811 73 3817 79
<< m5 >>
rect 84 5723 92 5760
rect 84 5717 85 5723
rect 91 5717 92 5723
rect 84 5483 92 5717
rect 84 5477 85 5483
rect 91 5477 92 5483
rect 84 5139 92 5477
rect 84 5133 85 5139
rect 91 5133 92 5139
rect 84 4915 92 5133
rect 84 4909 85 4915
rect 91 4909 92 4915
rect 84 4675 92 4909
rect 84 4669 85 4675
rect 91 4669 92 4675
rect 84 4439 92 4669
rect 84 4433 85 4439
rect 91 4433 92 4439
rect 84 4195 92 4433
rect 84 4189 85 4195
rect 91 4189 92 4195
rect 84 3947 92 4189
rect 84 3941 85 3947
rect 91 3941 92 3947
rect 84 3703 92 3941
rect 84 3697 85 3703
rect 91 3697 92 3703
rect 84 3439 92 3697
rect 84 3433 85 3439
rect 91 3433 92 3439
rect 84 3183 92 3433
rect 84 3177 85 3183
rect 91 3177 92 3183
rect 84 2959 92 3177
rect 84 2953 85 2959
rect 91 2953 92 2959
rect 84 2719 92 2953
rect 84 2713 85 2719
rect 91 2713 92 2719
rect 84 2483 92 2713
rect 84 2477 85 2483
rect 91 2477 92 2483
rect 84 2247 92 2477
rect 84 2241 85 2247
rect 91 2241 92 2247
rect 84 2019 92 2241
rect 84 2013 85 2019
rect 91 2013 92 2019
rect 84 1791 92 2013
rect 84 1785 85 1791
rect 91 1785 92 1791
rect 84 1567 92 1785
rect 84 1561 85 1567
rect 91 1561 92 1567
rect 84 1323 92 1561
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 823 92 1069
rect 84 817 85 823
rect 91 817 92 823
rect 84 599 92 817
rect 84 593 85 599
rect 91 593 92 599
rect 84 363 92 593
rect 84 357 85 363
rect 91 357 92 363
rect 84 99 92 357
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 5607 104 5760
rect 96 5601 97 5607
rect 103 5601 104 5607
rect 96 5267 104 5601
rect 96 5261 97 5267
rect 103 5261 104 5267
rect 96 5027 104 5261
rect 96 5021 97 5027
rect 103 5021 104 5027
rect 96 4791 104 5021
rect 96 4785 97 4791
rect 103 4785 104 4791
rect 96 4551 104 4785
rect 96 4545 97 4551
rect 103 4545 104 4551
rect 96 4319 104 4545
rect 96 4313 97 4319
rect 103 4313 104 4319
rect 96 4071 104 4313
rect 96 4065 97 4071
rect 103 4065 104 4071
rect 96 3827 104 4065
rect 96 3821 97 3827
rect 103 3821 104 3827
rect 96 3571 104 3821
rect 96 3565 97 3571
rect 103 3565 104 3571
rect 96 3311 104 3565
rect 96 3305 97 3311
rect 103 3305 104 3311
rect 96 3071 104 3305
rect 96 3065 97 3071
rect 103 3065 104 3071
rect 96 2835 104 3065
rect 96 2829 97 2835
rect 103 2829 104 2835
rect 96 2603 104 2829
rect 96 2597 97 2603
rect 103 2597 104 2603
rect 96 2359 104 2597
rect 96 2353 97 2359
rect 103 2353 104 2359
rect 96 2135 104 2353
rect 96 2129 97 2135
rect 103 2129 104 2135
rect 96 1907 104 2129
rect 96 1901 97 1907
rect 103 1901 104 1907
rect 96 1679 104 1901
rect 96 1673 97 1679
rect 103 1673 104 1679
rect 96 1435 104 1673
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1199 104 1429
rect 96 1193 97 1199
rect 103 1193 104 1199
rect 96 951 104 1193
rect 96 945 97 951
rect 103 945 104 951
rect 96 711 104 945
rect 96 705 97 711
rect 103 705 104 711
rect 96 487 104 705
rect 96 481 97 487
rect 103 481 104 487
rect 96 211 104 481
rect 96 205 97 211
rect 103 205 104 211
rect 96 72 104 205
rect 1946 5723 1954 5760
rect 1946 5717 1947 5723
rect 1953 5717 1954 5723
rect 1946 5583 1954 5717
rect 1946 5577 1947 5583
rect 1953 5577 1954 5583
rect 1946 5483 1954 5577
rect 1946 5477 1947 5483
rect 1953 5477 1954 5483
rect 1946 5351 1954 5477
rect 1946 5345 1947 5351
rect 1953 5345 1954 5351
rect 1946 5139 1954 5345
rect 1946 5133 1947 5139
rect 1953 5133 1954 5139
rect 1946 5103 1954 5133
rect 1946 5097 1947 5103
rect 1953 5097 1954 5103
rect 1946 4915 1954 5097
rect 1946 4909 1947 4915
rect 1953 4909 1954 4915
rect 1946 4831 1954 4909
rect 1946 4825 1947 4831
rect 1953 4825 1954 4831
rect 1946 4675 1954 4825
rect 1946 4669 1947 4675
rect 1953 4669 1954 4675
rect 1946 4599 1954 4669
rect 1946 4593 1947 4599
rect 1953 4593 1954 4599
rect 1946 4439 1954 4593
rect 1946 4433 1947 4439
rect 1953 4433 1954 4439
rect 1946 4331 1954 4433
rect 1946 4325 1947 4331
rect 1953 4325 1954 4331
rect 1946 4195 1954 4325
rect 1946 4189 1947 4195
rect 1953 4189 1954 4195
rect 1946 4091 1954 4189
rect 1946 4085 1947 4091
rect 1953 4085 1954 4091
rect 1946 3947 1954 4085
rect 1946 3941 1947 3947
rect 1953 3941 1954 3947
rect 1946 3863 1954 3941
rect 1946 3857 1947 3863
rect 1953 3857 1954 3863
rect 1946 3703 1954 3857
rect 1946 3697 1947 3703
rect 1953 3697 1954 3703
rect 1946 3627 1954 3697
rect 1946 3621 1947 3627
rect 1953 3621 1954 3627
rect 1946 3439 1954 3621
rect 1946 3433 1947 3439
rect 1953 3433 1954 3439
rect 1946 3367 1954 3433
rect 1946 3361 1947 3367
rect 1953 3361 1954 3367
rect 1946 3183 1954 3361
rect 1946 3177 1947 3183
rect 1953 3177 1954 3183
rect 1946 3139 1954 3177
rect 1946 3133 1947 3139
rect 1953 3133 1954 3139
rect 1946 2959 1954 3133
rect 1946 2953 1947 2959
rect 1953 2953 1954 2959
rect 1946 2719 1954 2953
rect 1946 2713 1947 2719
rect 1953 2713 1954 2719
rect 1946 2639 1954 2713
rect 1946 2633 1947 2639
rect 1953 2633 1954 2639
rect 1946 2483 1954 2633
rect 1946 2477 1947 2483
rect 1953 2477 1954 2483
rect 1946 2415 1954 2477
rect 1946 2409 1947 2415
rect 1953 2409 1954 2415
rect 1946 2247 1954 2409
rect 1946 2241 1947 2247
rect 1953 2241 1954 2247
rect 1946 2179 1954 2241
rect 1946 2173 1947 2179
rect 1953 2173 1954 2179
rect 1946 2019 1954 2173
rect 1946 2013 1947 2019
rect 1953 2013 1954 2019
rect 1946 1939 1954 2013
rect 1946 1933 1947 1939
rect 1953 1933 1954 1939
rect 1946 1791 1954 1933
rect 1946 1785 1947 1791
rect 1953 1785 1954 1791
rect 1946 1689 1954 1785
rect 1946 1683 1947 1689
rect 1953 1683 1954 1689
rect 1946 1567 1954 1683
rect 1946 1561 1947 1567
rect 1953 1561 1954 1567
rect 1946 1445 1954 1561
rect 1946 1439 1947 1445
rect 1953 1439 1954 1445
rect 1946 1323 1954 1439
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1209 1954 1317
rect 1946 1203 1947 1209
rect 1953 1203 1954 1209
rect 1946 1075 1954 1203
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 967 1954 1069
rect 1946 961 1947 967
rect 1953 961 1954 967
rect 1946 823 1954 961
rect 1946 817 1947 823
rect 1953 817 1954 823
rect 1946 739 1954 817
rect 1946 733 1947 739
rect 1953 733 1954 739
rect 1946 599 1954 733
rect 1946 593 1947 599
rect 1953 593 1954 599
rect 1946 363 1954 593
rect 1946 357 1947 363
rect 1953 357 1954 363
rect 1946 339 1954 357
rect 1946 333 1947 339
rect 1953 333 1954 339
rect 1946 99 1954 333
rect 1946 93 1947 99
rect 1953 93 1954 99
rect 1946 79 1954 93
rect 1946 73 1947 79
rect 1953 73 1954 79
rect 1946 72 1954 73
rect 1958 5695 1966 5760
rect 1958 5689 1959 5695
rect 1965 5689 1966 5695
rect 1958 5607 1966 5689
rect 1958 5601 1959 5607
rect 1965 5601 1966 5607
rect 1958 5463 1966 5601
rect 1958 5457 1959 5463
rect 1965 5457 1966 5463
rect 1958 5267 1966 5457
rect 1958 5261 1959 5267
rect 1965 5261 1966 5267
rect 1958 5239 1966 5261
rect 1958 5233 1959 5239
rect 1965 5233 1966 5239
rect 1958 5027 1966 5233
rect 1958 5021 1959 5027
rect 1965 5021 1966 5027
rect 1958 4971 1966 5021
rect 1958 4965 1959 4971
rect 1965 4965 1966 4971
rect 1958 4791 1966 4965
rect 1958 4785 1959 4791
rect 1965 4785 1966 4791
rect 1958 4711 1966 4785
rect 1958 4705 1959 4711
rect 1965 4705 1966 4711
rect 1958 4551 1966 4705
rect 1958 4545 1959 4551
rect 1965 4545 1966 4551
rect 1958 4447 1966 4545
rect 1958 4441 1959 4447
rect 1965 4441 1966 4447
rect 1958 4319 1966 4441
rect 1958 4313 1959 4319
rect 1965 4313 1966 4319
rect 1958 4207 1966 4313
rect 1958 4201 1959 4207
rect 1965 4201 1966 4207
rect 1958 4071 1966 4201
rect 1958 4065 1959 4071
rect 1965 4065 1966 4071
rect 1958 3979 1966 4065
rect 1958 3973 1959 3979
rect 1965 3973 1966 3979
rect 1958 3827 1966 3973
rect 1958 3821 1959 3827
rect 1965 3821 1966 3827
rect 1958 3743 1966 3821
rect 1958 3737 1959 3743
rect 1965 3737 1966 3743
rect 1958 3571 1966 3737
rect 1958 3565 1959 3571
rect 1965 3565 1966 3571
rect 1958 3491 1966 3565
rect 1958 3485 1959 3491
rect 1965 3485 1966 3491
rect 1958 3311 1966 3485
rect 1958 3305 1959 3311
rect 1965 3305 1966 3311
rect 1958 3251 1966 3305
rect 1958 3245 1959 3251
rect 1965 3245 1966 3251
rect 1958 3071 1966 3245
rect 1958 3065 1959 3071
rect 1965 3065 1966 3071
rect 1958 3019 1966 3065
rect 1958 3013 1959 3019
rect 1965 3013 1966 3019
rect 1958 2835 1966 3013
rect 1958 2829 1959 2835
rect 1965 2829 1966 2835
rect 1958 2603 1966 2829
rect 1958 2597 1959 2603
rect 1965 2597 1966 2603
rect 1958 2527 1966 2597
rect 1958 2521 1959 2527
rect 1965 2521 1966 2527
rect 1958 2359 1966 2521
rect 1958 2353 1959 2359
rect 1965 2353 1966 2359
rect 1958 2295 1966 2353
rect 1958 2289 1959 2295
rect 1965 2289 1966 2295
rect 1958 2135 1966 2289
rect 1958 2129 1959 2135
rect 1965 2129 1966 2135
rect 1958 2059 1966 2129
rect 1958 2053 1959 2059
rect 1965 2053 1966 2059
rect 1958 1907 1966 2053
rect 1958 1901 1959 1907
rect 1965 1901 1966 1907
rect 1958 1827 1966 1901
rect 1958 1821 1959 1827
rect 1965 1821 1966 1827
rect 1958 1679 1966 1821
rect 1958 1673 1959 1679
rect 1965 1673 1966 1679
rect 1958 1547 1966 1673
rect 1958 1541 1959 1547
rect 1965 1541 1966 1547
rect 1958 1435 1966 1541
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1303 1966 1429
rect 1958 1297 1959 1303
rect 1965 1297 1966 1303
rect 1958 1199 1966 1297
rect 1958 1193 1959 1199
rect 1965 1193 1966 1199
rect 1958 1079 1966 1193
rect 1958 1073 1959 1079
rect 1965 1073 1966 1079
rect 1958 951 1966 1073
rect 1958 945 1959 951
rect 1965 945 1966 951
rect 1958 855 1966 945
rect 1958 849 1959 855
rect 1965 849 1966 855
rect 1958 711 1966 849
rect 1958 705 1959 711
rect 1965 705 1966 711
rect 1958 487 1966 705
rect 1958 481 1959 487
rect 1965 481 1966 487
rect 1958 467 1966 481
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 211 1966 461
rect 1958 205 1959 211
rect 1965 205 1966 211
rect 1958 191 1966 205
rect 1958 185 1959 191
rect 1965 185 1966 191
rect 1958 72 1966 185
rect 3810 5583 3818 5760
rect 3810 5577 3811 5583
rect 3817 5577 3818 5583
rect 3810 5539 3818 5577
rect 3810 5533 3811 5539
rect 3817 5533 3818 5539
rect 3810 5351 3818 5533
rect 3810 5345 3811 5351
rect 3817 5345 3818 5351
rect 3810 5295 3818 5345
rect 3810 5289 3811 5295
rect 3817 5289 3818 5295
rect 3810 5103 3818 5289
rect 3810 5097 3811 5103
rect 3817 5097 3818 5103
rect 3810 5047 3818 5097
rect 3810 5041 3811 5047
rect 3817 5041 3818 5047
rect 3810 4831 3818 5041
rect 3810 4825 3811 4831
rect 3817 4825 3818 4831
rect 3810 4787 3818 4825
rect 3810 4781 3811 4787
rect 3817 4781 3818 4787
rect 3810 4599 3818 4781
rect 3810 4593 3811 4599
rect 3817 4593 3818 4599
rect 3810 4519 3818 4593
rect 3810 4513 3811 4519
rect 3817 4513 3818 4519
rect 3810 4331 3818 4513
rect 3810 4325 3811 4331
rect 3817 4325 3818 4331
rect 3810 4295 3818 4325
rect 3810 4289 3811 4295
rect 3817 4289 3818 4295
rect 3810 4091 3818 4289
rect 3810 4085 3811 4091
rect 3817 4085 3818 4091
rect 3810 3989 3818 4085
rect 3810 3983 3811 3989
rect 3817 3983 3818 3989
rect 3810 3863 3818 3983
rect 3810 3857 3811 3863
rect 3817 3857 3818 3863
rect 3810 3703 3818 3857
rect 3810 3697 3811 3703
rect 3817 3697 3818 3703
rect 3810 3627 3818 3697
rect 3810 3621 3811 3627
rect 3817 3621 3818 3627
rect 3810 3439 3818 3621
rect 3810 3433 3811 3439
rect 3817 3433 3818 3439
rect 3810 3367 3818 3433
rect 3810 3361 3811 3367
rect 3817 3361 3818 3367
rect 3810 3207 3818 3361
rect 3810 3201 3811 3207
rect 3817 3201 3818 3207
rect 3810 3139 3818 3201
rect 3810 3133 3811 3139
rect 3817 3133 3818 3139
rect 3810 2975 3818 3133
rect 3810 2969 3811 2975
rect 3817 2969 3818 2975
rect 3810 2735 3818 2969
rect 3810 2729 3811 2735
rect 3817 2729 3818 2735
rect 3810 2639 3818 2729
rect 3810 2633 3811 2639
rect 3817 2633 3818 2639
rect 3810 2495 3818 2633
rect 3810 2489 3811 2495
rect 3817 2489 3818 2495
rect 3810 2415 3818 2489
rect 3810 2409 3811 2415
rect 3817 2409 3818 2415
rect 3810 2259 3818 2409
rect 3810 2253 3811 2259
rect 3817 2253 3818 2259
rect 3810 2179 3818 2253
rect 3810 2173 3811 2179
rect 3817 2173 3818 2179
rect 3810 2023 3818 2173
rect 3810 2017 3811 2023
rect 3817 2017 3818 2023
rect 3810 1939 3818 2017
rect 3810 1933 3811 1939
rect 3817 1933 3818 1939
rect 3810 1791 3818 1933
rect 3810 1785 3811 1791
rect 3817 1785 3818 1791
rect 3810 1671 3818 1785
rect 3810 1665 3811 1671
rect 3817 1665 3818 1671
rect 3810 1567 3818 1665
rect 3810 1561 3811 1567
rect 3817 1561 3818 1567
rect 3810 1435 3818 1561
rect 3810 1429 3811 1435
rect 3817 1429 3818 1435
rect 3810 1323 3818 1429
rect 3810 1317 3811 1323
rect 3817 1317 3818 1323
rect 3810 1191 3818 1317
rect 3810 1185 3811 1191
rect 3817 1185 3818 1191
rect 3810 1089 3818 1185
rect 3810 1083 3811 1089
rect 3817 1083 3818 1089
rect 3810 967 3818 1083
rect 3810 961 3811 967
rect 3817 961 3818 967
rect 3810 827 3818 961
rect 3810 821 3811 827
rect 3817 821 3818 827
rect 3810 739 3818 821
rect 3810 733 3811 739
rect 3817 733 3818 739
rect 3810 579 3818 733
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 355 3818 573
rect 3810 349 3811 355
rect 3817 349 3818 355
rect 3810 339 3818 349
rect 3810 333 3811 339
rect 3817 333 3818 339
rect 3810 103 3818 333
rect 3810 97 3811 103
rect 3817 97 3818 103
rect 3810 79 3818 97
rect 3810 73 3811 79
rect 3817 73 3818 79
rect 3810 72 3818 73
rect 3822 5695 3830 5760
rect 3822 5689 3823 5695
rect 3829 5689 3830 5695
rect 3822 5651 3830 5689
rect 3822 5645 3823 5651
rect 3829 5645 3830 5651
rect 3822 5463 3830 5645
rect 3822 5457 3823 5463
rect 3829 5457 3830 5463
rect 3822 5423 3830 5457
rect 3822 5417 3823 5423
rect 3829 5417 3830 5423
rect 3822 5239 3830 5417
rect 3822 5233 3823 5239
rect 3829 5233 3830 5239
rect 3822 5175 3830 5233
rect 3822 5169 3823 5175
rect 3829 5169 3830 5175
rect 3822 4971 3830 5169
rect 3822 4965 3823 4971
rect 3829 4965 3830 4971
rect 3822 4919 3830 4965
rect 3822 4913 3823 4919
rect 3829 4913 3830 4919
rect 3822 4711 3830 4913
rect 3822 4705 3823 4711
rect 3829 4705 3830 4711
rect 3822 4655 3830 4705
rect 3822 4649 3823 4655
rect 3829 4649 3830 4655
rect 3822 4447 3830 4649
rect 3822 4441 3823 4447
rect 3829 4441 3830 4447
rect 3822 4407 3830 4441
rect 3822 4401 3823 4407
rect 3829 4401 3830 4407
rect 3822 4207 3830 4401
rect 3822 4201 3823 4207
rect 3829 4201 3830 4207
rect 3822 4099 3830 4201
rect 3822 4093 3823 4099
rect 3829 4093 3830 4099
rect 3822 3979 3830 4093
rect 3822 3973 3823 3979
rect 3829 3973 3830 3979
rect 3822 3835 3830 3973
rect 3822 3829 3823 3835
rect 3829 3829 3830 3835
rect 3822 3743 3830 3829
rect 3822 3737 3823 3743
rect 3829 3737 3830 3743
rect 3822 3563 3830 3737
rect 3822 3557 3823 3563
rect 3829 3557 3830 3563
rect 3822 3491 3830 3557
rect 3822 3485 3823 3491
rect 3829 3485 3830 3491
rect 3822 3327 3830 3485
rect 3822 3321 3823 3327
rect 3829 3321 3830 3327
rect 3822 3251 3830 3321
rect 3822 3245 3823 3251
rect 3829 3245 3830 3251
rect 3822 3091 3830 3245
rect 3822 3085 3823 3091
rect 3829 3085 3830 3091
rect 3822 3019 3830 3085
rect 3822 3013 3823 3019
rect 3829 3013 3830 3019
rect 3822 2863 3830 3013
rect 3822 2857 3823 2863
rect 3829 2857 3830 2863
rect 3822 2607 3830 2857
rect 3822 2601 3823 2607
rect 3829 2601 3830 2607
rect 3822 2527 3830 2601
rect 3822 2521 3823 2527
rect 3829 2521 3830 2527
rect 3822 2383 3830 2521
rect 3822 2377 3823 2383
rect 3829 2377 3830 2383
rect 3822 2295 3830 2377
rect 3822 2289 3823 2295
rect 3829 2289 3830 2295
rect 3822 2139 3830 2289
rect 3822 2133 3823 2139
rect 3829 2133 3830 2139
rect 3822 2059 3830 2133
rect 3822 2053 3823 2059
rect 3829 2053 3830 2059
rect 3822 1907 3830 2053
rect 3822 1901 3823 1907
rect 3829 1901 3830 1907
rect 3822 1827 3830 1901
rect 3822 1821 3823 1827
rect 3829 1821 3830 1827
rect 3822 1679 3830 1821
rect 3822 1673 3823 1679
rect 3829 1673 3830 1679
rect 3822 1547 3830 1673
rect 3822 1541 3823 1547
rect 3829 1541 3830 1547
rect 3822 1439 3830 1541
rect 3822 1433 3823 1439
rect 3829 1433 3830 1439
rect 3822 1303 3830 1433
rect 3822 1297 3823 1303
rect 3829 1297 3830 1303
rect 3822 1203 3830 1297
rect 3822 1197 3823 1203
rect 3829 1197 3830 1203
rect 3822 1079 3830 1197
rect 3822 1073 3823 1079
rect 3829 1073 3830 1079
rect 3822 947 3830 1073
rect 3822 941 3823 947
rect 3829 941 3830 947
rect 3822 855 3830 941
rect 3822 849 3823 855
rect 3829 849 3830 855
rect 3822 691 3830 849
rect 3822 685 3823 691
rect 3829 685 3830 691
rect 3822 467 3830 685
rect 3822 461 3823 467
rect 3829 461 3830 467
rect 3822 215 3830 461
rect 3822 209 3823 215
rect 3829 209 3830 215
rect 3822 191 3830 209
rect 3822 185 3823 191
rect 3829 185 3830 191
rect 3822 72 3830 185
rect 5694 5539 5702 5760
rect 5694 5533 5695 5539
rect 5701 5533 5702 5539
rect 5694 5295 5702 5533
rect 5694 5289 5695 5295
rect 5701 5289 5702 5295
rect 5694 5047 5702 5289
rect 5694 5041 5695 5047
rect 5701 5041 5702 5047
rect 5694 4787 5702 5041
rect 5694 4781 5695 4787
rect 5701 4781 5702 4787
rect 5694 4519 5702 4781
rect 5694 4513 5695 4519
rect 5701 4513 5702 4519
rect 5694 4295 5702 4513
rect 5694 4289 5695 4295
rect 5701 4289 5702 4295
rect 5694 3979 5702 4289
rect 5694 3973 5695 3979
rect 5701 3973 5702 3979
rect 5694 3703 5702 3973
rect 5694 3697 5695 3703
rect 5701 3697 5702 3703
rect 5694 3439 5702 3697
rect 5694 3433 5695 3439
rect 5701 3433 5702 3439
rect 5694 3207 5702 3433
rect 5694 3201 5695 3207
rect 5701 3201 5702 3207
rect 5694 2975 5702 3201
rect 5694 2969 5695 2975
rect 5701 2969 5702 2975
rect 5694 2735 5702 2969
rect 5694 2729 5695 2735
rect 5701 2729 5702 2735
rect 5694 2495 5702 2729
rect 5694 2489 5695 2495
rect 5701 2489 5702 2495
rect 5694 2259 5702 2489
rect 5694 2253 5695 2259
rect 5701 2253 5702 2259
rect 5694 2023 5702 2253
rect 5694 2017 5695 2023
rect 5701 2017 5702 2023
rect 5694 1791 5702 2017
rect 5694 1785 5695 1791
rect 5701 1785 5702 1791
rect 5694 1567 5702 1785
rect 5694 1561 5695 1567
rect 5701 1561 5702 1567
rect 5694 1323 5702 1561
rect 5694 1317 5695 1323
rect 5701 1317 5702 1323
rect 5694 1071 5702 1317
rect 5694 1065 5695 1071
rect 5701 1065 5702 1071
rect 5694 827 5702 1065
rect 5694 821 5695 827
rect 5701 821 5702 827
rect 5694 579 5702 821
rect 5694 573 5695 579
rect 5701 573 5702 579
rect 5694 355 5702 573
rect 5694 349 5695 355
rect 5701 349 5702 355
rect 5694 103 5702 349
rect 5694 97 5695 103
rect 5701 97 5702 103
rect 5694 72 5702 97
rect 5706 5651 5714 5760
rect 5706 5645 5707 5651
rect 5713 5645 5714 5651
rect 5706 5423 5714 5645
rect 5706 5417 5707 5423
rect 5713 5417 5714 5423
rect 5706 5175 5714 5417
rect 5706 5169 5707 5175
rect 5713 5169 5714 5175
rect 5706 4919 5714 5169
rect 5706 4913 5707 4919
rect 5713 4913 5714 4919
rect 5706 4655 5714 4913
rect 5706 4649 5707 4655
rect 5713 4649 5714 4655
rect 5706 4407 5714 4649
rect 5706 4401 5707 4407
rect 5713 4401 5714 4407
rect 5706 4099 5714 4401
rect 5706 4093 5707 4099
rect 5713 4093 5714 4099
rect 5706 3835 5714 4093
rect 5706 3829 5707 3835
rect 5713 3829 5714 3835
rect 5706 3563 5714 3829
rect 5706 3557 5707 3563
rect 5713 3557 5714 3563
rect 5706 3327 5714 3557
rect 5706 3321 5707 3327
rect 5713 3321 5714 3327
rect 5706 3091 5714 3321
rect 5706 3085 5707 3091
rect 5713 3085 5714 3091
rect 5706 2863 5714 3085
rect 5706 2857 5707 2863
rect 5713 2857 5714 2863
rect 5706 2607 5714 2857
rect 5706 2601 5707 2607
rect 5713 2601 5714 2607
rect 5706 2383 5714 2601
rect 5706 2377 5707 2383
rect 5713 2377 5714 2383
rect 5706 2139 5714 2377
rect 5706 2133 5707 2139
rect 5713 2133 5714 2139
rect 5706 1907 5714 2133
rect 5706 1901 5707 1907
rect 5713 1901 5714 1907
rect 5706 1679 5714 1901
rect 5706 1673 5707 1679
rect 5713 1673 5714 1679
rect 5706 1439 5714 1673
rect 5706 1433 5707 1439
rect 5713 1433 5714 1439
rect 5706 1203 5714 1433
rect 5706 1197 5707 1203
rect 5713 1197 5714 1203
rect 5706 947 5714 1197
rect 5706 941 5707 947
rect 5713 941 5714 947
rect 5706 691 5714 941
rect 5706 685 5707 691
rect 5713 685 5714 691
rect 5706 215 5714 685
rect 5706 209 5707 215
rect 5713 209 5714 215
rect 5706 72 5714 209
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__267
timestamp 1731220429
transform 1 0 5656 0 1 5560
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220429
transform 1 0 3832 0 1 5560
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220429
transform 1 0 5656 0 -1 5512
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220429
transform 1 0 3832 0 -1 5512
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220429
transform 1 0 5656 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220429
transform 1 0 3832 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220429
transform 1 0 5656 0 -1 5268
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220429
transform 1 0 3832 0 -1 5268
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220429
transform 1 0 5656 0 1 5084
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220429
transform 1 0 3832 0 1 5084
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220429
transform 1 0 5656 0 -1 5020
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220429
transform 1 0 3832 0 -1 5020
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220429
transform 1 0 5656 0 1 4828
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220429
transform 1 0 3832 0 1 4828
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220429
transform 1 0 5656 0 -1 4760
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220429
transform 1 0 3832 0 -1 4760
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220429
transform 1 0 5656 0 1 4564
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220429
transform 1 0 3832 0 1 4564
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220429
transform 1 0 5656 0 -1 4492
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220429
transform 1 0 3832 0 -1 4492
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220429
transform 1 0 5656 0 1 4316
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220429
transform 1 0 3832 0 1 4316
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220429
transform 1 0 5656 0 -1 4268
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220429
transform 1 0 3832 0 -1 4268
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220429
transform 1 0 5656 0 1 4008
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220429
transform 1 0 3832 0 1 4008
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220429
transform 1 0 5656 0 -1 3952
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220429
transform 1 0 3832 0 -1 3952
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220429
transform 1 0 5656 0 1 3744
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220429
transform 1 0 3832 0 1 3744
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220429
transform 1 0 5656 0 -1 3676
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220429
transform 1 0 3832 0 -1 3676
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220429
transform 1 0 5656 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220429
transform 1 0 3832 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220429
transform 1 0 5656 0 -1 3412
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220429
transform 1 0 3832 0 -1 3412
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220429
transform 1 0 5656 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220429
transform 1 0 3832 0 1 3236
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220429
transform 1 0 5656 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220429
transform 1 0 3832 0 -1 3180
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220429
transform 1 0 5656 0 1 3000
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220429
transform 1 0 3832 0 1 3000
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220429
transform 1 0 5656 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220429
transform 1 0 3832 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220429
transform 1 0 5656 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220429
transform 1 0 3832 0 1 2772
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220429
transform 1 0 5656 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220429
transform 1 0 3832 0 -1 2708
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220429
transform 1 0 5656 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220429
transform 1 0 3832 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220429
transform 1 0 5656 0 -1 2468
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220429
transform 1 0 3832 0 -1 2468
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220429
transform 1 0 5656 0 1 2292
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220429
transform 1 0 3832 0 1 2292
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220429
transform 1 0 5656 0 -1 2232
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220429
transform 1 0 3832 0 -1 2232
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220429
transform 1 0 5656 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220429
transform 1 0 3832 0 1 2048
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220429
transform 1 0 5656 0 -1 1996
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220429
transform 1 0 3832 0 -1 1996
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220429
transform 1 0 5656 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220429
transform 1 0 3832 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220429
transform 1 0 5656 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220429
transform 1 0 3832 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220429
transform 1 0 5656 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220429
transform 1 0 3832 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220429
transform 1 0 5656 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220429
transform 1 0 3832 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220429
transform 1 0 5656 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220429
transform 1 0 3832 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220429
transform 1 0 5656 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220429
transform 1 0 3832 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220429
transform 1 0 5656 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220429
transform 1 0 3832 0 1 1112
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220429
transform 1 0 5656 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220429
transform 1 0 3832 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220429
transform 1 0 5656 0 1 856
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220429
transform 1 0 3832 0 1 856
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220429
transform 1 0 5656 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220429
transform 1 0 3832 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220429
transform 1 0 5656 0 1 600
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220429
transform 1 0 3832 0 1 600
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220429
transform 1 0 5656 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220429
transform 1 0 3832 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220429
transform 1 0 5656 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220429
transform 1 0 3832 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220429
transform 1 0 5656 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220429
transform 1 0 3832 0 -1 328
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220429
transform 1 0 5656 0 1 124
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220429
transform 1 0 3832 0 1 124
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220429
transform 1 0 3792 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220429
transform 1 0 1968 0 1 5604
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220429
transform 1 0 3792 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220429
transform 1 0 1968 0 -1 5556
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220429
transform 1 0 3792 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220429
transform 1 0 1968 0 1 5372
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220429
transform 1 0 3792 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220429
transform 1 0 1968 0 -1 5324
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220429
transform 1 0 3792 0 1 5148
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220429
transform 1 0 1968 0 1 5148
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220429
transform 1 0 3792 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220429
transform 1 0 1968 0 -1 5076
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220429
transform 1 0 3792 0 1 4880
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220429
transform 1 0 1968 0 1 4880
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220429
transform 1 0 3792 0 -1 4804
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220429
transform 1 0 1968 0 -1 4804
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220429
transform 1 0 3792 0 1 4620
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220429
transform 1 0 1968 0 1 4620
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220429
transform 1 0 3792 0 -1 4572
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220429
transform 1 0 1968 0 -1 4572
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220429
transform 1 0 3792 0 1 4356
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220429
transform 1 0 1968 0 1 4356
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220429
transform 1 0 3792 0 -1 4304
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220429
transform 1 0 1968 0 -1 4304
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220429
transform 1 0 3792 0 1 4116
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220429
transform 1 0 1968 0 1 4116
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220429
transform 1 0 3792 0 -1 4064
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220429
transform 1 0 1968 0 -1 4064
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220429
transform 1 0 3792 0 1 3888
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220429
transform 1 0 1968 0 1 3888
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220429
transform 1 0 3792 0 -1 3836
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220429
transform 1 0 1968 0 -1 3836
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220429
transform 1 0 3792 0 1 3652
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220429
transform 1 0 1968 0 1 3652
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220429
transform 1 0 3792 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220429
transform 1 0 1968 0 -1 3600
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220429
transform 1 0 3792 0 1 3400
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220429
transform 1 0 1968 0 1 3400
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220429
transform 1 0 3792 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220429
transform 1 0 1968 0 -1 3340
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220429
transform 1 0 3792 0 1 3160
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220429
transform 1 0 1968 0 1 3160
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220429
transform 1 0 3792 0 -1 3112
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220429
transform 1 0 1968 0 -1 3112
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220429
transform 1 0 3792 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220429
transform 1 0 1968 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220429
transform 1 0 3792 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220429
transform 1 0 1968 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220429
transform 1 0 3792 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220429
transform 1 0 1968 0 1 2436
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220429
transform 1 0 3792 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220429
transform 1 0 1968 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220429
transform 1 0 3792 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220429
transform 1 0 1968 0 1 2204
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220429
transform 1 0 3792 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220429
transform 1 0 1968 0 -1 2152
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220429
transform 1 0 3792 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220429
transform 1 0 1968 0 1 1968
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220429
transform 1 0 3792 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220429
transform 1 0 1968 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220429
transform 1 0 3792 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220429
transform 1 0 1968 0 1 1736
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220429
transform 1 0 3792 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220429
transform 1 0 1968 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220429
transform 1 0 3792 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220429
transform 1 0 1968 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220429
transform 1 0 3792 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220429
transform 1 0 1968 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220429
transform 1 0 3792 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220429
transform 1 0 1968 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220429
transform 1 0 3792 0 -1 1164
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220429
transform 1 0 1968 0 -1 1164
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220429
transform 1 0 3792 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220429
transform 1 0 1968 0 1 988
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220429
transform 1 0 3792 0 -1 940
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220429
transform 1 0 1968 0 -1 940
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220429
transform 1 0 3792 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220429
transform 1 0 1968 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220429
transform 1 0 3792 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220429
transform 1 0 1968 0 -1 712
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220429
transform 1 0 3792 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220429
transform 1 0 1968 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220429
transform 1 0 3792 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220429
transform 1 0 1968 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220429
transform 1 0 3792 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220429
transform 1 0 1968 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220429
transform 1 0 1928 0 -1 5696
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220429
transform 1 0 104 0 -1 5696
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220429
transform 1 0 1928 0 1 5516
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220429
transform 1 0 104 0 1 5516
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220429
transform 1 0 1928 0 -1 5456
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220429
transform 1 0 104 0 -1 5456
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220429
transform 1 0 1928 0 1 5176
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220429
transform 1 0 104 0 1 5176
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220429
transform 1 0 1928 0 -1 5112
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220429
transform 1 0 104 0 -1 5112
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220429
transform 1 0 1928 0 1 4936
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220429
transform 1 0 104 0 1 4936
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220429
transform 1 0 1928 0 -1 4888
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220429
transform 1 0 104 0 -1 4888
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220429
transform 1 0 1928 0 1 4700
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220429
transform 1 0 104 0 1 4700
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220429
transform 1 0 1928 0 -1 4648
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220429
transform 1 0 104 0 -1 4648
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220429
transform 1 0 1928 0 1 4460
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220429
transform 1 0 104 0 1 4460
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220429
transform 1 0 1928 0 -1 4412
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220429
transform 1 0 104 0 -1 4412
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220429
transform 1 0 1928 0 1 4228
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220429
transform 1 0 104 0 1 4228
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220429
transform 1 0 1928 0 -1 4168
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220429
transform 1 0 104 0 -1 4168
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220429
transform 1 0 1928 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220429
transform 1 0 104 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220429
transform 1 0 1928 0 -1 3920
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220429
transform 1 0 104 0 -1 3920
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220429
transform 1 0 1928 0 1 3736
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220429
transform 1 0 104 0 1 3736
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220429
transform 1 0 1928 0 -1 3676
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220429
transform 1 0 104 0 -1 3676
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220429
transform 1 0 1928 0 1 3480
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220429
transform 1 0 104 0 1 3480
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220429
transform 1 0 1928 0 -1 3412
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220429
transform 1 0 104 0 -1 3412
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220429
transform 1 0 1928 0 1 3220
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220429
transform 1 0 104 0 1 3220
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220429
transform 1 0 1928 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220429
transform 1 0 104 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220429
transform 1 0 1928 0 1 2980
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220429
transform 1 0 104 0 1 2980
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220429
transform 1 0 1928 0 -1 2932
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220429
transform 1 0 104 0 -1 2932
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220429
transform 1 0 1928 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220429
transform 1 0 104 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220429
transform 1 0 1928 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220429
transform 1 0 104 0 -1 2692
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220429
transform 1 0 1928 0 1 2512
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220429
transform 1 0 104 0 1 2512
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220429
transform 1 0 1928 0 -1 2456
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220429
transform 1 0 104 0 -1 2456
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220429
transform 1 0 1928 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220429
transform 1 0 104 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220429
transform 1 0 1928 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220429
transform 1 0 104 0 -1 2220
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220429
transform 1 0 1928 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220429
transform 1 0 104 0 1 2044
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220429
transform 1 0 1928 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220429
transform 1 0 104 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220429
transform 1 0 1928 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220429
transform 1 0 104 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220429
transform 1 0 1928 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220429
transform 1 0 104 0 -1 1764
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220429
transform 1 0 1928 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220429
transform 1 0 104 0 1 1588
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220429
transform 1 0 1928 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220429
transform 1 0 104 0 -1 1540
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220429
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220429
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220429
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220429
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220429
transform 1 0 1928 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220429
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220429
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220429
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220429
transform 1 0 1928 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220429
transform 1 0 104 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220429
transform 1 0 1928 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220429
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220429
transform 1 0 1928 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220429
transform 1 0 104 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220429
transform 1 0 1928 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220429
transform 1 0 104 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220429
transform 1 0 1928 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220429
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220429
transform 1 0 1928 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220429
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220429
transform 1 0 1928 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220429
transform 1 0 104 0 1 120
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220429
transform 1 0 5512 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220429
transform 1 0 5376 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220429
transform 1 0 5512 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220429
transform 1 0 5496 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220429
transform 1 0 5496 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220429
transform 1 0 5512 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220429
transform 1 0 5512 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220429
transform 1 0 5512 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220429
transform 1 0 5464 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220429
transform 1 0 5512 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220429
transform 1 0 5240 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220429
transform 1 0 5288 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220429
transform 1 0 5280 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220429
transform 1 0 5136 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220429
transform 1 0 5328 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220429
transform 1 0 5240 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220429
transform 1 0 5104 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220429
transform 1 0 4968 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220429
transform 1 0 4832 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220429
transform 1 0 4696 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220429
transform 1 0 4560 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220429
transform 1 0 4424 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220429
transform 1 0 4288 0 1 100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220429
transform 1 0 4608 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220429
transform 1 0 4776 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220429
transform 1 0 4952 0 -1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220429
transform 1 0 5048 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220429
transform 1 0 4816 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220429
transform 1 0 4592 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220429
transform 1 0 4376 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220429
transform 1 0 5088 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220429
transform 1 0 4896 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220429
transform 1 0 4712 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220429
transform 1 0 4544 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220429
transform 1 0 4992 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220429
transform 1 0 4752 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220429
transform 1 0 4528 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220429
transform 1 0 4320 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220429
transform 1 0 4136 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220429
transform 1 0 3952 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220429
transform 1 0 4208 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220429
transform 1 0 4504 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220429
transform 1 0 4832 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220429
transform 1 0 5184 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220429
transform 1 0 4936 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220429
transform 1 0 4752 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220429
transform 1 0 4584 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220429
transform 1 0 5128 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220429
transform 1 0 5328 0 1 832
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220429
transform 1 0 5376 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220429
transform 1 0 5240 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220429
transform 1 0 5104 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220429
transform 1 0 4968 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220429
transform 1 0 4832 0 -1 1068
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220429
transform 1 0 5272 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220429
transform 1 0 5040 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220429
transform 1 0 4808 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220429
transform 1 0 4576 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220429
transform 1 0 4336 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220429
transform 1 0 5192 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220429
transform 1 0 4920 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220429
transform 1 0 4664 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220429
transform 1 0 4424 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220429
transform 1 0 4208 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220429
transform 1 0 5160 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220429
transform 1 0 4864 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220429
transform 1 0 4592 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220429
transform 1 0 4352 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220429
transform 1 0 4144 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220429
transform 1 0 5160 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220429
transform 1 0 4824 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220429
transform 1 0 4512 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220429
transform 1 0 4480 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220429
transform 1 0 4280 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220429
transform 1 0 5256 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220429
transform 1 0 4976 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220429
transform 1 0 4712 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220429
transform 1 0 4528 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220429
transform 1 0 4336 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220429
transform 1 0 4736 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220429
transform 1 0 5184 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220429
transform 1 0 4952 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220429
transform 1 0 4840 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220429
transform 1 0 4680 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220429
transform 1 0 5176 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220429
transform 1 0 5008 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220429
transform 1 0 4968 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220429
transform 1 0 4832 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220429
transform 1 0 5104 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220429
transform 1 0 5376 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220429
transform 1 0 5240 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220429
transform 1 0 5376 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220429
transform 1 0 5352 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220429
transform 1 0 5416 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220429
transform 1 0 5456 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220429
transform 1 0 5496 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220429
transform 1 0 5512 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220429
transform 1 0 5512 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220429
transform 1 0 5512 0 -1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220429
transform 1 0 5512 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220429
transform 1 0 5512 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220429
transform 1 0 5512 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220429
transform 1 0 5464 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220429
transform 1 0 5416 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220429
transform 1 0 5416 0 -1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220429
transform 1 0 5184 0 -1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220429
transform 1 0 5024 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220429
transform 1 0 5184 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220429
transform 1 0 5344 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220429
transform 1 0 5360 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220429
transform 1 0 5184 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220429
transform 1 0 4920 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220429
transform 1 0 4784 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220429
transform 1 0 5216 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220429
transform 1 0 5064 0 1 2024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220429
transform 1 0 5016 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220429
transform 1 0 4856 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220429
transform 1 0 4704 0 -1 2256
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220429
transform 1 0 4704 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220429
transform 1 0 4864 0 1 2268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220429
transform 1 0 4728 0 -1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220429
transform 1 0 4504 0 -1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220429
transform 1 0 4952 0 -1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220429
transform 1 0 5184 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220429
transform 1 0 4904 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220429
transform 1 0 4640 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220429
transform 1 0 4392 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220429
transform 1 0 4176 0 1 2492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220429
transform 1 0 5224 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220429
transform 1 0 5032 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220429
transform 1 0 4848 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220429
transform 1 0 4680 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220429
transform 1 0 4536 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220429
transform 1 0 4536 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220429
transform 1 0 4400 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220429
transform 1 0 4808 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220429
transform 1 0 4672 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220429
transform 1 0 4608 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220429
transform 1 0 4360 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220429
transform 1 0 4144 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220429
transform 1 0 5192 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220429
transform 1 0 4888 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220429
transform 1 0 4480 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220429
transform 1 0 4304 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220429
transform 1 0 5088 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220429
transform 1 0 4872 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220429
transform 1 0 4672 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220429
transform 1 0 4536 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220429
transform 1 0 4712 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220429
transform 1 0 5320 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220429
transform 1 0 5104 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220429
transform 1 0 4904 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220429
transform 1 0 4832 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220429
transform 1 0 4696 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220429
transform 1 0 4968 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220429
transform 1 0 5104 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220429
transform 1 0 5376 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220429
transform 1 0 5416 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220429
transform 1 0 5280 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220429
transform 1 0 5144 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220429
transform 1 0 5008 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220429
transform 1 0 4872 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220429
transform 1 0 5176 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220429
transform 1 0 5008 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220429
transform 1 0 4848 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220429
transform 1 0 4696 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220429
transform 1 0 4552 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220429
transform 1 0 5072 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220429
transform 1 0 4848 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220429
transform 1 0 4640 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220429
transform 1 0 4448 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220429
transform 1 0 4272 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220429
transform 1 0 5008 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220429
transform 1 0 4760 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220429
transform 1 0 4528 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220429
transform 1 0 4320 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220429
transform 1 0 4136 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220429
transform 1 0 4152 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220429
transform 1 0 4288 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220429
transform 1 0 4424 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220429
transform 1 0 4560 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220429
transform 1 0 4696 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220429
transform 1 0 4832 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220429
transform 1 0 4968 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220429
transform 1 0 5104 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220429
transform 1 0 5240 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220429
transform 1 0 5376 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220429
transform 1 0 5272 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220429
transform 1 0 5304 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220429
transform 1 0 5352 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220429
transform 1 0 5240 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220429
transform 1 0 5312 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220429
transform 1 0 5496 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220429
transform 1 0 5512 0 1 2976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220429
transform 1 0 5512 0 -1 3204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220429
transform 1 0 5512 0 1 3212
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220429
transform 1 0 5512 0 1 3448
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220429
transform 1 0 5512 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220429
transform 1 0 5512 0 1 3720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220429
transform 1 0 5512 0 -1 3976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220429
transform 1 0 5512 0 1 3984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220429
transform 1 0 5512 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220429
transform 1 0 5512 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220429
transform 1 0 5512 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220429
transform 1 0 5512 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220429
transform 1 0 5504 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220429
transform 1 0 5496 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220429
transform 1 0 5480 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220429
transform 1 0 5464 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220429
transform 1 0 5184 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220429
transform 1 0 5496 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220429
transform 1 0 5512 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220429
transform 1 0 5336 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220429
transform 1 0 5136 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220429
transform 1 0 4936 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220429
transform 1 0 4736 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220429
transform 1 0 5280 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220429
transform 1 0 5048 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220429
transform 1 0 4816 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220429
transform 1 0 4584 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220429
transform 1 0 5104 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220429
transform 1 0 4968 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220429
transform 1 0 4832 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220429
transform 1 0 4696 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220429
transform 1 0 4560 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220429
transform 1 0 4424 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220429
transform 1 0 4288 0 1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220429
transform 1 0 4096 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220429
transform 1 0 4344 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220429
transform 1 0 4304 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220429
transform 1 0 4528 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220429
transform 1 0 4312 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220429
transform 1 0 4584 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220429
transform 1 0 4880 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220429
transform 1 0 4608 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220429
transform 1 0 4360 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220429
transform 1 0 4152 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220429
transform 1 0 5168 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220429
transform 1 0 4880 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220429
transform 1 0 4800 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220429
transform 1 0 4600 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220429
transform 1 0 4416 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220429
transform 1 0 5248 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220429
transform 1 0 5016 0 -1 5044
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220429
transform 1 0 4984 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220429
transform 1 0 4824 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220429
transform 1 0 4672 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220429
transform 1 0 5320 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220429
transform 1 0 5152 0 1 4804
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220429
transform 1 0 5096 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220429
transform 1 0 4960 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220429
transform 1 0 4824 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220429
transform 1 0 5232 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220429
transform 1 0 5368 0 -1 4784
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220429
transform 1 0 5336 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220429
transform 1 0 5168 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220429
transform 1 0 5008 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220429
transform 1 0 4856 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220429
transform 1 0 4712 0 1 4540
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220429
transform 1 0 5240 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220429
transform 1 0 4976 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220429
transform 1 0 4720 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220429
transform 1 0 4472 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220429
transform 1 0 4792 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220429
transform 1 0 5024 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220429
transform 1 0 5272 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220429
transform 1 0 5224 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220429
transform 1 0 4928 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220429
transform 1 0 4648 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220429
transform 1 0 4400 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220429
transform 1 0 4192 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220429
transform 1 0 4016 0 -1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220429
transform 1 0 4584 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220429
transform 1 0 4400 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220429
transform 1 0 4264 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220429
transform 1 0 4128 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220429
transform 1 0 3992 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220429
transform 1 0 4248 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220429
transform 1 0 4032 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220429
transform 1 0 3856 0 -1 4516
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220429
transform 1 0 3856 0 1 4292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220429
transform 1 0 3648 0 1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220429
transform 1 0 3648 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220429
transform 1 0 3488 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220429
transform 1 0 3312 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220429
transform 1 0 3136 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220429
transform 1 0 2952 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220429
transform 1 0 2832 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220429
transform 1 0 3048 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220429
transform 1 0 3648 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220429
transform 1 0 3464 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220429
transform 1 0 3256 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220429
transform 1 0 3248 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220429
transform 1 0 3040 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220429
transform 1 0 2824 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220429
transform 1 0 3456 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220429
transform 1 0 3648 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220429
transform 1 0 3648 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220429
transform 1 0 3456 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220429
transform 1 0 3240 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220429
transform 1 0 3024 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220429
transform 1 0 2800 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220429
transform 1 0 3648 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220429
transform 1 0 3472 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220429
transform 1 0 3280 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220429
transform 1 0 3088 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220429
transform 1 0 2888 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220429
transform 1 0 3472 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220429
transform 1 0 3272 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220429
transform 1 0 3072 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220429
transform 1 0 2872 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220429
transform 1 0 2664 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220429
transform 1 0 3272 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220429
transform 1 0 3104 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220429
transform 1 0 2936 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220429
transform 1 0 2776 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220429
transform 1 0 2616 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220429
transform 1 0 3096 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220429
transform 1 0 2944 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220429
transform 1 0 2792 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220429
transform 1 0 2640 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220429
transform 1 0 2488 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220429
transform 1 0 2520 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220429
transform 1 0 2696 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220429
transform 1 0 2864 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220429
transform 1 0 3040 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220429
transform 1 0 3216 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220429
transform 1 0 3048 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220429
transform 1 0 2848 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220429
transform 1 0 2648 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220429
transform 1 0 3448 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220429
transform 1 0 3248 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220429
transform 1 0 3144 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220429
transform 1 0 2880 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220429
transform 1 0 2600 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220429
transform 1 0 3648 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220429
transform 1 0 3408 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220429
transform 1 0 3376 0 1 2904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220429
transform 1 0 3240 0 1 2904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220429
transform 1 0 3104 0 1 2904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220429
transform 1 0 3512 0 1 2904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220429
transform 1 0 3648 0 1 2904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220429
transform 1 0 3856 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220429
transform 1 0 3992 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220429
transform 1 0 3856 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220429
transform 1 0 3992 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220429
transform 1 0 4128 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220429
transform 1 0 4264 0 1 2748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220429
transform 1 0 4400 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220429
transform 1 0 4264 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220429
transform 1 0 4128 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220429
transform 1 0 3992 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220429
transform 1 0 3856 0 -1 2732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220429
transform 1 0 3648 0 -1 2636
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220429
transform 1 0 3512 0 -1 2636
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220429
transform 1 0 3376 0 -1 2636
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220429
transform 1 0 3240 0 -1 2636
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220429
transform 1 0 3648 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220429
transform 1 0 3448 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220429
transform 1 0 3224 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220429
transform 1 0 3000 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220429
transform 1 0 2768 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220429
transform 1 0 3496 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220429
transform 1 0 3328 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220429
transform 1 0 3160 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220429
transform 1 0 3000 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220429
transform 1 0 2840 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220429
transform 1 0 3360 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220429
transform 1 0 3224 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220429
transform 1 0 3088 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220429
transform 1 0 2952 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220429
transform 1 0 2816 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220429
transform 1 0 2808 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220429
transform 1 0 2672 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220429
transform 1 0 2944 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220429
transform 1 0 3080 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220429
transform 1 0 3216 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220429
transform 1 0 3088 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220429
transform 1 0 3240 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220429
transform 1 0 3392 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220429
transform 1 0 3320 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220429
transform 1 0 3176 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220429
transform 1 0 3192 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220429
transform 1 0 3040 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220429
transform 1 0 2888 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220429
transform 1 0 2768 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220429
transform 1 0 2904 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220429
transform 1 0 3040 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220429
transform 1 0 2944 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220429
transform 1 0 2808 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220429
transform 1 0 2672 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220429
transform 1 0 2536 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220429
transform 1 0 2680 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220429
transform 1 0 2544 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220429
transform 1 0 2408 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220429
transform 1 0 2272 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220429
transform 1 0 2136 0 1 2180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220429
transform 1 0 2680 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220429
transform 1 0 2512 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220429
transform 1 0 2344 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220429
transform 1 0 2184 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220429
transform 1 0 2024 0 -1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220429
transform 1 0 2520 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220429
transform 1 0 2248 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220429
transform 1 0 1992 0 1 2412
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220429
transform 1 0 1784 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220429
transform 1 0 1640 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220429
transform 1 0 1480 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220429
transform 1 0 1320 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220429
transform 1 0 1152 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220429
transform 1 0 1784 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220429
transform 1 0 1648 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220429
transform 1 0 1504 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220429
transform 1 0 1352 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220429
transform 1 0 1208 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220429
transform 1 0 1280 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220429
transform 1 0 1448 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220429
transform 1 0 1616 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220429
transform 1 0 1784 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220429
transform 1 0 1784 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220429
transform 1 0 1632 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220429
transform 1 0 1456 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220429
transform 1 0 1352 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220429
transform 1 0 1576 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220429
transform 1 0 1784 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220429
transform 1 0 1992 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220429
transform 1 0 2296 0 -1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220429
transform 1 0 2432 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220429
transform 1 0 2208 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220429
transform 1 0 1992 0 1 3136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220429
transform 1 0 1992 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220429
transform 1 0 2160 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220429
transform 1 0 2344 0 -1 3364
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220429
transform 1 0 2336 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220429
transform 1 0 2184 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220429
transform 1 0 2032 0 1 3376
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220429
transform 1 0 2104 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220429
transform 1 0 2280 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220429
transform 1 0 2448 0 -1 3624
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220429
transform 1 0 2448 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220429
transform 1 0 2224 0 1 3628
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220429
transform 1 0 2208 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220429
transform 1 0 2672 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220429
transform 1 0 2448 0 -1 3860
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220429
transform 1 0 2320 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220429
transform 1 0 2568 0 1 3864
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220429
transform 1 0 2592 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220429
transform 1 0 2344 0 -1 4088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220429
transform 1 0 2368 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220429
transform 1 0 2608 0 1 4092
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220429
transform 1 0 2760 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220429
transform 1 0 2568 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220429
transform 1 0 2368 0 -1 4328
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220429
transform 1 0 2568 0 1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220429
transform 1 0 3120 0 1 4332
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220429
transform 1 0 3016 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220429
transform 1 0 2840 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220429
transform 1 0 2664 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220429
transform 1 0 2496 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220429
transform 1 0 2744 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220429
transform 1 0 2904 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220429
transform 1 0 3064 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220429
transform 1 0 3232 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220429
transform 1 0 3208 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220429
transform 1 0 3064 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220429
transform 1 0 3496 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220429
transform 1 0 3352 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220429
transform 1 0 3320 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220429
transform 1 0 3648 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220429
transform 1 0 3496 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220429
transform 1 0 3408 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220429
transform 1 0 3648 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220429
transform 1 0 3856 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220429
transform 1 0 3992 0 1 5060
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220429
transform 1 0 3856 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220429
transform 1 0 4064 0 -1 5292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220429
transform 1 0 4072 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220429
transform 1 0 3856 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220429
transform 1 0 3856 0 -1 5536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220429
transform 1 0 3648 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220429
transform 1 0 3432 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220429
transform 1 0 3648 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220429
transform 1 0 3496 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220429
transform 1 0 3320 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220429
transform 1 0 3144 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220429
transform 1 0 2960 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220429
transform 1 0 2776 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220429
transform 1 0 2952 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220429
transform 1 0 3192 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220429
transform 1 0 3072 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220429
transform 1 0 3288 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220429
transform 1 0 3256 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220429
transform 1 0 3256 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220429
transform 1 0 3144 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220429
transform 1 0 2880 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220429
transform 1 0 2816 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220429
transform 1 0 3152 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220429
transform 1 0 2984 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220429
transform 1 0 2920 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220429
transform 1 0 2776 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220429
transform 1 0 2632 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220429
transform 1 0 2496 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220429
transform 1 0 2360 0 -1 4828
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220429
transform 1 0 2584 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220429
transform 1 0 2424 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220429
transform 1 0 2264 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220429
transform 1 0 2128 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220429
transform 1 0 1992 0 1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220429
transform 1 0 2320 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220429
transform 1 0 2144 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220429
transform 1 0 1992 0 -1 4596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220429
transform 1 0 1784 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220429
transform 1 0 1576 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220429
transform 1 0 1344 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220429
transform 1 0 1408 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220429
transform 1 0 1600 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220429
transform 1 0 1784 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220429
transform 1 0 1696 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220429
transform 1 0 1560 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220429
transform 1 0 1424 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220429
transform 1 0 1512 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220429
transform 1 0 1784 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220429
transform 1 0 1648 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220429
transform 1 0 1576 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220429
transform 1 0 1440 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220429
transform 1 0 1712 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220429
transform 1 0 1648 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220429
transform 1 0 1488 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220429
transform 1 0 1328 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220429
transform 1 0 1272 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220429
transform 1 0 1456 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220429
transform 1 0 1640 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220429
transform 1 0 1624 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220429
transform 1 0 1424 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220429
transform 1 0 1224 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220429
transform 1 0 1160 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220429
transform 1 0 1376 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220429
transform 1 0 1592 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220429
transform 1 0 1560 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220429
transform 1 0 1336 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220429
transform 1 0 1112 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220429
transform 1 0 1072 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220429
transform 1 0 1296 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220429
transform 1 0 1520 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220429
transform 1 0 1480 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220429
transform 1 0 1232 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220429
transform 1 0 992 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220429
transform 1 0 880 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220429
transform 1 0 1120 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220429
transform 1 0 1280 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220429
transform 1 0 1104 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220429
transform 1 0 920 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220429
transform 1 0 936 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220429
transform 1 0 1112 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220429
transform 1 0 1056 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220429
transform 1 0 904 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220429
transform 1 0 744 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220429
transform 1 0 808 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220429
transform 1 0 984 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220429
transform 1 0 1184 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220429
transform 1 0 984 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220429
transform 1 0 784 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220429
transform 1 0 592 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220429
transform 1 0 480 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220429
transform 1 0 672 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220429
transform 1 0 864 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220429
transform 1 0 712 0 -1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220429
transform 1 0 560 0 -1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220429
transform 1 0 552 0 1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220429
transform 1 0 1008 0 1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220429
transform 1 0 776 0 1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220429
transform 1 0 768 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220429
transform 1 0 1112 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220429
transform 1 0 1456 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220429
transform 1 0 1152 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220429
transform 1 0 928 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220429
transform 1 0 696 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220429
transform 1 0 448 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220429
transform 1 0 640 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220429
transform 1 0 864 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220429
transform 1 0 1088 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220429
transform 1 0 1112 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220429
transform 1 0 880 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220429
transform 1 0 664 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220429
transform 1 0 736 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220429
transform 1 0 840 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220429
transform 1 0 584 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220429
transform 1 0 520 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220429
transform 1 0 696 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220429
transform 1 0 520 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220429
transform 1 0 432 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220429
transform 1 0 632 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220429
transform 1 0 544 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220429
transform 1 0 368 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220429
transform 1 0 720 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220429
transform 1 0 904 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220429
transform 1 0 1088 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220429
transform 1 0 1048 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220429
transform 1 0 840 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220429
transform 1 0 808 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220429
transform 1 0 664 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220429
transform 1 0 944 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220429
transform 1 0 864 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220429
transform 1 0 1032 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220429
transform 1 0 1360 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220429
transform 1 0 1096 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220429
transform 1 0 920 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220429
transform 1 0 1096 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220429
transform 1 0 1272 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220429
transform 1 0 1632 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220429
transform 1 0 1448 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220429
transform 1 0 1352 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220429
transform 1 0 1592 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220429
transform 1 0 1768 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220429
transform 1 0 1536 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220429
transform 1 0 1312 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220429
transform 1 0 1368 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220429
transform 1 0 1584 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220429
transform 1 0 1784 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220429
transform 1 0 1784 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220429
transform 1 0 1992 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220429
transform 1 0 2128 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220429
transform 1 0 2128 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220429
transform 1 0 1992 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220429
transform 1 0 2264 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220429
transform 1 0 2400 0 -1 2176
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220429
transform 1 0 2264 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220429
transform 1 0 2400 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220429
transform 1 0 2536 0 1 1944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220429
transform 1 0 2496 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220429
transform 1 0 2632 0 -1 1936
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220429
transform 1 0 2584 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220429
transform 1 0 2440 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220429
transform 1 0 2736 0 1 1712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220429
transform 1 0 2936 0 -1 1668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220429
transform 1 0 2568 0 -1 1668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220429
transform 1 0 2200 0 -1 1668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220429
transform 1 0 1992 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220429
transform 1 0 2272 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220429
transform 1 0 2536 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220429
transform 1 0 2800 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220429
transform 1 0 2584 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220429
transform 1 0 2368 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220429
transform 1 0 2160 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220429
transform 1 0 1992 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220429
transform 1 0 1784 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220429
transform 1 0 1648 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220429
transform 1 0 1496 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220429
transform 1 0 1344 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220429
transform 1 0 1192 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220429
transform 1 0 1088 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220429
transform 1 0 1232 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220429
transform 1 0 1376 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220429
transform 1 0 1512 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220429
transform 1 0 1648 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220429
transform 1 0 1784 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220429
transform 1 0 1992 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220429
transform 1 0 2128 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220429
transform 1 0 2272 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220429
transform 1 0 2624 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220429
transform 1 0 2440 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220429
transform 1 0 2336 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220429
transform 1 0 2200 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220429
transform 1 0 2064 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220429
transform 1 0 2304 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220429
transform 1 0 2480 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220429
transform 1 0 2824 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220429
transform 1 0 2656 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220429
transform 1 0 2624 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220429
transform 1 0 2472 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220429
transform 1 0 2800 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220429
transform 1 0 3424 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220429
transform 1 0 3200 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220429
transform 1 0 2992 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220429
transform 1 0 2816 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220429
transform 1 0 3024 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220429
transform 1 0 3232 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220429
transform 1 0 3224 0 -1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220429
transform 1 0 3088 0 -1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220429
transform 1 0 2952 0 -1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220429
transform 1 0 3088 0 1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220429
transform 1 0 3224 0 1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220429
transform 1 0 3360 0 1 1188
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220429
transform 1 0 3496 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220429
transform 1 0 3256 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220429
transform 1 0 3024 0 -1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220429
transform 1 0 3008 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220429
transform 1 0 2776 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220429
transform 1 0 3232 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220429
transform 1 0 3648 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220429
transform 1 0 3448 0 1 1432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220429
transform 1 0 3304 0 -1 1668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220429
transform 1 0 3648 0 -1 1668
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220429
transform 1 0 3856 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220429
transform 1 0 3856 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220429
transform 1 0 3992 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220429
transform 1 0 4160 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220429
transform 1 0 4128 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220429
transform 1 0 3992 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220429
transform 1 0 4240 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220429
transform 1 0 4016 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220429
transform 1 0 3856 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220429
transform 1 0 3856 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220429
transform 1 0 3992 0 1 1324
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220429
transform 1 0 3856 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220429
transform 1 0 4016 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220429
transform 1 0 4088 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220429
transform 1 0 3856 0 1 1088
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220429
transform 1 0 3648 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220429
transform 1 0 3448 0 1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220429
transform 1 0 3648 0 -1 964
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220429
transform 1 0 3648 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220429
transform 1 0 3496 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220429
transform 1 0 3328 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220429
transform 1 0 3160 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220429
transform 1 0 2992 0 1 740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220429
transform 1 0 3104 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220429
transform 1 0 3240 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220429
transform 1 0 3376 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220429
transform 1 0 3512 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220429
transform 1 0 3648 0 -1 736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220429
transform 1 0 3856 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220429
transform 1 0 3992 0 1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220429
transform 1 0 4400 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220429
transform 1 0 4264 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220429
transform 1 0 4128 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220429
transform 1 0 3992 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220429
transform 1 0 3856 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220429
transform 1 0 3648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220429
transform 1 0 3472 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220429
transform 1 0 3272 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220429
transform 1 0 3072 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220429
transform 1 0 2864 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220429
transform 1 0 3624 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220429
transform 1 0 3488 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220429
transform 1 0 3352 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220429
transform 1 0 3216 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220429
transform 1 0 3080 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220429
transform 1 0 2944 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220429
transform 1 0 3624 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220429
transform 1 0 3488 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220429
transform 1 0 3352 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220429
transform 1 0 3216 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220429
transform 1 0 3080 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220429
transform 1 0 2944 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220429
transform 1 0 2808 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220429
transform 1 0 2672 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220429
transform 1 0 2536 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220429
transform 1 0 2536 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220429
transform 1 0 2400 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220429
transform 1 0 2264 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220429
transform 1 0 2128 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220429
transform 1 0 1992 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220429
transform 1 0 2808 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220429
transform 1 0 2672 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220429
transform 1 0 2400 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220429
transform 1 0 2264 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220429
transform 1 0 2128 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220429
transform 1 0 1992 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220429
transform 1 0 2648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220429
transform 1 0 2424 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220429
transform 1 0 2200 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220429
transform 1 0 1992 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220429
transform 1 0 1784 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220429
transform 1 0 1616 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220429
transform 1 0 1432 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220429
transform 1 0 1432 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220429
transform 1 0 1616 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220429
transform 1 0 1784 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220429
transform 1 0 1656 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220429
transform 1 0 1368 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220429
transform 1 0 1248 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220429
transform 1 0 1056 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220429
transform 1 0 1064 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220429
transform 1 0 1248 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220429
transform 1 0 1408 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220429
transform 1 0 1192 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220429
transform 1 0 1136 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220429
transform 1 0 1312 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220429
transform 1 0 1488 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220429
transform 1 0 1352 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220429
transform 1 0 1216 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220429
transform 1 0 1080 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220429
transform 1 0 944 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220429
transform 1 0 808 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220429
transform 1 0 672 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220429
transform 1 0 536 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220429
transform 1 0 616 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220429
transform 1 0 784 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220429
transform 1 0 960 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220429
transform 1 0 984 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220429
transform 1 0 784 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220429
transform 1 0 584 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220429
transform 1 0 392 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220429
transform 1 0 872 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220429
transform 1 0 680 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220429
transform 1 0 488 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220429
transform 1 0 296 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220429
transform 1 0 128 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220429
transform 1 0 864 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220429
transform 1 0 672 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220429
transform 1 0 480 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220429
transform 1 0 288 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220429
transform 1 0 128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220429
transform 1 0 128 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220429
transform 1 0 320 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220429
transform 1 0 1080 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220429
transform 1 0 808 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220429
transform 1 0 552 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220429
transform 1 0 192 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220429
transform 1 0 232 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220429
transform 1 0 232 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220429
transform 1 0 376 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220429
transform 1 0 336 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220429
transform 1 0 328 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220429
transform 1 0 352 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220429
transform 1 0 544 0 -1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220429
transform 1 0 456 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220429
transform 1 0 272 0 1 1564
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220429
transform 1 0 416 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220429
transform 1 0 200 0 -1 1788
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220429
transform 1 0 192 0 1 1792
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220429
transform 1 0 128 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220429
transform 1 0 432 0 -1 2016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220429
transform 1 0 328 0 1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220429
transform 1 0 128 0 1 2020
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220429
transform 1 0 128 0 -1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220429
transform 1 0 408 0 -1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220429
transform 1 0 264 0 -1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220429
transform 1 0 128 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220429
transform 1 0 288 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220429
transform 1 0 192 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220429
transform 1 0 392 0 -1 2480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220429
transform 1 0 232 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220429
transform 1 0 432 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220429
transform 1 0 624 0 1 2488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220429
transform 1 0 584 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220429
transform 1 0 416 0 -1 2716
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220429
transform 1 0 360 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220429
transform 1 0 560 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220429
transform 1 0 752 0 1 2720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220429
transform 1 0 728 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220429
transform 1 0 520 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220429
transform 1 0 312 0 -1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220429
transform 1 0 352 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220429
transform 1 0 624 0 1 2956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220429
transform 1 0 752 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220429
transform 1 0 512 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220429
transform 1 0 272 0 -1 3180
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220429
transform 1 0 208 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220429
transform 1 0 848 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220429
transform 1 0 632 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220429
transform 1 0 416 0 1 3196
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220429
transform 1 0 224 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220429
transform 1 0 888 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220429
transform 1 0 664 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220429
transform 1 0 440 0 -1 3436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220429
transform 1 0 376 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220429
transform 1 0 200 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220429
transform 1 0 952 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220429
transform 1 0 752 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220429
transform 1 0 560 0 1 3456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220429
transform 1 0 464 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220429
transform 1 0 296 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220429
transform 1 0 1024 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220429
transform 1 0 832 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220429
transform 1 0 648 0 -1 3700
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220429
transform 1 0 584 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220429
transform 1 0 424 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220429
transform 1 0 1096 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220429
transform 1 0 920 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220429
transform 1 0 752 0 1 3712
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220429
transform 1 0 712 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220429
transform 1 0 568 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220429
transform 1 0 1168 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220429
transform 1 0 1016 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220429
transform 1 0 864 0 -1 3944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220429
transform 1 0 760 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220429
transform 1 0 624 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220429
transform 1 0 896 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220429
transform 1 0 1304 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220429
transform 1 0 1168 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220429
transform 1 0 1032 0 1 3956
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220429
transform 1 0 968 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220429
transform 1 0 832 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220429
transform 1 0 696 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220429
transform 1 0 1104 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220429
transform 1 0 1240 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220429
transform 1 0 1376 0 -1 4192
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220429
transform 1 0 1288 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220429
transform 1 0 1152 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220429
transform 1 0 1016 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220429
transform 1 0 880 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220429
transform 1 0 744 0 1 4204
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220429
transform 1 0 1216 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220429
transform 1 0 1032 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220429
transform 1 0 856 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220429
transform 1 0 688 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220429
transform 1 0 528 0 -1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220429
transform 1 0 1120 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220429
transform 1 0 904 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220429
transform 1 0 688 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220429
transform 1 0 488 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220429
transform 1 0 296 0 1 4436
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220429
transform 1 0 672 0 -1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220429
transform 1 0 536 0 -1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220429
transform 1 0 400 0 -1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220429
transform 1 0 264 0 -1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220429
transform 1 0 128 0 -1 4672
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220429
transform 1 0 672 0 1 4676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220429
transform 1 0 536 0 1 4676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220429
transform 1 0 400 0 1 4676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220429
transform 1 0 264 0 1 4676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220429
transform 1 0 128 0 1 4676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220429
transform 1 0 128 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220429
transform 1 0 384 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220429
transform 1 0 1432 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220429
transform 1 0 1056 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220429
transform 1 0 704 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220429
transform 1 0 408 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220429
transform 1 0 136 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220429
transform 1 0 960 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220429
transform 1 0 680 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220429
transform 1 0 472 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220429
transform 1 0 288 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220429
transform 1 0 1120 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220429
transform 1 0 888 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220429
transform 1 0 672 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220429
transform 1 0 592 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220429
transform 1 0 456 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220429
transform 1 0 728 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220429
transform 1 0 864 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220429
transform 1 0 1000 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220429
transform 1 0 1136 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220429
transform 1 0 1272 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220429
transform 1 0 1544 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220429
transform 1 0 1408 0 1 5152
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220429
transform 1 0 1360 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220429
transform 1 0 1600 0 -1 5136
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220429
transform 1 0 1520 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220429
transform 1 0 1240 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220429
transform 1 0 1784 0 1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220429
transform 1 0 1784 0 -1 4912
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220429
transform 1 0 1992 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220429
transform 1 0 2128 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220429
transform 1 0 2296 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220429
transform 1 0 2464 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220429
transform 1 0 2640 0 1 4856
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220429
transform 1 0 2608 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220429
transform 1 0 2328 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220429
transform 1 0 2048 0 -1 5100
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220429
transform 1 0 2096 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220429
transform 1 0 2232 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220429
transform 1 0 2376 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220429
transform 1 0 2528 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220429
transform 1 0 2696 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220429
transform 1 0 2880 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220429
transform 1 0 3064 0 1 5124
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220429
transform 1 0 3104 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220429
transform 1 0 2960 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220429
transform 1 0 2824 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220429
transform 1 0 2688 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220429
transform 1 0 2552 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220429
transform 1 0 2416 0 -1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220429
transform 1 0 2424 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220429
transform 1 0 2640 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220429
transform 1 0 2856 0 1 5348
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220429
transform 1 0 2712 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220429
transform 1 0 2472 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220429
transform 1 0 2232 0 -1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220429
transform 1 0 2584 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220429
transform 1 0 2384 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220429
transform 1 0 2176 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220429
transform 1 0 1992 0 1 5580
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220429
transform 1 0 1784 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220429
transform 1 0 1512 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220429
transform 1 0 1400 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220429
transform 1 0 1576 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220429
transform 1 0 1760 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220429
transform 1 0 1784 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220429
transform 1 0 1648 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220429
transform 1 0 1512 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220429
transform 1 0 1376 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220429
transform 1 0 1240 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220429
transform 1 0 1104 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220429
transform 1 0 968 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220429
transform 1 0 832 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220429
transform 1 0 696 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220429
transform 1 0 560 0 -1 5480
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220429
transform 1 0 1224 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220429
transform 1 0 1048 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220429
transform 1 0 880 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220429
transform 1 0 720 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220429
transform 1 0 560 0 1 5492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220429
transform 1 0 1224 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220429
transform 1 0 952 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220429
transform 1 0 696 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220429
transform 1 0 472 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220429
transform 1 0 272 0 -1 5720
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220429
transform 1 0 128 0 -1 5720
box 3 5 132 108
<< end >>
