magic
tech sky130l
timestamp 1730768468
<< m1 >>
rect 1656 1363 1660 1505
rect 336 1279 340 1303
rect 216 1135 220 1273
rect 408 615 412 639
rect 616 615 620 639
rect 848 615 852 639
<< m2c >>
rect 232 1729 236 1733
rect 368 1729 372 1733
rect 504 1729 508 1733
rect 640 1729 644 1733
rect 776 1729 780 1733
rect 111 1725 115 1729
rect 1719 1725 1723 1729
rect 111 1707 115 1711
rect 1719 1707 1723 1711
rect 111 1637 115 1641
rect 1719 1637 1723 1641
rect 111 1619 115 1623
rect 1719 1619 1723 1623
rect 304 1615 308 1619
rect 440 1615 444 1619
rect 576 1615 580 1619
rect 712 1615 716 1619
rect 848 1615 852 1619
rect 584 1505 588 1509
rect 720 1505 724 1509
rect 856 1505 860 1509
rect 992 1505 996 1509
rect 1128 1505 1132 1509
rect 1264 1505 1268 1509
rect 1400 1505 1404 1509
rect 1536 1505 1540 1509
rect 1656 1505 1660 1509
rect 1672 1505 1676 1509
rect 111 1501 115 1505
rect 111 1483 115 1487
rect 111 1409 115 1413
rect 111 1391 115 1395
rect 696 1387 700 1391
rect 832 1387 836 1391
rect 968 1387 972 1391
rect 1112 1387 1116 1391
rect 1256 1387 1260 1391
rect 1400 1387 1404 1391
rect 1536 1387 1540 1391
rect 1719 1501 1723 1505
rect 1719 1483 1723 1487
rect 1719 1409 1723 1413
rect 1719 1391 1723 1395
rect 1672 1387 1676 1391
rect 1656 1359 1660 1363
rect 336 1303 340 1307
rect 216 1273 220 1277
rect 232 1273 236 1277
rect 336 1275 340 1279
rect 440 1273 444 1277
rect 704 1273 708 1277
rect 992 1273 996 1277
rect 1304 1273 1308 1277
rect 1616 1273 1620 1277
rect 111 1269 115 1273
rect 111 1251 115 1255
rect 111 1181 115 1185
rect 111 1163 115 1167
rect 1719 1269 1723 1273
rect 1719 1251 1723 1255
rect 1719 1181 1723 1185
rect 1719 1163 1723 1167
rect 232 1159 236 1163
rect 400 1159 404 1163
rect 616 1159 620 1163
rect 848 1159 852 1163
rect 1096 1159 1100 1163
rect 1360 1159 1364 1163
rect 1624 1159 1628 1163
rect 216 1131 220 1135
rect 408 1041 412 1045
rect 632 1041 636 1045
rect 872 1041 876 1045
rect 1120 1041 1124 1045
rect 1376 1041 1380 1045
rect 1640 1041 1644 1045
rect 111 1037 115 1041
rect 1719 1037 1723 1041
rect 111 1019 115 1023
rect 1719 1019 1723 1023
rect 111 961 115 965
rect 1719 961 1723 965
rect 111 943 115 947
rect 1719 943 1723 947
rect 600 939 604 943
rect 784 939 788 943
rect 992 939 996 943
rect 1208 939 1212 943
rect 1440 939 1444 943
rect 1672 939 1676 943
rect 840 825 844 829
rect 976 825 980 829
rect 1112 825 1116 829
rect 1248 825 1252 829
rect 1384 825 1388 829
rect 1528 825 1532 829
rect 1672 825 1676 829
rect 111 821 115 825
rect 1719 821 1723 825
rect 111 803 115 807
rect 1719 803 1723 807
rect 111 729 115 733
rect 1719 729 1723 733
rect 111 711 115 715
rect 1719 711 1723 715
rect 776 707 780 711
rect 936 707 940 711
rect 1104 707 1108 711
rect 1288 707 1292 711
rect 1472 707 1476 711
rect 1664 707 1668 711
rect 408 639 412 643
rect 320 609 324 613
rect 408 611 412 615
rect 616 639 620 643
rect 512 609 516 613
rect 616 611 620 615
rect 848 639 852 643
rect 720 609 724 613
rect 848 611 852 615
rect 952 609 956 613
rect 1192 609 1196 613
rect 1432 609 1436 613
rect 111 605 115 609
rect 1719 605 1723 609
rect 111 587 115 591
rect 1719 587 1723 591
rect 111 517 115 521
rect 1719 517 1723 521
rect 111 499 115 503
rect 1719 499 1723 503
rect 232 495 236 499
rect 400 495 404 499
rect 616 495 620 499
rect 856 495 860 499
rect 1112 495 1116 499
rect 1376 495 1380 499
rect 1640 495 1644 499
rect 296 381 300 385
rect 528 381 532 385
rect 760 381 764 385
rect 984 381 988 385
rect 1208 381 1212 385
rect 1432 381 1436 385
rect 1656 381 1660 385
rect 111 377 115 381
rect 1719 377 1723 381
rect 111 359 115 363
rect 1719 359 1723 363
rect 111 289 115 293
rect 1719 289 1723 293
rect 111 271 115 275
rect 1719 271 1723 275
rect 512 267 516 271
rect 728 267 732 271
rect 952 267 956 271
rect 1192 267 1196 271
rect 1440 267 1444 271
rect 1672 267 1676 271
rect 584 157 588 161
rect 720 157 724 161
rect 856 157 860 161
rect 992 157 996 161
rect 1128 157 1132 161
rect 1264 157 1268 161
rect 1400 157 1404 161
rect 1672 157 1676 161
rect 111 153 115 157
rect 1719 153 1723 157
rect 111 135 115 139
rect 1719 135 1723 139
<< m2 >>
rect 246 1759 252 1760
rect 246 1755 247 1759
rect 251 1758 252 1759
rect 386 1759 392 1760
rect 251 1756 281 1758
rect 251 1755 252 1756
rect 246 1754 252 1755
rect 386 1755 387 1759
rect 391 1758 392 1759
rect 522 1759 528 1760
rect 391 1756 417 1758
rect 391 1755 392 1756
rect 386 1754 392 1755
rect 522 1755 523 1759
rect 527 1758 528 1759
rect 658 1759 664 1760
rect 527 1756 553 1758
rect 527 1755 528 1756
rect 522 1754 528 1755
rect 658 1755 659 1759
rect 663 1758 664 1759
rect 663 1756 689 1758
rect 663 1755 664 1756
rect 658 1754 664 1755
rect 231 1733 237 1734
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 231 1729 232 1733
rect 236 1732 237 1733
rect 246 1733 252 1734
rect 246 1732 247 1733
rect 236 1730 247 1732
rect 236 1729 237 1730
rect 231 1728 237 1729
rect 246 1729 247 1730
rect 251 1729 252 1733
rect 246 1728 252 1729
rect 367 1733 373 1734
rect 367 1729 368 1733
rect 372 1732 373 1733
rect 386 1733 392 1734
rect 386 1732 387 1733
rect 372 1730 387 1732
rect 372 1729 373 1730
rect 367 1728 373 1729
rect 386 1729 387 1730
rect 391 1729 392 1733
rect 386 1728 392 1729
rect 503 1733 509 1734
rect 503 1729 504 1733
rect 508 1732 509 1733
rect 522 1733 528 1734
rect 522 1732 523 1733
rect 508 1730 523 1732
rect 508 1729 509 1730
rect 503 1728 509 1729
rect 522 1729 523 1730
rect 527 1729 528 1733
rect 522 1728 528 1729
rect 639 1733 645 1734
rect 639 1729 640 1733
rect 644 1732 645 1733
rect 658 1733 664 1734
rect 658 1732 659 1733
rect 644 1730 659 1732
rect 644 1729 645 1730
rect 639 1728 645 1729
rect 658 1729 659 1730
rect 663 1729 664 1733
rect 658 1728 664 1729
rect 766 1733 772 1734
rect 766 1729 767 1733
rect 771 1732 772 1733
rect 775 1733 781 1734
rect 775 1732 776 1733
rect 771 1730 776 1732
rect 771 1729 772 1730
rect 766 1728 772 1729
rect 775 1729 776 1730
rect 780 1729 781 1733
rect 775 1728 781 1729
rect 1718 1729 1724 1730
rect 110 1724 116 1725
rect 134 1727 140 1728
rect 134 1723 135 1727
rect 139 1723 140 1727
rect 134 1722 140 1723
rect 270 1727 276 1728
rect 270 1723 271 1727
rect 275 1723 276 1727
rect 270 1722 276 1723
rect 406 1727 412 1728
rect 406 1723 407 1727
rect 411 1723 412 1727
rect 406 1722 412 1723
rect 542 1727 548 1728
rect 542 1723 543 1727
rect 547 1723 548 1727
rect 542 1722 548 1723
rect 678 1727 684 1728
rect 678 1723 679 1727
rect 683 1723 684 1727
rect 1718 1725 1719 1729
rect 1723 1725 1724 1729
rect 1718 1724 1724 1725
rect 678 1722 684 1723
rect 158 1712 164 1713
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 158 1708 159 1712
rect 163 1708 164 1712
rect 158 1707 164 1708
rect 294 1712 300 1713
rect 294 1708 295 1712
rect 299 1708 300 1712
rect 294 1707 300 1708
rect 430 1712 436 1713
rect 430 1708 431 1712
rect 435 1708 436 1712
rect 430 1707 436 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 702 1712 708 1713
rect 702 1708 703 1712
rect 707 1708 708 1712
rect 702 1707 708 1708
rect 1718 1711 1724 1712
rect 1718 1707 1719 1711
rect 1723 1707 1724 1711
rect 110 1706 116 1707
rect 1718 1706 1724 1707
rect 110 1641 116 1642
rect 1718 1641 1724 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 110 1636 116 1637
rect 230 1640 236 1641
rect 230 1636 231 1640
rect 235 1636 236 1640
rect 230 1635 236 1636
rect 366 1640 372 1641
rect 366 1636 367 1640
rect 371 1636 372 1640
rect 366 1635 372 1636
rect 502 1640 508 1641
rect 502 1636 503 1640
rect 507 1636 508 1640
rect 502 1635 508 1636
rect 638 1640 644 1641
rect 638 1636 639 1640
rect 643 1636 644 1640
rect 638 1635 644 1636
rect 774 1640 780 1641
rect 774 1636 775 1640
rect 779 1636 780 1640
rect 1718 1637 1719 1641
rect 1723 1637 1724 1641
rect 1718 1636 1724 1637
rect 774 1635 780 1636
rect 206 1625 212 1626
rect 110 1623 116 1624
rect 110 1619 111 1623
rect 115 1619 116 1623
rect 206 1621 207 1625
rect 211 1621 212 1625
rect 206 1620 212 1621
rect 342 1625 348 1626
rect 342 1621 343 1625
rect 347 1621 348 1625
rect 342 1620 348 1621
rect 478 1625 484 1626
rect 478 1621 479 1625
rect 483 1621 484 1625
rect 478 1620 484 1621
rect 614 1625 620 1626
rect 614 1621 615 1625
rect 619 1621 620 1625
rect 614 1620 620 1621
rect 750 1625 756 1626
rect 750 1621 751 1625
rect 755 1621 756 1625
rect 750 1620 756 1621
rect 1718 1623 1724 1624
rect 110 1618 116 1619
rect 303 1619 309 1620
rect 303 1615 304 1619
rect 308 1618 309 1619
rect 350 1619 356 1620
rect 350 1618 351 1619
rect 308 1616 351 1618
rect 308 1615 309 1616
rect 303 1614 309 1615
rect 350 1615 351 1616
rect 355 1615 356 1619
rect 350 1614 356 1615
rect 439 1619 445 1620
rect 439 1615 440 1619
rect 444 1618 445 1619
rect 486 1619 492 1620
rect 486 1618 487 1619
rect 444 1616 487 1618
rect 444 1615 445 1616
rect 439 1614 445 1615
rect 486 1615 487 1616
rect 491 1615 492 1619
rect 486 1614 492 1615
rect 575 1619 581 1620
rect 575 1615 576 1619
rect 580 1618 581 1619
rect 622 1619 628 1620
rect 622 1618 623 1619
rect 580 1616 623 1618
rect 580 1615 581 1616
rect 575 1614 581 1615
rect 622 1615 623 1616
rect 627 1615 628 1619
rect 622 1614 628 1615
rect 711 1619 717 1620
rect 711 1615 712 1619
rect 716 1618 717 1619
rect 758 1619 764 1620
rect 758 1618 759 1619
rect 716 1616 759 1618
rect 716 1615 717 1616
rect 711 1614 717 1615
rect 758 1615 759 1616
rect 763 1615 764 1619
rect 847 1619 853 1620
rect 847 1618 848 1619
rect 758 1614 764 1615
rect 768 1616 848 1618
rect 594 1611 600 1612
rect 594 1607 595 1611
rect 599 1610 600 1611
rect 768 1610 770 1616
rect 847 1615 848 1616
rect 852 1615 853 1619
rect 1718 1619 1719 1623
rect 1723 1619 1724 1623
rect 1718 1618 1724 1619
rect 847 1614 853 1615
rect 599 1608 770 1610
rect 599 1607 600 1608
rect 594 1606 600 1607
rect 766 1599 772 1600
rect 766 1598 767 1599
rect 284 1596 767 1598
rect 284 1589 286 1596
rect 766 1595 767 1596
rect 771 1595 772 1599
rect 766 1594 772 1595
rect 350 1591 356 1592
rect 350 1587 351 1591
rect 355 1587 356 1591
rect 350 1586 356 1587
rect 486 1591 492 1592
rect 486 1587 487 1591
rect 491 1587 492 1591
rect 486 1586 492 1587
rect 622 1591 628 1592
rect 622 1587 623 1591
rect 627 1587 628 1591
rect 622 1586 628 1587
rect 758 1591 764 1592
rect 758 1587 759 1591
rect 763 1587 764 1591
rect 758 1586 764 1587
rect 594 1539 600 1540
rect 594 1538 595 1539
rect 565 1536 595 1538
rect 594 1535 595 1536
rect 599 1535 600 1539
rect 1274 1539 1280 1540
rect 1274 1538 1275 1539
rect 1245 1536 1275 1538
rect 594 1534 600 1535
rect 602 1535 608 1536
rect 602 1531 603 1535
rect 607 1534 608 1535
rect 738 1535 744 1536
rect 607 1532 633 1534
rect 607 1531 608 1532
rect 602 1530 608 1531
rect 738 1531 739 1535
rect 743 1534 744 1535
rect 874 1535 880 1536
rect 743 1532 769 1534
rect 743 1531 744 1532
rect 738 1530 744 1531
rect 874 1531 875 1535
rect 879 1534 880 1535
rect 1010 1535 1016 1536
rect 879 1532 905 1534
rect 879 1531 880 1532
rect 874 1530 880 1531
rect 1010 1531 1011 1535
rect 1015 1534 1016 1535
rect 1274 1535 1275 1536
rect 1279 1535 1280 1539
rect 1274 1534 1280 1535
rect 1282 1535 1288 1536
rect 1015 1532 1041 1534
rect 1015 1531 1016 1532
rect 1010 1530 1016 1531
rect 1282 1531 1283 1535
rect 1287 1534 1288 1535
rect 1418 1535 1424 1536
rect 1287 1532 1313 1534
rect 1287 1531 1288 1532
rect 1282 1530 1288 1531
rect 1418 1531 1419 1535
rect 1423 1534 1424 1535
rect 1554 1535 1560 1536
rect 1423 1532 1449 1534
rect 1423 1531 1424 1532
rect 1418 1530 1424 1531
rect 1554 1531 1555 1535
rect 1559 1534 1560 1535
rect 1559 1532 1585 1534
rect 1559 1531 1560 1532
rect 1554 1530 1560 1531
rect 583 1509 589 1510
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 583 1505 584 1509
rect 588 1508 589 1509
rect 602 1509 608 1510
rect 602 1508 603 1509
rect 588 1506 603 1508
rect 588 1505 589 1506
rect 583 1504 589 1505
rect 602 1505 603 1506
rect 607 1505 608 1509
rect 602 1504 608 1505
rect 719 1509 725 1510
rect 719 1505 720 1509
rect 724 1508 725 1509
rect 738 1509 744 1510
rect 738 1508 739 1509
rect 724 1506 739 1508
rect 724 1505 725 1506
rect 719 1504 725 1505
rect 738 1505 739 1506
rect 743 1505 744 1509
rect 738 1504 744 1505
rect 855 1509 861 1510
rect 855 1505 856 1509
rect 860 1508 861 1509
rect 874 1509 880 1510
rect 874 1508 875 1509
rect 860 1506 875 1508
rect 860 1505 861 1506
rect 855 1504 861 1505
rect 874 1505 875 1506
rect 879 1505 880 1509
rect 874 1504 880 1505
rect 991 1509 997 1510
rect 991 1505 992 1509
rect 996 1508 997 1509
rect 1010 1509 1016 1510
rect 1010 1508 1011 1509
rect 996 1506 1011 1508
rect 996 1505 997 1506
rect 991 1504 997 1505
rect 1010 1505 1011 1506
rect 1015 1505 1016 1509
rect 1010 1504 1016 1505
rect 1110 1509 1116 1510
rect 1110 1505 1111 1509
rect 1115 1508 1116 1509
rect 1127 1509 1133 1510
rect 1127 1508 1128 1509
rect 1115 1506 1128 1508
rect 1115 1505 1116 1506
rect 1110 1504 1116 1505
rect 1127 1505 1128 1506
rect 1132 1505 1133 1509
rect 1127 1504 1133 1505
rect 1263 1509 1269 1510
rect 1263 1505 1264 1509
rect 1268 1508 1269 1509
rect 1282 1509 1288 1510
rect 1282 1508 1283 1509
rect 1268 1506 1283 1508
rect 1268 1505 1269 1506
rect 1263 1504 1269 1505
rect 1282 1505 1283 1506
rect 1287 1505 1288 1509
rect 1282 1504 1288 1505
rect 1399 1509 1405 1510
rect 1399 1505 1400 1509
rect 1404 1508 1405 1509
rect 1418 1509 1424 1510
rect 1418 1508 1419 1509
rect 1404 1506 1419 1508
rect 1404 1505 1405 1506
rect 1399 1504 1405 1505
rect 1418 1505 1419 1506
rect 1423 1505 1424 1509
rect 1418 1504 1424 1505
rect 1535 1509 1541 1510
rect 1535 1505 1536 1509
rect 1540 1508 1541 1509
rect 1554 1509 1560 1510
rect 1554 1508 1555 1509
rect 1540 1506 1555 1508
rect 1540 1505 1541 1506
rect 1535 1504 1541 1505
rect 1554 1505 1555 1506
rect 1559 1505 1560 1509
rect 1554 1504 1560 1505
rect 1655 1509 1661 1510
rect 1655 1505 1656 1509
rect 1660 1508 1661 1509
rect 1671 1509 1677 1510
rect 1671 1508 1672 1509
rect 1660 1506 1672 1508
rect 1660 1505 1661 1506
rect 1655 1504 1661 1505
rect 1671 1505 1672 1506
rect 1676 1505 1677 1509
rect 1671 1504 1677 1505
rect 1718 1505 1724 1506
rect 110 1500 116 1501
rect 486 1503 492 1504
rect 486 1499 487 1503
rect 491 1499 492 1503
rect 486 1498 492 1499
rect 622 1503 628 1504
rect 622 1499 623 1503
rect 627 1499 628 1503
rect 622 1498 628 1499
rect 758 1503 764 1504
rect 758 1499 759 1503
rect 763 1499 764 1503
rect 758 1498 764 1499
rect 894 1503 900 1504
rect 894 1499 895 1503
rect 899 1499 900 1503
rect 894 1498 900 1499
rect 1030 1503 1036 1504
rect 1030 1499 1031 1503
rect 1035 1499 1036 1503
rect 1030 1498 1036 1499
rect 1166 1503 1172 1504
rect 1166 1499 1167 1503
rect 1171 1499 1172 1503
rect 1166 1498 1172 1499
rect 1302 1503 1308 1504
rect 1302 1499 1303 1503
rect 1307 1499 1308 1503
rect 1302 1498 1308 1499
rect 1438 1503 1444 1504
rect 1438 1499 1439 1503
rect 1443 1499 1444 1503
rect 1438 1498 1444 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1499 1580 1503
rect 1718 1501 1719 1505
rect 1723 1501 1724 1505
rect 1718 1500 1724 1501
rect 1574 1498 1580 1499
rect 510 1488 516 1489
rect 110 1487 116 1488
rect 110 1483 111 1487
rect 115 1483 116 1487
rect 510 1484 511 1488
rect 515 1484 516 1488
rect 510 1483 516 1484
rect 646 1488 652 1489
rect 646 1484 647 1488
rect 651 1484 652 1488
rect 646 1483 652 1484
rect 782 1488 788 1489
rect 782 1484 783 1488
rect 787 1484 788 1488
rect 782 1483 788 1484
rect 918 1488 924 1489
rect 918 1484 919 1488
rect 923 1484 924 1488
rect 918 1483 924 1484
rect 1054 1488 1060 1489
rect 1054 1484 1055 1488
rect 1059 1484 1060 1488
rect 1054 1483 1060 1484
rect 1190 1488 1196 1489
rect 1190 1484 1191 1488
rect 1195 1484 1196 1488
rect 1190 1483 1196 1484
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1462 1483 1468 1484
rect 1598 1488 1604 1489
rect 1598 1484 1599 1488
rect 1603 1484 1604 1488
rect 1598 1483 1604 1484
rect 1718 1487 1724 1488
rect 1718 1483 1719 1487
rect 1723 1483 1724 1487
rect 110 1482 116 1483
rect 1718 1482 1724 1483
rect 110 1413 116 1414
rect 1718 1413 1724 1414
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 110 1408 116 1409
rect 622 1412 628 1413
rect 622 1408 623 1412
rect 627 1408 628 1412
rect 622 1407 628 1408
rect 758 1412 764 1413
rect 758 1408 759 1412
rect 763 1408 764 1412
rect 758 1407 764 1408
rect 894 1412 900 1413
rect 894 1408 895 1412
rect 899 1408 900 1412
rect 894 1407 900 1408
rect 1038 1412 1044 1413
rect 1038 1408 1039 1412
rect 1043 1408 1044 1412
rect 1038 1407 1044 1408
rect 1182 1412 1188 1413
rect 1182 1408 1183 1412
rect 1187 1408 1188 1412
rect 1182 1407 1188 1408
rect 1326 1412 1332 1413
rect 1326 1408 1327 1412
rect 1331 1408 1332 1412
rect 1326 1407 1332 1408
rect 1462 1412 1468 1413
rect 1462 1408 1463 1412
rect 1467 1408 1468 1412
rect 1462 1407 1468 1408
rect 1598 1412 1604 1413
rect 1598 1408 1599 1412
rect 1603 1408 1604 1412
rect 1718 1409 1719 1413
rect 1723 1409 1724 1413
rect 1718 1408 1724 1409
rect 1598 1407 1604 1408
rect 598 1397 604 1398
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 598 1393 599 1397
rect 603 1393 604 1397
rect 598 1392 604 1393
rect 734 1397 740 1398
rect 734 1393 735 1397
rect 739 1393 740 1397
rect 734 1392 740 1393
rect 870 1397 876 1398
rect 870 1393 871 1397
rect 875 1393 876 1397
rect 870 1392 876 1393
rect 1014 1397 1020 1398
rect 1014 1393 1015 1397
rect 1019 1393 1020 1397
rect 1014 1392 1020 1393
rect 1158 1397 1164 1398
rect 1158 1393 1159 1397
rect 1163 1393 1164 1397
rect 1158 1392 1164 1393
rect 1302 1397 1308 1398
rect 1302 1393 1303 1397
rect 1307 1393 1308 1397
rect 1302 1392 1308 1393
rect 1438 1397 1444 1398
rect 1438 1393 1439 1397
rect 1443 1393 1444 1397
rect 1438 1392 1444 1393
rect 1574 1397 1580 1398
rect 1574 1393 1575 1397
rect 1579 1393 1580 1397
rect 1574 1392 1580 1393
rect 1718 1395 1724 1396
rect 110 1390 116 1391
rect 695 1391 701 1392
rect 695 1387 696 1391
rect 700 1390 701 1391
rect 742 1391 748 1392
rect 742 1390 743 1391
rect 700 1388 743 1390
rect 700 1387 701 1388
rect 695 1386 701 1387
rect 742 1387 743 1388
rect 747 1387 748 1391
rect 742 1386 748 1387
rect 831 1391 837 1392
rect 831 1387 832 1391
rect 836 1390 837 1391
rect 878 1391 884 1392
rect 878 1390 879 1391
rect 836 1388 879 1390
rect 836 1387 837 1388
rect 831 1386 837 1387
rect 878 1387 879 1388
rect 883 1387 884 1391
rect 878 1386 884 1387
rect 967 1391 976 1392
rect 967 1387 968 1391
rect 975 1387 976 1391
rect 1111 1391 1117 1392
rect 1111 1390 1112 1391
rect 967 1386 976 1387
rect 980 1388 1112 1390
rect 674 1383 680 1384
rect 674 1379 675 1383
rect 679 1382 680 1383
rect 980 1382 982 1388
rect 1111 1387 1112 1388
rect 1116 1387 1117 1391
rect 1111 1386 1117 1387
rect 1254 1391 1261 1392
rect 1254 1387 1255 1391
rect 1260 1387 1261 1391
rect 1254 1386 1261 1387
rect 1278 1391 1284 1392
rect 1278 1387 1279 1391
rect 1283 1390 1284 1391
rect 1399 1391 1405 1392
rect 1399 1390 1400 1391
rect 1283 1388 1400 1390
rect 1283 1387 1284 1388
rect 1278 1386 1284 1387
rect 1399 1387 1400 1388
rect 1404 1387 1405 1391
rect 1399 1386 1405 1387
rect 1534 1391 1541 1392
rect 1534 1387 1535 1391
rect 1540 1387 1541 1391
rect 1534 1386 1541 1387
rect 1558 1391 1564 1392
rect 1558 1387 1559 1391
rect 1563 1390 1564 1391
rect 1671 1391 1677 1392
rect 1671 1390 1672 1391
rect 1563 1388 1672 1390
rect 1563 1387 1564 1388
rect 1558 1386 1564 1387
rect 1671 1387 1672 1388
rect 1676 1387 1677 1391
rect 1718 1391 1719 1395
rect 1723 1391 1724 1395
rect 1718 1390 1724 1391
rect 1671 1386 1677 1387
rect 679 1380 982 1382
rect 679 1379 680 1380
rect 674 1378 680 1379
rect 970 1371 976 1372
rect 970 1367 971 1371
rect 975 1370 976 1371
rect 975 1368 1161 1370
rect 975 1367 976 1368
rect 970 1366 976 1367
rect 674 1363 680 1364
rect 674 1359 675 1363
rect 679 1359 680 1363
rect 674 1358 680 1359
rect 742 1363 748 1364
rect 742 1359 743 1363
rect 747 1359 748 1363
rect 742 1358 748 1359
rect 878 1363 884 1364
rect 878 1359 879 1363
rect 883 1359 884 1363
rect 1110 1363 1116 1364
rect 1110 1362 1111 1363
rect 1093 1360 1111 1362
rect 878 1358 884 1359
rect 1110 1359 1111 1360
rect 1115 1359 1116 1363
rect 1159 1362 1161 1368
rect 1358 1363 1364 1364
rect 1159 1360 1169 1362
rect 1110 1358 1116 1359
rect 1358 1359 1359 1363
rect 1363 1359 1364 1363
rect 1558 1363 1564 1364
rect 1558 1362 1559 1363
rect 1517 1360 1559 1362
rect 1358 1358 1364 1359
rect 1558 1359 1559 1360
rect 1563 1359 1564 1363
rect 1655 1363 1661 1364
rect 1655 1362 1656 1363
rect 1653 1360 1656 1362
rect 1558 1358 1564 1359
rect 1655 1359 1656 1360
rect 1660 1359 1661 1363
rect 1655 1358 1661 1359
rect 335 1307 341 1308
rect 335 1306 336 1307
rect 213 1304 336 1306
rect 335 1303 336 1304
rect 340 1303 341 1307
rect 526 1307 532 1308
rect 526 1306 527 1307
rect 421 1304 527 1306
rect 335 1302 341 1303
rect 526 1303 527 1304
rect 531 1303 532 1307
rect 886 1307 892 1308
rect 886 1306 887 1307
rect 685 1304 887 1306
rect 526 1302 532 1303
rect 886 1303 887 1304
rect 891 1303 892 1307
rect 1198 1307 1204 1308
rect 1198 1306 1199 1307
rect 973 1304 1199 1306
rect 886 1302 892 1303
rect 1198 1303 1199 1304
rect 1203 1303 1204 1307
rect 1198 1302 1204 1303
rect 1254 1303 1260 1304
rect 1254 1299 1255 1303
rect 1259 1299 1260 1303
rect 1254 1298 1260 1299
rect 1534 1303 1540 1304
rect 1534 1299 1535 1303
rect 1539 1299 1540 1303
rect 1534 1298 1540 1299
rect 335 1279 341 1280
rect 215 1277 221 1278
rect 110 1273 116 1274
rect 110 1269 111 1273
rect 115 1269 116 1273
rect 215 1273 216 1277
rect 220 1276 221 1277
rect 231 1277 237 1278
rect 231 1276 232 1277
rect 220 1274 232 1276
rect 220 1273 221 1274
rect 215 1272 221 1273
rect 231 1273 232 1274
rect 236 1273 237 1277
rect 335 1275 336 1279
rect 340 1278 341 1279
rect 526 1279 532 1280
rect 340 1276 422 1278
rect 439 1277 445 1278
rect 439 1276 440 1277
rect 340 1275 341 1276
rect 335 1274 341 1275
rect 420 1274 440 1276
rect 231 1272 237 1273
rect 439 1273 440 1274
rect 444 1273 445 1277
rect 526 1275 527 1279
rect 531 1278 532 1279
rect 886 1279 892 1280
rect 531 1276 686 1278
rect 703 1277 709 1278
rect 703 1276 704 1277
rect 531 1275 532 1276
rect 526 1274 532 1275
rect 684 1274 704 1276
rect 439 1272 445 1273
rect 703 1273 704 1274
rect 708 1273 709 1277
rect 886 1275 887 1279
rect 891 1278 892 1279
rect 1198 1279 1204 1280
rect 891 1276 974 1278
rect 991 1277 997 1278
rect 991 1276 992 1277
rect 891 1275 892 1276
rect 886 1274 892 1275
rect 972 1274 992 1276
rect 703 1272 709 1273
rect 991 1273 992 1274
rect 996 1273 997 1277
rect 1198 1275 1199 1279
rect 1203 1278 1204 1279
rect 1203 1276 1286 1278
rect 1303 1277 1309 1278
rect 1303 1276 1304 1277
rect 1203 1275 1204 1276
rect 1198 1274 1204 1275
rect 1284 1274 1304 1276
rect 991 1272 997 1273
rect 1303 1273 1304 1274
rect 1308 1273 1309 1277
rect 1303 1272 1309 1273
rect 1602 1277 1608 1278
rect 1602 1273 1603 1277
rect 1607 1276 1608 1277
rect 1615 1277 1621 1278
rect 1615 1276 1616 1277
rect 1607 1274 1616 1276
rect 1607 1273 1608 1274
rect 1602 1272 1608 1273
rect 1615 1273 1616 1274
rect 1620 1273 1621 1277
rect 1615 1272 1621 1273
rect 1718 1273 1724 1274
rect 110 1268 116 1269
rect 134 1271 140 1272
rect 134 1267 135 1271
rect 139 1267 140 1271
rect 134 1266 140 1267
rect 342 1271 348 1272
rect 342 1267 343 1271
rect 347 1267 348 1271
rect 342 1266 348 1267
rect 606 1271 612 1272
rect 606 1267 607 1271
rect 611 1267 612 1271
rect 606 1266 612 1267
rect 894 1271 900 1272
rect 894 1267 895 1271
rect 899 1267 900 1271
rect 894 1266 900 1267
rect 1206 1271 1212 1272
rect 1206 1267 1207 1271
rect 1211 1267 1212 1271
rect 1206 1266 1212 1267
rect 1518 1271 1524 1272
rect 1518 1267 1519 1271
rect 1523 1267 1524 1271
rect 1718 1269 1719 1273
rect 1723 1269 1724 1273
rect 1718 1268 1724 1269
rect 1518 1266 1524 1267
rect 158 1256 164 1257
rect 110 1255 116 1256
rect 110 1251 111 1255
rect 115 1251 116 1255
rect 158 1252 159 1256
rect 163 1252 164 1256
rect 158 1251 164 1252
rect 366 1256 372 1257
rect 366 1252 367 1256
rect 371 1252 372 1256
rect 366 1251 372 1252
rect 630 1256 636 1257
rect 630 1252 631 1256
rect 635 1252 636 1256
rect 630 1251 636 1252
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 1230 1256 1236 1257
rect 1230 1252 1231 1256
rect 1235 1252 1236 1256
rect 1230 1251 1236 1252
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1718 1255 1724 1256
rect 1718 1251 1719 1255
rect 1723 1251 1724 1255
rect 110 1250 116 1251
rect 1718 1250 1724 1251
rect 110 1185 116 1186
rect 1718 1185 1724 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 158 1184 164 1185
rect 158 1180 159 1184
rect 163 1180 164 1184
rect 158 1179 164 1180
rect 326 1184 332 1185
rect 326 1180 327 1184
rect 331 1180 332 1184
rect 326 1179 332 1180
rect 542 1184 548 1185
rect 542 1180 543 1184
rect 547 1180 548 1184
rect 542 1179 548 1180
rect 774 1184 780 1185
rect 774 1180 775 1184
rect 779 1180 780 1184
rect 774 1179 780 1180
rect 1022 1184 1028 1185
rect 1022 1180 1023 1184
rect 1027 1180 1028 1184
rect 1022 1179 1028 1180
rect 1286 1184 1292 1185
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 1550 1184 1556 1185
rect 1550 1180 1551 1184
rect 1555 1180 1556 1184
rect 1718 1181 1719 1185
rect 1723 1181 1724 1185
rect 1718 1180 1724 1181
rect 1550 1179 1556 1180
rect 134 1169 140 1170
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 134 1165 135 1169
rect 139 1165 140 1169
rect 134 1164 140 1165
rect 302 1169 308 1170
rect 302 1165 303 1169
rect 307 1165 308 1169
rect 302 1164 308 1165
rect 518 1169 524 1170
rect 518 1165 519 1169
rect 523 1165 524 1169
rect 518 1164 524 1165
rect 750 1169 756 1170
rect 750 1165 751 1169
rect 755 1165 756 1169
rect 750 1164 756 1165
rect 998 1169 1004 1170
rect 998 1165 999 1169
rect 1003 1165 1004 1169
rect 998 1164 1004 1165
rect 1262 1169 1268 1170
rect 1262 1165 1263 1169
rect 1267 1165 1268 1169
rect 1262 1164 1268 1165
rect 1526 1169 1532 1170
rect 1526 1165 1527 1169
rect 1531 1165 1532 1169
rect 1526 1164 1532 1165
rect 1718 1167 1724 1168
rect 110 1162 116 1163
rect 231 1163 237 1164
rect 231 1159 232 1163
rect 236 1162 237 1163
rect 310 1163 316 1164
rect 310 1162 311 1163
rect 236 1160 311 1162
rect 236 1159 237 1160
rect 231 1158 237 1159
rect 310 1159 311 1160
rect 315 1159 316 1163
rect 310 1158 316 1159
rect 399 1163 405 1164
rect 399 1159 400 1163
rect 404 1162 405 1163
rect 526 1163 532 1164
rect 526 1162 527 1163
rect 404 1160 527 1162
rect 404 1159 405 1160
rect 399 1158 405 1159
rect 526 1159 527 1160
rect 531 1159 532 1163
rect 526 1158 532 1159
rect 615 1163 621 1164
rect 615 1159 616 1163
rect 620 1162 621 1163
rect 758 1163 764 1164
rect 758 1162 759 1163
rect 620 1160 759 1162
rect 620 1159 621 1160
rect 615 1158 621 1159
rect 758 1159 759 1160
rect 763 1159 764 1163
rect 758 1158 764 1159
rect 847 1163 853 1164
rect 847 1159 848 1163
rect 852 1162 853 1163
rect 1006 1163 1012 1164
rect 1006 1162 1007 1163
rect 852 1160 1007 1162
rect 852 1159 853 1160
rect 847 1158 853 1159
rect 1006 1159 1007 1160
rect 1011 1159 1012 1163
rect 1095 1163 1101 1164
rect 1095 1162 1096 1163
rect 1006 1158 1012 1159
rect 1020 1160 1096 1162
rect 418 1151 424 1152
rect 418 1147 419 1151
rect 423 1150 424 1151
rect 1020 1150 1022 1160
rect 1095 1159 1096 1160
rect 1100 1159 1101 1163
rect 1095 1158 1101 1159
rect 1358 1163 1365 1164
rect 1358 1159 1359 1163
rect 1364 1159 1365 1163
rect 1358 1158 1365 1159
rect 1618 1163 1629 1164
rect 1618 1159 1619 1163
rect 1623 1159 1624 1163
rect 1628 1159 1629 1163
rect 1718 1163 1719 1167
rect 1723 1163 1724 1167
rect 1718 1162 1724 1163
rect 1618 1158 1629 1159
rect 423 1148 1022 1150
rect 423 1147 424 1148
rect 418 1146 424 1147
rect 215 1135 221 1136
rect 215 1134 216 1135
rect 213 1132 216 1134
rect 215 1131 216 1132
rect 220 1131 221 1135
rect 215 1130 221 1131
rect 310 1135 316 1136
rect 310 1131 311 1135
rect 315 1131 316 1135
rect 310 1130 316 1131
rect 526 1135 532 1136
rect 526 1131 527 1135
rect 531 1131 532 1135
rect 526 1130 532 1131
rect 758 1135 764 1136
rect 758 1131 759 1135
rect 763 1131 764 1135
rect 758 1130 764 1131
rect 1006 1135 1012 1136
rect 1006 1131 1007 1135
rect 1011 1131 1012 1135
rect 1358 1135 1364 1136
rect 1358 1134 1359 1135
rect 1341 1132 1359 1134
rect 1006 1130 1012 1131
rect 1358 1131 1359 1132
rect 1363 1131 1364 1135
rect 1358 1130 1364 1131
rect 1602 1135 1608 1136
rect 1602 1131 1603 1135
rect 1607 1131 1608 1135
rect 1602 1130 1608 1131
rect 418 1075 424 1076
rect 418 1074 419 1075
rect 389 1072 419 1074
rect 418 1071 419 1072
rect 423 1071 424 1075
rect 1526 1075 1532 1076
rect 1526 1074 1527 1075
rect 1357 1072 1527 1074
rect 418 1070 424 1071
rect 426 1071 432 1072
rect 426 1067 427 1071
rect 431 1070 432 1071
rect 650 1071 656 1072
rect 431 1068 545 1070
rect 431 1067 432 1068
rect 426 1066 432 1067
rect 650 1067 651 1071
rect 655 1070 656 1071
rect 890 1071 896 1072
rect 655 1068 785 1070
rect 655 1067 656 1068
rect 650 1066 656 1067
rect 890 1067 891 1071
rect 895 1070 896 1071
rect 1526 1071 1527 1072
rect 1531 1071 1532 1075
rect 1526 1070 1532 1071
rect 1618 1071 1624 1072
rect 895 1068 1033 1070
rect 895 1067 896 1068
rect 890 1066 896 1067
rect 1618 1067 1619 1071
rect 1623 1067 1624 1071
rect 1618 1066 1624 1067
rect 407 1045 413 1046
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 407 1041 408 1045
rect 412 1044 413 1045
rect 426 1045 432 1046
rect 426 1044 427 1045
rect 412 1042 427 1044
rect 412 1041 413 1042
rect 407 1040 413 1041
rect 426 1041 427 1042
rect 431 1041 432 1045
rect 426 1040 432 1041
rect 631 1045 637 1046
rect 631 1041 632 1045
rect 636 1044 637 1045
rect 650 1045 656 1046
rect 650 1044 651 1045
rect 636 1042 651 1044
rect 636 1041 637 1042
rect 631 1040 637 1041
rect 650 1041 651 1042
rect 655 1041 656 1045
rect 650 1040 656 1041
rect 871 1045 877 1046
rect 871 1041 872 1045
rect 876 1044 877 1045
rect 890 1045 896 1046
rect 890 1044 891 1045
rect 876 1042 891 1044
rect 876 1041 877 1042
rect 871 1040 877 1041
rect 890 1041 891 1042
rect 895 1041 896 1045
rect 890 1040 896 1041
rect 1102 1045 1108 1046
rect 1102 1041 1103 1045
rect 1107 1044 1108 1045
rect 1119 1045 1125 1046
rect 1119 1044 1120 1045
rect 1107 1042 1120 1044
rect 1107 1041 1108 1042
rect 1102 1040 1108 1041
rect 1119 1041 1120 1042
rect 1124 1041 1125 1045
rect 1119 1040 1125 1041
rect 1358 1045 1364 1046
rect 1358 1041 1359 1045
rect 1363 1044 1364 1045
rect 1375 1045 1381 1046
rect 1375 1044 1376 1045
rect 1363 1042 1376 1044
rect 1363 1041 1364 1042
rect 1358 1040 1364 1041
rect 1375 1041 1376 1042
rect 1380 1041 1381 1045
rect 1375 1040 1381 1041
rect 1638 1045 1645 1046
rect 1638 1041 1639 1045
rect 1644 1041 1645 1045
rect 1638 1040 1645 1041
rect 1718 1041 1724 1042
rect 110 1036 116 1037
rect 310 1039 316 1040
rect 310 1035 311 1039
rect 315 1035 316 1039
rect 310 1034 316 1035
rect 534 1039 540 1040
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 774 1039 780 1040
rect 774 1035 775 1039
rect 779 1035 780 1039
rect 774 1034 780 1035
rect 1022 1039 1028 1040
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1022 1034 1028 1035
rect 1278 1039 1284 1040
rect 1278 1035 1279 1039
rect 1283 1035 1284 1039
rect 1278 1034 1284 1035
rect 1542 1039 1548 1040
rect 1542 1035 1543 1039
rect 1547 1035 1548 1039
rect 1718 1037 1719 1041
rect 1723 1037 1724 1041
rect 1718 1036 1724 1037
rect 1542 1034 1548 1035
rect 334 1024 340 1025
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 334 1020 335 1024
rect 339 1020 340 1024
rect 334 1019 340 1020
rect 558 1024 564 1025
rect 558 1020 559 1024
rect 563 1020 564 1024
rect 558 1019 564 1020
rect 798 1024 804 1025
rect 798 1020 799 1024
rect 803 1020 804 1024
rect 798 1019 804 1020
rect 1046 1024 1052 1025
rect 1046 1020 1047 1024
rect 1051 1020 1052 1024
rect 1046 1019 1052 1020
rect 1302 1024 1308 1025
rect 1302 1020 1303 1024
rect 1307 1020 1308 1024
rect 1302 1019 1308 1020
rect 1566 1024 1572 1025
rect 1566 1020 1567 1024
rect 1571 1020 1572 1024
rect 1566 1019 1572 1020
rect 1718 1023 1724 1024
rect 1718 1019 1719 1023
rect 1723 1019 1724 1023
rect 110 1018 116 1019
rect 1718 1018 1724 1019
rect 110 965 116 966
rect 1718 965 1724 966
rect 110 961 111 965
rect 115 961 116 965
rect 110 960 116 961
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 710 964 716 965
rect 710 960 711 964
rect 715 960 716 964
rect 710 959 716 960
rect 918 964 924 965
rect 918 960 919 964
rect 923 960 924 964
rect 918 959 924 960
rect 1134 964 1140 965
rect 1134 960 1135 964
rect 1139 960 1140 964
rect 1134 959 1140 960
rect 1366 964 1372 965
rect 1366 960 1367 964
rect 1371 960 1372 964
rect 1366 959 1372 960
rect 1598 964 1604 965
rect 1598 960 1599 964
rect 1603 960 1604 964
rect 1718 961 1719 965
rect 1723 961 1724 965
rect 1718 960 1724 961
rect 1598 959 1604 960
rect 502 949 508 950
rect 110 947 116 948
rect 110 943 111 947
rect 115 943 116 947
rect 502 945 503 949
rect 507 945 508 949
rect 502 944 508 945
rect 686 949 692 950
rect 686 945 687 949
rect 691 945 692 949
rect 686 944 692 945
rect 894 949 900 950
rect 894 945 895 949
rect 899 945 900 949
rect 894 944 900 945
rect 1110 949 1116 950
rect 1110 945 1111 949
rect 1115 945 1116 949
rect 1110 944 1116 945
rect 1342 949 1348 950
rect 1342 945 1343 949
rect 1347 945 1348 949
rect 1342 944 1348 945
rect 1574 949 1580 950
rect 1574 945 1575 949
rect 1579 945 1580 949
rect 1574 944 1580 945
rect 1718 947 1724 948
rect 110 942 116 943
rect 599 943 605 944
rect 599 939 600 943
rect 604 942 605 943
rect 694 943 700 944
rect 694 942 695 943
rect 604 940 695 942
rect 604 939 605 940
rect 599 938 605 939
rect 694 939 695 940
rect 699 939 700 943
rect 694 938 700 939
rect 783 943 789 944
rect 783 939 784 943
rect 788 942 789 943
rect 902 943 908 944
rect 902 942 903 943
rect 788 940 903 942
rect 788 939 789 940
rect 783 938 789 939
rect 902 939 903 940
rect 907 939 908 943
rect 902 938 908 939
rect 991 943 997 944
rect 991 939 992 943
rect 996 942 997 943
rect 1118 943 1124 944
rect 1118 942 1119 943
rect 996 940 1119 942
rect 996 939 997 940
rect 991 938 997 939
rect 1118 939 1119 940
rect 1123 939 1124 943
rect 1118 938 1124 939
rect 1207 943 1213 944
rect 1207 939 1208 943
rect 1212 942 1213 943
rect 1350 943 1356 944
rect 1350 942 1351 943
rect 1212 940 1351 942
rect 1212 939 1213 940
rect 1207 938 1213 939
rect 1350 939 1351 940
rect 1355 939 1356 943
rect 1439 943 1445 944
rect 1439 942 1440 943
rect 1350 938 1356 939
rect 1360 940 1440 942
rect 850 935 856 936
rect 850 931 851 935
rect 855 934 856 935
rect 1360 934 1362 940
rect 1439 939 1440 940
rect 1444 939 1445 943
rect 1439 938 1445 939
rect 1666 943 1677 944
rect 1666 939 1667 943
rect 1671 939 1672 943
rect 1676 939 1677 943
rect 1718 943 1719 947
rect 1723 943 1724 947
rect 1718 942 1724 943
rect 1666 938 1677 939
rect 855 932 1362 934
rect 855 931 856 932
rect 850 930 856 931
rect 1102 923 1108 924
rect 1102 922 1103 923
rect 688 920 1103 922
rect 688 914 690 920
rect 1102 919 1103 920
rect 1107 919 1108 923
rect 1102 918 1108 919
rect 581 912 690 914
rect 694 915 700 916
rect 694 911 695 915
rect 699 911 700 915
rect 694 910 700 911
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 1118 915 1124 916
rect 1118 911 1119 915
rect 1123 911 1124 915
rect 1118 910 1124 911
rect 1350 915 1356 916
rect 1350 911 1351 915
rect 1355 911 1356 915
rect 1350 910 1356 911
rect 1638 915 1644 916
rect 1638 911 1639 915
rect 1643 911 1644 915
rect 1638 910 1644 911
rect 850 859 856 860
rect 850 858 851 859
rect 821 856 851 858
rect 850 855 851 856
rect 855 855 856 859
rect 1666 859 1672 860
rect 1666 858 1667 859
rect 1653 856 1667 858
rect 850 854 856 855
rect 858 855 864 856
rect 858 851 859 855
rect 863 854 864 855
rect 994 855 1000 856
rect 863 852 889 854
rect 863 851 864 852
rect 858 850 864 851
rect 994 851 995 855
rect 999 854 1000 855
rect 1114 855 1120 856
rect 999 852 1025 854
rect 999 851 1000 852
rect 994 850 1000 851
rect 1114 851 1115 855
rect 1119 854 1120 855
rect 1250 855 1256 856
rect 1119 852 1161 854
rect 1119 851 1120 852
rect 1114 850 1120 851
rect 1250 851 1251 855
rect 1255 854 1256 855
rect 1438 855 1444 856
rect 1255 852 1297 854
rect 1255 851 1256 852
rect 1250 850 1256 851
rect 1438 851 1439 855
rect 1443 851 1444 855
rect 1666 855 1667 856
rect 1671 855 1672 859
rect 1666 854 1672 855
rect 1438 850 1444 851
rect 839 829 845 830
rect 110 825 116 826
rect 110 821 111 825
rect 115 821 116 825
rect 839 825 840 829
rect 844 828 845 829
rect 858 829 864 830
rect 858 828 859 829
rect 844 826 859 828
rect 844 825 845 826
rect 839 824 845 825
rect 858 825 859 826
rect 863 825 864 829
rect 858 824 864 825
rect 975 829 981 830
rect 975 825 976 829
rect 980 828 981 829
rect 994 829 1000 830
rect 994 828 995 829
rect 980 826 995 828
rect 980 825 981 826
rect 975 824 981 825
rect 994 825 995 826
rect 999 825 1000 829
rect 994 824 1000 825
rect 1111 829 1120 830
rect 1111 825 1112 829
rect 1119 825 1120 829
rect 1111 824 1120 825
rect 1247 829 1256 830
rect 1247 825 1248 829
rect 1255 825 1256 829
rect 1247 824 1256 825
rect 1382 829 1389 830
rect 1382 825 1383 829
rect 1388 825 1389 829
rect 1382 824 1389 825
rect 1526 829 1533 830
rect 1526 825 1527 829
rect 1532 825 1533 829
rect 1526 824 1533 825
rect 1654 829 1660 830
rect 1654 825 1655 829
rect 1659 828 1660 829
rect 1671 829 1677 830
rect 1671 828 1672 829
rect 1659 826 1672 828
rect 1659 825 1660 826
rect 1654 824 1660 825
rect 1671 825 1672 826
rect 1676 825 1677 829
rect 1671 824 1677 825
rect 1718 825 1724 826
rect 110 820 116 821
rect 742 823 748 824
rect 742 819 743 823
rect 747 819 748 823
rect 742 818 748 819
rect 878 823 884 824
rect 878 819 879 823
rect 883 819 884 823
rect 878 818 884 819
rect 1014 823 1020 824
rect 1014 819 1015 823
rect 1019 819 1020 823
rect 1014 818 1020 819
rect 1150 823 1156 824
rect 1150 819 1151 823
rect 1155 819 1156 823
rect 1150 818 1156 819
rect 1286 823 1292 824
rect 1286 819 1287 823
rect 1291 819 1292 823
rect 1286 818 1292 819
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1574 823 1580 824
rect 1574 819 1575 823
rect 1579 819 1580 823
rect 1718 821 1719 825
rect 1723 821 1724 825
rect 1718 820 1724 821
rect 1574 818 1580 819
rect 766 808 772 809
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 766 804 767 808
rect 771 804 772 808
rect 766 803 772 804
rect 902 808 908 809
rect 902 804 903 808
rect 907 804 908 808
rect 902 803 908 804
rect 1038 808 1044 809
rect 1038 804 1039 808
rect 1043 804 1044 808
rect 1038 803 1044 804
rect 1174 808 1180 809
rect 1174 804 1175 808
rect 1179 804 1180 808
rect 1174 803 1180 804
rect 1310 808 1316 809
rect 1310 804 1311 808
rect 1315 804 1316 808
rect 1310 803 1316 804
rect 1454 808 1460 809
rect 1454 804 1455 808
rect 1459 804 1460 808
rect 1454 803 1460 804
rect 1598 808 1604 809
rect 1598 804 1599 808
rect 1603 804 1604 808
rect 1598 803 1604 804
rect 1718 807 1724 808
rect 1718 803 1719 807
rect 1723 803 1724 807
rect 110 802 116 803
rect 1718 802 1724 803
rect 110 733 116 734
rect 1718 733 1724 734
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 702 732 708 733
rect 702 728 703 732
rect 707 728 708 732
rect 702 727 708 728
rect 862 732 868 733
rect 862 728 863 732
rect 867 728 868 732
rect 862 727 868 728
rect 1030 732 1036 733
rect 1030 728 1031 732
rect 1035 728 1036 732
rect 1030 727 1036 728
rect 1214 732 1220 733
rect 1214 728 1215 732
rect 1219 728 1220 732
rect 1214 727 1220 728
rect 1398 732 1404 733
rect 1398 728 1399 732
rect 1403 728 1404 732
rect 1398 727 1404 728
rect 1590 732 1596 733
rect 1590 728 1591 732
rect 1595 728 1596 732
rect 1718 729 1719 733
rect 1723 729 1724 733
rect 1718 728 1724 729
rect 1590 727 1596 728
rect 678 717 684 718
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 678 713 679 717
rect 683 713 684 717
rect 678 712 684 713
rect 838 717 844 718
rect 838 713 839 717
rect 843 713 844 717
rect 838 712 844 713
rect 1006 717 1012 718
rect 1006 713 1007 717
rect 1011 713 1012 717
rect 1006 712 1012 713
rect 1190 717 1196 718
rect 1190 713 1191 717
rect 1195 713 1196 717
rect 1190 712 1196 713
rect 1374 717 1380 718
rect 1374 713 1375 717
rect 1379 713 1380 717
rect 1374 712 1380 713
rect 1566 717 1572 718
rect 1566 713 1567 717
rect 1571 713 1572 717
rect 1566 712 1572 713
rect 1718 715 1724 716
rect 110 710 116 711
rect 775 711 781 712
rect 775 707 776 711
rect 780 710 781 711
rect 846 711 852 712
rect 846 710 847 711
rect 780 708 847 710
rect 780 707 781 708
rect 775 706 781 707
rect 846 707 847 708
rect 851 707 852 711
rect 846 706 852 707
rect 935 711 941 712
rect 935 707 936 711
rect 940 710 941 711
rect 1014 711 1020 712
rect 1014 710 1015 711
rect 940 708 1015 710
rect 940 707 941 708
rect 935 706 941 707
rect 1014 707 1015 708
rect 1019 707 1020 711
rect 1014 706 1020 707
rect 1102 711 1109 712
rect 1102 707 1103 711
rect 1108 707 1109 711
rect 1287 711 1293 712
rect 1287 710 1288 711
rect 1102 706 1109 707
rect 1159 708 1288 710
rect 754 703 760 704
rect 754 699 755 703
rect 759 702 760 703
rect 1159 702 1161 708
rect 1287 707 1288 708
rect 1292 707 1293 711
rect 1287 706 1293 707
rect 1334 711 1340 712
rect 1334 707 1335 711
rect 1339 710 1340 711
rect 1471 711 1477 712
rect 1471 710 1472 711
rect 1339 708 1472 710
rect 1339 707 1340 708
rect 1334 706 1340 707
rect 1471 707 1472 708
rect 1476 707 1477 711
rect 1471 706 1477 707
rect 1618 711 1624 712
rect 1618 707 1619 711
rect 1623 710 1624 711
rect 1663 711 1669 712
rect 1663 710 1664 711
rect 1623 708 1664 710
rect 1623 707 1624 708
rect 1618 706 1624 707
rect 1663 707 1664 708
rect 1668 707 1669 711
rect 1718 711 1719 715
rect 1723 711 1724 715
rect 1718 710 1724 711
rect 1663 706 1669 707
rect 759 700 1161 702
rect 759 699 760 700
rect 754 698 760 699
rect 754 683 760 684
rect 754 679 755 683
rect 759 679 760 683
rect 754 678 760 679
rect 846 683 852 684
rect 846 679 847 683
rect 851 679 852 683
rect 846 678 852 679
rect 1014 683 1020 684
rect 1014 679 1015 683
rect 1019 679 1020 683
rect 1334 683 1340 684
rect 1334 682 1335 683
rect 1269 680 1335 682
rect 1014 678 1020 679
rect 1334 679 1335 680
rect 1339 679 1340 683
rect 1334 678 1340 679
rect 1382 683 1388 684
rect 1382 679 1383 683
rect 1387 679 1388 683
rect 1654 683 1660 684
rect 1654 682 1655 683
rect 1645 680 1655 682
rect 1382 678 1388 679
rect 1654 679 1655 680
rect 1659 679 1660 683
rect 1654 678 1660 679
rect 407 643 413 644
rect 407 642 408 643
rect 301 640 408 642
rect 407 639 408 640
rect 412 639 413 643
rect 615 643 621 644
rect 615 642 616 643
rect 493 640 616 642
rect 407 638 413 639
rect 615 639 616 640
rect 620 639 621 643
rect 847 643 853 644
rect 847 642 848 643
rect 701 640 848 642
rect 615 638 621 639
rect 847 639 848 640
rect 852 639 853 643
rect 1010 643 1016 644
rect 1010 642 1011 643
rect 933 640 1011 642
rect 847 638 853 639
rect 1010 639 1011 640
rect 1015 639 1016 643
rect 1010 638 1016 639
rect 1102 639 1108 640
rect 1102 635 1103 639
rect 1107 635 1108 639
rect 1102 634 1108 635
rect 1374 639 1380 640
rect 1374 635 1375 639
rect 1379 635 1380 639
rect 1374 634 1380 635
rect 210 615 216 616
rect 210 611 211 615
rect 215 614 216 615
rect 407 615 413 616
rect 215 613 325 614
rect 215 612 320 613
rect 215 611 216 612
rect 210 610 216 611
rect 110 609 116 610
rect 110 605 111 609
rect 115 605 116 609
rect 319 609 320 612
rect 324 609 325 613
rect 407 611 408 615
rect 412 614 413 615
rect 615 615 621 616
rect 412 612 494 614
rect 511 613 517 614
rect 511 612 512 613
rect 412 611 413 612
rect 407 610 413 611
rect 492 610 512 612
rect 319 608 325 609
rect 511 609 512 610
rect 516 609 517 613
rect 615 611 616 615
rect 620 614 621 615
rect 847 615 853 616
rect 620 612 702 614
rect 719 613 725 614
rect 719 612 720 613
rect 620 611 621 612
rect 615 610 621 611
rect 700 610 720 612
rect 511 608 517 609
rect 719 609 720 610
rect 724 609 725 613
rect 847 611 848 615
rect 852 614 853 615
rect 1010 615 1016 616
rect 852 612 934 614
rect 951 613 957 614
rect 951 612 952 613
rect 852 611 853 612
rect 847 610 853 611
rect 932 610 952 612
rect 719 608 725 609
rect 951 609 952 610
rect 956 609 957 613
rect 1010 611 1011 615
rect 1015 614 1016 615
rect 1015 612 1178 614
rect 1191 613 1197 614
rect 1191 612 1192 613
rect 1015 611 1016 612
rect 1010 610 1016 611
rect 1176 610 1192 612
rect 951 608 957 609
rect 1191 609 1192 610
rect 1196 609 1197 613
rect 1191 608 1197 609
rect 1431 613 1437 614
rect 1431 609 1432 613
rect 1436 609 1437 613
rect 1431 608 1437 609
rect 1718 609 1724 610
rect 110 604 116 605
rect 222 607 228 608
rect 222 603 223 607
rect 227 603 228 607
rect 222 602 228 603
rect 414 607 420 608
rect 414 603 415 607
rect 419 603 420 607
rect 414 602 420 603
rect 622 607 628 608
rect 622 603 623 607
rect 627 603 628 607
rect 622 602 628 603
rect 854 607 860 608
rect 854 603 855 607
rect 859 603 860 607
rect 854 602 860 603
rect 1094 607 1100 608
rect 1094 603 1095 607
rect 1099 603 1100 607
rect 1094 602 1100 603
rect 1334 607 1340 608
rect 1334 603 1335 607
rect 1339 603 1340 607
rect 1718 605 1719 609
rect 1723 605 1724 609
rect 1718 604 1724 605
rect 1334 602 1340 603
rect 246 592 252 593
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 246 588 247 592
rect 251 588 252 592
rect 246 587 252 588
rect 438 592 444 593
rect 438 588 439 592
rect 443 588 444 592
rect 438 587 444 588
rect 646 592 652 593
rect 646 588 647 592
rect 651 588 652 592
rect 646 587 652 588
rect 878 592 884 593
rect 878 588 879 592
rect 883 588 884 592
rect 878 587 884 588
rect 1118 592 1124 593
rect 1118 588 1119 592
rect 1123 588 1124 592
rect 1118 587 1124 588
rect 1358 592 1364 593
rect 1358 588 1359 592
rect 1363 588 1364 592
rect 1358 587 1364 588
rect 1718 591 1724 592
rect 1718 587 1719 591
rect 1723 587 1724 591
rect 110 586 116 587
rect 1718 586 1724 587
rect 110 521 116 522
rect 1718 521 1724 522
rect 110 517 111 521
rect 115 517 116 521
rect 110 516 116 517
rect 158 520 164 521
rect 158 516 159 520
rect 163 516 164 520
rect 158 515 164 516
rect 326 520 332 521
rect 326 516 327 520
rect 331 516 332 520
rect 326 515 332 516
rect 542 520 548 521
rect 542 516 543 520
rect 547 516 548 520
rect 542 515 548 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 1038 520 1044 521
rect 1038 516 1039 520
rect 1043 516 1044 520
rect 1038 515 1044 516
rect 1302 520 1308 521
rect 1302 516 1303 520
rect 1307 516 1308 520
rect 1302 515 1308 516
rect 1566 520 1572 521
rect 1566 516 1567 520
rect 1571 516 1572 520
rect 1718 517 1719 521
rect 1723 517 1724 521
rect 1718 516 1724 517
rect 1566 515 1572 516
rect 134 505 140 506
rect 110 503 116 504
rect 110 499 111 503
rect 115 499 116 503
rect 134 501 135 505
rect 139 501 140 505
rect 134 500 140 501
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 518 505 524 506
rect 518 501 519 505
rect 523 501 524 505
rect 518 500 524 501
rect 758 505 764 506
rect 758 501 759 505
rect 763 501 764 505
rect 758 500 764 501
rect 1014 505 1020 506
rect 1014 501 1015 505
rect 1019 501 1020 505
rect 1014 500 1020 501
rect 1278 505 1284 506
rect 1278 501 1279 505
rect 1283 501 1284 505
rect 1278 500 1284 501
rect 1542 505 1548 506
rect 1542 501 1543 505
rect 1547 501 1548 505
rect 1542 500 1548 501
rect 1718 503 1724 504
rect 110 498 116 499
rect 231 499 237 500
rect 231 495 232 499
rect 236 498 237 499
rect 310 499 316 500
rect 310 498 311 499
rect 236 496 311 498
rect 236 495 237 496
rect 231 494 237 495
rect 310 495 311 496
rect 315 495 316 499
rect 310 494 316 495
rect 399 499 405 500
rect 399 495 400 499
rect 404 498 405 499
rect 526 499 532 500
rect 526 498 527 499
rect 404 496 527 498
rect 404 495 405 496
rect 399 494 405 495
rect 526 495 527 496
rect 531 495 532 499
rect 526 494 532 495
rect 615 499 621 500
rect 615 495 616 499
rect 620 498 621 499
rect 766 499 772 500
rect 766 498 767 499
rect 620 496 767 498
rect 620 495 621 496
rect 615 494 621 495
rect 766 495 767 496
rect 771 495 772 499
rect 766 494 772 495
rect 855 499 861 500
rect 855 495 856 499
rect 860 498 861 499
rect 1022 499 1028 500
rect 1022 498 1023 499
rect 860 496 1023 498
rect 860 495 861 496
rect 855 494 861 495
rect 1022 495 1023 496
rect 1027 495 1028 499
rect 1111 499 1117 500
rect 1111 498 1112 499
rect 1022 494 1028 495
rect 1040 496 1112 498
rect 290 491 296 492
rect 290 487 291 491
rect 295 490 296 491
rect 1040 490 1042 496
rect 1111 495 1112 496
rect 1116 495 1117 499
rect 1111 494 1117 495
rect 1374 499 1381 500
rect 1374 495 1375 499
rect 1380 495 1381 499
rect 1374 494 1381 495
rect 1634 499 1645 500
rect 1634 495 1635 499
rect 1639 495 1640 499
rect 1644 495 1645 499
rect 1718 499 1719 503
rect 1723 499 1724 503
rect 1718 498 1724 499
rect 1634 494 1645 495
rect 295 488 1042 490
rect 295 487 296 488
rect 290 486 296 487
rect 210 471 216 472
rect 210 467 211 471
rect 215 467 216 471
rect 210 466 216 467
rect 310 471 316 472
rect 310 467 311 471
rect 315 467 316 471
rect 310 466 316 467
rect 526 471 532 472
rect 526 467 527 471
rect 531 467 532 471
rect 526 466 532 467
rect 766 471 772 472
rect 766 467 767 471
rect 771 467 772 471
rect 766 466 772 467
rect 1022 471 1028 472
rect 1022 467 1023 471
rect 1027 467 1028 471
rect 1414 471 1420 472
rect 1414 470 1415 471
rect 1357 468 1415 470
rect 1022 466 1028 467
rect 1414 467 1415 468
rect 1419 467 1420 471
rect 1414 466 1420 467
rect 1618 471 1624 472
rect 1618 467 1619 471
rect 1623 467 1624 471
rect 1618 466 1624 467
rect 290 415 296 416
rect 290 414 291 415
rect 277 412 291 414
rect 290 411 291 412
rect 295 411 296 415
rect 290 410 296 411
rect 298 411 304 412
rect 298 407 299 411
rect 303 410 304 411
rect 546 411 552 412
rect 303 408 441 410
rect 303 407 304 408
rect 298 406 304 407
rect 546 407 547 411
rect 551 410 552 411
rect 1002 411 1008 412
rect 551 408 673 410
rect 551 407 552 408
rect 546 406 552 407
rect 960 402 962 409
rect 1002 407 1003 411
rect 1007 410 1008 411
rect 1226 411 1232 412
rect 1007 408 1121 410
rect 1007 407 1008 408
rect 1002 406 1008 407
rect 1226 407 1227 411
rect 1231 410 1232 411
rect 1634 411 1640 412
rect 1231 408 1345 410
rect 1231 407 1232 408
rect 1226 406 1232 407
rect 1634 407 1635 411
rect 1639 407 1640 411
rect 1634 406 1640 407
rect 1190 403 1196 404
rect 1190 402 1191 403
rect 960 400 1191 402
rect 1190 399 1191 400
rect 1195 399 1196 403
rect 1190 398 1196 399
rect 295 385 304 386
rect 110 381 116 382
rect 110 377 111 381
rect 115 377 116 381
rect 295 381 296 385
rect 303 381 304 385
rect 295 380 304 381
rect 527 385 533 386
rect 527 381 528 385
rect 532 384 533 385
rect 546 385 552 386
rect 546 384 547 385
rect 532 382 547 384
rect 532 381 533 382
rect 527 380 533 381
rect 546 381 547 382
rect 551 381 552 385
rect 546 380 552 381
rect 759 385 768 386
rect 759 381 760 385
rect 767 381 768 385
rect 759 380 768 381
rect 983 385 989 386
rect 983 381 984 385
rect 988 384 989 385
rect 1002 385 1008 386
rect 1002 384 1003 385
rect 988 382 1003 384
rect 988 381 989 382
rect 983 380 989 381
rect 1002 381 1003 382
rect 1007 381 1008 385
rect 1002 380 1008 381
rect 1207 385 1213 386
rect 1207 381 1208 385
rect 1212 384 1213 385
rect 1226 385 1232 386
rect 1226 384 1227 385
rect 1212 382 1227 384
rect 1212 381 1213 382
rect 1207 380 1213 381
rect 1226 381 1227 382
rect 1231 381 1232 385
rect 1226 380 1232 381
rect 1414 385 1420 386
rect 1414 381 1415 385
rect 1419 384 1420 385
rect 1431 385 1437 386
rect 1431 384 1432 385
rect 1419 382 1432 384
rect 1419 381 1420 382
rect 1414 380 1420 381
rect 1431 381 1432 382
rect 1436 381 1437 385
rect 1431 380 1437 381
rect 1650 385 1661 386
rect 1650 381 1651 385
rect 1655 381 1656 385
rect 1660 381 1661 385
rect 1650 380 1661 381
rect 1718 381 1724 382
rect 110 376 116 377
rect 198 379 204 380
rect 198 375 199 379
rect 203 375 204 379
rect 198 374 204 375
rect 430 379 436 380
rect 430 375 431 379
rect 435 375 436 379
rect 430 374 436 375
rect 662 379 668 380
rect 662 375 663 379
rect 667 375 668 379
rect 662 374 668 375
rect 886 379 892 380
rect 886 375 887 379
rect 891 375 892 379
rect 886 374 892 375
rect 1110 379 1116 380
rect 1110 375 1111 379
rect 1115 375 1116 379
rect 1110 374 1116 375
rect 1334 379 1340 380
rect 1334 375 1335 379
rect 1339 375 1340 379
rect 1334 374 1340 375
rect 1558 379 1564 380
rect 1558 375 1559 379
rect 1563 375 1564 379
rect 1718 377 1719 381
rect 1723 377 1724 381
rect 1718 376 1724 377
rect 1558 374 1564 375
rect 222 364 228 365
rect 110 363 116 364
rect 110 359 111 363
rect 115 359 116 363
rect 222 360 223 364
rect 227 360 228 364
rect 222 359 228 360
rect 454 364 460 365
rect 454 360 455 364
rect 459 360 460 364
rect 454 359 460 360
rect 686 364 692 365
rect 686 360 687 364
rect 691 360 692 364
rect 686 359 692 360
rect 910 364 916 365
rect 910 360 911 364
rect 915 360 916 364
rect 910 359 916 360
rect 1134 364 1140 365
rect 1134 360 1135 364
rect 1139 360 1140 364
rect 1134 359 1140 360
rect 1358 364 1364 365
rect 1358 360 1359 364
rect 1363 360 1364 364
rect 1358 359 1364 360
rect 1582 364 1588 365
rect 1582 360 1583 364
rect 1587 360 1588 364
rect 1582 359 1588 360
rect 1718 363 1724 364
rect 1718 359 1719 363
rect 1723 359 1724 363
rect 110 358 116 359
rect 1718 358 1724 359
rect 110 293 116 294
rect 1718 293 1724 294
rect 110 289 111 293
rect 115 289 116 293
rect 110 288 116 289
rect 438 292 444 293
rect 438 288 439 292
rect 443 288 444 292
rect 438 287 444 288
rect 654 292 660 293
rect 654 288 655 292
rect 659 288 660 292
rect 654 287 660 288
rect 878 292 884 293
rect 878 288 879 292
rect 883 288 884 292
rect 878 287 884 288
rect 1118 292 1124 293
rect 1118 288 1119 292
rect 1123 288 1124 292
rect 1118 287 1124 288
rect 1366 292 1372 293
rect 1366 288 1367 292
rect 1371 288 1372 292
rect 1366 287 1372 288
rect 1598 292 1604 293
rect 1598 288 1599 292
rect 1603 288 1604 292
rect 1718 289 1719 293
rect 1723 289 1724 293
rect 1718 288 1724 289
rect 1598 287 1604 288
rect 414 277 420 278
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 414 273 415 277
rect 419 273 420 277
rect 414 272 420 273
rect 630 277 636 278
rect 630 273 631 277
rect 635 273 636 277
rect 630 272 636 273
rect 854 277 860 278
rect 854 273 855 277
rect 859 273 860 277
rect 854 272 860 273
rect 1094 277 1100 278
rect 1094 273 1095 277
rect 1099 273 1100 277
rect 1094 272 1100 273
rect 1342 277 1348 278
rect 1342 273 1343 277
rect 1347 273 1348 277
rect 1342 272 1348 273
rect 1574 277 1580 278
rect 1574 273 1575 277
rect 1579 273 1580 277
rect 1574 272 1580 273
rect 1718 275 1724 276
rect 110 270 116 271
rect 510 271 517 272
rect 510 267 511 271
rect 516 267 517 271
rect 510 266 517 267
rect 574 271 580 272
rect 574 267 575 271
rect 579 270 580 271
rect 727 271 733 272
rect 727 270 728 271
rect 579 268 728 270
rect 579 267 580 268
rect 574 266 580 267
rect 727 267 728 268
rect 732 267 733 271
rect 727 266 733 267
rect 754 271 760 272
rect 754 267 755 271
rect 759 270 760 271
rect 951 271 957 272
rect 951 270 952 271
rect 759 268 952 270
rect 759 267 760 268
rect 754 266 760 267
rect 951 267 952 268
rect 956 267 957 271
rect 951 266 957 267
rect 1190 271 1197 272
rect 1190 267 1191 271
rect 1196 267 1197 271
rect 1190 266 1197 267
rect 1298 271 1304 272
rect 1298 267 1299 271
rect 1303 270 1304 271
rect 1439 271 1445 272
rect 1439 270 1440 271
rect 1303 268 1440 270
rect 1303 267 1304 268
rect 1298 266 1304 267
rect 1439 267 1440 268
rect 1444 267 1445 271
rect 1439 266 1445 267
rect 1666 271 1677 272
rect 1666 267 1667 271
rect 1671 267 1672 271
rect 1676 267 1677 271
rect 1718 271 1719 275
rect 1723 271 1724 275
rect 1718 270 1724 271
rect 1666 266 1677 267
rect 574 243 580 244
rect 574 242 575 243
rect 493 240 575 242
rect 574 239 575 240
rect 579 239 580 243
rect 754 243 760 244
rect 754 242 755 243
rect 709 240 755 242
rect 574 238 580 239
rect 754 239 755 240
rect 759 239 760 243
rect 754 238 760 239
rect 762 243 768 244
rect 762 239 763 243
rect 767 242 768 243
rect 1298 243 1304 244
rect 1298 242 1299 243
rect 767 240 865 242
rect 1173 240 1299 242
rect 767 239 768 240
rect 762 238 768 239
rect 1298 239 1299 240
rect 1303 239 1304 243
rect 1298 238 1304 239
rect 1398 243 1404 244
rect 1398 239 1399 243
rect 1403 239 1404 243
rect 1398 238 1404 239
rect 1650 243 1656 244
rect 1650 239 1651 243
rect 1655 239 1656 243
rect 1650 238 1656 239
rect 1666 191 1672 192
rect 1666 190 1667 191
rect 1653 188 1667 190
rect 510 187 516 188
rect 510 183 511 187
rect 515 183 516 187
rect 510 182 516 183
rect 602 187 608 188
rect 602 183 603 187
rect 607 186 608 187
rect 738 187 744 188
rect 607 184 633 186
rect 607 183 608 184
rect 602 182 608 183
rect 738 183 739 187
rect 743 186 744 187
rect 874 187 880 188
rect 743 184 769 186
rect 743 183 744 184
rect 738 182 744 183
rect 874 183 875 187
rect 879 186 880 187
rect 1010 187 1016 188
rect 879 184 905 186
rect 879 183 880 184
rect 874 182 880 183
rect 1010 183 1011 187
rect 1015 186 1016 187
rect 1146 187 1152 188
rect 1015 184 1041 186
rect 1015 183 1016 184
rect 1010 182 1016 183
rect 1146 183 1147 187
rect 1151 186 1152 187
rect 1266 187 1272 188
rect 1151 184 1177 186
rect 1151 183 1152 184
rect 1146 182 1152 183
rect 1266 183 1267 187
rect 1271 186 1272 187
rect 1514 187 1520 188
rect 1271 184 1313 186
rect 1271 183 1272 184
rect 1266 182 1272 183
rect 1514 183 1515 187
rect 1519 183 1520 187
rect 1666 187 1667 188
rect 1671 187 1672 191
rect 1666 186 1672 187
rect 1514 182 1520 183
rect 1514 163 1520 164
rect 583 161 589 162
rect 110 157 116 158
rect 110 153 111 157
rect 115 153 116 157
rect 583 157 584 161
rect 588 160 589 161
rect 602 161 608 162
rect 602 160 603 161
rect 588 158 603 160
rect 588 157 589 158
rect 583 156 589 157
rect 602 157 603 158
rect 607 157 608 161
rect 602 156 608 157
rect 719 161 725 162
rect 719 157 720 161
rect 724 160 725 161
rect 738 161 744 162
rect 738 160 739 161
rect 724 158 739 160
rect 724 157 725 158
rect 719 156 725 157
rect 738 157 739 158
rect 743 157 744 161
rect 738 156 744 157
rect 855 161 861 162
rect 855 157 856 161
rect 860 160 861 161
rect 874 161 880 162
rect 874 160 875 161
rect 860 158 875 160
rect 860 157 861 158
rect 855 156 861 157
rect 874 157 875 158
rect 879 157 880 161
rect 874 156 880 157
rect 991 161 997 162
rect 991 157 992 161
rect 996 160 997 161
rect 1010 161 1016 162
rect 1010 160 1011 161
rect 996 158 1011 160
rect 996 157 997 158
rect 991 156 997 157
rect 1010 157 1011 158
rect 1015 157 1016 161
rect 1010 156 1016 157
rect 1127 161 1133 162
rect 1127 157 1128 161
rect 1132 160 1133 161
rect 1146 161 1152 162
rect 1146 160 1147 161
rect 1132 158 1147 160
rect 1132 157 1133 158
rect 1127 156 1133 157
rect 1146 157 1147 158
rect 1151 157 1152 161
rect 1146 156 1152 157
rect 1263 161 1272 162
rect 1263 157 1264 161
rect 1271 157 1272 161
rect 1263 156 1272 157
rect 1398 161 1405 162
rect 1398 157 1399 161
rect 1404 157 1405 161
rect 1514 159 1515 163
rect 1519 162 1520 163
rect 1519 160 1654 162
rect 1671 161 1677 162
rect 1671 160 1672 161
rect 1519 159 1520 160
rect 1514 158 1520 159
rect 1652 158 1672 160
rect 1398 156 1405 157
rect 1671 157 1672 158
rect 1676 157 1677 161
rect 1671 156 1677 157
rect 1718 157 1724 158
rect 110 152 116 153
rect 486 155 492 156
rect 486 151 487 155
rect 491 151 492 155
rect 486 150 492 151
rect 622 155 628 156
rect 622 151 623 155
rect 627 151 628 155
rect 622 150 628 151
rect 758 155 764 156
rect 758 151 759 155
rect 763 151 764 155
rect 758 150 764 151
rect 894 155 900 156
rect 894 151 895 155
rect 899 151 900 155
rect 894 150 900 151
rect 1030 155 1036 156
rect 1030 151 1031 155
rect 1035 151 1036 155
rect 1030 150 1036 151
rect 1166 155 1172 156
rect 1166 151 1167 155
rect 1171 151 1172 155
rect 1166 150 1172 151
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1302 150 1308 151
rect 1438 155 1444 156
rect 1438 151 1439 155
rect 1443 151 1444 155
rect 1438 150 1444 151
rect 1574 155 1580 156
rect 1574 151 1575 155
rect 1579 151 1580 155
rect 1718 153 1719 157
rect 1723 153 1724 157
rect 1718 152 1724 153
rect 1574 150 1580 151
rect 510 140 516 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 510 136 511 140
rect 515 136 516 140
rect 510 135 516 136
rect 646 140 652 141
rect 646 136 647 140
rect 651 136 652 140
rect 646 135 652 136
rect 782 140 788 141
rect 782 136 783 140
rect 787 136 788 140
rect 782 135 788 136
rect 918 140 924 141
rect 918 136 919 140
rect 923 136 924 140
rect 918 135 924 136
rect 1054 140 1060 141
rect 1054 136 1055 140
rect 1059 136 1060 140
rect 1054 135 1060 136
rect 1190 140 1196 141
rect 1190 136 1191 140
rect 1195 136 1196 140
rect 1190 135 1196 136
rect 1326 140 1332 141
rect 1326 136 1327 140
rect 1331 136 1332 140
rect 1326 135 1332 136
rect 1462 140 1468 141
rect 1462 136 1463 140
rect 1467 136 1468 140
rect 1462 135 1468 136
rect 1598 140 1604 141
rect 1598 136 1599 140
rect 1603 136 1604 140
rect 1598 135 1604 136
rect 1718 139 1724 140
rect 1718 135 1719 139
rect 1723 135 1724 139
rect 110 134 116 135
rect 1718 134 1724 135
<< m3c >>
rect 247 1755 251 1759
rect 387 1755 391 1759
rect 523 1755 527 1759
rect 659 1755 663 1759
rect 111 1725 115 1729
rect 247 1729 251 1733
rect 387 1729 391 1733
rect 523 1729 527 1733
rect 659 1729 663 1733
rect 767 1729 771 1733
rect 135 1723 139 1727
rect 271 1723 275 1727
rect 407 1723 411 1727
rect 543 1723 547 1727
rect 679 1723 683 1727
rect 1719 1725 1723 1729
rect 111 1707 115 1711
rect 159 1708 163 1712
rect 295 1708 299 1712
rect 431 1708 435 1712
rect 567 1708 571 1712
rect 703 1708 707 1712
rect 1719 1707 1723 1711
rect 111 1637 115 1641
rect 231 1636 235 1640
rect 367 1636 371 1640
rect 503 1636 507 1640
rect 639 1636 643 1640
rect 775 1636 779 1640
rect 1719 1637 1723 1641
rect 111 1619 115 1623
rect 207 1621 211 1625
rect 343 1621 347 1625
rect 479 1621 483 1625
rect 615 1621 619 1625
rect 751 1621 755 1625
rect 351 1615 355 1619
rect 487 1615 491 1619
rect 623 1615 627 1619
rect 759 1615 763 1619
rect 595 1607 599 1611
rect 1719 1619 1723 1623
rect 767 1595 771 1599
rect 351 1587 355 1591
rect 487 1587 491 1591
rect 623 1587 627 1591
rect 759 1587 763 1591
rect 595 1535 599 1539
rect 603 1531 607 1535
rect 739 1531 743 1535
rect 875 1531 879 1535
rect 1011 1531 1015 1535
rect 1275 1535 1279 1539
rect 1283 1531 1287 1535
rect 1419 1531 1423 1535
rect 1555 1531 1559 1535
rect 111 1501 115 1505
rect 603 1505 607 1509
rect 739 1505 743 1509
rect 875 1505 879 1509
rect 1011 1505 1015 1509
rect 1111 1505 1115 1509
rect 1283 1505 1287 1509
rect 1419 1505 1423 1509
rect 1555 1505 1559 1509
rect 487 1499 491 1503
rect 623 1499 627 1503
rect 759 1499 763 1503
rect 895 1499 899 1503
rect 1031 1499 1035 1503
rect 1167 1499 1171 1503
rect 1303 1499 1307 1503
rect 1439 1499 1443 1503
rect 1575 1499 1579 1503
rect 1719 1501 1723 1505
rect 111 1483 115 1487
rect 511 1484 515 1488
rect 647 1484 651 1488
rect 783 1484 787 1488
rect 919 1484 923 1488
rect 1055 1484 1059 1488
rect 1191 1484 1195 1488
rect 1327 1484 1331 1488
rect 1463 1484 1467 1488
rect 1599 1484 1603 1488
rect 1719 1483 1723 1487
rect 111 1409 115 1413
rect 623 1408 627 1412
rect 759 1408 763 1412
rect 895 1408 899 1412
rect 1039 1408 1043 1412
rect 1183 1408 1187 1412
rect 1327 1408 1331 1412
rect 1463 1408 1467 1412
rect 1599 1408 1603 1412
rect 1719 1409 1723 1413
rect 111 1391 115 1395
rect 599 1393 603 1397
rect 735 1393 739 1397
rect 871 1393 875 1397
rect 1015 1393 1019 1397
rect 1159 1393 1163 1397
rect 1303 1393 1307 1397
rect 1439 1393 1443 1397
rect 1575 1393 1579 1397
rect 743 1387 747 1391
rect 879 1387 883 1391
rect 971 1387 972 1391
rect 972 1387 975 1391
rect 675 1379 679 1383
rect 1255 1387 1256 1391
rect 1256 1387 1259 1391
rect 1279 1387 1283 1391
rect 1535 1387 1536 1391
rect 1536 1387 1539 1391
rect 1559 1387 1563 1391
rect 1719 1391 1723 1395
rect 971 1367 975 1371
rect 675 1359 679 1363
rect 743 1359 747 1363
rect 879 1359 883 1363
rect 1111 1359 1115 1363
rect 1359 1359 1363 1363
rect 1559 1359 1563 1363
rect 527 1303 531 1307
rect 887 1303 891 1307
rect 1199 1303 1203 1307
rect 1255 1299 1259 1303
rect 1535 1299 1539 1303
rect 111 1269 115 1273
rect 527 1275 531 1279
rect 887 1275 891 1279
rect 1199 1275 1203 1279
rect 1603 1273 1607 1277
rect 135 1267 139 1271
rect 343 1267 347 1271
rect 607 1267 611 1271
rect 895 1267 899 1271
rect 1207 1267 1211 1271
rect 1519 1267 1523 1271
rect 1719 1269 1723 1273
rect 111 1251 115 1255
rect 159 1252 163 1256
rect 367 1252 371 1256
rect 631 1252 635 1256
rect 919 1252 923 1256
rect 1231 1252 1235 1256
rect 1543 1252 1547 1256
rect 1719 1251 1723 1255
rect 111 1181 115 1185
rect 159 1180 163 1184
rect 327 1180 331 1184
rect 543 1180 547 1184
rect 775 1180 779 1184
rect 1023 1180 1027 1184
rect 1287 1180 1291 1184
rect 1551 1180 1555 1184
rect 1719 1181 1723 1185
rect 111 1163 115 1167
rect 135 1165 139 1169
rect 303 1165 307 1169
rect 519 1165 523 1169
rect 751 1165 755 1169
rect 999 1165 1003 1169
rect 1263 1165 1267 1169
rect 1527 1165 1531 1169
rect 311 1159 315 1163
rect 527 1159 531 1163
rect 759 1159 763 1163
rect 1007 1159 1011 1163
rect 419 1147 423 1151
rect 1359 1159 1360 1163
rect 1360 1159 1363 1163
rect 1619 1159 1623 1163
rect 1719 1163 1723 1167
rect 311 1131 315 1135
rect 527 1131 531 1135
rect 759 1131 763 1135
rect 1007 1131 1011 1135
rect 1359 1131 1363 1135
rect 1603 1131 1607 1135
rect 419 1071 423 1075
rect 427 1067 431 1071
rect 651 1067 655 1071
rect 891 1067 895 1071
rect 1527 1071 1531 1075
rect 1619 1067 1623 1071
rect 111 1037 115 1041
rect 427 1041 431 1045
rect 651 1041 655 1045
rect 891 1041 895 1045
rect 1103 1041 1107 1045
rect 1359 1041 1363 1045
rect 1639 1041 1640 1045
rect 1640 1041 1643 1045
rect 311 1035 315 1039
rect 535 1035 539 1039
rect 775 1035 779 1039
rect 1023 1035 1027 1039
rect 1279 1035 1283 1039
rect 1543 1035 1547 1039
rect 1719 1037 1723 1041
rect 111 1019 115 1023
rect 335 1020 339 1024
rect 559 1020 563 1024
rect 799 1020 803 1024
rect 1047 1020 1051 1024
rect 1303 1020 1307 1024
rect 1567 1020 1571 1024
rect 1719 1019 1723 1023
rect 111 961 115 965
rect 527 960 531 964
rect 711 960 715 964
rect 919 960 923 964
rect 1135 960 1139 964
rect 1367 960 1371 964
rect 1599 960 1603 964
rect 1719 961 1723 965
rect 111 943 115 947
rect 503 945 507 949
rect 687 945 691 949
rect 895 945 899 949
rect 1111 945 1115 949
rect 1343 945 1347 949
rect 1575 945 1579 949
rect 695 939 699 943
rect 903 939 907 943
rect 1119 939 1123 943
rect 1351 939 1355 943
rect 851 931 855 935
rect 1667 939 1671 943
rect 1719 943 1723 947
rect 1103 919 1107 923
rect 695 911 699 915
rect 903 911 907 915
rect 1119 911 1123 915
rect 1351 911 1355 915
rect 1639 911 1643 915
rect 851 855 855 859
rect 859 851 863 855
rect 995 851 999 855
rect 1115 851 1119 855
rect 1251 851 1255 855
rect 1439 851 1443 855
rect 1667 855 1671 859
rect 111 821 115 825
rect 859 825 863 829
rect 995 825 999 829
rect 1115 825 1116 829
rect 1116 825 1119 829
rect 1251 825 1252 829
rect 1252 825 1255 829
rect 1383 825 1384 829
rect 1384 825 1387 829
rect 1527 825 1528 829
rect 1528 825 1531 829
rect 1655 825 1659 829
rect 743 819 747 823
rect 879 819 883 823
rect 1015 819 1019 823
rect 1151 819 1155 823
rect 1287 819 1291 823
rect 1431 819 1435 823
rect 1575 819 1579 823
rect 1719 821 1723 825
rect 111 803 115 807
rect 767 804 771 808
rect 903 804 907 808
rect 1039 804 1043 808
rect 1175 804 1179 808
rect 1311 804 1315 808
rect 1455 804 1459 808
rect 1599 804 1603 808
rect 1719 803 1723 807
rect 111 729 115 733
rect 703 728 707 732
rect 863 728 867 732
rect 1031 728 1035 732
rect 1215 728 1219 732
rect 1399 728 1403 732
rect 1591 728 1595 732
rect 1719 729 1723 733
rect 111 711 115 715
rect 679 713 683 717
rect 839 713 843 717
rect 1007 713 1011 717
rect 1191 713 1195 717
rect 1375 713 1379 717
rect 1567 713 1571 717
rect 847 707 851 711
rect 1015 707 1019 711
rect 1103 707 1104 711
rect 1104 707 1107 711
rect 755 699 759 703
rect 1335 707 1339 711
rect 1619 707 1623 711
rect 1719 711 1723 715
rect 755 679 759 683
rect 847 679 851 683
rect 1015 679 1019 683
rect 1335 679 1339 683
rect 1383 679 1387 683
rect 1655 679 1659 683
rect 1011 639 1015 643
rect 1103 635 1107 639
rect 1375 635 1379 639
rect 211 611 215 615
rect 111 605 115 609
rect 1011 611 1015 615
rect 1432 609 1436 613
rect 223 603 227 607
rect 415 603 419 607
rect 623 603 627 607
rect 855 603 859 607
rect 1095 603 1099 607
rect 1335 603 1339 607
rect 1719 605 1723 609
rect 111 587 115 591
rect 247 588 251 592
rect 439 588 443 592
rect 647 588 651 592
rect 879 588 883 592
rect 1119 588 1123 592
rect 1359 588 1363 592
rect 1719 587 1723 591
rect 111 517 115 521
rect 159 516 163 520
rect 327 516 331 520
rect 543 516 547 520
rect 783 516 787 520
rect 1039 516 1043 520
rect 1303 516 1307 520
rect 1567 516 1571 520
rect 1719 517 1723 521
rect 111 499 115 503
rect 135 501 139 505
rect 303 501 307 505
rect 519 501 523 505
rect 759 501 763 505
rect 1015 501 1019 505
rect 1279 501 1283 505
rect 1543 501 1547 505
rect 311 495 315 499
rect 527 495 531 499
rect 767 495 771 499
rect 1023 495 1027 499
rect 291 487 295 491
rect 1375 495 1376 499
rect 1376 495 1379 499
rect 1635 495 1639 499
rect 1719 499 1723 503
rect 211 467 215 471
rect 311 467 315 471
rect 527 467 531 471
rect 767 467 771 471
rect 1023 467 1027 471
rect 1415 467 1419 471
rect 1619 467 1623 471
rect 291 411 295 415
rect 299 407 303 411
rect 547 407 551 411
rect 1003 407 1007 411
rect 1227 407 1231 411
rect 1635 407 1639 411
rect 1191 399 1195 403
rect 111 377 115 381
rect 299 381 300 385
rect 300 381 303 385
rect 547 381 551 385
rect 763 381 764 385
rect 764 381 767 385
rect 1003 381 1007 385
rect 1227 381 1231 385
rect 1415 381 1419 385
rect 1651 381 1655 385
rect 199 375 203 379
rect 431 375 435 379
rect 663 375 667 379
rect 887 375 891 379
rect 1111 375 1115 379
rect 1335 375 1339 379
rect 1559 375 1563 379
rect 1719 377 1723 381
rect 111 359 115 363
rect 223 360 227 364
rect 455 360 459 364
rect 687 360 691 364
rect 911 360 915 364
rect 1135 360 1139 364
rect 1359 360 1363 364
rect 1583 360 1587 364
rect 1719 359 1723 363
rect 111 289 115 293
rect 439 288 443 292
rect 655 288 659 292
rect 879 288 883 292
rect 1119 288 1123 292
rect 1367 288 1371 292
rect 1599 288 1603 292
rect 1719 289 1723 293
rect 111 271 115 275
rect 415 273 419 277
rect 631 273 635 277
rect 855 273 859 277
rect 1095 273 1099 277
rect 1343 273 1347 277
rect 1575 273 1579 277
rect 511 267 512 271
rect 512 267 515 271
rect 575 267 579 271
rect 755 267 759 271
rect 1191 267 1192 271
rect 1192 267 1195 271
rect 1299 267 1303 271
rect 1667 267 1671 271
rect 1719 271 1723 275
rect 575 239 579 243
rect 755 239 759 243
rect 763 239 767 243
rect 1299 239 1303 243
rect 1399 239 1403 243
rect 1651 239 1655 243
rect 511 183 515 187
rect 603 183 607 187
rect 739 183 743 187
rect 875 183 879 187
rect 1011 183 1015 187
rect 1147 183 1151 187
rect 1267 183 1271 187
rect 1515 183 1519 187
rect 1667 187 1671 191
rect 111 153 115 157
rect 603 157 607 161
rect 739 157 743 161
rect 875 157 879 161
rect 1011 157 1015 161
rect 1147 157 1151 161
rect 1267 157 1268 161
rect 1268 157 1271 161
rect 1399 157 1400 161
rect 1400 157 1403 161
rect 1515 159 1519 163
rect 487 151 491 155
rect 623 151 627 155
rect 759 151 763 155
rect 895 151 899 155
rect 1031 151 1035 155
rect 1167 151 1171 155
rect 1303 151 1307 155
rect 1439 151 1443 155
rect 1575 151 1579 155
rect 1719 153 1723 157
rect 111 135 115 139
rect 511 136 515 140
rect 647 136 651 140
rect 783 136 787 140
rect 919 136 923 140
rect 1055 136 1059 140
rect 1191 136 1195 140
rect 1327 136 1331 140
rect 1463 136 1467 140
rect 1599 136 1603 140
rect 1719 135 1723 139
<< m3 >>
rect 111 1782 115 1783
rect 111 1777 115 1778
rect 135 1782 139 1783
rect 135 1777 139 1778
rect 271 1782 275 1783
rect 271 1777 275 1778
rect 407 1782 411 1783
rect 407 1777 411 1778
rect 543 1782 547 1783
rect 543 1777 547 1778
rect 679 1782 683 1783
rect 679 1777 683 1778
rect 1719 1782 1723 1783
rect 1719 1777 1723 1778
rect 112 1730 114 1777
rect 110 1729 116 1730
rect 110 1725 111 1729
rect 115 1725 116 1729
rect 136 1728 138 1777
rect 246 1759 252 1760
rect 246 1755 247 1759
rect 251 1755 252 1759
rect 246 1754 252 1755
rect 248 1734 250 1754
rect 246 1733 252 1734
rect 246 1729 247 1733
rect 251 1729 252 1733
rect 246 1728 252 1729
rect 272 1728 274 1777
rect 386 1759 392 1760
rect 386 1755 387 1759
rect 391 1755 392 1759
rect 386 1754 392 1755
rect 388 1734 390 1754
rect 386 1733 392 1734
rect 386 1729 387 1733
rect 391 1729 392 1733
rect 386 1728 392 1729
rect 408 1728 410 1777
rect 522 1759 528 1760
rect 522 1755 523 1759
rect 527 1755 528 1759
rect 522 1754 528 1755
rect 524 1734 526 1754
rect 522 1733 528 1734
rect 522 1729 523 1733
rect 527 1729 528 1733
rect 522 1728 528 1729
rect 544 1728 546 1777
rect 658 1759 664 1760
rect 658 1755 659 1759
rect 663 1755 664 1759
rect 658 1754 664 1755
rect 660 1734 662 1754
rect 658 1733 664 1734
rect 658 1729 659 1733
rect 663 1729 664 1733
rect 658 1728 664 1729
rect 680 1728 682 1777
rect 766 1733 772 1734
rect 766 1729 767 1733
rect 771 1729 772 1733
rect 1720 1730 1722 1777
rect 766 1728 772 1729
rect 1718 1729 1724 1730
rect 110 1724 116 1725
rect 134 1727 140 1728
rect 134 1723 135 1727
rect 139 1723 140 1727
rect 134 1722 140 1723
rect 270 1727 276 1728
rect 270 1723 271 1727
rect 275 1723 276 1727
rect 270 1722 276 1723
rect 406 1727 412 1728
rect 406 1723 407 1727
rect 411 1723 412 1727
rect 406 1722 412 1723
rect 542 1727 548 1728
rect 542 1723 543 1727
rect 547 1723 548 1727
rect 542 1722 548 1723
rect 678 1727 684 1728
rect 678 1723 679 1727
rect 683 1723 684 1727
rect 678 1722 684 1723
rect 158 1712 164 1713
rect 110 1711 116 1712
rect 110 1707 111 1711
rect 115 1707 116 1711
rect 158 1708 159 1712
rect 163 1708 164 1712
rect 158 1707 164 1708
rect 294 1712 300 1713
rect 294 1708 295 1712
rect 299 1708 300 1712
rect 294 1707 300 1708
rect 430 1712 436 1713
rect 430 1708 431 1712
rect 435 1708 436 1712
rect 430 1707 436 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 702 1712 708 1713
rect 702 1708 703 1712
rect 707 1708 708 1712
rect 702 1707 708 1708
rect 110 1706 116 1707
rect 112 1671 114 1706
rect 160 1671 162 1707
rect 296 1671 298 1707
rect 432 1671 434 1707
rect 568 1671 570 1707
rect 704 1671 706 1707
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 159 1670 163 1671
rect 159 1665 163 1666
rect 231 1670 235 1671
rect 231 1665 235 1666
rect 295 1670 299 1671
rect 295 1665 299 1666
rect 367 1670 371 1671
rect 367 1665 371 1666
rect 431 1670 435 1671
rect 431 1665 435 1666
rect 503 1670 507 1671
rect 503 1665 507 1666
rect 567 1670 571 1671
rect 567 1665 571 1666
rect 639 1670 643 1671
rect 639 1665 643 1666
rect 703 1670 707 1671
rect 703 1665 707 1666
rect 112 1642 114 1665
rect 110 1641 116 1642
rect 232 1641 234 1665
rect 368 1641 370 1665
rect 504 1641 506 1665
rect 640 1641 642 1665
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 110 1636 116 1637
rect 230 1640 236 1641
rect 230 1636 231 1640
rect 235 1636 236 1640
rect 230 1635 236 1636
rect 366 1640 372 1641
rect 366 1636 367 1640
rect 371 1636 372 1640
rect 366 1635 372 1636
rect 502 1640 508 1641
rect 502 1636 503 1640
rect 507 1636 508 1640
rect 502 1635 508 1636
rect 638 1640 644 1641
rect 638 1636 639 1640
rect 643 1636 644 1640
rect 638 1635 644 1636
rect 206 1625 212 1626
rect 110 1623 116 1624
rect 110 1619 111 1623
rect 115 1619 116 1623
rect 206 1621 207 1625
rect 211 1621 212 1625
rect 206 1620 212 1621
rect 342 1625 348 1626
rect 342 1621 343 1625
rect 347 1621 348 1625
rect 342 1620 348 1621
rect 478 1625 484 1626
rect 478 1621 479 1625
rect 483 1621 484 1625
rect 478 1620 484 1621
rect 614 1625 620 1626
rect 614 1621 615 1625
rect 619 1621 620 1625
rect 614 1620 620 1621
rect 750 1625 756 1626
rect 750 1621 751 1625
rect 755 1621 756 1625
rect 750 1620 756 1621
rect 110 1618 116 1619
rect 112 1559 114 1618
rect 208 1559 210 1620
rect 344 1559 346 1620
rect 350 1619 356 1620
rect 350 1615 351 1619
rect 355 1615 356 1619
rect 350 1614 356 1615
rect 352 1592 354 1614
rect 350 1591 356 1592
rect 350 1587 351 1591
rect 355 1587 356 1591
rect 350 1586 356 1587
rect 480 1559 482 1620
rect 486 1619 492 1620
rect 486 1615 487 1619
rect 491 1615 492 1619
rect 486 1614 492 1615
rect 488 1592 490 1614
rect 594 1611 600 1612
rect 594 1607 595 1611
rect 599 1607 600 1611
rect 594 1606 600 1607
rect 486 1591 492 1592
rect 486 1587 487 1591
rect 491 1587 492 1591
rect 486 1586 492 1587
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 207 1558 211 1559
rect 207 1553 211 1554
rect 343 1558 347 1559
rect 343 1553 347 1554
rect 479 1558 483 1559
rect 479 1553 483 1554
rect 487 1558 491 1559
rect 487 1553 491 1554
rect 112 1506 114 1553
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 488 1504 490 1553
rect 596 1540 598 1606
rect 616 1559 618 1620
rect 622 1619 628 1620
rect 622 1615 623 1619
rect 627 1615 628 1619
rect 622 1614 628 1615
rect 624 1592 626 1614
rect 622 1591 628 1592
rect 622 1587 623 1591
rect 627 1587 628 1591
rect 622 1586 628 1587
rect 752 1559 754 1620
rect 758 1619 764 1620
rect 758 1615 759 1619
rect 763 1615 764 1619
rect 758 1614 764 1615
rect 760 1592 762 1614
rect 768 1600 770 1728
rect 1718 1725 1719 1729
rect 1723 1725 1724 1729
rect 1718 1724 1724 1725
rect 1718 1711 1724 1712
rect 1718 1707 1719 1711
rect 1723 1707 1724 1711
rect 1718 1706 1724 1707
rect 1720 1671 1722 1706
rect 775 1670 779 1671
rect 775 1665 779 1666
rect 1719 1670 1723 1671
rect 1719 1665 1723 1666
rect 776 1641 778 1665
rect 1720 1642 1722 1665
rect 1718 1641 1724 1642
rect 774 1640 780 1641
rect 774 1636 775 1640
rect 779 1636 780 1640
rect 1718 1637 1719 1641
rect 1723 1637 1724 1641
rect 1718 1636 1724 1637
rect 774 1635 780 1636
rect 1718 1623 1724 1624
rect 1718 1619 1719 1623
rect 1723 1619 1724 1623
rect 1718 1618 1724 1619
rect 766 1599 772 1600
rect 766 1595 767 1599
rect 771 1595 772 1599
rect 766 1594 772 1595
rect 758 1591 764 1592
rect 758 1587 759 1591
rect 763 1587 764 1591
rect 758 1586 764 1587
rect 1720 1559 1722 1618
rect 615 1558 619 1559
rect 615 1553 619 1554
rect 623 1558 627 1559
rect 623 1553 627 1554
rect 751 1558 755 1559
rect 751 1553 755 1554
rect 759 1558 763 1559
rect 759 1553 763 1554
rect 895 1558 899 1559
rect 895 1553 899 1554
rect 1031 1558 1035 1559
rect 1031 1553 1035 1554
rect 1167 1558 1171 1559
rect 1167 1553 1171 1554
rect 1303 1558 1307 1559
rect 1303 1553 1307 1554
rect 1439 1558 1443 1559
rect 1439 1553 1443 1554
rect 1575 1558 1579 1559
rect 1575 1553 1579 1554
rect 1719 1558 1723 1559
rect 1719 1553 1723 1554
rect 594 1539 600 1540
rect 594 1535 595 1539
rect 599 1535 600 1539
rect 594 1534 600 1535
rect 602 1535 608 1536
rect 602 1531 603 1535
rect 607 1531 608 1535
rect 602 1530 608 1531
rect 604 1510 606 1530
rect 602 1509 608 1510
rect 602 1505 603 1509
rect 607 1505 608 1509
rect 602 1504 608 1505
rect 624 1504 626 1553
rect 738 1535 744 1536
rect 738 1531 739 1535
rect 743 1531 744 1535
rect 738 1530 744 1531
rect 740 1510 742 1530
rect 738 1509 744 1510
rect 738 1505 739 1509
rect 743 1505 744 1509
rect 738 1504 744 1505
rect 760 1504 762 1553
rect 874 1535 880 1536
rect 874 1531 875 1535
rect 879 1531 880 1535
rect 874 1530 880 1531
rect 876 1510 878 1530
rect 874 1509 880 1510
rect 874 1505 875 1509
rect 879 1505 880 1509
rect 874 1504 880 1505
rect 896 1504 898 1553
rect 1010 1535 1016 1536
rect 1010 1531 1011 1535
rect 1015 1531 1016 1535
rect 1010 1530 1016 1531
rect 1012 1510 1014 1530
rect 1010 1509 1016 1510
rect 1010 1505 1011 1509
rect 1015 1505 1016 1509
rect 1010 1504 1016 1505
rect 1032 1504 1034 1553
rect 1110 1509 1116 1510
rect 1110 1505 1111 1509
rect 1115 1505 1116 1509
rect 1110 1504 1116 1505
rect 1168 1504 1170 1553
rect 1274 1539 1280 1540
rect 1274 1535 1275 1539
rect 1279 1535 1280 1539
rect 1274 1534 1280 1535
rect 1282 1535 1288 1536
rect 110 1500 116 1501
rect 486 1503 492 1504
rect 486 1499 487 1503
rect 491 1499 492 1503
rect 486 1498 492 1499
rect 622 1503 628 1504
rect 622 1499 623 1503
rect 627 1499 628 1503
rect 622 1498 628 1499
rect 758 1503 764 1504
rect 758 1499 759 1503
rect 763 1499 764 1503
rect 758 1498 764 1499
rect 894 1503 900 1504
rect 894 1499 895 1503
rect 899 1499 900 1503
rect 894 1498 900 1499
rect 1030 1503 1036 1504
rect 1030 1499 1031 1503
rect 1035 1499 1036 1503
rect 1030 1498 1036 1499
rect 510 1488 516 1489
rect 110 1487 116 1488
rect 110 1483 111 1487
rect 115 1483 116 1487
rect 510 1484 511 1488
rect 515 1484 516 1488
rect 510 1483 516 1484
rect 646 1488 652 1489
rect 646 1484 647 1488
rect 651 1484 652 1488
rect 646 1483 652 1484
rect 782 1488 788 1489
rect 782 1484 783 1488
rect 787 1484 788 1488
rect 782 1483 788 1484
rect 918 1488 924 1489
rect 918 1484 919 1488
rect 923 1484 924 1488
rect 918 1483 924 1484
rect 1054 1488 1060 1489
rect 1054 1484 1055 1488
rect 1059 1484 1060 1488
rect 1054 1483 1060 1484
rect 110 1482 116 1483
rect 112 1443 114 1482
rect 512 1443 514 1483
rect 648 1443 650 1483
rect 784 1443 786 1483
rect 920 1443 922 1483
rect 1056 1443 1058 1483
rect 111 1442 115 1443
rect 111 1437 115 1438
rect 511 1442 515 1443
rect 511 1437 515 1438
rect 623 1442 627 1443
rect 623 1437 627 1438
rect 647 1442 651 1443
rect 647 1437 651 1438
rect 759 1442 763 1443
rect 759 1437 763 1438
rect 783 1442 787 1443
rect 783 1437 787 1438
rect 895 1442 899 1443
rect 895 1437 899 1438
rect 919 1442 923 1443
rect 919 1437 923 1438
rect 1039 1442 1043 1443
rect 1039 1437 1043 1438
rect 1055 1442 1059 1443
rect 1055 1437 1059 1438
rect 112 1414 114 1437
rect 110 1413 116 1414
rect 624 1413 626 1437
rect 760 1413 762 1437
rect 896 1413 898 1437
rect 1040 1413 1042 1437
rect 110 1409 111 1413
rect 115 1409 116 1413
rect 110 1408 116 1409
rect 622 1412 628 1413
rect 622 1408 623 1412
rect 627 1408 628 1412
rect 622 1407 628 1408
rect 758 1412 764 1413
rect 758 1408 759 1412
rect 763 1408 764 1412
rect 758 1407 764 1408
rect 894 1412 900 1413
rect 894 1408 895 1412
rect 899 1408 900 1412
rect 894 1407 900 1408
rect 1038 1412 1044 1413
rect 1038 1408 1039 1412
rect 1043 1408 1044 1412
rect 1038 1407 1044 1408
rect 598 1397 604 1398
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 598 1393 599 1397
rect 603 1393 604 1397
rect 598 1392 604 1393
rect 734 1397 740 1398
rect 734 1393 735 1397
rect 739 1393 740 1397
rect 734 1392 740 1393
rect 870 1397 876 1398
rect 870 1393 871 1397
rect 875 1393 876 1397
rect 870 1392 876 1393
rect 1014 1397 1020 1398
rect 1014 1393 1015 1397
rect 1019 1393 1020 1397
rect 1014 1392 1020 1393
rect 110 1390 116 1391
rect 112 1327 114 1390
rect 600 1327 602 1392
rect 674 1383 680 1384
rect 674 1379 675 1383
rect 679 1379 680 1383
rect 674 1378 680 1379
rect 676 1364 678 1378
rect 674 1363 680 1364
rect 674 1359 675 1363
rect 679 1359 680 1363
rect 674 1358 680 1359
rect 736 1327 738 1392
rect 742 1391 748 1392
rect 742 1387 743 1391
rect 747 1387 748 1391
rect 742 1386 748 1387
rect 744 1364 746 1386
rect 742 1363 748 1364
rect 742 1359 743 1363
rect 747 1359 748 1363
rect 742 1358 748 1359
rect 872 1327 874 1392
rect 878 1391 884 1392
rect 878 1387 879 1391
rect 883 1387 884 1391
rect 878 1386 884 1387
rect 970 1391 976 1392
rect 970 1387 971 1391
rect 975 1387 976 1391
rect 970 1386 976 1387
rect 880 1364 882 1386
rect 972 1372 974 1386
rect 970 1371 976 1372
rect 970 1367 971 1371
rect 975 1367 976 1371
rect 970 1366 976 1367
rect 878 1363 884 1364
rect 878 1359 879 1363
rect 883 1359 884 1363
rect 878 1358 884 1359
rect 1016 1327 1018 1392
rect 1112 1364 1114 1504
rect 1166 1503 1172 1504
rect 1166 1499 1167 1503
rect 1171 1499 1172 1503
rect 1166 1498 1172 1499
rect 1190 1488 1196 1489
rect 1190 1484 1191 1488
rect 1195 1484 1196 1488
rect 1190 1483 1196 1484
rect 1192 1443 1194 1483
rect 1276 1459 1278 1534
rect 1282 1531 1283 1535
rect 1287 1531 1288 1535
rect 1282 1530 1288 1531
rect 1284 1510 1286 1530
rect 1282 1509 1288 1510
rect 1282 1505 1283 1509
rect 1287 1505 1288 1509
rect 1282 1504 1288 1505
rect 1304 1504 1306 1553
rect 1418 1535 1424 1536
rect 1418 1531 1419 1535
rect 1423 1531 1424 1535
rect 1418 1530 1424 1531
rect 1420 1510 1422 1530
rect 1418 1509 1424 1510
rect 1418 1505 1419 1509
rect 1423 1505 1424 1509
rect 1418 1504 1424 1505
rect 1440 1504 1442 1553
rect 1554 1535 1560 1536
rect 1554 1531 1555 1535
rect 1559 1531 1560 1535
rect 1554 1530 1560 1531
rect 1556 1510 1558 1530
rect 1554 1509 1560 1510
rect 1554 1505 1555 1509
rect 1559 1505 1560 1509
rect 1554 1504 1560 1505
rect 1576 1504 1578 1553
rect 1720 1506 1722 1553
rect 1718 1505 1724 1506
rect 1302 1503 1308 1504
rect 1302 1499 1303 1503
rect 1307 1499 1308 1503
rect 1302 1498 1308 1499
rect 1438 1503 1444 1504
rect 1438 1499 1439 1503
rect 1443 1499 1444 1503
rect 1438 1498 1444 1499
rect 1574 1503 1580 1504
rect 1574 1499 1575 1503
rect 1579 1499 1580 1503
rect 1718 1501 1719 1505
rect 1723 1501 1724 1505
rect 1718 1500 1724 1501
rect 1574 1498 1580 1499
rect 1326 1488 1332 1489
rect 1326 1484 1327 1488
rect 1331 1484 1332 1488
rect 1326 1483 1332 1484
rect 1462 1488 1468 1489
rect 1462 1484 1463 1488
rect 1467 1484 1468 1488
rect 1462 1483 1468 1484
rect 1598 1488 1604 1489
rect 1598 1484 1599 1488
rect 1603 1484 1604 1488
rect 1598 1483 1604 1484
rect 1718 1487 1724 1488
rect 1718 1483 1719 1487
rect 1723 1483 1724 1487
rect 1276 1457 1282 1459
rect 1183 1442 1187 1443
rect 1183 1437 1187 1438
rect 1191 1442 1195 1443
rect 1191 1437 1195 1438
rect 1184 1413 1186 1437
rect 1182 1412 1188 1413
rect 1182 1408 1183 1412
rect 1187 1408 1188 1412
rect 1182 1407 1188 1408
rect 1158 1397 1164 1398
rect 1158 1393 1159 1397
rect 1163 1393 1164 1397
rect 1158 1392 1164 1393
rect 1280 1392 1282 1457
rect 1328 1443 1330 1483
rect 1464 1443 1466 1483
rect 1600 1443 1602 1483
rect 1718 1482 1724 1483
rect 1720 1443 1722 1482
rect 1327 1442 1331 1443
rect 1327 1437 1331 1438
rect 1463 1442 1467 1443
rect 1463 1437 1467 1438
rect 1599 1442 1603 1443
rect 1599 1437 1603 1438
rect 1719 1442 1723 1443
rect 1719 1437 1723 1438
rect 1328 1413 1330 1437
rect 1464 1413 1466 1437
rect 1600 1413 1602 1437
rect 1720 1414 1722 1437
rect 1718 1413 1724 1414
rect 1326 1412 1332 1413
rect 1326 1408 1327 1412
rect 1331 1408 1332 1412
rect 1326 1407 1332 1408
rect 1462 1412 1468 1413
rect 1462 1408 1463 1412
rect 1467 1408 1468 1412
rect 1462 1407 1468 1408
rect 1598 1412 1604 1413
rect 1598 1408 1599 1412
rect 1603 1408 1604 1412
rect 1718 1409 1719 1413
rect 1723 1409 1724 1413
rect 1718 1408 1724 1409
rect 1598 1407 1604 1408
rect 1302 1397 1308 1398
rect 1302 1393 1303 1397
rect 1307 1393 1308 1397
rect 1302 1392 1308 1393
rect 1438 1397 1444 1398
rect 1438 1393 1439 1397
rect 1443 1393 1444 1397
rect 1438 1392 1444 1393
rect 1574 1397 1580 1398
rect 1574 1393 1575 1397
rect 1579 1393 1580 1397
rect 1574 1392 1580 1393
rect 1718 1395 1724 1396
rect 1110 1363 1116 1364
rect 1110 1359 1111 1363
rect 1115 1359 1116 1363
rect 1110 1358 1116 1359
rect 1160 1327 1162 1392
rect 1254 1391 1260 1392
rect 1254 1387 1255 1391
rect 1259 1387 1260 1391
rect 1254 1386 1260 1387
rect 1278 1391 1284 1392
rect 1278 1387 1279 1391
rect 1283 1387 1284 1391
rect 1278 1386 1284 1387
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 135 1326 139 1327
rect 135 1321 139 1322
rect 343 1326 347 1327
rect 343 1321 347 1322
rect 599 1326 603 1327
rect 599 1321 603 1322
rect 607 1326 611 1327
rect 607 1321 611 1322
rect 735 1326 739 1327
rect 735 1321 739 1322
rect 871 1326 875 1327
rect 871 1321 875 1322
rect 895 1326 899 1327
rect 895 1321 899 1322
rect 1015 1326 1019 1327
rect 1015 1321 1019 1322
rect 1159 1326 1163 1327
rect 1159 1321 1163 1322
rect 1207 1326 1211 1327
rect 1207 1321 1211 1322
rect 112 1274 114 1321
rect 110 1273 116 1274
rect 110 1269 111 1273
rect 115 1269 116 1273
rect 136 1272 138 1321
rect 344 1272 346 1321
rect 526 1307 532 1308
rect 526 1303 527 1307
rect 531 1303 532 1307
rect 526 1302 532 1303
rect 528 1280 530 1302
rect 526 1279 532 1280
rect 526 1275 527 1279
rect 531 1275 532 1279
rect 526 1274 532 1275
rect 608 1272 610 1321
rect 886 1307 892 1308
rect 886 1303 887 1307
rect 891 1303 892 1307
rect 886 1302 892 1303
rect 888 1280 890 1302
rect 886 1279 892 1280
rect 886 1275 887 1279
rect 891 1275 892 1279
rect 886 1274 892 1275
rect 896 1272 898 1321
rect 1198 1307 1204 1308
rect 1198 1303 1199 1307
rect 1203 1303 1204 1307
rect 1198 1302 1204 1303
rect 1200 1280 1202 1302
rect 1198 1279 1204 1280
rect 1198 1275 1199 1279
rect 1203 1275 1204 1279
rect 1198 1274 1204 1275
rect 1208 1272 1210 1321
rect 1256 1304 1258 1386
rect 1304 1327 1306 1392
rect 1358 1363 1364 1364
rect 1358 1359 1359 1363
rect 1363 1359 1364 1363
rect 1358 1358 1364 1359
rect 1303 1326 1307 1327
rect 1303 1321 1307 1322
rect 1254 1303 1260 1304
rect 1254 1299 1255 1303
rect 1259 1299 1260 1303
rect 1254 1298 1260 1299
rect 110 1268 116 1269
rect 134 1271 140 1272
rect 134 1267 135 1271
rect 139 1267 140 1271
rect 134 1266 140 1267
rect 342 1271 348 1272
rect 342 1267 343 1271
rect 347 1267 348 1271
rect 342 1266 348 1267
rect 606 1271 612 1272
rect 606 1267 607 1271
rect 611 1267 612 1271
rect 606 1266 612 1267
rect 894 1271 900 1272
rect 894 1267 895 1271
rect 899 1267 900 1271
rect 894 1266 900 1267
rect 1206 1271 1212 1272
rect 1206 1267 1207 1271
rect 1211 1267 1212 1271
rect 1206 1266 1212 1267
rect 158 1256 164 1257
rect 110 1255 116 1256
rect 110 1251 111 1255
rect 115 1251 116 1255
rect 158 1252 159 1256
rect 163 1252 164 1256
rect 158 1251 164 1252
rect 366 1256 372 1257
rect 366 1252 367 1256
rect 371 1252 372 1256
rect 366 1251 372 1252
rect 630 1256 636 1257
rect 630 1252 631 1256
rect 635 1252 636 1256
rect 630 1251 636 1252
rect 918 1256 924 1257
rect 918 1252 919 1256
rect 923 1252 924 1256
rect 918 1251 924 1252
rect 1230 1256 1236 1257
rect 1230 1252 1231 1256
rect 1235 1252 1236 1256
rect 1230 1251 1236 1252
rect 110 1250 116 1251
rect 112 1215 114 1250
rect 160 1215 162 1251
rect 368 1215 370 1251
rect 632 1215 634 1251
rect 920 1215 922 1251
rect 1232 1215 1234 1251
rect 111 1214 115 1215
rect 111 1209 115 1210
rect 159 1214 163 1215
rect 159 1209 163 1210
rect 327 1214 331 1215
rect 327 1209 331 1210
rect 367 1214 371 1215
rect 367 1209 371 1210
rect 543 1214 547 1215
rect 543 1209 547 1210
rect 631 1214 635 1215
rect 631 1209 635 1210
rect 775 1214 779 1215
rect 775 1209 779 1210
rect 919 1214 923 1215
rect 919 1209 923 1210
rect 1023 1214 1027 1215
rect 1023 1209 1027 1210
rect 1231 1214 1235 1215
rect 1231 1209 1235 1210
rect 1287 1214 1291 1215
rect 1287 1209 1291 1210
rect 112 1186 114 1209
rect 110 1185 116 1186
rect 160 1185 162 1209
rect 328 1185 330 1209
rect 544 1185 546 1209
rect 776 1185 778 1209
rect 1024 1185 1026 1209
rect 1288 1185 1290 1209
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 158 1184 164 1185
rect 158 1180 159 1184
rect 163 1180 164 1184
rect 158 1179 164 1180
rect 326 1184 332 1185
rect 326 1180 327 1184
rect 331 1180 332 1184
rect 326 1179 332 1180
rect 542 1184 548 1185
rect 542 1180 543 1184
rect 547 1180 548 1184
rect 542 1179 548 1180
rect 774 1184 780 1185
rect 774 1180 775 1184
rect 779 1180 780 1184
rect 774 1179 780 1180
rect 1022 1184 1028 1185
rect 1022 1180 1023 1184
rect 1027 1180 1028 1184
rect 1022 1179 1028 1180
rect 1286 1184 1292 1185
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 134 1169 140 1170
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 134 1165 135 1169
rect 139 1165 140 1169
rect 134 1164 140 1165
rect 302 1169 308 1170
rect 302 1165 303 1169
rect 307 1165 308 1169
rect 302 1164 308 1165
rect 518 1169 524 1170
rect 518 1165 519 1169
rect 523 1165 524 1169
rect 518 1164 524 1165
rect 750 1169 756 1170
rect 750 1165 751 1169
rect 755 1165 756 1169
rect 750 1164 756 1165
rect 998 1169 1004 1170
rect 998 1165 999 1169
rect 1003 1165 1004 1169
rect 998 1164 1004 1165
rect 1262 1169 1268 1170
rect 1262 1165 1263 1169
rect 1267 1165 1268 1169
rect 1262 1164 1268 1165
rect 1360 1164 1362 1358
rect 1440 1327 1442 1392
rect 1534 1391 1540 1392
rect 1534 1387 1535 1391
rect 1539 1387 1540 1391
rect 1534 1386 1540 1387
rect 1558 1391 1564 1392
rect 1558 1387 1559 1391
rect 1563 1387 1564 1391
rect 1558 1386 1564 1387
rect 1439 1326 1443 1327
rect 1439 1321 1443 1322
rect 1519 1326 1523 1327
rect 1519 1321 1523 1322
rect 1520 1272 1522 1321
rect 1536 1304 1538 1386
rect 1560 1364 1562 1386
rect 1558 1363 1564 1364
rect 1558 1359 1559 1363
rect 1563 1359 1564 1363
rect 1558 1358 1564 1359
rect 1576 1327 1578 1392
rect 1718 1391 1719 1395
rect 1723 1391 1724 1395
rect 1718 1390 1724 1391
rect 1720 1327 1722 1390
rect 1575 1326 1579 1327
rect 1575 1321 1579 1322
rect 1719 1326 1723 1327
rect 1719 1321 1723 1322
rect 1534 1303 1540 1304
rect 1534 1299 1535 1303
rect 1539 1299 1540 1303
rect 1534 1298 1540 1299
rect 1602 1277 1608 1278
rect 1602 1273 1603 1277
rect 1607 1273 1608 1277
rect 1720 1274 1722 1321
rect 1602 1272 1608 1273
rect 1718 1273 1724 1274
rect 1518 1271 1524 1272
rect 1518 1267 1519 1271
rect 1523 1267 1524 1271
rect 1518 1266 1524 1267
rect 1542 1256 1548 1257
rect 1542 1252 1543 1256
rect 1547 1252 1548 1256
rect 1542 1251 1548 1252
rect 1544 1215 1546 1251
rect 1543 1214 1547 1215
rect 1543 1209 1547 1210
rect 1551 1214 1555 1215
rect 1551 1209 1555 1210
rect 1552 1185 1554 1209
rect 1550 1184 1556 1185
rect 1550 1180 1551 1184
rect 1555 1180 1556 1184
rect 1550 1179 1556 1180
rect 1526 1169 1532 1170
rect 1526 1165 1527 1169
rect 1531 1165 1532 1169
rect 1526 1164 1532 1165
rect 110 1162 116 1163
rect 112 1095 114 1162
rect 136 1095 138 1164
rect 304 1095 306 1164
rect 310 1163 316 1164
rect 310 1159 311 1163
rect 315 1159 316 1163
rect 310 1158 316 1159
rect 312 1136 314 1158
rect 418 1151 424 1152
rect 418 1147 419 1151
rect 423 1147 424 1151
rect 418 1146 424 1147
rect 310 1135 316 1136
rect 310 1131 311 1135
rect 315 1131 316 1135
rect 310 1130 316 1131
rect 111 1094 115 1095
rect 111 1089 115 1090
rect 135 1094 139 1095
rect 135 1089 139 1090
rect 303 1094 307 1095
rect 303 1089 307 1090
rect 311 1094 315 1095
rect 311 1089 315 1090
rect 112 1042 114 1089
rect 110 1041 116 1042
rect 110 1037 111 1041
rect 115 1037 116 1041
rect 312 1040 314 1089
rect 420 1076 422 1146
rect 520 1095 522 1164
rect 526 1163 532 1164
rect 526 1159 527 1163
rect 531 1159 532 1163
rect 526 1158 532 1159
rect 528 1136 530 1158
rect 526 1135 532 1136
rect 526 1131 527 1135
rect 531 1131 532 1135
rect 526 1130 532 1131
rect 752 1095 754 1164
rect 758 1163 764 1164
rect 758 1159 759 1163
rect 763 1159 764 1163
rect 758 1158 764 1159
rect 760 1136 762 1158
rect 758 1135 764 1136
rect 758 1131 759 1135
rect 763 1131 764 1135
rect 758 1130 764 1131
rect 1000 1095 1002 1164
rect 1006 1163 1012 1164
rect 1006 1159 1007 1163
rect 1011 1159 1012 1163
rect 1006 1158 1012 1159
rect 1008 1136 1010 1158
rect 1006 1135 1012 1136
rect 1006 1131 1007 1135
rect 1011 1131 1012 1135
rect 1006 1130 1012 1131
rect 1264 1095 1266 1164
rect 1358 1163 1364 1164
rect 1358 1159 1359 1163
rect 1363 1159 1364 1163
rect 1358 1158 1364 1159
rect 1358 1135 1364 1136
rect 1358 1131 1359 1135
rect 1363 1131 1364 1135
rect 1358 1130 1364 1131
rect 519 1094 523 1095
rect 519 1089 523 1090
rect 535 1094 539 1095
rect 535 1089 539 1090
rect 751 1094 755 1095
rect 751 1089 755 1090
rect 775 1094 779 1095
rect 775 1089 779 1090
rect 999 1094 1003 1095
rect 999 1089 1003 1090
rect 1023 1094 1027 1095
rect 1023 1089 1027 1090
rect 1263 1094 1267 1095
rect 1263 1089 1267 1090
rect 1279 1094 1283 1095
rect 1279 1089 1283 1090
rect 418 1075 424 1076
rect 418 1071 419 1075
rect 423 1071 424 1075
rect 418 1070 424 1071
rect 426 1071 432 1072
rect 426 1067 427 1071
rect 431 1067 432 1071
rect 426 1066 432 1067
rect 428 1046 430 1066
rect 426 1045 432 1046
rect 426 1041 427 1045
rect 431 1041 432 1045
rect 426 1040 432 1041
rect 536 1040 538 1089
rect 650 1071 656 1072
rect 650 1067 651 1071
rect 655 1067 656 1071
rect 650 1066 656 1067
rect 652 1046 654 1066
rect 650 1045 656 1046
rect 650 1041 651 1045
rect 655 1041 656 1045
rect 650 1040 656 1041
rect 776 1040 778 1089
rect 890 1071 896 1072
rect 890 1067 891 1071
rect 895 1067 896 1071
rect 890 1066 896 1067
rect 892 1046 894 1066
rect 890 1045 896 1046
rect 890 1041 891 1045
rect 895 1041 896 1045
rect 890 1040 896 1041
rect 1024 1040 1026 1089
rect 1102 1045 1108 1046
rect 1102 1041 1103 1045
rect 1107 1041 1108 1045
rect 1102 1040 1108 1041
rect 1280 1040 1282 1089
rect 1360 1046 1362 1130
rect 1528 1095 1530 1164
rect 1604 1136 1606 1272
rect 1718 1269 1719 1273
rect 1723 1269 1724 1273
rect 1718 1268 1724 1269
rect 1718 1255 1724 1256
rect 1718 1251 1719 1255
rect 1723 1251 1724 1255
rect 1718 1250 1724 1251
rect 1720 1215 1722 1250
rect 1719 1214 1723 1215
rect 1719 1209 1723 1210
rect 1720 1186 1722 1209
rect 1718 1185 1724 1186
rect 1718 1181 1719 1185
rect 1723 1181 1724 1185
rect 1718 1180 1724 1181
rect 1718 1167 1724 1168
rect 1618 1163 1624 1164
rect 1618 1159 1619 1163
rect 1623 1159 1624 1163
rect 1718 1163 1719 1167
rect 1723 1163 1724 1167
rect 1718 1162 1724 1163
rect 1618 1158 1624 1159
rect 1602 1135 1608 1136
rect 1602 1131 1603 1135
rect 1607 1131 1608 1135
rect 1602 1130 1608 1131
rect 1527 1094 1531 1095
rect 1527 1089 1531 1090
rect 1543 1094 1547 1095
rect 1543 1089 1547 1090
rect 1526 1075 1532 1076
rect 1526 1071 1527 1075
rect 1531 1071 1532 1075
rect 1526 1070 1532 1071
rect 1358 1045 1364 1046
rect 1358 1041 1359 1045
rect 1363 1041 1364 1045
rect 1358 1040 1364 1041
rect 110 1036 116 1037
rect 310 1039 316 1040
rect 310 1035 311 1039
rect 315 1035 316 1039
rect 310 1034 316 1035
rect 534 1039 540 1040
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 774 1039 780 1040
rect 774 1035 775 1039
rect 779 1035 780 1039
rect 774 1034 780 1035
rect 1022 1039 1028 1040
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1022 1034 1028 1035
rect 334 1024 340 1025
rect 110 1023 116 1024
rect 110 1019 111 1023
rect 115 1019 116 1023
rect 334 1020 335 1024
rect 339 1020 340 1024
rect 334 1019 340 1020
rect 558 1024 564 1025
rect 558 1020 559 1024
rect 563 1020 564 1024
rect 558 1019 564 1020
rect 798 1024 804 1025
rect 798 1020 799 1024
rect 803 1020 804 1024
rect 798 1019 804 1020
rect 1046 1024 1052 1025
rect 1046 1020 1047 1024
rect 1051 1020 1052 1024
rect 1046 1019 1052 1020
rect 110 1018 116 1019
rect 112 995 114 1018
rect 336 995 338 1019
rect 560 995 562 1019
rect 800 995 802 1019
rect 1048 995 1050 1019
rect 111 994 115 995
rect 111 989 115 990
rect 335 994 339 995
rect 335 989 339 990
rect 527 994 531 995
rect 527 989 531 990
rect 559 994 563 995
rect 559 989 563 990
rect 711 994 715 995
rect 711 989 715 990
rect 799 994 803 995
rect 799 989 803 990
rect 919 994 923 995
rect 919 989 923 990
rect 1047 994 1051 995
rect 1047 989 1051 990
rect 112 966 114 989
rect 110 965 116 966
rect 528 965 530 989
rect 712 965 714 989
rect 920 965 922 989
rect 110 961 111 965
rect 115 961 116 965
rect 110 960 116 961
rect 526 964 532 965
rect 526 960 527 964
rect 531 960 532 964
rect 526 959 532 960
rect 710 964 716 965
rect 710 960 711 964
rect 715 960 716 964
rect 710 959 716 960
rect 918 964 924 965
rect 918 960 919 964
rect 923 960 924 964
rect 918 959 924 960
rect 502 949 508 950
rect 110 947 116 948
rect 110 943 111 947
rect 115 943 116 947
rect 502 945 503 949
rect 507 945 508 949
rect 502 944 508 945
rect 686 949 692 950
rect 686 945 687 949
rect 691 945 692 949
rect 686 944 692 945
rect 894 949 900 950
rect 894 945 895 949
rect 899 945 900 949
rect 894 944 900 945
rect 110 942 116 943
rect 112 879 114 942
rect 504 879 506 944
rect 688 879 690 944
rect 694 943 700 944
rect 694 939 695 943
rect 699 939 700 943
rect 694 938 700 939
rect 696 916 698 938
rect 850 935 856 936
rect 850 931 851 935
rect 855 931 856 935
rect 850 930 856 931
rect 694 915 700 916
rect 694 911 695 915
rect 699 911 700 915
rect 694 910 700 911
rect 111 878 115 879
rect 111 873 115 874
rect 503 878 507 879
rect 503 873 507 874
rect 687 878 691 879
rect 687 873 691 874
rect 743 878 747 879
rect 743 873 747 874
rect 112 826 114 873
rect 110 825 116 826
rect 110 821 111 825
rect 115 821 116 825
rect 744 824 746 873
rect 852 860 854 930
rect 896 879 898 944
rect 902 943 908 944
rect 902 939 903 943
rect 907 939 908 943
rect 902 938 908 939
rect 904 916 906 938
rect 1104 924 1106 1040
rect 1278 1039 1284 1040
rect 1278 1035 1279 1039
rect 1283 1035 1284 1039
rect 1278 1034 1284 1035
rect 1302 1024 1308 1025
rect 1302 1020 1303 1024
rect 1307 1020 1308 1024
rect 1302 1019 1308 1020
rect 1304 995 1306 1019
rect 1135 994 1139 995
rect 1135 989 1139 990
rect 1303 994 1307 995
rect 1303 989 1307 990
rect 1367 994 1371 995
rect 1367 989 1371 990
rect 1136 965 1138 989
rect 1368 965 1370 989
rect 1134 964 1140 965
rect 1134 960 1135 964
rect 1139 960 1140 964
rect 1134 959 1140 960
rect 1366 964 1372 965
rect 1366 960 1367 964
rect 1371 960 1372 964
rect 1366 959 1372 960
rect 1110 949 1116 950
rect 1110 945 1111 949
rect 1115 945 1116 949
rect 1110 944 1116 945
rect 1342 949 1348 950
rect 1342 945 1343 949
rect 1347 945 1348 949
rect 1342 944 1348 945
rect 1102 923 1108 924
rect 1102 919 1103 923
rect 1107 919 1108 923
rect 1102 918 1108 919
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 1112 879 1114 944
rect 1118 943 1124 944
rect 1118 939 1119 943
rect 1123 939 1124 943
rect 1118 938 1124 939
rect 1120 916 1122 938
rect 1118 915 1124 916
rect 1118 911 1119 915
rect 1123 911 1124 915
rect 1118 910 1124 911
rect 1344 879 1346 944
rect 1350 943 1356 944
rect 1350 939 1351 943
rect 1355 939 1356 943
rect 1350 938 1356 939
rect 1352 916 1354 938
rect 1350 915 1356 916
rect 1350 911 1351 915
rect 1355 911 1356 915
rect 1350 910 1356 911
rect 879 878 883 879
rect 879 873 883 874
rect 895 878 899 879
rect 895 873 899 874
rect 1015 878 1019 879
rect 1015 873 1019 874
rect 1111 878 1115 879
rect 1111 873 1115 874
rect 1151 878 1155 879
rect 1151 873 1155 874
rect 1287 878 1291 879
rect 1287 873 1291 874
rect 1343 878 1347 879
rect 1343 873 1347 874
rect 1431 878 1435 879
rect 1431 873 1435 874
rect 850 859 856 860
rect 850 855 851 859
rect 855 855 856 859
rect 850 854 856 855
rect 858 855 864 856
rect 858 851 859 855
rect 863 851 864 855
rect 858 850 864 851
rect 860 830 862 850
rect 858 829 864 830
rect 858 825 859 829
rect 863 825 864 829
rect 858 824 864 825
rect 880 824 882 873
rect 994 855 1000 856
rect 994 851 995 855
rect 999 851 1000 855
rect 994 850 1000 851
rect 996 830 998 850
rect 994 829 1000 830
rect 994 825 995 829
rect 999 825 1000 829
rect 994 824 1000 825
rect 1016 824 1018 873
rect 1114 855 1120 856
rect 1114 851 1115 855
rect 1119 851 1120 855
rect 1114 850 1120 851
rect 1116 830 1118 850
rect 1114 829 1120 830
rect 1114 825 1115 829
rect 1119 825 1120 829
rect 1114 824 1120 825
rect 1152 824 1154 873
rect 1250 855 1256 856
rect 1250 851 1251 855
rect 1255 851 1256 855
rect 1250 850 1256 851
rect 1252 830 1254 850
rect 1250 829 1256 830
rect 1250 825 1251 829
rect 1255 825 1256 829
rect 1250 824 1256 825
rect 1288 824 1290 873
rect 1382 829 1388 830
rect 1382 825 1383 829
rect 1387 825 1388 829
rect 1382 824 1388 825
rect 1432 824 1434 873
rect 1438 855 1444 856
rect 1438 851 1439 855
rect 1443 851 1444 855
rect 1438 850 1444 851
rect 110 820 116 821
rect 742 823 748 824
rect 742 819 743 823
rect 747 819 748 823
rect 742 818 748 819
rect 878 823 884 824
rect 878 819 879 823
rect 883 819 884 823
rect 878 818 884 819
rect 1014 823 1020 824
rect 1014 819 1015 823
rect 1019 819 1020 823
rect 1014 818 1020 819
rect 1150 823 1156 824
rect 1150 819 1151 823
rect 1155 819 1156 823
rect 1150 818 1156 819
rect 1286 823 1292 824
rect 1286 819 1287 823
rect 1291 819 1292 823
rect 1286 818 1292 819
rect 766 808 772 809
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 766 804 767 808
rect 771 804 772 808
rect 766 803 772 804
rect 902 808 908 809
rect 902 804 903 808
rect 907 804 908 808
rect 902 803 908 804
rect 1038 808 1044 809
rect 1038 804 1039 808
rect 1043 804 1044 808
rect 1038 803 1044 804
rect 1174 808 1180 809
rect 1174 804 1175 808
rect 1179 804 1180 808
rect 1174 803 1180 804
rect 1310 808 1316 809
rect 1310 804 1311 808
rect 1315 804 1316 808
rect 1310 803 1316 804
rect 110 802 116 803
rect 112 763 114 802
rect 768 763 770 803
rect 904 763 906 803
rect 1040 763 1042 803
rect 1176 763 1178 803
rect 1312 763 1314 803
rect 111 762 115 763
rect 111 757 115 758
rect 703 762 707 763
rect 703 757 707 758
rect 767 762 771 763
rect 767 757 771 758
rect 863 762 867 763
rect 863 757 867 758
rect 903 762 907 763
rect 903 757 907 758
rect 1031 762 1035 763
rect 1031 757 1035 758
rect 1039 762 1043 763
rect 1039 757 1043 758
rect 1175 762 1179 763
rect 1175 757 1179 758
rect 1215 762 1219 763
rect 1215 757 1219 758
rect 1311 762 1315 763
rect 1311 757 1315 758
rect 112 734 114 757
rect 110 733 116 734
rect 704 733 706 757
rect 864 733 866 757
rect 1032 733 1034 757
rect 1216 733 1218 757
rect 110 729 111 733
rect 115 729 116 733
rect 110 728 116 729
rect 702 732 708 733
rect 702 728 703 732
rect 707 728 708 732
rect 702 727 708 728
rect 862 732 868 733
rect 862 728 863 732
rect 867 728 868 732
rect 862 727 868 728
rect 1030 732 1036 733
rect 1030 728 1031 732
rect 1035 728 1036 732
rect 1030 727 1036 728
rect 1214 732 1220 733
rect 1214 728 1215 732
rect 1219 728 1220 732
rect 1214 727 1220 728
rect 678 717 684 718
rect 110 715 116 716
rect 110 711 111 715
rect 115 711 116 715
rect 678 713 679 717
rect 683 713 684 717
rect 678 712 684 713
rect 838 717 844 718
rect 838 713 839 717
rect 843 713 844 717
rect 838 712 844 713
rect 1006 717 1012 718
rect 1006 713 1007 717
rect 1011 713 1012 717
rect 1006 712 1012 713
rect 1190 717 1196 718
rect 1190 713 1191 717
rect 1195 713 1196 717
rect 1190 712 1196 713
rect 1374 717 1380 718
rect 1374 713 1375 717
rect 1379 713 1380 717
rect 1374 712 1380 713
rect 110 710 116 711
rect 112 663 114 710
rect 680 663 682 712
rect 754 703 760 704
rect 754 699 755 703
rect 759 699 760 703
rect 754 698 760 699
rect 756 684 758 698
rect 754 683 760 684
rect 754 679 755 683
rect 759 679 760 683
rect 754 678 760 679
rect 840 663 842 712
rect 846 711 852 712
rect 846 707 847 711
rect 851 707 852 711
rect 846 706 852 707
rect 848 684 850 706
rect 846 683 852 684
rect 846 679 847 683
rect 851 679 852 683
rect 846 678 852 679
rect 1008 663 1010 712
rect 1014 711 1020 712
rect 1014 707 1015 711
rect 1019 707 1020 711
rect 1014 706 1020 707
rect 1102 711 1108 712
rect 1102 707 1103 711
rect 1107 707 1108 711
rect 1102 706 1108 707
rect 1016 684 1018 706
rect 1014 683 1020 684
rect 1014 679 1015 683
rect 1019 679 1020 683
rect 1014 678 1020 679
rect 111 662 115 663
rect 111 657 115 658
rect 223 662 227 663
rect 223 657 227 658
rect 415 662 419 663
rect 415 657 419 658
rect 623 662 627 663
rect 623 657 627 658
rect 679 662 683 663
rect 679 657 683 658
rect 839 662 843 663
rect 839 657 843 658
rect 855 662 859 663
rect 855 657 859 658
rect 1007 662 1011 663
rect 1007 657 1011 658
rect 1095 662 1099 663
rect 1095 657 1099 658
rect 112 610 114 657
rect 210 615 216 616
rect 210 611 211 615
rect 215 611 216 615
rect 210 610 216 611
rect 110 609 116 610
rect 110 605 111 609
rect 115 605 116 609
rect 110 604 116 605
rect 110 591 116 592
rect 110 587 111 591
rect 115 587 116 591
rect 110 586 116 587
rect 112 551 114 586
rect 111 550 115 551
rect 111 545 115 546
rect 159 550 163 551
rect 159 545 163 546
rect 112 522 114 545
rect 110 521 116 522
rect 160 521 162 545
rect 110 517 111 521
rect 115 517 116 521
rect 110 516 116 517
rect 158 520 164 521
rect 158 516 159 520
rect 163 516 164 520
rect 158 515 164 516
rect 134 505 140 506
rect 110 503 116 504
rect 110 499 111 503
rect 115 499 116 503
rect 134 501 135 505
rect 139 501 140 505
rect 134 500 140 501
rect 110 498 116 499
rect 112 435 114 498
rect 136 435 138 500
rect 212 472 214 610
rect 224 608 226 657
rect 416 608 418 657
rect 624 608 626 657
rect 856 608 858 657
rect 1010 643 1016 644
rect 1010 639 1011 643
rect 1015 639 1016 643
rect 1010 638 1016 639
rect 1012 616 1014 638
rect 1010 615 1016 616
rect 1010 611 1011 615
rect 1015 611 1016 615
rect 1010 610 1016 611
rect 1096 608 1098 657
rect 1104 640 1106 706
rect 1192 663 1194 712
rect 1334 711 1340 712
rect 1334 707 1335 711
rect 1339 707 1340 711
rect 1334 706 1340 707
rect 1336 684 1338 706
rect 1334 683 1340 684
rect 1334 679 1335 683
rect 1339 679 1340 683
rect 1334 678 1340 679
rect 1376 663 1378 712
rect 1384 684 1386 824
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1399 762 1403 763
rect 1399 757 1403 758
rect 1400 733 1402 757
rect 1398 732 1404 733
rect 1398 728 1399 732
rect 1403 728 1404 732
rect 1398 727 1404 728
rect 1382 683 1388 684
rect 1382 679 1383 683
rect 1387 679 1388 683
rect 1382 678 1388 679
rect 1191 662 1195 663
rect 1191 657 1195 658
rect 1335 662 1339 663
rect 1335 657 1339 658
rect 1375 662 1379 663
rect 1375 657 1379 658
rect 1102 639 1108 640
rect 1102 635 1103 639
rect 1107 635 1108 639
rect 1102 634 1108 635
rect 1336 608 1338 657
rect 1374 639 1380 640
rect 1374 635 1375 639
rect 1379 635 1380 639
rect 1374 634 1380 635
rect 222 607 228 608
rect 222 603 223 607
rect 227 603 228 607
rect 222 602 228 603
rect 414 607 420 608
rect 414 603 415 607
rect 419 603 420 607
rect 414 602 420 603
rect 622 607 628 608
rect 622 603 623 607
rect 627 603 628 607
rect 622 602 628 603
rect 854 607 860 608
rect 854 603 855 607
rect 859 603 860 607
rect 854 602 860 603
rect 1094 607 1100 608
rect 1094 603 1095 607
rect 1099 603 1100 607
rect 1094 602 1100 603
rect 1334 607 1340 608
rect 1334 603 1335 607
rect 1339 603 1340 607
rect 1334 602 1340 603
rect 246 592 252 593
rect 246 588 247 592
rect 251 588 252 592
rect 246 587 252 588
rect 438 592 444 593
rect 438 588 439 592
rect 443 588 444 592
rect 438 587 444 588
rect 646 592 652 593
rect 646 588 647 592
rect 651 588 652 592
rect 646 587 652 588
rect 878 592 884 593
rect 878 588 879 592
rect 883 588 884 592
rect 878 587 884 588
rect 1118 592 1124 593
rect 1118 588 1119 592
rect 1123 588 1124 592
rect 1118 587 1124 588
rect 1358 592 1364 593
rect 1358 588 1359 592
rect 1363 588 1364 592
rect 1358 587 1364 588
rect 248 551 250 587
rect 440 551 442 587
rect 648 551 650 587
rect 880 551 882 587
rect 1120 551 1122 587
rect 1360 551 1362 587
rect 247 550 251 551
rect 247 545 251 546
rect 327 550 331 551
rect 327 545 331 546
rect 439 550 443 551
rect 439 545 443 546
rect 543 550 547 551
rect 543 545 547 546
rect 647 550 651 551
rect 647 545 651 546
rect 783 550 787 551
rect 783 545 787 546
rect 879 550 883 551
rect 879 545 883 546
rect 1039 550 1043 551
rect 1039 545 1043 546
rect 1119 550 1123 551
rect 1119 545 1123 546
rect 1303 550 1307 551
rect 1303 545 1307 546
rect 1359 550 1363 551
rect 1359 545 1363 546
rect 328 521 330 545
rect 544 521 546 545
rect 784 521 786 545
rect 1040 521 1042 545
rect 1304 521 1306 545
rect 326 520 332 521
rect 326 516 327 520
rect 331 516 332 520
rect 326 515 332 516
rect 542 520 548 521
rect 542 516 543 520
rect 547 516 548 520
rect 542 515 548 516
rect 782 520 788 521
rect 782 516 783 520
rect 787 516 788 520
rect 782 515 788 516
rect 1038 520 1044 521
rect 1038 516 1039 520
rect 1043 516 1044 520
rect 1038 515 1044 516
rect 1302 520 1308 521
rect 1302 516 1303 520
rect 1307 516 1308 520
rect 1302 515 1308 516
rect 302 505 308 506
rect 302 501 303 505
rect 307 501 308 505
rect 302 500 308 501
rect 518 505 524 506
rect 518 501 519 505
rect 523 501 524 505
rect 518 500 524 501
rect 758 505 764 506
rect 758 501 759 505
rect 763 501 764 505
rect 758 500 764 501
rect 1014 505 1020 506
rect 1014 501 1015 505
rect 1019 501 1020 505
rect 1014 500 1020 501
rect 1278 505 1284 506
rect 1278 501 1279 505
rect 1283 501 1284 505
rect 1278 500 1284 501
rect 1376 500 1378 634
rect 1440 614 1442 850
rect 1528 830 1530 1070
rect 1544 1040 1546 1089
rect 1620 1072 1622 1158
rect 1720 1095 1722 1162
rect 1719 1094 1723 1095
rect 1719 1089 1723 1090
rect 1618 1071 1624 1072
rect 1618 1067 1619 1071
rect 1623 1067 1624 1071
rect 1618 1066 1624 1067
rect 1638 1045 1644 1046
rect 1638 1041 1639 1045
rect 1643 1041 1644 1045
rect 1720 1042 1722 1089
rect 1638 1040 1644 1041
rect 1718 1041 1724 1042
rect 1542 1039 1548 1040
rect 1542 1035 1543 1039
rect 1547 1035 1548 1039
rect 1542 1034 1548 1035
rect 1566 1024 1572 1025
rect 1566 1020 1567 1024
rect 1571 1020 1572 1024
rect 1566 1019 1572 1020
rect 1568 995 1570 1019
rect 1567 994 1571 995
rect 1567 989 1571 990
rect 1599 994 1603 995
rect 1599 989 1603 990
rect 1600 965 1602 989
rect 1598 964 1604 965
rect 1598 960 1599 964
rect 1603 960 1604 964
rect 1598 959 1604 960
rect 1574 949 1580 950
rect 1574 945 1575 949
rect 1579 945 1580 949
rect 1574 944 1580 945
rect 1576 879 1578 944
rect 1640 916 1642 1040
rect 1718 1037 1719 1041
rect 1723 1037 1724 1041
rect 1718 1036 1724 1037
rect 1718 1023 1724 1024
rect 1718 1019 1719 1023
rect 1723 1019 1724 1023
rect 1718 1018 1724 1019
rect 1720 995 1722 1018
rect 1719 994 1723 995
rect 1719 989 1723 990
rect 1720 966 1722 989
rect 1718 965 1724 966
rect 1718 961 1719 965
rect 1723 961 1724 965
rect 1718 960 1724 961
rect 1718 947 1724 948
rect 1666 943 1672 944
rect 1666 939 1667 943
rect 1671 939 1672 943
rect 1718 943 1719 947
rect 1723 943 1724 947
rect 1718 942 1724 943
rect 1666 938 1672 939
rect 1638 915 1644 916
rect 1638 911 1639 915
rect 1643 911 1644 915
rect 1638 910 1644 911
rect 1575 878 1579 879
rect 1575 873 1579 874
rect 1526 829 1532 830
rect 1526 825 1527 829
rect 1531 825 1532 829
rect 1526 824 1532 825
rect 1576 824 1578 873
rect 1668 860 1670 938
rect 1720 879 1722 942
rect 1719 878 1723 879
rect 1719 873 1723 874
rect 1666 859 1672 860
rect 1666 855 1667 859
rect 1671 855 1672 859
rect 1666 854 1672 855
rect 1654 829 1660 830
rect 1654 825 1655 829
rect 1659 825 1660 829
rect 1720 826 1722 873
rect 1654 824 1660 825
rect 1718 825 1724 826
rect 1574 823 1580 824
rect 1574 819 1575 823
rect 1579 819 1580 823
rect 1574 818 1580 819
rect 1454 808 1460 809
rect 1454 804 1455 808
rect 1459 804 1460 808
rect 1454 803 1460 804
rect 1598 808 1604 809
rect 1598 804 1599 808
rect 1603 804 1604 808
rect 1598 803 1604 804
rect 1456 763 1458 803
rect 1600 763 1602 803
rect 1455 762 1459 763
rect 1455 757 1459 758
rect 1591 762 1595 763
rect 1591 757 1595 758
rect 1599 762 1603 763
rect 1599 757 1603 758
rect 1592 733 1594 757
rect 1590 732 1596 733
rect 1590 728 1591 732
rect 1595 728 1596 732
rect 1590 727 1596 728
rect 1566 717 1572 718
rect 1566 713 1567 717
rect 1571 713 1572 717
rect 1566 712 1572 713
rect 1568 663 1570 712
rect 1618 711 1624 712
rect 1618 707 1619 711
rect 1623 707 1624 711
rect 1618 706 1624 707
rect 1567 662 1571 663
rect 1567 657 1571 658
rect 1431 613 1442 614
rect 1431 609 1432 613
rect 1436 612 1442 613
rect 1436 609 1437 612
rect 1431 608 1437 609
rect 1567 550 1571 551
rect 1567 545 1571 546
rect 1568 521 1570 545
rect 1566 520 1572 521
rect 1566 516 1567 520
rect 1571 516 1572 520
rect 1566 515 1572 516
rect 1542 505 1548 506
rect 1542 501 1543 505
rect 1547 501 1548 505
rect 1542 500 1548 501
rect 290 491 296 492
rect 290 487 291 491
rect 295 487 296 491
rect 290 486 296 487
rect 210 471 216 472
rect 210 467 211 471
rect 215 467 216 471
rect 210 466 216 467
rect 111 434 115 435
rect 111 429 115 430
rect 135 434 139 435
rect 135 429 139 430
rect 199 434 203 435
rect 199 429 203 430
rect 112 382 114 429
rect 110 381 116 382
rect 110 377 111 381
rect 115 377 116 381
rect 200 380 202 429
rect 292 416 294 486
rect 304 435 306 500
rect 310 499 316 500
rect 310 495 311 499
rect 315 495 316 499
rect 310 494 316 495
rect 312 472 314 494
rect 310 471 316 472
rect 310 467 311 471
rect 315 467 316 471
rect 310 466 316 467
rect 520 435 522 500
rect 526 499 532 500
rect 526 495 527 499
rect 531 495 532 499
rect 526 494 532 495
rect 528 472 530 494
rect 526 471 532 472
rect 526 467 527 471
rect 531 467 532 471
rect 526 466 532 467
rect 760 435 762 500
rect 766 499 772 500
rect 766 495 767 499
rect 771 495 772 499
rect 766 494 772 495
rect 768 472 770 494
rect 766 471 772 472
rect 766 467 767 471
rect 771 467 772 471
rect 766 466 772 467
rect 1016 435 1018 500
rect 1022 499 1028 500
rect 1022 495 1023 499
rect 1027 495 1028 499
rect 1022 494 1028 495
rect 1024 472 1026 494
rect 1022 471 1028 472
rect 1022 467 1023 471
rect 1027 467 1028 471
rect 1022 466 1028 467
rect 1280 435 1282 500
rect 1374 499 1380 500
rect 1374 495 1375 499
rect 1379 495 1380 499
rect 1374 494 1380 495
rect 1414 471 1420 472
rect 1414 467 1415 471
rect 1419 467 1420 471
rect 1414 466 1420 467
rect 303 434 307 435
rect 303 429 307 430
rect 431 434 435 435
rect 431 429 435 430
rect 519 434 523 435
rect 519 429 523 430
rect 663 434 667 435
rect 663 429 667 430
rect 759 434 763 435
rect 759 429 763 430
rect 887 434 891 435
rect 887 429 891 430
rect 1015 434 1019 435
rect 1015 429 1019 430
rect 1111 434 1115 435
rect 1111 429 1115 430
rect 1279 434 1283 435
rect 1279 429 1283 430
rect 1335 434 1339 435
rect 1335 429 1339 430
rect 290 415 296 416
rect 290 411 291 415
rect 295 411 296 415
rect 290 410 296 411
rect 298 411 304 412
rect 298 407 299 411
rect 303 407 304 411
rect 298 406 304 407
rect 300 386 302 406
rect 298 385 304 386
rect 298 381 299 385
rect 303 381 304 385
rect 298 380 304 381
rect 432 380 434 429
rect 546 411 552 412
rect 546 407 547 411
rect 551 407 552 411
rect 546 406 552 407
rect 548 386 550 406
rect 546 385 552 386
rect 546 381 547 385
rect 551 381 552 385
rect 546 380 552 381
rect 664 380 666 429
rect 762 385 768 386
rect 762 381 763 385
rect 767 381 768 385
rect 762 380 768 381
rect 888 380 890 429
rect 1002 411 1008 412
rect 1002 407 1003 411
rect 1007 407 1008 411
rect 1002 406 1008 407
rect 1004 386 1006 406
rect 1002 385 1008 386
rect 1002 381 1003 385
rect 1007 381 1008 385
rect 1002 380 1008 381
rect 1112 380 1114 429
rect 1226 411 1232 412
rect 1226 407 1227 411
rect 1231 407 1232 411
rect 1226 406 1232 407
rect 1190 403 1196 404
rect 1190 399 1191 403
rect 1195 399 1196 403
rect 1190 398 1196 399
rect 110 376 116 377
rect 198 379 204 380
rect 198 375 199 379
rect 203 375 204 379
rect 198 374 204 375
rect 430 379 436 380
rect 430 375 431 379
rect 435 375 436 379
rect 430 374 436 375
rect 662 379 668 380
rect 662 375 663 379
rect 667 375 668 379
rect 662 374 668 375
rect 222 364 228 365
rect 110 363 116 364
rect 110 359 111 363
rect 115 359 116 363
rect 222 360 223 364
rect 227 360 228 364
rect 222 359 228 360
rect 454 364 460 365
rect 454 360 455 364
rect 459 360 460 364
rect 454 359 460 360
rect 686 364 692 365
rect 686 360 687 364
rect 691 360 692 364
rect 686 359 692 360
rect 110 358 116 359
rect 112 323 114 358
rect 224 323 226 359
rect 456 323 458 359
rect 688 323 690 359
rect 111 322 115 323
rect 111 317 115 318
rect 223 322 227 323
rect 223 317 227 318
rect 439 322 443 323
rect 439 317 443 318
rect 455 322 459 323
rect 455 317 459 318
rect 655 322 659 323
rect 655 317 659 318
rect 687 322 691 323
rect 687 317 691 318
rect 112 294 114 317
rect 110 293 116 294
rect 440 293 442 317
rect 656 293 658 317
rect 110 289 111 293
rect 115 289 116 293
rect 110 288 116 289
rect 438 292 444 293
rect 438 288 439 292
rect 443 288 444 292
rect 438 287 444 288
rect 654 292 660 293
rect 654 288 655 292
rect 659 288 660 292
rect 654 287 660 288
rect 414 277 420 278
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 414 273 415 277
rect 419 273 420 277
rect 414 272 420 273
rect 630 277 636 278
rect 630 273 631 277
rect 635 273 636 277
rect 630 272 636 273
rect 110 270 116 271
rect 112 211 114 270
rect 416 211 418 272
rect 510 271 516 272
rect 510 267 511 271
rect 515 267 516 271
rect 510 266 516 267
rect 574 271 580 272
rect 574 267 575 271
rect 579 267 580 271
rect 574 266 580 267
rect 111 210 115 211
rect 111 205 115 206
rect 415 210 419 211
rect 415 205 419 206
rect 487 210 491 211
rect 487 205 491 206
rect 112 158 114 205
rect 110 157 116 158
rect 110 153 111 157
rect 115 153 116 157
rect 488 156 490 205
rect 512 188 514 266
rect 576 244 578 266
rect 574 243 580 244
rect 574 239 575 243
rect 579 239 580 243
rect 574 238 580 239
rect 632 211 634 272
rect 754 271 760 272
rect 754 267 755 271
rect 759 267 760 271
rect 754 266 760 267
rect 756 244 758 266
rect 764 244 766 380
rect 886 379 892 380
rect 886 375 887 379
rect 891 375 892 379
rect 886 374 892 375
rect 1110 379 1116 380
rect 1110 375 1111 379
rect 1115 375 1116 379
rect 1110 374 1116 375
rect 910 364 916 365
rect 910 360 911 364
rect 915 360 916 364
rect 910 359 916 360
rect 1134 364 1140 365
rect 1134 360 1135 364
rect 1139 360 1140 364
rect 1134 359 1140 360
rect 912 323 914 359
rect 1136 323 1138 359
rect 879 322 883 323
rect 879 317 883 318
rect 911 322 915 323
rect 911 317 915 318
rect 1119 322 1123 323
rect 1119 317 1123 318
rect 1135 322 1139 323
rect 1135 317 1139 318
rect 880 293 882 317
rect 1120 293 1122 317
rect 878 292 884 293
rect 878 288 879 292
rect 883 288 884 292
rect 878 287 884 288
rect 1118 292 1124 293
rect 1118 288 1119 292
rect 1123 288 1124 292
rect 1118 287 1124 288
rect 854 277 860 278
rect 854 273 855 277
rect 859 273 860 277
rect 854 272 860 273
rect 1094 277 1100 278
rect 1094 273 1095 277
rect 1099 273 1100 277
rect 1094 272 1100 273
rect 1192 272 1194 398
rect 1228 386 1230 406
rect 1226 385 1232 386
rect 1226 381 1227 385
rect 1231 381 1232 385
rect 1226 380 1232 381
rect 1336 380 1338 429
rect 1416 386 1418 466
rect 1544 435 1546 500
rect 1620 472 1622 706
rect 1656 684 1658 824
rect 1718 821 1719 825
rect 1723 821 1724 825
rect 1718 820 1724 821
rect 1718 807 1724 808
rect 1718 803 1719 807
rect 1723 803 1724 807
rect 1718 802 1724 803
rect 1720 763 1722 802
rect 1719 762 1723 763
rect 1719 757 1723 758
rect 1720 734 1722 757
rect 1718 733 1724 734
rect 1718 729 1719 733
rect 1723 729 1724 733
rect 1718 728 1724 729
rect 1718 715 1724 716
rect 1718 711 1719 715
rect 1723 711 1724 715
rect 1718 710 1724 711
rect 1654 683 1660 684
rect 1654 679 1655 683
rect 1659 679 1660 683
rect 1654 678 1660 679
rect 1720 663 1722 710
rect 1719 662 1723 663
rect 1719 657 1723 658
rect 1720 610 1722 657
rect 1718 609 1724 610
rect 1718 605 1719 609
rect 1723 605 1724 609
rect 1718 604 1724 605
rect 1718 591 1724 592
rect 1718 587 1719 591
rect 1723 587 1724 591
rect 1718 586 1724 587
rect 1720 551 1722 586
rect 1719 550 1723 551
rect 1719 545 1723 546
rect 1720 522 1722 545
rect 1718 521 1724 522
rect 1718 517 1719 521
rect 1723 517 1724 521
rect 1718 516 1724 517
rect 1718 503 1724 504
rect 1634 499 1640 500
rect 1634 495 1635 499
rect 1639 495 1640 499
rect 1718 499 1719 503
rect 1723 499 1724 503
rect 1718 498 1724 499
rect 1634 494 1640 495
rect 1618 471 1624 472
rect 1618 467 1619 471
rect 1623 467 1624 471
rect 1618 466 1624 467
rect 1543 434 1547 435
rect 1543 429 1547 430
rect 1559 434 1563 435
rect 1559 429 1563 430
rect 1414 385 1420 386
rect 1414 381 1415 385
rect 1419 381 1420 385
rect 1414 380 1420 381
rect 1560 380 1562 429
rect 1636 412 1638 494
rect 1720 435 1722 498
rect 1719 434 1723 435
rect 1719 429 1723 430
rect 1634 411 1640 412
rect 1634 407 1635 411
rect 1639 407 1640 411
rect 1634 406 1640 407
rect 1650 385 1656 386
rect 1650 381 1651 385
rect 1655 381 1656 385
rect 1720 382 1722 429
rect 1650 380 1656 381
rect 1718 381 1724 382
rect 1334 379 1340 380
rect 1334 375 1335 379
rect 1339 375 1340 379
rect 1334 374 1340 375
rect 1558 379 1564 380
rect 1558 375 1559 379
rect 1563 375 1564 379
rect 1558 374 1564 375
rect 1358 364 1364 365
rect 1358 360 1359 364
rect 1363 360 1364 364
rect 1358 359 1364 360
rect 1582 364 1588 365
rect 1582 360 1583 364
rect 1587 360 1588 364
rect 1582 359 1588 360
rect 1360 323 1362 359
rect 1584 323 1586 359
rect 1359 322 1363 323
rect 1359 317 1363 318
rect 1367 322 1371 323
rect 1367 317 1371 318
rect 1583 322 1587 323
rect 1583 317 1587 318
rect 1599 322 1603 323
rect 1599 317 1603 318
rect 1368 293 1370 317
rect 1600 293 1602 317
rect 1366 292 1372 293
rect 1366 288 1367 292
rect 1371 288 1372 292
rect 1366 287 1372 288
rect 1598 292 1604 293
rect 1598 288 1599 292
rect 1603 288 1604 292
rect 1598 287 1604 288
rect 1342 277 1348 278
rect 1342 273 1343 277
rect 1347 273 1348 277
rect 1342 272 1348 273
rect 1574 277 1580 278
rect 1574 273 1575 277
rect 1579 273 1580 277
rect 1574 272 1580 273
rect 754 243 760 244
rect 754 239 755 243
rect 759 239 760 243
rect 754 238 760 239
rect 762 243 768 244
rect 762 239 763 243
rect 767 239 768 243
rect 762 238 768 239
rect 856 211 858 272
rect 1096 211 1098 272
rect 1190 271 1196 272
rect 1190 267 1191 271
rect 1195 267 1196 271
rect 1190 266 1196 267
rect 1298 271 1304 272
rect 1298 267 1299 271
rect 1303 267 1304 271
rect 1298 266 1304 267
rect 1300 244 1302 266
rect 1298 243 1304 244
rect 1298 239 1299 243
rect 1303 239 1304 243
rect 1298 238 1304 239
rect 1344 211 1346 272
rect 1398 243 1404 244
rect 1398 239 1399 243
rect 1403 239 1404 243
rect 1398 238 1404 239
rect 623 210 627 211
rect 623 205 627 206
rect 631 210 635 211
rect 631 205 635 206
rect 759 210 763 211
rect 759 205 763 206
rect 855 210 859 211
rect 855 205 859 206
rect 895 210 899 211
rect 895 205 899 206
rect 1031 210 1035 211
rect 1031 205 1035 206
rect 1095 210 1099 211
rect 1095 205 1099 206
rect 1167 210 1171 211
rect 1167 205 1171 206
rect 1303 210 1307 211
rect 1303 205 1307 206
rect 1343 210 1347 211
rect 1343 205 1347 206
rect 510 187 516 188
rect 510 183 511 187
rect 515 183 516 187
rect 510 182 516 183
rect 602 187 608 188
rect 602 183 603 187
rect 607 183 608 187
rect 602 182 608 183
rect 604 162 606 182
rect 602 161 608 162
rect 602 157 603 161
rect 607 157 608 161
rect 602 156 608 157
rect 624 156 626 205
rect 738 187 744 188
rect 738 183 739 187
rect 743 183 744 187
rect 738 182 744 183
rect 740 162 742 182
rect 738 161 744 162
rect 738 157 739 161
rect 743 157 744 161
rect 738 156 744 157
rect 760 156 762 205
rect 874 187 880 188
rect 874 183 875 187
rect 879 183 880 187
rect 874 182 880 183
rect 876 162 878 182
rect 874 161 880 162
rect 874 157 875 161
rect 879 157 880 161
rect 874 156 880 157
rect 896 156 898 205
rect 1010 187 1016 188
rect 1010 183 1011 187
rect 1015 183 1016 187
rect 1010 182 1016 183
rect 1012 162 1014 182
rect 1010 161 1016 162
rect 1010 157 1011 161
rect 1015 157 1016 161
rect 1010 156 1016 157
rect 1032 156 1034 205
rect 1146 187 1152 188
rect 1146 183 1147 187
rect 1151 183 1152 187
rect 1146 182 1152 183
rect 1148 162 1150 182
rect 1146 161 1152 162
rect 1146 157 1147 161
rect 1151 157 1152 161
rect 1146 156 1152 157
rect 1168 156 1170 205
rect 1266 187 1272 188
rect 1266 183 1267 187
rect 1271 183 1272 187
rect 1266 182 1272 183
rect 1268 162 1270 182
rect 1266 161 1272 162
rect 1266 157 1267 161
rect 1271 157 1272 161
rect 1266 156 1272 157
rect 1304 156 1306 205
rect 1400 162 1402 238
rect 1576 211 1578 272
rect 1652 244 1654 380
rect 1718 377 1719 381
rect 1723 377 1724 381
rect 1718 376 1724 377
rect 1718 363 1724 364
rect 1718 359 1719 363
rect 1723 359 1724 363
rect 1718 358 1724 359
rect 1720 323 1722 358
rect 1719 322 1723 323
rect 1719 317 1723 318
rect 1720 294 1722 317
rect 1718 293 1724 294
rect 1718 289 1719 293
rect 1723 289 1724 293
rect 1718 288 1724 289
rect 1718 275 1724 276
rect 1666 271 1672 272
rect 1666 267 1667 271
rect 1671 267 1672 271
rect 1718 271 1719 275
rect 1723 271 1724 275
rect 1718 270 1724 271
rect 1666 266 1672 267
rect 1650 243 1656 244
rect 1650 239 1651 243
rect 1655 239 1656 243
rect 1650 238 1656 239
rect 1439 210 1443 211
rect 1439 205 1443 206
rect 1575 210 1579 211
rect 1575 205 1579 206
rect 1398 161 1404 162
rect 1398 157 1399 161
rect 1403 157 1404 161
rect 1398 156 1404 157
rect 1440 156 1442 205
rect 1514 187 1520 188
rect 1514 183 1515 187
rect 1519 183 1520 187
rect 1514 182 1520 183
rect 1516 164 1518 182
rect 1514 163 1520 164
rect 1514 159 1515 163
rect 1519 159 1520 163
rect 1514 158 1520 159
rect 1576 156 1578 205
rect 1668 192 1670 266
rect 1720 211 1722 270
rect 1719 210 1723 211
rect 1719 205 1723 206
rect 1666 191 1672 192
rect 1666 187 1667 191
rect 1671 187 1672 191
rect 1666 186 1672 187
rect 1720 158 1722 205
rect 1718 157 1724 158
rect 110 152 116 153
rect 486 155 492 156
rect 486 151 487 155
rect 491 151 492 155
rect 486 150 492 151
rect 622 155 628 156
rect 622 151 623 155
rect 627 151 628 155
rect 622 150 628 151
rect 758 155 764 156
rect 758 151 759 155
rect 763 151 764 155
rect 758 150 764 151
rect 894 155 900 156
rect 894 151 895 155
rect 899 151 900 155
rect 894 150 900 151
rect 1030 155 1036 156
rect 1030 151 1031 155
rect 1035 151 1036 155
rect 1030 150 1036 151
rect 1166 155 1172 156
rect 1166 151 1167 155
rect 1171 151 1172 155
rect 1166 150 1172 151
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1302 150 1308 151
rect 1438 155 1444 156
rect 1438 151 1439 155
rect 1443 151 1444 155
rect 1438 150 1444 151
rect 1574 155 1580 156
rect 1574 151 1575 155
rect 1579 151 1580 155
rect 1718 153 1719 157
rect 1723 153 1724 157
rect 1718 152 1724 153
rect 1574 150 1580 151
rect 510 140 516 141
rect 110 139 116 140
rect 110 135 111 139
rect 115 135 116 139
rect 510 136 511 140
rect 515 136 516 140
rect 510 135 516 136
rect 646 140 652 141
rect 646 136 647 140
rect 651 136 652 140
rect 646 135 652 136
rect 782 140 788 141
rect 782 136 783 140
rect 787 136 788 140
rect 782 135 788 136
rect 918 140 924 141
rect 918 136 919 140
rect 923 136 924 140
rect 918 135 924 136
rect 1054 140 1060 141
rect 1054 136 1055 140
rect 1059 136 1060 140
rect 1054 135 1060 136
rect 1190 140 1196 141
rect 1190 136 1191 140
rect 1195 136 1196 140
rect 1190 135 1196 136
rect 1326 140 1332 141
rect 1326 136 1327 140
rect 1331 136 1332 140
rect 1326 135 1332 136
rect 1462 140 1468 141
rect 1462 136 1463 140
rect 1467 136 1468 140
rect 1462 135 1468 136
rect 1598 140 1604 141
rect 1598 136 1599 140
rect 1603 136 1604 140
rect 1598 135 1604 136
rect 1718 139 1724 140
rect 1718 135 1719 139
rect 1723 135 1724 139
rect 110 134 116 135
rect 112 111 114 134
rect 512 111 514 135
rect 648 111 650 135
rect 784 111 786 135
rect 920 111 922 135
rect 1056 111 1058 135
rect 1192 111 1194 135
rect 1328 111 1330 135
rect 1464 111 1466 135
rect 1600 111 1602 135
rect 1718 134 1724 135
rect 1720 111 1722 134
rect 111 110 115 111
rect 111 105 115 106
rect 511 110 515 111
rect 511 105 515 106
rect 647 110 651 111
rect 647 105 651 106
rect 783 110 787 111
rect 783 105 787 106
rect 919 110 923 111
rect 919 105 923 106
rect 1055 110 1059 111
rect 1055 105 1059 106
rect 1191 110 1195 111
rect 1191 105 1195 106
rect 1327 110 1331 111
rect 1327 105 1331 106
rect 1463 110 1467 111
rect 1463 105 1467 106
rect 1599 110 1603 111
rect 1599 105 1603 106
rect 1719 110 1723 111
rect 1719 105 1723 106
<< m4c >>
rect 111 1778 115 1782
rect 135 1778 139 1782
rect 271 1778 275 1782
rect 407 1778 411 1782
rect 543 1778 547 1782
rect 679 1778 683 1782
rect 1719 1778 1723 1782
rect 111 1666 115 1670
rect 159 1666 163 1670
rect 231 1666 235 1670
rect 295 1666 299 1670
rect 367 1666 371 1670
rect 431 1666 435 1670
rect 503 1666 507 1670
rect 567 1666 571 1670
rect 639 1666 643 1670
rect 703 1666 707 1670
rect 111 1554 115 1558
rect 207 1554 211 1558
rect 343 1554 347 1558
rect 479 1554 483 1558
rect 487 1554 491 1558
rect 775 1666 779 1670
rect 1719 1666 1723 1670
rect 615 1554 619 1558
rect 623 1554 627 1558
rect 751 1554 755 1558
rect 759 1554 763 1558
rect 895 1554 899 1558
rect 1031 1554 1035 1558
rect 1167 1554 1171 1558
rect 1303 1554 1307 1558
rect 1439 1554 1443 1558
rect 1575 1554 1579 1558
rect 1719 1554 1723 1558
rect 111 1438 115 1442
rect 511 1438 515 1442
rect 623 1438 627 1442
rect 647 1438 651 1442
rect 759 1438 763 1442
rect 783 1438 787 1442
rect 895 1438 899 1442
rect 919 1438 923 1442
rect 1039 1438 1043 1442
rect 1055 1438 1059 1442
rect 1183 1438 1187 1442
rect 1191 1438 1195 1442
rect 1327 1438 1331 1442
rect 1463 1438 1467 1442
rect 1599 1438 1603 1442
rect 1719 1438 1723 1442
rect 111 1322 115 1326
rect 135 1322 139 1326
rect 343 1322 347 1326
rect 599 1322 603 1326
rect 607 1322 611 1326
rect 735 1322 739 1326
rect 871 1322 875 1326
rect 895 1322 899 1326
rect 1015 1322 1019 1326
rect 1159 1322 1163 1326
rect 1207 1322 1211 1326
rect 1303 1322 1307 1326
rect 111 1210 115 1214
rect 159 1210 163 1214
rect 327 1210 331 1214
rect 367 1210 371 1214
rect 543 1210 547 1214
rect 631 1210 635 1214
rect 775 1210 779 1214
rect 919 1210 923 1214
rect 1023 1210 1027 1214
rect 1231 1210 1235 1214
rect 1287 1210 1291 1214
rect 1439 1322 1443 1326
rect 1519 1322 1523 1326
rect 1575 1322 1579 1326
rect 1719 1322 1723 1326
rect 1543 1210 1547 1214
rect 1551 1210 1555 1214
rect 111 1090 115 1094
rect 135 1090 139 1094
rect 303 1090 307 1094
rect 311 1090 315 1094
rect 519 1090 523 1094
rect 535 1090 539 1094
rect 751 1090 755 1094
rect 775 1090 779 1094
rect 999 1090 1003 1094
rect 1023 1090 1027 1094
rect 1263 1090 1267 1094
rect 1279 1090 1283 1094
rect 1719 1210 1723 1214
rect 1527 1090 1531 1094
rect 1543 1090 1547 1094
rect 111 990 115 994
rect 335 990 339 994
rect 527 990 531 994
rect 559 990 563 994
rect 711 990 715 994
rect 799 990 803 994
rect 919 990 923 994
rect 1047 990 1051 994
rect 111 874 115 878
rect 503 874 507 878
rect 687 874 691 878
rect 743 874 747 878
rect 1135 990 1139 994
rect 1303 990 1307 994
rect 1367 990 1371 994
rect 879 874 883 878
rect 895 874 899 878
rect 1015 874 1019 878
rect 1111 874 1115 878
rect 1151 874 1155 878
rect 1287 874 1291 878
rect 1343 874 1347 878
rect 1431 874 1435 878
rect 111 758 115 762
rect 703 758 707 762
rect 767 758 771 762
rect 863 758 867 762
rect 903 758 907 762
rect 1031 758 1035 762
rect 1039 758 1043 762
rect 1175 758 1179 762
rect 1215 758 1219 762
rect 1311 758 1315 762
rect 111 658 115 662
rect 223 658 227 662
rect 415 658 419 662
rect 623 658 627 662
rect 679 658 683 662
rect 839 658 843 662
rect 855 658 859 662
rect 1007 658 1011 662
rect 1095 658 1099 662
rect 111 546 115 550
rect 159 546 163 550
rect 1399 758 1403 762
rect 1191 658 1195 662
rect 1335 658 1339 662
rect 1375 658 1379 662
rect 247 546 251 550
rect 327 546 331 550
rect 439 546 443 550
rect 543 546 547 550
rect 647 546 651 550
rect 783 546 787 550
rect 879 546 883 550
rect 1039 546 1043 550
rect 1119 546 1123 550
rect 1303 546 1307 550
rect 1359 546 1363 550
rect 1719 1090 1723 1094
rect 1567 990 1571 994
rect 1599 990 1603 994
rect 1719 990 1723 994
rect 1575 874 1579 878
rect 1719 874 1723 878
rect 1455 758 1459 762
rect 1591 758 1595 762
rect 1599 758 1603 762
rect 1567 658 1571 662
rect 1567 546 1571 550
rect 111 430 115 434
rect 135 430 139 434
rect 199 430 203 434
rect 303 430 307 434
rect 431 430 435 434
rect 519 430 523 434
rect 663 430 667 434
rect 759 430 763 434
rect 887 430 891 434
rect 1015 430 1019 434
rect 1111 430 1115 434
rect 1279 430 1283 434
rect 1335 430 1339 434
rect 111 318 115 322
rect 223 318 227 322
rect 439 318 443 322
rect 455 318 459 322
rect 655 318 659 322
rect 687 318 691 322
rect 111 206 115 210
rect 415 206 419 210
rect 487 206 491 210
rect 879 318 883 322
rect 911 318 915 322
rect 1119 318 1123 322
rect 1135 318 1139 322
rect 1719 758 1723 762
rect 1719 658 1723 662
rect 1719 546 1723 550
rect 1543 430 1547 434
rect 1559 430 1563 434
rect 1719 430 1723 434
rect 1359 318 1363 322
rect 1367 318 1371 322
rect 1583 318 1587 322
rect 1599 318 1603 322
rect 623 206 627 210
rect 631 206 635 210
rect 759 206 763 210
rect 855 206 859 210
rect 895 206 899 210
rect 1031 206 1035 210
rect 1095 206 1099 210
rect 1167 206 1171 210
rect 1303 206 1307 210
rect 1343 206 1347 210
rect 1719 318 1723 322
rect 1439 206 1443 210
rect 1575 206 1579 210
rect 1719 206 1723 210
rect 111 106 115 110
rect 511 106 515 110
rect 647 106 651 110
rect 783 106 787 110
rect 919 106 923 110
rect 1055 106 1059 110
rect 1191 106 1195 110
rect 1327 106 1331 110
rect 1463 106 1467 110
rect 1599 106 1603 110
rect 1719 106 1723 110
<< m4 >>
rect 96 1777 97 1783
rect 103 1782 1755 1783
rect 103 1778 111 1782
rect 115 1778 135 1782
rect 139 1778 271 1782
rect 275 1778 407 1782
rect 411 1778 543 1782
rect 547 1778 679 1782
rect 683 1778 1719 1782
rect 1723 1778 1755 1782
rect 103 1777 1755 1778
rect 1761 1777 1762 1783
rect 84 1665 85 1671
rect 91 1670 1743 1671
rect 91 1666 111 1670
rect 115 1666 159 1670
rect 163 1666 231 1670
rect 235 1666 295 1670
rect 299 1666 367 1670
rect 371 1666 431 1670
rect 435 1666 503 1670
rect 507 1666 567 1670
rect 571 1666 639 1670
rect 643 1666 703 1670
rect 707 1666 775 1670
rect 779 1666 1719 1670
rect 1723 1666 1743 1670
rect 91 1665 1743 1666
rect 1749 1665 1750 1671
rect 96 1553 97 1559
rect 103 1558 1755 1559
rect 103 1554 111 1558
rect 115 1554 207 1558
rect 211 1554 343 1558
rect 347 1554 479 1558
rect 483 1554 487 1558
rect 491 1554 615 1558
rect 619 1554 623 1558
rect 627 1554 751 1558
rect 755 1554 759 1558
rect 763 1554 895 1558
rect 899 1554 1031 1558
rect 1035 1554 1167 1558
rect 1171 1554 1303 1558
rect 1307 1554 1439 1558
rect 1443 1554 1575 1558
rect 1579 1554 1719 1558
rect 1723 1554 1755 1558
rect 103 1553 1755 1554
rect 1761 1553 1762 1559
rect 84 1437 85 1443
rect 91 1442 1743 1443
rect 91 1438 111 1442
rect 115 1438 511 1442
rect 515 1438 623 1442
rect 627 1438 647 1442
rect 651 1438 759 1442
rect 763 1438 783 1442
rect 787 1438 895 1442
rect 899 1438 919 1442
rect 923 1438 1039 1442
rect 1043 1438 1055 1442
rect 1059 1438 1183 1442
rect 1187 1438 1191 1442
rect 1195 1438 1327 1442
rect 1331 1438 1463 1442
rect 1467 1438 1599 1442
rect 1603 1438 1719 1442
rect 1723 1438 1743 1442
rect 91 1437 1743 1438
rect 1749 1437 1750 1443
rect 96 1321 97 1327
rect 103 1326 1755 1327
rect 103 1322 111 1326
rect 115 1322 135 1326
rect 139 1322 343 1326
rect 347 1322 599 1326
rect 603 1322 607 1326
rect 611 1322 735 1326
rect 739 1322 871 1326
rect 875 1322 895 1326
rect 899 1322 1015 1326
rect 1019 1322 1159 1326
rect 1163 1322 1207 1326
rect 1211 1322 1303 1326
rect 1307 1322 1439 1326
rect 1443 1322 1519 1326
rect 1523 1322 1575 1326
rect 1579 1322 1719 1326
rect 1723 1322 1755 1326
rect 103 1321 1755 1322
rect 1761 1321 1762 1327
rect 84 1209 85 1215
rect 91 1214 1743 1215
rect 91 1210 111 1214
rect 115 1210 159 1214
rect 163 1210 327 1214
rect 331 1210 367 1214
rect 371 1210 543 1214
rect 547 1210 631 1214
rect 635 1210 775 1214
rect 779 1210 919 1214
rect 923 1210 1023 1214
rect 1027 1210 1231 1214
rect 1235 1210 1287 1214
rect 1291 1210 1543 1214
rect 1547 1210 1551 1214
rect 1555 1210 1719 1214
rect 1723 1210 1743 1214
rect 91 1209 1743 1210
rect 1749 1209 1750 1215
rect 96 1089 97 1095
rect 103 1094 1755 1095
rect 103 1090 111 1094
rect 115 1090 135 1094
rect 139 1090 303 1094
rect 307 1090 311 1094
rect 315 1090 519 1094
rect 523 1090 535 1094
rect 539 1090 751 1094
rect 755 1090 775 1094
rect 779 1090 999 1094
rect 1003 1090 1023 1094
rect 1027 1090 1263 1094
rect 1267 1090 1279 1094
rect 1283 1090 1527 1094
rect 1531 1090 1543 1094
rect 1547 1090 1719 1094
rect 1723 1090 1755 1094
rect 103 1089 1755 1090
rect 1761 1089 1762 1095
rect 84 989 85 995
rect 91 994 1743 995
rect 91 990 111 994
rect 115 990 335 994
rect 339 990 527 994
rect 531 990 559 994
rect 563 990 711 994
rect 715 990 799 994
rect 803 990 919 994
rect 923 990 1047 994
rect 1051 990 1135 994
rect 1139 990 1303 994
rect 1307 990 1367 994
rect 1371 990 1567 994
rect 1571 990 1599 994
rect 1603 990 1719 994
rect 1723 990 1743 994
rect 91 989 1743 990
rect 1749 989 1750 995
rect 96 873 97 879
rect 103 878 1755 879
rect 103 874 111 878
rect 115 874 503 878
rect 507 874 687 878
rect 691 874 743 878
rect 747 874 879 878
rect 883 874 895 878
rect 899 874 1015 878
rect 1019 874 1111 878
rect 1115 874 1151 878
rect 1155 874 1287 878
rect 1291 874 1343 878
rect 1347 874 1431 878
rect 1435 874 1575 878
rect 1579 874 1719 878
rect 1723 874 1755 878
rect 103 873 1755 874
rect 1761 873 1762 879
rect 84 757 85 763
rect 91 762 1743 763
rect 91 758 111 762
rect 115 758 703 762
rect 707 758 767 762
rect 771 758 863 762
rect 867 758 903 762
rect 907 758 1031 762
rect 1035 758 1039 762
rect 1043 758 1175 762
rect 1179 758 1215 762
rect 1219 758 1311 762
rect 1315 758 1399 762
rect 1403 758 1455 762
rect 1459 758 1591 762
rect 1595 758 1599 762
rect 1603 758 1719 762
rect 1723 758 1743 762
rect 91 757 1743 758
rect 1749 757 1750 763
rect 96 657 97 663
rect 103 662 1755 663
rect 103 658 111 662
rect 115 658 223 662
rect 227 658 415 662
rect 419 658 623 662
rect 627 658 679 662
rect 683 658 839 662
rect 843 658 855 662
rect 859 658 1007 662
rect 1011 658 1095 662
rect 1099 658 1191 662
rect 1195 658 1335 662
rect 1339 658 1375 662
rect 1379 658 1567 662
rect 1571 658 1719 662
rect 1723 658 1755 662
rect 103 657 1755 658
rect 1761 657 1762 663
rect 84 545 85 551
rect 91 550 1743 551
rect 91 546 111 550
rect 115 546 159 550
rect 163 546 247 550
rect 251 546 327 550
rect 331 546 439 550
rect 443 546 543 550
rect 547 546 647 550
rect 651 546 783 550
rect 787 546 879 550
rect 883 546 1039 550
rect 1043 546 1119 550
rect 1123 546 1303 550
rect 1307 546 1359 550
rect 1363 546 1567 550
rect 1571 546 1719 550
rect 1723 546 1743 550
rect 91 545 1743 546
rect 1749 545 1750 551
rect 96 429 97 435
rect 103 434 1755 435
rect 103 430 111 434
rect 115 430 135 434
rect 139 430 199 434
rect 203 430 303 434
rect 307 430 431 434
rect 435 430 519 434
rect 523 430 663 434
rect 667 430 759 434
rect 763 430 887 434
rect 891 430 1015 434
rect 1019 430 1111 434
rect 1115 430 1279 434
rect 1283 430 1335 434
rect 1339 430 1543 434
rect 1547 430 1559 434
rect 1563 430 1719 434
rect 1723 430 1755 434
rect 103 429 1755 430
rect 1761 429 1762 435
rect 84 317 85 323
rect 91 322 1743 323
rect 91 318 111 322
rect 115 318 223 322
rect 227 318 439 322
rect 443 318 455 322
rect 459 318 655 322
rect 659 318 687 322
rect 691 318 879 322
rect 883 318 911 322
rect 915 318 1119 322
rect 1123 318 1135 322
rect 1139 318 1359 322
rect 1363 318 1367 322
rect 1371 318 1583 322
rect 1587 318 1599 322
rect 1603 318 1719 322
rect 1723 318 1743 322
rect 91 317 1743 318
rect 1749 317 1750 323
rect 96 205 97 211
rect 103 210 1755 211
rect 103 206 111 210
rect 115 206 415 210
rect 419 206 487 210
rect 491 206 623 210
rect 627 206 631 210
rect 635 206 759 210
rect 763 206 855 210
rect 859 206 895 210
rect 899 206 1031 210
rect 1035 206 1095 210
rect 1099 206 1167 210
rect 1171 206 1303 210
rect 1307 206 1343 210
rect 1347 206 1439 210
rect 1443 206 1575 210
rect 1579 206 1719 210
rect 1723 206 1755 210
rect 103 205 1755 206
rect 1761 205 1762 211
rect 84 105 85 111
rect 91 110 1743 111
rect 91 106 111 110
rect 115 106 511 110
rect 515 106 647 110
rect 651 106 783 110
rect 787 106 919 110
rect 923 106 1055 110
rect 1059 106 1191 110
rect 1195 106 1327 110
rect 1331 106 1463 110
rect 1467 106 1599 110
rect 1603 106 1719 110
rect 1723 106 1743 110
rect 91 105 1743 106
rect 1749 105 1750 111
<< m5c >>
rect 97 1777 103 1783
rect 1755 1777 1761 1783
rect 85 1665 91 1671
rect 1743 1665 1749 1671
rect 97 1553 103 1559
rect 1755 1553 1761 1559
rect 85 1437 91 1443
rect 1743 1437 1749 1443
rect 97 1321 103 1327
rect 1755 1321 1761 1327
rect 85 1209 91 1215
rect 1743 1209 1749 1215
rect 97 1089 103 1095
rect 1755 1089 1761 1095
rect 85 989 91 995
rect 1743 989 1749 995
rect 97 873 103 879
rect 1755 873 1761 879
rect 85 757 91 763
rect 1743 757 1749 763
rect 97 657 103 663
rect 1755 657 1761 663
rect 85 545 91 551
rect 1743 545 1749 551
rect 97 429 103 435
rect 1755 429 1761 435
rect 85 317 91 323
rect 1743 317 1749 323
rect 97 205 103 211
rect 1755 205 1761 211
rect 85 105 91 111
rect 1743 105 1749 111
<< m5 >>
rect 84 1671 92 1800
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1443 92 1665
rect 84 1437 85 1443
rect 91 1437 92 1443
rect 84 1215 92 1437
rect 84 1209 85 1215
rect 91 1209 92 1215
rect 84 995 92 1209
rect 84 989 85 995
rect 91 989 92 995
rect 84 763 92 989
rect 84 757 85 763
rect 91 757 92 763
rect 84 551 92 757
rect 84 545 85 551
rect 91 545 92 551
rect 84 323 92 545
rect 84 317 85 323
rect 91 317 92 323
rect 84 111 92 317
rect 84 105 85 111
rect 91 105 92 111
rect 84 72 92 105
rect 96 1783 104 1800
rect 96 1777 97 1783
rect 103 1777 104 1783
rect 96 1559 104 1777
rect 96 1553 97 1559
rect 103 1553 104 1559
rect 96 1327 104 1553
rect 96 1321 97 1327
rect 103 1321 104 1327
rect 96 1095 104 1321
rect 96 1089 97 1095
rect 103 1089 104 1095
rect 96 879 104 1089
rect 96 873 97 879
rect 103 873 104 879
rect 96 663 104 873
rect 96 657 97 663
rect 103 657 104 663
rect 96 435 104 657
rect 96 429 97 435
rect 103 429 104 435
rect 96 211 104 429
rect 96 205 97 211
rect 103 205 104 211
rect 96 72 104 205
rect 1742 1671 1750 1800
rect 1742 1665 1743 1671
rect 1749 1665 1750 1671
rect 1742 1443 1750 1665
rect 1742 1437 1743 1443
rect 1749 1437 1750 1443
rect 1742 1215 1750 1437
rect 1742 1209 1743 1215
rect 1749 1209 1750 1215
rect 1742 995 1750 1209
rect 1742 989 1743 995
rect 1749 989 1750 995
rect 1742 763 1750 989
rect 1742 757 1743 763
rect 1749 757 1750 763
rect 1742 551 1750 757
rect 1742 545 1743 551
rect 1749 545 1750 551
rect 1742 323 1750 545
rect 1742 317 1743 323
rect 1749 317 1750 323
rect 1742 111 1750 317
rect 1742 105 1743 111
rect 1749 105 1750 111
rect 1742 72 1750 105
rect 1754 1783 1762 1800
rect 1754 1777 1755 1783
rect 1761 1777 1762 1783
rect 1754 1559 1762 1777
rect 1754 1553 1755 1559
rect 1761 1553 1762 1559
rect 1754 1327 1762 1553
rect 1754 1321 1755 1327
rect 1761 1321 1762 1327
rect 1754 1095 1762 1321
rect 1754 1089 1755 1095
rect 1761 1089 1762 1095
rect 1754 879 1762 1089
rect 1754 873 1755 879
rect 1761 873 1762 879
rect 1754 663 1762 873
rect 1754 657 1755 663
rect 1761 657 1762 663
rect 1754 435 1762 657
rect 1754 429 1755 435
rect 1761 429 1762 435
rect 1754 211 1762 429
rect 1754 205 1755 211
rect 1761 205 1762 211
rect 1754 72 1762 205
use welltap_svt  __well_tap__0
timestamp 1730768468
transform 1 0 104 0 1 132
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730768468
transform 1 0 104 0 1 132
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768468
transform 1 0 480 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768468
transform 1 0 480 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768468
transform 1 0 616 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768468
transform 1 0 616 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768468
transform 1 0 752 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768468
transform 1 0 752 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768468
transform 1 0 888 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768468
transform 1 0 888 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768468
transform 1 0 1024 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768468
transform 1 0 1024 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768468
transform 1 0 1160 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768468
transform 1 0 1160 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768468
transform 1 0 1296 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768468
transform 1 0 1296 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768468
transform 1 0 1432 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768468
transform 1 0 1432 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768468
transform 1 0 1568 0 1 108
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768468
transform 1 0 1568 0 1 108
box 8 5 126 98
use welltap_svt  __well_tap__1
timestamp 1730768468
transform 1 0 1712 0 1 132
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730768468
transform 1 0 1712 0 1 132
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768468
transform 1 0 408 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768468
transform 1 0 408 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768468
transform 1 0 624 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768468
transform 1 0 624 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768468
transform 1 0 848 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768468
transform 1 0 848 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768468
transform 1 0 1088 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768468
transform 1 0 1088 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768468
transform 1 0 1336 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768468
transform 1 0 1336 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768468
transform 1 0 1568 0 -1 320
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768468
transform 1 0 1568 0 -1 320
box 8 5 126 98
use welltap_svt  __well_tap__2
timestamp 1730768468
transform 1 0 104 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730768468
transform 1 0 104 0 -1 296
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768468
transform 1 0 192 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768468
transform 1 0 192 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768468
transform 1 0 424 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768468
transform 1 0 424 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768468
transform 1 0 656 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768468
transform 1 0 656 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768468
transform 1 0 880 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768468
transform 1 0 880 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768468
transform 1 0 1104 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768468
transform 1 0 1104 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768468
transform 1 0 1328 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768468
transform 1 0 1328 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768468
transform 1 0 1552 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768468
transform 1 0 1552 0 1 332
box 8 5 126 98
use welltap_svt  __well_tap__3
timestamp 1730768468
transform 1 0 1712 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730768468
transform 1 0 1712 0 -1 296
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768468
transform 1 0 104 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768468
transform 1 0 104 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768468
transform 1 0 1712 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768468
transform 1 0 1712 0 1 356
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768468
transform 1 0 128 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768468
transform 1 0 104 0 -1 524
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768468
transform 1 0 128 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768468
transform 1 0 104 0 -1 524
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768468
transform 1 0 296 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768468
transform 1 0 296 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768468
transform 1 0 512 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768468
transform 1 0 512 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768468
transform 1 0 752 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768468
transform 1 0 752 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768468
transform 1 0 1008 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768468
transform 1 0 1008 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768468
transform 1 0 1272 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768468
transform 1 0 1272 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768468
transform 1 0 1536 0 -1 548
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768468
transform 1 0 1536 0 -1 548
box 8 5 126 98
use welltap_svt  __well_tap__7
timestamp 1730768468
transform 1 0 1712 0 -1 524
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730768468
transform 1 0 1712 0 -1 524
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768468
transform 1 0 104 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768468
transform 1 0 104 0 1 584
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768468
transform 1 0 216 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768468
transform 1 0 216 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768468
transform 1 0 408 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768468
transform 1 0 408 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768468
transform 1 0 616 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768468
transform 1 0 616 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768468
transform 1 0 848 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768468
transform 1 0 848 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768468
transform 1 0 1088 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768468
transform 1 0 1088 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768468
transform 1 0 1328 0 1 560
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768468
transform 1 0 1328 0 1 560
box 8 5 126 98
use welltap_svt  __well_tap__9
timestamp 1730768468
transform 1 0 1712 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730768468
transform 1 0 1712 0 1 584
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730768468
transform 1 0 104 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730768468
transform 1 0 104 0 -1 736
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768468
transform 1 0 672 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768468
transform 1 0 672 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768468
transform 1 0 832 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768468
transform 1 0 832 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768468
transform 1 0 1000 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768468
transform 1 0 1000 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768468
transform 1 0 1184 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768468
transform 1 0 1184 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768468
transform 1 0 1368 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768468
transform 1 0 1368 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768468
transform 1 0 1560 0 -1 760
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768468
transform 1 0 1560 0 -1 760
box 8 5 126 98
use welltap_svt  __well_tap__11
timestamp 1730768468
transform 1 0 1712 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730768468
transform 1 0 1712 0 -1 736
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768468
transform 1 0 104 0 1 800
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768468
transform 1 0 104 0 1 800
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768468
transform 1 0 736 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768468
transform 1 0 736 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768468
transform 1 0 872 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768468
transform 1 0 872 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768468
transform 1 0 1008 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768468
transform 1 0 1008 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768468
transform 1 0 1144 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768468
transform 1 0 1144 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768468
transform 1 0 1280 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768468
transform 1 0 1280 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768468
transform 1 0 1424 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768468
transform 1 0 1424 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768468
transform 1 0 1568 0 1 776
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768468
transform 1 0 1568 0 1 776
box 8 5 126 98
use welltap_svt  __well_tap__13
timestamp 1730768468
transform 1 0 1712 0 1 800
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730768468
transform 1 0 1712 0 1 800
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768468
transform 1 0 496 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768468
transform 1 0 496 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768468
transform 1 0 680 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768468
transform 1 0 680 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768468
transform 1 0 888 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768468
transform 1 0 888 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768468
transform 1 0 1104 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768468
transform 1 0 1104 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768468
transform 1 0 1336 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768468
transform 1 0 1336 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768468
transform 1 0 1568 0 -1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768468
transform 1 0 1568 0 -1 992
box 8 5 126 98
use welltap_svt  __well_tap__14
timestamp 1730768468
transform 1 0 104 0 -1 968
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730768468
transform 1 0 104 0 -1 968
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768468
transform 1 0 304 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768468
transform 1 0 304 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768468
transform 1 0 528 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768468
transform 1 0 528 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768468
transform 1 0 768 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768468
transform 1 0 768 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768468
transform 1 0 1016 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768468
transform 1 0 1016 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768468
transform 1 0 1272 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768468
transform 1 0 1272 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768468
transform 1 0 1536 0 1 992
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768468
transform 1 0 1536 0 1 992
box 8 5 126 98
use welltap_svt  __well_tap__15
timestamp 1730768468
transform 1 0 1712 0 -1 968
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730768468
transform 1 0 1712 0 -1 968
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730768468
transform 1 0 104 0 1 1016
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730768468
transform 1 0 104 0 1 1016
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730768468
transform 1 0 1712 0 1 1016
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730768468
transform 1 0 1712 0 1 1016
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768468
transform 1 0 128 0 -1 1212
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768468
transform 1 0 104 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768468
transform 1 0 128 0 -1 1212
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768468
transform 1 0 104 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768468
transform 1 0 296 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768468
transform 1 0 296 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768468
transform 1 0 512 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768468
transform 1 0 512 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768468
transform 1 0 744 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768468
transform 1 0 744 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768468
transform 1 0 992 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768468
transform 1 0 992 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768468
transform 1 0 1256 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768468
transform 1 0 1256 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768468
transform 1 0 1520 0 -1 1212
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768468
transform 1 0 1520 0 -1 1212
box 8 5 126 98
use welltap_svt  __well_tap__19
timestamp 1730768468
transform 1 0 1712 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730768468
transform 1 0 1712 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768468
transform 1 0 128 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768468
transform 1 0 104 0 1 1248
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768468
transform 1 0 128 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768468
transform 1 0 104 0 1 1248
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768468
transform 1 0 336 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768468
transform 1 0 336 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768468
transform 1 0 600 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768468
transform 1 0 600 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768468
transform 1 0 888 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768468
transform 1 0 888 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768468
transform 1 0 1200 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768468
transform 1 0 1200 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768468
transform 1 0 1512 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768468
transform 1 0 1512 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__21
timestamp 1730768468
transform 1 0 1712 0 1 1248
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730768468
transform 1 0 1712 0 1 1248
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768468
transform 1 0 592 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768468
transform 1 0 592 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768468
transform 1 0 728 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768468
transform 1 0 728 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768468
transform 1 0 864 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768468
transform 1 0 864 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768468
transform 1 0 1008 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768468
transform 1 0 1008 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768468
transform 1 0 1152 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768468
transform 1 0 1152 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768468
transform 1 0 1296 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768468
transform 1 0 1296 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768468
transform 1 0 1432 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768468
transform 1 0 1432 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768468
transform 1 0 1568 0 -1 1440
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768468
transform 1 0 1568 0 -1 1440
box 8 5 126 98
use welltap_svt  __well_tap__22
timestamp 1730768468
transform 1 0 104 0 -1 1416
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730768468
transform 1 0 104 0 -1 1416
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768468
transform 1 0 480 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768468
transform 1 0 480 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768468
transform 1 0 616 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768468
transform 1 0 616 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768468
transform 1 0 752 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768468
transform 1 0 752 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768468
transform 1 0 888 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768468
transform 1 0 888 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768468
transform 1 0 1024 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768468
transform 1 0 1024 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768468
transform 1 0 1160 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768468
transform 1 0 1160 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768468
transform 1 0 1296 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768468
transform 1 0 1296 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768468
transform 1 0 1432 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768468
transform 1 0 1432 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768468
transform 1 0 1568 0 1 1456
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768468
transform 1 0 1568 0 1 1456
box 8 5 126 98
use welltap_svt  __well_tap__23
timestamp 1730768468
transform 1 0 1712 0 -1 1416
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730768468
transform 1 0 1712 0 -1 1416
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768468
transform 1 0 104 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768468
transform 1 0 104 0 1 1480
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768468
transform 1 0 200 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768468
transform 1 0 200 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768468
transform 1 0 336 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768468
transform 1 0 336 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768468
transform 1 0 472 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768468
transform 1 0 472 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768468
transform 1 0 608 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768468
transform 1 0 608 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768468
transform 1 0 744 0 -1 1668
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768468
transform 1 0 744 0 -1 1668
box 8 5 126 98
use welltap_svt  __well_tap__25
timestamp 1730768468
transform 1 0 1712 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730768468
transform 1 0 1712 0 1 1480
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730768468
transform 1 0 104 0 -1 1644
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730768468
transform 1 0 104 0 -1 1644
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768468
transform 1 0 1712 0 -1 1644
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768468
transform 1 0 1712 0 -1 1644
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768468
transform 1 0 128 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768468
transform 1 0 104 0 1 1704
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768468
transform 1 0 128 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768468
transform 1 0 104 0 1 1704
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768468
transform 1 0 264 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768468
transform 1 0 264 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768468
transform 1 0 400 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768468
transform 1 0 400 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768468
transform 1 0 536 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768468
transform 1 0 536 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768468
transform 1 0 672 0 1 1680
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768468
transform 1 0 672 0 1 1680
box 8 5 126 98
use welltap_svt  __well_tap__29
timestamp 1730768468
transform 1 0 1712 0 1 1704
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730768468
transform 1 0 1712 0 1 1704
box 8 4 12 24
<< end >>
