magic
tech sky130l
timestamp 1731220536
<< m2 >>
rect 3398 4067 3404 4068
rect 3398 4063 3399 4067
rect 3403 4063 3404 4067
rect 3398 4062 3404 4063
rect 3502 4067 3508 4068
rect 3502 4063 3503 4067
rect 3507 4063 3508 4067
rect 3502 4062 3508 4063
rect 3606 4067 3612 4068
rect 3606 4063 3607 4067
rect 3611 4063 3612 4067
rect 3606 4062 3612 4063
rect 3710 4067 3716 4068
rect 3710 4063 3711 4067
rect 3715 4063 3716 4067
rect 3710 4062 3716 4063
rect 2070 4048 2076 4049
rect 2070 4044 2071 4048
rect 2075 4044 2076 4048
rect 2070 4043 2076 4044
rect 3990 4048 3996 4049
rect 3990 4044 3991 4048
rect 3995 4044 3996 4048
rect 3990 4043 3996 4044
rect 494 4031 500 4032
rect 494 4027 495 4031
rect 499 4027 500 4031
rect 494 4026 500 4027
rect 598 4031 604 4032
rect 598 4027 599 4031
rect 603 4027 604 4031
rect 598 4026 604 4027
rect 702 4031 708 4032
rect 702 4027 703 4031
rect 707 4027 708 4031
rect 702 4026 708 4027
rect 806 4031 812 4032
rect 806 4027 807 4031
rect 811 4027 812 4031
rect 806 4026 812 4027
rect 910 4031 916 4032
rect 910 4027 911 4031
rect 915 4027 916 4031
rect 910 4026 916 4027
rect 1014 4031 1020 4032
rect 1014 4027 1015 4031
rect 1019 4027 1020 4031
rect 1014 4026 1020 4027
rect 1118 4031 1124 4032
rect 1118 4027 1119 4031
rect 1123 4027 1124 4031
rect 1118 4026 1124 4027
rect 1222 4031 1228 4032
rect 1222 4027 1223 4031
rect 1227 4027 1228 4031
rect 1222 4026 1228 4027
rect 1326 4031 1332 4032
rect 1326 4027 1327 4031
rect 1331 4027 1332 4031
rect 1326 4026 1332 4027
rect 1430 4031 1436 4032
rect 1430 4027 1431 4031
rect 1435 4027 1436 4031
rect 1430 4026 1436 4027
rect 2070 4031 2076 4032
rect 2070 4027 2071 4031
rect 2075 4027 2076 4031
rect 3990 4031 3996 4032
rect 3990 4027 3991 4031
rect 3995 4027 3996 4031
rect 2070 4026 2076 4027
rect 3398 4026 3404 4027
rect 3398 4022 3399 4026
rect 3403 4022 3404 4026
rect 3398 4021 3404 4022
rect 3502 4026 3508 4027
rect 3502 4022 3503 4026
rect 3507 4022 3508 4026
rect 3502 4021 3508 4022
rect 3606 4026 3612 4027
rect 3606 4022 3607 4026
rect 3611 4022 3612 4026
rect 3606 4021 3612 4022
rect 3710 4026 3716 4027
rect 3990 4026 3996 4027
rect 3710 4022 3711 4026
rect 3715 4022 3716 4026
rect 3710 4021 3716 4022
rect 110 4012 116 4013
rect 110 4008 111 4012
rect 115 4008 116 4012
rect 110 4007 116 4008
rect 2030 4012 2036 4013
rect 2030 4008 2031 4012
rect 2035 4008 2036 4012
rect 2030 4007 2036 4008
rect 110 3995 116 3996
rect 110 3991 111 3995
rect 115 3991 116 3995
rect 2030 3995 2036 3996
rect 2030 3991 2031 3995
rect 2035 3991 2036 3995
rect 110 3990 116 3991
rect 494 3990 500 3991
rect 494 3986 495 3990
rect 499 3986 500 3990
rect 494 3985 500 3986
rect 598 3990 604 3991
rect 598 3986 599 3990
rect 603 3986 604 3990
rect 598 3985 604 3986
rect 702 3990 708 3991
rect 702 3986 703 3990
rect 707 3986 708 3990
rect 702 3985 708 3986
rect 806 3990 812 3991
rect 806 3986 807 3990
rect 811 3986 812 3990
rect 806 3985 812 3986
rect 910 3990 916 3991
rect 910 3986 911 3990
rect 915 3986 916 3990
rect 910 3985 916 3986
rect 1014 3990 1020 3991
rect 1014 3986 1015 3990
rect 1019 3986 1020 3990
rect 1014 3985 1020 3986
rect 1118 3990 1124 3991
rect 1118 3986 1119 3990
rect 1123 3986 1124 3990
rect 1118 3985 1124 3986
rect 1222 3990 1228 3991
rect 1222 3986 1223 3990
rect 1227 3986 1228 3990
rect 1222 3985 1228 3986
rect 1326 3990 1332 3991
rect 1326 3986 1327 3990
rect 1331 3986 1332 3990
rect 1326 3985 1332 3986
rect 1430 3990 1436 3991
rect 2030 3990 2036 3991
rect 2110 3994 2116 3995
rect 2110 3990 2111 3994
rect 2115 3990 2116 3994
rect 1430 3986 1431 3990
rect 1435 3986 1436 3990
rect 1430 3985 1436 3986
rect 2070 3989 2076 3990
rect 2110 3989 2116 3990
rect 2214 3994 2220 3995
rect 2214 3990 2215 3994
rect 2219 3990 2220 3994
rect 2214 3989 2220 3990
rect 2318 3994 2324 3995
rect 2318 3990 2319 3994
rect 2323 3990 2324 3994
rect 2318 3989 2324 3990
rect 2422 3994 2428 3995
rect 2422 3990 2423 3994
rect 2427 3990 2428 3994
rect 2422 3989 2428 3990
rect 2526 3994 2532 3995
rect 2526 3990 2527 3994
rect 2531 3990 2532 3994
rect 2526 3989 2532 3990
rect 2646 3994 2652 3995
rect 2646 3990 2647 3994
rect 2651 3990 2652 3994
rect 2646 3989 2652 3990
rect 2774 3994 2780 3995
rect 2774 3990 2775 3994
rect 2779 3990 2780 3994
rect 2774 3989 2780 3990
rect 2902 3994 2908 3995
rect 2902 3990 2903 3994
rect 2907 3990 2908 3994
rect 2902 3989 2908 3990
rect 3030 3994 3036 3995
rect 3030 3990 3031 3994
rect 3035 3990 3036 3994
rect 3030 3989 3036 3990
rect 3158 3994 3164 3995
rect 3158 3990 3159 3994
rect 3163 3990 3164 3994
rect 3158 3989 3164 3990
rect 3286 3994 3292 3995
rect 3286 3990 3287 3994
rect 3291 3990 3292 3994
rect 3286 3989 3292 3990
rect 3414 3994 3420 3995
rect 3414 3990 3415 3994
rect 3419 3990 3420 3994
rect 3414 3989 3420 3990
rect 3550 3994 3556 3995
rect 3550 3990 3551 3994
rect 3555 3990 3556 3994
rect 3550 3989 3556 3990
rect 3990 3989 3996 3990
rect 2070 3985 2071 3989
rect 2075 3985 2076 3989
rect 2070 3984 2076 3985
rect 3990 3985 3991 3989
rect 3995 3985 3996 3989
rect 3990 3984 3996 3985
rect 2070 3972 2076 3973
rect 2070 3968 2071 3972
rect 2075 3968 2076 3972
rect 2070 3967 2076 3968
rect 3990 3972 3996 3973
rect 3990 3968 3991 3972
rect 3995 3968 3996 3972
rect 3990 3967 3996 3968
rect 390 3958 396 3959
rect 390 3954 391 3958
rect 395 3954 396 3958
rect 110 3953 116 3954
rect 390 3953 396 3954
rect 494 3958 500 3959
rect 494 3954 495 3958
rect 499 3954 500 3958
rect 494 3953 500 3954
rect 598 3958 604 3959
rect 598 3954 599 3958
rect 603 3954 604 3958
rect 598 3953 604 3954
rect 702 3958 708 3959
rect 702 3954 703 3958
rect 707 3954 708 3958
rect 702 3953 708 3954
rect 806 3958 812 3959
rect 806 3954 807 3958
rect 811 3954 812 3958
rect 806 3953 812 3954
rect 910 3958 916 3959
rect 910 3954 911 3958
rect 915 3954 916 3958
rect 910 3953 916 3954
rect 1014 3958 1020 3959
rect 1014 3954 1015 3958
rect 1019 3954 1020 3958
rect 1014 3953 1020 3954
rect 1118 3958 1124 3959
rect 1118 3954 1119 3958
rect 1123 3954 1124 3958
rect 1118 3953 1124 3954
rect 1222 3958 1228 3959
rect 1222 3954 1223 3958
rect 1227 3954 1228 3958
rect 1222 3953 1228 3954
rect 1326 3958 1332 3959
rect 1326 3954 1327 3958
rect 1331 3954 1332 3958
rect 1326 3953 1332 3954
rect 1430 3958 1436 3959
rect 1430 3954 1431 3958
rect 1435 3954 1436 3958
rect 1430 3953 1436 3954
rect 1534 3958 1540 3959
rect 1534 3954 1535 3958
rect 1539 3954 1540 3958
rect 1534 3953 1540 3954
rect 2030 3953 2036 3954
rect 110 3949 111 3953
rect 115 3949 116 3953
rect 110 3948 116 3949
rect 2030 3949 2031 3953
rect 2035 3949 2036 3953
rect 2030 3948 2036 3949
rect 2110 3953 2116 3954
rect 2110 3949 2111 3953
rect 2115 3949 2116 3953
rect 2110 3948 2116 3949
rect 2214 3953 2220 3954
rect 2214 3949 2215 3953
rect 2219 3949 2220 3953
rect 2214 3948 2220 3949
rect 2318 3953 2324 3954
rect 2318 3949 2319 3953
rect 2323 3949 2324 3953
rect 2318 3948 2324 3949
rect 2422 3953 2428 3954
rect 2422 3949 2423 3953
rect 2427 3949 2428 3953
rect 2422 3948 2428 3949
rect 2526 3953 2532 3954
rect 2526 3949 2527 3953
rect 2531 3949 2532 3953
rect 2526 3948 2532 3949
rect 2646 3953 2652 3954
rect 2646 3949 2647 3953
rect 2651 3949 2652 3953
rect 2646 3948 2652 3949
rect 2774 3953 2780 3954
rect 2774 3949 2775 3953
rect 2779 3949 2780 3953
rect 2774 3948 2780 3949
rect 2902 3953 2908 3954
rect 2902 3949 2903 3953
rect 2907 3949 2908 3953
rect 2902 3948 2908 3949
rect 3030 3953 3036 3954
rect 3030 3949 3031 3953
rect 3035 3949 3036 3953
rect 3030 3948 3036 3949
rect 3158 3953 3164 3954
rect 3158 3949 3159 3953
rect 3163 3949 3164 3953
rect 3158 3948 3164 3949
rect 3286 3953 3292 3954
rect 3286 3949 3287 3953
rect 3291 3949 3292 3953
rect 3286 3948 3292 3949
rect 3414 3953 3420 3954
rect 3414 3949 3415 3953
rect 3419 3949 3420 3953
rect 3414 3948 3420 3949
rect 3550 3953 3556 3954
rect 3550 3949 3551 3953
rect 3555 3949 3556 3953
rect 3550 3948 3556 3949
rect 110 3936 116 3937
rect 110 3932 111 3936
rect 115 3932 116 3936
rect 110 3931 116 3932
rect 2030 3936 2036 3937
rect 2030 3932 2031 3936
rect 2035 3932 2036 3936
rect 2030 3931 2036 3932
rect 2142 3919 2148 3920
rect 390 3917 396 3918
rect 390 3913 391 3917
rect 395 3913 396 3917
rect 390 3912 396 3913
rect 494 3917 500 3918
rect 494 3913 495 3917
rect 499 3913 500 3917
rect 494 3912 500 3913
rect 598 3917 604 3918
rect 598 3913 599 3917
rect 603 3913 604 3917
rect 598 3912 604 3913
rect 702 3917 708 3918
rect 702 3913 703 3917
rect 707 3913 708 3917
rect 702 3912 708 3913
rect 806 3917 812 3918
rect 806 3913 807 3917
rect 811 3913 812 3917
rect 806 3912 812 3913
rect 910 3917 916 3918
rect 910 3913 911 3917
rect 915 3913 916 3917
rect 910 3912 916 3913
rect 1014 3917 1020 3918
rect 1014 3913 1015 3917
rect 1019 3913 1020 3917
rect 1014 3912 1020 3913
rect 1118 3917 1124 3918
rect 1118 3913 1119 3917
rect 1123 3913 1124 3917
rect 1118 3912 1124 3913
rect 1222 3917 1228 3918
rect 1222 3913 1223 3917
rect 1227 3913 1228 3917
rect 1222 3912 1228 3913
rect 1326 3917 1332 3918
rect 1326 3913 1327 3917
rect 1331 3913 1332 3917
rect 1326 3912 1332 3913
rect 1430 3917 1436 3918
rect 1430 3913 1431 3917
rect 1435 3913 1436 3917
rect 1430 3912 1436 3913
rect 1534 3917 1540 3918
rect 1534 3913 1535 3917
rect 1539 3913 1540 3917
rect 2142 3915 2143 3919
rect 2147 3915 2148 3919
rect 2142 3914 2148 3915
rect 2318 3919 2324 3920
rect 2318 3915 2319 3919
rect 2323 3915 2324 3919
rect 2318 3914 2324 3915
rect 2486 3919 2492 3920
rect 2486 3915 2487 3919
rect 2491 3915 2492 3919
rect 2486 3914 2492 3915
rect 2646 3919 2652 3920
rect 2646 3915 2647 3919
rect 2651 3915 2652 3919
rect 2646 3914 2652 3915
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2950 3919 2956 3920
rect 2950 3915 2951 3919
rect 2955 3915 2956 3919
rect 2950 3914 2956 3915
rect 3102 3919 3108 3920
rect 3102 3915 3103 3919
rect 3107 3915 3108 3919
rect 3102 3914 3108 3915
rect 3254 3919 3260 3920
rect 3254 3915 3255 3919
rect 3259 3915 3260 3919
rect 3254 3914 3260 3915
rect 1534 3912 1540 3913
rect 2070 3900 2076 3901
rect 2070 3896 2071 3900
rect 2075 3896 2076 3900
rect 2070 3895 2076 3896
rect 3990 3900 3996 3901
rect 3990 3896 3991 3900
rect 3995 3896 3996 3900
rect 3990 3895 3996 3896
rect 374 3883 380 3884
rect 374 3879 375 3883
rect 379 3879 380 3883
rect 374 3878 380 3879
rect 494 3883 500 3884
rect 494 3879 495 3883
rect 499 3879 500 3883
rect 494 3878 500 3879
rect 622 3883 628 3884
rect 622 3879 623 3883
rect 627 3879 628 3883
rect 622 3878 628 3879
rect 758 3883 764 3884
rect 758 3879 759 3883
rect 763 3879 764 3883
rect 758 3878 764 3879
rect 894 3883 900 3884
rect 894 3879 895 3883
rect 899 3879 900 3883
rect 894 3878 900 3879
rect 1022 3883 1028 3884
rect 1022 3879 1023 3883
rect 1027 3879 1028 3883
rect 1022 3878 1028 3879
rect 1150 3883 1156 3884
rect 1150 3879 1151 3883
rect 1155 3879 1156 3883
rect 1150 3878 1156 3879
rect 1278 3883 1284 3884
rect 1278 3879 1279 3883
rect 1283 3879 1284 3883
rect 1278 3878 1284 3879
rect 1414 3883 1420 3884
rect 1414 3879 1415 3883
rect 1419 3879 1420 3883
rect 1414 3878 1420 3879
rect 1550 3883 1556 3884
rect 1550 3879 1551 3883
rect 1555 3879 1556 3883
rect 1550 3878 1556 3879
rect 2070 3883 2076 3884
rect 2070 3879 2071 3883
rect 2075 3879 2076 3883
rect 3990 3883 3996 3884
rect 3990 3879 3991 3883
rect 3995 3879 3996 3883
rect 2070 3878 2076 3879
rect 2142 3878 2148 3879
rect 2142 3874 2143 3878
rect 2147 3874 2148 3878
rect 2142 3873 2148 3874
rect 2318 3878 2324 3879
rect 2318 3874 2319 3878
rect 2323 3874 2324 3878
rect 2318 3873 2324 3874
rect 2486 3878 2492 3879
rect 2486 3874 2487 3878
rect 2491 3874 2492 3878
rect 2486 3873 2492 3874
rect 2646 3878 2652 3879
rect 2646 3874 2647 3878
rect 2651 3874 2652 3878
rect 2646 3873 2652 3874
rect 2798 3878 2804 3879
rect 2798 3874 2799 3878
rect 2803 3874 2804 3878
rect 2798 3873 2804 3874
rect 2950 3878 2956 3879
rect 2950 3874 2951 3878
rect 2955 3874 2956 3878
rect 2950 3873 2956 3874
rect 3102 3878 3108 3879
rect 3102 3874 3103 3878
rect 3107 3874 3108 3878
rect 3102 3873 3108 3874
rect 3254 3878 3260 3879
rect 3990 3878 3996 3879
rect 3254 3874 3255 3878
rect 3259 3874 3260 3878
rect 3254 3873 3260 3874
rect 110 3864 116 3865
rect 110 3860 111 3864
rect 115 3860 116 3864
rect 110 3859 116 3860
rect 2030 3864 2036 3865
rect 2030 3860 2031 3864
rect 2035 3860 2036 3864
rect 2030 3859 2036 3860
rect 110 3847 116 3848
rect 110 3843 111 3847
rect 115 3843 116 3847
rect 2030 3847 2036 3848
rect 2030 3843 2031 3847
rect 2035 3843 2036 3847
rect 110 3842 116 3843
rect 374 3842 380 3843
rect 374 3838 375 3842
rect 379 3838 380 3842
rect 374 3837 380 3838
rect 494 3842 500 3843
rect 494 3838 495 3842
rect 499 3838 500 3842
rect 494 3837 500 3838
rect 622 3842 628 3843
rect 622 3838 623 3842
rect 627 3838 628 3842
rect 622 3837 628 3838
rect 758 3842 764 3843
rect 758 3838 759 3842
rect 763 3838 764 3842
rect 758 3837 764 3838
rect 894 3842 900 3843
rect 894 3838 895 3842
rect 899 3838 900 3842
rect 894 3837 900 3838
rect 1022 3842 1028 3843
rect 1022 3838 1023 3842
rect 1027 3838 1028 3842
rect 1022 3837 1028 3838
rect 1150 3842 1156 3843
rect 1150 3838 1151 3842
rect 1155 3838 1156 3842
rect 1150 3837 1156 3838
rect 1278 3842 1284 3843
rect 1278 3838 1279 3842
rect 1283 3838 1284 3842
rect 1278 3837 1284 3838
rect 1414 3842 1420 3843
rect 1414 3838 1415 3842
rect 1419 3838 1420 3842
rect 1414 3837 1420 3838
rect 1550 3842 1556 3843
rect 2030 3842 2036 3843
rect 2118 3846 2124 3847
rect 2118 3842 2119 3846
rect 2123 3842 2124 3846
rect 1550 3838 1551 3842
rect 1555 3838 1556 3842
rect 1550 3837 1556 3838
rect 2070 3841 2076 3842
rect 2118 3841 2124 3842
rect 2286 3846 2292 3847
rect 2286 3842 2287 3846
rect 2291 3842 2292 3846
rect 2286 3841 2292 3842
rect 2446 3846 2452 3847
rect 2446 3842 2447 3846
rect 2451 3842 2452 3846
rect 2446 3841 2452 3842
rect 2598 3846 2604 3847
rect 2598 3842 2599 3846
rect 2603 3842 2604 3846
rect 2598 3841 2604 3842
rect 2742 3846 2748 3847
rect 2742 3842 2743 3846
rect 2747 3842 2748 3846
rect 2742 3841 2748 3842
rect 2878 3846 2884 3847
rect 2878 3842 2879 3846
rect 2883 3842 2884 3846
rect 2878 3841 2884 3842
rect 3022 3846 3028 3847
rect 3022 3842 3023 3846
rect 3027 3842 3028 3846
rect 3022 3841 3028 3842
rect 3166 3846 3172 3847
rect 3166 3842 3167 3846
rect 3171 3842 3172 3846
rect 3166 3841 3172 3842
rect 3990 3841 3996 3842
rect 2070 3837 2071 3841
rect 2075 3837 2076 3841
rect 2070 3836 2076 3837
rect 3990 3837 3991 3841
rect 3995 3837 3996 3841
rect 3990 3836 3996 3837
rect 2070 3824 2076 3825
rect 2070 3820 2071 3824
rect 2075 3820 2076 3824
rect 2070 3819 2076 3820
rect 3990 3824 3996 3825
rect 3990 3820 3991 3824
rect 3995 3820 3996 3824
rect 3990 3819 3996 3820
rect 2118 3805 2124 3806
rect 430 3802 436 3803
rect 430 3798 431 3802
rect 435 3798 436 3802
rect 110 3797 116 3798
rect 430 3797 436 3798
rect 574 3802 580 3803
rect 574 3798 575 3802
rect 579 3798 580 3802
rect 574 3797 580 3798
rect 718 3802 724 3803
rect 718 3798 719 3802
rect 723 3798 724 3802
rect 718 3797 724 3798
rect 862 3802 868 3803
rect 862 3798 863 3802
rect 867 3798 868 3802
rect 862 3797 868 3798
rect 998 3802 1004 3803
rect 998 3798 999 3802
rect 1003 3798 1004 3802
rect 998 3797 1004 3798
rect 1134 3802 1140 3803
rect 1134 3798 1135 3802
rect 1139 3798 1140 3802
rect 1134 3797 1140 3798
rect 1270 3802 1276 3803
rect 1270 3798 1271 3802
rect 1275 3798 1276 3802
rect 1270 3797 1276 3798
rect 1406 3802 1412 3803
rect 1406 3798 1407 3802
rect 1411 3798 1412 3802
rect 1406 3797 1412 3798
rect 1550 3802 1556 3803
rect 1550 3798 1551 3802
rect 1555 3798 1556 3802
rect 2118 3801 2119 3805
rect 2123 3801 2124 3805
rect 2118 3800 2124 3801
rect 2286 3805 2292 3806
rect 2286 3801 2287 3805
rect 2291 3801 2292 3805
rect 2286 3800 2292 3801
rect 2446 3805 2452 3806
rect 2446 3801 2447 3805
rect 2451 3801 2452 3805
rect 2446 3800 2452 3801
rect 2598 3805 2604 3806
rect 2598 3801 2599 3805
rect 2603 3801 2604 3805
rect 2598 3800 2604 3801
rect 2742 3805 2748 3806
rect 2742 3801 2743 3805
rect 2747 3801 2748 3805
rect 2742 3800 2748 3801
rect 2878 3805 2884 3806
rect 2878 3801 2879 3805
rect 2883 3801 2884 3805
rect 2878 3800 2884 3801
rect 3022 3805 3028 3806
rect 3022 3801 3023 3805
rect 3027 3801 3028 3805
rect 3022 3800 3028 3801
rect 3166 3805 3172 3806
rect 3166 3801 3167 3805
rect 3171 3801 3172 3805
rect 3166 3800 3172 3801
rect 1550 3797 1556 3798
rect 2030 3797 2036 3798
rect 110 3793 111 3797
rect 115 3793 116 3797
rect 110 3792 116 3793
rect 2030 3793 2031 3797
rect 2035 3793 2036 3797
rect 2030 3792 2036 3793
rect 110 3780 116 3781
rect 110 3776 111 3780
rect 115 3776 116 3780
rect 110 3775 116 3776
rect 2030 3780 2036 3781
rect 2030 3776 2031 3780
rect 2035 3776 2036 3780
rect 2030 3775 2036 3776
rect 2110 3771 2116 3772
rect 2110 3767 2111 3771
rect 2115 3767 2116 3771
rect 2110 3766 2116 3767
rect 2238 3771 2244 3772
rect 2238 3767 2239 3771
rect 2243 3767 2244 3771
rect 2238 3766 2244 3767
rect 2390 3771 2396 3772
rect 2390 3767 2391 3771
rect 2395 3767 2396 3771
rect 2390 3766 2396 3767
rect 2542 3771 2548 3772
rect 2542 3767 2543 3771
rect 2547 3767 2548 3771
rect 2542 3766 2548 3767
rect 2686 3771 2692 3772
rect 2686 3767 2687 3771
rect 2691 3767 2692 3771
rect 2686 3766 2692 3767
rect 2822 3771 2828 3772
rect 2822 3767 2823 3771
rect 2827 3767 2828 3771
rect 2822 3766 2828 3767
rect 2950 3771 2956 3772
rect 2950 3767 2951 3771
rect 2955 3767 2956 3771
rect 2950 3766 2956 3767
rect 3086 3771 3092 3772
rect 3086 3767 3087 3771
rect 3091 3767 3092 3771
rect 3086 3766 3092 3767
rect 3222 3771 3228 3772
rect 3222 3767 3223 3771
rect 3227 3767 3228 3771
rect 3222 3766 3228 3767
rect 430 3761 436 3762
rect 430 3757 431 3761
rect 435 3757 436 3761
rect 430 3756 436 3757
rect 574 3761 580 3762
rect 574 3757 575 3761
rect 579 3757 580 3761
rect 574 3756 580 3757
rect 718 3761 724 3762
rect 718 3757 719 3761
rect 723 3757 724 3761
rect 718 3756 724 3757
rect 862 3761 868 3762
rect 862 3757 863 3761
rect 867 3757 868 3761
rect 862 3756 868 3757
rect 998 3761 1004 3762
rect 998 3757 999 3761
rect 1003 3757 1004 3761
rect 998 3756 1004 3757
rect 1134 3761 1140 3762
rect 1134 3757 1135 3761
rect 1139 3757 1140 3761
rect 1134 3756 1140 3757
rect 1270 3761 1276 3762
rect 1270 3757 1271 3761
rect 1275 3757 1276 3761
rect 1270 3756 1276 3757
rect 1406 3761 1412 3762
rect 1406 3757 1407 3761
rect 1411 3757 1412 3761
rect 1406 3756 1412 3757
rect 1550 3761 1556 3762
rect 1550 3757 1551 3761
rect 1555 3757 1556 3761
rect 1550 3756 1556 3757
rect 2070 3752 2076 3753
rect 2070 3748 2071 3752
rect 2075 3748 2076 3752
rect 2070 3747 2076 3748
rect 3990 3752 3996 3753
rect 3990 3748 3991 3752
rect 3995 3748 3996 3752
rect 3990 3747 3996 3748
rect 2070 3735 2076 3736
rect 2070 3731 2071 3735
rect 2075 3731 2076 3735
rect 3990 3735 3996 3736
rect 3990 3731 3991 3735
rect 3995 3731 3996 3735
rect 2070 3730 2076 3731
rect 2110 3730 2116 3731
rect 2110 3726 2111 3730
rect 2115 3726 2116 3730
rect 2110 3725 2116 3726
rect 2238 3730 2244 3731
rect 2238 3726 2239 3730
rect 2243 3726 2244 3730
rect 2238 3725 2244 3726
rect 2390 3730 2396 3731
rect 2390 3726 2391 3730
rect 2395 3726 2396 3730
rect 2390 3725 2396 3726
rect 2542 3730 2548 3731
rect 2542 3726 2543 3730
rect 2547 3726 2548 3730
rect 2542 3725 2548 3726
rect 2686 3730 2692 3731
rect 2686 3726 2687 3730
rect 2691 3726 2692 3730
rect 2686 3725 2692 3726
rect 2822 3730 2828 3731
rect 2822 3726 2823 3730
rect 2827 3726 2828 3730
rect 2822 3725 2828 3726
rect 2950 3730 2956 3731
rect 2950 3726 2951 3730
rect 2955 3726 2956 3730
rect 2950 3725 2956 3726
rect 3086 3730 3092 3731
rect 3086 3726 3087 3730
rect 3091 3726 3092 3730
rect 3086 3725 3092 3726
rect 3222 3730 3228 3731
rect 3990 3730 3996 3731
rect 3222 3726 3223 3730
rect 3227 3726 3228 3730
rect 3222 3725 3228 3726
rect 358 3723 364 3724
rect 358 3719 359 3723
rect 363 3719 364 3723
rect 358 3718 364 3719
rect 494 3723 500 3724
rect 494 3719 495 3723
rect 499 3719 500 3723
rect 494 3718 500 3719
rect 630 3723 636 3724
rect 630 3719 631 3723
rect 635 3719 636 3723
rect 630 3718 636 3719
rect 774 3723 780 3724
rect 774 3719 775 3723
rect 779 3719 780 3723
rect 774 3718 780 3719
rect 918 3723 924 3724
rect 918 3719 919 3723
rect 923 3719 924 3723
rect 918 3718 924 3719
rect 1070 3723 1076 3724
rect 1070 3719 1071 3723
rect 1075 3719 1076 3723
rect 1070 3718 1076 3719
rect 1222 3723 1228 3724
rect 1222 3719 1223 3723
rect 1227 3719 1228 3723
rect 1222 3718 1228 3719
rect 1374 3723 1380 3724
rect 1374 3719 1375 3723
rect 1379 3719 1380 3723
rect 1374 3718 1380 3719
rect 1526 3723 1532 3724
rect 1526 3719 1527 3723
rect 1531 3719 1532 3723
rect 1526 3718 1532 3719
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 110 3699 116 3700
rect 2030 3704 2036 3705
rect 2030 3700 2031 3704
rect 2035 3700 2036 3704
rect 2030 3699 2036 3700
rect 2110 3690 2116 3691
rect 110 3687 116 3688
rect 110 3683 111 3687
rect 115 3683 116 3687
rect 2030 3687 2036 3688
rect 2030 3683 2031 3687
rect 2035 3683 2036 3687
rect 2110 3686 2111 3690
rect 2115 3686 2116 3690
rect 110 3682 116 3683
rect 358 3682 364 3683
rect 358 3678 359 3682
rect 363 3678 364 3682
rect 358 3677 364 3678
rect 494 3682 500 3683
rect 494 3678 495 3682
rect 499 3678 500 3682
rect 494 3677 500 3678
rect 630 3682 636 3683
rect 630 3678 631 3682
rect 635 3678 636 3682
rect 630 3677 636 3678
rect 774 3682 780 3683
rect 774 3678 775 3682
rect 779 3678 780 3682
rect 774 3677 780 3678
rect 918 3682 924 3683
rect 918 3678 919 3682
rect 923 3678 924 3682
rect 918 3677 924 3678
rect 1070 3682 1076 3683
rect 1070 3678 1071 3682
rect 1075 3678 1076 3682
rect 1070 3677 1076 3678
rect 1222 3682 1228 3683
rect 1222 3678 1223 3682
rect 1227 3678 1228 3682
rect 1222 3677 1228 3678
rect 1374 3682 1380 3683
rect 1374 3678 1375 3682
rect 1379 3678 1380 3682
rect 1374 3677 1380 3678
rect 1526 3682 1532 3683
rect 2030 3682 2036 3683
rect 2070 3685 2076 3686
rect 2110 3685 2116 3686
rect 2294 3690 2300 3691
rect 2294 3686 2295 3690
rect 2299 3686 2300 3690
rect 2294 3685 2300 3686
rect 2486 3690 2492 3691
rect 2486 3686 2487 3690
rect 2491 3686 2492 3690
rect 2486 3685 2492 3686
rect 2670 3690 2676 3691
rect 2670 3686 2671 3690
rect 2675 3686 2676 3690
rect 2670 3685 2676 3686
rect 2846 3690 2852 3691
rect 2846 3686 2847 3690
rect 2851 3686 2852 3690
rect 2846 3685 2852 3686
rect 3014 3690 3020 3691
rect 3014 3686 3015 3690
rect 3019 3686 3020 3690
rect 3014 3685 3020 3686
rect 3182 3690 3188 3691
rect 3182 3686 3183 3690
rect 3187 3686 3188 3690
rect 3182 3685 3188 3686
rect 3358 3690 3364 3691
rect 3358 3686 3359 3690
rect 3363 3686 3364 3690
rect 3358 3685 3364 3686
rect 3990 3685 3996 3686
rect 1526 3678 1527 3682
rect 1531 3678 1532 3682
rect 2070 3681 2071 3685
rect 2075 3681 2076 3685
rect 2070 3680 2076 3681
rect 3990 3681 3991 3685
rect 3995 3681 3996 3685
rect 3990 3680 3996 3681
rect 1526 3677 1532 3678
rect 2070 3668 2076 3669
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 3990 3668 3996 3669
rect 3990 3664 3991 3668
rect 3995 3664 3996 3668
rect 3990 3663 3996 3664
rect 342 3650 348 3651
rect 342 3646 343 3650
rect 347 3646 348 3650
rect 110 3645 116 3646
rect 342 3645 348 3646
rect 518 3650 524 3651
rect 518 3646 519 3650
rect 523 3646 524 3650
rect 518 3645 524 3646
rect 694 3650 700 3651
rect 694 3646 695 3650
rect 699 3646 700 3650
rect 694 3645 700 3646
rect 862 3650 868 3651
rect 862 3646 863 3650
rect 867 3646 868 3650
rect 862 3645 868 3646
rect 1030 3650 1036 3651
rect 1030 3646 1031 3650
rect 1035 3646 1036 3650
rect 1030 3645 1036 3646
rect 1190 3650 1196 3651
rect 1190 3646 1191 3650
rect 1195 3646 1196 3650
rect 1190 3645 1196 3646
rect 1342 3650 1348 3651
rect 1342 3646 1343 3650
rect 1347 3646 1348 3650
rect 1342 3645 1348 3646
rect 1494 3650 1500 3651
rect 1494 3646 1495 3650
rect 1499 3646 1500 3650
rect 1494 3645 1500 3646
rect 1654 3650 1660 3651
rect 1654 3646 1655 3650
rect 1659 3646 1660 3650
rect 2110 3649 2116 3650
rect 1654 3645 1660 3646
rect 2030 3645 2036 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 110 3640 116 3641
rect 2030 3641 2031 3645
rect 2035 3641 2036 3645
rect 2110 3645 2111 3649
rect 2115 3645 2116 3649
rect 2110 3644 2116 3645
rect 2294 3649 2300 3650
rect 2294 3645 2295 3649
rect 2299 3645 2300 3649
rect 2294 3644 2300 3645
rect 2486 3649 2492 3650
rect 2486 3645 2487 3649
rect 2491 3645 2492 3649
rect 2486 3644 2492 3645
rect 2670 3649 2676 3650
rect 2670 3645 2671 3649
rect 2675 3645 2676 3649
rect 2670 3644 2676 3645
rect 2846 3649 2852 3650
rect 2846 3645 2847 3649
rect 2851 3645 2852 3649
rect 2846 3644 2852 3645
rect 3014 3649 3020 3650
rect 3014 3645 3015 3649
rect 3019 3645 3020 3649
rect 3014 3644 3020 3645
rect 3182 3649 3188 3650
rect 3182 3645 3183 3649
rect 3187 3645 3188 3649
rect 3182 3644 3188 3645
rect 3358 3649 3364 3650
rect 3358 3645 3359 3649
rect 3363 3645 3364 3649
rect 3358 3644 3364 3645
rect 2030 3640 2036 3641
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 2030 3628 2036 3629
rect 2030 3624 2031 3628
rect 2035 3624 2036 3628
rect 2030 3623 2036 3624
rect 2110 3611 2116 3612
rect 342 3609 348 3610
rect 342 3605 343 3609
rect 347 3605 348 3609
rect 342 3604 348 3605
rect 518 3609 524 3610
rect 518 3605 519 3609
rect 523 3605 524 3609
rect 518 3604 524 3605
rect 694 3609 700 3610
rect 694 3605 695 3609
rect 699 3605 700 3609
rect 694 3604 700 3605
rect 862 3609 868 3610
rect 862 3605 863 3609
rect 867 3605 868 3609
rect 862 3604 868 3605
rect 1030 3609 1036 3610
rect 1030 3605 1031 3609
rect 1035 3605 1036 3609
rect 1030 3604 1036 3605
rect 1190 3609 1196 3610
rect 1190 3605 1191 3609
rect 1195 3605 1196 3609
rect 1190 3604 1196 3605
rect 1342 3609 1348 3610
rect 1342 3605 1343 3609
rect 1347 3605 1348 3609
rect 1342 3604 1348 3605
rect 1494 3609 1500 3610
rect 1494 3605 1495 3609
rect 1499 3605 1500 3609
rect 1494 3604 1500 3605
rect 1654 3609 1660 3610
rect 1654 3605 1655 3609
rect 1659 3605 1660 3609
rect 2110 3607 2111 3611
rect 2115 3607 2116 3611
rect 2110 3606 2116 3607
rect 2294 3611 2300 3612
rect 2294 3607 2295 3611
rect 2299 3607 2300 3611
rect 2294 3606 2300 3607
rect 2494 3611 2500 3612
rect 2494 3607 2495 3611
rect 2499 3607 2500 3611
rect 2494 3606 2500 3607
rect 2686 3611 2692 3612
rect 2686 3607 2687 3611
rect 2691 3607 2692 3611
rect 2686 3606 2692 3607
rect 2862 3611 2868 3612
rect 2862 3607 2863 3611
rect 2867 3607 2868 3611
rect 2862 3606 2868 3607
rect 3022 3611 3028 3612
rect 3022 3607 3023 3611
rect 3027 3607 3028 3611
rect 3022 3606 3028 3607
rect 3166 3611 3172 3612
rect 3166 3607 3167 3611
rect 3171 3607 3172 3611
rect 3166 3606 3172 3607
rect 3302 3611 3308 3612
rect 3302 3607 3303 3611
rect 3307 3607 3308 3611
rect 3302 3606 3308 3607
rect 3430 3611 3436 3612
rect 3430 3607 3431 3611
rect 3435 3607 3436 3611
rect 3430 3606 3436 3607
rect 3550 3611 3556 3612
rect 3550 3607 3551 3611
rect 3555 3607 3556 3611
rect 3550 3606 3556 3607
rect 3670 3611 3676 3612
rect 3670 3607 3671 3611
rect 3675 3607 3676 3611
rect 3670 3606 3676 3607
rect 3790 3611 3796 3612
rect 3790 3607 3791 3611
rect 3795 3607 3796 3611
rect 3790 3606 3796 3607
rect 3894 3611 3900 3612
rect 3894 3607 3895 3611
rect 3899 3607 3900 3611
rect 3894 3606 3900 3607
rect 1654 3604 1660 3605
rect 2070 3592 2076 3593
rect 2070 3588 2071 3592
rect 2075 3588 2076 3592
rect 2070 3587 2076 3588
rect 3990 3592 3996 3593
rect 3990 3588 3991 3592
rect 3995 3588 3996 3592
rect 3990 3587 3996 3588
rect 238 3579 244 3580
rect 238 3575 239 3579
rect 243 3575 244 3579
rect 238 3574 244 3575
rect 398 3579 404 3580
rect 398 3575 399 3579
rect 403 3575 404 3579
rect 398 3574 404 3575
rect 550 3579 556 3580
rect 550 3575 551 3579
rect 555 3575 556 3579
rect 550 3574 556 3575
rect 702 3579 708 3580
rect 702 3575 703 3579
rect 707 3575 708 3579
rect 702 3574 708 3575
rect 854 3579 860 3580
rect 854 3575 855 3579
rect 859 3575 860 3579
rect 854 3574 860 3575
rect 998 3579 1004 3580
rect 998 3575 999 3579
rect 1003 3575 1004 3579
rect 998 3574 1004 3575
rect 1134 3579 1140 3580
rect 1134 3575 1135 3579
rect 1139 3575 1140 3579
rect 1134 3574 1140 3575
rect 1262 3579 1268 3580
rect 1262 3575 1263 3579
rect 1267 3575 1268 3579
rect 1262 3574 1268 3575
rect 1382 3579 1388 3580
rect 1382 3575 1383 3579
rect 1387 3575 1388 3579
rect 1382 3574 1388 3575
rect 1494 3579 1500 3580
rect 1494 3575 1495 3579
rect 1499 3575 1500 3579
rect 1494 3574 1500 3575
rect 1606 3579 1612 3580
rect 1606 3575 1607 3579
rect 1611 3575 1612 3579
rect 1606 3574 1612 3575
rect 1718 3579 1724 3580
rect 1718 3575 1719 3579
rect 1723 3575 1724 3579
rect 1718 3574 1724 3575
rect 1830 3579 1836 3580
rect 1830 3575 1831 3579
rect 1835 3575 1836 3579
rect 1830 3574 1836 3575
rect 1934 3579 1940 3580
rect 1934 3575 1935 3579
rect 1939 3575 1940 3579
rect 1934 3574 1940 3575
rect 2070 3575 2076 3576
rect 2070 3571 2071 3575
rect 2075 3571 2076 3575
rect 3990 3575 3996 3576
rect 3990 3571 3991 3575
rect 3995 3571 3996 3575
rect 2070 3570 2076 3571
rect 2110 3570 2116 3571
rect 2110 3566 2111 3570
rect 2115 3566 2116 3570
rect 2110 3565 2116 3566
rect 2294 3570 2300 3571
rect 2294 3566 2295 3570
rect 2299 3566 2300 3570
rect 2294 3565 2300 3566
rect 2494 3570 2500 3571
rect 2494 3566 2495 3570
rect 2499 3566 2500 3570
rect 2494 3565 2500 3566
rect 2686 3570 2692 3571
rect 2686 3566 2687 3570
rect 2691 3566 2692 3570
rect 2686 3565 2692 3566
rect 2862 3570 2868 3571
rect 2862 3566 2863 3570
rect 2867 3566 2868 3570
rect 2862 3565 2868 3566
rect 3022 3570 3028 3571
rect 3022 3566 3023 3570
rect 3027 3566 3028 3570
rect 3022 3565 3028 3566
rect 3166 3570 3172 3571
rect 3166 3566 3167 3570
rect 3171 3566 3172 3570
rect 3166 3565 3172 3566
rect 3302 3570 3308 3571
rect 3302 3566 3303 3570
rect 3307 3566 3308 3570
rect 3302 3565 3308 3566
rect 3430 3570 3436 3571
rect 3430 3566 3431 3570
rect 3435 3566 3436 3570
rect 3430 3565 3436 3566
rect 3550 3570 3556 3571
rect 3550 3566 3551 3570
rect 3555 3566 3556 3570
rect 3550 3565 3556 3566
rect 3670 3570 3676 3571
rect 3670 3566 3671 3570
rect 3675 3566 3676 3570
rect 3670 3565 3676 3566
rect 3790 3570 3796 3571
rect 3790 3566 3791 3570
rect 3795 3566 3796 3570
rect 3790 3565 3796 3566
rect 3894 3570 3900 3571
rect 3990 3570 3996 3571
rect 3894 3566 3895 3570
rect 3899 3566 3900 3570
rect 3894 3565 3900 3566
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 2030 3560 2036 3561
rect 2030 3556 2031 3560
rect 2035 3556 2036 3560
rect 2030 3555 2036 3556
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 2030 3543 2036 3544
rect 2030 3539 2031 3543
rect 2035 3539 2036 3543
rect 110 3538 116 3539
rect 238 3538 244 3539
rect 238 3534 239 3538
rect 243 3534 244 3538
rect 238 3533 244 3534
rect 398 3538 404 3539
rect 398 3534 399 3538
rect 403 3534 404 3538
rect 398 3533 404 3534
rect 550 3538 556 3539
rect 550 3534 551 3538
rect 555 3534 556 3538
rect 550 3533 556 3534
rect 702 3538 708 3539
rect 702 3534 703 3538
rect 707 3534 708 3538
rect 702 3533 708 3534
rect 854 3538 860 3539
rect 854 3534 855 3538
rect 859 3534 860 3538
rect 854 3533 860 3534
rect 998 3538 1004 3539
rect 998 3534 999 3538
rect 1003 3534 1004 3538
rect 998 3533 1004 3534
rect 1134 3538 1140 3539
rect 1134 3534 1135 3538
rect 1139 3534 1140 3538
rect 1134 3533 1140 3534
rect 1262 3538 1268 3539
rect 1262 3534 1263 3538
rect 1267 3534 1268 3538
rect 1262 3533 1268 3534
rect 1382 3538 1388 3539
rect 1382 3534 1383 3538
rect 1387 3534 1388 3538
rect 1382 3533 1388 3534
rect 1494 3538 1500 3539
rect 1494 3534 1495 3538
rect 1499 3534 1500 3538
rect 1494 3533 1500 3534
rect 1606 3538 1612 3539
rect 1606 3534 1607 3538
rect 1611 3534 1612 3538
rect 1606 3533 1612 3534
rect 1718 3538 1724 3539
rect 1718 3534 1719 3538
rect 1723 3534 1724 3538
rect 1718 3533 1724 3534
rect 1830 3538 1836 3539
rect 1830 3534 1831 3538
rect 1835 3534 1836 3538
rect 1830 3533 1836 3534
rect 1934 3538 1940 3539
rect 2030 3538 2036 3539
rect 1934 3534 1935 3538
rect 1939 3534 1940 3538
rect 1934 3533 1940 3534
rect 2446 3526 2452 3527
rect 2446 3522 2447 3526
rect 2451 3522 2452 3526
rect 2070 3521 2076 3522
rect 2446 3521 2452 3522
rect 2590 3526 2596 3527
rect 2590 3522 2591 3526
rect 2595 3522 2596 3526
rect 2590 3521 2596 3522
rect 2726 3526 2732 3527
rect 2726 3522 2727 3526
rect 2731 3522 2732 3526
rect 2726 3521 2732 3522
rect 2862 3526 2868 3527
rect 2862 3522 2863 3526
rect 2867 3522 2868 3526
rect 2862 3521 2868 3522
rect 2990 3526 2996 3527
rect 2990 3522 2991 3526
rect 2995 3522 2996 3526
rect 2990 3521 2996 3522
rect 3118 3526 3124 3527
rect 3118 3522 3119 3526
rect 3123 3522 3124 3526
rect 3118 3521 3124 3522
rect 3238 3526 3244 3527
rect 3238 3522 3239 3526
rect 3243 3522 3244 3526
rect 3238 3521 3244 3522
rect 3350 3526 3356 3527
rect 3350 3522 3351 3526
rect 3355 3522 3356 3526
rect 3350 3521 3356 3522
rect 3462 3526 3468 3527
rect 3462 3522 3463 3526
rect 3467 3522 3468 3526
rect 3462 3521 3468 3522
rect 3574 3526 3580 3527
rect 3574 3522 3575 3526
rect 3579 3522 3580 3526
rect 3574 3521 3580 3522
rect 3686 3526 3692 3527
rect 3686 3522 3687 3526
rect 3691 3522 3692 3526
rect 3686 3521 3692 3522
rect 3790 3526 3796 3527
rect 3790 3522 3791 3526
rect 3795 3522 3796 3526
rect 3790 3521 3796 3522
rect 3894 3526 3900 3527
rect 3894 3522 3895 3526
rect 3899 3522 3900 3526
rect 3894 3521 3900 3522
rect 3990 3521 3996 3522
rect 2070 3517 2071 3521
rect 2075 3517 2076 3521
rect 2070 3516 2076 3517
rect 3990 3517 3991 3521
rect 3995 3517 3996 3521
rect 3990 3516 3996 3517
rect 150 3506 156 3507
rect 150 3502 151 3506
rect 155 3502 156 3506
rect 110 3501 116 3502
rect 150 3501 156 3502
rect 374 3506 380 3507
rect 374 3502 375 3506
rect 379 3502 380 3506
rect 374 3501 380 3502
rect 614 3506 620 3507
rect 614 3502 615 3506
rect 619 3502 620 3506
rect 614 3501 620 3502
rect 846 3506 852 3507
rect 846 3502 847 3506
rect 851 3502 852 3506
rect 846 3501 852 3502
rect 1062 3506 1068 3507
rect 1062 3502 1063 3506
rect 1067 3502 1068 3506
rect 1062 3501 1068 3502
rect 1254 3506 1260 3507
rect 1254 3502 1255 3506
rect 1259 3502 1260 3506
rect 1254 3501 1260 3502
rect 1438 3506 1444 3507
rect 1438 3502 1439 3506
rect 1443 3502 1444 3506
rect 1438 3501 1444 3502
rect 1614 3506 1620 3507
rect 1614 3502 1615 3506
rect 1619 3502 1620 3506
rect 1614 3501 1620 3502
rect 1782 3506 1788 3507
rect 1782 3502 1783 3506
rect 1787 3502 1788 3506
rect 1782 3501 1788 3502
rect 1934 3506 1940 3507
rect 1934 3502 1935 3506
rect 1939 3502 1940 3506
rect 2070 3504 2076 3505
rect 1934 3501 1940 3502
rect 2030 3501 2036 3502
rect 110 3497 111 3501
rect 115 3497 116 3501
rect 110 3496 116 3497
rect 2030 3497 2031 3501
rect 2035 3497 2036 3501
rect 2070 3500 2071 3504
rect 2075 3500 2076 3504
rect 2070 3499 2076 3500
rect 3990 3504 3996 3505
rect 3990 3500 3991 3504
rect 3995 3500 3996 3504
rect 3990 3499 3996 3500
rect 2030 3496 2036 3497
rect 2446 3485 2452 3486
rect 110 3484 116 3485
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 2030 3484 2036 3485
rect 2030 3480 2031 3484
rect 2035 3480 2036 3484
rect 2446 3481 2447 3485
rect 2451 3481 2452 3485
rect 2446 3480 2452 3481
rect 2590 3485 2596 3486
rect 2590 3481 2591 3485
rect 2595 3481 2596 3485
rect 2590 3480 2596 3481
rect 2726 3485 2732 3486
rect 2726 3481 2727 3485
rect 2731 3481 2732 3485
rect 2726 3480 2732 3481
rect 2862 3485 2868 3486
rect 2862 3481 2863 3485
rect 2867 3481 2868 3485
rect 2862 3480 2868 3481
rect 2990 3485 2996 3486
rect 2990 3481 2991 3485
rect 2995 3481 2996 3485
rect 2990 3480 2996 3481
rect 3118 3485 3124 3486
rect 3118 3481 3119 3485
rect 3123 3481 3124 3485
rect 3118 3480 3124 3481
rect 3238 3485 3244 3486
rect 3238 3481 3239 3485
rect 3243 3481 3244 3485
rect 3238 3480 3244 3481
rect 3350 3485 3356 3486
rect 3350 3481 3351 3485
rect 3355 3481 3356 3485
rect 3350 3480 3356 3481
rect 3462 3485 3468 3486
rect 3462 3481 3463 3485
rect 3467 3481 3468 3485
rect 3462 3480 3468 3481
rect 3574 3485 3580 3486
rect 3574 3481 3575 3485
rect 3579 3481 3580 3485
rect 3574 3480 3580 3481
rect 3686 3485 3692 3486
rect 3686 3481 3687 3485
rect 3691 3481 3692 3485
rect 3686 3480 3692 3481
rect 3790 3485 3796 3486
rect 3790 3481 3791 3485
rect 3795 3481 3796 3485
rect 3790 3480 3796 3481
rect 3894 3485 3900 3486
rect 3894 3481 3895 3485
rect 3899 3481 3900 3485
rect 3894 3480 3900 3481
rect 2030 3479 2036 3480
rect 150 3465 156 3466
rect 150 3461 151 3465
rect 155 3461 156 3465
rect 150 3460 156 3461
rect 374 3465 380 3466
rect 374 3461 375 3465
rect 379 3461 380 3465
rect 374 3460 380 3461
rect 614 3465 620 3466
rect 614 3461 615 3465
rect 619 3461 620 3465
rect 614 3460 620 3461
rect 846 3465 852 3466
rect 846 3461 847 3465
rect 851 3461 852 3465
rect 846 3460 852 3461
rect 1062 3465 1068 3466
rect 1062 3461 1063 3465
rect 1067 3461 1068 3465
rect 1062 3460 1068 3461
rect 1254 3465 1260 3466
rect 1254 3461 1255 3465
rect 1259 3461 1260 3465
rect 1254 3460 1260 3461
rect 1438 3465 1444 3466
rect 1438 3461 1439 3465
rect 1443 3461 1444 3465
rect 1438 3460 1444 3461
rect 1614 3465 1620 3466
rect 1614 3461 1615 3465
rect 1619 3461 1620 3465
rect 1614 3460 1620 3461
rect 1782 3465 1788 3466
rect 1782 3461 1783 3465
rect 1787 3461 1788 3465
rect 1782 3460 1788 3461
rect 1934 3465 1940 3466
rect 1934 3461 1935 3465
rect 1939 3461 1940 3465
rect 1934 3460 1940 3461
rect 2342 3455 2348 3456
rect 2342 3451 2343 3455
rect 2347 3451 2348 3455
rect 2342 3450 2348 3451
rect 2854 3455 2860 3456
rect 2854 3451 2855 3455
rect 2859 3451 2860 3455
rect 2854 3450 2860 3451
rect 3374 3455 3380 3456
rect 3374 3451 3375 3455
rect 3379 3451 3380 3455
rect 3374 3450 3380 3451
rect 3894 3455 3900 3456
rect 3894 3451 3895 3455
rect 3899 3451 3900 3455
rect 3894 3450 3900 3451
rect 2070 3436 2076 3437
rect 2070 3432 2071 3436
rect 2075 3432 2076 3436
rect 2070 3431 2076 3432
rect 3990 3436 3996 3437
rect 3990 3432 3991 3436
rect 3995 3432 3996 3436
rect 3990 3431 3996 3432
rect 2070 3419 2076 3420
rect 2070 3415 2071 3419
rect 2075 3415 2076 3419
rect 3990 3419 3996 3420
rect 3990 3415 3991 3419
rect 3995 3415 3996 3419
rect 2070 3414 2076 3415
rect 2342 3414 2348 3415
rect 150 3411 156 3412
rect 150 3407 151 3411
rect 155 3407 156 3411
rect 150 3406 156 3407
rect 334 3411 340 3412
rect 334 3407 335 3411
rect 339 3407 340 3411
rect 334 3406 340 3407
rect 582 3411 588 3412
rect 582 3407 583 3411
rect 587 3407 588 3411
rect 582 3406 588 3407
rect 862 3411 868 3412
rect 862 3407 863 3411
rect 867 3407 868 3411
rect 862 3406 868 3407
rect 1158 3411 1164 3412
rect 1158 3407 1159 3411
rect 1163 3407 1164 3411
rect 1158 3406 1164 3407
rect 1462 3411 1468 3412
rect 1462 3407 1463 3411
rect 1467 3407 1468 3411
rect 2342 3410 2343 3414
rect 2347 3410 2348 3414
rect 2342 3409 2348 3410
rect 2854 3414 2860 3415
rect 2854 3410 2855 3414
rect 2859 3410 2860 3414
rect 2854 3409 2860 3410
rect 3374 3414 3380 3415
rect 3374 3410 3375 3414
rect 3379 3410 3380 3414
rect 3374 3409 3380 3410
rect 3894 3414 3900 3415
rect 3990 3414 3996 3415
rect 3894 3410 3895 3414
rect 3899 3410 3900 3414
rect 3894 3409 3900 3410
rect 1462 3406 1468 3407
rect 110 3392 116 3393
rect 110 3388 111 3392
rect 115 3388 116 3392
rect 110 3387 116 3388
rect 2030 3392 2036 3393
rect 2030 3388 2031 3392
rect 2035 3388 2036 3392
rect 2030 3387 2036 3388
rect 2182 3378 2188 3379
rect 110 3375 116 3376
rect 110 3371 111 3375
rect 115 3371 116 3375
rect 2030 3375 2036 3376
rect 2030 3371 2031 3375
rect 2035 3371 2036 3375
rect 2182 3374 2183 3378
rect 2187 3374 2188 3378
rect 110 3370 116 3371
rect 150 3370 156 3371
rect 150 3366 151 3370
rect 155 3366 156 3370
rect 150 3365 156 3366
rect 334 3370 340 3371
rect 334 3366 335 3370
rect 339 3366 340 3370
rect 334 3365 340 3366
rect 582 3370 588 3371
rect 582 3366 583 3370
rect 587 3366 588 3370
rect 582 3365 588 3366
rect 862 3370 868 3371
rect 862 3366 863 3370
rect 867 3366 868 3370
rect 862 3365 868 3366
rect 1158 3370 1164 3371
rect 1158 3366 1159 3370
rect 1163 3366 1164 3370
rect 1158 3365 1164 3366
rect 1462 3370 1468 3371
rect 2030 3370 2036 3371
rect 2070 3373 2076 3374
rect 2182 3373 2188 3374
rect 2582 3378 2588 3379
rect 2582 3374 2583 3378
rect 2587 3374 2588 3378
rect 2582 3373 2588 3374
rect 3006 3378 3012 3379
rect 3006 3374 3007 3378
rect 3011 3374 3012 3378
rect 3006 3373 3012 3374
rect 3446 3378 3452 3379
rect 3446 3374 3447 3378
rect 3451 3374 3452 3378
rect 3446 3373 3452 3374
rect 3894 3378 3900 3379
rect 3894 3374 3895 3378
rect 3899 3374 3900 3378
rect 3894 3373 3900 3374
rect 3990 3373 3996 3374
rect 1462 3366 1463 3370
rect 1467 3366 1468 3370
rect 2070 3369 2071 3373
rect 2075 3369 2076 3373
rect 2070 3368 2076 3369
rect 3990 3369 3991 3373
rect 3995 3369 3996 3373
rect 3990 3368 3996 3369
rect 1462 3365 1468 3366
rect 2070 3356 2076 3357
rect 2070 3352 2071 3356
rect 2075 3352 2076 3356
rect 2070 3351 2076 3352
rect 3990 3356 3996 3357
rect 3990 3352 3991 3356
rect 3995 3352 3996 3356
rect 3990 3351 3996 3352
rect 2182 3337 2188 3338
rect 2182 3333 2183 3337
rect 2187 3333 2188 3337
rect 2182 3332 2188 3333
rect 2582 3337 2588 3338
rect 2582 3333 2583 3337
rect 2587 3333 2588 3337
rect 2582 3332 2588 3333
rect 3006 3337 3012 3338
rect 3006 3333 3007 3337
rect 3011 3333 3012 3337
rect 3006 3332 3012 3333
rect 3446 3337 3452 3338
rect 3446 3333 3447 3337
rect 3451 3333 3452 3337
rect 3446 3332 3452 3333
rect 3894 3337 3900 3338
rect 3894 3333 3895 3337
rect 3899 3333 3900 3337
rect 3894 3332 3900 3333
rect 150 3330 156 3331
rect 150 3326 151 3330
rect 155 3326 156 3330
rect 110 3325 116 3326
rect 150 3325 156 3326
rect 286 3330 292 3331
rect 286 3326 287 3330
rect 291 3326 292 3330
rect 286 3325 292 3326
rect 462 3330 468 3331
rect 462 3326 463 3330
rect 467 3326 468 3330
rect 462 3325 468 3326
rect 638 3330 644 3331
rect 638 3326 639 3330
rect 643 3326 644 3330
rect 638 3325 644 3326
rect 814 3330 820 3331
rect 814 3326 815 3330
rect 819 3326 820 3330
rect 814 3325 820 3326
rect 990 3330 996 3331
rect 990 3326 991 3330
rect 995 3326 996 3330
rect 990 3325 996 3326
rect 1158 3330 1164 3331
rect 1158 3326 1159 3330
rect 1163 3326 1164 3330
rect 1158 3325 1164 3326
rect 1318 3330 1324 3331
rect 1318 3326 1319 3330
rect 1323 3326 1324 3330
rect 1318 3325 1324 3326
rect 1486 3330 1492 3331
rect 1486 3326 1487 3330
rect 1491 3326 1492 3330
rect 1486 3325 1492 3326
rect 1654 3330 1660 3331
rect 1654 3326 1655 3330
rect 1659 3326 1660 3330
rect 1654 3325 1660 3326
rect 2030 3325 2036 3326
rect 110 3321 111 3325
rect 115 3321 116 3325
rect 110 3320 116 3321
rect 2030 3321 2031 3325
rect 2035 3321 2036 3325
rect 2030 3320 2036 3321
rect 110 3308 116 3309
rect 110 3304 111 3308
rect 115 3304 116 3308
rect 110 3303 116 3304
rect 2030 3308 2036 3309
rect 2030 3304 2031 3308
rect 2035 3304 2036 3308
rect 2030 3303 2036 3304
rect 2110 3291 2116 3292
rect 150 3289 156 3290
rect 150 3285 151 3289
rect 155 3285 156 3289
rect 150 3284 156 3285
rect 286 3289 292 3290
rect 286 3285 287 3289
rect 291 3285 292 3289
rect 286 3284 292 3285
rect 462 3289 468 3290
rect 462 3285 463 3289
rect 467 3285 468 3289
rect 462 3284 468 3285
rect 638 3289 644 3290
rect 638 3285 639 3289
rect 643 3285 644 3289
rect 638 3284 644 3285
rect 814 3289 820 3290
rect 814 3285 815 3289
rect 819 3285 820 3289
rect 814 3284 820 3285
rect 990 3289 996 3290
rect 990 3285 991 3289
rect 995 3285 996 3289
rect 990 3284 996 3285
rect 1158 3289 1164 3290
rect 1158 3285 1159 3289
rect 1163 3285 1164 3289
rect 1158 3284 1164 3285
rect 1318 3289 1324 3290
rect 1318 3285 1319 3289
rect 1323 3285 1324 3289
rect 1318 3284 1324 3285
rect 1486 3289 1492 3290
rect 1486 3285 1487 3289
rect 1491 3285 1492 3289
rect 1486 3284 1492 3285
rect 1654 3289 1660 3290
rect 1654 3285 1655 3289
rect 1659 3285 1660 3289
rect 2110 3287 2111 3291
rect 2115 3287 2116 3291
rect 2110 3286 2116 3287
rect 2294 3291 2300 3292
rect 2294 3287 2295 3291
rect 2299 3287 2300 3291
rect 2294 3286 2300 3287
rect 2502 3291 2508 3292
rect 2502 3287 2503 3291
rect 2507 3287 2508 3291
rect 2502 3286 2508 3287
rect 2702 3291 2708 3292
rect 2702 3287 2703 3291
rect 2707 3287 2708 3291
rect 2702 3286 2708 3287
rect 2894 3291 2900 3292
rect 2894 3287 2895 3291
rect 2899 3287 2900 3291
rect 2894 3286 2900 3287
rect 3070 3291 3076 3292
rect 3070 3287 3071 3291
rect 3075 3287 3076 3291
rect 3070 3286 3076 3287
rect 3230 3291 3236 3292
rect 3230 3287 3231 3291
rect 3235 3287 3236 3291
rect 3230 3286 3236 3287
rect 3374 3291 3380 3292
rect 3374 3287 3375 3291
rect 3379 3287 3380 3291
rect 3374 3286 3380 3287
rect 3510 3291 3516 3292
rect 3510 3287 3511 3291
rect 3515 3287 3516 3291
rect 3510 3286 3516 3287
rect 3646 3291 3652 3292
rect 3646 3287 3647 3291
rect 3651 3287 3652 3291
rect 3646 3286 3652 3287
rect 3782 3291 3788 3292
rect 3782 3287 3783 3291
rect 3787 3287 3788 3291
rect 3782 3286 3788 3287
rect 3894 3291 3900 3292
rect 3894 3287 3895 3291
rect 3899 3287 3900 3291
rect 3894 3286 3900 3287
rect 1654 3284 1660 3285
rect 2070 3272 2076 3273
rect 2070 3268 2071 3272
rect 2075 3268 2076 3272
rect 2070 3267 2076 3268
rect 3990 3272 3996 3273
rect 3990 3268 3991 3272
rect 3995 3268 3996 3272
rect 3990 3267 3996 3268
rect 2070 3255 2076 3256
rect 2070 3251 2071 3255
rect 2075 3251 2076 3255
rect 3990 3255 3996 3256
rect 3990 3251 3991 3255
rect 3995 3251 3996 3255
rect 2070 3250 2076 3251
rect 2110 3250 2116 3251
rect 150 3247 156 3248
rect 150 3243 151 3247
rect 155 3243 156 3247
rect 150 3242 156 3243
rect 294 3247 300 3248
rect 294 3243 295 3247
rect 299 3243 300 3247
rect 294 3242 300 3243
rect 478 3247 484 3248
rect 478 3243 479 3247
rect 483 3243 484 3247
rect 478 3242 484 3243
rect 670 3247 676 3248
rect 670 3243 671 3247
rect 675 3243 676 3247
rect 670 3242 676 3243
rect 862 3247 868 3248
rect 862 3243 863 3247
rect 867 3243 868 3247
rect 862 3242 868 3243
rect 1054 3247 1060 3248
rect 1054 3243 1055 3247
rect 1059 3243 1060 3247
rect 1054 3242 1060 3243
rect 1246 3247 1252 3248
rect 1246 3243 1247 3247
rect 1251 3243 1252 3247
rect 1246 3242 1252 3243
rect 1430 3247 1436 3248
rect 1430 3243 1431 3247
rect 1435 3243 1436 3247
rect 1430 3242 1436 3243
rect 1614 3247 1620 3248
rect 1614 3243 1615 3247
rect 1619 3243 1620 3247
rect 1614 3242 1620 3243
rect 1806 3247 1812 3248
rect 1806 3243 1807 3247
rect 1811 3243 1812 3247
rect 2110 3246 2111 3250
rect 2115 3246 2116 3250
rect 2110 3245 2116 3246
rect 2294 3250 2300 3251
rect 2294 3246 2295 3250
rect 2299 3246 2300 3250
rect 2294 3245 2300 3246
rect 2502 3250 2508 3251
rect 2502 3246 2503 3250
rect 2507 3246 2508 3250
rect 2502 3245 2508 3246
rect 2702 3250 2708 3251
rect 2702 3246 2703 3250
rect 2707 3246 2708 3250
rect 2702 3245 2708 3246
rect 2894 3250 2900 3251
rect 2894 3246 2895 3250
rect 2899 3246 2900 3250
rect 2894 3245 2900 3246
rect 3070 3250 3076 3251
rect 3070 3246 3071 3250
rect 3075 3246 3076 3250
rect 3070 3245 3076 3246
rect 3230 3250 3236 3251
rect 3230 3246 3231 3250
rect 3235 3246 3236 3250
rect 3230 3245 3236 3246
rect 3374 3250 3380 3251
rect 3374 3246 3375 3250
rect 3379 3246 3380 3250
rect 3374 3245 3380 3246
rect 3510 3250 3516 3251
rect 3510 3246 3511 3250
rect 3515 3246 3516 3250
rect 3510 3245 3516 3246
rect 3646 3250 3652 3251
rect 3646 3246 3647 3250
rect 3651 3246 3652 3250
rect 3646 3245 3652 3246
rect 3782 3250 3788 3251
rect 3782 3246 3783 3250
rect 3787 3246 3788 3250
rect 3782 3245 3788 3246
rect 3894 3250 3900 3251
rect 3990 3250 3996 3251
rect 3894 3246 3895 3250
rect 3899 3246 3900 3250
rect 3894 3245 3900 3246
rect 1806 3242 1812 3243
rect 110 3228 116 3229
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 2030 3228 2036 3229
rect 2030 3224 2031 3228
rect 2035 3224 2036 3228
rect 2030 3223 2036 3224
rect 2110 3218 2116 3219
rect 2110 3214 2111 3218
rect 2115 3214 2116 3218
rect 2070 3213 2076 3214
rect 2110 3213 2116 3214
rect 2238 3218 2244 3219
rect 2238 3214 2239 3218
rect 2243 3214 2244 3218
rect 2238 3213 2244 3214
rect 2398 3218 2404 3219
rect 2398 3214 2399 3218
rect 2403 3214 2404 3218
rect 2398 3213 2404 3214
rect 2558 3218 2564 3219
rect 2558 3214 2559 3218
rect 2563 3214 2564 3218
rect 2558 3213 2564 3214
rect 2718 3218 2724 3219
rect 2718 3214 2719 3218
rect 2723 3214 2724 3218
rect 2718 3213 2724 3214
rect 2878 3218 2884 3219
rect 2878 3214 2879 3218
rect 2883 3214 2884 3218
rect 2878 3213 2884 3214
rect 3030 3218 3036 3219
rect 3030 3214 3031 3218
rect 3035 3214 3036 3218
rect 3030 3213 3036 3214
rect 3166 3218 3172 3219
rect 3166 3214 3167 3218
rect 3171 3214 3172 3218
rect 3166 3213 3172 3214
rect 3302 3218 3308 3219
rect 3302 3214 3303 3218
rect 3307 3214 3308 3218
rect 3302 3213 3308 3214
rect 3430 3218 3436 3219
rect 3430 3214 3431 3218
rect 3435 3214 3436 3218
rect 3430 3213 3436 3214
rect 3550 3218 3556 3219
rect 3550 3214 3551 3218
rect 3555 3214 3556 3218
rect 3550 3213 3556 3214
rect 3670 3218 3676 3219
rect 3670 3214 3671 3218
rect 3675 3214 3676 3218
rect 3670 3213 3676 3214
rect 3790 3218 3796 3219
rect 3790 3214 3791 3218
rect 3795 3214 3796 3218
rect 3790 3213 3796 3214
rect 3894 3218 3900 3219
rect 3894 3214 3895 3218
rect 3899 3214 3900 3218
rect 3894 3213 3900 3214
rect 3990 3213 3996 3214
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 2030 3211 2036 3212
rect 2030 3207 2031 3211
rect 2035 3207 2036 3211
rect 2070 3209 2071 3213
rect 2075 3209 2076 3213
rect 2070 3208 2076 3209
rect 3990 3209 3991 3213
rect 3995 3209 3996 3213
rect 3990 3208 3996 3209
rect 110 3206 116 3207
rect 150 3206 156 3207
rect 150 3202 151 3206
rect 155 3202 156 3206
rect 150 3201 156 3202
rect 294 3206 300 3207
rect 294 3202 295 3206
rect 299 3202 300 3206
rect 294 3201 300 3202
rect 478 3206 484 3207
rect 478 3202 479 3206
rect 483 3202 484 3206
rect 478 3201 484 3202
rect 670 3206 676 3207
rect 670 3202 671 3206
rect 675 3202 676 3206
rect 670 3201 676 3202
rect 862 3206 868 3207
rect 862 3202 863 3206
rect 867 3202 868 3206
rect 862 3201 868 3202
rect 1054 3206 1060 3207
rect 1054 3202 1055 3206
rect 1059 3202 1060 3206
rect 1054 3201 1060 3202
rect 1246 3206 1252 3207
rect 1246 3202 1247 3206
rect 1251 3202 1252 3206
rect 1246 3201 1252 3202
rect 1430 3206 1436 3207
rect 1430 3202 1431 3206
rect 1435 3202 1436 3206
rect 1430 3201 1436 3202
rect 1614 3206 1620 3207
rect 1614 3202 1615 3206
rect 1619 3202 1620 3206
rect 1614 3201 1620 3202
rect 1806 3206 1812 3207
rect 2030 3206 2036 3207
rect 1806 3202 1807 3206
rect 1811 3202 1812 3206
rect 1806 3201 1812 3202
rect 2070 3196 2076 3197
rect 2070 3192 2071 3196
rect 2075 3192 2076 3196
rect 2070 3191 2076 3192
rect 3990 3196 3996 3197
rect 3990 3192 3991 3196
rect 3995 3192 3996 3196
rect 3990 3191 3996 3192
rect 2110 3177 2116 3178
rect 2110 3173 2111 3177
rect 2115 3173 2116 3177
rect 2110 3172 2116 3173
rect 2238 3177 2244 3178
rect 2238 3173 2239 3177
rect 2243 3173 2244 3177
rect 2238 3172 2244 3173
rect 2398 3177 2404 3178
rect 2398 3173 2399 3177
rect 2403 3173 2404 3177
rect 2398 3172 2404 3173
rect 2558 3177 2564 3178
rect 2558 3173 2559 3177
rect 2563 3173 2564 3177
rect 2558 3172 2564 3173
rect 2718 3177 2724 3178
rect 2718 3173 2719 3177
rect 2723 3173 2724 3177
rect 2718 3172 2724 3173
rect 2878 3177 2884 3178
rect 2878 3173 2879 3177
rect 2883 3173 2884 3177
rect 2878 3172 2884 3173
rect 3030 3177 3036 3178
rect 3030 3173 3031 3177
rect 3035 3173 3036 3177
rect 3030 3172 3036 3173
rect 3166 3177 3172 3178
rect 3166 3173 3167 3177
rect 3171 3173 3172 3177
rect 3166 3172 3172 3173
rect 3302 3177 3308 3178
rect 3302 3173 3303 3177
rect 3307 3173 3308 3177
rect 3302 3172 3308 3173
rect 3430 3177 3436 3178
rect 3430 3173 3431 3177
rect 3435 3173 3436 3177
rect 3430 3172 3436 3173
rect 3550 3177 3556 3178
rect 3550 3173 3551 3177
rect 3555 3173 3556 3177
rect 3550 3172 3556 3173
rect 3670 3177 3676 3178
rect 3670 3173 3671 3177
rect 3675 3173 3676 3177
rect 3670 3172 3676 3173
rect 3790 3177 3796 3178
rect 3790 3173 3791 3177
rect 3795 3173 3796 3177
rect 3790 3172 3796 3173
rect 3894 3177 3900 3178
rect 3894 3173 3895 3177
rect 3899 3173 3900 3177
rect 3894 3172 3900 3173
rect 286 3162 292 3163
rect 286 3158 287 3162
rect 291 3158 292 3162
rect 110 3157 116 3158
rect 286 3157 292 3158
rect 422 3162 428 3163
rect 422 3158 423 3162
rect 427 3158 428 3162
rect 422 3157 428 3158
rect 566 3162 572 3163
rect 566 3158 567 3162
rect 571 3158 572 3162
rect 566 3157 572 3158
rect 726 3162 732 3163
rect 726 3158 727 3162
rect 731 3158 732 3162
rect 726 3157 732 3158
rect 902 3162 908 3163
rect 902 3158 903 3162
rect 907 3158 908 3162
rect 902 3157 908 3158
rect 1094 3162 1100 3163
rect 1094 3158 1095 3162
rect 1099 3158 1100 3162
rect 1094 3157 1100 3158
rect 1294 3162 1300 3163
rect 1294 3158 1295 3162
rect 1299 3158 1300 3162
rect 1294 3157 1300 3158
rect 1494 3162 1500 3163
rect 1494 3158 1495 3162
rect 1499 3158 1500 3162
rect 1494 3157 1500 3158
rect 1702 3162 1708 3163
rect 1702 3158 1703 3162
rect 1707 3158 1708 3162
rect 1702 3157 1708 3158
rect 1918 3162 1924 3163
rect 1918 3158 1919 3162
rect 1923 3158 1924 3162
rect 1918 3157 1924 3158
rect 2030 3157 2036 3158
rect 110 3153 111 3157
rect 115 3153 116 3157
rect 110 3152 116 3153
rect 2030 3153 2031 3157
rect 2035 3153 2036 3157
rect 2030 3152 2036 3153
rect 110 3140 116 3141
rect 110 3136 111 3140
rect 115 3136 116 3140
rect 110 3135 116 3136
rect 2030 3140 2036 3141
rect 2030 3136 2031 3140
rect 2035 3136 2036 3140
rect 2030 3135 2036 3136
rect 2182 3131 2188 3132
rect 2182 3127 2183 3131
rect 2187 3127 2188 3131
rect 2182 3126 2188 3127
rect 2366 3131 2372 3132
rect 2366 3127 2367 3131
rect 2371 3127 2372 3131
rect 2366 3126 2372 3127
rect 2550 3131 2556 3132
rect 2550 3127 2551 3131
rect 2555 3127 2556 3131
rect 2550 3126 2556 3127
rect 2734 3131 2740 3132
rect 2734 3127 2735 3131
rect 2739 3127 2740 3131
rect 2734 3126 2740 3127
rect 2910 3131 2916 3132
rect 2910 3127 2911 3131
rect 2915 3127 2916 3131
rect 2910 3126 2916 3127
rect 3086 3131 3092 3132
rect 3086 3127 3087 3131
rect 3091 3127 3092 3131
rect 3086 3126 3092 3127
rect 3262 3131 3268 3132
rect 3262 3127 3263 3131
rect 3267 3127 3268 3131
rect 3262 3126 3268 3127
rect 3446 3131 3452 3132
rect 3446 3127 3447 3131
rect 3451 3127 3452 3131
rect 3446 3126 3452 3127
rect 286 3121 292 3122
rect 286 3117 287 3121
rect 291 3117 292 3121
rect 286 3116 292 3117
rect 422 3121 428 3122
rect 422 3117 423 3121
rect 427 3117 428 3121
rect 422 3116 428 3117
rect 566 3121 572 3122
rect 566 3117 567 3121
rect 571 3117 572 3121
rect 566 3116 572 3117
rect 726 3121 732 3122
rect 726 3117 727 3121
rect 731 3117 732 3121
rect 726 3116 732 3117
rect 902 3121 908 3122
rect 902 3117 903 3121
rect 907 3117 908 3121
rect 902 3116 908 3117
rect 1094 3121 1100 3122
rect 1094 3117 1095 3121
rect 1099 3117 1100 3121
rect 1094 3116 1100 3117
rect 1294 3121 1300 3122
rect 1294 3117 1295 3121
rect 1299 3117 1300 3121
rect 1294 3116 1300 3117
rect 1494 3121 1500 3122
rect 1494 3117 1495 3121
rect 1499 3117 1500 3121
rect 1494 3116 1500 3117
rect 1702 3121 1708 3122
rect 1702 3117 1703 3121
rect 1707 3117 1708 3121
rect 1702 3116 1708 3117
rect 1918 3121 1924 3122
rect 1918 3117 1919 3121
rect 1923 3117 1924 3121
rect 1918 3116 1924 3117
rect 2070 3112 2076 3113
rect 2070 3108 2071 3112
rect 2075 3108 2076 3112
rect 2070 3107 2076 3108
rect 3990 3112 3996 3113
rect 3990 3108 3991 3112
rect 3995 3108 3996 3112
rect 3990 3107 3996 3108
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 3990 3095 3996 3096
rect 3990 3091 3991 3095
rect 3995 3091 3996 3095
rect 2070 3090 2076 3091
rect 2182 3090 2188 3091
rect 2182 3086 2183 3090
rect 2187 3086 2188 3090
rect 2182 3085 2188 3086
rect 2366 3090 2372 3091
rect 2366 3086 2367 3090
rect 2371 3086 2372 3090
rect 2366 3085 2372 3086
rect 2550 3090 2556 3091
rect 2550 3086 2551 3090
rect 2555 3086 2556 3090
rect 2550 3085 2556 3086
rect 2734 3090 2740 3091
rect 2734 3086 2735 3090
rect 2739 3086 2740 3090
rect 2734 3085 2740 3086
rect 2910 3090 2916 3091
rect 2910 3086 2911 3090
rect 2915 3086 2916 3090
rect 2910 3085 2916 3086
rect 3086 3090 3092 3091
rect 3086 3086 3087 3090
rect 3091 3086 3092 3090
rect 3086 3085 3092 3086
rect 3262 3090 3268 3091
rect 3262 3086 3263 3090
rect 3267 3086 3268 3090
rect 3262 3085 3268 3086
rect 3446 3090 3452 3091
rect 3990 3090 3996 3091
rect 3446 3086 3447 3090
rect 3451 3086 3452 3090
rect 3446 3085 3452 3086
rect 574 3075 580 3076
rect 574 3071 575 3075
rect 579 3071 580 3075
rect 574 3070 580 3071
rect 678 3075 684 3076
rect 678 3071 679 3075
rect 683 3071 684 3075
rect 678 3070 684 3071
rect 798 3075 804 3076
rect 798 3071 799 3075
rect 803 3071 804 3075
rect 798 3070 804 3071
rect 934 3075 940 3076
rect 934 3071 935 3075
rect 939 3071 940 3075
rect 934 3070 940 3071
rect 1078 3075 1084 3076
rect 1078 3071 1079 3075
rect 1083 3071 1084 3075
rect 1078 3070 1084 3071
rect 1230 3075 1236 3076
rect 1230 3071 1231 3075
rect 1235 3071 1236 3075
rect 1230 3070 1236 3071
rect 1390 3075 1396 3076
rect 1390 3071 1391 3075
rect 1395 3071 1396 3075
rect 1390 3070 1396 3071
rect 1558 3075 1564 3076
rect 1558 3071 1559 3075
rect 1563 3071 1564 3075
rect 1558 3070 1564 3071
rect 1726 3075 1732 3076
rect 1726 3071 1727 3075
rect 1731 3071 1732 3075
rect 1726 3070 1732 3071
rect 1902 3075 1908 3076
rect 1902 3071 1903 3075
rect 1907 3071 1908 3075
rect 1902 3070 1908 3071
rect 110 3056 116 3057
rect 110 3052 111 3056
rect 115 3052 116 3056
rect 110 3051 116 3052
rect 2030 3056 2036 3057
rect 2030 3052 2031 3056
rect 2035 3052 2036 3056
rect 2030 3051 2036 3052
rect 2350 3050 2356 3051
rect 2350 3046 2351 3050
rect 2355 3046 2356 3050
rect 2070 3045 2076 3046
rect 2350 3045 2356 3046
rect 2454 3050 2460 3051
rect 2454 3046 2455 3050
rect 2459 3046 2460 3050
rect 2454 3045 2460 3046
rect 2566 3050 2572 3051
rect 2566 3046 2567 3050
rect 2571 3046 2572 3050
rect 2566 3045 2572 3046
rect 2686 3050 2692 3051
rect 2686 3046 2687 3050
rect 2691 3046 2692 3050
rect 2686 3045 2692 3046
rect 2806 3050 2812 3051
rect 2806 3046 2807 3050
rect 2811 3046 2812 3050
rect 2806 3045 2812 3046
rect 2926 3050 2932 3051
rect 2926 3046 2927 3050
rect 2931 3046 2932 3050
rect 2926 3045 2932 3046
rect 3046 3050 3052 3051
rect 3046 3046 3047 3050
rect 3051 3046 3052 3050
rect 3046 3045 3052 3046
rect 3166 3050 3172 3051
rect 3166 3046 3167 3050
rect 3171 3046 3172 3050
rect 3166 3045 3172 3046
rect 3294 3050 3300 3051
rect 3294 3046 3295 3050
rect 3299 3046 3300 3050
rect 3294 3045 3300 3046
rect 3990 3045 3996 3046
rect 2070 3041 2071 3045
rect 2075 3041 2076 3045
rect 2070 3040 2076 3041
rect 3990 3041 3991 3045
rect 3995 3041 3996 3045
rect 3990 3040 3996 3041
rect 110 3039 116 3040
rect 110 3035 111 3039
rect 115 3035 116 3039
rect 2030 3039 2036 3040
rect 2030 3035 2031 3039
rect 2035 3035 2036 3039
rect 110 3034 116 3035
rect 574 3034 580 3035
rect 574 3030 575 3034
rect 579 3030 580 3034
rect 574 3029 580 3030
rect 678 3034 684 3035
rect 678 3030 679 3034
rect 683 3030 684 3034
rect 678 3029 684 3030
rect 798 3034 804 3035
rect 798 3030 799 3034
rect 803 3030 804 3034
rect 798 3029 804 3030
rect 934 3034 940 3035
rect 934 3030 935 3034
rect 939 3030 940 3034
rect 934 3029 940 3030
rect 1078 3034 1084 3035
rect 1078 3030 1079 3034
rect 1083 3030 1084 3034
rect 1078 3029 1084 3030
rect 1230 3034 1236 3035
rect 1230 3030 1231 3034
rect 1235 3030 1236 3034
rect 1230 3029 1236 3030
rect 1390 3034 1396 3035
rect 1390 3030 1391 3034
rect 1395 3030 1396 3034
rect 1390 3029 1396 3030
rect 1558 3034 1564 3035
rect 1558 3030 1559 3034
rect 1563 3030 1564 3034
rect 1558 3029 1564 3030
rect 1726 3034 1732 3035
rect 1726 3030 1727 3034
rect 1731 3030 1732 3034
rect 1726 3029 1732 3030
rect 1902 3034 1908 3035
rect 2030 3034 2036 3035
rect 1902 3030 1903 3034
rect 1907 3030 1908 3034
rect 1902 3029 1908 3030
rect 2070 3028 2076 3029
rect 2070 3024 2071 3028
rect 2075 3024 2076 3028
rect 2070 3023 2076 3024
rect 3990 3028 3996 3029
rect 3990 3024 3991 3028
rect 3995 3024 3996 3028
rect 3990 3023 3996 3024
rect 2350 3009 2356 3010
rect 2350 3005 2351 3009
rect 2355 3005 2356 3009
rect 2350 3004 2356 3005
rect 2454 3009 2460 3010
rect 2454 3005 2455 3009
rect 2459 3005 2460 3009
rect 2454 3004 2460 3005
rect 2566 3009 2572 3010
rect 2566 3005 2567 3009
rect 2571 3005 2572 3009
rect 2566 3004 2572 3005
rect 2686 3009 2692 3010
rect 2686 3005 2687 3009
rect 2691 3005 2692 3009
rect 2686 3004 2692 3005
rect 2806 3009 2812 3010
rect 2806 3005 2807 3009
rect 2811 3005 2812 3009
rect 2806 3004 2812 3005
rect 2926 3009 2932 3010
rect 2926 3005 2927 3009
rect 2931 3005 2932 3009
rect 2926 3004 2932 3005
rect 3046 3009 3052 3010
rect 3046 3005 3047 3009
rect 3051 3005 3052 3009
rect 3046 3004 3052 3005
rect 3166 3009 3172 3010
rect 3166 3005 3167 3009
rect 3171 3005 3172 3009
rect 3166 3004 3172 3005
rect 3294 3009 3300 3010
rect 3294 3005 3295 3009
rect 3299 3005 3300 3009
rect 3294 3004 3300 3005
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 110 2985 116 2986
rect 550 2985 556 2986
rect 654 2990 660 2991
rect 654 2986 655 2990
rect 659 2986 660 2990
rect 654 2985 660 2986
rect 758 2990 764 2991
rect 758 2986 759 2990
rect 763 2986 764 2990
rect 758 2985 764 2986
rect 870 2990 876 2991
rect 870 2986 871 2990
rect 875 2986 876 2990
rect 870 2985 876 2986
rect 990 2990 996 2991
rect 990 2986 991 2990
rect 995 2986 996 2990
rect 990 2985 996 2986
rect 1118 2990 1124 2991
rect 1118 2986 1119 2990
rect 1123 2986 1124 2990
rect 1118 2985 1124 2986
rect 1254 2990 1260 2991
rect 1254 2986 1255 2990
rect 1259 2986 1260 2990
rect 1254 2985 1260 2986
rect 1390 2990 1396 2991
rect 1390 2986 1391 2990
rect 1395 2986 1396 2990
rect 1390 2985 1396 2986
rect 1534 2990 1540 2991
rect 1534 2986 1535 2990
rect 1539 2986 1540 2990
rect 1534 2985 1540 2986
rect 1686 2990 1692 2991
rect 1686 2986 1687 2990
rect 1691 2986 1692 2990
rect 1686 2985 1692 2986
rect 2030 2985 2036 2986
rect 110 2981 111 2985
rect 115 2981 116 2985
rect 110 2980 116 2981
rect 2030 2981 2031 2985
rect 2035 2981 2036 2985
rect 2030 2980 2036 2981
rect 2494 2979 2500 2980
rect 2494 2975 2495 2979
rect 2499 2975 2500 2979
rect 2494 2974 2500 2975
rect 2598 2979 2604 2980
rect 2598 2975 2599 2979
rect 2603 2975 2604 2979
rect 2598 2974 2604 2975
rect 2702 2979 2708 2980
rect 2702 2975 2703 2979
rect 2707 2975 2708 2979
rect 2702 2974 2708 2975
rect 2806 2979 2812 2980
rect 2806 2975 2807 2979
rect 2811 2975 2812 2979
rect 2806 2974 2812 2975
rect 2910 2979 2916 2980
rect 2910 2975 2911 2979
rect 2915 2975 2916 2979
rect 2910 2974 2916 2975
rect 3014 2979 3020 2980
rect 3014 2975 3015 2979
rect 3019 2975 3020 2979
rect 3014 2974 3020 2975
rect 3118 2979 3124 2980
rect 3118 2975 3119 2979
rect 3123 2975 3124 2979
rect 3118 2974 3124 2975
rect 3222 2979 3228 2980
rect 3222 2975 3223 2979
rect 3227 2975 3228 2979
rect 3222 2974 3228 2975
rect 110 2968 116 2969
rect 110 2964 111 2968
rect 115 2964 116 2968
rect 110 2963 116 2964
rect 2030 2968 2036 2969
rect 2030 2964 2031 2968
rect 2035 2964 2036 2968
rect 2030 2963 2036 2964
rect 2070 2960 2076 2961
rect 2070 2956 2071 2960
rect 2075 2956 2076 2960
rect 2070 2955 2076 2956
rect 3990 2960 3996 2961
rect 3990 2956 3991 2960
rect 3995 2956 3996 2960
rect 3990 2955 3996 2956
rect 550 2949 556 2950
rect 550 2945 551 2949
rect 555 2945 556 2949
rect 550 2944 556 2945
rect 654 2949 660 2950
rect 654 2945 655 2949
rect 659 2945 660 2949
rect 654 2944 660 2945
rect 758 2949 764 2950
rect 758 2945 759 2949
rect 763 2945 764 2949
rect 758 2944 764 2945
rect 870 2949 876 2950
rect 870 2945 871 2949
rect 875 2945 876 2949
rect 870 2944 876 2945
rect 990 2949 996 2950
rect 990 2945 991 2949
rect 995 2945 996 2949
rect 990 2944 996 2945
rect 1118 2949 1124 2950
rect 1118 2945 1119 2949
rect 1123 2945 1124 2949
rect 1118 2944 1124 2945
rect 1254 2949 1260 2950
rect 1254 2945 1255 2949
rect 1259 2945 1260 2949
rect 1254 2944 1260 2945
rect 1390 2949 1396 2950
rect 1390 2945 1391 2949
rect 1395 2945 1396 2949
rect 1390 2944 1396 2945
rect 1534 2949 1540 2950
rect 1534 2945 1535 2949
rect 1539 2945 1540 2949
rect 1534 2944 1540 2945
rect 1686 2949 1692 2950
rect 1686 2945 1687 2949
rect 1691 2945 1692 2949
rect 1686 2944 1692 2945
rect 2070 2943 2076 2944
rect 2070 2939 2071 2943
rect 2075 2939 2076 2943
rect 3990 2943 3996 2944
rect 3990 2939 3991 2943
rect 3995 2939 3996 2943
rect 2070 2938 2076 2939
rect 2494 2938 2500 2939
rect 2494 2934 2495 2938
rect 2499 2934 2500 2938
rect 2494 2933 2500 2934
rect 2598 2938 2604 2939
rect 2598 2934 2599 2938
rect 2603 2934 2604 2938
rect 2598 2933 2604 2934
rect 2702 2938 2708 2939
rect 2702 2934 2703 2938
rect 2707 2934 2708 2938
rect 2702 2933 2708 2934
rect 2806 2938 2812 2939
rect 2806 2934 2807 2938
rect 2811 2934 2812 2938
rect 2806 2933 2812 2934
rect 2910 2938 2916 2939
rect 2910 2934 2911 2938
rect 2915 2934 2916 2938
rect 2910 2933 2916 2934
rect 3014 2938 3020 2939
rect 3014 2934 3015 2938
rect 3019 2934 3020 2938
rect 3014 2933 3020 2934
rect 3118 2938 3124 2939
rect 3118 2934 3119 2938
rect 3123 2934 3124 2938
rect 3118 2933 3124 2934
rect 3222 2938 3228 2939
rect 3990 2938 3996 2939
rect 3222 2934 3223 2938
rect 3227 2934 3228 2938
rect 3222 2933 3228 2934
rect 310 2907 316 2908
rect 310 2903 311 2907
rect 315 2903 316 2907
rect 310 2902 316 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 558 2907 564 2908
rect 558 2903 559 2907
rect 563 2903 564 2907
rect 558 2902 564 2903
rect 694 2907 700 2908
rect 694 2903 695 2907
rect 699 2903 700 2907
rect 694 2902 700 2903
rect 830 2907 836 2908
rect 830 2903 831 2907
rect 835 2903 836 2907
rect 830 2902 836 2903
rect 974 2907 980 2908
rect 974 2903 975 2907
rect 979 2903 980 2907
rect 974 2902 980 2903
rect 1118 2907 1124 2908
rect 1118 2903 1119 2907
rect 1123 2903 1124 2907
rect 1118 2902 1124 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1422 2907 1428 2908
rect 1422 2903 1423 2907
rect 1427 2903 1428 2907
rect 1422 2902 1428 2903
rect 1574 2907 1580 2908
rect 1574 2903 1575 2907
rect 1579 2903 1580 2907
rect 1574 2902 1580 2903
rect 2414 2906 2420 2907
rect 2414 2902 2415 2906
rect 2419 2902 2420 2906
rect 2070 2901 2076 2902
rect 2414 2901 2420 2902
rect 2518 2906 2524 2907
rect 2518 2902 2519 2906
rect 2523 2902 2524 2906
rect 2518 2901 2524 2902
rect 2622 2906 2628 2907
rect 2622 2902 2623 2906
rect 2627 2902 2628 2906
rect 2622 2901 2628 2902
rect 2726 2906 2732 2907
rect 2726 2902 2727 2906
rect 2731 2902 2732 2906
rect 2726 2901 2732 2902
rect 2830 2906 2836 2907
rect 2830 2902 2831 2906
rect 2835 2902 2836 2906
rect 2830 2901 2836 2902
rect 2934 2906 2940 2907
rect 2934 2902 2935 2906
rect 2939 2902 2940 2906
rect 2934 2901 2940 2902
rect 3038 2906 3044 2907
rect 3038 2902 3039 2906
rect 3043 2902 3044 2906
rect 3038 2901 3044 2902
rect 3142 2906 3148 2907
rect 3142 2902 3143 2906
rect 3147 2902 3148 2906
rect 3142 2901 3148 2902
rect 3246 2906 3252 2907
rect 3246 2902 3247 2906
rect 3251 2902 3252 2906
rect 3246 2901 3252 2902
rect 3990 2901 3996 2902
rect 2070 2897 2071 2901
rect 2075 2897 2076 2901
rect 2070 2896 2076 2897
rect 3990 2897 3991 2901
rect 3995 2897 3996 2901
rect 3990 2896 3996 2897
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 110 2883 116 2884
rect 2030 2888 2036 2889
rect 2030 2884 2031 2888
rect 2035 2884 2036 2888
rect 2030 2883 2036 2884
rect 2070 2884 2076 2885
rect 2070 2880 2071 2884
rect 2075 2880 2076 2884
rect 2070 2879 2076 2880
rect 3990 2884 3996 2885
rect 3990 2880 3991 2884
rect 3995 2880 3996 2884
rect 3990 2879 3996 2880
rect 110 2871 116 2872
rect 110 2867 111 2871
rect 115 2867 116 2871
rect 2030 2871 2036 2872
rect 2030 2867 2031 2871
rect 2035 2867 2036 2871
rect 110 2866 116 2867
rect 310 2866 316 2867
rect 310 2862 311 2866
rect 315 2862 316 2866
rect 310 2861 316 2862
rect 430 2866 436 2867
rect 430 2862 431 2866
rect 435 2862 436 2866
rect 430 2861 436 2862
rect 558 2866 564 2867
rect 558 2862 559 2866
rect 563 2862 564 2866
rect 558 2861 564 2862
rect 694 2866 700 2867
rect 694 2862 695 2866
rect 699 2862 700 2866
rect 694 2861 700 2862
rect 830 2866 836 2867
rect 830 2862 831 2866
rect 835 2862 836 2866
rect 830 2861 836 2862
rect 974 2866 980 2867
rect 974 2862 975 2866
rect 979 2862 980 2866
rect 974 2861 980 2862
rect 1118 2866 1124 2867
rect 1118 2862 1119 2866
rect 1123 2862 1124 2866
rect 1118 2861 1124 2862
rect 1270 2866 1276 2867
rect 1270 2862 1271 2866
rect 1275 2862 1276 2866
rect 1270 2861 1276 2862
rect 1422 2866 1428 2867
rect 1422 2862 1423 2866
rect 1427 2862 1428 2866
rect 1422 2861 1428 2862
rect 1574 2866 1580 2867
rect 2030 2866 2036 2867
rect 1574 2862 1575 2866
rect 1579 2862 1580 2866
rect 1574 2861 1580 2862
rect 2414 2865 2420 2866
rect 2414 2861 2415 2865
rect 2419 2861 2420 2865
rect 2414 2860 2420 2861
rect 2518 2865 2524 2866
rect 2518 2861 2519 2865
rect 2523 2861 2524 2865
rect 2518 2860 2524 2861
rect 2622 2865 2628 2866
rect 2622 2861 2623 2865
rect 2627 2861 2628 2865
rect 2622 2860 2628 2861
rect 2726 2865 2732 2866
rect 2726 2861 2727 2865
rect 2731 2861 2732 2865
rect 2726 2860 2732 2861
rect 2830 2865 2836 2866
rect 2830 2861 2831 2865
rect 2835 2861 2836 2865
rect 2830 2860 2836 2861
rect 2934 2865 2940 2866
rect 2934 2861 2935 2865
rect 2939 2861 2940 2865
rect 2934 2860 2940 2861
rect 3038 2865 3044 2866
rect 3038 2861 3039 2865
rect 3043 2861 3044 2865
rect 3038 2860 3044 2861
rect 3142 2865 3148 2866
rect 3142 2861 3143 2865
rect 3147 2861 3148 2865
rect 3142 2860 3148 2861
rect 3246 2865 3252 2866
rect 3246 2861 3247 2865
rect 3251 2861 3252 2865
rect 3246 2860 3252 2861
rect 2406 2831 2412 2832
rect 2406 2827 2407 2831
rect 2411 2827 2412 2831
rect 2406 2826 2412 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2614 2831 2620 2832
rect 2614 2827 2615 2831
rect 2619 2827 2620 2831
rect 2614 2826 2620 2827
rect 2718 2831 2724 2832
rect 2718 2827 2719 2831
rect 2723 2827 2724 2831
rect 2718 2826 2724 2827
rect 2822 2831 2828 2832
rect 2822 2827 2823 2831
rect 2827 2827 2828 2831
rect 2822 2826 2828 2827
rect 2926 2831 2932 2832
rect 2926 2827 2927 2831
rect 2931 2827 2932 2831
rect 2926 2826 2932 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3134 2831 3140 2832
rect 3134 2827 3135 2831
rect 3139 2827 3140 2831
rect 3134 2826 3140 2827
rect 3238 2831 3244 2832
rect 3238 2827 3239 2831
rect 3243 2827 3244 2831
rect 3238 2826 3244 2827
rect 150 2818 156 2819
rect 150 2814 151 2818
rect 155 2814 156 2818
rect 110 2813 116 2814
rect 150 2813 156 2814
rect 310 2818 316 2819
rect 310 2814 311 2818
rect 315 2814 316 2818
rect 310 2813 316 2814
rect 470 2818 476 2819
rect 470 2814 471 2818
rect 475 2814 476 2818
rect 470 2813 476 2814
rect 622 2818 628 2819
rect 622 2814 623 2818
rect 627 2814 628 2818
rect 622 2813 628 2814
rect 766 2818 772 2819
rect 766 2814 767 2818
rect 771 2814 772 2818
rect 766 2813 772 2814
rect 902 2818 908 2819
rect 902 2814 903 2818
rect 907 2814 908 2818
rect 902 2813 908 2814
rect 1030 2818 1036 2819
rect 1030 2814 1031 2818
rect 1035 2814 1036 2818
rect 1030 2813 1036 2814
rect 1158 2818 1164 2819
rect 1158 2814 1159 2818
rect 1163 2814 1164 2818
rect 1158 2813 1164 2814
rect 1286 2818 1292 2819
rect 1286 2814 1287 2818
rect 1291 2814 1292 2818
rect 1286 2813 1292 2814
rect 1414 2818 1420 2819
rect 1414 2814 1415 2818
rect 1419 2814 1420 2818
rect 1414 2813 1420 2814
rect 2030 2813 2036 2814
rect 110 2809 111 2813
rect 115 2809 116 2813
rect 110 2808 116 2809
rect 2030 2809 2031 2813
rect 2035 2809 2036 2813
rect 2030 2808 2036 2809
rect 2070 2812 2076 2813
rect 2070 2808 2071 2812
rect 2075 2808 2076 2812
rect 2070 2807 2076 2808
rect 3990 2812 3996 2813
rect 3990 2808 3991 2812
rect 3995 2808 3996 2812
rect 3990 2807 3996 2808
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 2030 2796 2036 2797
rect 2030 2792 2031 2796
rect 2035 2792 2036 2796
rect 2030 2791 2036 2792
rect 2070 2795 2076 2796
rect 2070 2791 2071 2795
rect 2075 2791 2076 2795
rect 3990 2795 3996 2796
rect 3990 2791 3991 2795
rect 3995 2791 3996 2795
rect 2070 2790 2076 2791
rect 2406 2790 2412 2791
rect 2406 2786 2407 2790
rect 2411 2786 2412 2790
rect 2406 2785 2412 2786
rect 2510 2790 2516 2791
rect 2510 2786 2511 2790
rect 2515 2786 2516 2790
rect 2510 2785 2516 2786
rect 2614 2790 2620 2791
rect 2614 2786 2615 2790
rect 2619 2786 2620 2790
rect 2614 2785 2620 2786
rect 2718 2790 2724 2791
rect 2718 2786 2719 2790
rect 2723 2786 2724 2790
rect 2718 2785 2724 2786
rect 2822 2790 2828 2791
rect 2822 2786 2823 2790
rect 2827 2786 2828 2790
rect 2822 2785 2828 2786
rect 2926 2790 2932 2791
rect 2926 2786 2927 2790
rect 2931 2786 2932 2790
rect 2926 2785 2932 2786
rect 3030 2790 3036 2791
rect 3030 2786 3031 2790
rect 3035 2786 3036 2790
rect 3030 2785 3036 2786
rect 3134 2790 3140 2791
rect 3134 2786 3135 2790
rect 3139 2786 3140 2790
rect 3134 2785 3140 2786
rect 3238 2790 3244 2791
rect 3990 2790 3996 2791
rect 3238 2786 3239 2790
rect 3243 2786 3244 2790
rect 3238 2785 3244 2786
rect 150 2777 156 2778
rect 150 2773 151 2777
rect 155 2773 156 2777
rect 150 2772 156 2773
rect 310 2777 316 2778
rect 310 2773 311 2777
rect 315 2773 316 2777
rect 310 2772 316 2773
rect 470 2777 476 2778
rect 470 2773 471 2777
rect 475 2773 476 2777
rect 470 2772 476 2773
rect 622 2777 628 2778
rect 622 2773 623 2777
rect 627 2773 628 2777
rect 622 2772 628 2773
rect 766 2777 772 2778
rect 766 2773 767 2777
rect 771 2773 772 2777
rect 766 2772 772 2773
rect 902 2777 908 2778
rect 902 2773 903 2777
rect 907 2773 908 2777
rect 902 2772 908 2773
rect 1030 2777 1036 2778
rect 1030 2773 1031 2777
rect 1035 2773 1036 2777
rect 1030 2772 1036 2773
rect 1158 2777 1164 2778
rect 1158 2773 1159 2777
rect 1163 2773 1164 2777
rect 1158 2772 1164 2773
rect 1286 2777 1292 2778
rect 1286 2773 1287 2777
rect 1291 2773 1292 2777
rect 1286 2772 1292 2773
rect 1414 2777 1420 2778
rect 1414 2773 1415 2777
rect 1419 2773 1420 2777
rect 1414 2772 1420 2773
rect 2302 2750 2308 2751
rect 2302 2746 2303 2750
rect 2307 2746 2308 2750
rect 2070 2745 2076 2746
rect 2302 2745 2308 2746
rect 2414 2750 2420 2751
rect 2414 2746 2415 2750
rect 2419 2746 2420 2750
rect 2414 2745 2420 2746
rect 2534 2750 2540 2751
rect 2534 2746 2535 2750
rect 2539 2746 2540 2750
rect 2534 2745 2540 2746
rect 2654 2750 2660 2751
rect 2654 2746 2655 2750
rect 2659 2746 2660 2750
rect 2654 2745 2660 2746
rect 2774 2750 2780 2751
rect 2774 2746 2775 2750
rect 2779 2746 2780 2750
rect 2774 2745 2780 2746
rect 2894 2750 2900 2751
rect 2894 2746 2895 2750
rect 2899 2746 2900 2750
rect 2894 2745 2900 2746
rect 3014 2750 3020 2751
rect 3014 2746 3015 2750
rect 3019 2746 3020 2750
rect 3014 2745 3020 2746
rect 3142 2750 3148 2751
rect 3142 2746 3143 2750
rect 3147 2746 3148 2750
rect 3142 2745 3148 2746
rect 3270 2750 3276 2751
rect 3270 2746 3271 2750
rect 3275 2746 3276 2750
rect 3270 2745 3276 2746
rect 3398 2750 3404 2751
rect 3398 2746 3399 2750
rect 3403 2746 3404 2750
rect 3398 2745 3404 2746
rect 3990 2745 3996 2746
rect 2070 2741 2071 2745
rect 2075 2741 2076 2745
rect 2070 2740 2076 2741
rect 3990 2741 3991 2745
rect 3995 2741 3996 2745
rect 3990 2740 3996 2741
rect 150 2731 156 2732
rect 150 2727 151 2731
rect 155 2727 156 2731
rect 150 2726 156 2727
rect 302 2731 308 2732
rect 302 2727 303 2731
rect 307 2727 308 2731
rect 302 2726 308 2727
rect 470 2731 476 2732
rect 470 2727 471 2731
rect 475 2727 476 2731
rect 470 2726 476 2727
rect 622 2731 628 2732
rect 622 2727 623 2731
rect 627 2727 628 2731
rect 622 2726 628 2727
rect 766 2731 772 2732
rect 766 2727 767 2731
rect 771 2727 772 2731
rect 766 2726 772 2727
rect 902 2731 908 2732
rect 902 2727 903 2731
rect 907 2727 908 2731
rect 902 2726 908 2727
rect 1038 2731 1044 2732
rect 1038 2727 1039 2731
rect 1043 2727 1044 2731
rect 1038 2726 1044 2727
rect 1166 2731 1172 2732
rect 1166 2727 1167 2731
rect 1171 2727 1172 2731
rect 1166 2726 1172 2727
rect 1294 2731 1300 2732
rect 1294 2727 1295 2731
rect 1299 2727 1300 2731
rect 1294 2726 1300 2727
rect 1422 2731 1428 2732
rect 1422 2727 1423 2731
rect 1427 2727 1428 2731
rect 1422 2726 1428 2727
rect 2070 2728 2076 2729
rect 2070 2724 2071 2728
rect 2075 2724 2076 2728
rect 2070 2723 2076 2724
rect 3990 2728 3996 2729
rect 3990 2724 3991 2728
rect 3995 2724 3996 2728
rect 3990 2723 3996 2724
rect 110 2712 116 2713
rect 110 2708 111 2712
rect 115 2708 116 2712
rect 110 2707 116 2708
rect 2030 2712 2036 2713
rect 2030 2708 2031 2712
rect 2035 2708 2036 2712
rect 2030 2707 2036 2708
rect 2302 2709 2308 2710
rect 2302 2705 2303 2709
rect 2307 2705 2308 2709
rect 2302 2704 2308 2705
rect 2414 2709 2420 2710
rect 2414 2705 2415 2709
rect 2419 2705 2420 2709
rect 2414 2704 2420 2705
rect 2534 2709 2540 2710
rect 2534 2705 2535 2709
rect 2539 2705 2540 2709
rect 2534 2704 2540 2705
rect 2654 2709 2660 2710
rect 2654 2705 2655 2709
rect 2659 2705 2660 2709
rect 2654 2704 2660 2705
rect 2774 2709 2780 2710
rect 2774 2705 2775 2709
rect 2779 2705 2780 2709
rect 2774 2704 2780 2705
rect 2894 2709 2900 2710
rect 2894 2705 2895 2709
rect 2899 2705 2900 2709
rect 2894 2704 2900 2705
rect 3014 2709 3020 2710
rect 3014 2705 3015 2709
rect 3019 2705 3020 2709
rect 3014 2704 3020 2705
rect 3142 2709 3148 2710
rect 3142 2705 3143 2709
rect 3147 2705 3148 2709
rect 3142 2704 3148 2705
rect 3270 2709 3276 2710
rect 3270 2705 3271 2709
rect 3275 2705 3276 2709
rect 3270 2704 3276 2705
rect 3398 2709 3404 2710
rect 3398 2705 3399 2709
rect 3403 2705 3404 2709
rect 3398 2704 3404 2705
rect 110 2695 116 2696
rect 110 2691 111 2695
rect 115 2691 116 2695
rect 2030 2695 2036 2696
rect 2030 2691 2031 2695
rect 2035 2691 2036 2695
rect 110 2690 116 2691
rect 150 2690 156 2691
rect 150 2686 151 2690
rect 155 2686 156 2690
rect 150 2685 156 2686
rect 302 2690 308 2691
rect 302 2686 303 2690
rect 307 2686 308 2690
rect 302 2685 308 2686
rect 470 2690 476 2691
rect 470 2686 471 2690
rect 475 2686 476 2690
rect 470 2685 476 2686
rect 622 2690 628 2691
rect 622 2686 623 2690
rect 627 2686 628 2690
rect 622 2685 628 2686
rect 766 2690 772 2691
rect 766 2686 767 2690
rect 771 2686 772 2690
rect 766 2685 772 2686
rect 902 2690 908 2691
rect 902 2686 903 2690
rect 907 2686 908 2690
rect 902 2685 908 2686
rect 1038 2690 1044 2691
rect 1038 2686 1039 2690
rect 1043 2686 1044 2690
rect 1038 2685 1044 2686
rect 1166 2690 1172 2691
rect 1166 2686 1167 2690
rect 1171 2686 1172 2690
rect 1166 2685 1172 2686
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1422 2690 1428 2691
rect 2030 2690 2036 2691
rect 1422 2686 1423 2690
rect 1427 2686 1428 2690
rect 1422 2685 1428 2686
rect 2150 2663 2156 2664
rect 2150 2659 2151 2663
rect 2155 2659 2156 2663
rect 2150 2658 2156 2659
rect 2302 2663 2308 2664
rect 2302 2659 2303 2663
rect 2307 2659 2308 2663
rect 2302 2658 2308 2659
rect 2462 2663 2468 2664
rect 2462 2659 2463 2663
rect 2467 2659 2468 2663
rect 2462 2658 2468 2659
rect 2622 2663 2628 2664
rect 2622 2659 2623 2663
rect 2627 2659 2628 2663
rect 2622 2658 2628 2659
rect 2790 2663 2796 2664
rect 2790 2659 2791 2663
rect 2795 2659 2796 2663
rect 2790 2658 2796 2659
rect 2950 2663 2956 2664
rect 2950 2659 2951 2663
rect 2955 2659 2956 2663
rect 2950 2658 2956 2659
rect 3110 2663 3116 2664
rect 3110 2659 3111 2663
rect 3115 2659 3116 2663
rect 3110 2658 3116 2659
rect 3262 2663 3268 2664
rect 3262 2659 3263 2663
rect 3267 2659 3268 2663
rect 3262 2658 3268 2659
rect 3414 2663 3420 2664
rect 3414 2659 3415 2663
rect 3419 2659 3420 2663
rect 3414 2658 3420 2659
rect 3574 2663 3580 2664
rect 3574 2659 3575 2663
rect 3579 2659 3580 2663
rect 3574 2658 3580 2659
rect 150 2646 156 2647
rect 150 2642 151 2646
rect 155 2642 156 2646
rect 110 2641 116 2642
rect 150 2641 156 2642
rect 318 2646 324 2647
rect 318 2642 319 2646
rect 323 2642 324 2646
rect 318 2641 324 2642
rect 510 2646 516 2647
rect 510 2642 511 2646
rect 515 2642 516 2646
rect 510 2641 516 2642
rect 702 2646 708 2647
rect 702 2642 703 2646
rect 707 2642 708 2646
rect 702 2641 708 2642
rect 886 2646 892 2647
rect 886 2642 887 2646
rect 891 2642 892 2646
rect 886 2641 892 2642
rect 1062 2646 1068 2647
rect 1062 2642 1063 2646
rect 1067 2642 1068 2646
rect 1062 2641 1068 2642
rect 1230 2646 1236 2647
rect 1230 2642 1231 2646
rect 1235 2642 1236 2646
rect 1230 2641 1236 2642
rect 1390 2646 1396 2647
rect 1390 2642 1391 2646
rect 1395 2642 1396 2646
rect 1390 2641 1396 2642
rect 1550 2646 1556 2647
rect 1550 2642 1551 2646
rect 1555 2642 1556 2646
rect 1550 2641 1556 2642
rect 1710 2646 1716 2647
rect 1710 2642 1711 2646
rect 1715 2642 1716 2646
rect 2070 2644 2076 2645
rect 1710 2641 1716 2642
rect 2030 2641 2036 2642
rect 110 2637 111 2641
rect 115 2637 116 2641
rect 110 2636 116 2637
rect 2030 2637 2031 2641
rect 2035 2637 2036 2641
rect 2070 2640 2071 2644
rect 2075 2640 2076 2644
rect 2070 2639 2076 2640
rect 3990 2644 3996 2645
rect 3990 2640 3991 2644
rect 3995 2640 3996 2644
rect 3990 2639 3996 2640
rect 2030 2636 2036 2637
rect 2070 2627 2076 2628
rect 110 2624 116 2625
rect 110 2620 111 2624
rect 115 2620 116 2624
rect 110 2619 116 2620
rect 2030 2624 2036 2625
rect 2030 2620 2031 2624
rect 2035 2620 2036 2624
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 3990 2627 3996 2628
rect 3990 2623 3991 2627
rect 3995 2623 3996 2627
rect 2070 2622 2076 2623
rect 2150 2622 2156 2623
rect 2030 2619 2036 2620
rect 2150 2618 2151 2622
rect 2155 2618 2156 2622
rect 2150 2617 2156 2618
rect 2302 2622 2308 2623
rect 2302 2618 2303 2622
rect 2307 2618 2308 2622
rect 2302 2617 2308 2618
rect 2462 2622 2468 2623
rect 2462 2618 2463 2622
rect 2467 2618 2468 2622
rect 2462 2617 2468 2618
rect 2622 2622 2628 2623
rect 2622 2618 2623 2622
rect 2627 2618 2628 2622
rect 2622 2617 2628 2618
rect 2790 2622 2796 2623
rect 2790 2618 2791 2622
rect 2795 2618 2796 2622
rect 2790 2617 2796 2618
rect 2950 2622 2956 2623
rect 2950 2618 2951 2622
rect 2955 2618 2956 2622
rect 2950 2617 2956 2618
rect 3110 2622 3116 2623
rect 3110 2618 3111 2622
rect 3115 2618 3116 2622
rect 3110 2617 3116 2618
rect 3262 2622 3268 2623
rect 3262 2618 3263 2622
rect 3267 2618 3268 2622
rect 3262 2617 3268 2618
rect 3414 2622 3420 2623
rect 3414 2618 3415 2622
rect 3419 2618 3420 2622
rect 3414 2617 3420 2618
rect 3574 2622 3580 2623
rect 3990 2622 3996 2623
rect 3574 2618 3575 2622
rect 3579 2618 3580 2622
rect 3574 2617 3580 2618
rect 150 2605 156 2606
rect 150 2601 151 2605
rect 155 2601 156 2605
rect 150 2600 156 2601
rect 318 2605 324 2606
rect 318 2601 319 2605
rect 323 2601 324 2605
rect 318 2600 324 2601
rect 510 2605 516 2606
rect 510 2601 511 2605
rect 515 2601 516 2605
rect 510 2600 516 2601
rect 702 2605 708 2606
rect 702 2601 703 2605
rect 707 2601 708 2605
rect 702 2600 708 2601
rect 886 2605 892 2606
rect 886 2601 887 2605
rect 891 2601 892 2605
rect 886 2600 892 2601
rect 1062 2605 1068 2606
rect 1062 2601 1063 2605
rect 1067 2601 1068 2605
rect 1062 2600 1068 2601
rect 1230 2605 1236 2606
rect 1230 2601 1231 2605
rect 1235 2601 1236 2605
rect 1230 2600 1236 2601
rect 1390 2605 1396 2606
rect 1390 2601 1391 2605
rect 1395 2601 1396 2605
rect 1390 2600 1396 2601
rect 1550 2605 1556 2606
rect 1550 2601 1551 2605
rect 1555 2601 1556 2605
rect 1550 2600 1556 2601
rect 1710 2605 1716 2606
rect 1710 2601 1711 2605
rect 1715 2601 1716 2605
rect 1710 2600 1716 2601
rect 2110 2582 2116 2583
rect 2110 2578 2111 2582
rect 2115 2578 2116 2582
rect 2070 2577 2076 2578
rect 2110 2577 2116 2578
rect 2326 2582 2332 2583
rect 2326 2578 2327 2582
rect 2331 2578 2332 2582
rect 2326 2577 2332 2578
rect 2558 2582 2564 2583
rect 2558 2578 2559 2582
rect 2563 2578 2564 2582
rect 2558 2577 2564 2578
rect 2782 2582 2788 2583
rect 2782 2578 2783 2582
rect 2787 2578 2788 2582
rect 2782 2577 2788 2578
rect 2998 2582 3004 2583
rect 2998 2578 2999 2582
rect 3003 2578 3004 2582
rect 2998 2577 3004 2578
rect 3198 2582 3204 2583
rect 3198 2578 3199 2582
rect 3203 2578 3204 2582
rect 3198 2577 3204 2578
rect 3382 2582 3388 2583
rect 3382 2578 3383 2582
rect 3387 2578 3388 2582
rect 3382 2577 3388 2578
rect 3558 2582 3564 2583
rect 3558 2578 3559 2582
rect 3563 2578 3564 2582
rect 3558 2577 3564 2578
rect 3734 2582 3740 2583
rect 3734 2578 3735 2582
rect 3739 2578 3740 2582
rect 3734 2577 3740 2578
rect 3894 2582 3900 2583
rect 3894 2578 3895 2582
rect 3899 2578 3900 2582
rect 3894 2577 3900 2578
rect 3990 2577 3996 2578
rect 2070 2573 2071 2577
rect 2075 2573 2076 2577
rect 2070 2572 2076 2573
rect 3990 2573 3991 2577
rect 3995 2573 3996 2577
rect 3990 2572 3996 2573
rect 2070 2560 2076 2561
rect 278 2559 284 2560
rect 278 2555 279 2559
rect 283 2555 284 2559
rect 278 2554 284 2555
rect 462 2559 468 2560
rect 462 2555 463 2559
rect 467 2555 468 2559
rect 462 2554 468 2555
rect 662 2559 668 2560
rect 662 2555 663 2559
rect 667 2555 668 2559
rect 662 2554 668 2555
rect 862 2559 868 2560
rect 862 2555 863 2559
rect 867 2555 868 2559
rect 862 2554 868 2555
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1254 2559 1260 2560
rect 1254 2555 1255 2559
rect 1259 2555 1260 2559
rect 1254 2554 1260 2555
rect 1430 2559 1436 2560
rect 1430 2555 1431 2559
rect 1435 2555 1436 2559
rect 1430 2554 1436 2555
rect 1606 2559 1612 2560
rect 1606 2555 1607 2559
rect 1611 2555 1612 2559
rect 1606 2554 1612 2555
rect 1782 2559 1788 2560
rect 1782 2555 1783 2559
rect 1787 2555 1788 2559
rect 1782 2554 1788 2555
rect 1934 2559 1940 2560
rect 1934 2555 1935 2559
rect 1939 2555 1940 2559
rect 2070 2556 2071 2560
rect 2075 2556 2076 2560
rect 2070 2555 2076 2556
rect 3990 2560 3996 2561
rect 3990 2556 3991 2560
rect 3995 2556 3996 2560
rect 3990 2555 3996 2556
rect 1934 2554 1940 2555
rect 2110 2541 2116 2542
rect 110 2540 116 2541
rect 110 2536 111 2540
rect 115 2536 116 2540
rect 110 2535 116 2536
rect 2030 2540 2036 2541
rect 2030 2536 2031 2540
rect 2035 2536 2036 2540
rect 2110 2537 2111 2541
rect 2115 2537 2116 2541
rect 2110 2536 2116 2537
rect 2326 2541 2332 2542
rect 2326 2537 2327 2541
rect 2331 2537 2332 2541
rect 2326 2536 2332 2537
rect 2558 2541 2564 2542
rect 2558 2537 2559 2541
rect 2563 2537 2564 2541
rect 2558 2536 2564 2537
rect 2782 2541 2788 2542
rect 2782 2537 2783 2541
rect 2787 2537 2788 2541
rect 2782 2536 2788 2537
rect 2998 2541 3004 2542
rect 2998 2537 2999 2541
rect 3003 2537 3004 2541
rect 2998 2536 3004 2537
rect 3198 2541 3204 2542
rect 3198 2537 3199 2541
rect 3203 2537 3204 2541
rect 3198 2536 3204 2537
rect 3382 2541 3388 2542
rect 3382 2537 3383 2541
rect 3387 2537 3388 2541
rect 3382 2536 3388 2537
rect 3558 2541 3564 2542
rect 3558 2537 3559 2541
rect 3563 2537 3564 2541
rect 3558 2536 3564 2537
rect 3734 2541 3740 2542
rect 3734 2537 3735 2541
rect 3739 2537 3740 2541
rect 3734 2536 3740 2537
rect 3894 2541 3900 2542
rect 3894 2537 3895 2541
rect 3899 2537 3900 2541
rect 3894 2536 3900 2537
rect 2030 2535 2036 2536
rect 110 2523 116 2524
rect 110 2519 111 2523
rect 115 2519 116 2523
rect 2030 2523 2036 2524
rect 2030 2519 2031 2523
rect 2035 2519 2036 2523
rect 110 2518 116 2519
rect 278 2518 284 2519
rect 278 2514 279 2518
rect 283 2514 284 2518
rect 278 2513 284 2514
rect 462 2518 468 2519
rect 462 2514 463 2518
rect 467 2514 468 2518
rect 462 2513 468 2514
rect 662 2518 668 2519
rect 662 2514 663 2518
rect 667 2514 668 2518
rect 662 2513 668 2514
rect 862 2518 868 2519
rect 862 2514 863 2518
rect 867 2514 868 2518
rect 862 2513 868 2514
rect 1062 2518 1068 2519
rect 1062 2514 1063 2518
rect 1067 2514 1068 2518
rect 1062 2513 1068 2514
rect 1254 2518 1260 2519
rect 1254 2514 1255 2518
rect 1259 2514 1260 2518
rect 1254 2513 1260 2514
rect 1430 2518 1436 2519
rect 1430 2514 1431 2518
rect 1435 2514 1436 2518
rect 1430 2513 1436 2514
rect 1606 2518 1612 2519
rect 1606 2514 1607 2518
rect 1611 2514 1612 2518
rect 1606 2513 1612 2514
rect 1782 2518 1788 2519
rect 1782 2514 1783 2518
rect 1787 2514 1788 2518
rect 1782 2513 1788 2514
rect 1934 2518 1940 2519
rect 2030 2518 2036 2519
rect 1934 2514 1935 2518
rect 1939 2514 1940 2518
rect 1934 2513 1940 2514
rect 2110 2511 2116 2512
rect 2110 2507 2111 2511
rect 2115 2507 2116 2511
rect 2110 2506 2116 2507
rect 2254 2511 2260 2512
rect 2254 2507 2255 2511
rect 2259 2507 2260 2511
rect 2254 2506 2260 2507
rect 2438 2511 2444 2512
rect 2438 2507 2439 2511
rect 2443 2507 2444 2511
rect 2438 2506 2444 2507
rect 2630 2511 2636 2512
rect 2630 2507 2631 2511
rect 2635 2507 2636 2511
rect 2630 2506 2636 2507
rect 2822 2511 2828 2512
rect 2822 2507 2823 2511
rect 2827 2507 2828 2511
rect 2822 2506 2828 2507
rect 3006 2511 3012 2512
rect 3006 2507 3007 2511
rect 3011 2507 3012 2511
rect 3006 2506 3012 2507
rect 3174 2511 3180 2512
rect 3174 2507 3175 2511
rect 3179 2507 3180 2511
rect 3174 2506 3180 2507
rect 3334 2511 3340 2512
rect 3334 2507 3335 2511
rect 3339 2507 3340 2511
rect 3334 2506 3340 2507
rect 3486 2511 3492 2512
rect 3486 2507 3487 2511
rect 3491 2507 3492 2511
rect 3486 2506 3492 2507
rect 3630 2511 3636 2512
rect 3630 2507 3631 2511
rect 3635 2507 3636 2511
rect 3630 2506 3636 2507
rect 3774 2511 3780 2512
rect 3774 2507 3775 2511
rect 3779 2507 3780 2511
rect 3774 2506 3780 2507
rect 3894 2511 3900 2512
rect 3894 2507 3895 2511
rect 3899 2507 3900 2511
rect 3894 2506 3900 2507
rect 2070 2492 2076 2493
rect 2070 2488 2071 2492
rect 2075 2488 2076 2492
rect 2070 2487 2076 2488
rect 3990 2492 3996 2493
rect 3990 2488 3991 2492
rect 3995 2488 3996 2492
rect 3990 2487 3996 2488
rect 2070 2475 2076 2476
rect 2070 2471 2071 2475
rect 2075 2471 2076 2475
rect 3990 2475 3996 2476
rect 3990 2471 3991 2475
rect 3995 2471 3996 2475
rect 310 2470 316 2471
rect 310 2466 311 2470
rect 315 2466 316 2470
rect 110 2465 116 2466
rect 310 2465 316 2466
rect 470 2470 476 2471
rect 470 2466 471 2470
rect 475 2466 476 2470
rect 470 2465 476 2466
rect 646 2470 652 2471
rect 646 2466 647 2470
rect 651 2466 652 2470
rect 646 2465 652 2466
rect 830 2470 836 2471
rect 830 2466 831 2470
rect 835 2466 836 2470
rect 830 2465 836 2466
rect 1014 2470 1020 2471
rect 1014 2466 1015 2470
rect 1019 2466 1020 2470
rect 1014 2465 1020 2466
rect 1190 2470 1196 2471
rect 1190 2466 1191 2470
rect 1195 2466 1196 2470
rect 1190 2465 1196 2466
rect 1366 2470 1372 2471
rect 1366 2466 1367 2470
rect 1371 2466 1372 2470
rect 1366 2465 1372 2466
rect 1534 2470 1540 2471
rect 1534 2466 1535 2470
rect 1539 2466 1540 2470
rect 1534 2465 1540 2466
rect 1702 2470 1708 2471
rect 1702 2466 1703 2470
rect 1707 2466 1708 2470
rect 1702 2465 1708 2466
rect 1870 2470 1876 2471
rect 2070 2470 2076 2471
rect 2110 2470 2116 2471
rect 1870 2466 1871 2470
rect 1875 2466 1876 2470
rect 2110 2466 2111 2470
rect 2115 2466 2116 2470
rect 1870 2465 1876 2466
rect 2030 2465 2036 2466
rect 2110 2465 2116 2466
rect 2254 2470 2260 2471
rect 2254 2466 2255 2470
rect 2259 2466 2260 2470
rect 2254 2465 2260 2466
rect 2438 2470 2444 2471
rect 2438 2466 2439 2470
rect 2443 2466 2444 2470
rect 2438 2465 2444 2466
rect 2630 2470 2636 2471
rect 2630 2466 2631 2470
rect 2635 2466 2636 2470
rect 2630 2465 2636 2466
rect 2822 2470 2828 2471
rect 2822 2466 2823 2470
rect 2827 2466 2828 2470
rect 2822 2465 2828 2466
rect 3006 2470 3012 2471
rect 3006 2466 3007 2470
rect 3011 2466 3012 2470
rect 3006 2465 3012 2466
rect 3174 2470 3180 2471
rect 3174 2466 3175 2470
rect 3179 2466 3180 2470
rect 3174 2465 3180 2466
rect 3334 2470 3340 2471
rect 3334 2466 3335 2470
rect 3339 2466 3340 2470
rect 3334 2465 3340 2466
rect 3486 2470 3492 2471
rect 3486 2466 3487 2470
rect 3491 2466 3492 2470
rect 3486 2465 3492 2466
rect 3630 2470 3636 2471
rect 3630 2466 3631 2470
rect 3635 2466 3636 2470
rect 3630 2465 3636 2466
rect 3774 2470 3780 2471
rect 3774 2466 3775 2470
rect 3779 2466 3780 2470
rect 3774 2465 3780 2466
rect 3894 2470 3900 2471
rect 3990 2470 3996 2471
rect 3894 2466 3895 2470
rect 3899 2466 3900 2470
rect 3894 2465 3900 2466
rect 110 2461 111 2465
rect 115 2461 116 2465
rect 110 2460 116 2461
rect 2030 2461 2031 2465
rect 2035 2461 2036 2465
rect 2030 2460 2036 2461
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 110 2443 116 2444
rect 2030 2448 2036 2449
rect 2030 2444 2031 2448
rect 2035 2444 2036 2448
rect 2030 2443 2036 2444
rect 2110 2430 2116 2431
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 470 2429 476 2430
rect 470 2425 471 2429
rect 475 2425 476 2429
rect 470 2424 476 2425
rect 646 2429 652 2430
rect 646 2425 647 2429
rect 651 2425 652 2429
rect 646 2424 652 2425
rect 830 2429 836 2430
rect 830 2425 831 2429
rect 835 2425 836 2429
rect 830 2424 836 2425
rect 1014 2429 1020 2430
rect 1014 2425 1015 2429
rect 1019 2425 1020 2429
rect 1014 2424 1020 2425
rect 1190 2429 1196 2430
rect 1190 2425 1191 2429
rect 1195 2425 1196 2429
rect 1190 2424 1196 2425
rect 1366 2429 1372 2430
rect 1366 2425 1367 2429
rect 1371 2425 1372 2429
rect 1366 2424 1372 2425
rect 1534 2429 1540 2430
rect 1534 2425 1535 2429
rect 1539 2425 1540 2429
rect 1534 2424 1540 2425
rect 1702 2429 1708 2430
rect 1702 2425 1703 2429
rect 1707 2425 1708 2429
rect 1702 2424 1708 2425
rect 1870 2429 1876 2430
rect 1870 2425 1871 2429
rect 1875 2425 1876 2429
rect 2110 2426 2111 2430
rect 2115 2426 2116 2430
rect 1870 2424 1876 2425
rect 2070 2425 2076 2426
rect 2110 2425 2116 2426
rect 2310 2430 2316 2431
rect 2310 2426 2311 2430
rect 2315 2426 2316 2430
rect 2310 2425 2316 2426
rect 2534 2430 2540 2431
rect 2534 2426 2535 2430
rect 2539 2426 2540 2430
rect 2534 2425 2540 2426
rect 2750 2430 2756 2431
rect 2750 2426 2751 2430
rect 2755 2426 2756 2430
rect 2750 2425 2756 2426
rect 2950 2430 2956 2431
rect 2950 2426 2951 2430
rect 2955 2426 2956 2430
rect 2950 2425 2956 2426
rect 3134 2430 3140 2431
rect 3134 2426 3135 2430
rect 3139 2426 3140 2430
rect 3134 2425 3140 2426
rect 3310 2430 3316 2431
rect 3310 2426 3311 2430
rect 3315 2426 3316 2430
rect 3310 2425 3316 2426
rect 3470 2430 3476 2431
rect 3470 2426 3471 2430
rect 3475 2426 3476 2430
rect 3470 2425 3476 2426
rect 3622 2430 3628 2431
rect 3622 2426 3623 2430
rect 3627 2426 3628 2430
rect 3622 2425 3628 2426
rect 3766 2430 3772 2431
rect 3766 2426 3767 2430
rect 3771 2426 3772 2430
rect 3766 2425 3772 2426
rect 3894 2430 3900 2431
rect 3894 2426 3895 2430
rect 3899 2426 3900 2430
rect 3894 2425 3900 2426
rect 3990 2425 3996 2426
rect 2070 2421 2071 2425
rect 2075 2421 2076 2425
rect 2070 2420 2076 2421
rect 3990 2421 3991 2425
rect 3995 2421 3996 2425
rect 3990 2420 3996 2421
rect 2070 2408 2076 2409
rect 2070 2404 2071 2408
rect 2075 2404 2076 2408
rect 2070 2403 2076 2404
rect 3990 2408 3996 2409
rect 3990 2404 3991 2408
rect 3995 2404 3996 2408
rect 3990 2403 3996 2404
rect 2110 2389 2116 2390
rect 206 2387 212 2388
rect 206 2383 207 2387
rect 211 2383 212 2387
rect 206 2382 212 2383
rect 350 2387 356 2388
rect 350 2383 351 2387
rect 355 2383 356 2387
rect 350 2382 356 2383
rect 502 2387 508 2388
rect 502 2383 503 2387
rect 507 2383 508 2387
rect 502 2382 508 2383
rect 654 2387 660 2388
rect 654 2383 655 2387
rect 659 2383 660 2387
rect 654 2382 660 2383
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 966 2387 972 2388
rect 966 2383 967 2387
rect 971 2383 972 2387
rect 966 2382 972 2383
rect 1118 2387 1124 2388
rect 1118 2383 1119 2387
rect 1123 2383 1124 2387
rect 1118 2382 1124 2383
rect 1262 2387 1268 2388
rect 1262 2383 1263 2387
rect 1267 2383 1268 2387
rect 1262 2382 1268 2383
rect 1414 2387 1420 2388
rect 1414 2383 1415 2387
rect 1419 2383 1420 2387
rect 1414 2382 1420 2383
rect 1566 2387 1572 2388
rect 1566 2383 1567 2387
rect 1571 2383 1572 2387
rect 2110 2385 2111 2389
rect 2115 2385 2116 2389
rect 2110 2384 2116 2385
rect 2310 2389 2316 2390
rect 2310 2385 2311 2389
rect 2315 2385 2316 2389
rect 2310 2384 2316 2385
rect 2534 2389 2540 2390
rect 2534 2385 2535 2389
rect 2539 2385 2540 2389
rect 2534 2384 2540 2385
rect 2750 2389 2756 2390
rect 2750 2385 2751 2389
rect 2755 2385 2756 2389
rect 2750 2384 2756 2385
rect 2950 2389 2956 2390
rect 2950 2385 2951 2389
rect 2955 2385 2956 2389
rect 2950 2384 2956 2385
rect 3134 2389 3140 2390
rect 3134 2385 3135 2389
rect 3139 2385 3140 2389
rect 3134 2384 3140 2385
rect 3310 2389 3316 2390
rect 3310 2385 3311 2389
rect 3315 2385 3316 2389
rect 3310 2384 3316 2385
rect 3470 2389 3476 2390
rect 3470 2385 3471 2389
rect 3475 2385 3476 2389
rect 3470 2384 3476 2385
rect 3622 2389 3628 2390
rect 3622 2385 3623 2389
rect 3627 2385 3628 2389
rect 3622 2384 3628 2385
rect 3766 2389 3772 2390
rect 3766 2385 3767 2389
rect 3771 2385 3772 2389
rect 3766 2384 3772 2385
rect 3894 2389 3900 2390
rect 3894 2385 3895 2389
rect 3899 2385 3900 2389
rect 3894 2384 3900 2385
rect 1566 2382 1572 2383
rect 110 2368 116 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 2030 2368 2036 2369
rect 2030 2364 2031 2368
rect 2035 2364 2036 2368
rect 2030 2363 2036 2364
rect 2110 2359 2116 2360
rect 2110 2355 2111 2359
rect 2115 2355 2116 2359
rect 2110 2354 2116 2355
rect 2326 2359 2332 2360
rect 2326 2355 2327 2359
rect 2331 2355 2332 2359
rect 2326 2354 2332 2355
rect 2558 2359 2564 2360
rect 2558 2355 2559 2359
rect 2563 2355 2564 2359
rect 2558 2354 2564 2355
rect 2782 2359 2788 2360
rect 2782 2355 2783 2359
rect 2787 2355 2788 2359
rect 2782 2354 2788 2355
rect 2998 2359 3004 2360
rect 2998 2355 2999 2359
rect 3003 2355 3004 2359
rect 2998 2354 3004 2355
rect 3190 2359 3196 2360
rect 3190 2355 3191 2359
rect 3195 2355 3196 2359
rect 3190 2354 3196 2355
rect 3374 2359 3380 2360
rect 3374 2355 3375 2359
rect 3379 2355 3380 2359
rect 3374 2354 3380 2355
rect 3542 2359 3548 2360
rect 3542 2355 3543 2359
rect 3547 2355 3548 2359
rect 3542 2354 3548 2355
rect 3710 2359 3716 2360
rect 3710 2355 3711 2359
rect 3715 2355 3716 2359
rect 3710 2354 3716 2355
rect 3886 2359 3892 2360
rect 3886 2355 3887 2359
rect 3891 2355 3892 2359
rect 3886 2354 3892 2355
rect 110 2351 116 2352
rect 110 2347 111 2351
rect 115 2347 116 2351
rect 2030 2351 2036 2352
rect 2030 2347 2031 2351
rect 2035 2347 2036 2351
rect 110 2346 116 2347
rect 206 2346 212 2347
rect 206 2342 207 2346
rect 211 2342 212 2346
rect 206 2341 212 2342
rect 350 2346 356 2347
rect 350 2342 351 2346
rect 355 2342 356 2346
rect 350 2341 356 2342
rect 502 2346 508 2347
rect 502 2342 503 2346
rect 507 2342 508 2346
rect 502 2341 508 2342
rect 654 2346 660 2347
rect 654 2342 655 2346
rect 659 2342 660 2346
rect 654 2341 660 2342
rect 814 2346 820 2347
rect 814 2342 815 2346
rect 819 2342 820 2346
rect 814 2341 820 2342
rect 966 2346 972 2347
rect 966 2342 967 2346
rect 971 2342 972 2346
rect 966 2341 972 2342
rect 1118 2346 1124 2347
rect 1118 2342 1119 2346
rect 1123 2342 1124 2346
rect 1118 2341 1124 2342
rect 1262 2346 1268 2347
rect 1262 2342 1263 2346
rect 1267 2342 1268 2346
rect 1262 2341 1268 2342
rect 1414 2346 1420 2347
rect 1414 2342 1415 2346
rect 1419 2342 1420 2346
rect 1414 2341 1420 2342
rect 1566 2346 1572 2347
rect 2030 2346 2036 2347
rect 1566 2342 1567 2346
rect 1571 2342 1572 2346
rect 1566 2341 1572 2342
rect 2070 2340 2076 2341
rect 2070 2336 2071 2340
rect 2075 2336 2076 2340
rect 2070 2335 2076 2336
rect 3990 2340 3996 2341
rect 3990 2336 3991 2340
rect 3995 2336 3996 2340
rect 3990 2335 3996 2336
rect 2070 2323 2076 2324
rect 2070 2319 2071 2323
rect 2075 2319 2076 2323
rect 3990 2323 3996 2324
rect 3990 2319 3991 2323
rect 3995 2319 3996 2323
rect 2070 2318 2076 2319
rect 2110 2318 2116 2319
rect 2110 2314 2111 2318
rect 2115 2314 2116 2318
rect 2110 2313 2116 2314
rect 2326 2318 2332 2319
rect 2326 2314 2327 2318
rect 2331 2314 2332 2318
rect 2326 2313 2332 2314
rect 2558 2318 2564 2319
rect 2558 2314 2559 2318
rect 2563 2314 2564 2318
rect 2558 2313 2564 2314
rect 2782 2318 2788 2319
rect 2782 2314 2783 2318
rect 2787 2314 2788 2318
rect 2782 2313 2788 2314
rect 2998 2318 3004 2319
rect 2998 2314 2999 2318
rect 3003 2314 3004 2318
rect 2998 2313 3004 2314
rect 3190 2318 3196 2319
rect 3190 2314 3191 2318
rect 3195 2314 3196 2318
rect 3190 2313 3196 2314
rect 3374 2318 3380 2319
rect 3374 2314 3375 2318
rect 3379 2314 3380 2318
rect 3374 2313 3380 2314
rect 3542 2318 3548 2319
rect 3542 2314 3543 2318
rect 3547 2314 3548 2318
rect 3542 2313 3548 2314
rect 3710 2318 3716 2319
rect 3710 2314 3711 2318
rect 3715 2314 3716 2318
rect 3710 2313 3716 2314
rect 3886 2318 3892 2319
rect 3990 2318 3996 2319
rect 3886 2314 3887 2318
rect 3891 2314 3892 2318
rect 3886 2313 3892 2314
rect 254 2302 260 2303
rect 254 2298 255 2302
rect 259 2298 260 2302
rect 110 2297 116 2298
rect 254 2297 260 2298
rect 358 2302 364 2303
rect 358 2298 359 2302
rect 363 2298 364 2302
rect 358 2297 364 2298
rect 470 2302 476 2303
rect 470 2298 471 2302
rect 475 2298 476 2302
rect 470 2297 476 2298
rect 582 2302 588 2303
rect 582 2298 583 2302
rect 587 2298 588 2302
rect 582 2297 588 2298
rect 694 2302 700 2303
rect 694 2298 695 2302
rect 699 2298 700 2302
rect 694 2297 700 2298
rect 806 2302 812 2303
rect 806 2298 807 2302
rect 811 2298 812 2302
rect 806 2297 812 2298
rect 918 2302 924 2303
rect 918 2298 919 2302
rect 923 2298 924 2302
rect 918 2297 924 2298
rect 1030 2302 1036 2303
rect 1030 2298 1031 2302
rect 1035 2298 1036 2302
rect 1030 2297 1036 2298
rect 1150 2302 1156 2303
rect 1150 2298 1151 2302
rect 1155 2298 1156 2302
rect 1150 2297 1156 2298
rect 1270 2302 1276 2303
rect 1270 2298 1271 2302
rect 1275 2298 1276 2302
rect 1270 2297 1276 2298
rect 2030 2297 2036 2298
rect 110 2293 111 2297
rect 115 2293 116 2297
rect 110 2292 116 2293
rect 2030 2293 2031 2297
rect 2035 2293 2036 2297
rect 2030 2292 2036 2293
rect 2110 2286 2116 2287
rect 2110 2282 2111 2286
rect 2115 2282 2116 2286
rect 2070 2281 2076 2282
rect 2110 2281 2116 2282
rect 2294 2286 2300 2287
rect 2294 2282 2295 2286
rect 2299 2282 2300 2286
rect 2294 2281 2300 2282
rect 2526 2286 2532 2287
rect 2526 2282 2527 2286
rect 2531 2282 2532 2286
rect 2526 2281 2532 2282
rect 2774 2286 2780 2287
rect 2774 2282 2775 2286
rect 2779 2282 2780 2286
rect 2774 2281 2780 2282
rect 3038 2286 3044 2287
rect 3038 2282 3039 2286
rect 3043 2282 3044 2286
rect 3038 2281 3044 2282
rect 3318 2286 3324 2287
rect 3318 2282 3319 2286
rect 3323 2282 3324 2286
rect 3318 2281 3324 2282
rect 3606 2286 3612 2287
rect 3606 2282 3607 2286
rect 3611 2282 3612 2286
rect 3606 2281 3612 2282
rect 3894 2286 3900 2287
rect 3894 2282 3895 2286
rect 3899 2282 3900 2286
rect 3894 2281 3900 2282
rect 3990 2281 3996 2282
rect 110 2280 116 2281
rect 110 2276 111 2280
rect 115 2276 116 2280
rect 110 2275 116 2276
rect 2030 2280 2036 2281
rect 2030 2276 2031 2280
rect 2035 2276 2036 2280
rect 2070 2277 2071 2281
rect 2075 2277 2076 2281
rect 2070 2276 2076 2277
rect 3990 2277 3991 2281
rect 3995 2277 3996 2281
rect 3990 2276 3996 2277
rect 2030 2275 2036 2276
rect 2070 2264 2076 2265
rect 254 2261 260 2262
rect 254 2257 255 2261
rect 259 2257 260 2261
rect 254 2256 260 2257
rect 358 2261 364 2262
rect 358 2257 359 2261
rect 363 2257 364 2261
rect 358 2256 364 2257
rect 470 2261 476 2262
rect 470 2257 471 2261
rect 475 2257 476 2261
rect 470 2256 476 2257
rect 582 2261 588 2262
rect 582 2257 583 2261
rect 587 2257 588 2261
rect 582 2256 588 2257
rect 694 2261 700 2262
rect 694 2257 695 2261
rect 699 2257 700 2261
rect 694 2256 700 2257
rect 806 2261 812 2262
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 806 2256 812 2257
rect 918 2261 924 2262
rect 918 2257 919 2261
rect 923 2257 924 2261
rect 918 2256 924 2257
rect 1030 2261 1036 2262
rect 1030 2257 1031 2261
rect 1035 2257 1036 2261
rect 1030 2256 1036 2257
rect 1150 2261 1156 2262
rect 1150 2257 1151 2261
rect 1155 2257 1156 2261
rect 1150 2256 1156 2257
rect 1270 2261 1276 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 2070 2260 2071 2264
rect 2075 2260 2076 2264
rect 2070 2259 2076 2260
rect 3990 2264 3996 2265
rect 3990 2260 3991 2264
rect 3995 2260 3996 2264
rect 3990 2259 3996 2260
rect 1270 2256 1276 2257
rect 2110 2245 2116 2246
rect 2110 2241 2111 2245
rect 2115 2241 2116 2245
rect 2110 2240 2116 2241
rect 2294 2245 2300 2246
rect 2294 2241 2295 2245
rect 2299 2241 2300 2245
rect 2294 2240 2300 2241
rect 2526 2245 2532 2246
rect 2526 2241 2527 2245
rect 2531 2241 2532 2245
rect 2526 2240 2532 2241
rect 2774 2245 2780 2246
rect 2774 2241 2775 2245
rect 2779 2241 2780 2245
rect 2774 2240 2780 2241
rect 3038 2245 3044 2246
rect 3038 2241 3039 2245
rect 3043 2241 3044 2245
rect 3038 2240 3044 2241
rect 3318 2245 3324 2246
rect 3318 2241 3319 2245
rect 3323 2241 3324 2245
rect 3318 2240 3324 2241
rect 3606 2245 3612 2246
rect 3606 2241 3607 2245
rect 3611 2241 3612 2245
rect 3606 2240 3612 2241
rect 3894 2245 3900 2246
rect 3894 2241 3895 2245
rect 3899 2241 3900 2245
rect 3894 2240 3900 2241
rect 182 2219 188 2220
rect 182 2215 183 2219
rect 187 2215 188 2219
rect 182 2214 188 2215
rect 342 2219 348 2220
rect 342 2215 343 2219
rect 347 2215 348 2219
rect 342 2214 348 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 790 2219 796 2220
rect 790 2215 791 2219
rect 795 2215 796 2219
rect 790 2214 796 2215
rect 934 2219 940 2220
rect 934 2215 935 2219
rect 939 2215 940 2219
rect 934 2214 940 2215
rect 1070 2219 1076 2220
rect 1070 2215 1071 2219
rect 1075 2215 1076 2219
rect 1070 2214 1076 2215
rect 1198 2219 1204 2220
rect 1198 2215 1199 2219
rect 1203 2215 1204 2219
rect 1198 2214 1204 2215
rect 1334 2219 1340 2220
rect 1334 2215 1335 2219
rect 1339 2215 1340 2219
rect 1334 2214 1340 2215
rect 1470 2219 1476 2220
rect 1470 2215 1471 2219
rect 1475 2215 1476 2219
rect 1470 2214 1476 2215
rect 2278 2207 2284 2208
rect 2278 2203 2279 2207
rect 2283 2203 2284 2207
rect 2278 2202 2284 2203
rect 2438 2207 2444 2208
rect 2438 2203 2439 2207
rect 2443 2203 2444 2207
rect 2438 2202 2444 2203
rect 2622 2207 2628 2208
rect 2622 2203 2623 2207
rect 2627 2203 2628 2207
rect 2622 2202 2628 2203
rect 2838 2207 2844 2208
rect 2838 2203 2839 2207
rect 2843 2203 2844 2207
rect 2838 2202 2844 2203
rect 3078 2207 3084 2208
rect 3078 2203 3079 2207
rect 3083 2203 3084 2207
rect 3078 2202 3084 2203
rect 3342 2207 3348 2208
rect 3342 2203 3343 2207
rect 3347 2203 3348 2207
rect 3342 2202 3348 2203
rect 3622 2207 3628 2208
rect 3622 2203 3623 2207
rect 3627 2203 3628 2207
rect 3622 2202 3628 2203
rect 3894 2207 3900 2208
rect 3894 2203 3895 2207
rect 3899 2203 3900 2207
rect 3894 2202 3900 2203
rect 110 2200 116 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 2030 2200 2036 2201
rect 2030 2196 2031 2200
rect 2035 2196 2036 2200
rect 2030 2195 2036 2196
rect 2070 2188 2076 2189
rect 2070 2184 2071 2188
rect 2075 2184 2076 2188
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 2030 2183 2036 2184
rect 2070 2183 2076 2184
rect 3990 2188 3996 2189
rect 3990 2184 3991 2188
rect 3995 2184 3996 2188
rect 3990 2183 3996 2184
rect 2030 2179 2031 2183
rect 2035 2179 2036 2183
rect 110 2178 116 2179
rect 182 2178 188 2179
rect 182 2174 183 2178
rect 187 2174 188 2178
rect 182 2173 188 2174
rect 342 2178 348 2179
rect 342 2174 343 2178
rect 347 2174 348 2178
rect 342 2173 348 2174
rect 494 2178 500 2179
rect 494 2174 495 2178
rect 499 2174 500 2178
rect 494 2173 500 2174
rect 646 2178 652 2179
rect 646 2174 647 2178
rect 651 2174 652 2178
rect 646 2173 652 2174
rect 790 2178 796 2179
rect 790 2174 791 2178
rect 795 2174 796 2178
rect 790 2173 796 2174
rect 934 2178 940 2179
rect 934 2174 935 2178
rect 939 2174 940 2178
rect 934 2173 940 2174
rect 1070 2178 1076 2179
rect 1070 2174 1071 2178
rect 1075 2174 1076 2178
rect 1070 2173 1076 2174
rect 1198 2178 1204 2179
rect 1198 2174 1199 2178
rect 1203 2174 1204 2178
rect 1198 2173 1204 2174
rect 1334 2178 1340 2179
rect 1334 2174 1335 2178
rect 1339 2174 1340 2178
rect 1334 2173 1340 2174
rect 1470 2178 1476 2179
rect 2030 2178 2036 2179
rect 1470 2174 1471 2178
rect 1475 2174 1476 2178
rect 1470 2173 1476 2174
rect 2070 2171 2076 2172
rect 2070 2167 2071 2171
rect 2075 2167 2076 2171
rect 3990 2171 3996 2172
rect 3990 2167 3991 2171
rect 3995 2167 3996 2171
rect 2070 2166 2076 2167
rect 2278 2166 2284 2167
rect 2278 2162 2279 2166
rect 2283 2162 2284 2166
rect 2278 2161 2284 2162
rect 2438 2166 2444 2167
rect 2438 2162 2439 2166
rect 2443 2162 2444 2166
rect 2438 2161 2444 2162
rect 2622 2166 2628 2167
rect 2622 2162 2623 2166
rect 2627 2162 2628 2166
rect 2622 2161 2628 2162
rect 2838 2166 2844 2167
rect 2838 2162 2839 2166
rect 2843 2162 2844 2166
rect 2838 2161 2844 2162
rect 3078 2166 3084 2167
rect 3078 2162 3079 2166
rect 3083 2162 3084 2166
rect 3078 2161 3084 2162
rect 3342 2166 3348 2167
rect 3342 2162 3343 2166
rect 3347 2162 3348 2166
rect 3342 2161 3348 2162
rect 3622 2166 3628 2167
rect 3622 2162 3623 2166
rect 3627 2162 3628 2166
rect 3622 2161 3628 2162
rect 3894 2166 3900 2167
rect 3990 2166 3996 2167
rect 3894 2162 3895 2166
rect 3899 2162 3900 2166
rect 3894 2161 3900 2162
rect 2390 2134 2396 2135
rect 150 2130 156 2131
rect 150 2126 151 2130
rect 155 2126 156 2130
rect 110 2125 116 2126
rect 150 2125 156 2126
rect 326 2130 332 2131
rect 326 2126 327 2130
rect 331 2126 332 2130
rect 326 2125 332 2126
rect 534 2130 540 2131
rect 534 2126 535 2130
rect 539 2126 540 2130
rect 534 2125 540 2126
rect 734 2130 740 2131
rect 734 2126 735 2130
rect 739 2126 740 2130
rect 734 2125 740 2126
rect 926 2130 932 2131
rect 926 2126 927 2130
rect 931 2126 932 2130
rect 926 2125 932 2126
rect 1110 2130 1116 2131
rect 1110 2126 1111 2130
rect 1115 2126 1116 2130
rect 1110 2125 1116 2126
rect 1278 2130 1284 2131
rect 1278 2126 1279 2130
rect 1283 2126 1284 2130
rect 1278 2125 1284 2126
rect 1446 2130 1452 2131
rect 1446 2126 1447 2130
rect 1451 2126 1452 2130
rect 1446 2125 1452 2126
rect 1614 2130 1620 2131
rect 1614 2126 1615 2130
rect 1619 2126 1620 2130
rect 1614 2125 1620 2126
rect 1782 2130 1788 2131
rect 2390 2130 2391 2134
rect 2395 2130 2396 2134
rect 1782 2126 1783 2130
rect 1787 2126 1788 2130
rect 2070 2129 2076 2130
rect 2390 2129 2396 2130
rect 2494 2134 2500 2135
rect 2494 2130 2495 2134
rect 2499 2130 2500 2134
rect 2494 2129 2500 2130
rect 2598 2134 2604 2135
rect 2598 2130 2599 2134
rect 2603 2130 2604 2134
rect 2598 2129 2604 2130
rect 2702 2134 2708 2135
rect 2702 2130 2703 2134
rect 2707 2130 2708 2134
rect 2702 2129 2708 2130
rect 2806 2134 2812 2135
rect 2806 2130 2807 2134
rect 2811 2130 2812 2134
rect 2806 2129 2812 2130
rect 2910 2134 2916 2135
rect 2910 2130 2911 2134
rect 2915 2130 2916 2134
rect 2910 2129 2916 2130
rect 3030 2134 3036 2135
rect 3030 2130 3031 2134
rect 3035 2130 3036 2134
rect 3030 2129 3036 2130
rect 3174 2134 3180 2135
rect 3174 2130 3175 2134
rect 3179 2130 3180 2134
rect 3174 2129 3180 2130
rect 3342 2134 3348 2135
rect 3342 2130 3343 2134
rect 3347 2130 3348 2134
rect 3342 2129 3348 2130
rect 3526 2134 3532 2135
rect 3526 2130 3527 2134
rect 3531 2130 3532 2134
rect 3526 2129 3532 2130
rect 3718 2134 3724 2135
rect 3718 2130 3719 2134
rect 3723 2130 3724 2134
rect 3718 2129 3724 2130
rect 3894 2134 3900 2135
rect 3894 2130 3895 2134
rect 3899 2130 3900 2134
rect 3894 2129 3900 2130
rect 3990 2129 3996 2130
rect 1782 2125 1788 2126
rect 2030 2125 2036 2126
rect 110 2121 111 2125
rect 115 2121 116 2125
rect 110 2120 116 2121
rect 2030 2121 2031 2125
rect 2035 2121 2036 2125
rect 2070 2125 2071 2129
rect 2075 2125 2076 2129
rect 2070 2124 2076 2125
rect 3990 2125 3991 2129
rect 3995 2125 3996 2129
rect 3990 2124 3996 2125
rect 2030 2120 2036 2121
rect 2070 2112 2076 2113
rect 110 2108 116 2109
rect 110 2104 111 2108
rect 115 2104 116 2108
rect 110 2103 116 2104
rect 2030 2108 2036 2109
rect 2030 2104 2031 2108
rect 2035 2104 2036 2108
rect 2070 2108 2071 2112
rect 2075 2108 2076 2112
rect 2070 2107 2076 2108
rect 3990 2112 3996 2113
rect 3990 2108 3991 2112
rect 3995 2108 3996 2112
rect 3990 2107 3996 2108
rect 2030 2103 2036 2104
rect 2390 2093 2396 2094
rect 150 2089 156 2090
rect 150 2085 151 2089
rect 155 2085 156 2089
rect 150 2084 156 2085
rect 326 2089 332 2090
rect 326 2085 327 2089
rect 331 2085 332 2089
rect 326 2084 332 2085
rect 534 2089 540 2090
rect 534 2085 535 2089
rect 539 2085 540 2089
rect 534 2084 540 2085
rect 734 2089 740 2090
rect 734 2085 735 2089
rect 739 2085 740 2089
rect 734 2084 740 2085
rect 926 2089 932 2090
rect 926 2085 927 2089
rect 931 2085 932 2089
rect 926 2084 932 2085
rect 1110 2089 1116 2090
rect 1110 2085 1111 2089
rect 1115 2085 1116 2089
rect 1110 2084 1116 2085
rect 1278 2089 1284 2090
rect 1278 2085 1279 2089
rect 1283 2085 1284 2089
rect 1278 2084 1284 2085
rect 1446 2089 1452 2090
rect 1446 2085 1447 2089
rect 1451 2085 1452 2089
rect 1446 2084 1452 2085
rect 1614 2089 1620 2090
rect 1614 2085 1615 2089
rect 1619 2085 1620 2089
rect 1614 2084 1620 2085
rect 1782 2089 1788 2090
rect 1782 2085 1783 2089
rect 1787 2085 1788 2089
rect 2390 2089 2391 2093
rect 2395 2089 2396 2093
rect 2390 2088 2396 2089
rect 2494 2093 2500 2094
rect 2494 2089 2495 2093
rect 2499 2089 2500 2093
rect 2494 2088 2500 2089
rect 2598 2093 2604 2094
rect 2598 2089 2599 2093
rect 2603 2089 2604 2093
rect 2598 2088 2604 2089
rect 2702 2093 2708 2094
rect 2702 2089 2703 2093
rect 2707 2089 2708 2093
rect 2702 2088 2708 2089
rect 2806 2093 2812 2094
rect 2806 2089 2807 2093
rect 2811 2089 2812 2093
rect 2806 2088 2812 2089
rect 2910 2093 2916 2094
rect 2910 2089 2911 2093
rect 2915 2089 2916 2093
rect 2910 2088 2916 2089
rect 3030 2093 3036 2094
rect 3030 2089 3031 2093
rect 3035 2089 3036 2093
rect 3030 2088 3036 2089
rect 3174 2093 3180 2094
rect 3174 2089 3175 2093
rect 3179 2089 3180 2093
rect 3174 2088 3180 2089
rect 3342 2093 3348 2094
rect 3342 2089 3343 2093
rect 3347 2089 3348 2093
rect 3342 2088 3348 2089
rect 3526 2093 3532 2094
rect 3526 2089 3527 2093
rect 3531 2089 3532 2093
rect 3526 2088 3532 2089
rect 3718 2093 3724 2094
rect 3718 2089 3719 2093
rect 3723 2089 3724 2093
rect 3718 2088 3724 2089
rect 3894 2093 3900 2094
rect 3894 2089 3895 2093
rect 3899 2089 3900 2093
rect 3894 2088 3900 2089
rect 1782 2084 1788 2085
rect 2486 2059 2492 2060
rect 2486 2055 2487 2059
rect 2491 2055 2492 2059
rect 2486 2054 2492 2055
rect 2590 2059 2596 2060
rect 2590 2055 2591 2059
rect 2595 2055 2596 2059
rect 2590 2054 2596 2055
rect 2694 2059 2700 2060
rect 2694 2055 2695 2059
rect 2699 2055 2700 2059
rect 2694 2054 2700 2055
rect 2806 2059 2812 2060
rect 2806 2055 2807 2059
rect 2811 2055 2812 2059
rect 2806 2054 2812 2055
rect 2934 2059 2940 2060
rect 2934 2055 2935 2059
rect 2939 2055 2940 2059
rect 2934 2054 2940 2055
rect 3094 2059 3100 2060
rect 3094 2055 3095 2059
rect 3099 2055 3100 2059
rect 3094 2054 3100 2055
rect 3278 2059 3284 2060
rect 3278 2055 3279 2059
rect 3283 2055 3284 2059
rect 3278 2054 3284 2055
rect 3478 2059 3484 2060
rect 3478 2055 3479 2059
rect 3483 2055 3484 2059
rect 3478 2054 3484 2055
rect 3694 2059 3700 2060
rect 3694 2055 3695 2059
rect 3699 2055 3700 2059
rect 3694 2054 3700 2055
rect 3894 2059 3900 2060
rect 3894 2055 3895 2059
rect 3899 2055 3900 2059
rect 3894 2054 3900 2055
rect 150 2047 156 2048
rect 150 2043 151 2047
rect 155 2043 156 2047
rect 150 2042 156 2043
rect 382 2047 388 2048
rect 382 2043 383 2047
rect 387 2043 388 2047
rect 382 2042 388 2043
rect 630 2047 636 2048
rect 630 2043 631 2047
rect 635 2043 636 2047
rect 630 2042 636 2043
rect 862 2047 868 2048
rect 862 2043 863 2047
rect 867 2043 868 2047
rect 862 2042 868 2043
rect 1070 2047 1076 2048
rect 1070 2043 1071 2047
rect 1075 2043 1076 2047
rect 1070 2042 1076 2043
rect 1262 2047 1268 2048
rect 1262 2043 1263 2047
rect 1267 2043 1268 2047
rect 1262 2042 1268 2043
rect 1446 2047 1452 2048
rect 1446 2043 1447 2047
rect 1451 2043 1452 2047
rect 1446 2042 1452 2043
rect 1614 2047 1620 2048
rect 1614 2043 1615 2047
rect 1619 2043 1620 2047
rect 1614 2042 1620 2043
rect 1782 2047 1788 2048
rect 1782 2043 1783 2047
rect 1787 2043 1788 2047
rect 1782 2042 1788 2043
rect 1934 2047 1940 2048
rect 1934 2043 1935 2047
rect 1939 2043 1940 2047
rect 1934 2042 1940 2043
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 3990 2040 3996 2041
rect 3990 2036 3991 2040
rect 3995 2036 3996 2040
rect 3990 2035 3996 2036
rect 110 2028 116 2029
rect 110 2024 111 2028
rect 115 2024 116 2028
rect 110 2023 116 2024
rect 2030 2028 2036 2029
rect 2030 2024 2031 2028
rect 2035 2024 2036 2028
rect 2030 2023 2036 2024
rect 2070 2023 2076 2024
rect 2070 2019 2071 2023
rect 2075 2019 2076 2023
rect 3990 2023 3996 2024
rect 3990 2019 3991 2023
rect 3995 2019 3996 2023
rect 2070 2018 2076 2019
rect 2486 2018 2492 2019
rect 2486 2014 2487 2018
rect 2491 2014 2492 2018
rect 2486 2013 2492 2014
rect 2590 2018 2596 2019
rect 2590 2014 2591 2018
rect 2595 2014 2596 2018
rect 2590 2013 2596 2014
rect 2694 2018 2700 2019
rect 2694 2014 2695 2018
rect 2699 2014 2700 2018
rect 2694 2013 2700 2014
rect 2806 2018 2812 2019
rect 2806 2014 2807 2018
rect 2811 2014 2812 2018
rect 2806 2013 2812 2014
rect 2934 2018 2940 2019
rect 2934 2014 2935 2018
rect 2939 2014 2940 2018
rect 2934 2013 2940 2014
rect 3094 2018 3100 2019
rect 3094 2014 3095 2018
rect 3099 2014 3100 2018
rect 3094 2013 3100 2014
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3478 2018 3484 2019
rect 3478 2014 3479 2018
rect 3483 2014 3484 2018
rect 3478 2013 3484 2014
rect 3694 2018 3700 2019
rect 3694 2014 3695 2018
rect 3699 2014 3700 2018
rect 3694 2013 3700 2014
rect 3894 2018 3900 2019
rect 3990 2018 3996 2019
rect 3894 2014 3895 2018
rect 3899 2014 3900 2018
rect 3894 2013 3900 2014
rect 110 2011 116 2012
rect 110 2007 111 2011
rect 115 2007 116 2011
rect 2030 2011 2036 2012
rect 2030 2007 2031 2011
rect 2035 2007 2036 2011
rect 110 2006 116 2007
rect 150 2006 156 2007
rect 150 2002 151 2006
rect 155 2002 156 2006
rect 150 2001 156 2002
rect 382 2006 388 2007
rect 382 2002 383 2006
rect 387 2002 388 2006
rect 382 2001 388 2002
rect 630 2006 636 2007
rect 630 2002 631 2006
rect 635 2002 636 2006
rect 630 2001 636 2002
rect 862 2006 868 2007
rect 862 2002 863 2006
rect 867 2002 868 2006
rect 862 2001 868 2002
rect 1070 2006 1076 2007
rect 1070 2002 1071 2006
rect 1075 2002 1076 2006
rect 1070 2001 1076 2002
rect 1262 2006 1268 2007
rect 1262 2002 1263 2006
rect 1267 2002 1268 2006
rect 1262 2001 1268 2002
rect 1446 2006 1452 2007
rect 1446 2002 1447 2006
rect 1451 2002 1452 2006
rect 1446 2001 1452 2002
rect 1614 2006 1620 2007
rect 1614 2002 1615 2006
rect 1619 2002 1620 2006
rect 1614 2001 1620 2002
rect 1782 2006 1788 2007
rect 1782 2002 1783 2006
rect 1787 2002 1788 2006
rect 1782 2001 1788 2002
rect 1934 2006 1940 2007
rect 2030 2006 2036 2007
rect 1934 2002 1935 2006
rect 1939 2002 1940 2006
rect 1934 2001 1940 2002
rect 2526 1978 2532 1979
rect 2526 1974 2527 1978
rect 2531 1974 2532 1978
rect 2070 1973 2076 1974
rect 2526 1973 2532 1974
rect 2702 1978 2708 1979
rect 2702 1974 2703 1978
rect 2707 1974 2708 1978
rect 2702 1973 2708 1974
rect 2886 1978 2892 1979
rect 2886 1974 2887 1978
rect 2891 1974 2892 1978
rect 2886 1973 2892 1974
rect 3078 1978 3084 1979
rect 3078 1974 3079 1978
rect 3083 1974 3084 1978
rect 3078 1973 3084 1974
rect 3278 1978 3284 1979
rect 3278 1974 3279 1978
rect 3283 1974 3284 1978
rect 3278 1973 3284 1974
rect 3486 1978 3492 1979
rect 3486 1974 3487 1978
rect 3491 1974 3492 1978
rect 3486 1973 3492 1974
rect 3702 1978 3708 1979
rect 3702 1974 3703 1978
rect 3707 1974 3708 1978
rect 3702 1973 3708 1974
rect 3894 1978 3900 1979
rect 3894 1974 3895 1978
rect 3899 1974 3900 1978
rect 3894 1973 3900 1974
rect 3990 1973 3996 1974
rect 2070 1969 2071 1973
rect 2075 1969 2076 1973
rect 2070 1968 2076 1969
rect 3990 1969 3991 1973
rect 3995 1969 3996 1973
rect 3990 1968 3996 1969
rect 150 1962 156 1963
rect 150 1958 151 1962
rect 155 1958 156 1962
rect 110 1957 116 1958
rect 150 1957 156 1958
rect 326 1962 332 1963
rect 326 1958 327 1962
rect 331 1958 332 1962
rect 326 1957 332 1958
rect 534 1962 540 1963
rect 534 1958 535 1962
rect 539 1958 540 1962
rect 534 1957 540 1958
rect 734 1962 740 1963
rect 734 1958 735 1962
rect 739 1958 740 1962
rect 734 1957 740 1958
rect 934 1962 940 1963
rect 934 1958 935 1962
rect 939 1958 940 1962
rect 934 1957 940 1958
rect 1126 1962 1132 1963
rect 1126 1958 1127 1962
rect 1131 1958 1132 1962
rect 1126 1957 1132 1958
rect 1302 1962 1308 1963
rect 1302 1958 1303 1962
rect 1307 1958 1308 1962
rect 1302 1957 1308 1958
rect 1470 1962 1476 1963
rect 1470 1958 1471 1962
rect 1475 1958 1476 1962
rect 1470 1957 1476 1958
rect 1630 1962 1636 1963
rect 1630 1958 1631 1962
rect 1635 1958 1636 1962
rect 1630 1957 1636 1958
rect 1790 1962 1796 1963
rect 1790 1958 1791 1962
rect 1795 1958 1796 1962
rect 1790 1957 1796 1958
rect 1934 1962 1940 1963
rect 1934 1958 1935 1962
rect 1939 1958 1940 1962
rect 1934 1957 1940 1958
rect 2030 1957 2036 1958
rect 110 1953 111 1957
rect 115 1953 116 1957
rect 110 1952 116 1953
rect 2030 1953 2031 1957
rect 2035 1953 2036 1957
rect 2030 1952 2036 1953
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2070 1951 2076 1952
rect 3990 1956 3996 1957
rect 3990 1952 3991 1956
rect 3995 1952 3996 1956
rect 3990 1951 3996 1952
rect 110 1940 116 1941
rect 110 1936 111 1940
rect 115 1936 116 1940
rect 110 1935 116 1936
rect 2030 1940 2036 1941
rect 2030 1936 2031 1940
rect 2035 1936 2036 1940
rect 2030 1935 2036 1936
rect 2526 1937 2532 1938
rect 2526 1933 2527 1937
rect 2531 1933 2532 1937
rect 2526 1932 2532 1933
rect 2702 1937 2708 1938
rect 2702 1933 2703 1937
rect 2707 1933 2708 1937
rect 2702 1932 2708 1933
rect 2886 1937 2892 1938
rect 2886 1933 2887 1937
rect 2891 1933 2892 1937
rect 2886 1932 2892 1933
rect 3078 1937 3084 1938
rect 3078 1933 3079 1937
rect 3083 1933 3084 1937
rect 3078 1932 3084 1933
rect 3278 1937 3284 1938
rect 3278 1933 3279 1937
rect 3283 1933 3284 1937
rect 3278 1932 3284 1933
rect 3486 1937 3492 1938
rect 3486 1933 3487 1937
rect 3491 1933 3492 1937
rect 3486 1932 3492 1933
rect 3702 1937 3708 1938
rect 3702 1933 3703 1937
rect 3707 1933 3708 1937
rect 3702 1932 3708 1933
rect 3894 1937 3900 1938
rect 3894 1933 3895 1937
rect 3899 1933 3900 1937
rect 3894 1932 3900 1933
rect 150 1921 156 1922
rect 150 1917 151 1921
rect 155 1917 156 1921
rect 150 1916 156 1917
rect 326 1921 332 1922
rect 326 1917 327 1921
rect 331 1917 332 1921
rect 326 1916 332 1917
rect 534 1921 540 1922
rect 534 1917 535 1921
rect 539 1917 540 1921
rect 534 1916 540 1917
rect 734 1921 740 1922
rect 734 1917 735 1921
rect 739 1917 740 1921
rect 734 1916 740 1917
rect 934 1921 940 1922
rect 934 1917 935 1921
rect 939 1917 940 1921
rect 934 1916 940 1917
rect 1126 1921 1132 1922
rect 1126 1917 1127 1921
rect 1131 1917 1132 1921
rect 1126 1916 1132 1917
rect 1302 1921 1308 1922
rect 1302 1917 1303 1921
rect 1307 1917 1308 1921
rect 1302 1916 1308 1917
rect 1470 1921 1476 1922
rect 1470 1917 1471 1921
rect 1475 1917 1476 1921
rect 1470 1916 1476 1917
rect 1630 1921 1636 1922
rect 1630 1917 1631 1921
rect 1635 1917 1636 1921
rect 1630 1916 1636 1917
rect 1790 1921 1796 1922
rect 1790 1917 1791 1921
rect 1795 1917 1796 1921
rect 1790 1916 1796 1917
rect 1934 1921 1940 1922
rect 1934 1917 1935 1921
rect 1939 1917 1940 1921
rect 1934 1916 1940 1917
rect 2110 1903 2116 1904
rect 2110 1899 2111 1903
rect 2115 1899 2116 1903
rect 2110 1898 2116 1899
rect 2302 1903 2308 1904
rect 2302 1899 2303 1903
rect 2307 1899 2308 1903
rect 2302 1898 2308 1899
rect 2518 1903 2524 1904
rect 2518 1899 2519 1903
rect 2523 1899 2524 1903
rect 2518 1898 2524 1899
rect 2734 1903 2740 1904
rect 2734 1899 2735 1903
rect 2739 1899 2740 1903
rect 2734 1898 2740 1899
rect 2958 1903 2964 1904
rect 2958 1899 2959 1903
rect 2963 1899 2964 1903
rect 2958 1898 2964 1899
rect 3190 1903 3196 1904
rect 3190 1899 3191 1903
rect 3195 1899 3196 1903
rect 3190 1898 3196 1899
rect 3430 1903 3436 1904
rect 3430 1899 3431 1903
rect 3435 1899 3436 1903
rect 3430 1898 3436 1899
rect 3670 1903 3676 1904
rect 3670 1899 3671 1903
rect 3675 1899 3676 1903
rect 3670 1898 3676 1899
rect 3894 1903 3900 1904
rect 3894 1899 3895 1903
rect 3899 1899 3900 1903
rect 3894 1898 3900 1899
rect 150 1887 156 1888
rect 150 1883 151 1887
rect 155 1883 156 1887
rect 150 1882 156 1883
rect 302 1887 308 1888
rect 302 1883 303 1887
rect 307 1883 308 1887
rect 302 1882 308 1883
rect 462 1887 468 1888
rect 462 1883 463 1887
rect 467 1883 468 1887
rect 462 1882 468 1883
rect 614 1887 620 1888
rect 614 1883 615 1887
rect 619 1883 620 1887
rect 614 1882 620 1883
rect 766 1887 772 1888
rect 766 1883 767 1887
rect 771 1883 772 1887
rect 766 1882 772 1883
rect 926 1887 932 1888
rect 926 1883 927 1887
rect 931 1883 932 1887
rect 926 1882 932 1883
rect 1102 1887 1108 1888
rect 1102 1883 1103 1887
rect 1107 1883 1108 1887
rect 1102 1882 1108 1883
rect 1294 1887 1300 1888
rect 1294 1883 1295 1887
rect 1299 1883 1300 1887
rect 1294 1882 1300 1883
rect 1510 1887 1516 1888
rect 1510 1883 1511 1887
rect 1515 1883 1516 1887
rect 1510 1882 1516 1883
rect 1734 1887 1740 1888
rect 1734 1883 1735 1887
rect 1739 1883 1740 1887
rect 1734 1882 1740 1883
rect 1934 1887 1940 1888
rect 1934 1883 1935 1887
rect 1939 1883 1940 1887
rect 1934 1882 1940 1883
rect 2070 1884 2076 1885
rect 2070 1880 2071 1884
rect 2075 1880 2076 1884
rect 2070 1879 2076 1880
rect 3990 1884 3996 1885
rect 3990 1880 3991 1884
rect 3995 1880 3996 1884
rect 3990 1879 3996 1880
rect 110 1868 116 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2070 1867 2076 1868
rect 2070 1863 2071 1867
rect 2075 1863 2076 1867
rect 3990 1867 3996 1868
rect 3990 1863 3991 1867
rect 3995 1863 3996 1867
rect 2070 1862 2076 1863
rect 2110 1862 2116 1863
rect 2110 1858 2111 1862
rect 2115 1858 2116 1862
rect 2110 1857 2116 1858
rect 2302 1862 2308 1863
rect 2302 1858 2303 1862
rect 2307 1858 2308 1862
rect 2302 1857 2308 1858
rect 2518 1862 2524 1863
rect 2518 1858 2519 1862
rect 2523 1858 2524 1862
rect 2518 1857 2524 1858
rect 2734 1862 2740 1863
rect 2734 1858 2735 1862
rect 2739 1858 2740 1862
rect 2734 1857 2740 1858
rect 2958 1862 2964 1863
rect 2958 1858 2959 1862
rect 2963 1858 2964 1862
rect 2958 1857 2964 1858
rect 3190 1862 3196 1863
rect 3190 1858 3191 1862
rect 3195 1858 3196 1862
rect 3190 1857 3196 1858
rect 3430 1862 3436 1863
rect 3430 1858 3431 1862
rect 3435 1858 3436 1862
rect 3430 1857 3436 1858
rect 3670 1862 3676 1863
rect 3670 1858 3671 1862
rect 3675 1858 3676 1862
rect 3670 1857 3676 1858
rect 3894 1862 3900 1863
rect 3990 1862 3996 1863
rect 3894 1858 3895 1862
rect 3899 1858 3900 1862
rect 3894 1857 3900 1858
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 2030 1851 2036 1852
rect 2030 1847 2031 1851
rect 2035 1847 2036 1851
rect 110 1846 116 1847
rect 150 1846 156 1847
rect 150 1842 151 1846
rect 155 1842 156 1846
rect 150 1841 156 1842
rect 302 1846 308 1847
rect 302 1842 303 1846
rect 307 1842 308 1846
rect 302 1841 308 1842
rect 462 1846 468 1847
rect 462 1842 463 1846
rect 467 1842 468 1846
rect 462 1841 468 1842
rect 614 1846 620 1847
rect 614 1842 615 1846
rect 619 1842 620 1846
rect 614 1841 620 1842
rect 766 1846 772 1847
rect 766 1842 767 1846
rect 771 1842 772 1846
rect 766 1841 772 1842
rect 926 1846 932 1847
rect 926 1842 927 1846
rect 931 1842 932 1846
rect 926 1841 932 1842
rect 1102 1846 1108 1847
rect 1102 1842 1103 1846
rect 1107 1842 1108 1846
rect 1102 1841 1108 1842
rect 1294 1846 1300 1847
rect 1294 1842 1295 1846
rect 1299 1842 1300 1846
rect 1294 1841 1300 1842
rect 1510 1846 1516 1847
rect 1510 1842 1511 1846
rect 1515 1842 1516 1846
rect 1510 1841 1516 1842
rect 1734 1846 1740 1847
rect 1734 1842 1735 1846
rect 1739 1842 1740 1846
rect 1734 1841 1740 1842
rect 1934 1846 1940 1847
rect 2030 1846 2036 1847
rect 1934 1842 1935 1846
rect 1939 1842 1940 1846
rect 1934 1841 1940 1842
rect 2110 1830 2116 1831
rect 2110 1826 2111 1830
rect 2115 1826 2116 1830
rect 2070 1825 2076 1826
rect 2110 1825 2116 1826
rect 2230 1830 2236 1831
rect 2230 1826 2231 1830
rect 2235 1826 2236 1830
rect 2230 1825 2236 1826
rect 2398 1830 2404 1831
rect 2398 1826 2399 1830
rect 2403 1826 2404 1830
rect 2398 1825 2404 1826
rect 2598 1830 2604 1831
rect 2598 1826 2599 1830
rect 2603 1826 2604 1830
rect 2598 1825 2604 1826
rect 2830 1830 2836 1831
rect 2830 1826 2831 1830
rect 2835 1826 2836 1830
rect 2830 1825 2836 1826
rect 3078 1830 3084 1831
rect 3078 1826 3079 1830
rect 3083 1826 3084 1830
rect 3078 1825 3084 1826
rect 3350 1830 3356 1831
rect 3350 1826 3351 1830
rect 3355 1826 3356 1830
rect 3350 1825 3356 1826
rect 3630 1830 3636 1831
rect 3630 1826 3631 1830
rect 3635 1826 3636 1830
rect 3630 1825 3636 1826
rect 3894 1830 3900 1831
rect 3894 1826 3895 1830
rect 3899 1826 3900 1830
rect 3894 1825 3900 1826
rect 3990 1825 3996 1826
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 3990 1821 3991 1825
rect 3995 1821 3996 1825
rect 3990 1820 3996 1821
rect 2070 1808 2076 1809
rect 2070 1804 2071 1808
rect 2075 1804 2076 1808
rect 2070 1803 2076 1804
rect 3990 1808 3996 1809
rect 3990 1804 3991 1808
rect 3995 1804 3996 1808
rect 3990 1803 3996 1804
rect 150 1802 156 1803
rect 150 1798 151 1802
rect 155 1798 156 1802
rect 110 1797 116 1798
rect 150 1797 156 1798
rect 342 1802 348 1803
rect 342 1798 343 1802
rect 347 1798 348 1802
rect 342 1797 348 1798
rect 542 1802 548 1803
rect 542 1798 543 1802
rect 547 1798 548 1802
rect 542 1797 548 1798
rect 734 1802 740 1803
rect 734 1798 735 1802
rect 739 1798 740 1802
rect 734 1797 740 1798
rect 918 1802 924 1803
rect 918 1798 919 1802
rect 923 1798 924 1802
rect 918 1797 924 1798
rect 1094 1802 1100 1803
rect 1094 1798 1095 1802
rect 1099 1798 1100 1802
rect 1094 1797 1100 1798
rect 1270 1802 1276 1803
rect 1270 1798 1271 1802
rect 1275 1798 1276 1802
rect 1270 1797 1276 1798
rect 1446 1802 1452 1803
rect 1446 1798 1447 1802
rect 1451 1798 1452 1802
rect 1446 1797 1452 1798
rect 1622 1802 1628 1803
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1806 1802 1812 1803
rect 1806 1798 1807 1802
rect 1811 1798 1812 1802
rect 1806 1797 1812 1798
rect 2030 1797 2036 1798
rect 110 1793 111 1797
rect 115 1793 116 1797
rect 110 1792 116 1793
rect 2030 1793 2031 1797
rect 2035 1793 2036 1797
rect 2030 1792 2036 1793
rect 2110 1789 2116 1790
rect 2110 1785 2111 1789
rect 2115 1785 2116 1789
rect 2110 1784 2116 1785
rect 2230 1789 2236 1790
rect 2230 1785 2231 1789
rect 2235 1785 2236 1789
rect 2230 1784 2236 1785
rect 2398 1789 2404 1790
rect 2398 1785 2399 1789
rect 2403 1785 2404 1789
rect 2398 1784 2404 1785
rect 2598 1789 2604 1790
rect 2598 1785 2599 1789
rect 2603 1785 2604 1789
rect 2598 1784 2604 1785
rect 2830 1789 2836 1790
rect 2830 1785 2831 1789
rect 2835 1785 2836 1789
rect 2830 1784 2836 1785
rect 3078 1789 3084 1790
rect 3078 1785 3079 1789
rect 3083 1785 3084 1789
rect 3078 1784 3084 1785
rect 3350 1789 3356 1790
rect 3350 1785 3351 1789
rect 3355 1785 3356 1789
rect 3350 1784 3356 1785
rect 3630 1789 3636 1790
rect 3630 1785 3631 1789
rect 3635 1785 3636 1789
rect 3630 1784 3636 1785
rect 3894 1789 3900 1790
rect 3894 1785 3895 1789
rect 3899 1785 3900 1789
rect 3894 1784 3900 1785
rect 110 1780 116 1781
rect 110 1776 111 1780
rect 115 1776 116 1780
rect 110 1775 116 1776
rect 2030 1780 2036 1781
rect 2030 1776 2031 1780
rect 2035 1776 2036 1780
rect 2030 1775 2036 1776
rect 150 1761 156 1762
rect 150 1757 151 1761
rect 155 1757 156 1761
rect 150 1756 156 1757
rect 342 1761 348 1762
rect 342 1757 343 1761
rect 347 1757 348 1761
rect 342 1756 348 1757
rect 542 1761 548 1762
rect 542 1757 543 1761
rect 547 1757 548 1761
rect 542 1756 548 1757
rect 734 1761 740 1762
rect 734 1757 735 1761
rect 739 1757 740 1761
rect 734 1756 740 1757
rect 918 1761 924 1762
rect 918 1757 919 1761
rect 923 1757 924 1761
rect 918 1756 924 1757
rect 1094 1761 1100 1762
rect 1094 1757 1095 1761
rect 1099 1757 1100 1761
rect 1094 1756 1100 1757
rect 1270 1761 1276 1762
rect 1270 1757 1271 1761
rect 1275 1757 1276 1761
rect 1270 1756 1276 1757
rect 1446 1761 1452 1762
rect 1446 1757 1447 1761
rect 1451 1757 1452 1761
rect 1446 1756 1452 1757
rect 1622 1761 1628 1762
rect 1622 1757 1623 1761
rect 1627 1757 1628 1761
rect 1622 1756 1628 1757
rect 1806 1761 1812 1762
rect 1806 1757 1807 1761
rect 1811 1757 1812 1761
rect 1806 1756 1812 1757
rect 2110 1755 2116 1756
rect 2110 1751 2111 1755
rect 2115 1751 2116 1755
rect 2110 1750 2116 1751
rect 2238 1755 2244 1756
rect 2238 1751 2239 1755
rect 2243 1751 2244 1755
rect 2238 1750 2244 1751
rect 2398 1755 2404 1756
rect 2398 1751 2399 1755
rect 2403 1751 2404 1755
rect 2398 1750 2404 1751
rect 2574 1755 2580 1756
rect 2574 1751 2575 1755
rect 2579 1751 2580 1755
rect 2574 1750 2580 1751
rect 2750 1755 2756 1756
rect 2750 1751 2751 1755
rect 2755 1751 2756 1755
rect 2750 1750 2756 1751
rect 2934 1755 2940 1756
rect 2934 1751 2935 1755
rect 2939 1751 2940 1755
rect 2934 1750 2940 1751
rect 3126 1755 3132 1756
rect 3126 1751 3127 1755
rect 3131 1751 3132 1755
rect 3126 1750 3132 1751
rect 3318 1755 3324 1756
rect 3318 1751 3319 1755
rect 3323 1751 3324 1755
rect 3318 1750 3324 1751
rect 3510 1755 3516 1756
rect 3510 1751 3511 1755
rect 3515 1751 3516 1755
rect 3510 1750 3516 1751
rect 3710 1755 3716 1756
rect 3710 1751 3711 1755
rect 3715 1751 3716 1755
rect 3710 1750 3716 1751
rect 3894 1755 3900 1756
rect 3894 1751 3895 1755
rect 3899 1751 3900 1755
rect 3894 1750 3900 1751
rect 2070 1736 2076 1737
rect 2070 1732 2071 1736
rect 2075 1732 2076 1736
rect 2070 1731 2076 1732
rect 3990 1736 3996 1737
rect 3990 1732 3991 1736
rect 3995 1732 3996 1736
rect 3990 1731 3996 1732
rect 150 1727 156 1728
rect 150 1723 151 1727
rect 155 1723 156 1727
rect 150 1722 156 1723
rect 318 1727 324 1728
rect 318 1723 319 1727
rect 323 1723 324 1727
rect 318 1722 324 1723
rect 526 1727 532 1728
rect 526 1723 527 1727
rect 531 1723 532 1727
rect 526 1722 532 1723
rect 742 1727 748 1728
rect 742 1723 743 1727
rect 747 1723 748 1727
rect 742 1722 748 1723
rect 958 1727 964 1728
rect 958 1723 959 1727
rect 963 1723 964 1727
rect 958 1722 964 1723
rect 1166 1727 1172 1728
rect 1166 1723 1167 1727
rect 1171 1723 1172 1727
rect 1166 1722 1172 1723
rect 1366 1727 1372 1728
rect 1366 1723 1367 1727
rect 1371 1723 1372 1727
rect 1366 1722 1372 1723
rect 1558 1727 1564 1728
rect 1558 1723 1559 1727
rect 1563 1723 1564 1727
rect 1558 1722 1564 1723
rect 1758 1727 1764 1728
rect 1758 1723 1759 1727
rect 1763 1723 1764 1727
rect 1758 1722 1764 1723
rect 1934 1727 1940 1728
rect 1934 1723 1935 1727
rect 1939 1723 1940 1727
rect 1934 1722 1940 1723
rect 2070 1719 2076 1720
rect 2070 1715 2071 1719
rect 2075 1715 2076 1719
rect 3990 1719 3996 1720
rect 3990 1715 3991 1719
rect 3995 1715 3996 1719
rect 2070 1714 2076 1715
rect 2110 1714 2116 1715
rect 2110 1710 2111 1714
rect 2115 1710 2116 1714
rect 2110 1709 2116 1710
rect 2238 1714 2244 1715
rect 2238 1710 2239 1714
rect 2243 1710 2244 1714
rect 2238 1709 2244 1710
rect 2398 1714 2404 1715
rect 2398 1710 2399 1714
rect 2403 1710 2404 1714
rect 2398 1709 2404 1710
rect 2574 1714 2580 1715
rect 2574 1710 2575 1714
rect 2579 1710 2580 1714
rect 2574 1709 2580 1710
rect 2750 1714 2756 1715
rect 2750 1710 2751 1714
rect 2755 1710 2756 1714
rect 2750 1709 2756 1710
rect 2934 1714 2940 1715
rect 2934 1710 2935 1714
rect 2939 1710 2940 1714
rect 2934 1709 2940 1710
rect 3126 1714 3132 1715
rect 3126 1710 3127 1714
rect 3131 1710 3132 1714
rect 3126 1709 3132 1710
rect 3318 1714 3324 1715
rect 3318 1710 3319 1714
rect 3323 1710 3324 1714
rect 3318 1709 3324 1710
rect 3510 1714 3516 1715
rect 3510 1710 3511 1714
rect 3515 1710 3516 1714
rect 3510 1709 3516 1710
rect 3710 1714 3716 1715
rect 3710 1710 3711 1714
rect 3715 1710 3716 1714
rect 3710 1709 3716 1710
rect 3894 1714 3900 1715
rect 3990 1714 3996 1715
rect 3894 1710 3895 1714
rect 3899 1710 3900 1714
rect 3894 1709 3900 1710
rect 110 1708 116 1709
rect 110 1704 111 1708
rect 115 1704 116 1708
rect 110 1703 116 1704
rect 2030 1708 2036 1709
rect 2030 1704 2031 1708
rect 2035 1704 2036 1708
rect 2030 1703 2036 1704
rect 110 1691 116 1692
rect 110 1687 111 1691
rect 115 1687 116 1691
rect 2030 1691 2036 1692
rect 2030 1687 2031 1691
rect 2035 1687 2036 1691
rect 110 1686 116 1687
rect 150 1686 156 1687
rect 150 1682 151 1686
rect 155 1682 156 1686
rect 150 1681 156 1682
rect 318 1686 324 1687
rect 318 1682 319 1686
rect 323 1682 324 1686
rect 318 1681 324 1682
rect 526 1686 532 1687
rect 526 1682 527 1686
rect 531 1682 532 1686
rect 526 1681 532 1682
rect 742 1686 748 1687
rect 742 1682 743 1686
rect 747 1682 748 1686
rect 742 1681 748 1682
rect 958 1686 964 1687
rect 958 1682 959 1686
rect 963 1682 964 1686
rect 958 1681 964 1682
rect 1166 1686 1172 1687
rect 1166 1682 1167 1686
rect 1171 1682 1172 1686
rect 1166 1681 1172 1682
rect 1366 1686 1372 1687
rect 1366 1682 1367 1686
rect 1371 1682 1372 1686
rect 1366 1681 1372 1682
rect 1558 1686 1564 1687
rect 1558 1682 1559 1686
rect 1563 1682 1564 1686
rect 1558 1681 1564 1682
rect 1758 1686 1764 1687
rect 1758 1682 1759 1686
rect 1763 1682 1764 1686
rect 1758 1681 1764 1682
rect 1934 1686 1940 1687
rect 2030 1686 2036 1687
rect 1934 1682 1935 1686
rect 1939 1682 1940 1686
rect 1934 1681 1940 1682
rect 2110 1674 2116 1675
rect 2110 1670 2111 1674
rect 2115 1670 2116 1674
rect 2070 1669 2076 1670
rect 2110 1669 2116 1670
rect 2310 1674 2316 1675
rect 2310 1670 2311 1674
rect 2315 1670 2316 1674
rect 2310 1669 2316 1670
rect 2526 1674 2532 1675
rect 2526 1670 2527 1674
rect 2531 1670 2532 1674
rect 2526 1669 2532 1670
rect 2742 1674 2748 1675
rect 2742 1670 2743 1674
rect 2747 1670 2748 1674
rect 2742 1669 2748 1670
rect 2950 1674 2956 1675
rect 2950 1670 2951 1674
rect 2955 1670 2956 1674
rect 2950 1669 2956 1670
rect 3150 1674 3156 1675
rect 3150 1670 3151 1674
rect 3155 1670 3156 1674
rect 3150 1669 3156 1670
rect 3342 1674 3348 1675
rect 3342 1670 3343 1674
rect 3347 1670 3348 1674
rect 3342 1669 3348 1670
rect 3526 1674 3532 1675
rect 3526 1670 3527 1674
rect 3531 1670 3532 1674
rect 3526 1669 3532 1670
rect 3718 1674 3724 1675
rect 3718 1670 3719 1674
rect 3723 1670 3724 1674
rect 3718 1669 3724 1670
rect 3894 1674 3900 1675
rect 3894 1670 3895 1674
rect 3899 1670 3900 1674
rect 3894 1669 3900 1670
rect 3990 1669 3996 1670
rect 2070 1665 2071 1669
rect 2075 1665 2076 1669
rect 2070 1664 2076 1665
rect 3990 1665 3991 1669
rect 3995 1665 3996 1669
rect 3990 1664 3996 1665
rect 150 1654 156 1655
rect 150 1650 151 1654
rect 155 1650 156 1654
rect 110 1649 116 1650
rect 150 1649 156 1650
rect 318 1654 324 1655
rect 318 1650 319 1654
rect 323 1650 324 1654
rect 318 1649 324 1650
rect 502 1654 508 1655
rect 502 1650 503 1654
rect 507 1650 508 1654
rect 502 1649 508 1650
rect 694 1654 700 1655
rect 694 1650 695 1654
rect 699 1650 700 1654
rect 694 1649 700 1650
rect 886 1654 892 1655
rect 886 1650 887 1654
rect 891 1650 892 1654
rect 886 1649 892 1650
rect 1078 1654 1084 1655
rect 1078 1650 1079 1654
rect 1083 1650 1084 1654
rect 1078 1649 1084 1650
rect 1262 1654 1268 1655
rect 1262 1650 1263 1654
rect 1267 1650 1268 1654
rect 1262 1649 1268 1650
rect 1438 1654 1444 1655
rect 1438 1650 1439 1654
rect 1443 1650 1444 1654
rect 1438 1649 1444 1650
rect 1614 1654 1620 1655
rect 1614 1650 1615 1654
rect 1619 1650 1620 1654
rect 1614 1649 1620 1650
rect 1790 1654 1796 1655
rect 1790 1650 1791 1654
rect 1795 1650 1796 1654
rect 2070 1652 2076 1653
rect 1790 1649 1796 1650
rect 2030 1649 2036 1650
rect 110 1645 111 1649
rect 115 1645 116 1649
rect 110 1644 116 1645
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2070 1648 2071 1652
rect 2075 1648 2076 1652
rect 2070 1647 2076 1648
rect 3990 1652 3996 1653
rect 3990 1648 3991 1652
rect 3995 1648 3996 1652
rect 3990 1647 3996 1648
rect 2030 1644 2036 1645
rect 2110 1633 2116 1634
rect 110 1632 116 1633
rect 110 1628 111 1632
rect 115 1628 116 1632
rect 110 1627 116 1628
rect 2030 1632 2036 1633
rect 2030 1628 2031 1632
rect 2035 1628 2036 1632
rect 2110 1629 2111 1633
rect 2115 1629 2116 1633
rect 2110 1628 2116 1629
rect 2310 1633 2316 1634
rect 2310 1629 2311 1633
rect 2315 1629 2316 1633
rect 2310 1628 2316 1629
rect 2526 1633 2532 1634
rect 2526 1629 2527 1633
rect 2531 1629 2532 1633
rect 2526 1628 2532 1629
rect 2742 1633 2748 1634
rect 2742 1629 2743 1633
rect 2747 1629 2748 1633
rect 2742 1628 2748 1629
rect 2950 1633 2956 1634
rect 2950 1629 2951 1633
rect 2955 1629 2956 1633
rect 2950 1628 2956 1629
rect 3150 1633 3156 1634
rect 3150 1629 3151 1633
rect 3155 1629 3156 1633
rect 3150 1628 3156 1629
rect 3342 1633 3348 1634
rect 3342 1629 3343 1633
rect 3347 1629 3348 1633
rect 3342 1628 3348 1629
rect 3526 1633 3532 1634
rect 3526 1629 3527 1633
rect 3531 1629 3532 1633
rect 3526 1628 3532 1629
rect 3718 1633 3724 1634
rect 3718 1629 3719 1633
rect 3723 1629 3724 1633
rect 3718 1628 3724 1629
rect 3894 1633 3900 1634
rect 3894 1629 3895 1633
rect 3899 1629 3900 1633
rect 3894 1628 3900 1629
rect 2030 1627 2036 1628
rect 150 1613 156 1614
rect 150 1609 151 1613
rect 155 1609 156 1613
rect 150 1608 156 1609
rect 318 1613 324 1614
rect 318 1609 319 1613
rect 323 1609 324 1613
rect 318 1608 324 1609
rect 502 1613 508 1614
rect 502 1609 503 1613
rect 507 1609 508 1613
rect 502 1608 508 1609
rect 694 1613 700 1614
rect 694 1609 695 1613
rect 699 1609 700 1613
rect 694 1608 700 1609
rect 886 1613 892 1614
rect 886 1609 887 1613
rect 891 1609 892 1613
rect 886 1608 892 1609
rect 1078 1613 1084 1614
rect 1078 1609 1079 1613
rect 1083 1609 1084 1613
rect 1078 1608 1084 1609
rect 1262 1613 1268 1614
rect 1262 1609 1263 1613
rect 1267 1609 1268 1613
rect 1262 1608 1268 1609
rect 1438 1613 1444 1614
rect 1438 1609 1439 1613
rect 1443 1609 1444 1613
rect 1438 1608 1444 1609
rect 1614 1613 1620 1614
rect 1614 1609 1615 1613
rect 1619 1609 1620 1613
rect 1614 1608 1620 1609
rect 1790 1613 1796 1614
rect 1790 1609 1791 1613
rect 1795 1609 1796 1613
rect 1790 1608 1796 1609
rect 2478 1591 2484 1592
rect 2478 1587 2479 1591
rect 2483 1587 2484 1591
rect 2478 1586 2484 1587
rect 2582 1591 2588 1592
rect 2582 1587 2583 1591
rect 2587 1587 2588 1591
rect 2582 1586 2588 1587
rect 2694 1591 2700 1592
rect 2694 1587 2695 1591
rect 2699 1587 2700 1591
rect 2694 1586 2700 1587
rect 2814 1591 2820 1592
rect 2814 1587 2815 1591
rect 2819 1587 2820 1591
rect 2814 1586 2820 1587
rect 2942 1591 2948 1592
rect 2942 1587 2943 1591
rect 2947 1587 2948 1591
rect 2942 1586 2948 1587
rect 3078 1591 3084 1592
rect 3078 1587 3079 1591
rect 3083 1587 3084 1591
rect 3078 1586 3084 1587
rect 3222 1591 3228 1592
rect 3222 1587 3223 1591
rect 3227 1587 3228 1591
rect 3222 1586 3228 1587
rect 3382 1591 3388 1592
rect 3382 1587 3383 1591
rect 3387 1587 3388 1591
rect 3382 1586 3388 1587
rect 3550 1591 3556 1592
rect 3550 1587 3551 1591
rect 3555 1587 3556 1591
rect 3550 1586 3556 1587
rect 3726 1591 3732 1592
rect 3726 1587 3727 1591
rect 3731 1587 3732 1591
rect 3726 1586 3732 1587
rect 3894 1591 3900 1592
rect 3894 1587 3895 1591
rect 3899 1587 3900 1591
rect 3894 1586 3900 1587
rect 318 1575 324 1576
rect 318 1571 319 1575
rect 323 1571 324 1575
rect 318 1570 324 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 598 1575 604 1576
rect 598 1571 599 1575
rect 603 1571 604 1575
rect 598 1570 604 1571
rect 742 1575 748 1576
rect 742 1571 743 1575
rect 747 1571 748 1575
rect 742 1570 748 1571
rect 886 1575 892 1576
rect 886 1571 887 1575
rect 891 1571 892 1575
rect 886 1570 892 1571
rect 1030 1575 1036 1576
rect 1030 1571 1031 1575
rect 1035 1571 1036 1575
rect 1030 1570 1036 1571
rect 1174 1575 1180 1576
rect 1174 1571 1175 1575
rect 1179 1571 1180 1575
rect 1174 1570 1180 1571
rect 1318 1575 1324 1576
rect 1318 1571 1319 1575
rect 1323 1571 1324 1575
rect 1318 1570 1324 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1622 1575 1628 1576
rect 1622 1571 1623 1575
rect 1627 1571 1628 1575
rect 1622 1570 1628 1571
rect 2070 1572 2076 1573
rect 2070 1568 2071 1572
rect 2075 1568 2076 1572
rect 2070 1567 2076 1568
rect 3990 1572 3996 1573
rect 3990 1568 3991 1572
rect 3995 1568 3996 1572
rect 3990 1567 3996 1568
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 110 1551 116 1552
rect 2030 1556 2036 1557
rect 2030 1552 2031 1556
rect 2035 1552 2036 1556
rect 2030 1551 2036 1552
rect 2070 1555 2076 1556
rect 2070 1551 2071 1555
rect 2075 1551 2076 1555
rect 3990 1555 3996 1556
rect 3990 1551 3991 1555
rect 3995 1551 3996 1555
rect 2070 1550 2076 1551
rect 2478 1550 2484 1551
rect 2478 1546 2479 1550
rect 2483 1546 2484 1550
rect 2478 1545 2484 1546
rect 2582 1550 2588 1551
rect 2582 1546 2583 1550
rect 2587 1546 2588 1550
rect 2582 1545 2588 1546
rect 2694 1550 2700 1551
rect 2694 1546 2695 1550
rect 2699 1546 2700 1550
rect 2694 1545 2700 1546
rect 2814 1550 2820 1551
rect 2814 1546 2815 1550
rect 2819 1546 2820 1550
rect 2814 1545 2820 1546
rect 2942 1550 2948 1551
rect 2942 1546 2943 1550
rect 2947 1546 2948 1550
rect 2942 1545 2948 1546
rect 3078 1550 3084 1551
rect 3078 1546 3079 1550
rect 3083 1546 3084 1550
rect 3078 1545 3084 1546
rect 3222 1550 3228 1551
rect 3222 1546 3223 1550
rect 3227 1546 3228 1550
rect 3222 1545 3228 1546
rect 3382 1550 3388 1551
rect 3382 1546 3383 1550
rect 3387 1546 3388 1550
rect 3382 1545 3388 1546
rect 3550 1550 3556 1551
rect 3550 1546 3551 1550
rect 3555 1546 3556 1550
rect 3550 1545 3556 1546
rect 3726 1550 3732 1551
rect 3726 1546 3727 1550
rect 3731 1546 3732 1550
rect 3726 1545 3732 1546
rect 3894 1550 3900 1551
rect 3990 1550 3996 1551
rect 3894 1546 3895 1550
rect 3899 1546 3900 1550
rect 3894 1545 3900 1546
rect 110 1539 116 1540
rect 110 1535 111 1539
rect 115 1535 116 1539
rect 2030 1539 2036 1540
rect 2030 1535 2031 1539
rect 2035 1535 2036 1539
rect 110 1534 116 1535
rect 318 1534 324 1535
rect 318 1530 319 1534
rect 323 1530 324 1534
rect 318 1529 324 1530
rect 454 1534 460 1535
rect 454 1530 455 1534
rect 459 1530 460 1534
rect 454 1529 460 1530
rect 598 1534 604 1535
rect 598 1530 599 1534
rect 603 1530 604 1534
rect 598 1529 604 1530
rect 742 1534 748 1535
rect 742 1530 743 1534
rect 747 1530 748 1534
rect 742 1529 748 1530
rect 886 1534 892 1535
rect 886 1530 887 1534
rect 891 1530 892 1534
rect 886 1529 892 1530
rect 1030 1534 1036 1535
rect 1030 1530 1031 1534
rect 1035 1530 1036 1534
rect 1030 1529 1036 1530
rect 1174 1534 1180 1535
rect 1174 1530 1175 1534
rect 1179 1530 1180 1534
rect 1174 1529 1180 1530
rect 1318 1534 1324 1535
rect 1318 1530 1319 1534
rect 1323 1530 1324 1534
rect 1318 1529 1324 1530
rect 1470 1534 1476 1535
rect 1470 1530 1471 1534
rect 1475 1530 1476 1534
rect 1470 1529 1476 1530
rect 1622 1534 1628 1535
rect 2030 1534 2036 1535
rect 1622 1530 1623 1534
rect 1627 1530 1628 1534
rect 1622 1529 1628 1530
rect 2486 1506 2492 1507
rect 2486 1502 2487 1506
rect 2491 1502 2492 1506
rect 2070 1501 2076 1502
rect 2486 1501 2492 1502
rect 2590 1506 2596 1507
rect 2590 1502 2591 1506
rect 2595 1502 2596 1506
rect 2590 1501 2596 1502
rect 2694 1506 2700 1507
rect 2694 1502 2695 1506
rect 2699 1502 2700 1506
rect 2694 1501 2700 1502
rect 2806 1506 2812 1507
rect 2806 1502 2807 1506
rect 2811 1502 2812 1506
rect 2806 1501 2812 1502
rect 2934 1506 2940 1507
rect 2934 1502 2935 1506
rect 2939 1502 2940 1506
rect 2934 1501 2940 1502
rect 3070 1506 3076 1507
rect 3070 1502 3071 1506
rect 3075 1502 3076 1506
rect 3070 1501 3076 1502
rect 3222 1506 3228 1507
rect 3222 1502 3223 1506
rect 3227 1502 3228 1506
rect 3222 1501 3228 1502
rect 3382 1506 3388 1507
rect 3382 1502 3383 1506
rect 3387 1502 3388 1506
rect 3382 1501 3388 1502
rect 3550 1506 3556 1507
rect 3550 1502 3551 1506
rect 3555 1502 3556 1506
rect 3550 1501 3556 1502
rect 3718 1506 3724 1507
rect 3718 1502 3719 1506
rect 3723 1502 3724 1506
rect 3718 1501 3724 1502
rect 3894 1506 3900 1507
rect 3894 1502 3895 1506
rect 3899 1502 3900 1506
rect 3894 1501 3900 1502
rect 3990 1501 3996 1502
rect 2070 1497 2071 1501
rect 2075 1497 2076 1501
rect 2070 1496 2076 1497
rect 3990 1497 3991 1501
rect 3995 1497 3996 1501
rect 3990 1496 3996 1497
rect 358 1494 364 1495
rect 358 1490 359 1494
rect 363 1490 364 1494
rect 110 1489 116 1490
rect 358 1489 364 1490
rect 486 1494 492 1495
rect 486 1490 487 1494
rect 491 1490 492 1494
rect 486 1489 492 1490
rect 622 1494 628 1495
rect 622 1490 623 1494
rect 627 1490 628 1494
rect 622 1489 628 1490
rect 774 1494 780 1495
rect 774 1490 775 1494
rect 779 1490 780 1494
rect 774 1489 780 1490
rect 926 1494 932 1495
rect 926 1490 927 1494
rect 931 1490 932 1494
rect 926 1489 932 1490
rect 1086 1494 1092 1495
rect 1086 1490 1087 1494
rect 1091 1490 1092 1494
rect 1086 1489 1092 1490
rect 1254 1494 1260 1495
rect 1254 1490 1255 1494
rect 1259 1490 1260 1494
rect 1254 1489 1260 1490
rect 1422 1494 1428 1495
rect 1422 1490 1423 1494
rect 1427 1490 1428 1494
rect 1422 1489 1428 1490
rect 1590 1494 1596 1495
rect 1590 1490 1591 1494
rect 1595 1490 1596 1494
rect 1590 1489 1596 1490
rect 1766 1494 1772 1495
rect 1766 1490 1767 1494
rect 1771 1490 1772 1494
rect 1766 1489 1772 1490
rect 2030 1489 2036 1490
rect 110 1485 111 1489
rect 115 1485 116 1489
rect 110 1484 116 1485
rect 2030 1485 2031 1489
rect 2035 1485 2036 1489
rect 2030 1484 2036 1485
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 3990 1484 3996 1485
rect 3990 1480 3991 1484
rect 3995 1480 3996 1484
rect 3990 1479 3996 1480
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 110 1467 116 1468
rect 2030 1472 2036 1473
rect 2030 1468 2031 1472
rect 2035 1468 2036 1472
rect 2030 1467 2036 1468
rect 2486 1465 2492 1466
rect 2486 1461 2487 1465
rect 2491 1461 2492 1465
rect 2486 1460 2492 1461
rect 2590 1465 2596 1466
rect 2590 1461 2591 1465
rect 2595 1461 2596 1465
rect 2590 1460 2596 1461
rect 2694 1465 2700 1466
rect 2694 1461 2695 1465
rect 2699 1461 2700 1465
rect 2694 1460 2700 1461
rect 2806 1465 2812 1466
rect 2806 1461 2807 1465
rect 2811 1461 2812 1465
rect 2806 1460 2812 1461
rect 2934 1465 2940 1466
rect 2934 1461 2935 1465
rect 2939 1461 2940 1465
rect 2934 1460 2940 1461
rect 3070 1465 3076 1466
rect 3070 1461 3071 1465
rect 3075 1461 3076 1465
rect 3070 1460 3076 1461
rect 3222 1465 3228 1466
rect 3222 1461 3223 1465
rect 3227 1461 3228 1465
rect 3222 1460 3228 1461
rect 3382 1465 3388 1466
rect 3382 1461 3383 1465
rect 3387 1461 3388 1465
rect 3382 1460 3388 1461
rect 3550 1465 3556 1466
rect 3550 1461 3551 1465
rect 3555 1461 3556 1465
rect 3550 1460 3556 1461
rect 3718 1465 3724 1466
rect 3718 1461 3719 1465
rect 3723 1461 3724 1465
rect 3718 1460 3724 1461
rect 3894 1465 3900 1466
rect 3894 1461 3895 1465
rect 3899 1461 3900 1465
rect 3894 1460 3900 1461
rect 358 1453 364 1454
rect 358 1449 359 1453
rect 363 1449 364 1453
rect 358 1448 364 1449
rect 486 1453 492 1454
rect 486 1449 487 1453
rect 491 1449 492 1453
rect 486 1448 492 1449
rect 622 1453 628 1454
rect 622 1449 623 1453
rect 627 1449 628 1453
rect 622 1448 628 1449
rect 774 1453 780 1454
rect 774 1449 775 1453
rect 779 1449 780 1453
rect 774 1448 780 1449
rect 926 1453 932 1454
rect 926 1449 927 1453
rect 931 1449 932 1453
rect 926 1448 932 1449
rect 1086 1453 1092 1454
rect 1086 1449 1087 1453
rect 1091 1449 1092 1453
rect 1086 1448 1092 1449
rect 1254 1453 1260 1454
rect 1254 1449 1255 1453
rect 1259 1449 1260 1453
rect 1254 1448 1260 1449
rect 1422 1453 1428 1454
rect 1422 1449 1423 1453
rect 1427 1449 1428 1453
rect 1422 1448 1428 1449
rect 1590 1453 1596 1454
rect 1590 1449 1591 1453
rect 1595 1449 1596 1453
rect 1590 1448 1596 1449
rect 1766 1453 1772 1454
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 2238 1431 2244 1432
rect 2238 1427 2239 1431
rect 2243 1427 2244 1431
rect 2238 1426 2244 1427
rect 2350 1431 2356 1432
rect 2350 1427 2351 1431
rect 2355 1427 2356 1431
rect 2350 1426 2356 1427
rect 2470 1431 2476 1432
rect 2470 1427 2471 1431
rect 2475 1427 2476 1431
rect 2470 1426 2476 1427
rect 2590 1431 2596 1432
rect 2590 1427 2591 1431
rect 2595 1427 2596 1431
rect 2590 1426 2596 1427
rect 2726 1431 2732 1432
rect 2726 1427 2727 1431
rect 2731 1427 2732 1431
rect 2726 1426 2732 1427
rect 2878 1431 2884 1432
rect 2878 1427 2879 1431
rect 2883 1427 2884 1431
rect 2878 1426 2884 1427
rect 3054 1431 3060 1432
rect 3054 1427 3055 1431
rect 3059 1427 3060 1431
rect 3054 1426 3060 1427
rect 3246 1431 3252 1432
rect 3246 1427 3247 1431
rect 3251 1427 3252 1431
rect 3246 1426 3252 1427
rect 3454 1431 3460 1432
rect 3454 1427 3455 1431
rect 3459 1427 3460 1431
rect 3454 1426 3460 1427
rect 3670 1431 3676 1432
rect 3670 1427 3671 1431
rect 3675 1427 3676 1431
rect 3670 1426 3676 1427
rect 3886 1431 3892 1432
rect 3886 1427 3887 1431
rect 3891 1427 3892 1431
rect 3886 1426 3892 1427
rect 150 1415 156 1416
rect 150 1411 151 1415
rect 155 1411 156 1415
rect 150 1410 156 1411
rect 270 1415 276 1416
rect 270 1411 271 1415
rect 275 1411 276 1415
rect 270 1410 276 1411
rect 430 1415 436 1416
rect 430 1411 431 1415
rect 435 1411 436 1415
rect 430 1410 436 1411
rect 614 1415 620 1416
rect 614 1411 615 1415
rect 619 1411 620 1415
rect 614 1410 620 1411
rect 806 1415 812 1416
rect 806 1411 807 1415
rect 811 1411 812 1415
rect 806 1410 812 1411
rect 1006 1415 1012 1416
rect 1006 1411 1007 1415
rect 1011 1411 1012 1415
rect 1006 1410 1012 1411
rect 1214 1415 1220 1416
rect 1214 1411 1215 1415
rect 1219 1411 1220 1415
rect 1214 1410 1220 1411
rect 1422 1415 1428 1416
rect 1422 1411 1423 1415
rect 1427 1411 1428 1415
rect 1422 1410 1428 1411
rect 1630 1415 1636 1416
rect 1630 1411 1631 1415
rect 1635 1411 1636 1415
rect 1630 1410 1636 1411
rect 1846 1415 1852 1416
rect 1846 1411 1847 1415
rect 1851 1411 1852 1415
rect 1846 1410 1852 1411
rect 2070 1412 2076 1413
rect 2070 1408 2071 1412
rect 2075 1408 2076 1412
rect 2070 1407 2076 1408
rect 3990 1412 3996 1413
rect 3990 1408 3991 1412
rect 3995 1408 3996 1412
rect 3990 1407 3996 1408
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 110 1391 116 1392
rect 2030 1396 2036 1397
rect 2030 1392 2031 1396
rect 2035 1392 2036 1396
rect 2030 1391 2036 1392
rect 2070 1395 2076 1396
rect 2070 1391 2071 1395
rect 2075 1391 2076 1395
rect 3990 1395 3996 1396
rect 3990 1391 3991 1395
rect 3995 1391 3996 1395
rect 2070 1390 2076 1391
rect 2238 1390 2244 1391
rect 2238 1386 2239 1390
rect 2243 1386 2244 1390
rect 2238 1385 2244 1386
rect 2350 1390 2356 1391
rect 2350 1386 2351 1390
rect 2355 1386 2356 1390
rect 2350 1385 2356 1386
rect 2470 1390 2476 1391
rect 2470 1386 2471 1390
rect 2475 1386 2476 1390
rect 2470 1385 2476 1386
rect 2590 1390 2596 1391
rect 2590 1386 2591 1390
rect 2595 1386 2596 1390
rect 2590 1385 2596 1386
rect 2726 1390 2732 1391
rect 2726 1386 2727 1390
rect 2731 1386 2732 1390
rect 2726 1385 2732 1386
rect 2878 1390 2884 1391
rect 2878 1386 2879 1390
rect 2883 1386 2884 1390
rect 2878 1385 2884 1386
rect 3054 1390 3060 1391
rect 3054 1386 3055 1390
rect 3059 1386 3060 1390
rect 3054 1385 3060 1386
rect 3246 1390 3252 1391
rect 3246 1386 3247 1390
rect 3251 1386 3252 1390
rect 3246 1385 3252 1386
rect 3454 1390 3460 1391
rect 3454 1386 3455 1390
rect 3459 1386 3460 1390
rect 3454 1385 3460 1386
rect 3670 1390 3676 1391
rect 3670 1386 3671 1390
rect 3675 1386 3676 1390
rect 3670 1385 3676 1386
rect 3886 1390 3892 1391
rect 3990 1390 3996 1391
rect 3886 1386 3887 1390
rect 3891 1386 3892 1390
rect 3886 1385 3892 1386
rect 110 1379 116 1380
rect 110 1375 111 1379
rect 115 1375 116 1379
rect 2030 1379 2036 1380
rect 2030 1375 2031 1379
rect 2035 1375 2036 1379
rect 110 1374 116 1375
rect 150 1374 156 1375
rect 150 1370 151 1374
rect 155 1370 156 1374
rect 150 1369 156 1370
rect 270 1374 276 1375
rect 270 1370 271 1374
rect 275 1370 276 1374
rect 270 1369 276 1370
rect 430 1374 436 1375
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 614 1374 620 1375
rect 614 1370 615 1374
rect 619 1370 620 1374
rect 614 1369 620 1370
rect 806 1374 812 1375
rect 806 1370 807 1374
rect 811 1370 812 1374
rect 806 1369 812 1370
rect 1006 1374 1012 1375
rect 1006 1370 1007 1374
rect 1011 1370 1012 1374
rect 1006 1369 1012 1370
rect 1214 1374 1220 1375
rect 1214 1370 1215 1374
rect 1219 1370 1220 1374
rect 1214 1369 1220 1370
rect 1422 1374 1428 1375
rect 1422 1370 1423 1374
rect 1427 1370 1428 1374
rect 1422 1369 1428 1370
rect 1630 1374 1636 1375
rect 1630 1370 1631 1374
rect 1635 1370 1636 1374
rect 1630 1369 1636 1370
rect 1846 1374 1852 1375
rect 2030 1374 2036 1375
rect 1846 1370 1847 1374
rect 1851 1370 1852 1374
rect 1846 1369 1852 1370
rect 2390 1350 2396 1351
rect 2390 1346 2391 1350
rect 2395 1346 2396 1350
rect 2070 1345 2076 1346
rect 2390 1345 2396 1346
rect 2526 1350 2532 1351
rect 2526 1346 2527 1350
rect 2531 1346 2532 1350
rect 2526 1345 2532 1346
rect 2678 1350 2684 1351
rect 2678 1346 2679 1350
rect 2683 1346 2684 1350
rect 2678 1345 2684 1346
rect 2838 1350 2844 1351
rect 2838 1346 2839 1350
rect 2843 1346 2844 1350
rect 2838 1345 2844 1346
rect 2998 1350 3004 1351
rect 2998 1346 2999 1350
rect 3003 1346 3004 1350
rect 2998 1345 3004 1346
rect 3166 1350 3172 1351
rect 3166 1346 3167 1350
rect 3171 1346 3172 1350
rect 3166 1345 3172 1346
rect 3342 1350 3348 1351
rect 3342 1346 3343 1350
rect 3347 1346 3348 1350
rect 3342 1345 3348 1346
rect 3518 1350 3524 1351
rect 3518 1346 3519 1350
rect 3523 1346 3524 1350
rect 3518 1345 3524 1346
rect 3694 1350 3700 1351
rect 3694 1346 3695 1350
rect 3699 1346 3700 1350
rect 3694 1345 3700 1346
rect 3878 1350 3884 1351
rect 3878 1346 3879 1350
rect 3883 1346 3884 1350
rect 3878 1345 3884 1346
rect 3990 1345 3996 1346
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 2070 1340 2076 1341
rect 3990 1341 3991 1345
rect 3995 1341 3996 1345
rect 3990 1340 3996 1341
rect 150 1330 156 1331
rect 150 1326 151 1330
rect 155 1326 156 1330
rect 110 1325 116 1326
rect 150 1325 156 1326
rect 286 1330 292 1331
rect 286 1326 287 1330
rect 291 1326 292 1330
rect 286 1325 292 1326
rect 462 1330 468 1331
rect 462 1326 463 1330
rect 467 1326 468 1330
rect 462 1325 468 1326
rect 662 1330 668 1331
rect 662 1326 663 1330
rect 667 1326 668 1330
rect 662 1325 668 1326
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 862 1325 868 1326
rect 1062 1330 1068 1331
rect 1062 1326 1063 1330
rect 1067 1326 1068 1330
rect 1062 1325 1068 1326
rect 1254 1330 1260 1331
rect 1254 1326 1255 1330
rect 1259 1326 1260 1330
rect 1254 1325 1260 1326
rect 1430 1330 1436 1331
rect 1430 1326 1431 1330
rect 1435 1326 1436 1330
rect 1430 1325 1436 1326
rect 1606 1330 1612 1331
rect 1606 1326 1607 1330
rect 1611 1326 1612 1330
rect 1606 1325 1612 1326
rect 1782 1330 1788 1331
rect 1782 1326 1783 1330
rect 1787 1326 1788 1330
rect 1782 1325 1788 1326
rect 1934 1330 1940 1331
rect 1934 1326 1935 1330
rect 1939 1326 1940 1330
rect 2070 1328 2076 1329
rect 1934 1325 1940 1326
rect 2030 1325 2036 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 110 1320 116 1321
rect 2030 1321 2031 1325
rect 2035 1321 2036 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 3990 1328 3996 1329
rect 3990 1324 3991 1328
rect 3995 1324 3996 1328
rect 3990 1323 3996 1324
rect 2030 1320 2036 1321
rect 2390 1309 2396 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 110 1303 116 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2390 1305 2391 1309
rect 2395 1305 2396 1309
rect 2390 1304 2396 1305
rect 2526 1309 2532 1310
rect 2526 1305 2527 1309
rect 2531 1305 2532 1309
rect 2526 1304 2532 1305
rect 2678 1309 2684 1310
rect 2678 1305 2679 1309
rect 2683 1305 2684 1309
rect 2678 1304 2684 1305
rect 2838 1309 2844 1310
rect 2838 1305 2839 1309
rect 2843 1305 2844 1309
rect 2838 1304 2844 1305
rect 2998 1309 3004 1310
rect 2998 1305 2999 1309
rect 3003 1305 3004 1309
rect 2998 1304 3004 1305
rect 3166 1309 3172 1310
rect 3166 1305 3167 1309
rect 3171 1305 3172 1309
rect 3166 1304 3172 1305
rect 3342 1309 3348 1310
rect 3342 1305 3343 1309
rect 3347 1305 3348 1309
rect 3342 1304 3348 1305
rect 3518 1309 3524 1310
rect 3518 1305 3519 1309
rect 3523 1305 3524 1309
rect 3518 1304 3524 1305
rect 3694 1309 3700 1310
rect 3694 1305 3695 1309
rect 3699 1305 3700 1309
rect 3694 1304 3700 1305
rect 3878 1309 3884 1310
rect 3878 1305 3879 1309
rect 3883 1305 3884 1309
rect 3878 1304 3884 1305
rect 2030 1303 2036 1304
rect 150 1289 156 1290
rect 150 1285 151 1289
rect 155 1285 156 1289
rect 150 1284 156 1285
rect 286 1289 292 1290
rect 286 1285 287 1289
rect 291 1285 292 1289
rect 286 1284 292 1285
rect 462 1289 468 1290
rect 462 1285 463 1289
rect 467 1285 468 1289
rect 462 1284 468 1285
rect 662 1289 668 1290
rect 662 1285 663 1289
rect 667 1285 668 1289
rect 662 1284 668 1285
rect 862 1289 868 1290
rect 862 1285 863 1289
rect 867 1285 868 1289
rect 862 1284 868 1285
rect 1062 1289 1068 1290
rect 1062 1285 1063 1289
rect 1067 1285 1068 1289
rect 1062 1284 1068 1285
rect 1254 1289 1260 1290
rect 1254 1285 1255 1289
rect 1259 1285 1260 1289
rect 1254 1284 1260 1285
rect 1430 1289 1436 1290
rect 1430 1285 1431 1289
rect 1435 1285 1436 1289
rect 1430 1284 1436 1285
rect 1606 1289 1612 1290
rect 1606 1285 1607 1289
rect 1611 1285 1612 1289
rect 1606 1284 1612 1285
rect 1782 1289 1788 1290
rect 1782 1285 1783 1289
rect 1787 1285 1788 1289
rect 1782 1284 1788 1285
rect 1934 1289 1940 1290
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 1934 1284 1940 1285
rect 2110 1271 2116 1272
rect 2110 1267 2111 1271
rect 2115 1267 2116 1271
rect 2110 1266 2116 1267
rect 2342 1271 2348 1272
rect 2342 1267 2343 1271
rect 2347 1267 2348 1271
rect 2342 1266 2348 1267
rect 2582 1271 2588 1272
rect 2582 1267 2583 1271
rect 2587 1267 2588 1271
rect 2582 1266 2588 1267
rect 2798 1271 2804 1272
rect 2798 1267 2799 1271
rect 2803 1267 2804 1271
rect 2798 1266 2804 1267
rect 2998 1271 3004 1272
rect 2998 1267 2999 1271
rect 3003 1267 3004 1271
rect 2998 1266 3004 1267
rect 3182 1271 3188 1272
rect 3182 1267 3183 1271
rect 3187 1267 3188 1271
rect 3182 1266 3188 1267
rect 3342 1271 3348 1272
rect 3342 1267 3343 1271
rect 3347 1267 3348 1271
rect 3342 1266 3348 1267
rect 3494 1271 3500 1272
rect 3494 1267 3495 1271
rect 3499 1267 3500 1271
rect 3494 1266 3500 1267
rect 3638 1271 3644 1272
rect 3638 1267 3639 1271
rect 3643 1267 3644 1271
rect 3638 1266 3644 1267
rect 3774 1271 3780 1272
rect 3774 1267 3775 1271
rect 3779 1267 3780 1271
rect 3774 1266 3780 1267
rect 3894 1271 3900 1272
rect 3894 1267 3895 1271
rect 3899 1267 3900 1271
rect 3894 1266 3900 1267
rect 206 1259 212 1260
rect 206 1255 207 1259
rect 211 1255 212 1259
rect 206 1254 212 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 454 1259 460 1260
rect 454 1255 455 1259
rect 459 1255 460 1259
rect 454 1254 460 1255
rect 582 1259 588 1260
rect 582 1255 583 1259
rect 587 1255 588 1259
rect 582 1254 588 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 878 1259 884 1260
rect 878 1255 879 1259
rect 883 1255 884 1259
rect 878 1254 884 1255
rect 1054 1259 1060 1260
rect 1054 1255 1055 1259
rect 1059 1255 1060 1259
rect 1054 1254 1060 1255
rect 1262 1259 1268 1260
rect 1262 1255 1263 1259
rect 1267 1255 1268 1259
rect 1262 1254 1268 1255
rect 1486 1259 1492 1260
rect 1486 1255 1487 1259
rect 1491 1255 1492 1259
rect 1486 1254 1492 1255
rect 1718 1259 1724 1260
rect 1718 1255 1719 1259
rect 1723 1255 1724 1259
rect 1718 1254 1724 1255
rect 1934 1259 1940 1260
rect 1934 1255 1935 1259
rect 1939 1255 1940 1259
rect 1934 1254 1940 1255
rect 2070 1252 2076 1253
rect 2070 1248 2071 1252
rect 2075 1248 2076 1252
rect 2070 1247 2076 1248
rect 3990 1252 3996 1253
rect 3990 1248 3991 1252
rect 3995 1248 3996 1252
rect 3990 1247 3996 1248
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 2030 1240 2036 1241
rect 2030 1236 2031 1240
rect 2035 1236 2036 1240
rect 2030 1235 2036 1236
rect 2070 1235 2076 1236
rect 2070 1231 2071 1235
rect 2075 1231 2076 1235
rect 3990 1235 3996 1236
rect 3990 1231 3991 1235
rect 3995 1231 3996 1235
rect 2070 1230 2076 1231
rect 2110 1230 2116 1231
rect 2110 1226 2111 1230
rect 2115 1226 2116 1230
rect 2110 1225 2116 1226
rect 2342 1230 2348 1231
rect 2342 1226 2343 1230
rect 2347 1226 2348 1230
rect 2342 1225 2348 1226
rect 2582 1230 2588 1231
rect 2582 1226 2583 1230
rect 2587 1226 2588 1230
rect 2582 1225 2588 1226
rect 2798 1230 2804 1231
rect 2798 1226 2799 1230
rect 2803 1226 2804 1230
rect 2798 1225 2804 1226
rect 2998 1230 3004 1231
rect 2998 1226 2999 1230
rect 3003 1226 3004 1230
rect 2998 1225 3004 1226
rect 3182 1230 3188 1231
rect 3182 1226 3183 1230
rect 3187 1226 3188 1230
rect 3182 1225 3188 1226
rect 3342 1230 3348 1231
rect 3342 1226 3343 1230
rect 3347 1226 3348 1230
rect 3342 1225 3348 1226
rect 3494 1230 3500 1231
rect 3494 1226 3495 1230
rect 3499 1226 3500 1230
rect 3494 1225 3500 1226
rect 3638 1230 3644 1231
rect 3638 1226 3639 1230
rect 3643 1226 3644 1230
rect 3638 1225 3644 1226
rect 3774 1230 3780 1231
rect 3774 1226 3775 1230
rect 3779 1226 3780 1230
rect 3774 1225 3780 1226
rect 3894 1230 3900 1231
rect 3990 1230 3996 1231
rect 3894 1226 3895 1230
rect 3899 1226 3900 1230
rect 3894 1225 3900 1226
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 2030 1223 2036 1224
rect 2030 1219 2031 1223
rect 2035 1219 2036 1223
rect 110 1218 116 1219
rect 206 1218 212 1219
rect 206 1214 207 1218
rect 211 1214 212 1218
rect 206 1213 212 1214
rect 326 1218 332 1219
rect 326 1214 327 1218
rect 331 1214 332 1218
rect 326 1213 332 1214
rect 454 1218 460 1219
rect 454 1214 455 1218
rect 459 1214 460 1218
rect 454 1213 460 1214
rect 582 1218 588 1219
rect 582 1214 583 1218
rect 587 1214 588 1218
rect 582 1213 588 1214
rect 718 1218 724 1219
rect 718 1214 719 1218
rect 723 1214 724 1218
rect 718 1213 724 1214
rect 878 1218 884 1219
rect 878 1214 879 1218
rect 883 1214 884 1218
rect 878 1213 884 1214
rect 1054 1218 1060 1219
rect 1054 1214 1055 1218
rect 1059 1214 1060 1218
rect 1054 1213 1060 1214
rect 1262 1218 1268 1219
rect 1262 1214 1263 1218
rect 1267 1214 1268 1218
rect 1262 1213 1268 1214
rect 1486 1218 1492 1219
rect 1486 1214 1487 1218
rect 1491 1214 1492 1218
rect 1486 1213 1492 1214
rect 1718 1218 1724 1219
rect 1718 1214 1719 1218
rect 1723 1214 1724 1218
rect 1718 1213 1724 1214
rect 1934 1218 1940 1219
rect 2030 1218 2036 1219
rect 1934 1214 1935 1218
rect 1939 1214 1940 1218
rect 1934 1213 1940 1214
rect 2110 1194 2116 1195
rect 2110 1190 2111 1194
rect 2115 1190 2116 1194
rect 2070 1189 2076 1190
rect 2110 1189 2116 1190
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2470 1194 2476 1195
rect 2470 1190 2471 1194
rect 2475 1190 2476 1194
rect 2470 1189 2476 1190
rect 2654 1194 2660 1195
rect 2654 1190 2655 1194
rect 2659 1190 2660 1194
rect 2654 1189 2660 1190
rect 2830 1194 2836 1195
rect 2830 1190 2831 1194
rect 2835 1190 2836 1194
rect 2830 1189 2836 1190
rect 2998 1194 3004 1195
rect 2998 1190 2999 1194
rect 3003 1190 3004 1194
rect 2998 1189 3004 1190
rect 3158 1194 3164 1195
rect 3158 1190 3159 1194
rect 3163 1190 3164 1194
rect 3158 1189 3164 1190
rect 3326 1194 3332 1195
rect 3326 1190 3327 1194
rect 3331 1190 3332 1194
rect 3326 1189 3332 1190
rect 3494 1194 3500 1195
rect 3494 1190 3495 1194
rect 3499 1190 3500 1194
rect 3494 1189 3500 1190
rect 3990 1189 3996 1190
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 3990 1185 3991 1189
rect 3995 1185 3996 1189
rect 3990 1184 3996 1185
rect 470 1178 476 1179
rect 470 1174 471 1178
rect 475 1174 476 1178
rect 110 1173 116 1174
rect 470 1173 476 1174
rect 582 1178 588 1179
rect 582 1174 583 1178
rect 587 1174 588 1178
rect 582 1173 588 1174
rect 702 1178 708 1179
rect 702 1174 703 1178
rect 707 1174 708 1178
rect 702 1173 708 1174
rect 822 1178 828 1179
rect 822 1174 823 1178
rect 827 1174 828 1178
rect 822 1173 828 1174
rect 942 1178 948 1179
rect 942 1174 943 1178
rect 947 1174 948 1178
rect 942 1173 948 1174
rect 1062 1178 1068 1179
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1182 1178 1188 1179
rect 1182 1174 1183 1178
rect 1187 1174 1188 1178
rect 1182 1173 1188 1174
rect 1302 1178 1308 1179
rect 1302 1174 1303 1178
rect 1307 1174 1308 1178
rect 1302 1173 1308 1174
rect 1422 1178 1428 1179
rect 1422 1174 1423 1178
rect 1427 1174 1428 1178
rect 1422 1173 1428 1174
rect 1542 1178 1548 1179
rect 1542 1174 1543 1178
rect 1547 1174 1548 1178
rect 1542 1173 1548 1174
rect 2030 1173 2036 1174
rect 110 1169 111 1173
rect 115 1169 116 1173
rect 110 1168 116 1169
rect 2030 1169 2031 1173
rect 2035 1169 2036 1173
rect 2030 1168 2036 1169
rect 2070 1172 2076 1173
rect 2070 1168 2071 1172
rect 2075 1168 2076 1172
rect 2070 1167 2076 1168
rect 3990 1172 3996 1173
rect 3990 1168 3991 1172
rect 3995 1168 3996 1172
rect 3990 1167 3996 1168
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 2030 1156 2036 1157
rect 2030 1152 2031 1156
rect 2035 1152 2036 1156
rect 2030 1151 2036 1152
rect 2110 1153 2116 1154
rect 2110 1149 2111 1153
rect 2115 1149 2116 1153
rect 2110 1148 2116 1149
rect 2278 1153 2284 1154
rect 2278 1149 2279 1153
rect 2283 1149 2284 1153
rect 2278 1148 2284 1149
rect 2470 1153 2476 1154
rect 2470 1149 2471 1153
rect 2475 1149 2476 1153
rect 2470 1148 2476 1149
rect 2654 1153 2660 1154
rect 2654 1149 2655 1153
rect 2659 1149 2660 1153
rect 2654 1148 2660 1149
rect 2830 1153 2836 1154
rect 2830 1149 2831 1153
rect 2835 1149 2836 1153
rect 2830 1148 2836 1149
rect 2998 1153 3004 1154
rect 2998 1149 2999 1153
rect 3003 1149 3004 1153
rect 2998 1148 3004 1149
rect 3158 1153 3164 1154
rect 3158 1149 3159 1153
rect 3163 1149 3164 1153
rect 3158 1148 3164 1149
rect 3326 1153 3332 1154
rect 3326 1149 3327 1153
rect 3331 1149 3332 1153
rect 3326 1148 3332 1149
rect 3494 1153 3500 1154
rect 3494 1149 3495 1153
rect 3499 1149 3500 1153
rect 3494 1148 3500 1149
rect 470 1137 476 1138
rect 470 1133 471 1137
rect 475 1133 476 1137
rect 470 1132 476 1133
rect 582 1137 588 1138
rect 582 1133 583 1137
rect 587 1133 588 1137
rect 582 1132 588 1133
rect 702 1137 708 1138
rect 702 1133 703 1137
rect 707 1133 708 1137
rect 702 1132 708 1133
rect 822 1137 828 1138
rect 822 1133 823 1137
rect 827 1133 828 1137
rect 822 1132 828 1133
rect 942 1137 948 1138
rect 942 1133 943 1137
rect 947 1133 948 1137
rect 942 1132 948 1133
rect 1062 1137 1068 1138
rect 1062 1133 1063 1137
rect 1067 1133 1068 1137
rect 1062 1132 1068 1133
rect 1182 1137 1188 1138
rect 1182 1133 1183 1137
rect 1187 1133 1188 1137
rect 1182 1132 1188 1133
rect 1302 1137 1308 1138
rect 1302 1133 1303 1137
rect 1307 1133 1308 1137
rect 1302 1132 1308 1133
rect 1422 1137 1428 1138
rect 1422 1133 1423 1137
rect 1427 1133 1428 1137
rect 1422 1132 1428 1133
rect 1542 1137 1548 1138
rect 1542 1133 1543 1137
rect 1547 1133 1548 1137
rect 1542 1132 1548 1133
rect 2110 1119 2116 1120
rect 2110 1115 2111 1119
rect 2115 1115 2116 1119
rect 2110 1114 2116 1115
rect 2294 1119 2300 1120
rect 2294 1115 2295 1119
rect 2299 1115 2300 1119
rect 2294 1114 2300 1115
rect 2502 1119 2508 1120
rect 2502 1115 2503 1119
rect 2507 1115 2508 1119
rect 2502 1114 2508 1115
rect 2702 1119 2708 1120
rect 2702 1115 2703 1119
rect 2707 1115 2708 1119
rect 2702 1114 2708 1115
rect 2894 1119 2900 1120
rect 2894 1115 2895 1119
rect 2899 1115 2900 1119
rect 2894 1114 2900 1115
rect 3078 1119 3084 1120
rect 3078 1115 3079 1119
rect 3083 1115 3084 1119
rect 3078 1114 3084 1115
rect 3254 1119 3260 1120
rect 3254 1115 3255 1119
rect 3259 1115 3260 1119
rect 3254 1114 3260 1115
rect 3430 1119 3436 1120
rect 3430 1115 3431 1119
rect 3435 1115 3436 1119
rect 3430 1114 3436 1115
rect 3614 1119 3620 1120
rect 3614 1115 3615 1119
rect 3619 1115 3620 1119
rect 3614 1114 3620 1115
rect 2070 1100 2076 1101
rect 622 1099 628 1100
rect 622 1095 623 1099
rect 627 1095 628 1099
rect 622 1094 628 1095
rect 734 1099 740 1100
rect 734 1095 735 1099
rect 739 1095 740 1099
rect 734 1094 740 1095
rect 854 1099 860 1100
rect 854 1095 855 1099
rect 859 1095 860 1099
rect 854 1094 860 1095
rect 974 1099 980 1100
rect 974 1095 975 1099
rect 979 1095 980 1099
rect 974 1094 980 1095
rect 1094 1099 1100 1100
rect 1094 1095 1095 1099
rect 1099 1095 1100 1099
rect 1094 1094 1100 1095
rect 1214 1099 1220 1100
rect 1214 1095 1215 1099
rect 1219 1095 1220 1099
rect 1214 1094 1220 1095
rect 1334 1099 1340 1100
rect 1334 1095 1335 1099
rect 1339 1095 1340 1099
rect 1334 1094 1340 1095
rect 1454 1099 1460 1100
rect 1454 1095 1455 1099
rect 1459 1095 1460 1099
rect 1454 1094 1460 1095
rect 1574 1099 1580 1100
rect 1574 1095 1575 1099
rect 1579 1095 1580 1099
rect 1574 1094 1580 1095
rect 1702 1099 1708 1100
rect 1702 1095 1703 1099
rect 1707 1095 1708 1099
rect 2070 1096 2071 1100
rect 2075 1096 2076 1100
rect 2070 1095 2076 1096
rect 3990 1100 3996 1101
rect 3990 1096 3991 1100
rect 3995 1096 3996 1100
rect 3990 1095 3996 1096
rect 1702 1094 1708 1095
rect 2070 1083 2076 1084
rect 110 1080 116 1081
rect 110 1076 111 1080
rect 115 1076 116 1080
rect 110 1075 116 1076
rect 2030 1080 2036 1081
rect 2030 1076 2031 1080
rect 2035 1076 2036 1080
rect 2070 1079 2071 1083
rect 2075 1079 2076 1083
rect 3990 1083 3996 1084
rect 3990 1079 3991 1083
rect 3995 1079 3996 1083
rect 2070 1078 2076 1079
rect 2110 1078 2116 1079
rect 2030 1075 2036 1076
rect 2110 1074 2111 1078
rect 2115 1074 2116 1078
rect 2110 1073 2116 1074
rect 2294 1078 2300 1079
rect 2294 1074 2295 1078
rect 2299 1074 2300 1078
rect 2294 1073 2300 1074
rect 2502 1078 2508 1079
rect 2502 1074 2503 1078
rect 2507 1074 2508 1078
rect 2502 1073 2508 1074
rect 2702 1078 2708 1079
rect 2702 1074 2703 1078
rect 2707 1074 2708 1078
rect 2702 1073 2708 1074
rect 2894 1078 2900 1079
rect 2894 1074 2895 1078
rect 2899 1074 2900 1078
rect 2894 1073 2900 1074
rect 3078 1078 3084 1079
rect 3078 1074 3079 1078
rect 3083 1074 3084 1078
rect 3078 1073 3084 1074
rect 3254 1078 3260 1079
rect 3254 1074 3255 1078
rect 3259 1074 3260 1078
rect 3254 1073 3260 1074
rect 3430 1078 3436 1079
rect 3430 1074 3431 1078
rect 3435 1074 3436 1078
rect 3430 1073 3436 1074
rect 3614 1078 3620 1079
rect 3990 1078 3996 1079
rect 3614 1074 3615 1078
rect 3619 1074 3620 1078
rect 3614 1073 3620 1074
rect 110 1063 116 1064
rect 110 1059 111 1063
rect 115 1059 116 1063
rect 2030 1063 2036 1064
rect 2030 1059 2031 1063
rect 2035 1059 2036 1063
rect 110 1058 116 1059
rect 622 1058 628 1059
rect 622 1054 623 1058
rect 627 1054 628 1058
rect 622 1053 628 1054
rect 734 1058 740 1059
rect 734 1054 735 1058
rect 739 1054 740 1058
rect 734 1053 740 1054
rect 854 1058 860 1059
rect 854 1054 855 1058
rect 859 1054 860 1058
rect 854 1053 860 1054
rect 974 1058 980 1059
rect 974 1054 975 1058
rect 979 1054 980 1058
rect 974 1053 980 1054
rect 1094 1058 1100 1059
rect 1094 1054 1095 1058
rect 1099 1054 1100 1058
rect 1094 1053 1100 1054
rect 1214 1058 1220 1059
rect 1214 1054 1215 1058
rect 1219 1054 1220 1058
rect 1214 1053 1220 1054
rect 1334 1058 1340 1059
rect 1334 1054 1335 1058
rect 1339 1054 1340 1058
rect 1334 1053 1340 1054
rect 1454 1058 1460 1059
rect 1454 1054 1455 1058
rect 1459 1054 1460 1058
rect 1454 1053 1460 1054
rect 1574 1058 1580 1059
rect 1574 1054 1575 1058
rect 1579 1054 1580 1058
rect 1574 1053 1580 1054
rect 1702 1058 1708 1059
rect 2030 1058 2036 1059
rect 1702 1054 1703 1058
rect 1707 1054 1708 1058
rect 1702 1053 1708 1054
rect 2166 1038 2172 1039
rect 2166 1034 2167 1038
rect 2171 1034 2172 1038
rect 2070 1033 2076 1034
rect 2166 1033 2172 1034
rect 2286 1038 2292 1039
rect 2286 1034 2287 1038
rect 2291 1034 2292 1038
rect 2286 1033 2292 1034
rect 2422 1038 2428 1039
rect 2422 1034 2423 1038
rect 2427 1034 2428 1038
rect 2422 1033 2428 1034
rect 2574 1038 2580 1039
rect 2574 1034 2575 1038
rect 2579 1034 2580 1038
rect 2574 1033 2580 1034
rect 2742 1038 2748 1039
rect 2742 1034 2743 1038
rect 2747 1034 2748 1038
rect 2742 1033 2748 1034
rect 2918 1038 2924 1039
rect 2918 1034 2919 1038
rect 2923 1034 2924 1038
rect 2918 1033 2924 1034
rect 3094 1038 3100 1039
rect 3094 1034 3095 1038
rect 3099 1034 3100 1038
rect 3094 1033 3100 1034
rect 3278 1038 3284 1039
rect 3278 1034 3279 1038
rect 3283 1034 3284 1038
rect 3278 1033 3284 1034
rect 3462 1038 3468 1039
rect 3462 1034 3463 1038
rect 3467 1034 3468 1038
rect 3462 1033 3468 1034
rect 3654 1038 3660 1039
rect 3654 1034 3655 1038
rect 3659 1034 3660 1038
rect 3654 1033 3660 1034
rect 3990 1033 3996 1034
rect 2070 1029 2071 1033
rect 2075 1029 2076 1033
rect 2070 1028 2076 1029
rect 3990 1029 3991 1033
rect 3995 1029 3996 1033
rect 3990 1028 3996 1029
rect 726 1018 732 1019
rect 726 1014 727 1018
rect 731 1014 732 1018
rect 110 1013 116 1014
rect 726 1013 732 1014
rect 846 1018 852 1019
rect 846 1014 847 1018
rect 851 1014 852 1018
rect 846 1013 852 1014
rect 966 1018 972 1019
rect 966 1014 967 1018
rect 971 1014 972 1018
rect 966 1013 972 1014
rect 1094 1018 1100 1019
rect 1094 1014 1095 1018
rect 1099 1014 1100 1018
rect 1094 1013 1100 1014
rect 1222 1018 1228 1019
rect 1222 1014 1223 1018
rect 1227 1014 1228 1018
rect 1222 1013 1228 1014
rect 1350 1018 1356 1019
rect 1350 1014 1351 1018
rect 1355 1014 1356 1018
rect 1350 1013 1356 1014
rect 1478 1018 1484 1019
rect 1478 1014 1479 1018
rect 1483 1014 1484 1018
rect 1478 1013 1484 1014
rect 1606 1018 1612 1019
rect 1606 1014 1607 1018
rect 1611 1014 1612 1018
rect 1606 1013 1612 1014
rect 1734 1018 1740 1019
rect 1734 1014 1735 1018
rect 1739 1014 1740 1018
rect 1734 1013 1740 1014
rect 1862 1018 1868 1019
rect 1862 1014 1863 1018
rect 1867 1014 1868 1018
rect 2070 1016 2076 1017
rect 1862 1013 1868 1014
rect 2030 1013 2036 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 110 1008 116 1009
rect 2030 1009 2031 1013
rect 2035 1009 2036 1013
rect 2070 1012 2071 1016
rect 2075 1012 2076 1016
rect 2070 1011 2076 1012
rect 3990 1016 3996 1017
rect 3990 1012 3991 1016
rect 3995 1012 3996 1016
rect 3990 1011 3996 1012
rect 2030 1008 2036 1009
rect 2166 997 2172 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 2030 996 2036 997
rect 2030 992 2031 996
rect 2035 992 2036 996
rect 2166 993 2167 997
rect 2171 993 2172 997
rect 2166 992 2172 993
rect 2286 997 2292 998
rect 2286 993 2287 997
rect 2291 993 2292 997
rect 2286 992 2292 993
rect 2422 997 2428 998
rect 2422 993 2423 997
rect 2427 993 2428 997
rect 2422 992 2428 993
rect 2574 997 2580 998
rect 2574 993 2575 997
rect 2579 993 2580 997
rect 2574 992 2580 993
rect 2742 997 2748 998
rect 2742 993 2743 997
rect 2747 993 2748 997
rect 2742 992 2748 993
rect 2918 997 2924 998
rect 2918 993 2919 997
rect 2923 993 2924 997
rect 2918 992 2924 993
rect 3094 997 3100 998
rect 3094 993 3095 997
rect 3099 993 3100 997
rect 3094 992 3100 993
rect 3278 997 3284 998
rect 3278 993 3279 997
rect 3283 993 3284 997
rect 3278 992 3284 993
rect 3462 997 3468 998
rect 3462 993 3463 997
rect 3467 993 3468 997
rect 3462 992 3468 993
rect 3654 997 3660 998
rect 3654 993 3655 997
rect 3659 993 3660 997
rect 3654 992 3660 993
rect 2030 991 2036 992
rect 726 977 732 978
rect 726 973 727 977
rect 731 973 732 977
rect 726 972 732 973
rect 846 977 852 978
rect 846 973 847 977
rect 851 973 852 977
rect 846 972 852 973
rect 966 977 972 978
rect 966 973 967 977
rect 971 973 972 977
rect 966 972 972 973
rect 1094 977 1100 978
rect 1094 973 1095 977
rect 1099 973 1100 977
rect 1094 972 1100 973
rect 1222 977 1228 978
rect 1222 973 1223 977
rect 1227 973 1228 977
rect 1222 972 1228 973
rect 1350 977 1356 978
rect 1350 973 1351 977
rect 1355 973 1356 977
rect 1350 972 1356 973
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1606 977 1612 978
rect 1606 973 1607 977
rect 1611 973 1612 977
rect 1606 972 1612 973
rect 1734 977 1740 978
rect 1734 973 1735 977
rect 1739 973 1740 977
rect 1734 972 1740 973
rect 1862 977 1868 978
rect 1862 973 1863 977
rect 1867 973 1868 977
rect 1862 972 1868 973
rect 2526 959 2532 960
rect 2526 955 2527 959
rect 2531 955 2532 959
rect 2526 954 2532 955
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 2646 954 2652 955
rect 2774 959 2780 960
rect 2774 955 2775 959
rect 2779 955 2780 959
rect 2774 954 2780 955
rect 2918 959 2924 960
rect 2918 955 2919 959
rect 2923 955 2924 959
rect 2918 954 2924 955
rect 3070 959 3076 960
rect 3070 955 3071 959
rect 3075 955 3076 959
rect 3070 954 3076 955
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3398 959 3404 960
rect 3398 955 3399 959
rect 3403 955 3404 959
rect 3398 954 3404 955
rect 3566 959 3572 960
rect 3566 955 3567 959
rect 3571 955 3572 959
rect 3566 954 3572 955
rect 3734 959 3740 960
rect 3734 955 3735 959
rect 3739 955 3740 959
rect 3734 954 3740 955
rect 2070 940 2076 941
rect 590 939 596 940
rect 590 935 591 939
rect 595 935 596 939
rect 590 934 596 935
rect 734 939 740 940
rect 734 935 735 939
rect 739 935 740 939
rect 734 934 740 935
rect 886 939 892 940
rect 886 935 887 939
rect 891 935 892 939
rect 886 934 892 935
rect 1038 939 1044 940
rect 1038 935 1039 939
rect 1043 935 1044 939
rect 1038 934 1044 935
rect 1198 939 1204 940
rect 1198 935 1199 939
rect 1203 935 1204 939
rect 1198 934 1204 935
rect 1350 939 1356 940
rect 1350 935 1351 939
rect 1355 935 1356 939
rect 1350 934 1356 935
rect 1502 939 1508 940
rect 1502 935 1503 939
rect 1507 935 1508 939
rect 1502 934 1508 935
rect 1654 939 1660 940
rect 1654 935 1655 939
rect 1659 935 1660 939
rect 1654 934 1660 935
rect 1806 939 1812 940
rect 1806 935 1807 939
rect 1811 935 1812 939
rect 1806 934 1812 935
rect 1934 939 1940 940
rect 1934 935 1935 939
rect 1939 935 1940 939
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 3990 940 3996 941
rect 3990 936 3991 940
rect 3995 936 3996 940
rect 3990 935 3996 936
rect 1934 934 1940 935
rect 2070 923 2076 924
rect 110 920 116 921
rect 110 916 111 920
rect 115 916 116 920
rect 110 915 116 916
rect 2030 920 2036 921
rect 2030 916 2031 920
rect 2035 916 2036 920
rect 2070 919 2071 923
rect 2075 919 2076 923
rect 3990 923 3996 924
rect 3990 919 3991 923
rect 3995 919 3996 923
rect 2070 918 2076 919
rect 2526 918 2532 919
rect 2030 915 2036 916
rect 2526 914 2527 918
rect 2531 914 2532 918
rect 2526 913 2532 914
rect 2646 918 2652 919
rect 2646 914 2647 918
rect 2651 914 2652 918
rect 2646 913 2652 914
rect 2774 918 2780 919
rect 2774 914 2775 918
rect 2779 914 2780 918
rect 2774 913 2780 914
rect 2918 918 2924 919
rect 2918 914 2919 918
rect 2923 914 2924 918
rect 2918 913 2924 914
rect 3070 918 3076 919
rect 3070 914 3071 918
rect 3075 914 3076 918
rect 3070 913 3076 914
rect 3230 918 3236 919
rect 3230 914 3231 918
rect 3235 914 3236 918
rect 3230 913 3236 914
rect 3398 918 3404 919
rect 3398 914 3399 918
rect 3403 914 3404 918
rect 3398 913 3404 914
rect 3566 918 3572 919
rect 3566 914 3567 918
rect 3571 914 3572 918
rect 3566 913 3572 914
rect 3734 918 3740 919
rect 3990 918 3996 919
rect 3734 914 3735 918
rect 3739 914 3740 918
rect 3734 913 3740 914
rect 110 903 116 904
rect 110 899 111 903
rect 115 899 116 903
rect 2030 903 2036 904
rect 2030 899 2031 903
rect 2035 899 2036 903
rect 110 898 116 899
rect 590 898 596 899
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 734 898 740 899
rect 734 894 735 898
rect 739 894 740 898
rect 734 893 740 894
rect 886 898 892 899
rect 886 894 887 898
rect 891 894 892 898
rect 886 893 892 894
rect 1038 898 1044 899
rect 1038 894 1039 898
rect 1043 894 1044 898
rect 1038 893 1044 894
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1350 898 1356 899
rect 1350 894 1351 898
rect 1355 894 1356 898
rect 1350 893 1356 894
rect 1502 898 1508 899
rect 1502 894 1503 898
rect 1507 894 1508 898
rect 1502 893 1508 894
rect 1654 898 1660 899
rect 1654 894 1655 898
rect 1659 894 1660 898
rect 1654 893 1660 894
rect 1806 898 1812 899
rect 1806 894 1807 898
rect 1811 894 1812 898
rect 1806 893 1812 894
rect 1934 898 1940 899
rect 2030 898 2036 899
rect 1934 894 1935 898
rect 1939 894 1940 898
rect 1934 893 1940 894
rect 2454 874 2460 875
rect 2454 870 2455 874
rect 2459 870 2460 874
rect 2070 869 2076 870
rect 2454 869 2460 870
rect 2574 874 2580 875
rect 2574 870 2575 874
rect 2579 870 2580 874
rect 2574 869 2580 870
rect 2710 874 2716 875
rect 2710 870 2711 874
rect 2715 870 2716 874
rect 2710 869 2716 870
rect 2862 874 2868 875
rect 2862 870 2863 874
rect 2867 870 2868 874
rect 2862 869 2868 870
rect 3014 874 3020 875
rect 3014 870 3015 874
rect 3019 870 3020 874
rect 3014 869 3020 870
rect 3166 874 3172 875
rect 3166 870 3167 874
rect 3171 870 3172 874
rect 3166 869 3172 870
rect 3318 874 3324 875
rect 3318 870 3319 874
rect 3323 870 3324 874
rect 3318 869 3324 870
rect 3470 874 3476 875
rect 3470 870 3471 874
rect 3475 870 3476 874
rect 3470 869 3476 870
rect 3614 874 3620 875
rect 3614 870 3615 874
rect 3619 870 3620 874
rect 3614 869 3620 870
rect 3766 874 3772 875
rect 3766 870 3767 874
rect 3771 870 3772 874
rect 3766 869 3772 870
rect 3894 874 3900 875
rect 3894 870 3895 874
rect 3899 870 3900 874
rect 3894 869 3900 870
rect 3990 869 3996 870
rect 2070 865 2071 869
rect 2075 865 2076 869
rect 2070 864 2076 865
rect 3990 865 3991 869
rect 3995 865 3996 869
rect 3990 864 3996 865
rect 438 858 444 859
rect 438 854 439 858
rect 443 854 444 858
rect 110 853 116 854
rect 438 853 444 854
rect 582 858 588 859
rect 582 854 583 858
rect 587 854 588 858
rect 582 853 588 854
rect 734 858 740 859
rect 734 854 735 858
rect 739 854 740 858
rect 734 853 740 854
rect 886 858 892 859
rect 886 854 887 858
rect 891 854 892 858
rect 886 853 892 854
rect 1046 858 1052 859
rect 1046 854 1047 858
rect 1051 854 1052 858
rect 1046 853 1052 854
rect 1198 858 1204 859
rect 1198 854 1199 858
rect 1203 854 1204 858
rect 1198 853 1204 854
rect 1350 858 1356 859
rect 1350 854 1351 858
rect 1355 854 1356 858
rect 1350 853 1356 854
rect 1494 858 1500 859
rect 1494 854 1495 858
rect 1499 854 1500 858
rect 1494 853 1500 854
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 1646 853 1652 854
rect 1798 858 1804 859
rect 1798 854 1799 858
rect 1803 854 1804 858
rect 1798 853 1804 854
rect 2030 853 2036 854
rect 110 849 111 853
rect 115 849 116 853
rect 110 848 116 849
rect 2030 849 2031 853
rect 2035 849 2036 853
rect 2030 848 2036 849
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2070 847 2076 848
rect 3990 852 3996 853
rect 3990 848 3991 852
rect 3995 848 3996 852
rect 3990 847 3996 848
rect 110 836 116 837
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 2030 836 2036 837
rect 2030 832 2031 836
rect 2035 832 2036 836
rect 2030 831 2036 832
rect 2454 833 2460 834
rect 2454 829 2455 833
rect 2459 829 2460 833
rect 2454 828 2460 829
rect 2574 833 2580 834
rect 2574 829 2575 833
rect 2579 829 2580 833
rect 2574 828 2580 829
rect 2710 833 2716 834
rect 2710 829 2711 833
rect 2715 829 2716 833
rect 2710 828 2716 829
rect 2862 833 2868 834
rect 2862 829 2863 833
rect 2867 829 2868 833
rect 2862 828 2868 829
rect 3014 833 3020 834
rect 3014 829 3015 833
rect 3019 829 3020 833
rect 3014 828 3020 829
rect 3166 833 3172 834
rect 3166 829 3167 833
rect 3171 829 3172 833
rect 3166 828 3172 829
rect 3318 833 3324 834
rect 3318 829 3319 833
rect 3323 829 3324 833
rect 3318 828 3324 829
rect 3470 833 3476 834
rect 3470 829 3471 833
rect 3475 829 3476 833
rect 3470 828 3476 829
rect 3614 833 3620 834
rect 3614 829 3615 833
rect 3619 829 3620 833
rect 3614 828 3620 829
rect 3766 833 3772 834
rect 3766 829 3767 833
rect 3771 829 3772 833
rect 3766 828 3772 829
rect 3894 833 3900 834
rect 3894 829 3895 833
rect 3899 829 3900 833
rect 3894 828 3900 829
rect 438 817 444 818
rect 438 813 439 817
rect 443 813 444 817
rect 438 812 444 813
rect 582 817 588 818
rect 582 813 583 817
rect 587 813 588 817
rect 582 812 588 813
rect 734 817 740 818
rect 734 813 735 817
rect 739 813 740 817
rect 734 812 740 813
rect 886 817 892 818
rect 886 813 887 817
rect 891 813 892 817
rect 886 812 892 813
rect 1046 817 1052 818
rect 1046 813 1047 817
rect 1051 813 1052 817
rect 1046 812 1052 813
rect 1198 817 1204 818
rect 1198 813 1199 817
rect 1203 813 1204 817
rect 1198 812 1204 813
rect 1350 817 1356 818
rect 1350 813 1351 817
rect 1355 813 1356 817
rect 1350 812 1356 813
rect 1494 817 1500 818
rect 1494 813 1495 817
rect 1499 813 1500 817
rect 1494 812 1500 813
rect 1646 817 1652 818
rect 1646 813 1647 817
rect 1651 813 1652 817
rect 1646 812 1652 813
rect 1798 817 1804 818
rect 1798 813 1799 817
rect 1803 813 1804 817
rect 1798 812 1804 813
rect 2214 803 2220 804
rect 2214 799 2215 803
rect 2219 799 2220 803
rect 2214 798 2220 799
rect 2342 803 2348 804
rect 2342 799 2343 803
rect 2347 799 2348 803
rect 2342 798 2348 799
rect 2478 803 2484 804
rect 2478 799 2479 803
rect 2483 799 2484 803
rect 2478 798 2484 799
rect 2622 803 2628 804
rect 2622 799 2623 803
rect 2627 799 2628 803
rect 2622 798 2628 799
rect 2782 803 2788 804
rect 2782 799 2783 803
rect 2787 799 2788 803
rect 2782 798 2788 799
rect 2958 803 2964 804
rect 2958 799 2959 803
rect 2963 799 2964 803
rect 2958 798 2964 799
rect 3166 803 3172 804
rect 3166 799 3167 803
rect 3171 799 3172 803
rect 3166 798 3172 799
rect 3390 803 3396 804
rect 3390 799 3391 803
rect 3395 799 3396 803
rect 3390 798 3396 799
rect 3622 803 3628 804
rect 3622 799 3623 803
rect 3627 799 3628 803
rect 3622 798 3628 799
rect 3862 803 3868 804
rect 3862 799 3863 803
rect 3867 799 3868 803
rect 3862 798 3868 799
rect 278 787 284 788
rect 278 783 279 787
rect 283 783 284 787
rect 278 782 284 783
rect 430 787 436 788
rect 430 783 431 787
rect 435 783 436 787
rect 430 782 436 783
rect 590 787 596 788
rect 590 783 591 787
rect 595 783 596 787
rect 590 782 596 783
rect 750 787 756 788
rect 750 783 751 787
rect 755 783 756 787
rect 750 782 756 783
rect 918 787 924 788
rect 918 783 919 787
rect 923 783 924 787
rect 918 782 924 783
rect 1086 787 1092 788
rect 1086 783 1087 787
rect 1091 783 1092 787
rect 1086 782 1092 783
rect 1254 787 1260 788
rect 1254 783 1255 787
rect 1259 783 1260 787
rect 1254 782 1260 783
rect 1422 787 1428 788
rect 1422 783 1423 787
rect 1427 783 1428 787
rect 1422 782 1428 783
rect 1590 787 1596 788
rect 1590 783 1591 787
rect 1595 783 1596 787
rect 1590 782 1596 783
rect 2070 784 2076 785
rect 2070 780 2071 784
rect 2075 780 2076 784
rect 2070 779 2076 780
rect 3990 784 3996 785
rect 3990 780 3991 784
rect 3995 780 3996 784
rect 3990 779 3996 780
rect 110 768 116 769
rect 110 764 111 768
rect 115 764 116 768
rect 110 763 116 764
rect 2030 768 2036 769
rect 2030 764 2031 768
rect 2035 764 2036 768
rect 2030 763 2036 764
rect 2070 767 2076 768
rect 2070 763 2071 767
rect 2075 763 2076 767
rect 3990 767 3996 768
rect 3990 763 3991 767
rect 3995 763 3996 767
rect 2070 762 2076 763
rect 2214 762 2220 763
rect 2214 758 2215 762
rect 2219 758 2220 762
rect 2214 757 2220 758
rect 2342 762 2348 763
rect 2342 758 2343 762
rect 2347 758 2348 762
rect 2342 757 2348 758
rect 2478 762 2484 763
rect 2478 758 2479 762
rect 2483 758 2484 762
rect 2478 757 2484 758
rect 2622 762 2628 763
rect 2622 758 2623 762
rect 2627 758 2628 762
rect 2622 757 2628 758
rect 2782 762 2788 763
rect 2782 758 2783 762
rect 2787 758 2788 762
rect 2782 757 2788 758
rect 2958 762 2964 763
rect 2958 758 2959 762
rect 2963 758 2964 762
rect 2958 757 2964 758
rect 3166 762 3172 763
rect 3166 758 3167 762
rect 3171 758 3172 762
rect 3166 757 3172 758
rect 3390 762 3396 763
rect 3390 758 3391 762
rect 3395 758 3396 762
rect 3390 757 3396 758
rect 3622 762 3628 763
rect 3622 758 3623 762
rect 3627 758 3628 762
rect 3622 757 3628 758
rect 3862 762 3868 763
rect 3990 762 3996 763
rect 3862 758 3863 762
rect 3867 758 3868 762
rect 3862 757 3868 758
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 2030 751 2036 752
rect 2030 747 2031 751
rect 2035 747 2036 751
rect 110 746 116 747
rect 278 746 284 747
rect 278 742 279 746
rect 283 742 284 746
rect 278 741 284 742
rect 430 746 436 747
rect 430 742 431 746
rect 435 742 436 746
rect 430 741 436 742
rect 590 746 596 747
rect 590 742 591 746
rect 595 742 596 746
rect 590 741 596 742
rect 750 746 756 747
rect 750 742 751 746
rect 755 742 756 746
rect 750 741 756 742
rect 918 746 924 747
rect 918 742 919 746
rect 923 742 924 746
rect 918 741 924 742
rect 1086 746 1092 747
rect 1086 742 1087 746
rect 1091 742 1092 746
rect 1086 741 1092 742
rect 1254 746 1260 747
rect 1254 742 1255 746
rect 1259 742 1260 746
rect 1254 741 1260 742
rect 1422 746 1428 747
rect 1422 742 1423 746
rect 1427 742 1428 746
rect 1422 741 1428 742
rect 1590 746 1596 747
rect 2030 746 2036 747
rect 1590 742 1591 746
rect 1595 742 1596 746
rect 1590 741 1596 742
rect 2110 722 2116 723
rect 2110 718 2111 722
rect 2115 718 2116 722
rect 2070 717 2076 718
rect 2110 717 2116 718
rect 2246 722 2252 723
rect 2246 718 2247 722
rect 2251 718 2252 722
rect 2246 717 2252 718
rect 2422 722 2428 723
rect 2422 718 2423 722
rect 2427 718 2428 722
rect 2422 717 2428 718
rect 2598 722 2604 723
rect 2598 718 2599 722
rect 2603 718 2604 722
rect 2598 717 2604 718
rect 2782 722 2788 723
rect 2782 718 2783 722
rect 2787 718 2788 722
rect 2782 717 2788 718
rect 2966 722 2972 723
rect 2966 718 2967 722
rect 2971 718 2972 722
rect 2966 717 2972 718
rect 3150 722 3156 723
rect 3150 718 3151 722
rect 3155 718 3156 722
rect 3150 717 3156 718
rect 3334 722 3340 723
rect 3334 718 3335 722
rect 3339 718 3340 722
rect 3334 717 3340 718
rect 3518 722 3524 723
rect 3518 718 3519 722
rect 3523 718 3524 722
rect 3518 717 3524 718
rect 3702 722 3708 723
rect 3702 718 3703 722
rect 3707 718 3708 722
rect 3702 717 3708 718
rect 3894 722 3900 723
rect 3894 718 3895 722
rect 3899 718 3900 722
rect 3894 717 3900 718
rect 3990 717 3996 718
rect 2070 713 2071 717
rect 2075 713 2076 717
rect 2070 712 2076 713
rect 3990 713 3991 717
rect 3995 713 3996 717
rect 3990 712 3996 713
rect 150 710 156 711
rect 150 706 151 710
rect 155 706 156 710
rect 110 705 116 706
rect 150 705 156 706
rect 270 710 276 711
rect 270 706 271 710
rect 275 706 276 710
rect 270 705 276 706
rect 422 710 428 711
rect 422 706 423 710
rect 427 706 428 710
rect 422 705 428 706
rect 574 710 580 711
rect 574 706 575 710
rect 579 706 580 710
rect 574 705 580 706
rect 734 710 740 711
rect 734 706 735 710
rect 739 706 740 710
rect 734 705 740 706
rect 886 710 892 711
rect 886 706 887 710
rect 891 706 892 710
rect 886 705 892 706
rect 1038 710 1044 711
rect 1038 706 1039 710
rect 1043 706 1044 710
rect 1038 705 1044 706
rect 1190 710 1196 711
rect 1190 706 1191 710
rect 1195 706 1196 710
rect 1190 705 1196 706
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1494 710 1500 711
rect 1494 706 1495 710
rect 1499 706 1500 710
rect 1494 705 1500 706
rect 2030 705 2036 706
rect 110 701 111 705
rect 115 701 116 705
rect 110 700 116 701
rect 2030 701 2031 705
rect 2035 701 2036 705
rect 2030 700 2036 701
rect 2070 700 2076 701
rect 2070 696 2071 700
rect 2075 696 2076 700
rect 2070 695 2076 696
rect 3990 700 3996 701
rect 3990 696 3991 700
rect 3995 696 3996 700
rect 3990 695 3996 696
rect 110 688 116 689
rect 110 684 111 688
rect 115 684 116 688
rect 110 683 116 684
rect 2030 688 2036 689
rect 2030 684 2031 688
rect 2035 684 2036 688
rect 2030 683 2036 684
rect 2110 681 2116 682
rect 2110 677 2111 681
rect 2115 677 2116 681
rect 2110 676 2116 677
rect 2246 681 2252 682
rect 2246 677 2247 681
rect 2251 677 2252 681
rect 2246 676 2252 677
rect 2422 681 2428 682
rect 2422 677 2423 681
rect 2427 677 2428 681
rect 2422 676 2428 677
rect 2598 681 2604 682
rect 2598 677 2599 681
rect 2603 677 2604 681
rect 2598 676 2604 677
rect 2782 681 2788 682
rect 2782 677 2783 681
rect 2787 677 2788 681
rect 2782 676 2788 677
rect 2966 681 2972 682
rect 2966 677 2967 681
rect 2971 677 2972 681
rect 2966 676 2972 677
rect 3150 681 3156 682
rect 3150 677 3151 681
rect 3155 677 3156 681
rect 3150 676 3156 677
rect 3334 681 3340 682
rect 3334 677 3335 681
rect 3339 677 3340 681
rect 3334 676 3340 677
rect 3518 681 3524 682
rect 3518 677 3519 681
rect 3523 677 3524 681
rect 3518 676 3524 677
rect 3702 681 3708 682
rect 3702 677 3703 681
rect 3707 677 3708 681
rect 3702 676 3708 677
rect 3894 681 3900 682
rect 3894 677 3895 681
rect 3899 677 3900 681
rect 3894 676 3900 677
rect 150 669 156 670
rect 150 665 151 669
rect 155 665 156 669
rect 150 664 156 665
rect 270 669 276 670
rect 270 665 271 669
rect 275 665 276 669
rect 270 664 276 665
rect 422 669 428 670
rect 422 665 423 669
rect 427 665 428 669
rect 422 664 428 665
rect 574 669 580 670
rect 574 665 575 669
rect 579 665 580 669
rect 574 664 580 665
rect 734 669 740 670
rect 734 665 735 669
rect 739 665 740 669
rect 734 664 740 665
rect 886 669 892 670
rect 886 665 887 669
rect 891 665 892 669
rect 886 664 892 665
rect 1038 669 1044 670
rect 1038 665 1039 669
rect 1043 665 1044 669
rect 1038 664 1044 665
rect 1190 669 1196 670
rect 1190 665 1191 669
rect 1195 665 1196 669
rect 1190 664 1196 665
rect 1342 669 1348 670
rect 1342 665 1343 669
rect 1347 665 1348 669
rect 1342 664 1348 665
rect 1494 669 1500 670
rect 1494 665 1495 669
rect 1499 665 1500 669
rect 1494 664 1500 665
rect 2110 647 2116 648
rect 2110 643 2111 647
rect 2115 643 2116 647
rect 2110 642 2116 643
rect 2374 647 2380 648
rect 2374 643 2375 647
rect 2379 643 2380 647
rect 2374 642 2380 643
rect 2654 647 2660 648
rect 2654 643 2655 647
rect 2659 643 2660 647
rect 2654 642 2660 643
rect 2918 647 2924 648
rect 2918 643 2919 647
rect 2923 643 2924 647
rect 2918 642 2924 643
rect 3174 647 3180 648
rect 3174 643 3175 647
rect 3179 643 3180 647
rect 3174 642 3180 643
rect 3422 647 3428 648
rect 3422 643 3423 647
rect 3427 643 3428 647
rect 3422 642 3428 643
rect 3670 647 3676 648
rect 3670 643 3671 647
rect 3675 643 3676 647
rect 3670 642 3676 643
rect 3894 647 3900 648
rect 3894 643 3895 647
rect 3899 643 3900 647
rect 3894 642 3900 643
rect 150 631 156 632
rect 150 627 151 631
rect 155 627 156 631
rect 150 626 156 627
rect 254 631 260 632
rect 254 627 255 631
rect 259 627 260 631
rect 254 626 260 627
rect 390 631 396 632
rect 390 627 391 631
rect 395 627 396 631
rect 390 626 396 627
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 662 631 668 632
rect 662 627 663 631
rect 667 627 668 631
rect 662 626 668 627
rect 806 631 812 632
rect 806 627 807 631
rect 811 627 812 631
rect 806 626 812 627
rect 958 631 964 632
rect 958 627 959 631
rect 963 627 964 631
rect 958 626 964 627
rect 1118 631 1124 632
rect 1118 627 1119 631
rect 1123 627 1124 631
rect 1118 626 1124 627
rect 1286 631 1292 632
rect 1286 627 1287 631
rect 1291 627 1292 631
rect 1286 626 1292 627
rect 1454 631 1460 632
rect 1454 627 1455 631
rect 1459 627 1460 631
rect 1454 626 1460 627
rect 1622 631 1628 632
rect 1622 627 1623 631
rect 1627 627 1628 631
rect 1622 626 1628 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 1934 631 1940 632
rect 1934 627 1935 631
rect 1939 627 1940 631
rect 1934 626 1940 627
rect 2070 628 2076 629
rect 2070 624 2071 628
rect 2075 624 2076 628
rect 2070 623 2076 624
rect 3990 628 3996 629
rect 3990 624 3991 628
rect 3995 624 3996 628
rect 3990 623 3996 624
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 110 607 116 608
rect 2030 612 2036 613
rect 2030 608 2031 612
rect 2035 608 2036 612
rect 2030 607 2036 608
rect 2070 611 2076 612
rect 2070 607 2071 611
rect 2075 607 2076 611
rect 3990 611 3996 612
rect 3990 607 3991 611
rect 3995 607 3996 611
rect 2070 606 2076 607
rect 2110 606 2116 607
rect 2110 602 2111 606
rect 2115 602 2116 606
rect 2110 601 2116 602
rect 2374 606 2380 607
rect 2374 602 2375 606
rect 2379 602 2380 606
rect 2374 601 2380 602
rect 2654 606 2660 607
rect 2654 602 2655 606
rect 2659 602 2660 606
rect 2654 601 2660 602
rect 2918 606 2924 607
rect 2918 602 2919 606
rect 2923 602 2924 606
rect 2918 601 2924 602
rect 3174 606 3180 607
rect 3174 602 3175 606
rect 3179 602 3180 606
rect 3174 601 3180 602
rect 3422 606 3428 607
rect 3422 602 3423 606
rect 3427 602 3428 606
rect 3422 601 3428 602
rect 3670 606 3676 607
rect 3670 602 3671 606
rect 3675 602 3676 606
rect 3670 601 3676 602
rect 3894 606 3900 607
rect 3990 606 3996 607
rect 3894 602 3895 606
rect 3899 602 3900 606
rect 3894 601 3900 602
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 2030 595 2036 596
rect 2030 591 2031 595
rect 2035 591 2036 595
rect 110 590 116 591
rect 150 590 156 591
rect 150 586 151 590
rect 155 586 156 590
rect 150 585 156 586
rect 254 590 260 591
rect 254 586 255 590
rect 259 586 260 590
rect 254 585 260 586
rect 390 590 396 591
rect 390 586 391 590
rect 395 586 396 590
rect 390 585 396 586
rect 526 590 532 591
rect 526 586 527 590
rect 531 586 532 590
rect 526 585 532 586
rect 662 590 668 591
rect 662 586 663 590
rect 667 586 668 590
rect 662 585 668 586
rect 806 590 812 591
rect 806 586 807 590
rect 811 586 812 590
rect 806 585 812 586
rect 958 590 964 591
rect 958 586 959 590
rect 963 586 964 590
rect 958 585 964 586
rect 1118 590 1124 591
rect 1118 586 1119 590
rect 1123 586 1124 590
rect 1118 585 1124 586
rect 1286 590 1292 591
rect 1286 586 1287 590
rect 1291 586 1292 590
rect 1286 585 1292 586
rect 1454 590 1460 591
rect 1454 586 1455 590
rect 1459 586 1460 590
rect 1454 585 1460 586
rect 1622 590 1628 591
rect 1622 586 1623 590
rect 1627 586 1628 590
rect 1622 585 1628 586
rect 1790 590 1796 591
rect 1790 586 1791 590
rect 1795 586 1796 590
rect 1790 585 1796 586
rect 1934 590 1940 591
rect 2030 590 2036 591
rect 1934 586 1935 590
rect 1939 586 1940 590
rect 1934 585 1940 586
rect 2110 562 2116 563
rect 2110 558 2111 562
rect 2115 558 2116 562
rect 2070 557 2076 558
rect 2110 557 2116 558
rect 2214 562 2220 563
rect 2214 558 2215 562
rect 2219 558 2220 562
rect 2214 557 2220 558
rect 2350 562 2356 563
rect 2350 558 2351 562
rect 2355 558 2356 562
rect 2350 557 2356 558
rect 2486 562 2492 563
rect 2486 558 2487 562
rect 2491 558 2492 562
rect 2486 557 2492 558
rect 2630 562 2636 563
rect 2630 558 2631 562
rect 2635 558 2636 562
rect 2630 557 2636 558
rect 2790 562 2796 563
rect 2790 558 2791 562
rect 2795 558 2796 562
rect 2790 557 2796 558
rect 2974 562 2980 563
rect 2974 558 2975 562
rect 2979 558 2980 562
rect 2974 557 2980 558
rect 3190 562 3196 563
rect 3190 558 3191 562
rect 3195 558 3196 562
rect 3190 557 3196 558
rect 3422 562 3428 563
rect 3422 558 3423 562
rect 3427 558 3428 562
rect 3422 557 3428 558
rect 3670 562 3676 563
rect 3670 558 3671 562
rect 3675 558 3676 562
rect 3670 557 3676 558
rect 3894 562 3900 563
rect 3894 558 3895 562
rect 3899 558 3900 562
rect 3894 557 3900 558
rect 3990 557 3996 558
rect 2070 553 2071 557
rect 2075 553 2076 557
rect 2070 552 2076 553
rect 3990 553 3991 557
rect 3995 553 3996 557
rect 3990 552 3996 553
rect 206 546 212 547
rect 206 542 207 546
rect 211 542 212 546
rect 110 541 116 542
rect 206 541 212 542
rect 326 546 332 547
rect 326 542 327 546
rect 331 542 332 546
rect 326 541 332 542
rect 446 546 452 547
rect 446 542 447 546
rect 451 542 452 546
rect 446 541 452 542
rect 566 546 572 547
rect 566 542 567 546
rect 571 542 572 546
rect 566 541 572 542
rect 686 546 692 547
rect 686 542 687 546
rect 691 542 692 546
rect 686 541 692 542
rect 798 546 804 547
rect 798 542 799 546
rect 803 542 804 546
rect 798 541 804 542
rect 910 546 916 547
rect 910 542 911 546
rect 915 542 916 546
rect 910 541 916 542
rect 1030 546 1036 547
rect 1030 542 1031 546
rect 1035 542 1036 546
rect 1030 541 1036 542
rect 1150 546 1156 547
rect 1150 542 1151 546
rect 1155 542 1156 546
rect 1150 541 1156 542
rect 1270 546 1276 547
rect 1270 542 1271 546
rect 1275 542 1276 546
rect 1270 541 1276 542
rect 2030 541 2036 542
rect 110 537 111 541
rect 115 537 116 541
rect 110 536 116 537
rect 2030 537 2031 541
rect 2035 537 2036 541
rect 2030 536 2036 537
rect 2070 540 2076 541
rect 2070 536 2071 540
rect 2075 536 2076 540
rect 2070 535 2076 536
rect 3990 540 3996 541
rect 3990 536 3991 540
rect 3995 536 3996 540
rect 3990 535 3996 536
rect 110 524 116 525
rect 110 520 111 524
rect 115 520 116 524
rect 110 519 116 520
rect 2030 524 2036 525
rect 2030 520 2031 524
rect 2035 520 2036 524
rect 2030 519 2036 520
rect 2110 521 2116 522
rect 2110 517 2111 521
rect 2115 517 2116 521
rect 2110 516 2116 517
rect 2214 521 2220 522
rect 2214 517 2215 521
rect 2219 517 2220 521
rect 2214 516 2220 517
rect 2350 521 2356 522
rect 2350 517 2351 521
rect 2355 517 2356 521
rect 2350 516 2356 517
rect 2486 521 2492 522
rect 2486 517 2487 521
rect 2491 517 2492 521
rect 2486 516 2492 517
rect 2630 521 2636 522
rect 2630 517 2631 521
rect 2635 517 2636 521
rect 2630 516 2636 517
rect 2790 521 2796 522
rect 2790 517 2791 521
rect 2795 517 2796 521
rect 2790 516 2796 517
rect 2974 521 2980 522
rect 2974 517 2975 521
rect 2979 517 2980 521
rect 2974 516 2980 517
rect 3190 521 3196 522
rect 3190 517 3191 521
rect 3195 517 3196 521
rect 3190 516 3196 517
rect 3422 521 3428 522
rect 3422 517 3423 521
rect 3427 517 3428 521
rect 3422 516 3428 517
rect 3670 521 3676 522
rect 3670 517 3671 521
rect 3675 517 3676 521
rect 3670 516 3676 517
rect 3894 521 3900 522
rect 3894 517 3895 521
rect 3899 517 3900 521
rect 3894 516 3900 517
rect 206 505 212 506
rect 206 501 207 505
rect 211 501 212 505
rect 206 500 212 501
rect 326 505 332 506
rect 326 501 327 505
rect 331 501 332 505
rect 326 500 332 501
rect 446 505 452 506
rect 446 501 447 505
rect 451 501 452 505
rect 446 500 452 501
rect 566 505 572 506
rect 566 501 567 505
rect 571 501 572 505
rect 566 500 572 501
rect 686 505 692 506
rect 686 501 687 505
rect 691 501 692 505
rect 686 500 692 501
rect 798 505 804 506
rect 798 501 799 505
rect 803 501 804 505
rect 798 500 804 501
rect 910 505 916 506
rect 910 501 911 505
rect 915 501 916 505
rect 910 500 916 501
rect 1030 505 1036 506
rect 1030 501 1031 505
rect 1035 501 1036 505
rect 1030 500 1036 501
rect 1150 505 1156 506
rect 1150 501 1151 505
rect 1155 501 1156 505
rect 1150 500 1156 501
rect 1270 505 1276 506
rect 1270 501 1271 505
rect 1275 501 1276 505
rect 1270 500 1276 501
rect 2422 487 2428 488
rect 2422 483 2423 487
rect 2427 483 2428 487
rect 2422 482 2428 483
rect 2526 487 2532 488
rect 2526 483 2527 487
rect 2531 483 2532 487
rect 2526 482 2532 483
rect 2630 487 2636 488
rect 2630 483 2631 487
rect 2635 483 2636 487
rect 2630 482 2636 483
rect 2742 487 2748 488
rect 2742 483 2743 487
rect 2747 483 2748 487
rect 2742 482 2748 483
rect 2870 487 2876 488
rect 2870 483 2871 487
rect 2875 483 2876 487
rect 2870 482 2876 483
rect 3030 487 3036 488
rect 3030 483 3031 487
rect 3035 483 3036 487
rect 3030 482 3036 483
rect 3222 487 3228 488
rect 3222 483 3223 487
rect 3227 483 3228 487
rect 3222 482 3228 483
rect 3446 487 3452 488
rect 3446 483 3447 487
rect 3451 483 3452 487
rect 3446 482 3452 483
rect 3678 487 3684 488
rect 3678 483 3679 487
rect 3683 483 3684 487
rect 3678 482 3684 483
rect 3894 487 3900 488
rect 3894 483 3895 487
rect 3899 483 3900 487
rect 3894 482 3900 483
rect 2070 468 2076 469
rect 438 467 444 468
rect 438 463 439 467
rect 443 463 444 467
rect 438 462 444 463
rect 542 467 548 468
rect 542 463 543 467
rect 547 463 548 467
rect 542 462 548 463
rect 646 467 652 468
rect 646 463 647 467
rect 651 463 652 467
rect 646 462 652 463
rect 750 467 756 468
rect 750 463 751 467
rect 755 463 756 467
rect 750 462 756 463
rect 854 467 860 468
rect 854 463 855 467
rect 859 463 860 467
rect 854 462 860 463
rect 958 467 964 468
rect 958 463 959 467
rect 963 463 964 467
rect 958 462 964 463
rect 1062 467 1068 468
rect 1062 463 1063 467
rect 1067 463 1068 467
rect 1062 462 1068 463
rect 1166 467 1172 468
rect 1166 463 1167 467
rect 1171 463 1172 467
rect 1166 462 1172 463
rect 1270 467 1276 468
rect 1270 463 1271 467
rect 1275 463 1276 467
rect 1270 462 1276 463
rect 1374 467 1380 468
rect 1374 463 1375 467
rect 1379 463 1380 467
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 3990 468 3996 469
rect 3990 464 3991 468
rect 3995 464 3996 468
rect 3990 463 3996 464
rect 1374 462 1380 463
rect 2070 451 2076 452
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 110 443 116 444
rect 2030 448 2036 449
rect 2030 444 2031 448
rect 2035 444 2036 448
rect 2070 447 2071 451
rect 2075 447 2076 451
rect 3990 451 3996 452
rect 3990 447 3991 451
rect 3995 447 3996 451
rect 2070 446 2076 447
rect 2422 446 2428 447
rect 2030 443 2036 444
rect 2422 442 2423 446
rect 2427 442 2428 446
rect 2422 441 2428 442
rect 2526 446 2532 447
rect 2526 442 2527 446
rect 2531 442 2532 446
rect 2526 441 2532 442
rect 2630 446 2636 447
rect 2630 442 2631 446
rect 2635 442 2636 446
rect 2630 441 2636 442
rect 2742 446 2748 447
rect 2742 442 2743 446
rect 2747 442 2748 446
rect 2742 441 2748 442
rect 2870 446 2876 447
rect 2870 442 2871 446
rect 2875 442 2876 446
rect 2870 441 2876 442
rect 3030 446 3036 447
rect 3030 442 3031 446
rect 3035 442 3036 446
rect 3030 441 3036 442
rect 3222 446 3228 447
rect 3222 442 3223 446
rect 3227 442 3228 446
rect 3222 441 3228 442
rect 3446 446 3452 447
rect 3446 442 3447 446
rect 3451 442 3452 446
rect 3446 441 3452 442
rect 3678 446 3684 447
rect 3678 442 3679 446
rect 3683 442 3684 446
rect 3678 441 3684 442
rect 3894 446 3900 447
rect 3990 446 3996 447
rect 3894 442 3895 446
rect 3899 442 3900 446
rect 3894 441 3900 442
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 2030 431 2036 432
rect 2030 427 2031 431
rect 2035 427 2036 431
rect 110 426 116 427
rect 438 426 444 427
rect 438 422 439 426
rect 443 422 444 426
rect 438 421 444 422
rect 542 426 548 427
rect 542 422 543 426
rect 547 422 548 426
rect 542 421 548 422
rect 646 426 652 427
rect 646 422 647 426
rect 651 422 652 426
rect 646 421 652 422
rect 750 426 756 427
rect 750 422 751 426
rect 755 422 756 426
rect 750 421 756 422
rect 854 426 860 427
rect 854 422 855 426
rect 859 422 860 426
rect 854 421 860 422
rect 958 426 964 427
rect 958 422 959 426
rect 963 422 964 426
rect 958 421 964 422
rect 1062 426 1068 427
rect 1062 422 1063 426
rect 1067 422 1068 426
rect 1062 421 1068 422
rect 1166 426 1172 427
rect 1166 422 1167 426
rect 1171 422 1172 426
rect 1166 421 1172 422
rect 1270 426 1276 427
rect 1270 422 1271 426
rect 1275 422 1276 426
rect 1270 421 1276 422
rect 1374 426 1380 427
rect 2030 426 2036 427
rect 1374 422 1375 426
rect 1379 422 1380 426
rect 1374 421 1380 422
rect 2526 410 2532 411
rect 2526 406 2527 410
rect 2531 406 2532 410
rect 2070 405 2076 406
rect 2526 405 2532 406
rect 2638 410 2644 411
rect 2638 406 2639 410
rect 2643 406 2644 410
rect 2638 405 2644 406
rect 2774 410 2780 411
rect 2774 406 2775 410
rect 2779 406 2780 410
rect 2774 405 2780 406
rect 2950 410 2956 411
rect 2950 406 2951 410
rect 2955 406 2956 410
rect 2950 405 2956 406
rect 3158 410 3164 411
rect 3158 406 3159 410
rect 3163 406 3164 410
rect 3158 405 3164 406
rect 3398 410 3404 411
rect 3398 406 3399 410
rect 3403 406 3404 410
rect 3398 405 3404 406
rect 3654 410 3660 411
rect 3654 406 3655 410
rect 3659 406 3660 410
rect 3654 405 3660 406
rect 3894 410 3900 411
rect 3894 406 3895 410
rect 3899 406 3900 410
rect 3894 405 3900 406
rect 3990 405 3996 406
rect 2070 401 2071 405
rect 2075 401 2076 405
rect 2070 400 2076 401
rect 3990 401 3991 405
rect 3995 401 3996 405
rect 3990 400 3996 401
rect 2070 388 2076 389
rect 622 386 628 387
rect 622 382 623 386
rect 627 382 628 386
rect 110 381 116 382
rect 622 381 628 382
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 934 386 940 387
rect 934 382 935 386
rect 939 382 940 386
rect 934 381 940 382
rect 1038 386 1044 387
rect 1038 382 1039 386
rect 1043 382 1044 386
rect 1038 381 1044 382
rect 1142 386 1148 387
rect 1142 382 1143 386
rect 1147 382 1148 386
rect 1142 381 1148 382
rect 1246 386 1252 387
rect 1246 382 1247 386
rect 1251 382 1252 386
rect 1246 381 1252 382
rect 1350 386 1356 387
rect 1350 382 1351 386
rect 1355 382 1356 386
rect 1350 381 1356 382
rect 1454 386 1460 387
rect 1454 382 1455 386
rect 1459 382 1460 386
rect 1454 381 1460 382
rect 1558 386 1564 387
rect 1558 382 1559 386
rect 1563 382 1564 386
rect 2070 384 2071 388
rect 2075 384 2076 388
rect 2070 383 2076 384
rect 3990 388 3996 389
rect 3990 384 3991 388
rect 3995 384 3996 388
rect 3990 383 3996 384
rect 1558 381 1564 382
rect 2030 381 2036 382
rect 110 377 111 381
rect 115 377 116 381
rect 110 376 116 377
rect 2030 377 2031 381
rect 2035 377 2036 381
rect 2030 376 2036 377
rect 2526 369 2532 370
rect 2526 365 2527 369
rect 2531 365 2532 369
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 110 359 116 360
rect 2030 364 2036 365
rect 2526 364 2532 365
rect 2638 369 2644 370
rect 2638 365 2639 369
rect 2643 365 2644 369
rect 2638 364 2644 365
rect 2774 369 2780 370
rect 2774 365 2775 369
rect 2779 365 2780 369
rect 2774 364 2780 365
rect 2950 369 2956 370
rect 2950 365 2951 369
rect 2955 365 2956 369
rect 2950 364 2956 365
rect 3158 369 3164 370
rect 3158 365 3159 369
rect 3163 365 3164 369
rect 3158 364 3164 365
rect 3398 369 3404 370
rect 3398 365 3399 369
rect 3403 365 3404 369
rect 3398 364 3404 365
rect 3654 369 3660 370
rect 3654 365 3655 369
rect 3659 365 3660 369
rect 3654 364 3660 365
rect 3894 369 3900 370
rect 3894 365 3895 369
rect 3899 365 3900 369
rect 3894 364 3900 365
rect 2030 360 2031 364
rect 2035 360 2036 364
rect 2030 359 2036 360
rect 622 345 628 346
rect 622 341 623 345
rect 627 341 628 345
rect 622 340 628 341
rect 726 345 732 346
rect 726 341 727 345
rect 731 341 732 345
rect 726 340 732 341
rect 830 345 836 346
rect 830 341 831 345
rect 835 341 836 345
rect 830 340 836 341
rect 934 345 940 346
rect 934 341 935 345
rect 939 341 940 345
rect 934 340 940 341
rect 1038 345 1044 346
rect 1038 341 1039 345
rect 1043 341 1044 345
rect 1038 340 1044 341
rect 1142 345 1148 346
rect 1142 341 1143 345
rect 1147 341 1148 345
rect 1142 340 1148 341
rect 1246 345 1252 346
rect 1246 341 1247 345
rect 1251 341 1252 345
rect 1246 340 1252 341
rect 1350 345 1356 346
rect 1350 341 1351 345
rect 1355 341 1356 345
rect 1350 340 1356 341
rect 1454 345 1460 346
rect 1454 341 1455 345
rect 1459 341 1460 345
rect 1454 340 1460 341
rect 1558 345 1564 346
rect 1558 341 1559 345
rect 1563 341 1564 345
rect 1558 340 1564 341
rect 2270 327 2276 328
rect 2270 323 2271 327
rect 2275 323 2276 327
rect 2270 322 2276 323
rect 2422 327 2428 328
rect 2422 323 2423 327
rect 2427 323 2428 327
rect 2422 322 2428 323
rect 2582 327 2588 328
rect 2582 323 2583 327
rect 2587 323 2588 327
rect 2582 322 2588 323
rect 2742 327 2748 328
rect 2742 323 2743 327
rect 2747 323 2748 327
rect 2742 322 2748 323
rect 2910 327 2916 328
rect 2910 323 2911 327
rect 2915 323 2916 327
rect 2910 322 2916 323
rect 3070 327 3076 328
rect 3070 323 3071 327
rect 3075 323 3076 327
rect 3070 322 3076 323
rect 3222 327 3228 328
rect 3222 323 3223 327
rect 3227 323 3228 327
rect 3222 322 3228 323
rect 3366 327 3372 328
rect 3366 323 3367 327
rect 3371 323 3372 327
rect 3366 322 3372 323
rect 3502 327 3508 328
rect 3502 323 3503 327
rect 3507 323 3508 327
rect 3502 322 3508 323
rect 3638 327 3644 328
rect 3638 323 3639 327
rect 3643 323 3644 327
rect 3638 322 3644 323
rect 3774 327 3780 328
rect 3774 323 3775 327
rect 3779 323 3780 327
rect 3774 322 3780 323
rect 3894 327 3900 328
rect 3894 323 3895 327
rect 3899 323 3900 327
rect 3894 322 3900 323
rect 398 315 404 316
rect 398 311 399 315
rect 403 311 404 315
rect 398 310 404 311
rect 542 315 548 316
rect 542 311 543 315
rect 547 311 548 315
rect 542 310 548 311
rect 686 315 692 316
rect 686 311 687 315
rect 691 311 692 315
rect 686 310 692 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 990 315 996 316
rect 990 311 991 315
rect 995 311 996 315
rect 990 310 996 311
rect 1142 315 1148 316
rect 1142 311 1143 315
rect 1147 311 1148 315
rect 1142 310 1148 311
rect 1302 315 1308 316
rect 1302 311 1303 315
rect 1307 311 1308 315
rect 1302 310 1308 311
rect 1462 315 1468 316
rect 1462 311 1463 315
rect 1467 311 1468 315
rect 1462 310 1468 311
rect 1622 315 1628 316
rect 1622 311 1623 315
rect 1627 311 1628 315
rect 1622 310 1628 311
rect 2070 308 2076 309
rect 2070 304 2071 308
rect 2075 304 2076 308
rect 2070 303 2076 304
rect 3990 308 3996 309
rect 3990 304 3991 308
rect 3995 304 3996 308
rect 3990 303 3996 304
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 2030 296 2036 297
rect 2030 292 2031 296
rect 2035 292 2036 296
rect 2030 291 2036 292
rect 2070 291 2076 292
rect 2070 287 2071 291
rect 2075 287 2076 291
rect 3990 291 3996 292
rect 3990 287 3991 291
rect 3995 287 3996 291
rect 2070 286 2076 287
rect 2270 286 2276 287
rect 2270 282 2271 286
rect 2275 282 2276 286
rect 2270 281 2276 282
rect 2422 286 2428 287
rect 2422 282 2423 286
rect 2427 282 2428 286
rect 2422 281 2428 282
rect 2582 286 2588 287
rect 2582 282 2583 286
rect 2587 282 2588 286
rect 2582 281 2588 282
rect 2742 286 2748 287
rect 2742 282 2743 286
rect 2747 282 2748 286
rect 2742 281 2748 282
rect 2910 286 2916 287
rect 2910 282 2911 286
rect 2915 282 2916 286
rect 2910 281 2916 282
rect 3070 286 3076 287
rect 3070 282 3071 286
rect 3075 282 3076 286
rect 3070 281 3076 282
rect 3222 286 3228 287
rect 3222 282 3223 286
rect 3227 282 3228 286
rect 3222 281 3228 282
rect 3366 286 3372 287
rect 3366 282 3367 286
rect 3371 282 3372 286
rect 3366 281 3372 282
rect 3502 286 3508 287
rect 3502 282 3503 286
rect 3507 282 3508 286
rect 3502 281 3508 282
rect 3638 286 3644 287
rect 3638 282 3639 286
rect 3643 282 3644 286
rect 3638 281 3644 282
rect 3774 286 3780 287
rect 3774 282 3775 286
rect 3779 282 3780 286
rect 3774 281 3780 282
rect 3894 286 3900 287
rect 3990 286 3996 287
rect 3894 282 3895 286
rect 3899 282 3900 286
rect 3894 281 3900 282
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 2030 279 2036 280
rect 2030 275 2031 279
rect 2035 275 2036 279
rect 110 274 116 275
rect 398 274 404 275
rect 398 270 399 274
rect 403 270 404 274
rect 398 269 404 270
rect 542 274 548 275
rect 542 270 543 274
rect 547 270 548 274
rect 542 269 548 270
rect 686 274 692 275
rect 686 270 687 274
rect 691 270 692 274
rect 686 269 692 270
rect 838 274 844 275
rect 838 270 839 274
rect 843 270 844 274
rect 838 269 844 270
rect 990 274 996 275
rect 990 270 991 274
rect 995 270 996 274
rect 990 269 996 270
rect 1142 274 1148 275
rect 1142 270 1143 274
rect 1147 270 1148 274
rect 1142 269 1148 270
rect 1302 274 1308 275
rect 1302 270 1303 274
rect 1307 270 1308 274
rect 1302 269 1308 270
rect 1462 274 1468 275
rect 1462 270 1463 274
rect 1467 270 1468 274
rect 1462 269 1468 270
rect 1622 274 1628 275
rect 2030 274 2036 275
rect 1622 270 1623 274
rect 1627 270 1628 274
rect 1622 269 1628 270
rect 2110 246 2116 247
rect 2110 242 2111 246
rect 2115 242 2116 246
rect 2070 241 2076 242
rect 2110 241 2116 242
rect 2246 246 2252 247
rect 2246 242 2247 246
rect 2251 242 2252 246
rect 2246 241 2252 242
rect 2422 246 2428 247
rect 2422 242 2423 246
rect 2427 242 2428 246
rect 2422 241 2428 242
rect 2598 246 2604 247
rect 2598 242 2599 246
rect 2603 242 2604 246
rect 2598 241 2604 242
rect 2774 246 2780 247
rect 2774 242 2775 246
rect 2779 242 2780 246
rect 2774 241 2780 242
rect 2942 246 2948 247
rect 2942 242 2943 246
rect 2947 242 2948 246
rect 2942 241 2948 242
rect 3102 246 3108 247
rect 3102 242 3103 246
rect 3107 242 3108 246
rect 3102 241 3108 242
rect 3254 246 3260 247
rect 3254 242 3255 246
rect 3259 242 3260 246
rect 3254 241 3260 242
rect 3390 246 3396 247
rect 3390 242 3391 246
rect 3395 242 3396 246
rect 3390 241 3396 242
rect 3526 246 3532 247
rect 3526 242 3527 246
rect 3531 242 3532 246
rect 3526 241 3532 242
rect 3654 246 3660 247
rect 3654 242 3655 246
rect 3659 242 3660 246
rect 3654 241 3660 242
rect 3782 246 3788 247
rect 3782 242 3783 246
rect 3787 242 3788 246
rect 3782 241 3788 242
rect 3894 246 3900 247
rect 3894 242 3895 246
rect 3899 242 3900 246
rect 3894 241 3900 242
rect 3990 241 3996 242
rect 206 238 212 239
rect 206 234 207 238
rect 211 234 212 238
rect 110 233 116 234
rect 206 233 212 234
rect 430 238 436 239
rect 430 234 431 238
rect 435 234 436 238
rect 430 233 436 234
rect 654 238 660 239
rect 654 234 655 238
rect 659 234 660 238
rect 654 233 660 234
rect 870 238 876 239
rect 870 234 871 238
rect 875 234 876 238
rect 870 233 876 234
rect 1070 238 1076 239
rect 1070 234 1071 238
rect 1075 234 1076 238
rect 1070 233 1076 234
rect 1262 238 1268 239
rect 1262 234 1263 238
rect 1267 234 1268 238
rect 1262 233 1268 234
rect 1446 238 1452 239
rect 1446 234 1447 238
rect 1451 234 1452 238
rect 1446 233 1452 234
rect 1630 238 1636 239
rect 1630 234 1631 238
rect 1635 234 1636 238
rect 1630 233 1636 234
rect 1814 238 1820 239
rect 1814 234 1815 238
rect 1819 234 1820 238
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2070 236 2076 237
rect 3990 237 3991 241
rect 3995 237 3996 241
rect 3990 236 3996 237
rect 1814 233 1820 234
rect 2030 233 2036 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 2030 229 2031 233
rect 2035 229 2036 233
rect 2030 228 2036 229
rect 2070 224 2076 225
rect 2070 220 2071 224
rect 2075 220 2076 224
rect 2070 219 2076 220
rect 3990 224 3996 225
rect 3990 220 3991 224
rect 3995 220 3996 224
rect 3990 219 3996 220
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 110 211 116 212
rect 2030 216 2036 217
rect 2030 212 2031 216
rect 2035 212 2036 216
rect 2030 211 2036 212
rect 2110 205 2116 206
rect 2110 201 2111 205
rect 2115 201 2116 205
rect 2110 200 2116 201
rect 2246 205 2252 206
rect 2246 201 2247 205
rect 2251 201 2252 205
rect 2246 200 2252 201
rect 2422 205 2428 206
rect 2422 201 2423 205
rect 2427 201 2428 205
rect 2422 200 2428 201
rect 2598 205 2604 206
rect 2598 201 2599 205
rect 2603 201 2604 205
rect 2598 200 2604 201
rect 2774 205 2780 206
rect 2774 201 2775 205
rect 2779 201 2780 205
rect 2774 200 2780 201
rect 2942 205 2948 206
rect 2942 201 2943 205
rect 2947 201 2948 205
rect 2942 200 2948 201
rect 3102 205 3108 206
rect 3102 201 3103 205
rect 3107 201 3108 205
rect 3102 200 3108 201
rect 3254 205 3260 206
rect 3254 201 3255 205
rect 3259 201 3260 205
rect 3254 200 3260 201
rect 3390 205 3396 206
rect 3390 201 3391 205
rect 3395 201 3396 205
rect 3390 200 3396 201
rect 3526 205 3532 206
rect 3526 201 3527 205
rect 3531 201 3532 205
rect 3526 200 3532 201
rect 3654 205 3660 206
rect 3654 201 3655 205
rect 3659 201 3660 205
rect 3654 200 3660 201
rect 3782 205 3788 206
rect 3782 201 3783 205
rect 3787 201 3788 205
rect 3782 200 3788 201
rect 3894 205 3900 206
rect 3894 201 3895 205
rect 3899 201 3900 205
rect 3894 200 3900 201
rect 206 197 212 198
rect 206 193 207 197
rect 211 193 212 197
rect 206 192 212 193
rect 430 197 436 198
rect 430 193 431 197
rect 435 193 436 197
rect 430 192 436 193
rect 654 197 660 198
rect 654 193 655 197
rect 659 193 660 197
rect 654 192 660 193
rect 870 197 876 198
rect 870 193 871 197
rect 875 193 876 197
rect 870 192 876 193
rect 1070 197 1076 198
rect 1070 193 1071 197
rect 1075 193 1076 197
rect 1070 192 1076 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1446 197 1452 198
rect 1446 193 1447 197
rect 1451 193 1452 197
rect 1446 192 1452 193
rect 1630 197 1636 198
rect 1630 193 1631 197
rect 1635 193 1636 197
rect 1630 192 1636 193
rect 1814 197 1820 198
rect 1814 193 1815 197
rect 1819 193 1820 197
rect 1814 192 1820 193
rect 2110 163 2116 164
rect 2110 159 2111 163
rect 2115 159 2116 163
rect 2110 158 2116 159
rect 2238 163 2244 164
rect 2238 159 2239 163
rect 2243 159 2244 163
rect 2238 158 2244 159
rect 2398 163 2404 164
rect 2398 159 2399 163
rect 2403 159 2404 163
rect 2398 158 2404 159
rect 2566 163 2572 164
rect 2566 159 2567 163
rect 2571 159 2572 163
rect 2566 158 2572 159
rect 2734 163 2740 164
rect 2734 159 2735 163
rect 2739 159 2740 163
rect 2734 158 2740 159
rect 2894 163 2900 164
rect 2894 159 2895 163
rect 2899 159 2900 163
rect 2894 158 2900 159
rect 3046 163 3052 164
rect 3046 159 3047 163
rect 3051 159 3052 163
rect 3046 158 3052 159
rect 3190 163 3196 164
rect 3190 159 3191 163
rect 3195 159 3196 163
rect 3190 158 3196 159
rect 3326 163 3332 164
rect 3326 159 3327 163
rect 3331 159 3332 163
rect 3326 158 3332 159
rect 3454 163 3460 164
rect 3454 159 3455 163
rect 3459 159 3460 163
rect 3454 158 3460 159
rect 3590 163 3596 164
rect 3590 159 3591 163
rect 3595 159 3596 163
rect 3590 158 3596 159
rect 3726 163 3732 164
rect 3726 159 3727 163
rect 3731 159 3732 163
rect 3726 158 3732 159
rect 2070 144 2076 145
rect 2070 140 2071 144
rect 2075 140 2076 144
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 150 134 156 135
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 358 139 364 140
rect 358 135 359 139
rect 363 135 364 139
rect 358 134 364 135
rect 462 139 468 140
rect 462 135 463 139
rect 467 135 468 139
rect 462 134 468 135
rect 566 139 572 140
rect 566 135 567 139
rect 571 135 572 139
rect 566 134 572 135
rect 670 139 676 140
rect 670 135 671 139
rect 675 135 676 139
rect 670 134 676 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 878 139 884 140
rect 878 135 879 139
rect 883 135 884 139
rect 878 134 884 135
rect 982 139 988 140
rect 982 135 983 139
rect 987 135 988 139
rect 982 134 988 135
rect 1086 139 1092 140
rect 1086 135 1087 139
rect 1091 135 1092 139
rect 1086 134 1092 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1294 139 1300 140
rect 1294 135 1295 139
rect 1299 135 1300 139
rect 1294 134 1300 135
rect 1398 139 1404 140
rect 1398 135 1399 139
rect 1403 135 1404 139
rect 1398 134 1404 135
rect 1510 139 1516 140
rect 1510 135 1511 139
rect 1515 135 1516 139
rect 1510 134 1516 135
rect 1622 139 1628 140
rect 1622 135 1623 139
rect 1627 135 1628 139
rect 1622 134 1628 135
rect 1726 139 1732 140
rect 1726 135 1727 139
rect 1731 135 1732 139
rect 1726 134 1732 135
rect 1830 139 1836 140
rect 1830 135 1831 139
rect 1835 135 1836 139
rect 1830 134 1836 135
rect 1934 139 1940 140
rect 2070 139 2076 140
rect 3990 144 3996 145
rect 3990 140 3991 144
rect 3995 140 3996 144
rect 3990 139 3996 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 1934 134 1940 135
rect 2070 127 2076 128
rect 2070 123 2071 127
rect 2075 123 2076 127
rect 3990 127 3996 128
rect 3990 123 3991 127
rect 3995 123 3996 127
rect 2070 122 2076 123
rect 2110 122 2116 123
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2110 118 2111 122
rect 2115 118 2116 122
rect 2110 117 2116 118
rect 2238 122 2244 123
rect 2238 118 2239 122
rect 2243 118 2244 122
rect 2238 117 2244 118
rect 2398 122 2404 123
rect 2398 118 2399 122
rect 2403 118 2404 122
rect 2398 117 2404 118
rect 2566 122 2572 123
rect 2566 118 2567 122
rect 2571 118 2572 122
rect 2566 117 2572 118
rect 2734 122 2740 123
rect 2734 118 2735 122
rect 2739 118 2740 122
rect 2734 117 2740 118
rect 2894 122 2900 123
rect 2894 118 2895 122
rect 2899 118 2900 122
rect 2894 117 2900 118
rect 3046 122 3052 123
rect 3046 118 3047 122
rect 3051 118 3052 122
rect 3046 117 3052 118
rect 3190 122 3196 123
rect 3190 118 3191 122
rect 3195 118 3196 122
rect 3190 117 3196 118
rect 3326 122 3332 123
rect 3326 118 3327 122
rect 3331 118 3332 122
rect 3326 117 3332 118
rect 3454 122 3460 123
rect 3454 118 3455 122
rect 3459 118 3460 122
rect 3454 117 3460 118
rect 3590 122 3596 123
rect 3590 118 3591 122
rect 3595 118 3596 122
rect 3590 117 3596 118
rect 3726 122 3732 123
rect 3990 122 3996 123
rect 3726 118 3727 122
rect 3731 118 3732 122
rect 3726 117 3732 118
rect 2030 115 2036 116
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 2030 103 2036 104
rect 2030 99 2031 103
rect 2035 99 2036 103
rect 110 98 116 99
rect 150 98 156 99
rect 150 94 151 98
rect 155 94 156 98
rect 150 93 156 94
rect 254 98 260 99
rect 254 94 255 98
rect 259 94 260 98
rect 254 93 260 94
rect 358 98 364 99
rect 358 94 359 98
rect 363 94 364 98
rect 358 93 364 94
rect 462 98 468 99
rect 462 94 463 98
rect 467 94 468 98
rect 462 93 468 94
rect 566 98 572 99
rect 566 94 567 98
rect 571 94 572 98
rect 566 93 572 94
rect 670 98 676 99
rect 670 94 671 98
rect 675 94 676 98
rect 670 93 676 94
rect 774 98 780 99
rect 774 94 775 98
rect 779 94 780 98
rect 774 93 780 94
rect 878 98 884 99
rect 878 94 879 98
rect 883 94 884 98
rect 878 93 884 94
rect 982 98 988 99
rect 982 94 983 98
rect 987 94 988 98
rect 982 93 988 94
rect 1086 98 1092 99
rect 1086 94 1087 98
rect 1091 94 1092 98
rect 1086 93 1092 94
rect 1190 98 1196 99
rect 1190 94 1191 98
rect 1195 94 1196 98
rect 1190 93 1196 94
rect 1294 98 1300 99
rect 1294 94 1295 98
rect 1299 94 1300 98
rect 1294 93 1300 94
rect 1398 98 1404 99
rect 1398 94 1399 98
rect 1403 94 1404 98
rect 1398 93 1404 94
rect 1510 98 1516 99
rect 1510 94 1511 98
rect 1515 94 1516 98
rect 1510 93 1516 94
rect 1622 98 1628 99
rect 1622 94 1623 98
rect 1627 94 1628 98
rect 1622 93 1628 94
rect 1726 98 1732 99
rect 1726 94 1727 98
rect 1731 94 1732 98
rect 1726 93 1732 94
rect 1830 98 1836 99
rect 1830 94 1831 98
rect 1835 94 1836 98
rect 1830 93 1836 94
rect 1934 98 1940 99
rect 2030 98 2036 99
rect 1934 94 1935 98
rect 1939 94 1940 98
rect 1934 93 1940 94
<< m3c >>
rect 3399 4063 3403 4067
rect 3503 4063 3507 4067
rect 3607 4063 3611 4067
rect 3711 4063 3715 4067
rect 2071 4044 2075 4048
rect 3991 4044 3995 4048
rect 495 4027 499 4031
rect 599 4027 603 4031
rect 703 4027 707 4031
rect 807 4027 811 4031
rect 911 4027 915 4031
rect 1015 4027 1019 4031
rect 1119 4027 1123 4031
rect 1223 4027 1227 4031
rect 1327 4027 1331 4031
rect 1431 4027 1435 4031
rect 2071 4027 2075 4031
rect 3991 4027 3995 4031
rect 3399 4022 3403 4026
rect 3503 4022 3507 4026
rect 3607 4022 3611 4026
rect 3711 4022 3715 4026
rect 111 4008 115 4012
rect 2031 4008 2035 4012
rect 111 3991 115 3995
rect 2031 3991 2035 3995
rect 495 3986 499 3990
rect 599 3986 603 3990
rect 703 3986 707 3990
rect 807 3986 811 3990
rect 911 3986 915 3990
rect 1015 3986 1019 3990
rect 1119 3986 1123 3990
rect 1223 3986 1227 3990
rect 1327 3986 1331 3990
rect 2111 3990 2115 3994
rect 1431 3986 1435 3990
rect 2215 3990 2219 3994
rect 2319 3990 2323 3994
rect 2423 3990 2427 3994
rect 2527 3990 2531 3994
rect 2647 3990 2651 3994
rect 2775 3990 2779 3994
rect 2903 3990 2907 3994
rect 3031 3990 3035 3994
rect 3159 3990 3163 3994
rect 3287 3990 3291 3994
rect 3415 3990 3419 3994
rect 3551 3990 3555 3994
rect 2071 3985 2075 3989
rect 3991 3985 3995 3989
rect 2071 3968 2075 3972
rect 3991 3968 3995 3972
rect 391 3954 395 3958
rect 495 3954 499 3958
rect 599 3954 603 3958
rect 703 3954 707 3958
rect 807 3954 811 3958
rect 911 3954 915 3958
rect 1015 3954 1019 3958
rect 1119 3954 1123 3958
rect 1223 3954 1227 3958
rect 1327 3954 1331 3958
rect 1431 3954 1435 3958
rect 1535 3954 1539 3958
rect 111 3949 115 3953
rect 2031 3949 2035 3953
rect 2111 3949 2115 3953
rect 2215 3949 2219 3953
rect 2319 3949 2323 3953
rect 2423 3949 2427 3953
rect 2527 3949 2531 3953
rect 2647 3949 2651 3953
rect 2775 3949 2779 3953
rect 2903 3949 2907 3953
rect 3031 3949 3035 3953
rect 3159 3949 3163 3953
rect 3287 3949 3291 3953
rect 3415 3949 3419 3953
rect 3551 3949 3555 3953
rect 111 3932 115 3936
rect 2031 3932 2035 3936
rect 391 3913 395 3917
rect 495 3913 499 3917
rect 599 3913 603 3917
rect 703 3913 707 3917
rect 807 3913 811 3917
rect 911 3913 915 3917
rect 1015 3913 1019 3917
rect 1119 3913 1123 3917
rect 1223 3913 1227 3917
rect 1327 3913 1331 3917
rect 1431 3913 1435 3917
rect 1535 3913 1539 3917
rect 2143 3915 2147 3919
rect 2319 3915 2323 3919
rect 2487 3915 2491 3919
rect 2647 3915 2651 3919
rect 2799 3915 2803 3919
rect 2951 3915 2955 3919
rect 3103 3915 3107 3919
rect 3255 3915 3259 3919
rect 2071 3896 2075 3900
rect 3991 3896 3995 3900
rect 375 3879 379 3883
rect 495 3879 499 3883
rect 623 3879 627 3883
rect 759 3879 763 3883
rect 895 3879 899 3883
rect 1023 3879 1027 3883
rect 1151 3879 1155 3883
rect 1279 3879 1283 3883
rect 1415 3879 1419 3883
rect 1551 3879 1555 3883
rect 2071 3879 2075 3883
rect 3991 3879 3995 3883
rect 2143 3874 2147 3878
rect 2319 3874 2323 3878
rect 2487 3874 2491 3878
rect 2647 3874 2651 3878
rect 2799 3874 2803 3878
rect 2951 3874 2955 3878
rect 3103 3874 3107 3878
rect 3255 3874 3259 3878
rect 111 3860 115 3864
rect 2031 3860 2035 3864
rect 111 3843 115 3847
rect 2031 3843 2035 3847
rect 375 3838 379 3842
rect 495 3838 499 3842
rect 623 3838 627 3842
rect 759 3838 763 3842
rect 895 3838 899 3842
rect 1023 3838 1027 3842
rect 1151 3838 1155 3842
rect 1279 3838 1283 3842
rect 1415 3838 1419 3842
rect 2119 3842 2123 3846
rect 1551 3838 1555 3842
rect 2287 3842 2291 3846
rect 2447 3842 2451 3846
rect 2599 3842 2603 3846
rect 2743 3842 2747 3846
rect 2879 3842 2883 3846
rect 3023 3842 3027 3846
rect 3167 3842 3171 3846
rect 2071 3837 2075 3841
rect 3991 3837 3995 3841
rect 2071 3820 2075 3824
rect 3991 3820 3995 3824
rect 431 3798 435 3802
rect 575 3798 579 3802
rect 719 3798 723 3802
rect 863 3798 867 3802
rect 999 3798 1003 3802
rect 1135 3798 1139 3802
rect 1271 3798 1275 3802
rect 1407 3798 1411 3802
rect 1551 3798 1555 3802
rect 2119 3801 2123 3805
rect 2287 3801 2291 3805
rect 2447 3801 2451 3805
rect 2599 3801 2603 3805
rect 2743 3801 2747 3805
rect 2879 3801 2883 3805
rect 3023 3801 3027 3805
rect 3167 3801 3171 3805
rect 111 3793 115 3797
rect 2031 3793 2035 3797
rect 111 3776 115 3780
rect 2031 3776 2035 3780
rect 2111 3767 2115 3771
rect 2239 3767 2243 3771
rect 2391 3767 2395 3771
rect 2543 3767 2547 3771
rect 2687 3767 2691 3771
rect 2823 3767 2827 3771
rect 2951 3767 2955 3771
rect 3087 3767 3091 3771
rect 3223 3767 3227 3771
rect 431 3757 435 3761
rect 575 3757 579 3761
rect 719 3757 723 3761
rect 863 3757 867 3761
rect 999 3757 1003 3761
rect 1135 3757 1139 3761
rect 1271 3757 1275 3761
rect 1407 3757 1411 3761
rect 1551 3757 1555 3761
rect 2071 3748 2075 3752
rect 3991 3748 3995 3752
rect 2071 3731 2075 3735
rect 3991 3731 3995 3735
rect 2111 3726 2115 3730
rect 2239 3726 2243 3730
rect 2391 3726 2395 3730
rect 2543 3726 2547 3730
rect 2687 3726 2691 3730
rect 2823 3726 2827 3730
rect 2951 3726 2955 3730
rect 3087 3726 3091 3730
rect 3223 3726 3227 3730
rect 359 3719 363 3723
rect 495 3719 499 3723
rect 631 3719 635 3723
rect 775 3719 779 3723
rect 919 3719 923 3723
rect 1071 3719 1075 3723
rect 1223 3719 1227 3723
rect 1375 3719 1379 3723
rect 1527 3719 1531 3723
rect 111 3700 115 3704
rect 2031 3700 2035 3704
rect 111 3683 115 3687
rect 2031 3683 2035 3687
rect 2111 3686 2115 3690
rect 359 3678 363 3682
rect 495 3678 499 3682
rect 631 3678 635 3682
rect 775 3678 779 3682
rect 919 3678 923 3682
rect 1071 3678 1075 3682
rect 1223 3678 1227 3682
rect 1375 3678 1379 3682
rect 2295 3686 2299 3690
rect 2487 3686 2491 3690
rect 2671 3686 2675 3690
rect 2847 3686 2851 3690
rect 3015 3686 3019 3690
rect 3183 3686 3187 3690
rect 3359 3686 3363 3690
rect 1527 3678 1531 3682
rect 2071 3681 2075 3685
rect 3991 3681 3995 3685
rect 2071 3664 2075 3668
rect 3991 3664 3995 3668
rect 343 3646 347 3650
rect 519 3646 523 3650
rect 695 3646 699 3650
rect 863 3646 867 3650
rect 1031 3646 1035 3650
rect 1191 3646 1195 3650
rect 1343 3646 1347 3650
rect 1495 3646 1499 3650
rect 1655 3646 1659 3650
rect 111 3641 115 3645
rect 2031 3641 2035 3645
rect 2111 3645 2115 3649
rect 2295 3645 2299 3649
rect 2487 3645 2491 3649
rect 2671 3645 2675 3649
rect 2847 3645 2851 3649
rect 3015 3645 3019 3649
rect 3183 3645 3187 3649
rect 3359 3645 3363 3649
rect 111 3624 115 3628
rect 2031 3624 2035 3628
rect 343 3605 347 3609
rect 519 3605 523 3609
rect 695 3605 699 3609
rect 863 3605 867 3609
rect 1031 3605 1035 3609
rect 1191 3605 1195 3609
rect 1343 3605 1347 3609
rect 1495 3605 1499 3609
rect 1655 3605 1659 3609
rect 2111 3607 2115 3611
rect 2295 3607 2299 3611
rect 2495 3607 2499 3611
rect 2687 3607 2691 3611
rect 2863 3607 2867 3611
rect 3023 3607 3027 3611
rect 3167 3607 3171 3611
rect 3303 3607 3307 3611
rect 3431 3607 3435 3611
rect 3551 3607 3555 3611
rect 3671 3607 3675 3611
rect 3791 3607 3795 3611
rect 3895 3607 3899 3611
rect 2071 3588 2075 3592
rect 3991 3588 3995 3592
rect 239 3575 243 3579
rect 399 3575 403 3579
rect 551 3575 555 3579
rect 703 3575 707 3579
rect 855 3575 859 3579
rect 999 3575 1003 3579
rect 1135 3575 1139 3579
rect 1263 3575 1267 3579
rect 1383 3575 1387 3579
rect 1495 3575 1499 3579
rect 1607 3575 1611 3579
rect 1719 3575 1723 3579
rect 1831 3575 1835 3579
rect 1935 3575 1939 3579
rect 2071 3571 2075 3575
rect 3991 3571 3995 3575
rect 2111 3566 2115 3570
rect 2295 3566 2299 3570
rect 2495 3566 2499 3570
rect 2687 3566 2691 3570
rect 2863 3566 2867 3570
rect 3023 3566 3027 3570
rect 3167 3566 3171 3570
rect 3303 3566 3307 3570
rect 3431 3566 3435 3570
rect 3551 3566 3555 3570
rect 3671 3566 3675 3570
rect 3791 3566 3795 3570
rect 3895 3566 3899 3570
rect 111 3556 115 3560
rect 2031 3556 2035 3560
rect 111 3539 115 3543
rect 2031 3539 2035 3543
rect 239 3534 243 3538
rect 399 3534 403 3538
rect 551 3534 555 3538
rect 703 3534 707 3538
rect 855 3534 859 3538
rect 999 3534 1003 3538
rect 1135 3534 1139 3538
rect 1263 3534 1267 3538
rect 1383 3534 1387 3538
rect 1495 3534 1499 3538
rect 1607 3534 1611 3538
rect 1719 3534 1723 3538
rect 1831 3534 1835 3538
rect 1935 3534 1939 3538
rect 2447 3522 2451 3526
rect 2591 3522 2595 3526
rect 2727 3522 2731 3526
rect 2863 3522 2867 3526
rect 2991 3522 2995 3526
rect 3119 3522 3123 3526
rect 3239 3522 3243 3526
rect 3351 3522 3355 3526
rect 3463 3522 3467 3526
rect 3575 3522 3579 3526
rect 3687 3522 3691 3526
rect 3791 3522 3795 3526
rect 3895 3522 3899 3526
rect 2071 3517 2075 3521
rect 3991 3517 3995 3521
rect 151 3502 155 3506
rect 375 3502 379 3506
rect 615 3502 619 3506
rect 847 3502 851 3506
rect 1063 3502 1067 3506
rect 1255 3502 1259 3506
rect 1439 3502 1443 3506
rect 1615 3502 1619 3506
rect 1783 3502 1787 3506
rect 1935 3502 1939 3506
rect 111 3497 115 3501
rect 2031 3497 2035 3501
rect 2071 3500 2075 3504
rect 3991 3500 3995 3504
rect 111 3480 115 3484
rect 2031 3480 2035 3484
rect 2447 3481 2451 3485
rect 2591 3481 2595 3485
rect 2727 3481 2731 3485
rect 2863 3481 2867 3485
rect 2991 3481 2995 3485
rect 3119 3481 3123 3485
rect 3239 3481 3243 3485
rect 3351 3481 3355 3485
rect 3463 3481 3467 3485
rect 3575 3481 3579 3485
rect 3687 3481 3691 3485
rect 3791 3481 3795 3485
rect 3895 3481 3899 3485
rect 151 3461 155 3465
rect 375 3461 379 3465
rect 615 3461 619 3465
rect 847 3461 851 3465
rect 1063 3461 1067 3465
rect 1255 3461 1259 3465
rect 1439 3461 1443 3465
rect 1615 3461 1619 3465
rect 1783 3461 1787 3465
rect 1935 3461 1939 3465
rect 2343 3451 2347 3455
rect 2855 3451 2859 3455
rect 3375 3451 3379 3455
rect 3895 3451 3899 3455
rect 2071 3432 2075 3436
rect 3991 3432 3995 3436
rect 2071 3415 2075 3419
rect 3991 3415 3995 3419
rect 151 3407 155 3411
rect 335 3407 339 3411
rect 583 3407 587 3411
rect 863 3407 867 3411
rect 1159 3407 1163 3411
rect 1463 3407 1467 3411
rect 2343 3410 2347 3414
rect 2855 3410 2859 3414
rect 3375 3410 3379 3414
rect 3895 3410 3899 3414
rect 111 3388 115 3392
rect 2031 3388 2035 3392
rect 111 3371 115 3375
rect 2031 3371 2035 3375
rect 2183 3374 2187 3378
rect 151 3366 155 3370
rect 335 3366 339 3370
rect 583 3366 587 3370
rect 863 3366 867 3370
rect 1159 3366 1163 3370
rect 2583 3374 2587 3378
rect 3007 3374 3011 3378
rect 3447 3374 3451 3378
rect 3895 3374 3899 3378
rect 1463 3366 1467 3370
rect 2071 3369 2075 3373
rect 3991 3369 3995 3373
rect 2071 3352 2075 3356
rect 3991 3352 3995 3356
rect 2183 3333 2187 3337
rect 2583 3333 2587 3337
rect 3007 3333 3011 3337
rect 3447 3333 3451 3337
rect 3895 3333 3899 3337
rect 151 3326 155 3330
rect 287 3326 291 3330
rect 463 3326 467 3330
rect 639 3326 643 3330
rect 815 3326 819 3330
rect 991 3326 995 3330
rect 1159 3326 1163 3330
rect 1319 3326 1323 3330
rect 1487 3326 1491 3330
rect 1655 3326 1659 3330
rect 111 3321 115 3325
rect 2031 3321 2035 3325
rect 111 3304 115 3308
rect 2031 3304 2035 3308
rect 151 3285 155 3289
rect 287 3285 291 3289
rect 463 3285 467 3289
rect 639 3285 643 3289
rect 815 3285 819 3289
rect 991 3285 995 3289
rect 1159 3285 1163 3289
rect 1319 3285 1323 3289
rect 1487 3285 1491 3289
rect 1655 3285 1659 3289
rect 2111 3287 2115 3291
rect 2295 3287 2299 3291
rect 2503 3287 2507 3291
rect 2703 3287 2707 3291
rect 2895 3287 2899 3291
rect 3071 3287 3075 3291
rect 3231 3287 3235 3291
rect 3375 3287 3379 3291
rect 3511 3287 3515 3291
rect 3647 3287 3651 3291
rect 3783 3287 3787 3291
rect 3895 3287 3899 3291
rect 2071 3268 2075 3272
rect 3991 3268 3995 3272
rect 2071 3251 2075 3255
rect 3991 3251 3995 3255
rect 151 3243 155 3247
rect 295 3243 299 3247
rect 479 3243 483 3247
rect 671 3243 675 3247
rect 863 3243 867 3247
rect 1055 3243 1059 3247
rect 1247 3243 1251 3247
rect 1431 3243 1435 3247
rect 1615 3243 1619 3247
rect 1807 3243 1811 3247
rect 2111 3246 2115 3250
rect 2295 3246 2299 3250
rect 2503 3246 2507 3250
rect 2703 3246 2707 3250
rect 2895 3246 2899 3250
rect 3071 3246 3075 3250
rect 3231 3246 3235 3250
rect 3375 3246 3379 3250
rect 3511 3246 3515 3250
rect 3647 3246 3651 3250
rect 3783 3246 3787 3250
rect 3895 3246 3899 3250
rect 111 3224 115 3228
rect 2031 3224 2035 3228
rect 2111 3214 2115 3218
rect 2239 3214 2243 3218
rect 2399 3214 2403 3218
rect 2559 3214 2563 3218
rect 2719 3214 2723 3218
rect 2879 3214 2883 3218
rect 3031 3214 3035 3218
rect 3167 3214 3171 3218
rect 3303 3214 3307 3218
rect 3431 3214 3435 3218
rect 3551 3214 3555 3218
rect 3671 3214 3675 3218
rect 3791 3214 3795 3218
rect 3895 3214 3899 3218
rect 111 3207 115 3211
rect 2031 3207 2035 3211
rect 2071 3209 2075 3213
rect 3991 3209 3995 3213
rect 151 3202 155 3206
rect 295 3202 299 3206
rect 479 3202 483 3206
rect 671 3202 675 3206
rect 863 3202 867 3206
rect 1055 3202 1059 3206
rect 1247 3202 1251 3206
rect 1431 3202 1435 3206
rect 1615 3202 1619 3206
rect 1807 3202 1811 3206
rect 2071 3192 2075 3196
rect 3991 3192 3995 3196
rect 2111 3173 2115 3177
rect 2239 3173 2243 3177
rect 2399 3173 2403 3177
rect 2559 3173 2563 3177
rect 2719 3173 2723 3177
rect 2879 3173 2883 3177
rect 3031 3173 3035 3177
rect 3167 3173 3171 3177
rect 3303 3173 3307 3177
rect 3431 3173 3435 3177
rect 3551 3173 3555 3177
rect 3671 3173 3675 3177
rect 3791 3173 3795 3177
rect 3895 3173 3899 3177
rect 287 3158 291 3162
rect 423 3158 427 3162
rect 567 3158 571 3162
rect 727 3158 731 3162
rect 903 3158 907 3162
rect 1095 3158 1099 3162
rect 1295 3158 1299 3162
rect 1495 3158 1499 3162
rect 1703 3158 1707 3162
rect 1919 3158 1923 3162
rect 111 3153 115 3157
rect 2031 3153 2035 3157
rect 111 3136 115 3140
rect 2031 3136 2035 3140
rect 2183 3127 2187 3131
rect 2367 3127 2371 3131
rect 2551 3127 2555 3131
rect 2735 3127 2739 3131
rect 2911 3127 2915 3131
rect 3087 3127 3091 3131
rect 3263 3127 3267 3131
rect 3447 3127 3451 3131
rect 287 3117 291 3121
rect 423 3117 427 3121
rect 567 3117 571 3121
rect 727 3117 731 3121
rect 903 3117 907 3121
rect 1095 3117 1099 3121
rect 1295 3117 1299 3121
rect 1495 3117 1499 3121
rect 1703 3117 1707 3121
rect 1919 3117 1923 3121
rect 2071 3108 2075 3112
rect 3991 3108 3995 3112
rect 2071 3091 2075 3095
rect 3991 3091 3995 3095
rect 2183 3086 2187 3090
rect 2367 3086 2371 3090
rect 2551 3086 2555 3090
rect 2735 3086 2739 3090
rect 2911 3086 2915 3090
rect 3087 3086 3091 3090
rect 3263 3086 3267 3090
rect 3447 3086 3451 3090
rect 575 3071 579 3075
rect 679 3071 683 3075
rect 799 3071 803 3075
rect 935 3071 939 3075
rect 1079 3071 1083 3075
rect 1231 3071 1235 3075
rect 1391 3071 1395 3075
rect 1559 3071 1563 3075
rect 1727 3071 1731 3075
rect 1903 3071 1907 3075
rect 111 3052 115 3056
rect 2031 3052 2035 3056
rect 2351 3046 2355 3050
rect 2455 3046 2459 3050
rect 2567 3046 2571 3050
rect 2687 3046 2691 3050
rect 2807 3046 2811 3050
rect 2927 3046 2931 3050
rect 3047 3046 3051 3050
rect 3167 3046 3171 3050
rect 3295 3046 3299 3050
rect 2071 3041 2075 3045
rect 3991 3041 3995 3045
rect 111 3035 115 3039
rect 2031 3035 2035 3039
rect 575 3030 579 3034
rect 679 3030 683 3034
rect 799 3030 803 3034
rect 935 3030 939 3034
rect 1079 3030 1083 3034
rect 1231 3030 1235 3034
rect 1391 3030 1395 3034
rect 1559 3030 1563 3034
rect 1727 3030 1731 3034
rect 1903 3030 1907 3034
rect 2071 3024 2075 3028
rect 3991 3024 3995 3028
rect 2351 3005 2355 3009
rect 2455 3005 2459 3009
rect 2567 3005 2571 3009
rect 2687 3005 2691 3009
rect 2807 3005 2811 3009
rect 2927 3005 2931 3009
rect 3047 3005 3051 3009
rect 3167 3005 3171 3009
rect 3295 3005 3299 3009
rect 551 2986 555 2990
rect 655 2986 659 2990
rect 759 2986 763 2990
rect 871 2986 875 2990
rect 991 2986 995 2990
rect 1119 2986 1123 2990
rect 1255 2986 1259 2990
rect 1391 2986 1395 2990
rect 1535 2986 1539 2990
rect 1687 2986 1691 2990
rect 111 2981 115 2985
rect 2031 2981 2035 2985
rect 2495 2975 2499 2979
rect 2599 2975 2603 2979
rect 2703 2975 2707 2979
rect 2807 2975 2811 2979
rect 2911 2975 2915 2979
rect 3015 2975 3019 2979
rect 3119 2975 3123 2979
rect 3223 2975 3227 2979
rect 111 2964 115 2968
rect 2031 2964 2035 2968
rect 2071 2956 2075 2960
rect 3991 2956 3995 2960
rect 551 2945 555 2949
rect 655 2945 659 2949
rect 759 2945 763 2949
rect 871 2945 875 2949
rect 991 2945 995 2949
rect 1119 2945 1123 2949
rect 1255 2945 1259 2949
rect 1391 2945 1395 2949
rect 1535 2945 1539 2949
rect 1687 2945 1691 2949
rect 2071 2939 2075 2943
rect 3991 2939 3995 2943
rect 2495 2934 2499 2938
rect 2599 2934 2603 2938
rect 2703 2934 2707 2938
rect 2807 2934 2811 2938
rect 2911 2934 2915 2938
rect 3015 2934 3019 2938
rect 3119 2934 3123 2938
rect 3223 2934 3227 2938
rect 311 2903 315 2907
rect 431 2903 435 2907
rect 559 2903 563 2907
rect 695 2903 699 2907
rect 831 2903 835 2907
rect 975 2903 979 2907
rect 1119 2903 1123 2907
rect 1271 2903 1275 2907
rect 1423 2903 1427 2907
rect 1575 2903 1579 2907
rect 2415 2902 2419 2906
rect 2519 2902 2523 2906
rect 2623 2902 2627 2906
rect 2727 2902 2731 2906
rect 2831 2902 2835 2906
rect 2935 2902 2939 2906
rect 3039 2902 3043 2906
rect 3143 2902 3147 2906
rect 3247 2902 3251 2906
rect 2071 2897 2075 2901
rect 3991 2897 3995 2901
rect 111 2884 115 2888
rect 2031 2884 2035 2888
rect 2071 2880 2075 2884
rect 3991 2880 3995 2884
rect 111 2867 115 2871
rect 2031 2867 2035 2871
rect 311 2862 315 2866
rect 431 2862 435 2866
rect 559 2862 563 2866
rect 695 2862 699 2866
rect 831 2862 835 2866
rect 975 2862 979 2866
rect 1119 2862 1123 2866
rect 1271 2862 1275 2866
rect 1423 2862 1427 2866
rect 1575 2862 1579 2866
rect 2415 2861 2419 2865
rect 2519 2861 2523 2865
rect 2623 2861 2627 2865
rect 2727 2861 2731 2865
rect 2831 2861 2835 2865
rect 2935 2861 2939 2865
rect 3039 2861 3043 2865
rect 3143 2861 3147 2865
rect 3247 2861 3251 2865
rect 2407 2827 2411 2831
rect 2511 2827 2515 2831
rect 2615 2827 2619 2831
rect 2719 2827 2723 2831
rect 2823 2827 2827 2831
rect 2927 2827 2931 2831
rect 3031 2827 3035 2831
rect 3135 2827 3139 2831
rect 3239 2827 3243 2831
rect 151 2814 155 2818
rect 311 2814 315 2818
rect 471 2814 475 2818
rect 623 2814 627 2818
rect 767 2814 771 2818
rect 903 2814 907 2818
rect 1031 2814 1035 2818
rect 1159 2814 1163 2818
rect 1287 2814 1291 2818
rect 1415 2814 1419 2818
rect 111 2809 115 2813
rect 2031 2809 2035 2813
rect 2071 2808 2075 2812
rect 3991 2808 3995 2812
rect 111 2792 115 2796
rect 2031 2792 2035 2796
rect 2071 2791 2075 2795
rect 3991 2791 3995 2795
rect 2407 2786 2411 2790
rect 2511 2786 2515 2790
rect 2615 2786 2619 2790
rect 2719 2786 2723 2790
rect 2823 2786 2827 2790
rect 2927 2786 2931 2790
rect 3031 2786 3035 2790
rect 3135 2786 3139 2790
rect 3239 2786 3243 2790
rect 151 2773 155 2777
rect 311 2773 315 2777
rect 471 2773 475 2777
rect 623 2773 627 2777
rect 767 2773 771 2777
rect 903 2773 907 2777
rect 1031 2773 1035 2777
rect 1159 2773 1163 2777
rect 1287 2773 1291 2777
rect 1415 2773 1419 2777
rect 2303 2746 2307 2750
rect 2415 2746 2419 2750
rect 2535 2746 2539 2750
rect 2655 2746 2659 2750
rect 2775 2746 2779 2750
rect 2895 2746 2899 2750
rect 3015 2746 3019 2750
rect 3143 2746 3147 2750
rect 3271 2746 3275 2750
rect 3399 2746 3403 2750
rect 2071 2741 2075 2745
rect 3991 2741 3995 2745
rect 151 2727 155 2731
rect 303 2727 307 2731
rect 471 2727 475 2731
rect 623 2727 627 2731
rect 767 2727 771 2731
rect 903 2727 907 2731
rect 1039 2727 1043 2731
rect 1167 2727 1171 2731
rect 1295 2727 1299 2731
rect 1423 2727 1427 2731
rect 2071 2724 2075 2728
rect 3991 2724 3995 2728
rect 111 2708 115 2712
rect 2031 2708 2035 2712
rect 2303 2705 2307 2709
rect 2415 2705 2419 2709
rect 2535 2705 2539 2709
rect 2655 2705 2659 2709
rect 2775 2705 2779 2709
rect 2895 2705 2899 2709
rect 3015 2705 3019 2709
rect 3143 2705 3147 2709
rect 3271 2705 3275 2709
rect 3399 2705 3403 2709
rect 111 2691 115 2695
rect 2031 2691 2035 2695
rect 151 2686 155 2690
rect 303 2686 307 2690
rect 471 2686 475 2690
rect 623 2686 627 2690
rect 767 2686 771 2690
rect 903 2686 907 2690
rect 1039 2686 1043 2690
rect 1167 2686 1171 2690
rect 1295 2686 1299 2690
rect 1423 2686 1427 2690
rect 2151 2659 2155 2663
rect 2303 2659 2307 2663
rect 2463 2659 2467 2663
rect 2623 2659 2627 2663
rect 2791 2659 2795 2663
rect 2951 2659 2955 2663
rect 3111 2659 3115 2663
rect 3263 2659 3267 2663
rect 3415 2659 3419 2663
rect 3575 2659 3579 2663
rect 151 2642 155 2646
rect 319 2642 323 2646
rect 511 2642 515 2646
rect 703 2642 707 2646
rect 887 2642 891 2646
rect 1063 2642 1067 2646
rect 1231 2642 1235 2646
rect 1391 2642 1395 2646
rect 1551 2642 1555 2646
rect 1711 2642 1715 2646
rect 111 2637 115 2641
rect 2031 2637 2035 2641
rect 2071 2640 2075 2644
rect 3991 2640 3995 2644
rect 111 2620 115 2624
rect 2031 2620 2035 2624
rect 2071 2623 2075 2627
rect 3991 2623 3995 2627
rect 2151 2618 2155 2622
rect 2303 2618 2307 2622
rect 2463 2618 2467 2622
rect 2623 2618 2627 2622
rect 2791 2618 2795 2622
rect 2951 2618 2955 2622
rect 3111 2618 3115 2622
rect 3263 2618 3267 2622
rect 3415 2618 3419 2622
rect 3575 2618 3579 2622
rect 151 2601 155 2605
rect 319 2601 323 2605
rect 511 2601 515 2605
rect 703 2601 707 2605
rect 887 2601 891 2605
rect 1063 2601 1067 2605
rect 1231 2601 1235 2605
rect 1391 2601 1395 2605
rect 1551 2601 1555 2605
rect 1711 2601 1715 2605
rect 2111 2578 2115 2582
rect 2327 2578 2331 2582
rect 2559 2578 2563 2582
rect 2783 2578 2787 2582
rect 2999 2578 3003 2582
rect 3199 2578 3203 2582
rect 3383 2578 3387 2582
rect 3559 2578 3563 2582
rect 3735 2578 3739 2582
rect 3895 2578 3899 2582
rect 2071 2573 2075 2577
rect 3991 2573 3995 2577
rect 279 2555 283 2559
rect 463 2555 467 2559
rect 663 2555 667 2559
rect 863 2555 867 2559
rect 1063 2555 1067 2559
rect 1255 2555 1259 2559
rect 1431 2555 1435 2559
rect 1607 2555 1611 2559
rect 1783 2555 1787 2559
rect 1935 2555 1939 2559
rect 2071 2556 2075 2560
rect 3991 2556 3995 2560
rect 111 2536 115 2540
rect 2031 2536 2035 2540
rect 2111 2537 2115 2541
rect 2327 2537 2331 2541
rect 2559 2537 2563 2541
rect 2783 2537 2787 2541
rect 2999 2537 3003 2541
rect 3199 2537 3203 2541
rect 3383 2537 3387 2541
rect 3559 2537 3563 2541
rect 3735 2537 3739 2541
rect 3895 2537 3899 2541
rect 111 2519 115 2523
rect 2031 2519 2035 2523
rect 279 2514 283 2518
rect 463 2514 467 2518
rect 663 2514 667 2518
rect 863 2514 867 2518
rect 1063 2514 1067 2518
rect 1255 2514 1259 2518
rect 1431 2514 1435 2518
rect 1607 2514 1611 2518
rect 1783 2514 1787 2518
rect 1935 2514 1939 2518
rect 2111 2507 2115 2511
rect 2255 2507 2259 2511
rect 2439 2507 2443 2511
rect 2631 2507 2635 2511
rect 2823 2507 2827 2511
rect 3007 2507 3011 2511
rect 3175 2507 3179 2511
rect 3335 2507 3339 2511
rect 3487 2507 3491 2511
rect 3631 2507 3635 2511
rect 3775 2507 3779 2511
rect 3895 2507 3899 2511
rect 2071 2488 2075 2492
rect 3991 2488 3995 2492
rect 2071 2471 2075 2475
rect 3991 2471 3995 2475
rect 311 2466 315 2470
rect 471 2466 475 2470
rect 647 2466 651 2470
rect 831 2466 835 2470
rect 1015 2466 1019 2470
rect 1191 2466 1195 2470
rect 1367 2466 1371 2470
rect 1535 2466 1539 2470
rect 1703 2466 1707 2470
rect 1871 2466 1875 2470
rect 2111 2466 2115 2470
rect 2255 2466 2259 2470
rect 2439 2466 2443 2470
rect 2631 2466 2635 2470
rect 2823 2466 2827 2470
rect 3007 2466 3011 2470
rect 3175 2466 3179 2470
rect 3335 2466 3339 2470
rect 3487 2466 3491 2470
rect 3631 2466 3635 2470
rect 3775 2466 3779 2470
rect 3895 2466 3899 2470
rect 111 2461 115 2465
rect 2031 2461 2035 2465
rect 111 2444 115 2448
rect 2031 2444 2035 2448
rect 311 2425 315 2429
rect 471 2425 475 2429
rect 647 2425 651 2429
rect 831 2425 835 2429
rect 1015 2425 1019 2429
rect 1191 2425 1195 2429
rect 1367 2425 1371 2429
rect 1535 2425 1539 2429
rect 1703 2425 1707 2429
rect 1871 2425 1875 2429
rect 2111 2426 2115 2430
rect 2311 2426 2315 2430
rect 2535 2426 2539 2430
rect 2751 2426 2755 2430
rect 2951 2426 2955 2430
rect 3135 2426 3139 2430
rect 3311 2426 3315 2430
rect 3471 2426 3475 2430
rect 3623 2426 3627 2430
rect 3767 2426 3771 2430
rect 3895 2426 3899 2430
rect 2071 2421 2075 2425
rect 3991 2421 3995 2425
rect 2071 2404 2075 2408
rect 3991 2404 3995 2408
rect 207 2383 211 2387
rect 351 2383 355 2387
rect 503 2383 507 2387
rect 655 2383 659 2387
rect 815 2383 819 2387
rect 967 2383 971 2387
rect 1119 2383 1123 2387
rect 1263 2383 1267 2387
rect 1415 2383 1419 2387
rect 1567 2383 1571 2387
rect 2111 2385 2115 2389
rect 2311 2385 2315 2389
rect 2535 2385 2539 2389
rect 2751 2385 2755 2389
rect 2951 2385 2955 2389
rect 3135 2385 3139 2389
rect 3311 2385 3315 2389
rect 3471 2385 3475 2389
rect 3623 2385 3627 2389
rect 3767 2385 3771 2389
rect 3895 2385 3899 2389
rect 111 2364 115 2368
rect 2031 2364 2035 2368
rect 2111 2355 2115 2359
rect 2327 2355 2331 2359
rect 2559 2355 2563 2359
rect 2783 2355 2787 2359
rect 2999 2355 3003 2359
rect 3191 2355 3195 2359
rect 3375 2355 3379 2359
rect 3543 2355 3547 2359
rect 3711 2355 3715 2359
rect 3887 2355 3891 2359
rect 111 2347 115 2351
rect 2031 2347 2035 2351
rect 207 2342 211 2346
rect 351 2342 355 2346
rect 503 2342 507 2346
rect 655 2342 659 2346
rect 815 2342 819 2346
rect 967 2342 971 2346
rect 1119 2342 1123 2346
rect 1263 2342 1267 2346
rect 1415 2342 1419 2346
rect 1567 2342 1571 2346
rect 2071 2336 2075 2340
rect 3991 2336 3995 2340
rect 2071 2319 2075 2323
rect 3991 2319 3995 2323
rect 2111 2314 2115 2318
rect 2327 2314 2331 2318
rect 2559 2314 2563 2318
rect 2783 2314 2787 2318
rect 2999 2314 3003 2318
rect 3191 2314 3195 2318
rect 3375 2314 3379 2318
rect 3543 2314 3547 2318
rect 3711 2314 3715 2318
rect 3887 2314 3891 2318
rect 255 2298 259 2302
rect 359 2298 363 2302
rect 471 2298 475 2302
rect 583 2298 587 2302
rect 695 2298 699 2302
rect 807 2298 811 2302
rect 919 2298 923 2302
rect 1031 2298 1035 2302
rect 1151 2298 1155 2302
rect 1271 2298 1275 2302
rect 111 2293 115 2297
rect 2031 2293 2035 2297
rect 2111 2282 2115 2286
rect 2295 2282 2299 2286
rect 2527 2282 2531 2286
rect 2775 2282 2779 2286
rect 3039 2282 3043 2286
rect 3319 2282 3323 2286
rect 3607 2282 3611 2286
rect 3895 2282 3899 2286
rect 111 2276 115 2280
rect 2031 2276 2035 2280
rect 2071 2277 2075 2281
rect 3991 2277 3995 2281
rect 255 2257 259 2261
rect 359 2257 363 2261
rect 471 2257 475 2261
rect 583 2257 587 2261
rect 695 2257 699 2261
rect 807 2257 811 2261
rect 919 2257 923 2261
rect 1031 2257 1035 2261
rect 1151 2257 1155 2261
rect 1271 2257 1275 2261
rect 2071 2260 2075 2264
rect 3991 2260 3995 2264
rect 2111 2241 2115 2245
rect 2295 2241 2299 2245
rect 2527 2241 2531 2245
rect 2775 2241 2779 2245
rect 3039 2241 3043 2245
rect 3319 2241 3323 2245
rect 3607 2241 3611 2245
rect 3895 2241 3899 2245
rect 183 2215 187 2219
rect 343 2215 347 2219
rect 495 2215 499 2219
rect 647 2215 651 2219
rect 791 2215 795 2219
rect 935 2215 939 2219
rect 1071 2215 1075 2219
rect 1199 2215 1203 2219
rect 1335 2215 1339 2219
rect 1471 2215 1475 2219
rect 2279 2203 2283 2207
rect 2439 2203 2443 2207
rect 2623 2203 2627 2207
rect 2839 2203 2843 2207
rect 3079 2203 3083 2207
rect 3343 2203 3347 2207
rect 3623 2203 3627 2207
rect 3895 2203 3899 2207
rect 111 2196 115 2200
rect 2031 2196 2035 2200
rect 2071 2184 2075 2188
rect 111 2179 115 2183
rect 3991 2184 3995 2188
rect 2031 2179 2035 2183
rect 183 2174 187 2178
rect 343 2174 347 2178
rect 495 2174 499 2178
rect 647 2174 651 2178
rect 791 2174 795 2178
rect 935 2174 939 2178
rect 1071 2174 1075 2178
rect 1199 2174 1203 2178
rect 1335 2174 1339 2178
rect 1471 2174 1475 2178
rect 2071 2167 2075 2171
rect 3991 2167 3995 2171
rect 2279 2162 2283 2166
rect 2439 2162 2443 2166
rect 2623 2162 2627 2166
rect 2839 2162 2843 2166
rect 3079 2162 3083 2166
rect 3343 2162 3347 2166
rect 3623 2162 3627 2166
rect 3895 2162 3899 2166
rect 151 2126 155 2130
rect 327 2126 331 2130
rect 535 2126 539 2130
rect 735 2126 739 2130
rect 927 2126 931 2130
rect 1111 2126 1115 2130
rect 1279 2126 1283 2130
rect 1447 2126 1451 2130
rect 1615 2126 1619 2130
rect 2391 2130 2395 2134
rect 1783 2126 1787 2130
rect 2495 2130 2499 2134
rect 2599 2130 2603 2134
rect 2703 2130 2707 2134
rect 2807 2130 2811 2134
rect 2911 2130 2915 2134
rect 3031 2130 3035 2134
rect 3175 2130 3179 2134
rect 3343 2130 3347 2134
rect 3527 2130 3531 2134
rect 3719 2130 3723 2134
rect 3895 2130 3899 2134
rect 111 2121 115 2125
rect 2031 2121 2035 2125
rect 2071 2125 2075 2129
rect 3991 2125 3995 2129
rect 111 2104 115 2108
rect 2031 2104 2035 2108
rect 2071 2108 2075 2112
rect 3991 2108 3995 2112
rect 151 2085 155 2089
rect 327 2085 331 2089
rect 535 2085 539 2089
rect 735 2085 739 2089
rect 927 2085 931 2089
rect 1111 2085 1115 2089
rect 1279 2085 1283 2089
rect 1447 2085 1451 2089
rect 1615 2085 1619 2089
rect 1783 2085 1787 2089
rect 2391 2089 2395 2093
rect 2495 2089 2499 2093
rect 2599 2089 2603 2093
rect 2703 2089 2707 2093
rect 2807 2089 2811 2093
rect 2911 2089 2915 2093
rect 3031 2089 3035 2093
rect 3175 2089 3179 2093
rect 3343 2089 3347 2093
rect 3527 2089 3531 2093
rect 3719 2089 3723 2093
rect 3895 2089 3899 2093
rect 2487 2055 2491 2059
rect 2591 2055 2595 2059
rect 2695 2055 2699 2059
rect 2807 2055 2811 2059
rect 2935 2055 2939 2059
rect 3095 2055 3099 2059
rect 3279 2055 3283 2059
rect 3479 2055 3483 2059
rect 3695 2055 3699 2059
rect 3895 2055 3899 2059
rect 151 2043 155 2047
rect 383 2043 387 2047
rect 631 2043 635 2047
rect 863 2043 867 2047
rect 1071 2043 1075 2047
rect 1263 2043 1267 2047
rect 1447 2043 1451 2047
rect 1615 2043 1619 2047
rect 1783 2043 1787 2047
rect 1935 2043 1939 2047
rect 2071 2036 2075 2040
rect 3991 2036 3995 2040
rect 111 2024 115 2028
rect 2031 2024 2035 2028
rect 2071 2019 2075 2023
rect 3991 2019 3995 2023
rect 2487 2014 2491 2018
rect 2591 2014 2595 2018
rect 2695 2014 2699 2018
rect 2807 2014 2811 2018
rect 2935 2014 2939 2018
rect 3095 2014 3099 2018
rect 3279 2014 3283 2018
rect 3479 2014 3483 2018
rect 3695 2014 3699 2018
rect 3895 2014 3899 2018
rect 111 2007 115 2011
rect 2031 2007 2035 2011
rect 151 2002 155 2006
rect 383 2002 387 2006
rect 631 2002 635 2006
rect 863 2002 867 2006
rect 1071 2002 1075 2006
rect 1263 2002 1267 2006
rect 1447 2002 1451 2006
rect 1615 2002 1619 2006
rect 1783 2002 1787 2006
rect 1935 2002 1939 2006
rect 2527 1974 2531 1978
rect 2703 1974 2707 1978
rect 2887 1974 2891 1978
rect 3079 1974 3083 1978
rect 3279 1974 3283 1978
rect 3487 1974 3491 1978
rect 3703 1974 3707 1978
rect 3895 1974 3899 1978
rect 2071 1969 2075 1973
rect 3991 1969 3995 1973
rect 151 1958 155 1962
rect 327 1958 331 1962
rect 535 1958 539 1962
rect 735 1958 739 1962
rect 935 1958 939 1962
rect 1127 1958 1131 1962
rect 1303 1958 1307 1962
rect 1471 1958 1475 1962
rect 1631 1958 1635 1962
rect 1791 1958 1795 1962
rect 1935 1958 1939 1962
rect 111 1953 115 1957
rect 2031 1953 2035 1957
rect 2071 1952 2075 1956
rect 3991 1952 3995 1956
rect 111 1936 115 1940
rect 2031 1936 2035 1940
rect 2527 1933 2531 1937
rect 2703 1933 2707 1937
rect 2887 1933 2891 1937
rect 3079 1933 3083 1937
rect 3279 1933 3283 1937
rect 3487 1933 3491 1937
rect 3703 1933 3707 1937
rect 3895 1933 3899 1937
rect 151 1917 155 1921
rect 327 1917 331 1921
rect 535 1917 539 1921
rect 735 1917 739 1921
rect 935 1917 939 1921
rect 1127 1917 1131 1921
rect 1303 1917 1307 1921
rect 1471 1917 1475 1921
rect 1631 1917 1635 1921
rect 1791 1917 1795 1921
rect 1935 1917 1939 1921
rect 2111 1899 2115 1903
rect 2303 1899 2307 1903
rect 2519 1899 2523 1903
rect 2735 1899 2739 1903
rect 2959 1899 2963 1903
rect 3191 1899 3195 1903
rect 3431 1899 3435 1903
rect 3671 1899 3675 1903
rect 3895 1899 3899 1903
rect 151 1883 155 1887
rect 303 1883 307 1887
rect 463 1883 467 1887
rect 615 1883 619 1887
rect 767 1883 771 1887
rect 927 1883 931 1887
rect 1103 1883 1107 1887
rect 1295 1883 1299 1887
rect 1511 1883 1515 1887
rect 1735 1883 1739 1887
rect 1935 1883 1939 1887
rect 2071 1880 2075 1884
rect 3991 1880 3995 1884
rect 111 1864 115 1868
rect 2031 1864 2035 1868
rect 2071 1863 2075 1867
rect 3991 1863 3995 1867
rect 2111 1858 2115 1862
rect 2303 1858 2307 1862
rect 2519 1858 2523 1862
rect 2735 1858 2739 1862
rect 2959 1858 2963 1862
rect 3191 1858 3195 1862
rect 3431 1858 3435 1862
rect 3671 1858 3675 1862
rect 3895 1858 3899 1862
rect 111 1847 115 1851
rect 2031 1847 2035 1851
rect 151 1842 155 1846
rect 303 1842 307 1846
rect 463 1842 467 1846
rect 615 1842 619 1846
rect 767 1842 771 1846
rect 927 1842 931 1846
rect 1103 1842 1107 1846
rect 1295 1842 1299 1846
rect 1511 1842 1515 1846
rect 1735 1842 1739 1846
rect 1935 1842 1939 1846
rect 2111 1826 2115 1830
rect 2231 1826 2235 1830
rect 2399 1826 2403 1830
rect 2599 1826 2603 1830
rect 2831 1826 2835 1830
rect 3079 1826 3083 1830
rect 3351 1826 3355 1830
rect 3631 1826 3635 1830
rect 3895 1826 3899 1830
rect 2071 1821 2075 1825
rect 3991 1821 3995 1825
rect 2071 1804 2075 1808
rect 3991 1804 3995 1808
rect 151 1798 155 1802
rect 343 1798 347 1802
rect 543 1798 547 1802
rect 735 1798 739 1802
rect 919 1798 923 1802
rect 1095 1798 1099 1802
rect 1271 1798 1275 1802
rect 1447 1798 1451 1802
rect 1623 1798 1627 1802
rect 1807 1798 1811 1802
rect 111 1793 115 1797
rect 2031 1793 2035 1797
rect 2111 1785 2115 1789
rect 2231 1785 2235 1789
rect 2399 1785 2403 1789
rect 2599 1785 2603 1789
rect 2831 1785 2835 1789
rect 3079 1785 3083 1789
rect 3351 1785 3355 1789
rect 3631 1785 3635 1789
rect 3895 1785 3899 1789
rect 111 1776 115 1780
rect 2031 1776 2035 1780
rect 151 1757 155 1761
rect 343 1757 347 1761
rect 543 1757 547 1761
rect 735 1757 739 1761
rect 919 1757 923 1761
rect 1095 1757 1099 1761
rect 1271 1757 1275 1761
rect 1447 1757 1451 1761
rect 1623 1757 1627 1761
rect 1807 1757 1811 1761
rect 2111 1751 2115 1755
rect 2239 1751 2243 1755
rect 2399 1751 2403 1755
rect 2575 1751 2579 1755
rect 2751 1751 2755 1755
rect 2935 1751 2939 1755
rect 3127 1751 3131 1755
rect 3319 1751 3323 1755
rect 3511 1751 3515 1755
rect 3711 1751 3715 1755
rect 3895 1751 3899 1755
rect 2071 1732 2075 1736
rect 3991 1732 3995 1736
rect 151 1723 155 1727
rect 319 1723 323 1727
rect 527 1723 531 1727
rect 743 1723 747 1727
rect 959 1723 963 1727
rect 1167 1723 1171 1727
rect 1367 1723 1371 1727
rect 1559 1723 1563 1727
rect 1759 1723 1763 1727
rect 1935 1723 1939 1727
rect 2071 1715 2075 1719
rect 3991 1715 3995 1719
rect 2111 1710 2115 1714
rect 2239 1710 2243 1714
rect 2399 1710 2403 1714
rect 2575 1710 2579 1714
rect 2751 1710 2755 1714
rect 2935 1710 2939 1714
rect 3127 1710 3131 1714
rect 3319 1710 3323 1714
rect 3511 1710 3515 1714
rect 3711 1710 3715 1714
rect 3895 1710 3899 1714
rect 111 1704 115 1708
rect 2031 1704 2035 1708
rect 111 1687 115 1691
rect 2031 1687 2035 1691
rect 151 1682 155 1686
rect 319 1682 323 1686
rect 527 1682 531 1686
rect 743 1682 747 1686
rect 959 1682 963 1686
rect 1167 1682 1171 1686
rect 1367 1682 1371 1686
rect 1559 1682 1563 1686
rect 1759 1682 1763 1686
rect 1935 1682 1939 1686
rect 2111 1670 2115 1674
rect 2311 1670 2315 1674
rect 2527 1670 2531 1674
rect 2743 1670 2747 1674
rect 2951 1670 2955 1674
rect 3151 1670 3155 1674
rect 3343 1670 3347 1674
rect 3527 1670 3531 1674
rect 3719 1670 3723 1674
rect 3895 1670 3899 1674
rect 2071 1665 2075 1669
rect 3991 1665 3995 1669
rect 151 1650 155 1654
rect 319 1650 323 1654
rect 503 1650 507 1654
rect 695 1650 699 1654
rect 887 1650 891 1654
rect 1079 1650 1083 1654
rect 1263 1650 1267 1654
rect 1439 1650 1443 1654
rect 1615 1650 1619 1654
rect 1791 1650 1795 1654
rect 111 1645 115 1649
rect 2031 1645 2035 1649
rect 2071 1648 2075 1652
rect 3991 1648 3995 1652
rect 111 1628 115 1632
rect 2031 1628 2035 1632
rect 2111 1629 2115 1633
rect 2311 1629 2315 1633
rect 2527 1629 2531 1633
rect 2743 1629 2747 1633
rect 2951 1629 2955 1633
rect 3151 1629 3155 1633
rect 3343 1629 3347 1633
rect 3527 1629 3531 1633
rect 3719 1629 3723 1633
rect 3895 1629 3899 1633
rect 151 1609 155 1613
rect 319 1609 323 1613
rect 503 1609 507 1613
rect 695 1609 699 1613
rect 887 1609 891 1613
rect 1079 1609 1083 1613
rect 1263 1609 1267 1613
rect 1439 1609 1443 1613
rect 1615 1609 1619 1613
rect 1791 1609 1795 1613
rect 2479 1587 2483 1591
rect 2583 1587 2587 1591
rect 2695 1587 2699 1591
rect 2815 1587 2819 1591
rect 2943 1587 2947 1591
rect 3079 1587 3083 1591
rect 3223 1587 3227 1591
rect 3383 1587 3387 1591
rect 3551 1587 3555 1591
rect 3727 1587 3731 1591
rect 3895 1587 3899 1591
rect 319 1571 323 1575
rect 455 1571 459 1575
rect 599 1571 603 1575
rect 743 1571 747 1575
rect 887 1571 891 1575
rect 1031 1571 1035 1575
rect 1175 1571 1179 1575
rect 1319 1571 1323 1575
rect 1471 1571 1475 1575
rect 1623 1571 1627 1575
rect 2071 1568 2075 1572
rect 3991 1568 3995 1572
rect 111 1552 115 1556
rect 2031 1552 2035 1556
rect 2071 1551 2075 1555
rect 3991 1551 3995 1555
rect 2479 1546 2483 1550
rect 2583 1546 2587 1550
rect 2695 1546 2699 1550
rect 2815 1546 2819 1550
rect 2943 1546 2947 1550
rect 3079 1546 3083 1550
rect 3223 1546 3227 1550
rect 3383 1546 3387 1550
rect 3551 1546 3555 1550
rect 3727 1546 3731 1550
rect 3895 1546 3899 1550
rect 111 1535 115 1539
rect 2031 1535 2035 1539
rect 319 1530 323 1534
rect 455 1530 459 1534
rect 599 1530 603 1534
rect 743 1530 747 1534
rect 887 1530 891 1534
rect 1031 1530 1035 1534
rect 1175 1530 1179 1534
rect 1319 1530 1323 1534
rect 1471 1530 1475 1534
rect 1623 1530 1627 1534
rect 2487 1502 2491 1506
rect 2591 1502 2595 1506
rect 2695 1502 2699 1506
rect 2807 1502 2811 1506
rect 2935 1502 2939 1506
rect 3071 1502 3075 1506
rect 3223 1502 3227 1506
rect 3383 1502 3387 1506
rect 3551 1502 3555 1506
rect 3719 1502 3723 1506
rect 3895 1502 3899 1506
rect 2071 1497 2075 1501
rect 3991 1497 3995 1501
rect 359 1490 363 1494
rect 487 1490 491 1494
rect 623 1490 627 1494
rect 775 1490 779 1494
rect 927 1490 931 1494
rect 1087 1490 1091 1494
rect 1255 1490 1259 1494
rect 1423 1490 1427 1494
rect 1591 1490 1595 1494
rect 1767 1490 1771 1494
rect 111 1485 115 1489
rect 2031 1485 2035 1489
rect 2071 1480 2075 1484
rect 3991 1480 3995 1484
rect 111 1468 115 1472
rect 2031 1468 2035 1472
rect 2487 1461 2491 1465
rect 2591 1461 2595 1465
rect 2695 1461 2699 1465
rect 2807 1461 2811 1465
rect 2935 1461 2939 1465
rect 3071 1461 3075 1465
rect 3223 1461 3227 1465
rect 3383 1461 3387 1465
rect 3551 1461 3555 1465
rect 3719 1461 3723 1465
rect 3895 1461 3899 1465
rect 359 1449 363 1453
rect 487 1449 491 1453
rect 623 1449 627 1453
rect 775 1449 779 1453
rect 927 1449 931 1453
rect 1087 1449 1091 1453
rect 1255 1449 1259 1453
rect 1423 1449 1427 1453
rect 1591 1449 1595 1453
rect 1767 1449 1771 1453
rect 2239 1427 2243 1431
rect 2351 1427 2355 1431
rect 2471 1427 2475 1431
rect 2591 1427 2595 1431
rect 2727 1427 2731 1431
rect 2879 1427 2883 1431
rect 3055 1427 3059 1431
rect 3247 1427 3251 1431
rect 3455 1427 3459 1431
rect 3671 1427 3675 1431
rect 3887 1427 3891 1431
rect 151 1411 155 1415
rect 271 1411 275 1415
rect 431 1411 435 1415
rect 615 1411 619 1415
rect 807 1411 811 1415
rect 1007 1411 1011 1415
rect 1215 1411 1219 1415
rect 1423 1411 1427 1415
rect 1631 1411 1635 1415
rect 1847 1411 1851 1415
rect 2071 1408 2075 1412
rect 3991 1408 3995 1412
rect 111 1392 115 1396
rect 2031 1392 2035 1396
rect 2071 1391 2075 1395
rect 3991 1391 3995 1395
rect 2239 1386 2243 1390
rect 2351 1386 2355 1390
rect 2471 1386 2475 1390
rect 2591 1386 2595 1390
rect 2727 1386 2731 1390
rect 2879 1386 2883 1390
rect 3055 1386 3059 1390
rect 3247 1386 3251 1390
rect 3455 1386 3459 1390
rect 3671 1386 3675 1390
rect 3887 1386 3891 1390
rect 111 1375 115 1379
rect 2031 1375 2035 1379
rect 151 1370 155 1374
rect 271 1370 275 1374
rect 431 1370 435 1374
rect 615 1370 619 1374
rect 807 1370 811 1374
rect 1007 1370 1011 1374
rect 1215 1370 1219 1374
rect 1423 1370 1427 1374
rect 1631 1370 1635 1374
rect 1847 1370 1851 1374
rect 2391 1346 2395 1350
rect 2527 1346 2531 1350
rect 2679 1346 2683 1350
rect 2839 1346 2843 1350
rect 2999 1346 3003 1350
rect 3167 1346 3171 1350
rect 3343 1346 3347 1350
rect 3519 1346 3523 1350
rect 3695 1346 3699 1350
rect 3879 1346 3883 1350
rect 2071 1341 2075 1345
rect 3991 1341 3995 1345
rect 151 1326 155 1330
rect 287 1326 291 1330
rect 463 1326 467 1330
rect 663 1326 667 1330
rect 863 1326 867 1330
rect 1063 1326 1067 1330
rect 1255 1326 1259 1330
rect 1431 1326 1435 1330
rect 1607 1326 1611 1330
rect 1783 1326 1787 1330
rect 1935 1326 1939 1330
rect 111 1321 115 1325
rect 2031 1321 2035 1325
rect 2071 1324 2075 1328
rect 3991 1324 3995 1328
rect 111 1304 115 1308
rect 2031 1304 2035 1308
rect 2391 1305 2395 1309
rect 2527 1305 2531 1309
rect 2679 1305 2683 1309
rect 2839 1305 2843 1309
rect 2999 1305 3003 1309
rect 3167 1305 3171 1309
rect 3343 1305 3347 1309
rect 3519 1305 3523 1309
rect 3695 1305 3699 1309
rect 3879 1305 3883 1309
rect 151 1285 155 1289
rect 287 1285 291 1289
rect 463 1285 467 1289
rect 663 1285 667 1289
rect 863 1285 867 1289
rect 1063 1285 1067 1289
rect 1255 1285 1259 1289
rect 1431 1285 1435 1289
rect 1607 1285 1611 1289
rect 1783 1285 1787 1289
rect 1935 1285 1939 1289
rect 2111 1267 2115 1271
rect 2343 1267 2347 1271
rect 2583 1267 2587 1271
rect 2799 1267 2803 1271
rect 2999 1267 3003 1271
rect 3183 1267 3187 1271
rect 3343 1267 3347 1271
rect 3495 1267 3499 1271
rect 3639 1267 3643 1271
rect 3775 1267 3779 1271
rect 3895 1267 3899 1271
rect 207 1255 211 1259
rect 327 1255 331 1259
rect 455 1255 459 1259
rect 583 1255 587 1259
rect 719 1255 723 1259
rect 879 1255 883 1259
rect 1055 1255 1059 1259
rect 1263 1255 1267 1259
rect 1487 1255 1491 1259
rect 1719 1255 1723 1259
rect 1935 1255 1939 1259
rect 2071 1248 2075 1252
rect 3991 1248 3995 1252
rect 111 1236 115 1240
rect 2031 1236 2035 1240
rect 2071 1231 2075 1235
rect 3991 1231 3995 1235
rect 2111 1226 2115 1230
rect 2343 1226 2347 1230
rect 2583 1226 2587 1230
rect 2799 1226 2803 1230
rect 2999 1226 3003 1230
rect 3183 1226 3187 1230
rect 3343 1226 3347 1230
rect 3495 1226 3499 1230
rect 3639 1226 3643 1230
rect 3775 1226 3779 1230
rect 3895 1226 3899 1230
rect 111 1219 115 1223
rect 2031 1219 2035 1223
rect 207 1214 211 1218
rect 327 1214 331 1218
rect 455 1214 459 1218
rect 583 1214 587 1218
rect 719 1214 723 1218
rect 879 1214 883 1218
rect 1055 1214 1059 1218
rect 1263 1214 1267 1218
rect 1487 1214 1491 1218
rect 1719 1214 1723 1218
rect 1935 1214 1939 1218
rect 2111 1190 2115 1194
rect 2279 1190 2283 1194
rect 2471 1190 2475 1194
rect 2655 1190 2659 1194
rect 2831 1190 2835 1194
rect 2999 1190 3003 1194
rect 3159 1190 3163 1194
rect 3327 1190 3331 1194
rect 3495 1190 3499 1194
rect 2071 1185 2075 1189
rect 3991 1185 3995 1189
rect 471 1174 475 1178
rect 583 1174 587 1178
rect 703 1174 707 1178
rect 823 1174 827 1178
rect 943 1174 947 1178
rect 1063 1174 1067 1178
rect 1183 1174 1187 1178
rect 1303 1174 1307 1178
rect 1423 1174 1427 1178
rect 1543 1174 1547 1178
rect 111 1169 115 1173
rect 2031 1169 2035 1173
rect 2071 1168 2075 1172
rect 3991 1168 3995 1172
rect 111 1152 115 1156
rect 2031 1152 2035 1156
rect 2111 1149 2115 1153
rect 2279 1149 2283 1153
rect 2471 1149 2475 1153
rect 2655 1149 2659 1153
rect 2831 1149 2835 1153
rect 2999 1149 3003 1153
rect 3159 1149 3163 1153
rect 3327 1149 3331 1153
rect 3495 1149 3499 1153
rect 471 1133 475 1137
rect 583 1133 587 1137
rect 703 1133 707 1137
rect 823 1133 827 1137
rect 943 1133 947 1137
rect 1063 1133 1067 1137
rect 1183 1133 1187 1137
rect 1303 1133 1307 1137
rect 1423 1133 1427 1137
rect 1543 1133 1547 1137
rect 2111 1115 2115 1119
rect 2295 1115 2299 1119
rect 2503 1115 2507 1119
rect 2703 1115 2707 1119
rect 2895 1115 2899 1119
rect 3079 1115 3083 1119
rect 3255 1115 3259 1119
rect 3431 1115 3435 1119
rect 3615 1115 3619 1119
rect 623 1095 627 1099
rect 735 1095 739 1099
rect 855 1095 859 1099
rect 975 1095 979 1099
rect 1095 1095 1099 1099
rect 1215 1095 1219 1099
rect 1335 1095 1339 1099
rect 1455 1095 1459 1099
rect 1575 1095 1579 1099
rect 1703 1095 1707 1099
rect 2071 1096 2075 1100
rect 3991 1096 3995 1100
rect 111 1076 115 1080
rect 2031 1076 2035 1080
rect 2071 1079 2075 1083
rect 3991 1079 3995 1083
rect 2111 1074 2115 1078
rect 2295 1074 2299 1078
rect 2503 1074 2507 1078
rect 2703 1074 2707 1078
rect 2895 1074 2899 1078
rect 3079 1074 3083 1078
rect 3255 1074 3259 1078
rect 3431 1074 3435 1078
rect 3615 1074 3619 1078
rect 111 1059 115 1063
rect 2031 1059 2035 1063
rect 623 1054 627 1058
rect 735 1054 739 1058
rect 855 1054 859 1058
rect 975 1054 979 1058
rect 1095 1054 1099 1058
rect 1215 1054 1219 1058
rect 1335 1054 1339 1058
rect 1455 1054 1459 1058
rect 1575 1054 1579 1058
rect 1703 1054 1707 1058
rect 2167 1034 2171 1038
rect 2287 1034 2291 1038
rect 2423 1034 2427 1038
rect 2575 1034 2579 1038
rect 2743 1034 2747 1038
rect 2919 1034 2923 1038
rect 3095 1034 3099 1038
rect 3279 1034 3283 1038
rect 3463 1034 3467 1038
rect 3655 1034 3659 1038
rect 2071 1029 2075 1033
rect 3991 1029 3995 1033
rect 727 1014 731 1018
rect 847 1014 851 1018
rect 967 1014 971 1018
rect 1095 1014 1099 1018
rect 1223 1014 1227 1018
rect 1351 1014 1355 1018
rect 1479 1014 1483 1018
rect 1607 1014 1611 1018
rect 1735 1014 1739 1018
rect 1863 1014 1867 1018
rect 111 1009 115 1013
rect 2031 1009 2035 1013
rect 2071 1012 2075 1016
rect 3991 1012 3995 1016
rect 111 992 115 996
rect 2031 992 2035 996
rect 2167 993 2171 997
rect 2287 993 2291 997
rect 2423 993 2427 997
rect 2575 993 2579 997
rect 2743 993 2747 997
rect 2919 993 2923 997
rect 3095 993 3099 997
rect 3279 993 3283 997
rect 3463 993 3467 997
rect 3655 993 3659 997
rect 727 973 731 977
rect 847 973 851 977
rect 967 973 971 977
rect 1095 973 1099 977
rect 1223 973 1227 977
rect 1351 973 1355 977
rect 1479 973 1483 977
rect 1607 973 1611 977
rect 1735 973 1739 977
rect 1863 973 1867 977
rect 2527 955 2531 959
rect 2647 955 2651 959
rect 2775 955 2779 959
rect 2919 955 2923 959
rect 3071 955 3075 959
rect 3231 955 3235 959
rect 3399 955 3403 959
rect 3567 955 3571 959
rect 3735 955 3739 959
rect 591 935 595 939
rect 735 935 739 939
rect 887 935 891 939
rect 1039 935 1043 939
rect 1199 935 1203 939
rect 1351 935 1355 939
rect 1503 935 1507 939
rect 1655 935 1659 939
rect 1807 935 1811 939
rect 1935 935 1939 939
rect 2071 936 2075 940
rect 3991 936 3995 940
rect 111 916 115 920
rect 2031 916 2035 920
rect 2071 919 2075 923
rect 3991 919 3995 923
rect 2527 914 2531 918
rect 2647 914 2651 918
rect 2775 914 2779 918
rect 2919 914 2923 918
rect 3071 914 3075 918
rect 3231 914 3235 918
rect 3399 914 3403 918
rect 3567 914 3571 918
rect 3735 914 3739 918
rect 111 899 115 903
rect 2031 899 2035 903
rect 591 894 595 898
rect 735 894 739 898
rect 887 894 891 898
rect 1039 894 1043 898
rect 1199 894 1203 898
rect 1351 894 1355 898
rect 1503 894 1507 898
rect 1655 894 1659 898
rect 1807 894 1811 898
rect 1935 894 1939 898
rect 2455 870 2459 874
rect 2575 870 2579 874
rect 2711 870 2715 874
rect 2863 870 2867 874
rect 3015 870 3019 874
rect 3167 870 3171 874
rect 3319 870 3323 874
rect 3471 870 3475 874
rect 3615 870 3619 874
rect 3767 870 3771 874
rect 3895 870 3899 874
rect 2071 865 2075 869
rect 3991 865 3995 869
rect 439 854 443 858
rect 583 854 587 858
rect 735 854 739 858
rect 887 854 891 858
rect 1047 854 1051 858
rect 1199 854 1203 858
rect 1351 854 1355 858
rect 1495 854 1499 858
rect 1647 854 1651 858
rect 1799 854 1803 858
rect 111 849 115 853
rect 2031 849 2035 853
rect 2071 848 2075 852
rect 3991 848 3995 852
rect 111 832 115 836
rect 2031 832 2035 836
rect 2455 829 2459 833
rect 2575 829 2579 833
rect 2711 829 2715 833
rect 2863 829 2867 833
rect 3015 829 3019 833
rect 3167 829 3171 833
rect 3319 829 3323 833
rect 3471 829 3475 833
rect 3615 829 3619 833
rect 3767 829 3771 833
rect 3895 829 3899 833
rect 439 813 443 817
rect 583 813 587 817
rect 735 813 739 817
rect 887 813 891 817
rect 1047 813 1051 817
rect 1199 813 1203 817
rect 1351 813 1355 817
rect 1495 813 1499 817
rect 1647 813 1651 817
rect 1799 813 1803 817
rect 2215 799 2219 803
rect 2343 799 2347 803
rect 2479 799 2483 803
rect 2623 799 2627 803
rect 2783 799 2787 803
rect 2959 799 2963 803
rect 3167 799 3171 803
rect 3391 799 3395 803
rect 3623 799 3627 803
rect 3863 799 3867 803
rect 279 783 283 787
rect 431 783 435 787
rect 591 783 595 787
rect 751 783 755 787
rect 919 783 923 787
rect 1087 783 1091 787
rect 1255 783 1259 787
rect 1423 783 1427 787
rect 1591 783 1595 787
rect 2071 780 2075 784
rect 3991 780 3995 784
rect 111 764 115 768
rect 2031 764 2035 768
rect 2071 763 2075 767
rect 3991 763 3995 767
rect 2215 758 2219 762
rect 2343 758 2347 762
rect 2479 758 2483 762
rect 2623 758 2627 762
rect 2783 758 2787 762
rect 2959 758 2963 762
rect 3167 758 3171 762
rect 3391 758 3395 762
rect 3623 758 3627 762
rect 3863 758 3867 762
rect 111 747 115 751
rect 2031 747 2035 751
rect 279 742 283 746
rect 431 742 435 746
rect 591 742 595 746
rect 751 742 755 746
rect 919 742 923 746
rect 1087 742 1091 746
rect 1255 742 1259 746
rect 1423 742 1427 746
rect 1591 742 1595 746
rect 2111 718 2115 722
rect 2247 718 2251 722
rect 2423 718 2427 722
rect 2599 718 2603 722
rect 2783 718 2787 722
rect 2967 718 2971 722
rect 3151 718 3155 722
rect 3335 718 3339 722
rect 3519 718 3523 722
rect 3703 718 3707 722
rect 3895 718 3899 722
rect 2071 713 2075 717
rect 3991 713 3995 717
rect 151 706 155 710
rect 271 706 275 710
rect 423 706 427 710
rect 575 706 579 710
rect 735 706 739 710
rect 887 706 891 710
rect 1039 706 1043 710
rect 1191 706 1195 710
rect 1343 706 1347 710
rect 1495 706 1499 710
rect 111 701 115 705
rect 2031 701 2035 705
rect 2071 696 2075 700
rect 3991 696 3995 700
rect 111 684 115 688
rect 2031 684 2035 688
rect 2111 677 2115 681
rect 2247 677 2251 681
rect 2423 677 2427 681
rect 2599 677 2603 681
rect 2783 677 2787 681
rect 2967 677 2971 681
rect 3151 677 3155 681
rect 3335 677 3339 681
rect 3519 677 3523 681
rect 3703 677 3707 681
rect 3895 677 3899 681
rect 151 665 155 669
rect 271 665 275 669
rect 423 665 427 669
rect 575 665 579 669
rect 735 665 739 669
rect 887 665 891 669
rect 1039 665 1043 669
rect 1191 665 1195 669
rect 1343 665 1347 669
rect 1495 665 1499 669
rect 2111 643 2115 647
rect 2375 643 2379 647
rect 2655 643 2659 647
rect 2919 643 2923 647
rect 3175 643 3179 647
rect 3423 643 3427 647
rect 3671 643 3675 647
rect 3895 643 3899 647
rect 151 627 155 631
rect 255 627 259 631
rect 391 627 395 631
rect 527 627 531 631
rect 663 627 667 631
rect 807 627 811 631
rect 959 627 963 631
rect 1119 627 1123 631
rect 1287 627 1291 631
rect 1455 627 1459 631
rect 1623 627 1627 631
rect 1791 627 1795 631
rect 1935 627 1939 631
rect 2071 624 2075 628
rect 3991 624 3995 628
rect 111 608 115 612
rect 2031 608 2035 612
rect 2071 607 2075 611
rect 3991 607 3995 611
rect 2111 602 2115 606
rect 2375 602 2379 606
rect 2655 602 2659 606
rect 2919 602 2923 606
rect 3175 602 3179 606
rect 3423 602 3427 606
rect 3671 602 3675 606
rect 3895 602 3899 606
rect 111 591 115 595
rect 2031 591 2035 595
rect 151 586 155 590
rect 255 586 259 590
rect 391 586 395 590
rect 527 586 531 590
rect 663 586 667 590
rect 807 586 811 590
rect 959 586 963 590
rect 1119 586 1123 590
rect 1287 586 1291 590
rect 1455 586 1459 590
rect 1623 586 1627 590
rect 1791 586 1795 590
rect 1935 586 1939 590
rect 2111 558 2115 562
rect 2215 558 2219 562
rect 2351 558 2355 562
rect 2487 558 2491 562
rect 2631 558 2635 562
rect 2791 558 2795 562
rect 2975 558 2979 562
rect 3191 558 3195 562
rect 3423 558 3427 562
rect 3671 558 3675 562
rect 3895 558 3899 562
rect 2071 553 2075 557
rect 3991 553 3995 557
rect 207 542 211 546
rect 327 542 331 546
rect 447 542 451 546
rect 567 542 571 546
rect 687 542 691 546
rect 799 542 803 546
rect 911 542 915 546
rect 1031 542 1035 546
rect 1151 542 1155 546
rect 1271 542 1275 546
rect 111 537 115 541
rect 2031 537 2035 541
rect 2071 536 2075 540
rect 3991 536 3995 540
rect 111 520 115 524
rect 2031 520 2035 524
rect 2111 517 2115 521
rect 2215 517 2219 521
rect 2351 517 2355 521
rect 2487 517 2491 521
rect 2631 517 2635 521
rect 2791 517 2795 521
rect 2975 517 2979 521
rect 3191 517 3195 521
rect 3423 517 3427 521
rect 3671 517 3675 521
rect 3895 517 3899 521
rect 207 501 211 505
rect 327 501 331 505
rect 447 501 451 505
rect 567 501 571 505
rect 687 501 691 505
rect 799 501 803 505
rect 911 501 915 505
rect 1031 501 1035 505
rect 1151 501 1155 505
rect 1271 501 1275 505
rect 2423 483 2427 487
rect 2527 483 2531 487
rect 2631 483 2635 487
rect 2743 483 2747 487
rect 2871 483 2875 487
rect 3031 483 3035 487
rect 3223 483 3227 487
rect 3447 483 3451 487
rect 3679 483 3683 487
rect 3895 483 3899 487
rect 439 463 443 467
rect 543 463 547 467
rect 647 463 651 467
rect 751 463 755 467
rect 855 463 859 467
rect 959 463 963 467
rect 1063 463 1067 467
rect 1167 463 1171 467
rect 1271 463 1275 467
rect 1375 463 1379 467
rect 2071 464 2075 468
rect 3991 464 3995 468
rect 111 444 115 448
rect 2031 444 2035 448
rect 2071 447 2075 451
rect 3991 447 3995 451
rect 2423 442 2427 446
rect 2527 442 2531 446
rect 2631 442 2635 446
rect 2743 442 2747 446
rect 2871 442 2875 446
rect 3031 442 3035 446
rect 3223 442 3227 446
rect 3447 442 3451 446
rect 3679 442 3683 446
rect 3895 442 3899 446
rect 111 427 115 431
rect 2031 427 2035 431
rect 439 422 443 426
rect 543 422 547 426
rect 647 422 651 426
rect 751 422 755 426
rect 855 422 859 426
rect 959 422 963 426
rect 1063 422 1067 426
rect 1167 422 1171 426
rect 1271 422 1275 426
rect 1375 422 1379 426
rect 2527 406 2531 410
rect 2639 406 2643 410
rect 2775 406 2779 410
rect 2951 406 2955 410
rect 3159 406 3163 410
rect 3399 406 3403 410
rect 3655 406 3659 410
rect 3895 406 3899 410
rect 2071 401 2075 405
rect 3991 401 3995 405
rect 623 382 627 386
rect 727 382 731 386
rect 831 382 835 386
rect 935 382 939 386
rect 1039 382 1043 386
rect 1143 382 1147 386
rect 1247 382 1251 386
rect 1351 382 1355 386
rect 1455 382 1459 386
rect 1559 382 1563 386
rect 2071 384 2075 388
rect 3991 384 3995 388
rect 111 377 115 381
rect 2031 377 2035 381
rect 2527 365 2531 369
rect 111 360 115 364
rect 2639 365 2643 369
rect 2775 365 2779 369
rect 2951 365 2955 369
rect 3159 365 3163 369
rect 3399 365 3403 369
rect 3655 365 3659 369
rect 3895 365 3899 369
rect 2031 360 2035 364
rect 623 341 627 345
rect 727 341 731 345
rect 831 341 835 345
rect 935 341 939 345
rect 1039 341 1043 345
rect 1143 341 1147 345
rect 1247 341 1251 345
rect 1351 341 1355 345
rect 1455 341 1459 345
rect 1559 341 1563 345
rect 2271 323 2275 327
rect 2423 323 2427 327
rect 2583 323 2587 327
rect 2743 323 2747 327
rect 2911 323 2915 327
rect 3071 323 3075 327
rect 3223 323 3227 327
rect 3367 323 3371 327
rect 3503 323 3507 327
rect 3639 323 3643 327
rect 3775 323 3779 327
rect 3895 323 3899 327
rect 399 311 403 315
rect 543 311 547 315
rect 687 311 691 315
rect 839 311 843 315
rect 991 311 995 315
rect 1143 311 1147 315
rect 1303 311 1307 315
rect 1463 311 1467 315
rect 1623 311 1627 315
rect 2071 304 2075 308
rect 3991 304 3995 308
rect 111 292 115 296
rect 2031 292 2035 296
rect 2071 287 2075 291
rect 3991 287 3995 291
rect 2271 282 2275 286
rect 2423 282 2427 286
rect 2583 282 2587 286
rect 2743 282 2747 286
rect 2911 282 2915 286
rect 3071 282 3075 286
rect 3223 282 3227 286
rect 3367 282 3371 286
rect 3503 282 3507 286
rect 3639 282 3643 286
rect 3775 282 3779 286
rect 3895 282 3899 286
rect 111 275 115 279
rect 2031 275 2035 279
rect 399 270 403 274
rect 543 270 547 274
rect 687 270 691 274
rect 839 270 843 274
rect 991 270 995 274
rect 1143 270 1147 274
rect 1303 270 1307 274
rect 1463 270 1467 274
rect 1623 270 1627 274
rect 2111 242 2115 246
rect 2247 242 2251 246
rect 2423 242 2427 246
rect 2599 242 2603 246
rect 2775 242 2779 246
rect 2943 242 2947 246
rect 3103 242 3107 246
rect 3255 242 3259 246
rect 3391 242 3395 246
rect 3527 242 3531 246
rect 3655 242 3659 246
rect 3783 242 3787 246
rect 3895 242 3899 246
rect 207 234 211 238
rect 431 234 435 238
rect 655 234 659 238
rect 871 234 875 238
rect 1071 234 1075 238
rect 1263 234 1267 238
rect 1447 234 1451 238
rect 1631 234 1635 238
rect 1815 234 1819 238
rect 2071 237 2075 241
rect 3991 237 3995 241
rect 111 229 115 233
rect 2031 229 2035 233
rect 2071 220 2075 224
rect 3991 220 3995 224
rect 111 212 115 216
rect 2031 212 2035 216
rect 2111 201 2115 205
rect 2247 201 2251 205
rect 2423 201 2427 205
rect 2599 201 2603 205
rect 2775 201 2779 205
rect 2943 201 2947 205
rect 3103 201 3107 205
rect 3255 201 3259 205
rect 3391 201 3395 205
rect 3527 201 3531 205
rect 3655 201 3659 205
rect 3783 201 3787 205
rect 3895 201 3899 205
rect 207 193 211 197
rect 431 193 435 197
rect 655 193 659 197
rect 871 193 875 197
rect 1071 193 1075 197
rect 1263 193 1267 197
rect 1447 193 1451 197
rect 1631 193 1635 197
rect 1815 193 1819 197
rect 2111 159 2115 163
rect 2239 159 2243 163
rect 2399 159 2403 163
rect 2567 159 2571 163
rect 2735 159 2739 163
rect 2895 159 2899 163
rect 3047 159 3051 163
rect 3191 159 3195 163
rect 3327 159 3331 163
rect 3455 159 3459 163
rect 3591 159 3595 163
rect 3727 159 3731 163
rect 2071 140 2075 144
rect 151 135 155 139
rect 255 135 259 139
rect 359 135 363 139
rect 463 135 467 139
rect 567 135 571 139
rect 671 135 675 139
rect 775 135 779 139
rect 879 135 883 139
rect 983 135 987 139
rect 1087 135 1091 139
rect 1191 135 1195 139
rect 1295 135 1299 139
rect 1399 135 1403 139
rect 1511 135 1515 139
rect 1623 135 1627 139
rect 1727 135 1731 139
rect 1831 135 1835 139
rect 3991 140 3995 144
rect 1935 135 1939 139
rect 2071 123 2075 127
rect 3991 123 3995 127
rect 111 116 115 120
rect 2031 116 2035 120
rect 2111 118 2115 122
rect 2239 118 2243 122
rect 2399 118 2403 122
rect 2567 118 2571 122
rect 2735 118 2739 122
rect 2895 118 2899 122
rect 3047 118 3051 122
rect 3191 118 3195 122
rect 3327 118 3331 122
rect 3455 118 3459 122
rect 3591 118 3595 122
rect 3727 118 3731 122
rect 111 99 115 103
rect 2031 99 2035 103
rect 151 94 155 98
rect 255 94 259 98
rect 359 94 363 98
rect 463 94 467 98
rect 567 94 571 98
rect 671 94 675 98
rect 775 94 779 98
rect 879 94 883 98
rect 983 94 987 98
rect 1087 94 1091 98
rect 1191 94 1195 98
rect 1295 94 1299 98
rect 1399 94 1403 98
rect 1511 94 1515 98
rect 1623 94 1627 98
rect 1727 94 1731 98
rect 1831 94 1835 98
rect 1935 94 1939 98
<< m3 >>
rect 2071 4082 2075 4083
rect 2071 4077 2075 4078
rect 3399 4082 3403 4083
rect 3399 4077 3403 4078
rect 3503 4082 3507 4083
rect 3503 4077 3507 4078
rect 3607 4082 3611 4083
rect 3607 4077 3611 4078
rect 3711 4082 3715 4083
rect 3711 4077 3715 4078
rect 3991 4082 3995 4083
rect 3991 4077 3995 4078
rect 2072 4049 2074 4077
rect 3400 4068 3402 4077
rect 3504 4068 3506 4077
rect 3608 4068 3610 4077
rect 3712 4068 3714 4077
rect 3398 4067 3404 4068
rect 3398 4063 3399 4067
rect 3403 4063 3404 4067
rect 3398 4062 3404 4063
rect 3502 4067 3508 4068
rect 3502 4063 3503 4067
rect 3507 4063 3508 4067
rect 3502 4062 3508 4063
rect 3606 4067 3612 4068
rect 3606 4063 3607 4067
rect 3611 4063 3612 4067
rect 3606 4062 3612 4063
rect 3710 4067 3716 4068
rect 3710 4063 3711 4067
rect 3715 4063 3716 4067
rect 3710 4062 3716 4063
rect 3992 4049 3994 4077
rect 2070 4048 2076 4049
rect 111 4046 115 4047
rect 111 4041 115 4042
rect 495 4046 499 4047
rect 495 4041 499 4042
rect 599 4046 603 4047
rect 599 4041 603 4042
rect 703 4046 707 4047
rect 703 4041 707 4042
rect 807 4046 811 4047
rect 807 4041 811 4042
rect 911 4046 915 4047
rect 911 4041 915 4042
rect 1015 4046 1019 4047
rect 1015 4041 1019 4042
rect 1119 4046 1123 4047
rect 1119 4041 1123 4042
rect 1223 4046 1227 4047
rect 1223 4041 1227 4042
rect 1327 4046 1331 4047
rect 1327 4041 1331 4042
rect 1431 4046 1435 4047
rect 1431 4041 1435 4042
rect 2031 4046 2035 4047
rect 2070 4044 2071 4048
rect 2075 4044 2076 4048
rect 2070 4043 2076 4044
rect 3990 4048 3996 4049
rect 3990 4044 3991 4048
rect 3995 4044 3996 4048
rect 3990 4043 3996 4044
rect 2031 4041 2035 4042
rect 112 4013 114 4041
rect 496 4032 498 4041
rect 600 4032 602 4041
rect 704 4032 706 4041
rect 808 4032 810 4041
rect 912 4032 914 4041
rect 1016 4032 1018 4041
rect 1120 4032 1122 4041
rect 1224 4032 1226 4041
rect 1328 4032 1330 4041
rect 1432 4032 1434 4041
rect 494 4031 500 4032
rect 494 4027 495 4031
rect 499 4027 500 4031
rect 494 4026 500 4027
rect 598 4031 604 4032
rect 598 4027 599 4031
rect 603 4027 604 4031
rect 598 4026 604 4027
rect 702 4031 708 4032
rect 702 4027 703 4031
rect 707 4027 708 4031
rect 702 4026 708 4027
rect 806 4031 812 4032
rect 806 4027 807 4031
rect 811 4027 812 4031
rect 806 4026 812 4027
rect 910 4031 916 4032
rect 910 4027 911 4031
rect 915 4027 916 4031
rect 910 4026 916 4027
rect 1014 4031 1020 4032
rect 1014 4027 1015 4031
rect 1019 4027 1020 4031
rect 1014 4026 1020 4027
rect 1118 4031 1124 4032
rect 1118 4027 1119 4031
rect 1123 4027 1124 4031
rect 1118 4026 1124 4027
rect 1222 4031 1228 4032
rect 1222 4027 1223 4031
rect 1227 4027 1228 4031
rect 1222 4026 1228 4027
rect 1326 4031 1332 4032
rect 1326 4027 1327 4031
rect 1331 4027 1332 4031
rect 1326 4026 1332 4027
rect 1430 4031 1436 4032
rect 1430 4027 1431 4031
rect 1435 4027 1436 4031
rect 1430 4026 1436 4027
rect 2032 4013 2034 4041
rect 2070 4031 2076 4032
rect 2070 4027 2071 4031
rect 2075 4027 2076 4031
rect 3990 4031 3996 4032
rect 3990 4027 3991 4031
rect 3995 4027 3996 4031
rect 2070 4026 2076 4027
rect 3398 4026 3404 4027
rect 110 4012 116 4013
rect 110 4008 111 4012
rect 115 4008 116 4012
rect 110 4007 116 4008
rect 2030 4012 2036 4013
rect 2030 4008 2031 4012
rect 2035 4008 2036 4012
rect 2072 4011 2074 4026
rect 3398 4022 3399 4026
rect 3403 4022 3404 4026
rect 3398 4021 3404 4022
rect 3502 4026 3508 4027
rect 3502 4022 3503 4026
rect 3507 4022 3508 4026
rect 3502 4021 3508 4022
rect 3606 4026 3612 4027
rect 3606 4022 3607 4026
rect 3611 4022 3612 4026
rect 3606 4021 3612 4022
rect 3710 4026 3716 4027
rect 3990 4026 3996 4027
rect 3710 4022 3711 4026
rect 3715 4022 3716 4026
rect 3710 4021 3716 4022
rect 3400 4011 3402 4021
rect 3504 4011 3506 4021
rect 3608 4011 3610 4021
rect 3712 4011 3714 4021
rect 3992 4011 3994 4026
rect 2030 4007 2036 4008
rect 2071 4010 2075 4011
rect 2071 4005 2075 4006
rect 2111 4010 2115 4011
rect 2111 4005 2115 4006
rect 2215 4010 2219 4011
rect 2215 4005 2219 4006
rect 2319 4010 2323 4011
rect 2319 4005 2323 4006
rect 2423 4010 2427 4011
rect 2423 4005 2427 4006
rect 2527 4010 2531 4011
rect 2527 4005 2531 4006
rect 2647 4010 2651 4011
rect 2647 4005 2651 4006
rect 2775 4010 2779 4011
rect 2775 4005 2779 4006
rect 2903 4010 2907 4011
rect 2903 4005 2907 4006
rect 3031 4010 3035 4011
rect 3031 4005 3035 4006
rect 3159 4010 3163 4011
rect 3159 4005 3163 4006
rect 3287 4010 3291 4011
rect 3287 4005 3291 4006
rect 3399 4010 3403 4011
rect 3399 4005 3403 4006
rect 3415 4010 3419 4011
rect 3415 4005 3419 4006
rect 3503 4010 3507 4011
rect 3503 4005 3507 4006
rect 3551 4010 3555 4011
rect 3551 4005 3555 4006
rect 3607 4010 3611 4011
rect 3607 4005 3611 4006
rect 3711 4010 3715 4011
rect 3711 4005 3715 4006
rect 3991 4010 3995 4011
rect 3991 4005 3995 4006
rect 110 3995 116 3996
rect 110 3991 111 3995
rect 115 3991 116 3995
rect 2030 3995 2036 3996
rect 2030 3991 2031 3995
rect 2035 3991 2036 3995
rect 110 3990 116 3991
rect 494 3990 500 3991
rect 112 3975 114 3990
rect 494 3986 495 3990
rect 499 3986 500 3990
rect 494 3985 500 3986
rect 598 3990 604 3991
rect 598 3986 599 3990
rect 603 3986 604 3990
rect 598 3985 604 3986
rect 702 3990 708 3991
rect 702 3986 703 3990
rect 707 3986 708 3990
rect 702 3985 708 3986
rect 806 3990 812 3991
rect 806 3986 807 3990
rect 811 3986 812 3990
rect 806 3985 812 3986
rect 910 3990 916 3991
rect 910 3986 911 3990
rect 915 3986 916 3990
rect 910 3985 916 3986
rect 1014 3990 1020 3991
rect 1014 3986 1015 3990
rect 1019 3986 1020 3990
rect 1014 3985 1020 3986
rect 1118 3990 1124 3991
rect 1118 3986 1119 3990
rect 1123 3986 1124 3990
rect 1118 3985 1124 3986
rect 1222 3990 1228 3991
rect 1222 3986 1223 3990
rect 1227 3986 1228 3990
rect 1222 3985 1228 3986
rect 1326 3990 1332 3991
rect 1326 3986 1327 3990
rect 1331 3986 1332 3990
rect 1326 3985 1332 3986
rect 1430 3990 1436 3991
rect 2030 3990 2036 3991
rect 2072 3990 2074 4005
rect 2112 3995 2114 4005
rect 2216 3995 2218 4005
rect 2320 3995 2322 4005
rect 2424 3995 2426 4005
rect 2528 3995 2530 4005
rect 2648 3995 2650 4005
rect 2776 3995 2778 4005
rect 2904 3995 2906 4005
rect 3032 3995 3034 4005
rect 3160 3995 3162 4005
rect 3288 3995 3290 4005
rect 3416 3995 3418 4005
rect 3552 3995 3554 4005
rect 2110 3994 2116 3995
rect 2110 3990 2111 3994
rect 2115 3990 2116 3994
rect 1430 3986 1431 3990
rect 1435 3986 1436 3990
rect 1430 3985 1436 3986
rect 496 3975 498 3985
rect 600 3975 602 3985
rect 704 3975 706 3985
rect 808 3975 810 3985
rect 912 3975 914 3985
rect 1016 3975 1018 3985
rect 1120 3975 1122 3985
rect 1224 3975 1226 3985
rect 1328 3975 1330 3985
rect 1432 3975 1434 3985
rect 2032 3975 2034 3990
rect 2070 3989 2076 3990
rect 2110 3989 2116 3990
rect 2214 3994 2220 3995
rect 2214 3990 2215 3994
rect 2219 3990 2220 3994
rect 2214 3989 2220 3990
rect 2318 3994 2324 3995
rect 2318 3990 2319 3994
rect 2323 3990 2324 3994
rect 2318 3989 2324 3990
rect 2422 3994 2428 3995
rect 2422 3990 2423 3994
rect 2427 3990 2428 3994
rect 2422 3989 2428 3990
rect 2526 3994 2532 3995
rect 2526 3990 2527 3994
rect 2531 3990 2532 3994
rect 2526 3989 2532 3990
rect 2646 3994 2652 3995
rect 2646 3990 2647 3994
rect 2651 3990 2652 3994
rect 2646 3989 2652 3990
rect 2774 3994 2780 3995
rect 2774 3990 2775 3994
rect 2779 3990 2780 3994
rect 2774 3989 2780 3990
rect 2902 3994 2908 3995
rect 2902 3990 2903 3994
rect 2907 3990 2908 3994
rect 2902 3989 2908 3990
rect 3030 3994 3036 3995
rect 3030 3990 3031 3994
rect 3035 3990 3036 3994
rect 3030 3989 3036 3990
rect 3158 3994 3164 3995
rect 3158 3990 3159 3994
rect 3163 3990 3164 3994
rect 3158 3989 3164 3990
rect 3286 3994 3292 3995
rect 3286 3990 3287 3994
rect 3291 3990 3292 3994
rect 3286 3989 3292 3990
rect 3414 3994 3420 3995
rect 3414 3990 3415 3994
rect 3419 3990 3420 3994
rect 3414 3989 3420 3990
rect 3550 3994 3556 3995
rect 3550 3990 3551 3994
rect 3555 3990 3556 3994
rect 3992 3990 3994 4005
rect 3550 3989 3556 3990
rect 3990 3989 3996 3990
rect 2070 3985 2071 3989
rect 2075 3985 2076 3989
rect 2070 3984 2076 3985
rect 3990 3985 3991 3989
rect 3995 3985 3996 3989
rect 3990 3984 3996 3985
rect 111 3974 115 3975
rect 111 3969 115 3970
rect 391 3974 395 3975
rect 391 3969 395 3970
rect 495 3974 499 3975
rect 495 3969 499 3970
rect 599 3974 603 3975
rect 599 3969 603 3970
rect 703 3974 707 3975
rect 703 3969 707 3970
rect 807 3974 811 3975
rect 807 3969 811 3970
rect 911 3974 915 3975
rect 911 3969 915 3970
rect 1015 3974 1019 3975
rect 1015 3969 1019 3970
rect 1119 3974 1123 3975
rect 1119 3969 1123 3970
rect 1223 3974 1227 3975
rect 1223 3969 1227 3970
rect 1327 3974 1331 3975
rect 1327 3969 1331 3970
rect 1431 3974 1435 3975
rect 1431 3969 1435 3970
rect 1535 3974 1539 3975
rect 1535 3969 1539 3970
rect 2031 3974 2035 3975
rect 2031 3969 2035 3970
rect 2070 3972 2076 3973
rect 112 3954 114 3969
rect 392 3959 394 3969
rect 496 3959 498 3969
rect 600 3959 602 3969
rect 704 3959 706 3969
rect 808 3959 810 3969
rect 912 3959 914 3969
rect 1016 3959 1018 3969
rect 1120 3959 1122 3969
rect 1224 3959 1226 3969
rect 1328 3959 1330 3969
rect 1432 3959 1434 3969
rect 1536 3959 1538 3969
rect 390 3958 396 3959
rect 390 3954 391 3958
rect 395 3954 396 3958
rect 110 3953 116 3954
rect 390 3953 396 3954
rect 494 3958 500 3959
rect 494 3954 495 3958
rect 499 3954 500 3958
rect 494 3953 500 3954
rect 598 3958 604 3959
rect 598 3954 599 3958
rect 603 3954 604 3958
rect 598 3953 604 3954
rect 702 3958 708 3959
rect 702 3954 703 3958
rect 707 3954 708 3958
rect 702 3953 708 3954
rect 806 3958 812 3959
rect 806 3954 807 3958
rect 811 3954 812 3958
rect 806 3953 812 3954
rect 910 3958 916 3959
rect 910 3954 911 3958
rect 915 3954 916 3958
rect 910 3953 916 3954
rect 1014 3958 1020 3959
rect 1014 3954 1015 3958
rect 1019 3954 1020 3958
rect 1014 3953 1020 3954
rect 1118 3958 1124 3959
rect 1118 3954 1119 3958
rect 1123 3954 1124 3958
rect 1118 3953 1124 3954
rect 1222 3958 1228 3959
rect 1222 3954 1223 3958
rect 1227 3954 1228 3958
rect 1222 3953 1228 3954
rect 1326 3958 1332 3959
rect 1326 3954 1327 3958
rect 1331 3954 1332 3958
rect 1326 3953 1332 3954
rect 1430 3958 1436 3959
rect 1430 3954 1431 3958
rect 1435 3954 1436 3958
rect 1430 3953 1436 3954
rect 1534 3958 1540 3959
rect 1534 3954 1535 3958
rect 1539 3954 1540 3958
rect 2032 3954 2034 3969
rect 2070 3968 2071 3972
rect 2075 3968 2076 3972
rect 2070 3967 2076 3968
rect 3990 3972 3996 3973
rect 3990 3968 3991 3972
rect 3995 3968 3996 3972
rect 3990 3967 3996 3968
rect 1534 3953 1540 3954
rect 2030 3953 2036 3954
rect 110 3949 111 3953
rect 115 3949 116 3953
rect 110 3948 116 3949
rect 2030 3949 2031 3953
rect 2035 3949 2036 3953
rect 2030 3948 2036 3949
rect 110 3936 116 3937
rect 110 3932 111 3936
rect 115 3932 116 3936
rect 110 3931 116 3932
rect 2030 3936 2036 3937
rect 2030 3932 2031 3936
rect 2035 3932 2036 3936
rect 2072 3935 2074 3967
rect 2110 3953 2116 3954
rect 2110 3949 2111 3953
rect 2115 3949 2116 3953
rect 2110 3948 2116 3949
rect 2214 3953 2220 3954
rect 2214 3949 2215 3953
rect 2219 3949 2220 3953
rect 2214 3948 2220 3949
rect 2318 3953 2324 3954
rect 2318 3949 2319 3953
rect 2323 3949 2324 3953
rect 2318 3948 2324 3949
rect 2422 3953 2428 3954
rect 2422 3949 2423 3953
rect 2427 3949 2428 3953
rect 2422 3948 2428 3949
rect 2526 3953 2532 3954
rect 2526 3949 2527 3953
rect 2531 3949 2532 3953
rect 2526 3948 2532 3949
rect 2646 3953 2652 3954
rect 2646 3949 2647 3953
rect 2651 3949 2652 3953
rect 2646 3948 2652 3949
rect 2774 3953 2780 3954
rect 2774 3949 2775 3953
rect 2779 3949 2780 3953
rect 2774 3948 2780 3949
rect 2902 3953 2908 3954
rect 2902 3949 2903 3953
rect 2907 3949 2908 3953
rect 2902 3948 2908 3949
rect 3030 3953 3036 3954
rect 3030 3949 3031 3953
rect 3035 3949 3036 3953
rect 3030 3948 3036 3949
rect 3158 3953 3164 3954
rect 3158 3949 3159 3953
rect 3163 3949 3164 3953
rect 3158 3948 3164 3949
rect 3286 3953 3292 3954
rect 3286 3949 3287 3953
rect 3291 3949 3292 3953
rect 3286 3948 3292 3949
rect 3414 3953 3420 3954
rect 3414 3949 3415 3953
rect 3419 3949 3420 3953
rect 3414 3948 3420 3949
rect 3550 3953 3556 3954
rect 3550 3949 3551 3953
rect 3555 3949 3556 3953
rect 3550 3948 3556 3949
rect 2112 3935 2114 3948
rect 2216 3935 2218 3948
rect 2320 3935 2322 3948
rect 2424 3935 2426 3948
rect 2528 3935 2530 3948
rect 2648 3935 2650 3948
rect 2776 3935 2778 3948
rect 2904 3935 2906 3948
rect 3032 3935 3034 3948
rect 3160 3935 3162 3948
rect 3288 3935 3290 3948
rect 3416 3935 3418 3948
rect 3552 3935 3554 3948
rect 3992 3935 3994 3967
rect 2030 3931 2036 3932
rect 2071 3934 2075 3935
rect 112 3899 114 3931
rect 390 3917 396 3918
rect 390 3913 391 3917
rect 395 3913 396 3917
rect 390 3912 396 3913
rect 494 3917 500 3918
rect 494 3913 495 3917
rect 499 3913 500 3917
rect 494 3912 500 3913
rect 598 3917 604 3918
rect 598 3913 599 3917
rect 603 3913 604 3917
rect 598 3912 604 3913
rect 702 3917 708 3918
rect 702 3913 703 3917
rect 707 3913 708 3917
rect 702 3912 708 3913
rect 806 3917 812 3918
rect 806 3913 807 3917
rect 811 3913 812 3917
rect 806 3912 812 3913
rect 910 3917 916 3918
rect 910 3913 911 3917
rect 915 3913 916 3917
rect 910 3912 916 3913
rect 1014 3917 1020 3918
rect 1014 3913 1015 3917
rect 1019 3913 1020 3917
rect 1014 3912 1020 3913
rect 1118 3917 1124 3918
rect 1118 3913 1119 3917
rect 1123 3913 1124 3917
rect 1118 3912 1124 3913
rect 1222 3917 1228 3918
rect 1222 3913 1223 3917
rect 1227 3913 1228 3917
rect 1222 3912 1228 3913
rect 1326 3917 1332 3918
rect 1326 3913 1327 3917
rect 1331 3913 1332 3917
rect 1326 3912 1332 3913
rect 1430 3917 1436 3918
rect 1430 3913 1431 3917
rect 1435 3913 1436 3917
rect 1430 3912 1436 3913
rect 1534 3917 1540 3918
rect 1534 3913 1535 3917
rect 1539 3913 1540 3917
rect 1534 3912 1540 3913
rect 392 3899 394 3912
rect 496 3899 498 3912
rect 600 3899 602 3912
rect 704 3899 706 3912
rect 808 3899 810 3912
rect 912 3899 914 3912
rect 1016 3899 1018 3912
rect 1120 3899 1122 3912
rect 1224 3899 1226 3912
rect 1328 3899 1330 3912
rect 1432 3899 1434 3912
rect 1536 3899 1538 3912
rect 2032 3899 2034 3931
rect 2071 3929 2075 3930
rect 2111 3934 2115 3935
rect 2111 3929 2115 3930
rect 2143 3934 2147 3935
rect 2143 3929 2147 3930
rect 2215 3934 2219 3935
rect 2215 3929 2219 3930
rect 2319 3934 2323 3935
rect 2319 3929 2323 3930
rect 2423 3934 2427 3935
rect 2423 3929 2427 3930
rect 2487 3934 2491 3935
rect 2487 3929 2491 3930
rect 2527 3934 2531 3935
rect 2527 3929 2531 3930
rect 2647 3934 2651 3935
rect 2647 3929 2651 3930
rect 2775 3934 2779 3935
rect 2775 3929 2779 3930
rect 2799 3934 2803 3935
rect 2799 3929 2803 3930
rect 2903 3934 2907 3935
rect 2903 3929 2907 3930
rect 2951 3934 2955 3935
rect 2951 3929 2955 3930
rect 3031 3934 3035 3935
rect 3031 3929 3035 3930
rect 3103 3934 3107 3935
rect 3103 3929 3107 3930
rect 3159 3934 3163 3935
rect 3159 3929 3163 3930
rect 3255 3934 3259 3935
rect 3255 3929 3259 3930
rect 3287 3934 3291 3935
rect 3287 3929 3291 3930
rect 3415 3934 3419 3935
rect 3415 3929 3419 3930
rect 3551 3934 3555 3935
rect 3551 3929 3555 3930
rect 3991 3934 3995 3935
rect 3991 3929 3995 3930
rect 2072 3901 2074 3929
rect 2144 3920 2146 3929
rect 2320 3920 2322 3929
rect 2488 3920 2490 3929
rect 2648 3920 2650 3929
rect 2800 3920 2802 3929
rect 2952 3920 2954 3929
rect 3104 3920 3106 3929
rect 3256 3920 3258 3929
rect 2142 3919 2148 3920
rect 2142 3915 2143 3919
rect 2147 3915 2148 3919
rect 2142 3914 2148 3915
rect 2318 3919 2324 3920
rect 2318 3915 2319 3919
rect 2323 3915 2324 3919
rect 2318 3914 2324 3915
rect 2486 3919 2492 3920
rect 2486 3915 2487 3919
rect 2491 3915 2492 3919
rect 2486 3914 2492 3915
rect 2646 3919 2652 3920
rect 2646 3915 2647 3919
rect 2651 3915 2652 3919
rect 2646 3914 2652 3915
rect 2798 3919 2804 3920
rect 2798 3915 2799 3919
rect 2803 3915 2804 3919
rect 2798 3914 2804 3915
rect 2950 3919 2956 3920
rect 2950 3915 2951 3919
rect 2955 3915 2956 3919
rect 2950 3914 2956 3915
rect 3102 3919 3108 3920
rect 3102 3915 3103 3919
rect 3107 3915 3108 3919
rect 3102 3914 3108 3915
rect 3254 3919 3260 3920
rect 3254 3915 3255 3919
rect 3259 3915 3260 3919
rect 3254 3914 3260 3915
rect 3992 3901 3994 3929
rect 2070 3900 2076 3901
rect 111 3898 115 3899
rect 111 3893 115 3894
rect 375 3898 379 3899
rect 375 3893 379 3894
rect 391 3898 395 3899
rect 391 3893 395 3894
rect 495 3898 499 3899
rect 495 3893 499 3894
rect 599 3898 603 3899
rect 599 3893 603 3894
rect 623 3898 627 3899
rect 623 3893 627 3894
rect 703 3898 707 3899
rect 703 3893 707 3894
rect 759 3898 763 3899
rect 759 3893 763 3894
rect 807 3898 811 3899
rect 807 3893 811 3894
rect 895 3898 899 3899
rect 895 3893 899 3894
rect 911 3898 915 3899
rect 911 3893 915 3894
rect 1015 3898 1019 3899
rect 1015 3893 1019 3894
rect 1023 3898 1027 3899
rect 1023 3893 1027 3894
rect 1119 3898 1123 3899
rect 1119 3893 1123 3894
rect 1151 3898 1155 3899
rect 1151 3893 1155 3894
rect 1223 3898 1227 3899
rect 1223 3893 1227 3894
rect 1279 3898 1283 3899
rect 1279 3893 1283 3894
rect 1327 3898 1331 3899
rect 1327 3893 1331 3894
rect 1415 3898 1419 3899
rect 1415 3893 1419 3894
rect 1431 3898 1435 3899
rect 1431 3893 1435 3894
rect 1535 3898 1539 3899
rect 1535 3893 1539 3894
rect 1551 3898 1555 3899
rect 1551 3893 1555 3894
rect 2031 3898 2035 3899
rect 2070 3896 2071 3900
rect 2075 3896 2076 3900
rect 2070 3895 2076 3896
rect 3990 3900 3996 3901
rect 3990 3896 3991 3900
rect 3995 3896 3996 3900
rect 3990 3895 3996 3896
rect 2031 3893 2035 3894
rect 112 3865 114 3893
rect 376 3884 378 3893
rect 496 3884 498 3893
rect 624 3884 626 3893
rect 760 3884 762 3893
rect 896 3884 898 3893
rect 1024 3884 1026 3893
rect 1152 3884 1154 3893
rect 1280 3884 1282 3893
rect 1416 3884 1418 3893
rect 1552 3884 1554 3893
rect 374 3883 380 3884
rect 374 3879 375 3883
rect 379 3879 380 3883
rect 374 3878 380 3879
rect 494 3883 500 3884
rect 494 3879 495 3883
rect 499 3879 500 3883
rect 494 3878 500 3879
rect 622 3883 628 3884
rect 622 3879 623 3883
rect 627 3879 628 3883
rect 622 3878 628 3879
rect 758 3883 764 3884
rect 758 3879 759 3883
rect 763 3879 764 3883
rect 758 3878 764 3879
rect 894 3883 900 3884
rect 894 3879 895 3883
rect 899 3879 900 3883
rect 894 3878 900 3879
rect 1022 3883 1028 3884
rect 1022 3879 1023 3883
rect 1027 3879 1028 3883
rect 1022 3878 1028 3879
rect 1150 3883 1156 3884
rect 1150 3879 1151 3883
rect 1155 3879 1156 3883
rect 1150 3878 1156 3879
rect 1278 3883 1284 3884
rect 1278 3879 1279 3883
rect 1283 3879 1284 3883
rect 1278 3878 1284 3879
rect 1414 3883 1420 3884
rect 1414 3879 1415 3883
rect 1419 3879 1420 3883
rect 1414 3878 1420 3879
rect 1550 3883 1556 3884
rect 1550 3879 1551 3883
rect 1555 3879 1556 3883
rect 1550 3878 1556 3879
rect 2032 3865 2034 3893
rect 2070 3883 2076 3884
rect 2070 3879 2071 3883
rect 2075 3879 2076 3883
rect 3990 3883 3996 3884
rect 3990 3879 3991 3883
rect 3995 3879 3996 3883
rect 2070 3878 2076 3879
rect 2142 3878 2148 3879
rect 110 3864 116 3865
rect 110 3860 111 3864
rect 115 3860 116 3864
rect 110 3859 116 3860
rect 2030 3864 2036 3865
rect 2030 3860 2031 3864
rect 2035 3860 2036 3864
rect 2072 3863 2074 3878
rect 2142 3874 2143 3878
rect 2147 3874 2148 3878
rect 2142 3873 2148 3874
rect 2318 3878 2324 3879
rect 2318 3874 2319 3878
rect 2323 3874 2324 3878
rect 2318 3873 2324 3874
rect 2486 3878 2492 3879
rect 2486 3874 2487 3878
rect 2491 3874 2492 3878
rect 2486 3873 2492 3874
rect 2646 3878 2652 3879
rect 2646 3874 2647 3878
rect 2651 3874 2652 3878
rect 2646 3873 2652 3874
rect 2798 3878 2804 3879
rect 2798 3874 2799 3878
rect 2803 3874 2804 3878
rect 2798 3873 2804 3874
rect 2950 3878 2956 3879
rect 2950 3874 2951 3878
rect 2955 3874 2956 3878
rect 2950 3873 2956 3874
rect 3102 3878 3108 3879
rect 3102 3874 3103 3878
rect 3107 3874 3108 3878
rect 3102 3873 3108 3874
rect 3254 3878 3260 3879
rect 3990 3878 3996 3879
rect 3254 3874 3255 3878
rect 3259 3874 3260 3878
rect 3254 3873 3260 3874
rect 2144 3863 2146 3873
rect 2320 3863 2322 3873
rect 2488 3863 2490 3873
rect 2648 3863 2650 3873
rect 2800 3863 2802 3873
rect 2952 3863 2954 3873
rect 3104 3863 3106 3873
rect 3256 3863 3258 3873
rect 3992 3863 3994 3878
rect 2030 3859 2036 3860
rect 2071 3862 2075 3863
rect 2071 3857 2075 3858
rect 2119 3862 2123 3863
rect 2119 3857 2123 3858
rect 2143 3862 2147 3863
rect 2143 3857 2147 3858
rect 2287 3862 2291 3863
rect 2287 3857 2291 3858
rect 2319 3862 2323 3863
rect 2319 3857 2323 3858
rect 2447 3862 2451 3863
rect 2447 3857 2451 3858
rect 2487 3862 2491 3863
rect 2487 3857 2491 3858
rect 2599 3862 2603 3863
rect 2599 3857 2603 3858
rect 2647 3862 2651 3863
rect 2647 3857 2651 3858
rect 2743 3862 2747 3863
rect 2743 3857 2747 3858
rect 2799 3862 2803 3863
rect 2799 3857 2803 3858
rect 2879 3862 2883 3863
rect 2879 3857 2883 3858
rect 2951 3862 2955 3863
rect 2951 3857 2955 3858
rect 3023 3862 3027 3863
rect 3023 3857 3027 3858
rect 3103 3862 3107 3863
rect 3103 3857 3107 3858
rect 3167 3862 3171 3863
rect 3167 3857 3171 3858
rect 3255 3862 3259 3863
rect 3255 3857 3259 3858
rect 3991 3862 3995 3863
rect 3991 3857 3995 3858
rect 110 3847 116 3848
rect 110 3843 111 3847
rect 115 3843 116 3847
rect 2030 3847 2036 3848
rect 2030 3843 2031 3847
rect 2035 3843 2036 3847
rect 110 3842 116 3843
rect 374 3842 380 3843
rect 112 3819 114 3842
rect 374 3838 375 3842
rect 379 3838 380 3842
rect 374 3837 380 3838
rect 494 3842 500 3843
rect 494 3838 495 3842
rect 499 3838 500 3842
rect 494 3837 500 3838
rect 622 3842 628 3843
rect 622 3838 623 3842
rect 627 3838 628 3842
rect 622 3837 628 3838
rect 758 3842 764 3843
rect 758 3838 759 3842
rect 763 3838 764 3842
rect 758 3837 764 3838
rect 894 3842 900 3843
rect 894 3838 895 3842
rect 899 3838 900 3842
rect 894 3837 900 3838
rect 1022 3842 1028 3843
rect 1022 3838 1023 3842
rect 1027 3838 1028 3842
rect 1022 3837 1028 3838
rect 1150 3842 1156 3843
rect 1150 3838 1151 3842
rect 1155 3838 1156 3842
rect 1150 3837 1156 3838
rect 1278 3842 1284 3843
rect 1278 3838 1279 3842
rect 1283 3838 1284 3842
rect 1278 3837 1284 3838
rect 1414 3842 1420 3843
rect 1414 3838 1415 3842
rect 1419 3838 1420 3842
rect 1414 3837 1420 3838
rect 1550 3842 1556 3843
rect 2030 3842 2036 3843
rect 2072 3842 2074 3857
rect 2120 3847 2122 3857
rect 2288 3847 2290 3857
rect 2448 3847 2450 3857
rect 2600 3847 2602 3857
rect 2744 3847 2746 3857
rect 2880 3847 2882 3857
rect 3024 3847 3026 3857
rect 3168 3847 3170 3857
rect 2118 3846 2124 3847
rect 2118 3842 2119 3846
rect 2123 3842 2124 3846
rect 1550 3838 1551 3842
rect 1555 3838 1556 3842
rect 1550 3837 1556 3838
rect 376 3819 378 3837
rect 496 3819 498 3837
rect 624 3819 626 3837
rect 760 3819 762 3837
rect 896 3819 898 3837
rect 1024 3819 1026 3837
rect 1152 3819 1154 3837
rect 1280 3819 1282 3837
rect 1416 3819 1418 3837
rect 1552 3819 1554 3837
rect 2032 3819 2034 3842
rect 2070 3841 2076 3842
rect 2118 3841 2124 3842
rect 2286 3846 2292 3847
rect 2286 3842 2287 3846
rect 2291 3842 2292 3846
rect 2286 3841 2292 3842
rect 2446 3846 2452 3847
rect 2446 3842 2447 3846
rect 2451 3842 2452 3846
rect 2446 3841 2452 3842
rect 2598 3846 2604 3847
rect 2598 3842 2599 3846
rect 2603 3842 2604 3846
rect 2598 3841 2604 3842
rect 2742 3846 2748 3847
rect 2742 3842 2743 3846
rect 2747 3842 2748 3846
rect 2742 3841 2748 3842
rect 2878 3846 2884 3847
rect 2878 3842 2879 3846
rect 2883 3842 2884 3846
rect 2878 3841 2884 3842
rect 3022 3846 3028 3847
rect 3022 3842 3023 3846
rect 3027 3842 3028 3846
rect 3022 3841 3028 3842
rect 3166 3846 3172 3847
rect 3166 3842 3167 3846
rect 3171 3842 3172 3846
rect 3992 3842 3994 3857
rect 3166 3841 3172 3842
rect 3990 3841 3996 3842
rect 2070 3837 2071 3841
rect 2075 3837 2076 3841
rect 2070 3836 2076 3837
rect 3990 3837 3991 3841
rect 3995 3837 3996 3841
rect 3990 3836 3996 3837
rect 2070 3824 2076 3825
rect 2070 3820 2071 3824
rect 2075 3820 2076 3824
rect 2070 3819 2076 3820
rect 3990 3824 3996 3825
rect 3990 3820 3991 3824
rect 3995 3820 3996 3824
rect 3990 3819 3996 3820
rect 111 3818 115 3819
rect 111 3813 115 3814
rect 375 3818 379 3819
rect 375 3813 379 3814
rect 431 3818 435 3819
rect 431 3813 435 3814
rect 495 3818 499 3819
rect 495 3813 499 3814
rect 575 3818 579 3819
rect 575 3813 579 3814
rect 623 3818 627 3819
rect 623 3813 627 3814
rect 719 3818 723 3819
rect 719 3813 723 3814
rect 759 3818 763 3819
rect 759 3813 763 3814
rect 863 3818 867 3819
rect 863 3813 867 3814
rect 895 3818 899 3819
rect 895 3813 899 3814
rect 999 3818 1003 3819
rect 999 3813 1003 3814
rect 1023 3818 1027 3819
rect 1023 3813 1027 3814
rect 1135 3818 1139 3819
rect 1135 3813 1139 3814
rect 1151 3818 1155 3819
rect 1151 3813 1155 3814
rect 1271 3818 1275 3819
rect 1271 3813 1275 3814
rect 1279 3818 1283 3819
rect 1279 3813 1283 3814
rect 1407 3818 1411 3819
rect 1407 3813 1411 3814
rect 1415 3818 1419 3819
rect 1415 3813 1419 3814
rect 1551 3818 1555 3819
rect 1551 3813 1555 3814
rect 2031 3818 2035 3819
rect 2031 3813 2035 3814
rect 112 3798 114 3813
rect 432 3803 434 3813
rect 576 3803 578 3813
rect 720 3803 722 3813
rect 864 3803 866 3813
rect 1000 3803 1002 3813
rect 1136 3803 1138 3813
rect 1272 3803 1274 3813
rect 1408 3803 1410 3813
rect 1552 3803 1554 3813
rect 430 3802 436 3803
rect 430 3798 431 3802
rect 435 3798 436 3802
rect 110 3797 116 3798
rect 430 3797 436 3798
rect 574 3802 580 3803
rect 574 3798 575 3802
rect 579 3798 580 3802
rect 574 3797 580 3798
rect 718 3802 724 3803
rect 718 3798 719 3802
rect 723 3798 724 3802
rect 718 3797 724 3798
rect 862 3802 868 3803
rect 862 3798 863 3802
rect 867 3798 868 3802
rect 862 3797 868 3798
rect 998 3802 1004 3803
rect 998 3798 999 3802
rect 1003 3798 1004 3802
rect 998 3797 1004 3798
rect 1134 3802 1140 3803
rect 1134 3798 1135 3802
rect 1139 3798 1140 3802
rect 1134 3797 1140 3798
rect 1270 3802 1276 3803
rect 1270 3798 1271 3802
rect 1275 3798 1276 3802
rect 1270 3797 1276 3798
rect 1406 3802 1412 3803
rect 1406 3798 1407 3802
rect 1411 3798 1412 3802
rect 1406 3797 1412 3798
rect 1550 3802 1556 3803
rect 1550 3798 1551 3802
rect 1555 3798 1556 3802
rect 2032 3798 2034 3813
rect 1550 3797 1556 3798
rect 2030 3797 2036 3798
rect 110 3793 111 3797
rect 115 3793 116 3797
rect 110 3792 116 3793
rect 2030 3793 2031 3797
rect 2035 3793 2036 3797
rect 2030 3792 2036 3793
rect 2072 3787 2074 3819
rect 2118 3805 2124 3806
rect 2118 3801 2119 3805
rect 2123 3801 2124 3805
rect 2118 3800 2124 3801
rect 2286 3805 2292 3806
rect 2286 3801 2287 3805
rect 2291 3801 2292 3805
rect 2286 3800 2292 3801
rect 2446 3805 2452 3806
rect 2446 3801 2447 3805
rect 2451 3801 2452 3805
rect 2446 3800 2452 3801
rect 2598 3805 2604 3806
rect 2598 3801 2599 3805
rect 2603 3801 2604 3805
rect 2598 3800 2604 3801
rect 2742 3805 2748 3806
rect 2742 3801 2743 3805
rect 2747 3801 2748 3805
rect 2742 3800 2748 3801
rect 2878 3805 2884 3806
rect 2878 3801 2879 3805
rect 2883 3801 2884 3805
rect 2878 3800 2884 3801
rect 3022 3805 3028 3806
rect 3022 3801 3023 3805
rect 3027 3801 3028 3805
rect 3022 3800 3028 3801
rect 3166 3805 3172 3806
rect 3166 3801 3167 3805
rect 3171 3801 3172 3805
rect 3166 3800 3172 3801
rect 2120 3787 2122 3800
rect 2288 3787 2290 3800
rect 2448 3787 2450 3800
rect 2600 3787 2602 3800
rect 2744 3787 2746 3800
rect 2880 3787 2882 3800
rect 3024 3787 3026 3800
rect 3168 3787 3170 3800
rect 3992 3787 3994 3819
rect 2071 3786 2075 3787
rect 2071 3781 2075 3782
rect 2111 3786 2115 3787
rect 2111 3781 2115 3782
rect 2119 3786 2123 3787
rect 2119 3781 2123 3782
rect 2239 3786 2243 3787
rect 2239 3781 2243 3782
rect 2287 3786 2291 3787
rect 2287 3781 2291 3782
rect 2391 3786 2395 3787
rect 2391 3781 2395 3782
rect 2447 3786 2451 3787
rect 2447 3781 2451 3782
rect 2543 3786 2547 3787
rect 2543 3781 2547 3782
rect 2599 3786 2603 3787
rect 2599 3781 2603 3782
rect 2687 3786 2691 3787
rect 2687 3781 2691 3782
rect 2743 3786 2747 3787
rect 2743 3781 2747 3782
rect 2823 3786 2827 3787
rect 2823 3781 2827 3782
rect 2879 3786 2883 3787
rect 2879 3781 2883 3782
rect 2951 3786 2955 3787
rect 2951 3781 2955 3782
rect 3023 3786 3027 3787
rect 3023 3781 3027 3782
rect 3087 3786 3091 3787
rect 3087 3781 3091 3782
rect 3167 3786 3171 3787
rect 3167 3781 3171 3782
rect 3223 3786 3227 3787
rect 3223 3781 3227 3782
rect 3991 3786 3995 3787
rect 3991 3781 3995 3782
rect 110 3780 116 3781
rect 110 3776 111 3780
rect 115 3776 116 3780
rect 110 3775 116 3776
rect 2030 3780 2036 3781
rect 2030 3776 2031 3780
rect 2035 3776 2036 3780
rect 2030 3775 2036 3776
rect 112 3739 114 3775
rect 430 3761 436 3762
rect 430 3757 431 3761
rect 435 3757 436 3761
rect 430 3756 436 3757
rect 574 3761 580 3762
rect 574 3757 575 3761
rect 579 3757 580 3761
rect 574 3756 580 3757
rect 718 3761 724 3762
rect 718 3757 719 3761
rect 723 3757 724 3761
rect 718 3756 724 3757
rect 862 3761 868 3762
rect 862 3757 863 3761
rect 867 3757 868 3761
rect 862 3756 868 3757
rect 998 3761 1004 3762
rect 998 3757 999 3761
rect 1003 3757 1004 3761
rect 998 3756 1004 3757
rect 1134 3761 1140 3762
rect 1134 3757 1135 3761
rect 1139 3757 1140 3761
rect 1134 3756 1140 3757
rect 1270 3761 1276 3762
rect 1270 3757 1271 3761
rect 1275 3757 1276 3761
rect 1270 3756 1276 3757
rect 1406 3761 1412 3762
rect 1406 3757 1407 3761
rect 1411 3757 1412 3761
rect 1406 3756 1412 3757
rect 1550 3761 1556 3762
rect 1550 3757 1551 3761
rect 1555 3757 1556 3761
rect 1550 3756 1556 3757
rect 432 3739 434 3756
rect 576 3739 578 3756
rect 720 3739 722 3756
rect 864 3739 866 3756
rect 1000 3739 1002 3756
rect 1136 3739 1138 3756
rect 1272 3739 1274 3756
rect 1408 3739 1410 3756
rect 1552 3739 1554 3756
rect 2032 3739 2034 3775
rect 2072 3753 2074 3781
rect 2112 3772 2114 3781
rect 2240 3772 2242 3781
rect 2392 3772 2394 3781
rect 2544 3772 2546 3781
rect 2688 3772 2690 3781
rect 2824 3772 2826 3781
rect 2952 3772 2954 3781
rect 3088 3772 3090 3781
rect 3224 3772 3226 3781
rect 2110 3771 2116 3772
rect 2110 3767 2111 3771
rect 2115 3767 2116 3771
rect 2110 3766 2116 3767
rect 2238 3771 2244 3772
rect 2238 3767 2239 3771
rect 2243 3767 2244 3771
rect 2238 3766 2244 3767
rect 2390 3771 2396 3772
rect 2390 3767 2391 3771
rect 2395 3767 2396 3771
rect 2390 3766 2396 3767
rect 2542 3771 2548 3772
rect 2542 3767 2543 3771
rect 2547 3767 2548 3771
rect 2542 3766 2548 3767
rect 2686 3771 2692 3772
rect 2686 3767 2687 3771
rect 2691 3767 2692 3771
rect 2686 3766 2692 3767
rect 2822 3771 2828 3772
rect 2822 3767 2823 3771
rect 2827 3767 2828 3771
rect 2822 3766 2828 3767
rect 2950 3771 2956 3772
rect 2950 3767 2951 3771
rect 2955 3767 2956 3771
rect 2950 3766 2956 3767
rect 3086 3771 3092 3772
rect 3086 3767 3087 3771
rect 3091 3767 3092 3771
rect 3086 3766 3092 3767
rect 3222 3771 3228 3772
rect 3222 3767 3223 3771
rect 3227 3767 3228 3771
rect 3222 3766 3228 3767
rect 3992 3753 3994 3781
rect 2070 3752 2076 3753
rect 2070 3748 2071 3752
rect 2075 3748 2076 3752
rect 2070 3747 2076 3748
rect 3990 3752 3996 3753
rect 3990 3748 3991 3752
rect 3995 3748 3996 3752
rect 3990 3747 3996 3748
rect 111 3738 115 3739
rect 111 3733 115 3734
rect 359 3738 363 3739
rect 359 3733 363 3734
rect 431 3738 435 3739
rect 431 3733 435 3734
rect 495 3738 499 3739
rect 495 3733 499 3734
rect 575 3738 579 3739
rect 575 3733 579 3734
rect 631 3738 635 3739
rect 631 3733 635 3734
rect 719 3738 723 3739
rect 719 3733 723 3734
rect 775 3738 779 3739
rect 775 3733 779 3734
rect 863 3738 867 3739
rect 863 3733 867 3734
rect 919 3738 923 3739
rect 919 3733 923 3734
rect 999 3738 1003 3739
rect 999 3733 1003 3734
rect 1071 3738 1075 3739
rect 1071 3733 1075 3734
rect 1135 3738 1139 3739
rect 1135 3733 1139 3734
rect 1223 3738 1227 3739
rect 1223 3733 1227 3734
rect 1271 3738 1275 3739
rect 1271 3733 1275 3734
rect 1375 3738 1379 3739
rect 1375 3733 1379 3734
rect 1407 3738 1411 3739
rect 1407 3733 1411 3734
rect 1527 3738 1531 3739
rect 1527 3733 1531 3734
rect 1551 3738 1555 3739
rect 1551 3733 1555 3734
rect 2031 3738 2035 3739
rect 2031 3733 2035 3734
rect 2070 3735 2076 3736
rect 112 3705 114 3733
rect 360 3724 362 3733
rect 496 3724 498 3733
rect 632 3724 634 3733
rect 776 3724 778 3733
rect 920 3724 922 3733
rect 1072 3724 1074 3733
rect 1224 3724 1226 3733
rect 1376 3724 1378 3733
rect 1528 3724 1530 3733
rect 358 3723 364 3724
rect 358 3719 359 3723
rect 363 3719 364 3723
rect 358 3718 364 3719
rect 494 3723 500 3724
rect 494 3719 495 3723
rect 499 3719 500 3723
rect 494 3718 500 3719
rect 630 3723 636 3724
rect 630 3719 631 3723
rect 635 3719 636 3723
rect 630 3718 636 3719
rect 774 3723 780 3724
rect 774 3719 775 3723
rect 779 3719 780 3723
rect 774 3718 780 3719
rect 918 3723 924 3724
rect 918 3719 919 3723
rect 923 3719 924 3723
rect 918 3718 924 3719
rect 1070 3723 1076 3724
rect 1070 3719 1071 3723
rect 1075 3719 1076 3723
rect 1070 3718 1076 3719
rect 1222 3723 1228 3724
rect 1222 3719 1223 3723
rect 1227 3719 1228 3723
rect 1222 3718 1228 3719
rect 1374 3723 1380 3724
rect 1374 3719 1375 3723
rect 1379 3719 1380 3723
rect 1374 3718 1380 3719
rect 1526 3723 1532 3724
rect 1526 3719 1527 3723
rect 1531 3719 1532 3723
rect 1526 3718 1532 3719
rect 2032 3705 2034 3733
rect 2070 3731 2071 3735
rect 2075 3731 2076 3735
rect 3990 3735 3996 3736
rect 3990 3731 3991 3735
rect 3995 3731 3996 3735
rect 2070 3730 2076 3731
rect 2110 3730 2116 3731
rect 2072 3707 2074 3730
rect 2110 3726 2111 3730
rect 2115 3726 2116 3730
rect 2110 3725 2116 3726
rect 2238 3730 2244 3731
rect 2238 3726 2239 3730
rect 2243 3726 2244 3730
rect 2238 3725 2244 3726
rect 2390 3730 2396 3731
rect 2390 3726 2391 3730
rect 2395 3726 2396 3730
rect 2390 3725 2396 3726
rect 2542 3730 2548 3731
rect 2542 3726 2543 3730
rect 2547 3726 2548 3730
rect 2542 3725 2548 3726
rect 2686 3730 2692 3731
rect 2686 3726 2687 3730
rect 2691 3726 2692 3730
rect 2686 3725 2692 3726
rect 2822 3730 2828 3731
rect 2822 3726 2823 3730
rect 2827 3726 2828 3730
rect 2822 3725 2828 3726
rect 2950 3730 2956 3731
rect 2950 3726 2951 3730
rect 2955 3726 2956 3730
rect 2950 3725 2956 3726
rect 3086 3730 3092 3731
rect 3086 3726 3087 3730
rect 3091 3726 3092 3730
rect 3086 3725 3092 3726
rect 3222 3730 3228 3731
rect 3990 3730 3996 3731
rect 3222 3726 3223 3730
rect 3227 3726 3228 3730
rect 3222 3725 3228 3726
rect 2112 3707 2114 3725
rect 2240 3707 2242 3725
rect 2392 3707 2394 3725
rect 2544 3707 2546 3725
rect 2688 3707 2690 3725
rect 2824 3707 2826 3725
rect 2952 3707 2954 3725
rect 3088 3707 3090 3725
rect 3224 3707 3226 3725
rect 3992 3707 3994 3730
rect 2071 3706 2075 3707
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 110 3699 116 3700
rect 2030 3704 2036 3705
rect 2030 3700 2031 3704
rect 2035 3700 2036 3704
rect 2071 3701 2075 3702
rect 2111 3706 2115 3707
rect 2111 3701 2115 3702
rect 2239 3706 2243 3707
rect 2239 3701 2243 3702
rect 2295 3706 2299 3707
rect 2295 3701 2299 3702
rect 2391 3706 2395 3707
rect 2391 3701 2395 3702
rect 2487 3706 2491 3707
rect 2487 3701 2491 3702
rect 2543 3706 2547 3707
rect 2543 3701 2547 3702
rect 2671 3706 2675 3707
rect 2671 3701 2675 3702
rect 2687 3706 2691 3707
rect 2687 3701 2691 3702
rect 2823 3706 2827 3707
rect 2823 3701 2827 3702
rect 2847 3706 2851 3707
rect 2847 3701 2851 3702
rect 2951 3706 2955 3707
rect 2951 3701 2955 3702
rect 3015 3706 3019 3707
rect 3015 3701 3019 3702
rect 3087 3706 3091 3707
rect 3087 3701 3091 3702
rect 3183 3706 3187 3707
rect 3183 3701 3187 3702
rect 3223 3706 3227 3707
rect 3223 3701 3227 3702
rect 3359 3706 3363 3707
rect 3359 3701 3363 3702
rect 3991 3706 3995 3707
rect 3991 3701 3995 3702
rect 2030 3699 2036 3700
rect 110 3687 116 3688
rect 110 3683 111 3687
rect 115 3683 116 3687
rect 2030 3687 2036 3688
rect 2030 3683 2031 3687
rect 2035 3683 2036 3687
rect 2072 3686 2074 3701
rect 2112 3691 2114 3701
rect 2296 3691 2298 3701
rect 2488 3691 2490 3701
rect 2672 3691 2674 3701
rect 2848 3691 2850 3701
rect 3016 3691 3018 3701
rect 3184 3691 3186 3701
rect 3360 3691 3362 3701
rect 2110 3690 2116 3691
rect 2110 3686 2111 3690
rect 2115 3686 2116 3690
rect 110 3682 116 3683
rect 358 3682 364 3683
rect 112 3667 114 3682
rect 358 3678 359 3682
rect 363 3678 364 3682
rect 358 3677 364 3678
rect 494 3682 500 3683
rect 494 3678 495 3682
rect 499 3678 500 3682
rect 494 3677 500 3678
rect 630 3682 636 3683
rect 630 3678 631 3682
rect 635 3678 636 3682
rect 630 3677 636 3678
rect 774 3682 780 3683
rect 774 3678 775 3682
rect 779 3678 780 3682
rect 774 3677 780 3678
rect 918 3682 924 3683
rect 918 3678 919 3682
rect 923 3678 924 3682
rect 918 3677 924 3678
rect 1070 3682 1076 3683
rect 1070 3678 1071 3682
rect 1075 3678 1076 3682
rect 1070 3677 1076 3678
rect 1222 3682 1228 3683
rect 1222 3678 1223 3682
rect 1227 3678 1228 3682
rect 1222 3677 1228 3678
rect 1374 3682 1380 3683
rect 1374 3678 1375 3682
rect 1379 3678 1380 3682
rect 1374 3677 1380 3678
rect 1526 3682 1532 3683
rect 2030 3682 2036 3683
rect 2070 3685 2076 3686
rect 2110 3685 2116 3686
rect 2294 3690 2300 3691
rect 2294 3686 2295 3690
rect 2299 3686 2300 3690
rect 2294 3685 2300 3686
rect 2486 3690 2492 3691
rect 2486 3686 2487 3690
rect 2491 3686 2492 3690
rect 2486 3685 2492 3686
rect 2670 3690 2676 3691
rect 2670 3686 2671 3690
rect 2675 3686 2676 3690
rect 2670 3685 2676 3686
rect 2846 3690 2852 3691
rect 2846 3686 2847 3690
rect 2851 3686 2852 3690
rect 2846 3685 2852 3686
rect 3014 3690 3020 3691
rect 3014 3686 3015 3690
rect 3019 3686 3020 3690
rect 3014 3685 3020 3686
rect 3182 3690 3188 3691
rect 3182 3686 3183 3690
rect 3187 3686 3188 3690
rect 3182 3685 3188 3686
rect 3358 3690 3364 3691
rect 3358 3686 3359 3690
rect 3363 3686 3364 3690
rect 3992 3686 3994 3701
rect 3358 3685 3364 3686
rect 3990 3685 3996 3686
rect 1526 3678 1527 3682
rect 1531 3678 1532 3682
rect 1526 3677 1532 3678
rect 360 3667 362 3677
rect 496 3667 498 3677
rect 632 3667 634 3677
rect 776 3667 778 3677
rect 920 3667 922 3677
rect 1072 3667 1074 3677
rect 1224 3667 1226 3677
rect 1376 3667 1378 3677
rect 1528 3667 1530 3677
rect 2032 3667 2034 3682
rect 2070 3681 2071 3685
rect 2075 3681 2076 3685
rect 2070 3680 2076 3681
rect 3990 3681 3991 3685
rect 3995 3681 3996 3685
rect 3990 3680 3996 3681
rect 2070 3668 2076 3669
rect 111 3666 115 3667
rect 111 3661 115 3662
rect 343 3666 347 3667
rect 343 3661 347 3662
rect 359 3666 363 3667
rect 359 3661 363 3662
rect 495 3666 499 3667
rect 495 3661 499 3662
rect 519 3666 523 3667
rect 519 3661 523 3662
rect 631 3666 635 3667
rect 631 3661 635 3662
rect 695 3666 699 3667
rect 695 3661 699 3662
rect 775 3666 779 3667
rect 775 3661 779 3662
rect 863 3666 867 3667
rect 863 3661 867 3662
rect 919 3666 923 3667
rect 919 3661 923 3662
rect 1031 3666 1035 3667
rect 1031 3661 1035 3662
rect 1071 3666 1075 3667
rect 1071 3661 1075 3662
rect 1191 3666 1195 3667
rect 1191 3661 1195 3662
rect 1223 3666 1227 3667
rect 1223 3661 1227 3662
rect 1343 3666 1347 3667
rect 1343 3661 1347 3662
rect 1375 3666 1379 3667
rect 1375 3661 1379 3662
rect 1495 3666 1499 3667
rect 1495 3661 1499 3662
rect 1527 3666 1531 3667
rect 1527 3661 1531 3662
rect 1655 3666 1659 3667
rect 1655 3661 1659 3662
rect 2031 3666 2035 3667
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 3990 3668 3996 3669
rect 3990 3664 3991 3668
rect 3995 3664 3996 3668
rect 3990 3663 3996 3664
rect 2031 3661 2035 3662
rect 112 3646 114 3661
rect 344 3651 346 3661
rect 520 3651 522 3661
rect 696 3651 698 3661
rect 864 3651 866 3661
rect 1032 3651 1034 3661
rect 1192 3651 1194 3661
rect 1344 3651 1346 3661
rect 1496 3651 1498 3661
rect 1656 3651 1658 3661
rect 342 3650 348 3651
rect 342 3646 343 3650
rect 347 3646 348 3650
rect 110 3645 116 3646
rect 342 3645 348 3646
rect 518 3650 524 3651
rect 518 3646 519 3650
rect 523 3646 524 3650
rect 518 3645 524 3646
rect 694 3650 700 3651
rect 694 3646 695 3650
rect 699 3646 700 3650
rect 694 3645 700 3646
rect 862 3650 868 3651
rect 862 3646 863 3650
rect 867 3646 868 3650
rect 862 3645 868 3646
rect 1030 3650 1036 3651
rect 1030 3646 1031 3650
rect 1035 3646 1036 3650
rect 1030 3645 1036 3646
rect 1190 3650 1196 3651
rect 1190 3646 1191 3650
rect 1195 3646 1196 3650
rect 1190 3645 1196 3646
rect 1342 3650 1348 3651
rect 1342 3646 1343 3650
rect 1347 3646 1348 3650
rect 1342 3645 1348 3646
rect 1494 3650 1500 3651
rect 1494 3646 1495 3650
rect 1499 3646 1500 3650
rect 1494 3645 1500 3646
rect 1654 3650 1660 3651
rect 1654 3646 1655 3650
rect 1659 3646 1660 3650
rect 2032 3646 2034 3661
rect 1654 3645 1660 3646
rect 2030 3645 2036 3646
rect 110 3641 111 3645
rect 115 3641 116 3645
rect 110 3640 116 3641
rect 2030 3641 2031 3645
rect 2035 3641 2036 3645
rect 2030 3640 2036 3641
rect 110 3628 116 3629
rect 110 3624 111 3628
rect 115 3624 116 3628
rect 110 3623 116 3624
rect 2030 3628 2036 3629
rect 2030 3624 2031 3628
rect 2035 3624 2036 3628
rect 2072 3627 2074 3663
rect 2110 3649 2116 3650
rect 2110 3645 2111 3649
rect 2115 3645 2116 3649
rect 2110 3644 2116 3645
rect 2294 3649 2300 3650
rect 2294 3645 2295 3649
rect 2299 3645 2300 3649
rect 2294 3644 2300 3645
rect 2486 3649 2492 3650
rect 2486 3645 2487 3649
rect 2491 3645 2492 3649
rect 2486 3644 2492 3645
rect 2670 3649 2676 3650
rect 2670 3645 2671 3649
rect 2675 3645 2676 3649
rect 2670 3644 2676 3645
rect 2846 3649 2852 3650
rect 2846 3645 2847 3649
rect 2851 3645 2852 3649
rect 2846 3644 2852 3645
rect 3014 3649 3020 3650
rect 3014 3645 3015 3649
rect 3019 3645 3020 3649
rect 3014 3644 3020 3645
rect 3182 3649 3188 3650
rect 3182 3645 3183 3649
rect 3187 3645 3188 3649
rect 3182 3644 3188 3645
rect 3358 3649 3364 3650
rect 3358 3645 3359 3649
rect 3363 3645 3364 3649
rect 3358 3644 3364 3645
rect 2112 3627 2114 3644
rect 2296 3627 2298 3644
rect 2488 3627 2490 3644
rect 2672 3627 2674 3644
rect 2848 3627 2850 3644
rect 3016 3627 3018 3644
rect 3184 3627 3186 3644
rect 3360 3627 3362 3644
rect 3992 3627 3994 3663
rect 2030 3623 2036 3624
rect 2071 3626 2075 3627
rect 112 3595 114 3623
rect 342 3609 348 3610
rect 342 3605 343 3609
rect 347 3605 348 3609
rect 342 3604 348 3605
rect 518 3609 524 3610
rect 518 3605 519 3609
rect 523 3605 524 3609
rect 518 3604 524 3605
rect 694 3609 700 3610
rect 694 3605 695 3609
rect 699 3605 700 3609
rect 694 3604 700 3605
rect 862 3609 868 3610
rect 862 3605 863 3609
rect 867 3605 868 3609
rect 862 3604 868 3605
rect 1030 3609 1036 3610
rect 1030 3605 1031 3609
rect 1035 3605 1036 3609
rect 1030 3604 1036 3605
rect 1190 3609 1196 3610
rect 1190 3605 1191 3609
rect 1195 3605 1196 3609
rect 1190 3604 1196 3605
rect 1342 3609 1348 3610
rect 1342 3605 1343 3609
rect 1347 3605 1348 3609
rect 1342 3604 1348 3605
rect 1494 3609 1500 3610
rect 1494 3605 1495 3609
rect 1499 3605 1500 3609
rect 1494 3604 1500 3605
rect 1654 3609 1660 3610
rect 1654 3605 1655 3609
rect 1659 3605 1660 3609
rect 1654 3604 1660 3605
rect 344 3595 346 3604
rect 520 3595 522 3604
rect 696 3595 698 3604
rect 864 3595 866 3604
rect 1032 3595 1034 3604
rect 1192 3595 1194 3604
rect 1344 3595 1346 3604
rect 1496 3595 1498 3604
rect 1656 3595 1658 3604
rect 2032 3595 2034 3623
rect 2071 3621 2075 3622
rect 2111 3626 2115 3627
rect 2111 3621 2115 3622
rect 2295 3626 2299 3627
rect 2295 3621 2299 3622
rect 2487 3626 2491 3627
rect 2487 3621 2491 3622
rect 2495 3626 2499 3627
rect 2495 3621 2499 3622
rect 2671 3626 2675 3627
rect 2671 3621 2675 3622
rect 2687 3626 2691 3627
rect 2687 3621 2691 3622
rect 2847 3626 2851 3627
rect 2847 3621 2851 3622
rect 2863 3626 2867 3627
rect 2863 3621 2867 3622
rect 3015 3626 3019 3627
rect 3015 3621 3019 3622
rect 3023 3626 3027 3627
rect 3023 3621 3027 3622
rect 3167 3626 3171 3627
rect 3167 3621 3171 3622
rect 3183 3626 3187 3627
rect 3183 3621 3187 3622
rect 3303 3626 3307 3627
rect 3303 3621 3307 3622
rect 3359 3626 3363 3627
rect 3359 3621 3363 3622
rect 3431 3626 3435 3627
rect 3431 3621 3435 3622
rect 3551 3626 3555 3627
rect 3551 3621 3555 3622
rect 3671 3626 3675 3627
rect 3671 3621 3675 3622
rect 3791 3626 3795 3627
rect 3791 3621 3795 3622
rect 3895 3626 3899 3627
rect 3895 3621 3899 3622
rect 3991 3626 3995 3627
rect 3991 3621 3995 3622
rect 111 3594 115 3595
rect 111 3589 115 3590
rect 239 3594 243 3595
rect 239 3589 243 3590
rect 343 3594 347 3595
rect 343 3589 347 3590
rect 399 3594 403 3595
rect 399 3589 403 3590
rect 519 3594 523 3595
rect 519 3589 523 3590
rect 551 3594 555 3595
rect 551 3589 555 3590
rect 695 3594 699 3595
rect 695 3589 699 3590
rect 703 3594 707 3595
rect 703 3589 707 3590
rect 855 3594 859 3595
rect 855 3589 859 3590
rect 863 3594 867 3595
rect 863 3589 867 3590
rect 999 3594 1003 3595
rect 999 3589 1003 3590
rect 1031 3594 1035 3595
rect 1031 3589 1035 3590
rect 1135 3594 1139 3595
rect 1135 3589 1139 3590
rect 1191 3594 1195 3595
rect 1191 3589 1195 3590
rect 1263 3594 1267 3595
rect 1263 3589 1267 3590
rect 1343 3594 1347 3595
rect 1343 3589 1347 3590
rect 1383 3594 1387 3595
rect 1383 3589 1387 3590
rect 1495 3594 1499 3595
rect 1495 3589 1499 3590
rect 1607 3594 1611 3595
rect 1607 3589 1611 3590
rect 1655 3594 1659 3595
rect 1655 3589 1659 3590
rect 1719 3594 1723 3595
rect 1719 3589 1723 3590
rect 1831 3594 1835 3595
rect 1831 3589 1835 3590
rect 1935 3594 1939 3595
rect 1935 3589 1939 3590
rect 2031 3594 2035 3595
rect 2072 3593 2074 3621
rect 2112 3612 2114 3621
rect 2296 3612 2298 3621
rect 2496 3612 2498 3621
rect 2688 3612 2690 3621
rect 2864 3612 2866 3621
rect 3024 3612 3026 3621
rect 3168 3612 3170 3621
rect 3304 3612 3306 3621
rect 3432 3612 3434 3621
rect 3552 3612 3554 3621
rect 3672 3612 3674 3621
rect 3792 3612 3794 3621
rect 3896 3612 3898 3621
rect 2110 3611 2116 3612
rect 2110 3607 2111 3611
rect 2115 3607 2116 3611
rect 2110 3606 2116 3607
rect 2294 3611 2300 3612
rect 2294 3607 2295 3611
rect 2299 3607 2300 3611
rect 2294 3606 2300 3607
rect 2494 3611 2500 3612
rect 2494 3607 2495 3611
rect 2499 3607 2500 3611
rect 2494 3606 2500 3607
rect 2686 3611 2692 3612
rect 2686 3607 2687 3611
rect 2691 3607 2692 3611
rect 2686 3606 2692 3607
rect 2862 3611 2868 3612
rect 2862 3607 2863 3611
rect 2867 3607 2868 3611
rect 2862 3606 2868 3607
rect 3022 3611 3028 3612
rect 3022 3607 3023 3611
rect 3027 3607 3028 3611
rect 3022 3606 3028 3607
rect 3166 3611 3172 3612
rect 3166 3607 3167 3611
rect 3171 3607 3172 3611
rect 3166 3606 3172 3607
rect 3302 3611 3308 3612
rect 3302 3607 3303 3611
rect 3307 3607 3308 3611
rect 3302 3606 3308 3607
rect 3430 3611 3436 3612
rect 3430 3607 3431 3611
rect 3435 3607 3436 3611
rect 3430 3606 3436 3607
rect 3550 3611 3556 3612
rect 3550 3607 3551 3611
rect 3555 3607 3556 3611
rect 3550 3606 3556 3607
rect 3670 3611 3676 3612
rect 3670 3607 3671 3611
rect 3675 3607 3676 3611
rect 3670 3606 3676 3607
rect 3790 3611 3796 3612
rect 3790 3607 3791 3611
rect 3795 3607 3796 3611
rect 3790 3606 3796 3607
rect 3894 3611 3900 3612
rect 3894 3607 3895 3611
rect 3899 3607 3900 3611
rect 3894 3606 3900 3607
rect 3992 3593 3994 3621
rect 2031 3589 2035 3590
rect 2070 3592 2076 3593
rect 112 3561 114 3589
rect 240 3580 242 3589
rect 400 3580 402 3589
rect 552 3580 554 3589
rect 704 3580 706 3589
rect 856 3580 858 3589
rect 1000 3580 1002 3589
rect 1136 3580 1138 3589
rect 1264 3580 1266 3589
rect 1384 3580 1386 3589
rect 1496 3580 1498 3589
rect 1608 3580 1610 3589
rect 1720 3580 1722 3589
rect 1832 3580 1834 3589
rect 1936 3580 1938 3589
rect 238 3579 244 3580
rect 238 3575 239 3579
rect 243 3575 244 3579
rect 238 3574 244 3575
rect 398 3579 404 3580
rect 398 3575 399 3579
rect 403 3575 404 3579
rect 398 3574 404 3575
rect 550 3579 556 3580
rect 550 3575 551 3579
rect 555 3575 556 3579
rect 550 3574 556 3575
rect 702 3579 708 3580
rect 702 3575 703 3579
rect 707 3575 708 3579
rect 702 3574 708 3575
rect 854 3579 860 3580
rect 854 3575 855 3579
rect 859 3575 860 3579
rect 854 3574 860 3575
rect 998 3579 1004 3580
rect 998 3575 999 3579
rect 1003 3575 1004 3579
rect 998 3574 1004 3575
rect 1134 3579 1140 3580
rect 1134 3575 1135 3579
rect 1139 3575 1140 3579
rect 1134 3574 1140 3575
rect 1262 3579 1268 3580
rect 1262 3575 1263 3579
rect 1267 3575 1268 3579
rect 1262 3574 1268 3575
rect 1382 3579 1388 3580
rect 1382 3575 1383 3579
rect 1387 3575 1388 3579
rect 1382 3574 1388 3575
rect 1494 3579 1500 3580
rect 1494 3575 1495 3579
rect 1499 3575 1500 3579
rect 1494 3574 1500 3575
rect 1606 3579 1612 3580
rect 1606 3575 1607 3579
rect 1611 3575 1612 3579
rect 1606 3574 1612 3575
rect 1718 3579 1724 3580
rect 1718 3575 1719 3579
rect 1723 3575 1724 3579
rect 1718 3574 1724 3575
rect 1830 3579 1836 3580
rect 1830 3575 1831 3579
rect 1835 3575 1836 3579
rect 1830 3574 1836 3575
rect 1934 3579 1940 3580
rect 1934 3575 1935 3579
rect 1939 3575 1940 3579
rect 1934 3574 1940 3575
rect 2032 3561 2034 3589
rect 2070 3588 2071 3592
rect 2075 3588 2076 3592
rect 2070 3587 2076 3588
rect 3990 3592 3996 3593
rect 3990 3588 3991 3592
rect 3995 3588 3996 3592
rect 3990 3587 3996 3588
rect 2070 3575 2076 3576
rect 2070 3571 2071 3575
rect 2075 3571 2076 3575
rect 3990 3575 3996 3576
rect 3990 3571 3991 3575
rect 3995 3571 3996 3575
rect 2070 3570 2076 3571
rect 2110 3570 2116 3571
rect 110 3560 116 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 2030 3560 2036 3561
rect 2030 3556 2031 3560
rect 2035 3556 2036 3560
rect 2030 3555 2036 3556
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 2030 3543 2036 3544
rect 2072 3543 2074 3570
rect 2110 3566 2111 3570
rect 2115 3566 2116 3570
rect 2110 3565 2116 3566
rect 2294 3570 2300 3571
rect 2294 3566 2295 3570
rect 2299 3566 2300 3570
rect 2294 3565 2300 3566
rect 2494 3570 2500 3571
rect 2494 3566 2495 3570
rect 2499 3566 2500 3570
rect 2494 3565 2500 3566
rect 2686 3570 2692 3571
rect 2686 3566 2687 3570
rect 2691 3566 2692 3570
rect 2686 3565 2692 3566
rect 2862 3570 2868 3571
rect 2862 3566 2863 3570
rect 2867 3566 2868 3570
rect 2862 3565 2868 3566
rect 3022 3570 3028 3571
rect 3022 3566 3023 3570
rect 3027 3566 3028 3570
rect 3022 3565 3028 3566
rect 3166 3570 3172 3571
rect 3166 3566 3167 3570
rect 3171 3566 3172 3570
rect 3166 3565 3172 3566
rect 3302 3570 3308 3571
rect 3302 3566 3303 3570
rect 3307 3566 3308 3570
rect 3302 3565 3308 3566
rect 3430 3570 3436 3571
rect 3430 3566 3431 3570
rect 3435 3566 3436 3570
rect 3430 3565 3436 3566
rect 3550 3570 3556 3571
rect 3550 3566 3551 3570
rect 3555 3566 3556 3570
rect 3550 3565 3556 3566
rect 3670 3570 3676 3571
rect 3670 3566 3671 3570
rect 3675 3566 3676 3570
rect 3670 3565 3676 3566
rect 3790 3570 3796 3571
rect 3790 3566 3791 3570
rect 3795 3566 3796 3570
rect 3790 3565 3796 3566
rect 3894 3570 3900 3571
rect 3990 3570 3996 3571
rect 3894 3566 3895 3570
rect 3899 3566 3900 3570
rect 3894 3565 3900 3566
rect 2112 3543 2114 3565
rect 2296 3543 2298 3565
rect 2496 3543 2498 3565
rect 2688 3543 2690 3565
rect 2864 3543 2866 3565
rect 3024 3543 3026 3565
rect 3168 3543 3170 3565
rect 3304 3543 3306 3565
rect 3432 3543 3434 3565
rect 3552 3543 3554 3565
rect 3672 3543 3674 3565
rect 3792 3543 3794 3565
rect 3896 3543 3898 3565
rect 3992 3543 3994 3570
rect 2030 3539 2031 3543
rect 2035 3539 2036 3543
rect 110 3538 116 3539
rect 238 3538 244 3539
rect 112 3523 114 3538
rect 238 3534 239 3538
rect 243 3534 244 3538
rect 238 3533 244 3534
rect 398 3538 404 3539
rect 398 3534 399 3538
rect 403 3534 404 3538
rect 398 3533 404 3534
rect 550 3538 556 3539
rect 550 3534 551 3538
rect 555 3534 556 3538
rect 550 3533 556 3534
rect 702 3538 708 3539
rect 702 3534 703 3538
rect 707 3534 708 3538
rect 702 3533 708 3534
rect 854 3538 860 3539
rect 854 3534 855 3538
rect 859 3534 860 3538
rect 854 3533 860 3534
rect 998 3538 1004 3539
rect 998 3534 999 3538
rect 1003 3534 1004 3538
rect 998 3533 1004 3534
rect 1134 3538 1140 3539
rect 1134 3534 1135 3538
rect 1139 3534 1140 3538
rect 1134 3533 1140 3534
rect 1262 3538 1268 3539
rect 1262 3534 1263 3538
rect 1267 3534 1268 3538
rect 1262 3533 1268 3534
rect 1382 3538 1388 3539
rect 1382 3534 1383 3538
rect 1387 3534 1388 3538
rect 1382 3533 1388 3534
rect 1494 3538 1500 3539
rect 1494 3534 1495 3538
rect 1499 3534 1500 3538
rect 1494 3533 1500 3534
rect 1606 3538 1612 3539
rect 1606 3534 1607 3538
rect 1611 3534 1612 3538
rect 1606 3533 1612 3534
rect 1718 3538 1724 3539
rect 1718 3534 1719 3538
rect 1723 3534 1724 3538
rect 1718 3533 1724 3534
rect 1830 3538 1836 3539
rect 1830 3534 1831 3538
rect 1835 3534 1836 3538
rect 1830 3533 1836 3534
rect 1934 3538 1940 3539
rect 2030 3538 2036 3539
rect 2071 3542 2075 3543
rect 1934 3534 1935 3538
rect 1939 3534 1940 3538
rect 1934 3533 1940 3534
rect 240 3523 242 3533
rect 400 3523 402 3533
rect 552 3523 554 3533
rect 704 3523 706 3533
rect 856 3523 858 3533
rect 1000 3523 1002 3533
rect 1136 3523 1138 3533
rect 1264 3523 1266 3533
rect 1384 3523 1386 3533
rect 1496 3523 1498 3533
rect 1608 3523 1610 3533
rect 1720 3523 1722 3533
rect 1832 3523 1834 3533
rect 1936 3523 1938 3533
rect 2032 3523 2034 3538
rect 2071 3537 2075 3538
rect 2111 3542 2115 3543
rect 2111 3537 2115 3538
rect 2295 3542 2299 3543
rect 2295 3537 2299 3538
rect 2447 3542 2451 3543
rect 2447 3537 2451 3538
rect 2495 3542 2499 3543
rect 2495 3537 2499 3538
rect 2591 3542 2595 3543
rect 2591 3537 2595 3538
rect 2687 3542 2691 3543
rect 2687 3537 2691 3538
rect 2727 3542 2731 3543
rect 2727 3537 2731 3538
rect 2863 3542 2867 3543
rect 2863 3537 2867 3538
rect 2991 3542 2995 3543
rect 2991 3537 2995 3538
rect 3023 3542 3027 3543
rect 3023 3537 3027 3538
rect 3119 3542 3123 3543
rect 3119 3537 3123 3538
rect 3167 3542 3171 3543
rect 3167 3537 3171 3538
rect 3239 3542 3243 3543
rect 3239 3537 3243 3538
rect 3303 3542 3307 3543
rect 3303 3537 3307 3538
rect 3351 3542 3355 3543
rect 3351 3537 3355 3538
rect 3431 3542 3435 3543
rect 3431 3537 3435 3538
rect 3463 3542 3467 3543
rect 3463 3537 3467 3538
rect 3551 3542 3555 3543
rect 3551 3537 3555 3538
rect 3575 3542 3579 3543
rect 3575 3537 3579 3538
rect 3671 3542 3675 3543
rect 3671 3537 3675 3538
rect 3687 3542 3691 3543
rect 3687 3537 3691 3538
rect 3791 3542 3795 3543
rect 3791 3537 3795 3538
rect 3895 3542 3899 3543
rect 3895 3537 3899 3538
rect 3991 3542 3995 3543
rect 3991 3537 3995 3538
rect 111 3522 115 3523
rect 111 3517 115 3518
rect 151 3522 155 3523
rect 151 3517 155 3518
rect 239 3522 243 3523
rect 239 3517 243 3518
rect 375 3522 379 3523
rect 375 3517 379 3518
rect 399 3522 403 3523
rect 399 3517 403 3518
rect 551 3522 555 3523
rect 551 3517 555 3518
rect 615 3522 619 3523
rect 615 3517 619 3518
rect 703 3522 707 3523
rect 703 3517 707 3518
rect 847 3522 851 3523
rect 847 3517 851 3518
rect 855 3522 859 3523
rect 855 3517 859 3518
rect 999 3522 1003 3523
rect 999 3517 1003 3518
rect 1063 3522 1067 3523
rect 1063 3517 1067 3518
rect 1135 3522 1139 3523
rect 1135 3517 1139 3518
rect 1255 3522 1259 3523
rect 1255 3517 1259 3518
rect 1263 3522 1267 3523
rect 1263 3517 1267 3518
rect 1383 3522 1387 3523
rect 1383 3517 1387 3518
rect 1439 3522 1443 3523
rect 1439 3517 1443 3518
rect 1495 3522 1499 3523
rect 1495 3517 1499 3518
rect 1607 3522 1611 3523
rect 1607 3517 1611 3518
rect 1615 3522 1619 3523
rect 1615 3517 1619 3518
rect 1719 3522 1723 3523
rect 1719 3517 1723 3518
rect 1783 3522 1787 3523
rect 1783 3517 1787 3518
rect 1831 3522 1835 3523
rect 1831 3517 1835 3518
rect 1935 3522 1939 3523
rect 1935 3517 1939 3518
rect 2031 3522 2035 3523
rect 2072 3522 2074 3537
rect 2448 3527 2450 3537
rect 2592 3527 2594 3537
rect 2728 3527 2730 3537
rect 2864 3527 2866 3537
rect 2992 3527 2994 3537
rect 3120 3527 3122 3537
rect 3240 3527 3242 3537
rect 3352 3527 3354 3537
rect 3464 3527 3466 3537
rect 3576 3527 3578 3537
rect 3688 3527 3690 3537
rect 3792 3527 3794 3537
rect 3896 3527 3898 3537
rect 2446 3526 2452 3527
rect 2446 3522 2447 3526
rect 2451 3522 2452 3526
rect 2031 3517 2035 3518
rect 2070 3521 2076 3522
rect 2446 3521 2452 3522
rect 2590 3526 2596 3527
rect 2590 3522 2591 3526
rect 2595 3522 2596 3526
rect 2590 3521 2596 3522
rect 2726 3526 2732 3527
rect 2726 3522 2727 3526
rect 2731 3522 2732 3526
rect 2726 3521 2732 3522
rect 2862 3526 2868 3527
rect 2862 3522 2863 3526
rect 2867 3522 2868 3526
rect 2862 3521 2868 3522
rect 2990 3526 2996 3527
rect 2990 3522 2991 3526
rect 2995 3522 2996 3526
rect 2990 3521 2996 3522
rect 3118 3526 3124 3527
rect 3118 3522 3119 3526
rect 3123 3522 3124 3526
rect 3118 3521 3124 3522
rect 3238 3526 3244 3527
rect 3238 3522 3239 3526
rect 3243 3522 3244 3526
rect 3238 3521 3244 3522
rect 3350 3526 3356 3527
rect 3350 3522 3351 3526
rect 3355 3522 3356 3526
rect 3350 3521 3356 3522
rect 3462 3526 3468 3527
rect 3462 3522 3463 3526
rect 3467 3522 3468 3526
rect 3462 3521 3468 3522
rect 3574 3526 3580 3527
rect 3574 3522 3575 3526
rect 3579 3522 3580 3526
rect 3574 3521 3580 3522
rect 3686 3526 3692 3527
rect 3686 3522 3687 3526
rect 3691 3522 3692 3526
rect 3686 3521 3692 3522
rect 3790 3526 3796 3527
rect 3790 3522 3791 3526
rect 3795 3522 3796 3526
rect 3790 3521 3796 3522
rect 3894 3526 3900 3527
rect 3894 3522 3895 3526
rect 3899 3522 3900 3526
rect 3992 3522 3994 3537
rect 3894 3521 3900 3522
rect 3990 3521 3996 3522
rect 2070 3517 2071 3521
rect 2075 3517 2076 3521
rect 112 3502 114 3517
rect 152 3507 154 3517
rect 376 3507 378 3517
rect 616 3507 618 3517
rect 848 3507 850 3517
rect 1064 3507 1066 3517
rect 1256 3507 1258 3517
rect 1440 3507 1442 3517
rect 1616 3507 1618 3517
rect 1784 3507 1786 3517
rect 1936 3507 1938 3517
rect 150 3506 156 3507
rect 150 3502 151 3506
rect 155 3502 156 3506
rect 110 3501 116 3502
rect 150 3501 156 3502
rect 374 3506 380 3507
rect 374 3502 375 3506
rect 379 3502 380 3506
rect 374 3501 380 3502
rect 614 3506 620 3507
rect 614 3502 615 3506
rect 619 3502 620 3506
rect 614 3501 620 3502
rect 846 3506 852 3507
rect 846 3502 847 3506
rect 851 3502 852 3506
rect 846 3501 852 3502
rect 1062 3506 1068 3507
rect 1062 3502 1063 3506
rect 1067 3502 1068 3506
rect 1062 3501 1068 3502
rect 1254 3506 1260 3507
rect 1254 3502 1255 3506
rect 1259 3502 1260 3506
rect 1254 3501 1260 3502
rect 1438 3506 1444 3507
rect 1438 3502 1439 3506
rect 1443 3502 1444 3506
rect 1438 3501 1444 3502
rect 1614 3506 1620 3507
rect 1614 3502 1615 3506
rect 1619 3502 1620 3506
rect 1614 3501 1620 3502
rect 1782 3506 1788 3507
rect 1782 3502 1783 3506
rect 1787 3502 1788 3506
rect 1782 3501 1788 3502
rect 1934 3506 1940 3507
rect 1934 3502 1935 3506
rect 1939 3502 1940 3506
rect 2032 3502 2034 3517
rect 2070 3516 2076 3517
rect 3990 3517 3991 3521
rect 3995 3517 3996 3521
rect 3990 3516 3996 3517
rect 2070 3504 2076 3505
rect 1934 3501 1940 3502
rect 2030 3501 2036 3502
rect 110 3497 111 3501
rect 115 3497 116 3501
rect 110 3496 116 3497
rect 2030 3497 2031 3501
rect 2035 3497 2036 3501
rect 2070 3500 2071 3504
rect 2075 3500 2076 3504
rect 2070 3499 2076 3500
rect 3990 3504 3996 3505
rect 3990 3500 3991 3504
rect 3995 3500 3996 3504
rect 3990 3499 3996 3500
rect 2030 3496 2036 3497
rect 110 3484 116 3485
rect 110 3480 111 3484
rect 115 3480 116 3484
rect 110 3479 116 3480
rect 2030 3484 2036 3485
rect 2030 3480 2031 3484
rect 2035 3480 2036 3484
rect 2030 3479 2036 3480
rect 112 3427 114 3479
rect 150 3465 156 3466
rect 150 3461 151 3465
rect 155 3461 156 3465
rect 150 3460 156 3461
rect 374 3465 380 3466
rect 374 3461 375 3465
rect 379 3461 380 3465
rect 374 3460 380 3461
rect 614 3465 620 3466
rect 614 3461 615 3465
rect 619 3461 620 3465
rect 614 3460 620 3461
rect 846 3465 852 3466
rect 846 3461 847 3465
rect 851 3461 852 3465
rect 846 3460 852 3461
rect 1062 3465 1068 3466
rect 1062 3461 1063 3465
rect 1067 3461 1068 3465
rect 1062 3460 1068 3461
rect 1254 3465 1260 3466
rect 1254 3461 1255 3465
rect 1259 3461 1260 3465
rect 1254 3460 1260 3461
rect 1438 3465 1444 3466
rect 1438 3461 1439 3465
rect 1443 3461 1444 3465
rect 1438 3460 1444 3461
rect 1614 3465 1620 3466
rect 1614 3461 1615 3465
rect 1619 3461 1620 3465
rect 1614 3460 1620 3461
rect 1782 3465 1788 3466
rect 1782 3461 1783 3465
rect 1787 3461 1788 3465
rect 1782 3460 1788 3461
rect 1934 3465 1940 3466
rect 1934 3461 1935 3465
rect 1939 3461 1940 3465
rect 1934 3460 1940 3461
rect 152 3427 154 3460
rect 376 3427 378 3460
rect 616 3427 618 3460
rect 848 3427 850 3460
rect 1064 3427 1066 3460
rect 1256 3427 1258 3460
rect 1440 3427 1442 3460
rect 1616 3427 1618 3460
rect 1784 3427 1786 3460
rect 1936 3427 1938 3460
rect 2032 3427 2034 3479
rect 2072 3471 2074 3499
rect 2446 3485 2452 3486
rect 2446 3481 2447 3485
rect 2451 3481 2452 3485
rect 2446 3480 2452 3481
rect 2590 3485 2596 3486
rect 2590 3481 2591 3485
rect 2595 3481 2596 3485
rect 2590 3480 2596 3481
rect 2726 3485 2732 3486
rect 2726 3481 2727 3485
rect 2731 3481 2732 3485
rect 2726 3480 2732 3481
rect 2862 3485 2868 3486
rect 2862 3481 2863 3485
rect 2867 3481 2868 3485
rect 2862 3480 2868 3481
rect 2990 3485 2996 3486
rect 2990 3481 2991 3485
rect 2995 3481 2996 3485
rect 2990 3480 2996 3481
rect 3118 3485 3124 3486
rect 3118 3481 3119 3485
rect 3123 3481 3124 3485
rect 3118 3480 3124 3481
rect 3238 3485 3244 3486
rect 3238 3481 3239 3485
rect 3243 3481 3244 3485
rect 3238 3480 3244 3481
rect 3350 3485 3356 3486
rect 3350 3481 3351 3485
rect 3355 3481 3356 3485
rect 3350 3480 3356 3481
rect 3462 3485 3468 3486
rect 3462 3481 3463 3485
rect 3467 3481 3468 3485
rect 3462 3480 3468 3481
rect 3574 3485 3580 3486
rect 3574 3481 3575 3485
rect 3579 3481 3580 3485
rect 3574 3480 3580 3481
rect 3686 3485 3692 3486
rect 3686 3481 3687 3485
rect 3691 3481 3692 3485
rect 3686 3480 3692 3481
rect 3790 3485 3796 3486
rect 3790 3481 3791 3485
rect 3795 3481 3796 3485
rect 3790 3480 3796 3481
rect 3894 3485 3900 3486
rect 3894 3481 3895 3485
rect 3899 3481 3900 3485
rect 3894 3480 3900 3481
rect 2448 3471 2450 3480
rect 2592 3471 2594 3480
rect 2728 3471 2730 3480
rect 2864 3471 2866 3480
rect 2992 3471 2994 3480
rect 3120 3471 3122 3480
rect 3240 3471 3242 3480
rect 3352 3471 3354 3480
rect 3464 3471 3466 3480
rect 3576 3471 3578 3480
rect 3688 3471 3690 3480
rect 3792 3471 3794 3480
rect 3896 3471 3898 3480
rect 3992 3471 3994 3499
rect 2071 3470 2075 3471
rect 2071 3465 2075 3466
rect 2343 3470 2347 3471
rect 2343 3465 2347 3466
rect 2447 3470 2451 3471
rect 2447 3465 2451 3466
rect 2591 3470 2595 3471
rect 2591 3465 2595 3466
rect 2727 3470 2731 3471
rect 2727 3465 2731 3466
rect 2855 3470 2859 3471
rect 2855 3465 2859 3466
rect 2863 3470 2867 3471
rect 2863 3465 2867 3466
rect 2991 3470 2995 3471
rect 2991 3465 2995 3466
rect 3119 3470 3123 3471
rect 3119 3465 3123 3466
rect 3239 3470 3243 3471
rect 3239 3465 3243 3466
rect 3351 3470 3355 3471
rect 3351 3465 3355 3466
rect 3375 3470 3379 3471
rect 3375 3465 3379 3466
rect 3463 3470 3467 3471
rect 3463 3465 3467 3466
rect 3575 3470 3579 3471
rect 3575 3465 3579 3466
rect 3687 3470 3691 3471
rect 3687 3465 3691 3466
rect 3791 3470 3795 3471
rect 3791 3465 3795 3466
rect 3895 3470 3899 3471
rect 3895 3465 3899 3466
rect 3991 3470 3995 3471
rect 3991 3465 3995 3466
rect 2072 3437 2074 3465
rect 2344 3456 2346 3465
rect 2856 3456 2858 3465
rect 3376 3456 3378 3465
rect 3896 3456 3898 3465
rect 2342 3455 2348 3456
rect 2342 3451 2343 3455
rect 2347 3451 2348 3455
rect 2342 3450 2348 3451
rect 2854 3455 2860 3456
rect 2854 3451 2855 3455
rect 2859 3451 2860 3455
rect 2854 3450 2860 3451
rect 3374 3455 3380 3456
rect 3374 3451 3375 3455
rect 3379 3451 3380 3455
rect 3374 3450 3380 3451
rect 3894 3455 3900 3456
rect 3894 3451 3895 3455
rect 3899 3451 3900 3455
rect 3894 3450 3900 3451
rect 3992 3437 3994 3465
rect 2070 3436 2076 3437
rect 2070 3432 2071 3436
rect 2075 3432 2076 3436
rect 2070 3431 2076 3432
rect 3990 3436 3996 3437
rect 3990 3432 3991 3436
rect 3995 3432 3996 3436
rect 3990 3431 3996 3432
rect 111 3426 115 3427
rect 111 3421 115 3422
rect 151 3426 155 3427
rect 151 3421 155 3422
rect 335 3426 339 3427
rect 335 3421 339 3422
rect 375 3426 379 3427
rect 375 3421 379 3422
rect 583 3426 587 3427
rect 583 3421 587 3422
rect 615 3426 619 3427
rect 615 3421 619 3422
rect 847 3426 851 3427
rect 847 3421 851 3422
rect 863 3426 867 3427
rect 863 3421 867 3422
rect 1063 3426 1067 3427
rect 1063 3421 1067 3422
rect 1159 3426 1163 3427
rect 1159 3421 1163 3422
rect 1255 3426 1259 3427
rect 1255 3421 1259 3422
rect 1439 3426 1443 3427
rect 1439 3421 1443 3422
rect 1463 3426 1467 3427
rect 1463 3421 1467 3422
rect 1615 3426 1619 3427
rect 1615 3421 1619 3422
rect 1783 3426 1787 3427
rect 1783 3421 1787 3422
rect 1935 3426 1939 3427
rect 1935 3421 1939 3422
rect 2031 3426 2035 3427
rect 2031 3421 2035 3422
rect 112 3393 114 3421
rect 152 3412 154 3421
rect 336 3412 338 3421
rect 584 3412 586 3421
rect 864 3412 866 3421
rect 1160 3412 1162 3421
rect 1464 3412 1466 3421
rect 150 3411 156 3412
rect 150 3407 151 3411
rect 155 3407 156 3411
rect 150 3406 156 3407
rect 334 3411 340 3412
rect 334 3407 335 3411
rect 339 3407 340 3411
rect 334 3406 340 3407
rect 582 3411 588 3412
rect 582 3407 583 3411
rect 587 3407 588 3411
rect 582 3406 588 3407
rect 862 3411 868 3412
rect 862 3407 863 3411
rect 867 3407 868 3411
rect 862 3406 868 3407
rect 1158 3411 1164 3412
rect 1158 3407 1159 3411
rect 1163 3407 1164 3411
rect 1158 3406 1164 3407
rect 1462 3411 1468 3412
rect 1462 3407 1463 3411
rect 1467 3407 1468 3411
rect 1462 3406 1468 3407
rect 2032 3393 2034 3421
rect 2070 3419 2076 3420
rect 2070 3415 2071 3419
rect 2075 3415 2076 3419
rect 3990 3419 3996 3420
rect 3990 3415 3991 3419
rect 3995 3415 3996 3419
rect 2070 3414 2076 3415
rect 2342 3414 2348 3415
rect 2072 3395 2074 3414
rect 2342 3410 2343 3414
rect 2347 3410 2348 3414
rect 2342 3409 2348 3410
rect 2854 3414 2860 3415
rect 2854 3410 2855 3414
rect 2859 3410 2860 3414
rect 2854 3409 2860 3410
rect 3374 3414 3380 3415
rect 3374 3410 3375 3414
rect 3379 3410 3380 3414
rect 3374 3409 3380 3410
rect 3894 3414 3900 3415
rect 3990 3414 3996 3415
rect 3894 3410 3895 3414
rect 3899 3410 3900 3414
rect 3894 3409 3900 3410
rect 2344 3395 2346 3409
rect 2856 3395 2858 3409
rect 3376 3395 3378 3409
rect 3896 3395 3898 3409
rect 3992 3395 3994 3414
rect 2071 3394 2075 3395
rect 110 3392 116 3393
rect 110 3388 111 3392
rect 115 3388 116 3392
rect 110 3387 116 3388
rect 2030 3392 2036 3393
rect 2030 3388 2031 3392
rect 2035 3388 2036 3392
rect 2071 3389 2075 3390
rect 2183 3394 2187 3395
rect 2183 3389 2187 3390
rect 2343 3394 2347 3395
rect 2343 3389 2347 3390
rect 2583 3394 2587 3395
rect 2583 3389 2587 3390
rect 2855 3394 2859 3395
rect 2855 3389 2859 3390
rect 3007 3394 3011 3395
rect 3007 3389 3011 3390
rect 3375 3394 3379 3395
rect 3375 3389 3379 3390
rect 3447 3394 3451 3395
rect 3447 3389 3451 3390
rect 3895 3394 3899 3395
rect 3895 3389 3899 3390
rect 3991 3394 3995 3395
rect 3991 3389 3995 3390
rect 2030 3387 2036 3388
rect 110 3375 116 3376
rect 110 3371 111 3375
rect 115 3371 116 3375
rect 2030 3375 2036 3376
rect 2030 3371 2031 3375
rect 2035 3371 2036 3375
rect 2072 3374 2074 3389
rect 2184 3379 2186 3389
rect 2584 3379 2586 3389
rect 3008 3379 3010 3389
rect 3448 3379 3450 3389
rect 3896 3379 3898 3389
rect 2182 3378 2188 3379
rect 2182 3374 2183 3378
rect 2187 3374 2188 3378
rect 110 3370 116 3371
rect 150 3370 156 3371
rect 112 3347 114 3370
rect 150 3366 151 3370
rect 155 3366 156 3370
rect 150 3365 156 3366
rect 334 3370 340 3371
rect 334 3366 335 3370
rect 339 3366 340 3370
rect 334 3365 340 3366
rect 582 3370 588 3371
rect 582 3366 583 3370
rect 587 3366 588 3370
rect 582 3365 588 3366
rect 862 3370 868 3371
rect 862 3366 863 3370
rect 867 3366 868 3370
rect 862 3365 868 3366
rect 1158 3370 1164 3371
rect 1158 3366 1159 3370
rect 1163 3366 1164 3370
rect 1158 3365 1164 3366
rect 1462 3370 1468 3371
rect 2030 3370 2036 3371
rect 2070 3373 2076 3374
rect 2182 3373 2188 3374
rect 2582 3378 2588 3379
rect 2582 3374 2583 3378
rect 2587 3374 2588 3378
rect 2582 3373 2588 3374
rect 3006 3378 3012 3379
rect 3006 3374 3007 3378
rect 3011 3374 3012 3378
rect 3006 3373 3012 3374
rect 3446 3378 3452 3379
rect 3446 3374 3447 3378
rect 3451 3374 3452 3378
rect 3446 3373 3452 3374
rect 3894 3378 3900 3379
rect 3894 3374 3895 3378
rect 3899 3374 3900 3378
rect 3992 3374 3994 3389
rect 3894 3373 3900 3374
rect 3990 3373 3996 3374
rect 1462 3366 1463 3370
rect 1467 3366 1468 3370
rect 1462 3365 1468 3366
rect 152 3347 154 3365
rect 336 3347 338 3365
rect 584 3347 586 3365
rect 864 3347 866 3365
rect 1160 3347 1162 3365
rect 1464 3347 1466 3365
rect 2032 3347 2034 3370
rect 2070 3369 2071 3373
rect 2075 3369 2076 3373
rect 2070 3368 2076 3369
rect 3990 3369 3991 3373
rect 3995 3369 3996 3373
rect 3990 3368 3996 3369
rect 2070 3356 2076 3357
rect 2070 3352 2071 3356
rect 2075 3352 2076 3356
rect 2070 3351 2076 3352
rect 3990 3356 3996 3357
rect 3990 3352 3991 3356
rect 3995 3352 3996 3356
rect 3990 3351 3996 3352
rect 111 3346 115 3347
rect 111 3341 115 3342
rect 151 3346 155 3347
rect 151 3341 155 3342
rect 287 3346 291 3347
rect 287 3341 291 3342
rect 335 3346 339 3347
rect 335 3341 339 3342
rect 463 3346 467 3347
rect 463 3341 467 3342
rect 583 3346 587 3347
rect 583 3341 587 3342
rect 639 3346 643 3347
rect 639 3341 643 3342
rect 815 3346 819 3347
rect 815 3341 819 3342
rect 863 3346 867 3347
rect 863 3341 867 3342
rect 991 3346 995 3347
rect 991 3341 995 3342
rect 1159 3346 1163 3347
rect 1159 3341 1163 3342
rect 1319 3346 1323 3347
rect 1319 3341 1323 3342
rect 1463 3346 1467 3347
rect 1463 3341 1467 3342
rect 1487 3346 1491 3347
rect 1487 3341 1491 3342
rect 1655 3346 1659 3347
rect 1655 3341 1659 3342
rect 2031 3346 2035 3347
rect 2031 3341 2035 3342
rect 112 3326 114 3341
rect 152 3331 154 3341
rect 288 3331 290 3341
rect 464 3331 466 3341
rect 640 3331 642 3341
rect 816 3331 818 3341
rect 992 3331 994 3341
rect 1160 3331 1162 3341
rect 1320 3331 1322 3341
rect 1488 3331 1490 3341
rect 1656 3331 1658 3341
rect 150 3330 156 3331
rect 150 3326 151 3330
rect 155 3326 156 3330
rect 110 3325 116 3326
rect 150 3325 156 3326
rect 286 3330 292 3331
rect 286 3326 287 3330
rect 291 3326 292 3330
rect 286 3325 292 3326
rect 462 3330 468 3331
rect 462 3326 463 3330
rect 467 3326 468 3330
rect 462 3325 468 3326
rect 638 3330 644 3331
rect 638 3326 639 3330
rect 643 3326 644 3330
rect 638 3325 644 3326
rect 814 3330 820 3331
rect 814 3326 815 3330
rect 819 3326 820 3330
rect 814 3325 820 3326
rect 990 3330 996 3331
rect 990 3326 991 3330
rect 995 3326 996 3330
rect 990 3325 996 3326
rect 1158 3330 1164 3331
rect 1158 3326 1159 3330
rect 1163 3326 1164 3330
rect 1158 3325 1164 3326
rect 1318 3330 1324 3331
rect 1318 3326 1319 3330
rect 1323 3326 1324 3330
rect 1318 3325 1324 3326
rect 1486 3330 1492 3331
rect 1486 3326 1487 3330
rect 1491 3326 1492 3330
rect 1486 3325 1492 3326
rect 1654 3330 1660 3331
rect 1654 3326 1655 3330
rect 1659 3326 1660 3330
rect 2032 3326 2034 3341
rect 1654 3325 1660 3326
rect 2030 3325 2036 3326
rect 110 3321 111 3325
rect 115 3321 116 3325
rect 110 3320 116 3321
rect 2030 3321 2031 3325
rect 2035 3321 2036 3325
rect 2030 3320 2036 3321
rect 110 3308 116 3309
rect 110 3304 111 3308
rect 115 3304 116 3308
rect 110 3303 116 3304
rect 2030 3308 2036 3309
rect 2030 3304 2031 3308
rect 2035 3304 2036 3308
rect 2072 3307 2074 3351
rect 2182 3337 2188 3338
rect 2182 3333 2183 3337
rect 2187 3333 2188 3337
rect 2182 3332 2188 3333
rect 2582 3337 2588 3338
rect 2582 3333 2583 3337
rect 2587 3333 2588 3337
rect 2582 3332 2588 3333
rect 3006 3337 3012 3338
rect 3006 3333 3007 3337
rect 3011 3333 3012 3337
rect 3006 3332 3012 3333
rect 3446 3337 3452 3338
rect 3446 3333 3447 3337
rect 3451 3333 3452 3337
rect 3446 3332 3452 3333
rect 3894 3337 3900 3338
rect 3894 3333 3895 3337
rect 3899 3333 3900 3337
rect 3894 3332 3900 3333
rect 2184 3307 2186 3332
rect 2584 3307 2586 3332
rect 3008 3307 3010 3332
rect 3448 3307 3450 3332
rect 3896 3307 3898 3332
rect 3992 3307 3994 3351
rect 2030 3303 2036 3304
rect 2071 3306 2075 3307
rect 112 3263 114 3303
rect 150 3289 156 3290
rect 150 3285 151 3289
rect 155 3285 156 3289
rect 150 3284 156 3285
rect 286 3289 292 3290
rect 286 3285 287 3289
rect 291 3285 292 3289
rect 286 3284 292 3285
rect 462 3289 468 3290
rect 462 3285 463 3289
rect 467 3285 468 3289
rect 462 3284 468 3285
rect 638 3289 644 3290
rect 638 3285 639 3289
rect 643 3285 644 3289
rect 638 3284 644 3285
rect 814 3289 820 3290
rect 814 3285 815 3289
rect 819 3285 820 3289
rect 814 3284 820 3285
rect 990 3289 996 3290
rect 990 3285 991 3289
rect 995 3285 996 3289
rect 990 3284 996 3285
rect 1158 3289 1164 3290
rect 1158 3285 1159 3289
rect 1163 3285 1164 3289
rect 1158 3284 1164 3285
rect 1318 3289 1324 3290
rect 1318 3285 1319 3289
rect 1323 3285 1324 3289
rect 1318 3284 1324 3285
rect 1486 3289 1492 3290
rect 1486 3285 1487 3289
rect 1491 3285 1492 3289
rect 1486 3284 1492 3285
rect 1654 3289 1660 3290
rect 1654 3285 1655 3289
rect 1659 3285 1660 3289
rect 1654 3284 1660 3285
rect 152 3263 154 3284
rect 288 3263 290 3284
rect 464 3263 466 3284
rect 640 3263 642 3284
rect 816 3263 818 3284
rect 992 3263 994 3284
rect 1160 3263 1162 3284
rect 1320 3263 1322 3284
rect 1488 3263 1490 3284
rect 1656 3263 1658 3284
rect 2032 3263 2034 3303
rect 2071 3301 2075 3302
rect 2111 3306 2115 3307
rect 2111 3301 2115 3302
rect 2183 3306 2187 3307
rect 2183 3301 2187 3302
rect 2295 3306 2299 3307
rect 2295 3301 2299 3302
rect 2503 3306 2507 3307
rect 2503 3301 2507 3302
rect 2583 3306 2587 3307
rect 2583 3301 2587 3302
rect 2703 3306 2707 3307
rect 2703 3301 2707 3302
rect 2895 3306 2899 3307
rect 2895 3301 2899 3302
rect 3007 3306 3011 3307
rect 3007 3301 3011 3302
rect 3071 3306 3075 3307
rect 3071 3301 3075 3302
rect 3231 3306 3235 3307
rect 3231 3301 3235 3302
rect 3375 3306 3379 3307
rect 3375 3301 3379 3302
rect 3447 3306 3451 3307
rect 3447 3301 3451 3302
rect 3511 3306 3515 3307
rect 3511 3301 3515 3302
rect 3647 3306 3651 3307
rect 3647 3301 3651 3302
rect 3783 3306 3787 3307
rect 3783 3301 3787 3302
rect 3895 3306 3899 3307
rect 3895 3301 3899 3302
rect 3991 3306 3995 3307
rect 3991 3301 3995 3302
rect 2072 3273 2074 3301
rect 2112 3292 2114 3301
rect 2296 3292 2298 3301
rect 2504 3292 2506 3301
rect 2704 3292 2706 3301
rect 2896 3292 2898 3301
rect 3072 3292 3074 3301
rect 3232 3292 3234 3301
rect 3376 3292 3378 3301
rect 3512 3292 3514 3301
rect 3648 3292 3650 3301
rect 3784 3292 3786 3301
rect 3896 3292 3898 3301
rect 2110 3291 2116 3292
rect 2110 3287 2111 3291
rect 2115 3287 2116 3291
rect 2110 3286 2116 3287
rect 2294 3291 2300 3292
rect 2294 3287 2295 3291
rect 2299 3287 2300 3291
rect 2294 3286 2300 3287
rect 2502 3291 2508 3292
rect 2502 3287 2503 3291
rect 2507 3287 2508 3291
rect 2502 3286 2508 3287
rect 2702 3291 2708 3292
rect 2702 3287 2703 3291
rect 2707 3287 2708 3291
rect 2702 3286 2708 3287
rect 2894 3291 2900 3292
rect 2894 3287 2895 3291
rect 2899 3287 2900 3291
rect 2894 3286 2900 3287
rect 3070 3291 3076 3292
rect 3070 3287 3071 3291
rect 3075 3287 3076 3291
rect 3070 3286 3076 3287
rect 3230 3291 3236 3292
rect 3230 3287 3231 3291
rect 3235 3287 3236 3291
rect 3230 3286 3236 3287
rect 3374 3291 3380 3292
rect 3374 3287 3375 3291
rect 3379 3287 3380 3291
rect 3374 3286 3380 3287
rect 3510 3291 3516 3292
rect 3510 3287 3511 3291
rect 3515 3287 3516 3291
rect 3510 3286 3516 3287
rect 3646 3291 3652 3292
rect 3646 3287 3647 3291
rect 3651 3287 3652 3291
rect 3646 3286 3652 3287
rect 3782 3291 3788 3292
rect 3782 3287 3783 3291
rect 3787 3287 3788 3291
rect 3782 3286 3788 3287
rect 3894 3291 3900 3292
rect 3894 3287 3895 3291
rect 3899 3287 3900 3291
rect 3894 3286 3900 3287
rect 3992 3273 3994 3301
rect 2070 3272 2076 3273
rect 2070 3268 2071 3272
rect 2075 3268 2076 3272
rect 2070 3267 2076 3268
rect 3990 3272 3996 3273
rect 3990 3268 3991 3272
rect 3995 3268 3996 3272
rect 3990 3267 3996 3268
rect 111 3262 115 3263
rect 111 3257 115 3258
rect 151 3262 155 3263
rect 151 3257 155 3258
rect 287 3262 291 3263
rect 287 3257 291 3258
rect 295 3262 299 3263
rect 295 3257 299 3258
rect 463 3262 467 3263
rect 463 3257 467 3258
rect 479 3262 483 3263
rect 479 3257 483 3258
rect 639 3262 643 3263
rect 639 3257 643 3258
rect 671 3262 675 3263
rect 671 3257 675 3258
rect 815 3262 819 3263
rect 815 3257 819 3258
rect 863 3262 867 3263
rect 863 3257 867 3258
rect 991 3262 995 3263
rect 991 3257 995 3258
rect 1055 3262 1059 3263
rect 1055 3257 1059 3258
rect 1159 3262 1163 3263
rect 1159 3257 1163 3258
rect 1247 3262 1251 3263
rect 1247 3257 1251 3258
rect 1319 3262 1323 3263
rect 1319 3257 1323 3258
rect 1431 3262 1435 3263
rect 1431 3257 1435 3258
rect 1487 3262 1491 3263
rect 1487 3257 1491 3258
rect 1615 3262 1619 3263
rect 1615 3257 1619 3258
rect 1655 3262 1659 3263
rect 1655 3257 1659 3258
rect 1807 3262 1811 3263
rect 1807 3257 1811 3258
rect 2031 3262 2035 3263
rect 2031 3257 2035 3258
rect 112 3229 114 3257
rect 152 3248 154 3257
rect 296 3248 298 3257
rect 480 3248 482 3257
rect 672 3248 674 3257
rect 864 3248 866 3257
rect 1056 3248 1058 3257
rect 1248 3248 1250 3257
rect 1432 3248 1434 3257
rect 1616 3248 1618 3257
rect 1808 3248 1810 3257
rect 150 3247 156 3248
rect 150 3243 151 3247
rect 155 3243 156 3247
rect 150 3242 156 3243
rect 294 3247 300 3248
rect 294 3243 295 3247
rect 299 3243 300 3247
rect 294 3242 300 3243
rect 478 3247 484 3248
rect 478 3243 479 3247
rect 483 3243 484 3247
rect 478 3242 484 3243
rect 670 3247 676 3248
rect 670 3243 671 3247
rect 675 3243 676 3247
rect 670 3242 676 3243
rect 862 3247 868 3248
rect 862 3243 863 3247
rect 867 3243 868 3247
rect 862 3242 868 3243
rect 1054 3247 1060 3248
rect 1054 3243 1055 3247
rect 1059 3243 1060 3247
rect 1054 3242 1060 3243
rect 1246 3247 1252 3248
rect 1246 3243 1247 3247
rect 1251 3243 1252 3247
rect 1246 3242 1252 3243
rect 1430 3247 1436 3248
rect 1430 3243 1431 3247
rect 1435 3243 1436 3247
rect 1430 3242 1436 3243
rect 1614 3247 1620 3248
rect 1614 3243 1615 3247
rect 1619 3243 1620 3247
rect 1614 3242 1620 3243
rect 1806 3247 1812 3248
rect 1806 3243 1807 3247
rect 1811 3243 1812 3247
rect 1806 3242 1812 3243
rect 2032 3229 2034 3257
rect 2070 3255 2076 3256
rect 2070 3251 2071 3255
rect 2075 3251 2076 3255
rect 3990 3255 3996 3256
rect 3990 3251 3991 3255
rect 3995 3251 3996 3255
rect 2070 3250 2076 3251
rect 2110 3250 2116 3251
rect 2072 3235 2074 3250
rect 2110 3246 2111 3250
rect 2115 3246 2116 3250
rect 2110 3245 2116 3246
rect 2294 3250 2300 3251
rect 2294 3246 2295 3250
rect 2299 3246 2300 3250
rect 2294 3245 2300 3246
rect 2502 3250 2508 3251
rect 2502 3246 2503 3250
rect 2507 3246 2508 3250
rect 2502 3245 2508 3246
rect 2702 3250 2708 3251
rect 2702 3246 2703 3250
rect 2707 3246 2708 3250
rect 2702 3245 2708 3246
rect 2894 3250 2900 3251
rect 2894 3246 2895 3250
rect 2899 3246 2900 3250
rect 2894 3245 2900 3246
rect 3070 3250 3076 3251
rect 3070 3246 3071 3250
rect 3075 3246 3076 3250
rect 3070 3245 3076 3246
rect 3230 3250 3236 3251
rect 3230 3246 3231 3250
rect 3235 3246 3236 3250
rect 3230 3245 3236 3246
rect 3374 3250 3380 3251
rect 3374 3246 3375 3250
rect 3379 3246 3380 3250
rect 3374 3245 3380 3246
rect 3510 3250 3516 3251
rect 3510 3246 3511 3250
rect 3515 3246 3516 3250
rect 3510 3245 3516 3246
rect 3646 3250 3652 3251
rect 3646 3246 3647 3250
rect 3651 3246 3652 3250
rect 3646 3245 3652 3246
rect 3782 3250 3788 3251
rect 3782 3246 3783 3250
rect 3787 3246 3788 3250
rect 3782 3245 3788 3246
rect 3894 3250 3900 3251
rect 3990 3250 3996 3251
rect 3894 3246 3895 3250
rect 3899 3246 3900 3250
rect 3894 3245 3900 3246
rect 2112 3235 2114 3245
rect 2296 3235 2298 3245
rect 2504 3235 2506 3245
rect 2704 3235 2706 3245
rect 2896 3235 2898 3245
rect 3072 3235 3074 3245
rect 3232 3235 3234 3245
rect 3376 3235 3378 3245
rect 3512 3235 3514 3245
rect 3648 3235 3650 3245
rect 3784 3235 3786 3245
rect 3896 3235 3898 3245
rect 3992 3235 3994 3250
rect 2071 3234 2075 3235
rect 2071 3229 2075 3230
rect 2111 3234 2115 3235
rect 2111 3229 2115 3230
rect 2239 3234 2243 3235
rect 2239 3229 2243 3230
rect 2295 3234 2299 3235
rect 2295 3229 2299 3230
rect 2399 3234 2403 3235
rect 2399 3229 2403 3230
rect 2503 3234 2507 3235
rect 2503 3229 2507 3230
rect 2559 3234 2563 3235
rect 2559 3229 2563 3230
rect 2703 3234 2707 3235
rect 2703 3229 2707 3230
rect 2719 3234 2723 3235
rect 2719 3229 2723 3230
rect 2879 3234 2883 3235
rect 2879 3229 2883 3230
rect 2895 3234 2899 3235
rect 2895 3229 2899 3230
rect 3031 3234 3035 3235
rect 3031 3229 3035 3230
rect 3071 3234 3075 3235
rect 3071 3229 3075 3230
rect 3167 3234 3171 3235
rect 3167 3229 3171 3230
rect 3231 3234 3235 3235
rect 3231 3229 3235 3230
rect 3303 3234 3307 3235
rect 3303 3229 3307 3230
rect 3375 3234 3379 3235
rect 3375 3229 3379 3230
rect 3431 3234 3435 3235
rect 3431 3229 3435 3230
rect 3511 3234 3515 3235
rect 3511 3229 3515 3230
rect 3551 3234 3555 3235
rect 3551 3229 3555 3230
rect 3647 3234 3651 3235
rect 3647 3229 3651 3230
rect 3671 3234 3675 3235
rect 3671 3229 3675 3230
rect 3783 3234 3787 3235
rect 3783 3229 3787 3230
rect 3791 3234 3795 3235
rect 3791 3229 3795 3230
rect 3895 3234 3899 3235
rect 3895 3229 3899 3230
rect 3991 3234 3995 3235
rect 3991 3229 3995 3230
rect 110 3228 116 3229
rect 110 3224 111 3228
rect 115 3224 116 3228
rect 110 3223 116 3224
rect 2030 3228 2036 3229
rect 2030 3224 2031 3228
rect 2035 3224 2036 3228
rect 2030 3223 2036 3224
rect 2072 3214 2074 3229
rect 2112 3219 2114 3229
rect 2240 3219 2242 3229
rect 2400 3219 2402 3229
rect 2560 3219 2562 3229
rect 2720 3219 2722 3229
rect 2880 3219 2882 3229
rect 3032 3219 3034 3229
rect 3168 3219 3170 3229
rect 3304 3219 3306 3229
rect 3432 3219 3434 3229
rect 3552 3219 3554 3229
rect 3672 3219 3674 3229
rect 3792 3219 3794 3229
rect 3896 3219 3898 3229
rect 2110 3218 2116 3219
rect 2110 3214 2111 3218
rect 2115 3214 2116 3218
rect 2070 3213 2076 3214
rect 2110 3213 2116 3214
rect 2238 3218 2244 3219
rect 2238 3214 2239 3218
rect 2243 3214 2244 3218
rect 2238 3213 2244 3214
rect 2398 3218 2404 3219
rect 2398 3214 2399 3218
rect 2403 3214 2404 3218
rect 2398 3213 2404 3214
rect 2558 3218 2564 3219
rect 2558 3214 2559 3218
rect 2563 3214 2564 3218
rect 2558 3213 2564 3214
rect 2718 3218 2724 3219
rect 2718 3214 2719 3218
rect 2723 3214 2724 3218
rect 2718 3213 2724 3214
rect 2878 3218 2884 3219
rect 2878 3214 2879 3218
rect 2883 3214 2884 3218
rect 2878 3213 2884 3214
rect 3030 3218 3036 3219
rect 3030 3214 3031 3218
rect 3035 3214 3036 3218
rect 3030 3213 3036 3214
rect 3166 3218 3172 3219
rect 3166 3214 3167 3218
rect 3171 3214 3172 3218
rect 3166 3213 3172 3214
rect 3302 3218 3308 3219
rect 3302 3214 3303 3218
rect 3307 3214 3308 3218
rect 3302 3213 3308 3214
rect 3430 3218 3436 3219
rect 3430 3214 3431 3218
rect 3435 3214 3436 3218
rect 3430 3213 3436 3214
rect 3550 3218 3556 3219
rect 3550 3214 3551 3218
rect 3555 3214 3556 3218
rect 3550 3213 3556 3214
rect 3670 3218 3676 3219
rect 3670 3214 3671 3218
rect 3675 3214 3676 3218
rect 3670 3213 3676 3214
rect 3790 3218 3796 3219
rect 3790 3214 3791 3218
rect 3795 3214 3796 3218
rect 3790 3213 3796 3214
rect 3894 3218 3900 3219
rect 3894 3214 3895 3218
rect 3899 3214 3900 3218
rect 3992 3214 3994 3229
rect 3894 3213 3900 3214
rect 3990 3213 3996 3214
rect 110 3211 116 3212
rect 110 3207 111 3211
rect 115 3207 116 3211
rect 2030 3211 2036 3212
rect 2030 3207 2031 3211
rect 2035 3207 2036 3211
rect 2070 3209 2071 3213
rect 2075 3209 2076 3213
rect 2070 3208 2076 3209
rect 3990 3209 3991 3213
rect 3995 3209 3996 3213
rect 3990 3208 3996 3209
rect 110 3206 116 3207
rect 150 3206 156 3207
rect 112 3179 114 3206
rect 150 3202 151 3206
rect 155 3202 156 3206
rect 150 3201 156 3202
rect 294 3206 300 3207
rect 294 3202 295 3206
rect 299 3202 300 3206
rect 294 3201 300 3202
rect 478 3206 484 3207
rect 478 3202 479 3206
rect 483 3202 484 3206
rect 478 3201 484 3202
rect 670 3206 676 3207
rect 670 3202 671 3206
rect 675 3202 676 3206
rect 670 3201 676 3202
rect 862 3206 868 3207
rect 862 3202 863 3206
rect 867 3202 868 3206
rect 862 3201 868 3202
rect 1054 3206 1060 3207
rect 1054 3202 1055 3206
rect 1059 3202 1060 3206
rect 1054 3201 1060 3202
rect 1246 3206 1252 3207
rect 1246 3202 1247 3206
rect 1251 3202 1252 3206
rect 1246 3201 1252 3202
rect 1430 3206 1436 3207
rect 1430 3202 1431 3206
rect 1435 3202 1436 3206
rect 1430 3201 1436 3202
rect 1614 3206 1620 3207
rect 1614 3202 1615 3206
rect 1619 3202 1620 3206
rect 1614 3201 1620 3202
rect 1806 3206 1812 3207
rect 2030 3206 2036 3207
rect 1806 3202 1807 3206
rect 1811 3202 1812 3206
rect 1806 3201 1812 3202
rect 152 3179 154 3201
rect 296 3179 298 3201
rect 480 3179 482 3201
rect 672 3179 674 3201
rect 864 3179 866 3201
rect 1056 3179 1058 3201
rect 1248 3179 1250 3201
rect 1432 3179 1434 3201
rect 1616 3179 1618 3201
rect 1808 3179 1810 3201
rect 2032 3179 2034 3206
rect 2070 3196 2076 3197
rect 2070 3192 2071 3196
rect 2075 3192 2076 3196
rect 2070 3191 2076 3192
rect 3990 3196 3996 3197
rect 3990 3192 3991 3196
rect 3995 3192 3996 3196
rect 3990 3191 3996 3192
rect 111 3178 115 3179
rect 111 3173 115 3174
rect 151 3178 155 3179
rect 151 3173 155 3174
rect 287 3178 291 3179
rect 287 3173 291 3174
rect 295 3178 299 3179
rect 295 3173 299 3174
rect 423 3178 427 3179
rect 423 3173 427 3174
rect 479 3178 483 3179
rect 479 3173 483 3174
rect 567 3178 571 3179
rect 567 3173 571 3174
rect 671 3178 675 3179
rect 671 3173 675 3174
rect 727 3178 731 3179
rect 727 3173 731 3174
rect 863 3178 867 3179
rect 863 3173 867 3174
rect 903 3178 907 3179
rect 903 3173 907 3174
rect 1055 3178 1059 3179
rect 1055 3173 1059 3174
rect 1095 3178 1099 3179
rect 1095 3173 1099 3174
rect 1247 3178 1251 3179
rect 1247 3173 1251 3174
rect 1295 3178 1299 3179
rect 1295 3173 1299 3174
rect 1431 3178 1435 3179
rect 1431 3173 1435 3174
rect 1495 3178 1499 3179
rect 1495 3173 1499 3174
rect 1615 3178 1619 3179
rect 1615 3173 1619 3174
rect 1703 3178 1707 3179
rect 1703 3173 1707 3174
rect 1807 3178 1811 3179
rect 1807 3173 1811 3174
rect 1919 3178 1923 3179
rect 1919 3173 1923 3174
rect 2031 3178 2035 3179
rect 2031 3173 2035 3174
rect 112 3158 114 3173
rect 288 3163 290 3173
rect 424 3163 426 3173
rect 568 3163 570 3173
rect 728 3163 730 3173
rect 904 3163 906 3173
rect 1096 3163 1098 3173
rect 1296 3163 1298 3173
rect 1496 3163 1498 3173
rect 1704 3163 1706 3173
rect 1920 3163 1922 3173
rect 286 3162 292 3163
rect 286 3158 287 3162
rect 291 3158 292 3162
rect 110 3157 116 3158
rect 286 3157 292 3158
rect 422 3162 428 3163
rect 422 3158 423 3162
rect 427 3158 428 3162
rect 422 3157 428 3158
rect 566 3162 572 3163
rect 566 3158 567 3162
rect 571 3158 572 3162
rect 566 3157 572 3158
rect 726 3162 732 3163
rect 726 3158 727 3162
rect 731 3158 732 3162
rect 726 3157 732 3158
rect 902 3162 908 3163
rect 902 3158 903 3162
rect 907 3158 908 3162
rect 902 3157 908 3158
rect 1094 3162 1100 3163
rect 1094 3158 1095 3162
rect 1099 3158 1100 3162
rect 1094 3157 1100 3158
rect 1294 3162 1300 3163
rect 1294 3158 1295 3162
rect 1299 3158 1300 3162
rect 1294 3157 1300 3158
rect 1494 3162 1500 3163
rect 1494 3158 1495 3162
rect 1499 3158 1500 3162
rect 1494 3157 1500 3158
rect 1702 3162 1708 3163
rect 1702 3158 1703 3162
rect 1707 3158 1708 3162
rect 1702 3157 1708 3158
rect 1918 3162 1924 3163
rect 1918 3158 1919 3162
rect 1923 3158 1924 3162
rect 2032 3158 2034 3173
rect 1918 3157 1924 3158
rect 2030 3157 2036 3158
rect 110 3153 111 3157
rect 115 3153 116 3157
rect 110 3152 116 3153
rect 2030 3153 2031 3157
rect 2035 3153 2036 3157
rect 2030 3152 2036 3153
rect 2072 3147 2074 3191
rect 2110 3177 2116 3178
rect 2110 3173 2111 3177
rect 2115 3173 2116 3177
rect 2110 3172 2116 3173
rect 2238 3177 2244 3178
rect 2238 3173 2239 3177
rect 2243 3173 2244 3177
rect 2238 3172 2244 3173
rect 2398 3177 2404 3178
rect 2398 3173 2399 3177
rect 2403 3173 2404 3177
rect 2398 3172 2404 3173
rect 2558 3177 2564 3178
rect 2558 3173 2559 3177
rect 2563 3173 2564 3177
rect 2558 3172 2564 3173
rect 2718 3177 2724 3178
rect 2718 3173 2719 3177
rect 2723 3173 2724 3177
rect 2718 3172 2724 3173
rect 2878 3177 2884 3178
rect 2878 3173 2879 3177
rect 2883 3173 2884 3177
rect 2878 3172 2884 3173
rect 3030 3177 3036 3178
rect 3030 3173 3031 3177
rect 3035 3173 3036 3177
rect 3030 3172 3036 3173
rect 3166 3177 3172 3178
rect 3166 3173 3167 3177
rect 3171 3173 3172 3177
rect 3166 3172 3172 3173
rect 3302 3177 3308 3178
rect 3302 3173 3303 3177
rect 3307 3173 3308 3177
rect 3302 3172 3308 3173
rect 3430 3177 3436 3178
rect 3430 3173 3431 3177
rect 3435 3173 3436 3177
rect 3430 3172 3436 3173
rect 3550 3177 3556 3178
rect 3550 3173 3551 3177
rect 3555 3173 3556 3177
rect 3550 3172 3556 3173
rect 3670 3177 3676 3178
rect 3670 3173 3671 3177
rect 3675 3173 3676 3177
rect 3670 3172 3676 3173
rect 3790 3177 3796 3178
rect 3790 3173 3791 3177
rect 3795 3173 3796 3177
rect 3790 3172 3796 3173
rect 3894 3177 3900 3178
rect 3894 3173 3895 3177
rect 3899 3173 3900 3177
rect 3894 3172 3900 3173
rect 2112 3147 2114 3172
rect 2240 3147 2242 3172
rect 2400 3147 2402 3172
rect 2560 3147 2562 3172
rect 2720 3147 2722 3172
rect 2880 3147 2882 3172
rect 3032 3147 3034 3172
rect 3168 3147 3170 3172
rect 3304 3147 3306 3172
rect 3432 3147 3434 3172
rect 3552 3147 3554 3172
rect 3672 3147 3674 3172
rect 3792 3147 3794 3172
rect 3896 3147 3898 3172
rect 3992 3147 3994 3191
rect 2071 3146 2075 3147
rect 2071 3141 2075 3142
rect 2111 3146 2115 3147
rect 2111 3141 2115 3142
rect 2183 3146 2187 3147
rect 2183 3141 2187 3142
rect 2239 3146 2243 3147
rect 2239 3141 2243 3142
rect 2367 3146 2371 3147
rect 2367 3141 2371 3142
rect 2399 3146 2403 3147
rect 2399 3141 2403 3142
rect 2551 3146 2555 3147
rect 2551 3141 2555 3142
rect 2559 3146 2563 3147
rect 2559 3141 2563 3142
rect 2719 3146 2723 3147
rect 2719 3141 2723 3142
rect 2735 3146 2739 3147
rect 2735 3141 2739 3142
rect 2879 3146 2883 3147
rect 2879 3141 2883 3142
rect 2911 3146 2915 3147
rect 2911 3141 2915 3142
rect 3031 3146 3035 3147
rect 3031 3141 3035 3142
rect 3087 3146 3091 3147
rect 3087 3141 3091 3142
rect 3167 3146 3171 3147
rect 3167 3141 3171 3142
rect 3263 3146 3267 3147
rect 3263 3141 3267 3142
rect 3303 3146 3307 3147
rect 3303 3141 3307 3142
rect 3431 3146 3435 3147
rect 3431 3141 3435 3142
rect 3447 3146 3451 3147
rect 3447 3141 3451 3142
rect 3551 3146 3555 3147
rect 3551 3141 3555 3142
rect 3671 3146 3675 3147
rect 3671 3141 3675 3142
rect 3791 3146 3795 3147
rect 3791 3141 3795 3142
rect 3895 3146 3899 3147
rect 3895 3141 3899 3142
rect 3991 3146 3995 3147
rect 3991 3141 3995 3142
rect 110 3140 116 3141
rect 110 3136 111 3140
rect 115 3136 116 3140
rect 110 3135 116 3136
rect 2030 3140 2036 3141
rect 2030 3136 2031 3140
rect 2035 3136 2036 3140
rect 2030 3135 2036 3136
rect 112 3091 114 3135
rect 286 3121 292 3122
rect 286 3117 287 3121
rect 291 3117 292 3121
rect 286 3116 292 3117
rect 422 3121 428 3122
rect 422 3117 423 3121
rect 427 3117 428 3121
rect 422 3116 428 3117
rect 566 3121 572 3122
rect 566 3117 567 3121
rect 571 3117 572 3121
rect 566 3116 572 3117
rect 726 3121 732 3122
rect 726 3117 727 3121
rect 731 3117 732 3121
rect 726 3116 732 3117
rect 902 3121 908 3122
rect 902 3117 903 3121
rect 907 3117 908 3121
rect 902 3116 908 3117
rect 1094 3121 1100 3122
rect 1094 3117 1095 3121
rect 1099 3117 1100 3121
rect 1094 3116 1100 3117
rect 1294 3121 1300 3122
rect 1294 3117 1295 3121
rect 1299 3117 1300 3121
rect 1294 3116 1300 3117
rect 1494 3121 1500 3122
rect 1494 3117 1495 3121
rect 1499 3117 1500 3121
rect 1494 3116 1500 3117
rect 1702 3121 1708 3122
rect 1702 3117 1703 3121
rect 1707 3117 1708 3121
rect 1702 3116 1708 3117
rect 1918 3121 1924 3122
rect 1918 3117 1919 3121
rect 1923 3117 1924 3121
rect 1918 3116 1924 3117
rect 288 3091 290 3116
rect 424 3091 426 3116
rect 568 3091 570 3116
rect 728 3091 730 3116
rect 904 3091 906 3116
rect 1096 3091 1098 3116
rect 1296 3091 1298 3116
rect 1496 3091 1498 3116
rect 1704 3091 1706 3116
rect 1920 3091 1922 3116
rect 2032 3091 2034 3135
rect 2072 3113 2074 3141
rect 2184 3132 2186 3141
rect 2368 3132 2370 3141
rect 2552 3132 2554 3141
rect 2736 3132 2738 3141
rect 2912 3132 2914 3141
rect 3088 3132 3090 3141
rect 3264 3132 3266 3141
rect 3448 3132 3450 3141
rect 2182 3131 2188 3132
rect 2182 3127 2183 3131
rect 2187 3127 2188 3131
rect 2182 3126 2188 3127
rect 2366 3131 2372 3132
rect 2366 3127 2367 3131
rect 2371 3127 2372 3131
rect 2366 3126 2372 3127
rect 2550 3131 2556 3132
rect 2550 3127 2551 3131
rect 2555 3127 2556 3131
rect 2550 3126 2556 3127
rect 2734 3131 2740 3132
rect 2734 3127 2735 3131
rect 2739 3127 2740 3131
rect 2734 3126 2740 3127
rect 2910 3131 2916 3132
rect 2910 3127 2911 3131
rect 2915 3127 2916 3131
rect 2910 3126 2916 3127
rect 3086 3131 3092 3132
rect 3086 3127 3087 3131
rect 3091 3127 3092 3131
rect 3086 3126 3092 3127
rect 3262 3131 3268 3132
rect 3262 3127 3263 3131
rect 3267 3127 3268 3131
rect 3262 3126 3268 3127
rect 3446 3131 3452 3132
rect 3446 3127 3447 3131
rect 3451 3127 3452 3131
rect 3446 3126 3452 3127
rect 3992 3113 3994 3141
rect 2070 3112 2076 3113
rect 2070 3108 2071 3112
rect 2075 3108 2076 3112
rect 2070 3107 2076 3108
rect 3990 3112 3996 3113
rect 3990 3108 3991 3112
rect 3995 3108 3996 3112
rect 3990 3107 3996 3108
rect 2070 3095 2076 3096
rect 2070 3091 2071 3095
rect 2075 3091 2076 3095
rect 3990 3095 3996 3096
rect 3990 3091 3991 3095
rect 3995 3091 3996 3095
rect 111 3090 115 3091
rect 111 3085 115 3086
rect 287 3090 291 3091
rect 287 3085 291 3086
rect 423 3090 427 3091
rect 423 3085 427 3086
rect 567 3090 571 3091
rect 567 3085 571 3086
rect 575 3090 579 3091
rect 575 3085 579 3086
rect 679 3090 683 3091
rect 679 3085 683 3086
rect 727 3090 731 3091
rect 727 3085 731 3086
rect 799 3090 803 3091
rect 799 3085 803 3086
rect 903 3090 907 3091
rect 903 3085 907 3086
rect 935 3090 939 3091
rect 935 3085 939 3086
rect 1079 3090 1083 3091
rect 1079 3085 1083 3086
rect 1095 3090 1099 3091
rect 1095 3085 1099 3086
rect 1231 3090 1235 3091
rect 1231 3085 1235 3086
rect 1295 3090 1299 3091
rect 1295 3085 1299 3086
rect 1391 3090 1395 3091
rect 1391 3085 1395 3086
rect 1495 3090 1499 3091
rect 1495 3085 1499 3086
rect 1559 3090 1563 3091
rect 1559 3085 1563 3086
rect 1703 3090 1707 3091
rect 1703 3085 1707 3086
rect 1727 3090 1731 3091
rect 1727 3085 1731 3086
rect 1903 3090 1907 3091
rect 1903 3085 1907 3086
rect 1919 3090 1923 3091
rect 1919 3085 1923 3086
rect 2031 3090 2035 3091
rect 2070 3090 2076 3091
rect 2182 3090 2188 3091
rect 2031 3085 2035 3086
rect 112 3057 114 3085
rect 576 3076 578 3085
rect 680 3076 682 3085
rect 800 3076 802 3085
rect 936 3076 938 3085
rect 1080 3076 1082 3085
rect 1232 3076 1234 3085
rect 1392 3076 1394 3085
rect 1560 3076 1562 3085
rect 1728 3076 1730 3085
rect 1904 3076 1906 3085
rect 574 3075 580 3076
rect 574 3071 575 3075
rect 579 3071 580 3075
rect 574 3070 580 3071
rect 678 3075 684 3076
rect 678 3071 679 3075
rect 683 3071 684 3075
rect 678 3070 684 3071
rect 798 3075 804 3076
rect 798 3071 799 3075
rect 803 3071 804 3075
rect 798 3070 804 3071
rect 934 3075 940 3076
rect 934 3071 935 3075
rect 939 3071 940 3075
rect 934 3070 940 3071
rect 1078 3075 1084 3076
rect 1078 3071 1079 3075
rect 1083 3071 1084 3075
rect 1078 3070 1084 3071
rect 1230 3075 1236 3076
rect 1230 3071 1231 3075
rect 1235 3071 1236 3075
rect 1230 3070 1236 3071
rect 1390 3075 1396 3076
rect 1390 3071 1391 3075
rect 1395 3071 1396 3075
rect 1390 3070 1396 3071
rect 1558 3075 1564 3076
rect 1558 3071 1559 3075
rect 1563 3071 1564 3075
rect 1558 3070 1564 3071
rect 1726 3075 1732 3076
rect 1726 3071 1727 3075
rect 1731 3071 1732 3075
rect 1726 3070 1732 3071
rect 1902 3075 1908 3076
rect 1902 3071 1903 3075
rect 1907 3071 1908 3075
rect 1902 3070 1908 3071
rect 2032 3057 2034 3085
rect 2072 3067 2074 3090
rect 2182 3086 2183 3090
rect 2187 3086 2188 3090
rect 2182 3085 2188 3086
rect 2366 3090 2372 3091
rect 2366 3086 2367 3090
rect 2371 3086 2372 3090
rect 2366 3085 2372 3086
rect 2550 3090 2556 3091
rect 2550 3086 2551 3090
rect 2555 3086 2556 3090
rect 2550 3085 2556 3086
rect 2734 3090 2740 3091
rect 2734 3086 2735 3090
rect 2739 3086 2740 3090
rect 2734 3085 2740 3086
rect 2910 3090 2916 3091
rect 2910 3086 2911 3090
rect 2915 3086 2916 3090
rect 2910 3085 2916 3086
rect 3086 3090 3092 3091
rect 3086 3086 3087 3090
rect 3091 3086 3092 3090
rect 3086 3085 3092 3086
rect 3262 3090 3268 3091
rect 3262 3086 3263 3090
rect 3267 3086 3268 3090
rect 3262 3085 3268 3086
rect 3446 3090 3452 3091
rect 3990 3090 3996 3091
rect 3446 3086 3447 3090
rect 3451 3086 3452 3090
rect 3446 3085 3452 3086
rect 2184 3067 2186 3085
rect 2368 3067 2370 3085
rect 2552 3067 2554 3085
rect 2736 3067 2738 3085
rect 2912 3067 2914 3085
rect 3088 3067 3090 3085
rect 3264 3067 3266 3085
rect 3448 3067 3450 3085
rect 3992 3067 3994 3090
rect 2071 3066 2075 3067
rect 2071 3061 2075 3062
rect 2183 3066 2187 3067
rect 2183 3061 2187 3062
rect 2351 3066 2355 3067
rect 2351 3061 2355 3062
rect 2367 3066 2371 3067
rect 2367 3061 2371 3062
rect 2455 3066 2459 3067
rect 2455 3061 2459 3062
rect 2551 3066 2555 3067
rect 2551 3061 2555 3062
rect 2567 3066 2571 3067
rect 2567 3061 2571 3062
rect 2687 3066 2691 3067
rect 2687 3061 2691 3062
rect 2735 3066 2739 3067
rect 2735 3061 2739 3062
rect 2807 3066 2811 3067
rect 2807 3061 2811 3062
rect 2911 3066 2915 3067
rect 2911 3061 2915 3062
rect 2927 3066 2931 3067
rect 2927 3061 2931 3062
rect 3047 3066 3051 3067
rect 3047 3061 3051 3062
rect 3087 3066 3091 3067
rect 3087 3061 3091 3062
rect 3167 3066 3171 3067
rect 3167 3061 3171 3062
rect 3263 3066 3267 3067
rect 3263 3061 3267 3062
rect 3295 3066 3299 3067
rect 3295 3061 3299 3062
rect 3447 3066 3451 3067
rect 3447 3061 3451 3062
rect 3991 3066 3995 3067
rect 3991 3061 3995 3062
rect 110 3056 116 3057
rect 110 3052 111 3056
rect 115 3052 116 3056
rect 110 3051 116 3052
rect 2030 3056 2036 3057
rect 2030 3052 2031 3056
rect 2035 3052 2036 3056
rect 2030 3051 2036 3052
rect 2072 3046 2074 3061
rect 2352 3051 2354 3061
rect 2456 3051 2458 3061
rect 2568 3051 2570 3061
rect 2688 3051 2690 3061
rect 2808 3051 2810 3061
rect 2928 3051 2930 3061
rect 3048 3051 3050 3061
rect 3168 3051 3170 3061
rect 3296 3051 3298 3061
rect 2350 3050 2356 3051
rect 2350 3046 2351 3050
rect 2355 3046 2356 3050
rect 2070 3045 2076 3046
rect 2350 3045 2356 3046
rect 2454 3050 2460 3051
rect 2454 3046 2455 3050
rect 2459 3046 2460 3050
rect 2454 3045 2460 3046
rect 2566 3050 2572 3051
rect 2566 3046 2567 3050
rect 2571 3046 2572 3050
rect 2566 3045 2572 3046
rect 2686 3050 2692 3051
rect 2686 3046 2687 3050
rect 2691 3046 2692 3050
rect 2686 3045 2692 3046
rect 2806 3050 2812 3051
rect 2806 3046 2807 3050
rect 2811 3046 2812 3050
rect 2806 3045 2812 3046
rect 2926 3050 2932 3051
rect 2926 3046 2927 3050
rect 2931 3046 2932 3050
rect 2926 3045 2932 3046
rect 3046 3050 3052 3051
rect 3046 3046 3047 3050
rect 3051 3046 3052 3050
rect 3046 3045 3052 3046
rect 3166 3050 3172 3051
rect 3166 3046 3167 3050
rect 3171 3046 3172 3050
rect 3166 3045 3172 3046
rect 3294 3050 3300 3051
rect 3294 3046 3295 3050
rect 3299 3046 3300 3050
rect 3992 3046 3994 3061
rect 3294 3045 3300 3046
rect 3990 3045 3996 3046
rect 2070 3041 2071 3045
rect 2075 3041 2076 3045
rect 2070 3040 2076 3041
rect 3990 3041 3991 3045
rect 3995 3041 3996 3045
rect 3990 3040 3996 3041
rect 110 3039 116 3040
rect 110 3035 111 3039
rect 115 3035 116 3039
rect 2030 3039 2036 3040
rect 2030 3035 2031 3039
rect 2035 3035 2036 3039
rect 110 3034 116 3035
rect 574 3034 580 3035
rect 112 3007 114 3034
rect 574 3030 575 3034
rect 579 3030 580 3034
rect 574 3029 580 3030
rect 678 3034 684 3035
rect 678 3030 679 3034
rect 683 3030 684 3034
rect 678 3029 684 3030
rect 798 3034 804 3035
rect 798 3030 799 3034
rect 803 3030 804 3034
rect 798 3029 804 3030
rect 934 3034 940 3035
rect 934 3030 935 3034
rect 939 3030 940 3034
rect 934 3029 940 3030
rect 1078 3034 1084 3035
rect 1078 3030 1079 3034
rect 1083 3030 1084 3034
rect 1078 3029 1084 3030
rect 1230 3034 1236 3035
rect 1230 3030 1231 3034
rect 1235 3030 1236 3034
rect 1230 3029 1236 3030
rect 1390 3034 1396 3035
rect 1390 3030 1391 3034
rect 1395 3030 1396 3034
rect 1390 3029 1396 3030
rect 1558 3034 1564 3035
rect 1558 3030 1559 3034
rect 1563 3030 1564 3034
rect 1558 3029 1564 3030
rect 1726 3034 1732 3035
rect 1726 3030 1727 3034
rect 1731 3030 1732 3034
rect 1726 3029 1732 3030
rect 1902 3034 1908 3035
rect 2030 3034 2036 3035
rect 1902 3030 1903 3034
rect 1907 3030 1908 3034
rect 1902 3029 1908 3030
rect 576 3007 578 3029
rect 680 3007 682 3029
rect 800 3007 802 3029
rect 936 3007 938 3029
rect 1080 3007 1082 3029
rect 1232 3007 1234 3029
rect 1392 3007 1394 3029
rect 1560 3007 1562 3029
rect 1728 3007 1730 3029
rect 1904 3007 1906 3029
rect 2032 3007 2034 3034
rect 2070 3028 2076 3029
rect 2070 3024 2071 3028
rect 2075 3024 2076 3028
rect 2070 3023 2076 3024
rect 3990 3028 3996 3029
rect 3990 3024 3991 3028
rect 3995 3024 3996 3028
rect 3990 3023 3996 3024
rect 111 3006 115 3007
rect 111 3001 115 3002
rect 551 3006 555 3007
rect 551 3001 555 3002
rect 575 3006 579 3007
rect 575 3001 579 3002
rect 655 3006 659 3007
rect 655 3001 659 3002
rect 679 3006 683 3007
rect 679 3001 683 3002
rect 759 3006 763 3007
rect 759 3001 763 3002
rect 799 3006 803 3007
rect 799 3001 803 3002
rect 871 3006 875 3007
rect 871 3001 875 3002
rect 935 3006 939 3007
rect 935 3001 939 3002
rect 991 3006 995 3007
rect 991 3001 995 3002
rect 1079 3006 1083 3007
rect 1079 3001 1083 3002
rect 1119 3006 1123 3007
rect 1119 3001 1123 3002
rect 1231 3006 1235 3007
rect 1231 3001 1235 3002
rect 1255 3006 1259 3007
rect 1255 3001 1259 3002
rect 1391 3006 1395 3007
rect 1391 3001 1395 3002
rect 1535 3006 1539 3007
rect 1535 3001 1539 3002
rect 1559 3006 1563 3007
rect 1559 3001 1563 3002
rect 1687 3006 1691 3007
rect 1687 3001 1691 3002
rect 1727 3006 1731 3007
rect 1727 3001 1731 3002
rect 1903 3006 1907 3007
rect 1903 3001 1907 3002
rect 2031 3006 2035 3007
rect 2031 3001 2035 3002
rect 112 2986 114 3001
rect 552 2991 554 3001
rect 656 2991 658 3001
rect 760 2991 762 3001
rect 872 2991 874 3001
rect 992 2991 994 3001
rect 1120 2991 1122 3001
rect 1256 2991 1258 3001
rect 1392 2991 1394 3001
rect 1536 2991 1538 3001
rect 1688 2991 1690 3001
rect 550 2990 556 2991
rect 550 2986 551 2990
rect 555 2986 556 2990
rect 110 2985 116 2986
rect 550 2985 556 2986
rect 654 2990 660 2991
rect 654 2986 655 2990
rect 659 2986 660 2990
rect 654 2985 660 2986
rect 758 2990 764 2991
rect 758 2986 759 2990
rect 763 2986 764 2990
rect 758 2985 764 2986
rect 870 2990 876 2991
rect 870 2986 871 2990
rect 875 2986 876 2990
rect 870 2985 876 2986
rect 990 2990 996 2991
rect 990 2986 991 2990
rect 995 2986 996 2990
rect 990 2985 996 2986
rect 1118 2990 1124 2991
rect 1118 2986 1119 2990
rect 1123 2986 1124 2990
rect 1118 2985 1124 2986
rect 1254 2990 1260 2991
rect 1254 2986 1255 2990
rect 1259 2986 1260 2990
rect 1254 2985 1260 2986
rect 1390 2990 1396 2991
rect 1390 2986 1391 2990
rect 1395 2986 1396 2990
rect 1390 2985 1396 2986
rect 1534 2990 1540 2991
rect 1534 2986 1535 2990
rect 1539 2986 1540 2990
rect 1534 2985 1540 2986
rect 1686 2990 1692 2991
rect 1686 2986 1687 2990
rect 1691 2986 1692 2990
rect 2032 2986 2034 3001
rect 2072 2995 2074 3023
rect 2350 3009 2356 3010
rect 2350 3005 2351 3009
rect 2355 3005 2356 3009
rect 2350 3004 2356 3005
rect 2454 3009 2460 3010
rect 2454 3005 2455 3009
rect 2459 3005 2460 3009
rect 2454 3004 2460 3005
rect 2566 3009 2572 3010
rect 2566 3005 2567 3009
rect 2571 3005 2572 3009
rect 2566 3004 2572 3005
rect 2686 3009 2692 3010
rect 2686 3005 2687 3009
rect 2691 3005 2692 3009
rect 2686 3004 2692 3005
rect 2806 3009 2812 3010
rect 2806 3005 2807 3009
rect 2811 3005 2812 3009
rect 2806 3004 2812 3005
rect 2926 3009 2932 3010
rect 2926 3005 2927 3009
rect 2931 3005 2932 3009
rect 2926 3004 2932 3005
rect 3046 3009 3052 3010
rect 3046 3005 3047 3009
rect 3051 3005 3052 3009
rect 3046 3004 3052 3005
rect 3166 3009 3172 3010
rect 3166 3005 3167 3009
rect 3171 3005 3172 3009
rect 3166 3004 3172 3005
rect 3294 3009 3300 3010
rect 3294 3005 3295 3009
rect 3299 3005 3300 3009
rect 3294 3004 3300 3005
rect 2352 2995 2354 3004
rect 2456 2995 2458 3004
rect 2568 2995 2570 3004
rect 2688 2995 2690 3004
rect 2808 2995 2810 3004
rect 2928 2995 2930 3004
rect 3048 2995 3050 3004
rect 3168 2995 3170 3004
rect 3296 2995 3298 3004
rect 3992 2995 3994 3023
rect 2071 2994 2075 2995
rect 2071 2989 2075 2990
rect 2351 2994 2355 2995
rect 2351 2989 2355 2990
rect 2455 2994 2459 2995
rect 2455 2989 2459 2990
rect 2495 2994 2499 2995
rect 2495 2989 2499 2990
rect 2567 2994 2571 2995
rect 2567 2989 2571 2990
rect 2599 2994 2603 2995
rect 2599 2989 2603 2990
rect 2687 2994 2691 2995
rect 2687 2989 2691 2990
rect 2703 2994 2707 2995
rect 2703 2989 2707 2990
rect 2807 2994 2811 2995
rect 2807 2989 2811 2990
rect 2911 2994 2915 2995
rect 2911 2989 2915 2990
rect 2927 2994 2931 2995
rect 2927 2989 2931 2990
rect 3015 2994 3019 2995
rect 3015 2989 3019 2990
rect 3047 2994 3051 2995
rect 3047 2989 3051 2990
rect 3119 2994 3123 2995
rect 3119 2989 3123 2990
rect 3167 2994 3171 2995
rect 3167 2989 3171 2990
rect 3223 2994 3227 2995
rect 3223 2989 3227 2990
rect 3295 2994 3299 2995
rect 3295 2989 3299 2990
rect 3991 2994 3995 2995
rect 3991 2989 3995 2990
rect 1686 2985 1692 2986
rect 2030 2985 2036 2986
rect 110 2981 111 2985
rect 115 2981 116 2985
rect 110 2980 116 2981
rect 2030 2981 2031 2985
rect 2035 2981 2036 2985
rect 2030 2980 2036 2981
rect 110 2968 116 2969
rect 110 2964 111 2968
rect 115 2964 116 2968
rect 110 2963 116 2964
rect 2030 2968 2036 2969
rect 2030 2964 2031 2968
rect 2035 2964 2036 2968
rect 2030 2963 2036 2964
rect 112 2923 114 2963
rect 550 2949 556 2950
rect 550 2945 551 2949
rect 555 2945 556 2949
rect 550 2944 556 2945
rect 654 2949 660 2950
rect 654 2945 655 2949
rect 659 2945 660 2949
rect 654 2944 660 2945
rect 758 2949 764 2950
rect 758 2945 759 2949
rect 763 2945 764 2949
rect 758 2944 764 2945
rect 870 2949 876 2950
rect 870 2945 871 2949
rect 875 2945 876 2949
rect 870 2944 876 2945
rect 990 2949 996 2950
rect 990 2945 991 2949
rect 995 2945 996 2949
rect 990 2944 996 2945
rect 1118 2949 1124 2950
rect 1118 2945 1119 2949
rect 1123 2945 1124 2949
rect 1118 2944 1124 2945
rect 1254 2949 1260 2950
rect 1254 2945 1255 2949
rect 1259 2945 1260 2949
rect 1254 2944 1260 2945
rect 1390 2949 1396 2950
rect 1390 2945 1391 2949
rect 1395 2945 1396 2949
rect 1390 2944 1396 2945
rect 1534 2949 1540 2950
rect 1534 2945 1535 2949
rect 1539 2945 1540 2949
rect 1534 2944 1540 2945
rect 1686 2949 1692 2950
rect 1686 2945 1687 2949
rect 1691 2945 1692 2949
rect 1686 2944 1692 2945
rect 552 2923 554 2944
rect 656 2923 658 2944
rect 760 2923 762 2944
rect 872 2923 874 2944
rect 992 2923 994 2944
rect 1120 2923 1122 2944
rect 1256 2923 1258 2944
rect 1392 2923 1394 2944
rect 1536 2923 1538 2944
rect 1688 2923 1690 2944
rect 2032 2923 2034 2963
rect 2072 2961 2074 2989
rect 2496 2980 2498 2989
rect 2600 2980 2602 2989
rect 2704 2980 2706 2989
rect 2808 2980 2810 2989
rect 2912 2980 2914 2989
rect 3016 2980 3018 2989
rect 3120 2980 3122 2989
rect 3224 2980 3226 2989
rect 2494 2979 2500 2980
rect 2494 2975 2495 2979
rect 2499 2975 2500 2979
rect 2494 2974 2500 2975
rect 2598 2979 2604 2980
rect 2598 2975 2599 2979
rect 2603 2975 2604 2979
rect 2598 2974 2604 2975
rect 2702 2979 2708 2980
rect 2702 2975 2703 2979
rect 2707 2975 2708 2979
rect 2702 2974 2708 2975
rect 2806 2979 2812 2980
rect 2806 2975 2807 2979
rect 2811 2975 2812 2979
rect 2806 2974 2812 2975
rect 2910 2979 2916 2980
rect 2910 2975 2911 2979
rect 2915 2975 2916 2979
rect 2910 2974 2916 2975
rect 3014 2979 3020 2980
rect 3014 2975 3015 2979
rect 3019 2975 3020 2979
rect 3014 2974 3020 2975
rect 3118 2979 3124 2980
rect 3118 2975 3119 2979
rect 3123 2975 3124 2979
rect 3118 2974 3124 2975
rect 3222 2979 3228 2980
rect 3222 2975 3223 2979
rect 3227 2975 3228 2979
rect 3222 2974 3228 2975
rect 3992 2961 3994 2989
rect 2070 2960 2076 2961
rect 2070 2956 2071 2960
rect 2075 2956 2076 2960
rect 2070 2955 2076 2956
rect 3990 2960 3996 2961
rect 3990 2956 3991 2960
rect 3995 2956 3996 2960
rect 3990 2955 3996 2956
rect 2070 2943 2076 2944
rect 2070 2939 2071 2943
rect 2075 2939 2076 2943
rect 3990 2943 3996 2944
rect 3990 2939 3991 2943
rect 3995 2939 3996 2943
rect 2070 2938 2076 2939
rect 2494 2938 2500 2939
rect 2072 2923 2074 2938
rect 2494 2934 2495 2938
rect 2499 2934 2500 2938
rect 2494 2933 2500 2934
rect 2598 2938 2604 2939
rect 2598 2934 2599 2938
rect 2603 2934 2604 2938
rect 2598 2933 2604 2934
rect 2702 2938 2708 2939
rect 2702 2934 2703 2938
rect 2707 2934 2708 2938
rect 2702 2933 2708 2934
rect 2806 2938 2812 2939
rect 2806 2934 2807 2938
rect 2811 2934 2812 2938
rect 2806 2933 2812 2934
rect 2910 2938 2916 2939
rect 2910 2934 2911 2938
rect 2915 2934 2916 2938
rect 2910 2933 2916 2934
rect 3014 2938 3020 2939
rect 3014 2934 3015 2938
rect 3019 2934 3020 2938
rect 3014 2933 3020 2934
rect 3118 2938 3124 2939
rect 3118 2934 3119 2938
rect 3123 2934 3124 2938
rect 3118 2933 3124 2934
rect 3222 2938 3228 2939
rect 3990 2938 3996 2939
rect 3222 2934 3223 2938
rect 3227 2934 3228 2938
rect 3222 2933 3228 2934
rect 2496 2923 2498 2933
rect 2600 2923 2602 2933
rect 2704 2923 2706 2933
rect 2808 2923 2810 2933
rect 2912 2923 2914 2933
rect 3016 2923 3018 2933
rect 3120 2923 3122 2933
rect 3224 2923 3226 2933
rect 3992 2923 3994 2938
rect 111 2922 115 2923
rect 111 2917 115 2918
rect 311 2922 315 2923
rect 311 2917 315 2918
rect 431 2922 435 2923
rect 431 2917 435 2918
rect 551 2922 555 2923
rect 551 2917 555 2918
rect 559 2922 563 2923
rect 559 2917 563 2918
rect 655 2922 659 2923
rect 655 2917 659 2918
rect 695 2922 699 2923
rect 695 2917 699 2918
rect 759 2922 763 2923
rect 759 2917 763 2918
rect 831 2922 835 2923
rect 831 2917 835 2918
rect 871 2922 875 2923
rect 871 2917 875 2918
rect 975 2922 979 2923
rect 975 2917 979 2918
rect 991 2922 995 2923
rect 991 2917 995 2918
rect 1119 2922 1123 2923
rect 1119 2917 1123 2918
rect 1255 2922 1259 2923
rect 1255 2917 1259 2918
rect 1271 2922 1275 2923
rect 1271 2917 1275 2918
rect 1391 2922 1395 2923
rect 1391 2917 1395 2918
rect 1423 2922 1427 2923
rect 1423 2917 1427 2918
rect 1535 2922 1539 2923
rect 1535 2917 1539 2918
rect 1575 2922 1579 2923
rect 1575 2917 1579 2918
rect 1687 2922 1691 2923
rect 1687 2917 1691 2918
rect 2031 2922 2035 2923
rect 2031 2917 2035 2918
rect 2071 2922 2075 2923
rect 2071 2917 2075 2918
rect 2415 2922 2419 2923
rect 2415 2917 2419 2918
rect 2495 2922 2499 2923
rect 2495 2917 2499 2918
rect 2519 2922 2523 2923
rect 2519 2917 2523 2918
rect 2599 2922 2603 2923
rect 2599 2917 2603 2918
rect 2623 2922 2627 2923
rect 2623 2917 2627 2918
rect 2703 2922 2707 2923
rect 2703 2917 2707 2918
rect 2727 2922 2731 2923
rect 2727 2917 2731 2918
rect 2807 2922 2811 2923
rect 2807 2917 2811 2918
rect 2831 2922 2835 2923
rect 2831 2917 2835 2918
rect 2911 2922 2915 2923
rect 2911 2917 2915 2918
rect 2935 2922 2939 2923
rect 2935 2917 2939 2918
rect 3015 2922 3019 2923
rect 3015 2917 3019 2918
rect 3039 2922 3043 2923
rect 3039 2917 3043 2918
rect 3119 2922 3123 2923
rect 3119 2917 3123 2918
rect 3143 2922 3147 2923
rect 3143 2917 3147 2918
rect 3223 2922 3227 2923
rect 3223 2917 3227 2918
rect 3247 2922 3251 2923
rect 3247 2917 3251 2918
rect 3991 2922 3995 2923
rect 3991 2917 3995 2918
rect 112 2889 114 2917
rect 312 2908 314 2917
rect 432 2908 434 2917
rect 560 2908 562 2917
rect 696 2908 698 2917
rect 832 2908 834 2917
rect 976 2908 978 2917
rect 1120 2908 1122 2917
rect 1272 2908 1274 2917
rect 1424 2908 1426 2917
rect 1576 2908 1578 2917
rect 310 2907 316 2908
rect 310 2903 311 2907
rect 315 2903 316 2907
rect 310 2902 316 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 558 2907 564 2908
rect 558 2903 559 2907
rect 563 2903 564 2907
rect 558 2902 564 2903
rect 694 2907 700 2908
rect 694 2903 695 2907
rect 699 2903 700 2907
rect 694 2902 700 2903
rect 830 2907 836 2908
rect 830 2903 831 2907
rect 835 2903 836 2907
rect 830 2902 836 2903
rect 974 2907 980 2908
rect 974 2903 975 2907
rect 979 2903 980 2907
rect 974 2902 980 2903
rect 1118 2907 1124 2908
rect 1118 2903 1119 2907
rect 1123 2903 1124 2907
rect 1118 2902 1124 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1422 2907 1428 2908
rect 1422 2903 1423 2907
rect 1427 2903 1428 2907
rect 1422 2902 1428 2903
rect 1574 2907 1580 2908
rect 1574 2903 1575 2907
rect 1579 2903 1580 2907
rect 1574 2902 1580 2903
rect 2032 2889 2034 2917
rect 2072 2902 2074 2917
rect 2416 2907 2418 2917
rect 2520 2907 2522 2917
rect 2624 2907 2626 2917
rect 2728 2907 2730 2917
rect 2832 2907 2834 2917
rect 2936 2907 2938 2917
rect 3040 2907 3042 2917
rect 3144 2907 3146 2917
rect 3248 2907 3250 2917
rect 2414 2906 2420 2907
rect 2414 2902 2415 2906
rect 2419 2902 2420 2906
rect 2070 2901 2076 2902
rect 2414 2901 2420 2902
rect 2518 2906 2524 2907
rect 2518 2902 2519 2906
rect 2523 2902 2524 2906
rect 2518 2901 2524 2902
rect 2622 2906 2628 2907
rect 2622 2902 2623 2906
rect 2627 2902 2628 2906
rect 2622 2901 2628 2902
rect 2726 2906 2732 2907
rect 2726 2902 2727 2906
rect 2731 2902 2732 2906
rect 2726 2901 2732 2902
rect 2830 2906 2836 2907
rect 2830 2902 2831 2906
rect 2835 2902 2836 2906
rect 2830 2901 2836 2902
rect 2934 2906 2940 2907
rect 2934 2902 2935 2906
rect 2939 2902 2940 2906
rect 2934 2901 2940 2902
rect 3038 2906 3044 2907
rect 3038 2902 3039 2906
rect 3043 2902 3044 2906
rect 3038 2901 3044 2902
rect 3142 2906 3148 2907
rect 3142 2902 3143 2906
rect 3147 2902 3148 2906
rect 3142 2901 3148 2902
rect 3246 2906 3252 2907
rect 3246 2902 3247 2906
rect 3251 2902 3252 2906
rect 3992 2902 3994 2917
rect 3246 2901 3252 2902
rect 3990 2901 3996 2902
rect 2070 2897 2071 2901
rect 2075 2897 2076 2901
rect 2070 2896 2076 2897
rect 3990 2897 3991 2901
rect 3995 2897 3996 2901
rect 3990 2896 3996 2897
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 110 2883 116 2884
rect 2030 2888 2036 2889
rect 2030 2884 2031 2888
rect 2035 2884 2036 2888
rect 2030 2883 2036 2884
rect 2070 2884 2076 2885
rect 2070 2880 2071 2884
rect 2075 2880 2076 2884
rect 2070 2879 2076 2880
rect 3990 2884 3996 2885
rect 3990 2880 3991 2884
rect 3995 2880 3996 2884
rect 3990 2879 3996 2880
rect 110 2871 116 2872
rect 110 2867 111 2871
rect 115 2867 116 2871
rect 2030 2871 2036 2872
rect 2030 2867 2031 2871
rect 2035 2867 2036 2871
rect 110 2866 116 2867
rect 310 2866 316 2867
rect 112 2835 114 2866
rect 310 2862 311 2866
rect 315 2862 316 2866
rect 310 2861 316 2862
rect 430 2866 436 2867
rect 430 2862 431 2866
rect 435 2862 436 2866
rect 430 2861 436 2862
rect 558 2866 564 2867
rect 558 2862 559 2866
rect 563 2862 564 2866
rect 558 2861 564 2862
rect 694 2866 700 2867
rect 694 2862 695 2866
rect 699 2862 700 2866
rect 694 2861 700 2862
rect 830 2866 836 2867
rect 830 2862 831 2866
rect 835 2862 836 2866
rect 830 2861 836 2862
rect 974 2866 980 2867
rect 974 2862 975 2866
rect 979 2862 980 2866
rect 974 2861 980 2862
rect 1118 2866 1124 2867
rect 1118 2862 1119 2866
rect 1123 2862 1124 2866
rect 1118 2861 1124 2862
rect 1270 2866 1276 2867
rect 1270 2862 1271 2866
rect 1275 2862 1276 2866
rect 1270 2861 1276 2862
rect 1422 2866 1428 2867
rect 1422 2862 1423 2866
rect 1427 2862 1428 2866
rect 1422 2861 1428 2862
rect 1574 2866 1580 2867
rect 2030 2866 2036 2867
rect 1574 2862 1575 2866
rect 1579 2862 1580 2866
rect 1574 2861 1580 2862
rect 312 2835 314 2861
rect 432 2835 434 2861
rect 560 2835 562 2861
rect 696 2835 698 2861
rect 832 2835 834 2861
rect 976 2835 978 2861
rect 1120 2835 1122 2861
rect 1272 2835 1274 2861
rect 1424 2835 1426 2861
rect 1576 2835 1578 2861
rect 2032 2835 2034 2866
rect 2072 2847 2074 2879
rect 2414 2865 2420 2866
rect 2414 2861 2415 2865
rect 2419 2861 2420 2865
rect 2414 2860 2420 2861
rect 2518 2865 2524 2866
rect 2518 2861 2519 2865
rect 2523 2861 2524 2865
rect 2518 2860 2524 2861
rect 2622 2865 2628 2866
rect 2622 2861 2623 2865
rect 2627 2861 2628 2865
rect 2622 2860 2628 2861
rect 2726 2865 2732 2866
rect 2726 2861 2727 2865
rect 2731 2861 2732 2865
rect 2726 2860 2732 2861
rect 2830 2865 2836 2866
rect 2830 2861 2831 2865
rect 2835 2861 2836 2865
rect 2830 2860 2836 2861
rect 2934 2865 2940 2866
rect 2934 2861 2935 2865
rect 2939 2861 2940 2865
rect 2934 2860 2940 2861
rect 3038 2865 3044 2866
rect 3038 2861 3039 2865
rect 3043 2861 3044 2865
rect 3038 2860 3044 2861
rect 3142 2865 3148 2866
rect 3142 2861 3143 2865
rect 3147 2861 3148 2865
rect 3142 2860 3148 2861
rect 3246 2865 3252 2866
rect 3246 2861 3247 2865
rect 3251 2861 3252 2865
rect 3246 2860 3252 2861
rect 2416 2847 2418 2860
rect 2520 2847 2522 2860
rect 2624 2847 2626 2860
rect 2728 2847 2730 2860
rect 2832 2847 2834 2860
rect 2936 2847 2938 2860
rect 3040 2847 3042 2860
rect 3144 2847 3146 2860
rect 3248 2847 3250 2860
rect 3992 2847 3994 2879
rect 2071 2846 2075 2847
rect 2071 2841 2075 2842
rect 2407 2846 2411 2847
rect 2407 2841 2411 2842
rect 2415 2846 2419 2847
rect 2415 2841 2419 2842
rect 2511 2846 2515 2847
rect 2511 2841 2515 2842
rect 2519 2846 2523 2847
rect 2519 2841 2523 2842
rect 2615 2846 2619 2847
rect 2615 2841 2619 2842
rect 2623 2846 2627 2847
rect 2623 2841 2627 2842
rect 2719 2846 2723 2847
rect 2719 2841 2723 2842
rect 2727 2846 2731 2847
rect 2727 2841 2731 2842
rect 2823 2846 2827 2847
rect 2823 2841 2827 2842
rect 2831 2846 2835 2847
rect 2831 2841 2835 2842
rect 2927 2846 2931 2847
rect 2927 2841 2931 2842
rect 2935 2846 2939 2847
rect 2935 2841 2939 2842
rect 3031 2846 3035 2847
rect 3031 2841 3035 2842
rect 3039 2846 3043 2847
rect 3039 2841 3043 2842
rect 3135 2846 3139 2847
rect 3135 2841 3139 2842
rect 3143 2846 3147 2847
rect 3143 2841 3147 2842
rect 3239 2846 3243 2847
rect 3239 2841 3243 2842
rect 3247 2846 3251 2847
rect 3247 2841 3251 2842
rect 3991 2846 3995 2847
rect 3991 2841 3995 2842
rect 111 2834 115 2835
rect 111 2829 115 2830
rect 151 2834 155 2835
rect 151 2829 155 2830
rect 311 2834 315 2835
rect 311 2829 315 2830
rect 431 2834 435 2835
rect 431 2829 435 2830
rect 471 2834 475 2835
rect 471 2829 475 2830
rect 559 2834 563 2835
rect 559 2829 563 2830
rect 623 2834 627 2835
rect 623 2829 627 2830
rect 695 2834 699 2835
rect 695 2829 699 2830
rect 767 2834 771 2835
rect 767 2829 771 2830
rect 831 2834 835 2835
rect 831 2829 835 2830
rect 903 2834 907 2835
rect 903 2829 907 2830
rect 975 2834 979 2835
rect 975 2829 979 2830
rect 1031 2834 1035 2835
rect 1031 2829 1035 2830
rect 1119 2834 1123 2835
rect 1119 2829 1123 2830
rect 1159 2834 1163 2835
rect 1159 2829 1163 2830
rect 1271 2834 1275 2835
rect 1271 2829 1275 2830
rect 1287 2834 1291 2835
rect 1287 2829 1291 2830
rect 1415 2834 1419 2835
rect 1415 2829 1419 2830
rect 1423 2834 1427 2835
rect 1423 2829 1427 2830
rect 1575 2834 1579 2835
rect 1575 2829 1579 2830
rect 2031 2834 2035 2835
rect 2031 2829 2035 2830
rect 112 2814 114 2829
rect 152 2819 154 2829
rect 312 2819 314 2829
rect 472 2819 474 2829
rect 624 2819 626 2829
rect 768 2819 770 2829
rect 904 2819 906 2829
rect 1032 2819 1034 2829
rect 1160 2819 1162 2829
rect 1288 2819 1290 2829
rect 1416 2819 1418 2829
rect 150 2818 156 2819
rect 150 2814 151 2818
rect 155 2814 156 2818
rect 110 2813 116 2814
rect 150 2813 156 2814
rect 310 2818 316 2819
rect 310 2814 311 2818
rect 315 2814 316 2818
rect 310 2813 316 2814
rect 470 2818 476 2819
rect 470 2814 471 2818
rect 475 2814 476 2818
rect 470 2813 476 2814
rect 622 2818 628 2819
rect 622 2814 623 2818
rect 627 2814 628 2818
rect 622 2813 628 2814
rect 766 2818 772 2819
rect 766 2814 767 2818
rect 771 2814 772 2818
rect 766 2813 772 2814
rect 902 2818 908 2819
rect 902 2814 903 2818
rect 907 2814 908 2818
rect 902 2813 908 2814
rect 1030 2818 1036 2819
rect 1030 2814 1031 2818
rect 1035 2814 1036 2818
rect 1030 2813 1036 2814
rect 1158 2818 1164 2819
rect 1158 2814 1159 2818
rect 1163 2814 1164 2818
rect 1158 2813 1164 2814
rect 1286 2818 1292 2819
rect 1286 2814 1287 2818
rect 1291 2814 1292 2818
rect 1286 2813 1292 2814
rect 1414 2818 1420 2819
rect 1414 2814 1415 2818
rect 1419 2814 1420 2818
rect 2032 2814 2034 2829
rect 1414 2813 1420 2814
rect 2030 2813 2036 2814
rect 2072 2813 2074 2841
rect 2408 2832 2410 2841
rect 2512 2832 2514 2841
rect 2616 2832 2618 2841
rect 2720 2832 2722 2841
rect 2824 2832 2826 2841
rect 2928 2832 2930 2841
rect 3032 2832 3034 2841
rect 3136 2832 3138 2841
rect 3240 2832 3242 2841
rect 2406 2831 2412 2832
rect 2406 2827 2407 2831
rect 2411 2827 2412 2831
rect 2406 2826 2412 2827
rect 2510 2831 2516 2832
rect 2510 2827 2511 2831
rect 2515 2827 2516 2831
rect 2510 2826 2516 2827
rect 2614 2831 2620 2832
rect 2614 2827 2615 2831
rect 2619 2827 2620 2831
rect 2614 2826 2620 2827
rect 2718 2831 2724 2832
rect 2718 2827 2719 2831
rect 2723 2827 2724 2831
rect 2718 2826 2724 2827
rect 2822 2831 2828 2832
rect 2822 2827 2823 2831
rect 2827 2827 2828 2831
rect 2822 2826 2828 2827
rect 2926 2831 2932 2832
rect 2926 2827 2927 2831
rect 2931 2827 2932 2831
rect 2926 2826 2932 2827
rect 3030 2831 3036 2832
rect 3030 2827 3031 2831
rect 3035 2827 3036 2831
rect 3030 2826 3036 2827
rect 3134 2831 3140 2832
rect 3134 2827 3135 2831
rect 3139 2827 3140 2831
rect 3134 2826 3140 2827
rect 3238 2831 3244 2832
rect 3238 2827 3239 2831
rect 3243 2827 3244 2831
rect 3238 2826 3244 2827
rect 3992 2813 3994 2841
rect 110 2809 111 2813
rect 115 2809 116 2813
rect 110 2808 116 2809
rect 2030 2809 2031 2813
rect 2035 2809 2036 2813
rect 2030 2808 2036 2809
rect 2070 2812 2076 2813
rect 2070 2808 2071 2812
rect 2075 2808 2076 2812
rect 2070 2807 2076 2808
rect 3990 2812 3996 2813
rect 3990 2808 3991 2812
rect 3995 2808 3996 2812
rect 3990 2807 3996 2808
rect 110 2796 116 2797
rect 110 2792 111 2796
rect 115 2792 116 2796
rect 110 2791 116 2792
rect 2030 2796 2036 2797
rect 2030 2792 2031 2796
rect 2035 2792 2036 2796
rect 2030 2791 2036 2792
rect 2070 2795 2076 2796
rect 2070 2791 2071 2795
rect 2075 2791 2076 2795
rect 3990 2795 3996 2796
rect 3990 2791 3991 2795
rect 3995 2791 3996 2795
rect 112 2747 114 2791
rect 150 2777 156 2778
rect 150 2773 151 2777
rect 155 2773 156 2777
rect 150 2772 156 2773
rect 310 2777 316 2778
rect 310 2773 311 2777
rect 315 2773 316 2777
rect 310 2772 316 2773
rect 470 2777 476 2778
rect 470 2773 471 2777
rect 475 2773 476 2777
rect 470 2772 476 2773
rect 622 2777 628 2778
rect 622 2773 623 2777
rect 627 2773 628 2777
rect 622 2772 628 2773
rect 766 2777 772 2778
rect 766 2773 767 2777
rect 771 2773 772 2777
rect 766 2772 772 2773
rect 902 2777 908 2778
rect 902 2773 903 2777
rect 907 2773 908 2777
rect 902 2772 908 2773
rect 1030 2777 1036 2778
rect 1030 2773 1031 2777
rect 1035 2773 1036 2777
rect 1030 2772 1036 2773
rect 1158 2777 1164 2778
rect 1158 2773 1159 2777
rect 1163 2773 1164 2777
rect 1158 2772 1164 2773
rect 1286 2777 1292 2778
rect 1286 2773 1287 2777
rect 1291 2773 1292 2777
rect 1286 2772 1292 2773
rect 1414 2777 1420 2778
rect 1414 2773 1415 2777
rect 1419 2773 1420 2777
rect 1414 2772 1420 2773
rect 152 2747 154 2772
rect 312 2747 314 2772
rect 472 2747 474 2772
rect 624 2747 626 2772
rect 768 2747 770 2772
rect 904 2747 906 2772
rect 1032 2747 1034 2772
rect 1160 2747 1162 2772
rect 1288 2747 1290 2772
rect 1416 2747 1418 2772
rect 2032 2747 2034 2791
rect 2070 2790 2076 2791
rect 2406 2790 2412 2791
rect 2072 2767 2074 2790
rect 2406 2786 2407 2790
rect 2411 2786 2412 2790
rect 2406 2785 2412 2786
rect 2510 2790 2516 2791
rect 2510 2786 2511 2790
rect 2515 2786 2516 2790
rect 2510 2785 2516 2786
rect 2614 2790 2620 2791
rect 2614 2786 2615 2790
rect 2619 2786 2620 2790
rect 2614 2785 2620 2786
rect 2718 2790 2724 2791
rect 2718 2786 2719 2790
rect 2723 2786 2724 2790
rect 2718 2785 2724 2786
rect 2822 2790 2828 2791
rect 2822 2786 2823 2790
rect 2827 2786 2828 2790
rect 2822 2785 2828 2786
rect 2926 2790 2932 2791
rect 2926 2786 2927 2790
rect 2931 2786 2932 2790
rect 2926 2785 2932 2786
rect 3030 2790 3036 2791
rect 3030 2786 3031 2790
rect 3035 2786 3036 2790
rect 3030 2785 3036 2786
rect 3134 2790 3140 2791
rect 3134 2786 3135 2790
rect 3139 2786 3140 2790
rect 3134 2785 3140 2786
rect 3238 2790 3244 2791
rect 3990 2790 3996 2791
rect 3238 2786 3239 2790
rect 3243 2786 3244 2790
rect 3238 2785 3244 2786
rect 2408 2767 2410 2785
rect 2512 2767 2514 2785
rect 2616 2767 2618 2785
rect 2720 2767 2722 2785
rect 2824 2767 2826 2785
rect 2928 2767 2930 2785
rect 3032 2767 3034 2785
rect 3136 2767 3138 2785
rect 3240 2767 3242 2785
rect 3992 2767 3994 2790
rect 2071 2766 2075 2767
rect 2071 2761 2075 2762
rect 2303 2766 2307 2767
rect 2303 2761 2307 2762
rect 2407 2766 2411 2767
rect 2407 2761 2411 2762
rect 2415 2766 2419 2767
rect 2415 2761 2419 2762
rect 2511 2766 2515 2767
rect 2511 2761 2515 2762
rect 2535 2766 2539 2767
rect 2535 2761 2539 2762
rect 2615 2766 2619 2767
rect 2615 2761 2619 2762
rect 2655 2766 2659 2767
rect 2655 2761 2659 2762
rect 2719 2766 2723 2767
rect 2719 2761 2723 2762
rect 2775 2766 2779 2767
rect 2775 2761 2779 2762
rect 2823 2766 2827 2767
rect 2823 2761 2827 2762
rect 2895 2766 2899 2767
rect 2895 2761 2899 2762
rect 2927 2766 2931 2767
rect 2927 2761 2931 2762
rect 3015 2766 3019 2767
rect 3015 2761 3019 2762
rect 3031 2766 3035 2767
rect 3031 2761 3035 2762
rect 3135 2766 3139 2767
rect 3135 2761 3139 2762
rect 3143 2766 3147 2767
rect 3143 2761 3147 2762
rect 3239 2766 3243 2767
rect 3239 2761 3243 2762
rect 3271 2766 3275 2767
rect 3271 2761 3275 2762
rect 3399 2766 3403 2767
rect 3399 2761 3403 2762
rect 3991 2766 3995 2767
rect 3991 2761 3995 2762
rect 111 2746 115 2747
rect 111 2741 115 2742
rect 151 2746 155 2747
rect 151 2741 155 2742
rect 303 2746 307 2747
rect 303 2741 307 2742
rect 311 2746 315 2747
rect 311 2741 315 2742
rect 471 2746 475 2747
rect 471 2741 475 2742
rect 623 2746 627 2747
rect 623 2741 627 2742
rect 767 2746 771 2747
rect 767 2741 771 2742
rect 903 2746 907 2747
rect 903 2741 907 2742
rect 1031 2746 1035 2747
rect 1031 2741 1035 2742
rect 1039 2746 1043 2747
rect 1039 2741 1043 2742
rect 1159 2746 1163 2747
rect 1159 2741 1163 2742
rect 1167 2746 1171 2747
rect 1167 2741 1171 2742
rect 1287 2746 1291 2747
rect 1287 2741 1291 2742
rect 1295 2746 1299 2747
rect 1295 2741 1299 2742
rect 1415 2746 1419 2747
rect 1415 2741 1419 2742
rect 1423 2746 1427 2747
rect 1423 2741 1427 2742
rect 2031 2746 2035 2747
rect 2072 2746 2074 2761
rect 2304 2751 2306 2761
rect 2416 2751 2418 2761
rect 2536 2751 2538 2761
rect 2656 2751 2658 2761
rect 2776 2751 2778 2761
rect 2896 2751 2898 2761
rect 3016 2751 3018 2761
rect 3144 2751 3146 2761
rect 3272 2751 3274 2761
rect 3400 2751 3402 2761
rect 2302 2750 2308 2751
rect 2302 2746 2303 2750
rect 2307 2746 2308 2750
rect 2031 2741 2035 2742
rect 2070 2745 2076 2746
rect 2302 2745 2308 2746
rect 2414 2750 2420 2751
rect 2414 2746 2415 2750
rect 2419 2746 2420 2750
rect 2414 2745 2420 2746
rect 2534 2750 2540 2751
rect 2534 2746 2535 2750
rect 2539 2746 2540 2750
rect 2534 2745 2540 2746
rect 2654 2750 2660 2751
rect 2654 2746 2655 2750
rect 2659 2746 2660 2750
rect 2654 2745 2660 2746
rect 2774 2750 2780 2751
rect 2774 2746 2775 2750
rect 2779 2746 2780 2750
rect 2774 2745 2780 2746
rect 2894 2750 2900 2751
rect 2894 2746 2895 2750
rect 2899 2746 2900 2750
rect 2894 2745 2900 2746
rect 3014 2750 3020 2751
rect 3014 2746 3015 2750
rect 3019 2746 3020 2750
rect 3014 2745 3020 2746
rect 3142 2750 3148 2751
rect 3142 2746 3143 2750
rect 3147 2746 3148 2750
rect 3142 2745 3148 2746
rect 3270 2750 3276 2751
rect 3270 2746 3271 2750
rect 3275 2746 3276 2750
rect 3270 2745 3276 2746
rect 3398 2750 3404 2751
rect 3398 2746 3399 2750
rect 3403 2746 3404 2750
rect 3992 2746 3994 2761
rect 3398 2745 3404 2746
rect 3990 2745 3996 2746
rect 2070 2741 2071 2745
rect 2075 2741 2076 2745
rect 112 2713 114 2741
rect 152 2732 154 2741
rect 304 2732 306 2741
rect 472 2732 474 2741
rect 624 2732 626 2741
rect 768 2732 770 2741
rect 904 2732 906 2741
rect 1040 2732 1042 2741
rect 1168 2732 1170 2741
rect 1296 2732 1298 2741
rect 1424 2732 1426 2741
rect 150 2731 156 2732
rect 150 2727 151 2731
rect 155 2727 156 2731
rect 150 2726 156 2727
rect 302 2731 308 2732
rect 302 2727 303 2731
rect 307 2727 308 2731
rect 302 2726 308 2727
rect 470 2731 476 2732
rect 470 2727 471 2731
rect 475 2727 476 2731
rect 470 2726 476 2727
rect 622 2731 628 2732
rect 622 2727 623 2731
rect 627 2727 628 2731
rect 622 2726 628 2727
rect 766 2731 772 2732
rect 766 2727 767 2731
rect 771 2727 772 2731
rect 766 2726 772 2727
rect 902 2731 908 2732
rect 902 2727 903 2731
rect 907 2727 908 2731
rect 902 2726 908 2727
rect 1038 2731 1044 2732
rect 1038 2727 1039 2731
rect 1043 2727 1044 2731
rect 1038 2726 1044 2727
rect 1166 2731 1172 2732
rect 1166 2727 1167 2731
rect 1171 2727 1172 2731
rect 1166 2726 1172 2727
rect 1294 2731 1300 2732
rect 1294 2727 1295 2731
rect 1299 2727 1300 2731
rect 1294 2726 1300 2727
rect 1422 2731 1428 2732
rect 1422 2727 1423 2731
rect 1427 2727 1428 2731
rect 1422 2726 1428 2727
rect 2032 2713 2034 2741
rect 2070 2740 2076 2741
rect 3990 2741 3991 2745
rect 3995 2741 3996 2745
rect 3990 2740 3996 2741
rect 2070 2728 2076 2729
rect 2070 2724 2071 2728
rect 2075 2724 2076 2728
rect 2070 2723 2076 2724
rect 3990 2728 3996 2729
rect 3990 2724 3991 2728
rect 3995 2724 3996 2728
rect 3990 2723 3996 2724
rect 110 2712 116 2713
rect 110 2708 111 2712
rect 115 2708 116 2712
rect 110 2707 116 2708
rect 2030 2712 2036 2713
rect 2030 2708 2031 2712
rect 2035 2708 2036 2712
rect 2030 2707 2036 2708
rect 110 2695 116 2696
rect 110 2691 111 2695
rect 115 2691 116 2695
rect 2030 2695 2036 2696
rect 2030 2691 2031 2695
rect 2035 2691 2036 2695
rect 110 2690 116 2691
rect 150 2690 156 2691
rect 112 2663 114 2690
rect 150 2686 151 2690
rect 155 2686 156 2690
rect 150 2685 156 2686
rect 302 2690 308 2691
rect 302 2686 303 2690
rect 307 2686 308 2690
rect 302 2685 308 2686
rect 470 2690 476 2691
rect 470 2686 471 2690
rect 475 2686 476 2690
rect 470 2685 476 2686
rect 622 2690 628 2691
rect 622 2686 623 2690
rect 627 2686 628 2690
rect 622 2685 628 2686
rect 766 2690 772 2691
rect 766 2686 767 2690
rect 771 2686 772 2690
rect 766 2685 772 2686
rect 902 2690 908 2691
rect 902 2686 903 2690
rect 907 2686 908 2690
rect 902 2685 908 2686
rect 1038 2690 1044 2691
rect 1038 2686 1039 2690
rect 1043 2686 1044 2690
rect 1038 2685 1044 2686
rect 1166 2690 1172 2691
rect 1166 2686 1167 2690
rect 1171 2686 1172 2690
rect 1166 2685 1172 2686
rect 1294 2690 1300 2691
rect 1294 2686 1295 2690
rect 1299 2686 1300 2690
rect 1294 2685 1300 2686
rect 1422 2690 1428 2691
rect 2030 2690 2036 2691
rect 1422 2686 1423 2690
rect 1427 2686 1428 2690
rect 1422 2685 1428 2686
rect 152 2663 154 2685
rect 304 2663 306 2685
rect 472 2663 474 2685
rect 624 2663 626 2685
rect 768 2663 770 2685
rect 904 2663 906 2685
rect 1040 2663 1042 2685
rect 1168 2663 1170 2685
rect 1296 2663 1298 2685
rect 1424 2663 1426 2685
rect 2032 2663 2034 2690
rect 2072 2679 2074 2723
rect 2302 2709 2308 2710
rect 2302 2705 2303 2709
rect 2307 2705 2308 2709
rect 2302 2704 2308 2705
rect 2414 2709 2420 2710
rect 2414 2705 2415 2709
rect 2419 2705 2420 2709
rect 2414 2704 2420 2705
rect 2534 2709 2540 2710
rect 2534 2705 2535 2709
rect 2539 2705 2540 2709
rect 2534 2704 2540 2705
rect 2654 2709 2660 2710
rect 2654 2705 2655 2709
rect 2659 2705 2660 2709
rect 2654 2704 2660 2705
rect 2774 2709 2780 2710
rect 2774 2705 2775 2709
rect 2779 2705 2780 2709
rect 2774 2704 2780 2705
rect 2894 2709 2900 2710
rect 2894 2705 2895 2709
rect 2899 2705 2900 2709
rect 2894 2704 2900 2705
rect 3014 2709 3020 2710
rect 3014 2705 3015 2709
rect 3019 2705 3020 2709
rect 3014 2704 3020 2705
rect 3142 2709 3148 2710
rect 3142 2705 3143 2709
rect 3147 2705 3148 2709
rect 3142 2704 3148 2705
rect 3270 2709 3276 2710
rect 3270 2705 3271 2709
rect 3275 2705 3276 2709
rect 3270 2704 3276 2705
rect 3398 2709 3404 2710
rect 3398 2705 3399 2709
rect 3403 2705 3404 2709
rect 3398 2704 3404 2705
rect 2304 2679 2306 2704
rect 2416 2679 2418 2704
rect 2536 2679 2538 2704
rect 2656 2679 2658 2704
rect 2776 2679 2778 2704
rect 2896 2679 2898 2704
rect 3016 2679 3018 2704
rect 3144 2679 3146 2704
rect 3272 2679 3274 2704
rect 3400 2679 3402 2704
rect 3992 2679 3994 2723
rect 2071 2678 2075 2679
rect 2071 2673 2075 2674
rect 2151 2678 2155 2679
rect 2151 2673 2155 2674
rect 2303 2678 2307 2679
rect 2303 2673 2307 2674
rect 2415 2678 2419 2679
rect 2415 2673 2419 2674
rect 2463 2678 2467 2679
rect 2463 2673 2467 2674
rect 2535 2678 2539 2679
rect 2535 2673 2539 2674
rect 2623 2678 2627 2679
rect 2623 2673 2627 2674
rect 2655 2678 2659 2679
rect 2655 2673 2659 2674
rect 2775 2678 2779 2679
rect 2775 2673 2779 2674
rect 2791 2678 2795 2679
rect 2791 2673 2795 2674
rect 2895 2678 2899 2679
rect 2895 2673 2899 2674
rect 2951 2678 2955 2679
rect 2951 2673 2955 2674
rect 3015 2678 3019 2679
rect 3015 2673 3019 2674
rect 3111 2678 3115 2679
rect 3111 2673 3115 2674
rect 3143 2678 3147 2679
rect 3143 2673 3147 2674
rect 3263 2678 3267 2679
rect 3263 2673 3267 2674
rect 3271 2678 3275 2679
rect 3271 2673 3275 2674
rect 3399 2678 3403 2679
rect 3399 2673 3403 2674
rect 3415 2678 3419 2679
rect 3415 2673 3419 2674
rect 3575 2678 3579 2679
rect 3575 2673 3579 2674
rect 3991 2678 3995 2679
rect 3991 2673 3995 2674
rect 111 2662 115 2663
rect 111 2657 115 2658
rect 151 2662 155 2663
rect 151 2657 155 2658
rect 303 2662 307 2663
rect 303 2657 307 2658
rect 319 2662 323 2663
rect 319 2657 323 2658
rect 471 2662 475 2663
rect 471 2657 475 2658
rect 511 2662 515 2663
rect 511 2657 515 2658
rect 623 2662 627 2663
rect 623 2657 627 2658
rect 703 2662 707 2663
rect 703 2657 707 2658
rect 767 2662 771 2663
rect 767 2657 771 2658
rect 887 2662 891 2663
rect 887 2657 891 2658
rect 903 2662 907 2663
rect 903 2657 907 2658
rect 1039 2662 1043 2663
rect 1039 2657 1043 2658
rect 1063 2662 1067 2663
rect 1063 2657 1067 2658
rect 1167 2662 1171 2663
rect 1167 2657 1171 2658
rect 1231 2662 1235 2663
rect 1231 2657 1235 2658
rect 1295 2662 1299 2663
rect 1295 2657 1299 2658
rect 1391 2662 1395 2663
rect 1391 2657 1395 2658
rect 1423 2662 1427 2663
rect 1423 2657 1427 2658
rect 1551 2662 1555 2663
rect 1551 2657 1555 2658
rect 1711 2662 1715 2663
rect 1711 2657 1715 2658
rect 2031 2662 2035 2663
rect 2031 2657 2035 2658
rect 112 2642 114 2657
rect 152 2647 154 2657
rect 320 2647 322 2657
rect 512 2647 514 2657
rect 704 2647 706 2657
rect 888 2647 890 2657
rect 1064 2647 1066 2657
rect 1232 2647 1234 2657
rect 1392 2647 1394 2657
rect 1552 2647 1554 2657
rect 1712 2647 1714 2657
rect 150 2646 156 2647
rect 150 2642 151 2646
rect 155 2642 156 2646
rect 110 2641 116 2642
rect 150 2641 156 2642
rect 318 2646 324 2647
rect 318 2642 319 2646
rect 323 2642 324 2646
rect 318 2641 324 2642
rect 510 2646 516 2647
rect 510 2642 511 2646
rect 515 2642 516 2646
rect 510 2641 516 2642
rect 702 2646 708 2647
rect 702 2642 703 2646
rect 707 2642 708 2646
rect 702 2641 708 2642
rect 886 2646 892 2647
rect 886 2642 887 2646
rect 891 2642 892 2646
rect 886 2641 892 2642
rect 1062 2646 1068 2647
rect 1062 2642 1063 2646
rect 1067 2642 1068 2646
rect 1062 2641 1068 2642
rect 1230 2646 1236 2647
rect 1230 2642 1231 2646
rect 1235 2642 1236 2646
rect 1230 2641 1236 2642
rect 1390 2646 1396 2647
rect 1390 2642 1391 2646
rect 1395 2642 1396 2646
rect 1390 2641 1396 2642
rect 1550 2646 1556 2647
rect 1550 2642 1551 2646
rect 1555 2642 1556 2646
rect 1550 2641 1556 2642
rect 1710 2646 1716 2647
rect 1710 2642 1711 2646
rect 1715 2642 1716 2646
rect 2032 2642 2034 2657
rect 2072 2645 2074 2673
rect 2152 2664 2154 2673
rect 2304 2664 2306 2673
rect 2464 2664 2466 2673
rect 2624 2664 2626 2673
rect 2792 2664 2794 2673
rect 2952 2664 2954 2673
rect 3112 2664 3114 2673
rect 3264 2664 3266 2673
rect 3416 2664 3418 2673
rect 3576 2664 3578 2673
rect 2150 2663 2156 2664
rect 2150 2659 2151 2663
rect 2155 2659 2156 2663
rect 2150 2658 2156 2659
rect 2302 2663 2308 2664
rect 2302 2659 2303 2663
rect 2307 2659 2308 2663
rect 2302 2658 2308 2659
rect 2462 2663 2468 2664
rect 2462 2659 2463 2663
rect 2467 2659 2468 2663
rect 2462 2658 2468 2659
rect 2622 2663 2628 2664
rect 2622 2659 2623 2663
rect 2627 2659 2628 2663
rect 2622 2658 2628 2659
rect 2790 2663 2796 2664
rect 2790 2659 2791 2663
rect 2795 2659 2796 2663
rect 2790 2658 2796 2659
rect 2950 2663 2956 2664
rect 2950 2659 2951 2663
rect 2955 2659 2956 2663
rect 2950 2658 2956 2659
rect 3110 2663 3116 2664
rect 3110 2659 3111 2663
rect 3115 2659 3116 2663
rect 3110 2658 3116 2659
rect 3262 2663 3268 2664
rect 3262 2659 3263 2663
rect 3267 2659 3268 2663
rect 3262 2658 3268 2659
rect 3414 2663 3420 2664
rect 3414 2659 3415 2663
rect 3419 2659 3420 2663
rect 3414 2658 3420 2659
rect 3574 2663 3580 2664
rect 3574 2659 3575 2663
rect 3579 2659 3580 2663
rect 3574 2658 3580 2659
rect 3992 2645 3994 2673
rect 2070 2644 2076 2645
rect 1710 2641 1716 2642
rect 2030 2641 2036 2642
rect 110 2637 111 2641
rect 115 2637 116 2641
rect 110 2636 116 2637
rect 2030 2637 2031 2641
rect 2035 2637 2036 2641
rect 2070 2640 2071 2644
rect 2075 2640 2076 2644
rect 2070 2639 2076 2640
rect 3990 2644 3996 2645
rect 3990 2640 3991 2644
rect 3995 2640 3996 2644
rect 3990 2639 3996 2640
rect 2030 2636 2036 2637
rect 2070 2627 2076 2628
rect 110 2624 116 2625
rect 110 2620 111 2624
rect 115 2620 116 2624
rect 110 2619 116 2620
rect 2030 2624 2036 2625
rect 2030 2620 2031 2624
rect 2035 2620 2036 2624
rect 2070 2623 2071 2627
rect 2075 2623 2076 2627
rect 3990 2627 3996 2628
rect 3990 2623 3991 2627
rect 3995 2623 3996 2627
rect 2070 2622 2076 2623
rect 2150 2622 2156 2623
rect 2030 2619 2036 2620
rect 112 2575 114 2619
rect 150 2605 156 2606
rect 150 2601 151 2605
rect 155 2601 156 2605
rect 150 2600 156 2601
rect 318 2605 324 2606
rect 318 2601 319 2605
rect 323 2601 324 2605
rect 318 2600 324 2601
rect 510 2605 516 2606
rect 510 2601 511 2605
rect 515 2601 516 2605
rect 510 2600 516 2601
rect 702 2605 708 2606
rect 702 2601 703 2605
rect 707 2601 708 2605
rect 702 2600 708 2601
rect 886 2605 892 2606
rect 886 2601 887 2605
rect 891 2601 892 2605
rect 886 2600 892 2601
rect 1062 2605 1068 2606
rect 1062 2601 1063 2605
rect 1067 2601 1068 2605
rect 1062 2600 1068 2601
rect 1230 2605 1236 2606
rect 1230 2601 1231 2605
rect 1235 2601 1236 2605
rect 1230 2600 1236 2601
rect 1390 2605 1396 2606
rect 1390 2601 1391 2605
rect 1395 2601 1396 2605
rect 1390 2600 1396 2601
rect 1550 2605 1556 2606
rect 1550 2601 1551 2605
rect 1555 2601 1556 2605
rect 1550 2600 1556 2601
rect 1710 2605 1716 2606
rect 1710 2601 1711 2605
rect 1715 2601 1716 2605
rect 1710 2600 1716 2601
rect 152 2575 154 2600
rect 320 2575 322 2600
rect 512 2575 514 2600
rect 704 2575 706 2600
rect 888 2575 890 2600
rect 1064 2575 1066 2600
rect 1232 2575 1234 2600
rect 1392 2575 1394 2600
rect 1552 2575 1554 2600
rect 1712 2575 1714 2600
rect 2032 2575 2034 2619
rect 2072 2599 2074 2622
rect 2150 2618 2151 2622
rect 2155 2618 2156 2622
rect 2150 2617 2156 2618
rect 2302 2622 2308 2623
rect 2302 2618 2303 2622
rect 2307 2618 2308 2622
rect 2302 2617 2308 2618
rect 2462 2622 2468 2623
rect 2462 2618 2463 2622
rect 2467 2618 2468 2622
rect 2462 2617 2468 2618
rect 2622 2622 2628 2623
rect 2622 2618 2623 2622
rect 2627 2618 2628 2622
rect 2622 2617 2628 2618
rect 2790 2622 2796 2623
rect 2790 2618 2791 2622
rect 2795 2618 2796 2622
rect 2790 2617 2796 2618
rect 2950 2622 2956 2623
rect 2950 2618 2951 2622
rect 2955 2618 2956 2622
rect 2950 2617 2956 2618
rect 3110 2622 3116 2623
rect 3110 2618 3111 2622
rect 3115 2618 3116 2622
rect 3110 2617 3116 2618
rect 3262 2622 3268 2623
rect 3262 2618 3263 2622
rect 3267 2618 3268 2622
rect 3262 2617 3268 2618
rect 3414 2622 3420 2623
rect 3414 2618 3415 2622
rect 3419 2618 3420 2622
rect 3414 2617 3420 2618
rect 3574 2622 3580 2623
rect 3990 2622 3996 2623
rect 3574 2618 3575 2622
rect 3579 2618 3580 2622
rect 3574 2617 3580 2618
rect 2152 2599 2154 2617
rect 2304 2599 2306 2617
rect 2464 2599 2466 2617
rect 2624 2599 2626 2617
rect 2792 2599 2794 2617
rect 2952 2599 2954 2617
rect 3112 2599 3114 2617
rect 3264 2599 3266 2617
rect 3416 2599 3418 2617
rect 3576 2599 3578 2617
rect 3992 2599 3994 2622
rect 2071 2598 2075 2599
rect 2071 2593 2075 2594
rect 2111 2598 2115 2599
rect 2111 2593 2115 2594
rect 2151 2598 2155 2599
rect 2151 2593 2155 2594
rect 2303 2598 2307 2599
rect 2303 2593 2307 2594
rect 2327 2598 2331 2599
rect 2327 2593 2331 2594
rect 2463 2598 2467 2599
rect 2463 2593 2467 2594
rect 2559 2598 2563 2599
rect 2559 2593 2563 2594
rect 2623 2598 2627 2599
rect 2623 2593 2627 2594
rect 2783 2598 2787 2599
rect 2783 2593 2787 2594
rect 2791 2598 2795 2599
rect 2791 2593 2795 2594
rect 2951 2598 2955 2599
rect 2951 2593 2955 2594
rect 2999 2598 3003 2599
rect 2999 2593 3003 2594
rect 3111 2598 3115 2599
rect 3111 2593 3115 2594
rect 3199 2598 3203 2599
rect 3199 2593 3203 2594
rect 3263 2598 3267 2599
rect 3263 2593 3267 2594
rect 3383 2598 3387 2599
rect 3383 2593 3387 2594
rect 3415 2598 3419 2599
rect 3415 2593 3419 2594
rect 3559 2598 3563 2599
rect 3559 2593 3563 2594
rect 3575 2598 3579 2599
rect 3575 2593 3579 2594
rect 3735 2598 3739 2599
rect 3735 2593 3739 2594
rect 3895 2598 3899 2599
rect 3895 2593 3899 2594
rect 3991 2598 3995 2599
rect 3991 2593 3995 2594
rect 2072 2578 2074 2593
rect 2112 2583 2114 2593
rect 2328 2583 2330 2593
rect 2560 2583 2562 2593
rect 2784 2583 2786 2593
rect 3000 2583 3002 2593
rect 3200 2583 3202 2593
rect 3384 2583 3386 2593
rect 3560 2583 3562 2593
rect 3736 2583 3738 2593
rect 3896 2583 3898 2593
rect 2110 2582 2116 2583
rect 2110 2578 2111 2582
rect 2115 2578 2116 2582
rect 2070 2577 2076 2578
rect 2110 2577 2116 2578
rect 2326 2582 2332 2583
rect 2326 2578 2327 2582
rect 2331 2578 2332 2582
rect 2326 2577 2332 2578
rect 2558 2582 2564 2583
rect 2558 2578 2559 2582
rect 2563 2578 2564 2582
rect 2558 2577 2564 2578
rect 2782 2582 2788 2583
rect 2782 2578 2783 2582
rect 2787 2578 2788 2582
rect 2782 2577 2788 2578
rect 2998 2582 3004 2583
rect 2998 2578 2999 2582
rect 3003 2578 3004 2582
rect 2998 2577 3004 2578
rect 3198 2582 3204 2583
rect 3198 2578 3199 2582
rect 3203 2578 3204 2582
rect 3198 2577 3204 2578
rect 3382 2582 3388 2583
rect 3382 2578 3383 2582
rect 3387 2578 3388 2582
rect 3382 2577 3388 2578
rect 3558 2582 3564 2583
rect 3558 2578 3559 2582
rect 3563 2578 3564 2582
rect 3558 2577 3564 2578
rect 3734 2582 3740 2583
rect 3734 2578 3735 2582
rect 3739 2578 3740 2582
rect 3734 2577 3740 2578
rect 3894 2582 3900 2583
rect 3894 2578 3895 2582
rect 3899 2578 3900 2582
rect 3992 2578 3994 2593
rect 3894 2577 3900 2578
rect 3990 2577 3996 2578
rect 111 2574 115 2575
rect 111 2569 115 2570
rect 151 2574 155 2575
rect 151 2569 155 2570
rect 279 2574 283 2575
rect 279 2569 283 2570
rect 319 2574 323 2575
rect 319 2569 323 2570
rect 463 2574 467 2575
rect 463 2569 467 2570
rect 511 2574 515 2575
rect 511 2569 515 2570
rect 663 2574 667 2575
rect 663 2569 667 2570
rect 703 2574 707 2575
rect 703 2569 707 2570
rect 863 2574 867 2575
rect 863 2569 867 2570
rect 887 2574 891 2575
rect 887 2569 891 2570
rect 1063 2574 1067 2575
rect 1063 2569 1067 2570
rect 1231 2574 1235 2575
rect 1231 2569 1235 2570
rect 1255 2574 1259 2575
rect 1255 2569 1259 2570
rect 1391 2574 1395 2575
rect 1391 2569 1395 2570
rect 1431 2574 1435 2575
rect 1431 2569 1435 2570
rect 1551 2574 1555 2575
rect 1551 2569 1555 2570
rect 1607 2574 1611 2575
rect 1607 2569 1611 2570
rect 1711 2574 1715 2575
rect 1711 2569 1715 2570
rect 1783 2574 1787 2575
rect 1783 2569 1787 2570
rect 1935 2574 1939 2575
rect 1935 2569 1939 2570
rect 2031 2574 2035 2575
rect 2070 2573 2071 2577
rect 2075 2573 2076 2577
rect 2070 2572 2076 2573
rect 3990 2573 3991 2577
rect 3995 2573 3996 2577
rect 3990 2572 3996 2573
rect 2031 2569 2035 2570
rect 112 2541 114 2569
rect 280 2560 282 2569
rect 464 2560 466 2569
rect 664 2560 666 2569
rect 864 2560 866 2569
rect 1064 2560 1066 2569
rect 1256 2560 1258 2569
rect 1432 2560 1434 2569
rect 1608 2560 1610 2569
rect 1784 2560 1786 2569
rect 1936 2560 1938 2569
rect 278 2559 284 2560
rect 278 2555 279 2559
rect 283 2555 284 2559
rect 278 2554 284 2555
rect 462 2559 468 2560
rect 462 2555 463 2559
rect 467 2555 468 2559
rect 462 2554 468 2555
rect 662 2559 668 2560
rect 662 2555 663 2559
rect 667 2555 668 2559
rect 662 2554 668 2555
rect 862 2559 868 2560
rect 862 2555 863 2559
rect 867 2555 868 2559
rect 862 2554 868 2555
rect 1062 2559 1068 2560
rect 1062 2555 1063 2559
rect 1067 2555 1068 2559
rect 1062 2554 1068 2555
rect 1254 2559 1260 2560
rect 1254 2555 1255 2559
rect 1259 2555 1260 2559
rect 1254 2554 1260 2555
rect 1430 2559 1436 2560
rect 1430 2555 1431 2559
rect 1435 2555 1436 2559
rect 1430 2554 1436 2555
rect 1606 2559 1612 2560
rect 1606 2555 1607 2559
rect 1611 2555 1612 2559
rect 1606 2554 1612 2555
rect 1782 2559 1788 2560
rect 1782 2555 1783 2559
rect 1787 2555 1788 2559
rect 1782 2554 1788 2555
rect 1934 2559 1940 2560
rect 1934 2555 1935 2559
rect 1939 2555 1940 2559
rect 1934 2554 1940 2555
rect 2032 2541 2034 2569
rect 2070 2560 2076 2561
rect 2070 2556 2071 2560
rect 2075 2556 2076 2560
rect 2070 2555 2076 2556
rect 3990 2560 3996 2561
rect 3990 2556 3991 2560
rect 3995 2556 3996 2560
rect 3990 2555 3996 2556
rect 110 2540 116 2541
rect 110 2536 111 2540
rect 115 2536 116 2540
rect 110 2535 116 2536
rect 2030 2540 2036 2541
rect 2030 2536 2031 2540
rect 2035 2536 2036 2540
rect 2030 2535 2036 2536
rect 2072 2527 2074 2555
rect 2110 2541 2116 2542
rect 2110 2537 2111 2541
rect 2115 2537 2116 2541
rect 2110 2536 2116 2537
rect 2326 2541 2332 2542
rect 2326 2537 2327 2541
rect 2331 2537 2332 2541
rect 2326 2536 2332 2537
rect 2558 2541 2564 2542
rect 2558 2537 2559 2541
rect 2563 2537 2564 2541
rect 2558 2536 2564 2537
rect 2782 2541 2788 2542
rect 2782 2537 2783 2541
rect 2787 2537 2788 2541
rect 2782 2536 2788 2537
rect 2998 2541 3004 2542
rect 2998 2537 2999 2541
rect 3003 2537 3004 2541
rect 2998 2536 3004 2537
rect 3198 2541 3204 2542
rect 3198 2537 3199 2541
rect 3203 2537 3204 2541
rect 3198 2536 3204 2537
rect 3382 2541 3388 2542
rect 3382 2537 3383 2541
rect 3387 2537 3388 2541
rect 3382 2536 3388 2537
rect 3558 2541 3564 2542
rect 3558 2537 3559 2541
rect 3563 2537 3564 2541
rect 3558 2536 3564 2537
rect 3734 2541 3740 2542
rect 3734 2537 3735 2541
rect 3739 2537 3740 2541
rect 3734 2536 3740 2537
rect 3894 2541 3900 2542
rect 3894 2537 3895 2541
rect 3899 2537 3900 2541
rect 3894 2536 3900 2537
rect 2112 2527 2114 2536
rect 2328 2527 2330 2536
rect 2560 2527 2562 2536
rect 2784 2527 2786 2536
rect 3000 2527 3002 2536
rect 3200 2527 3202 2536
rect 3384 2527 3386 2536
rect 3560 2527 3562 2536
rect 3736 2527 3738 2536
rect 3896 2527 3898 2536
rect 3992 2527 3994 2555
rect 2071 2526 2075 2527
rect 110 2523 116 2524
rect 110 2519 111 2523
rect 115 2519 116 2523
rect 2030 2523 2036 2524
rect 2030 2519 2031 2523
rect 2035 2519 2036 2523
rect 2071 2521 2075 2522
rect 2111 2526 2115 2527
rect 2111 2521 2115 2522
rect 2255 2526 2259 2527
rect 2255 2521 2259 2522
rect 2327 2526 2331 2527
rect 2327 2521 2331 2522
rect 2439 2526 2443 2527
rect 2439 2521 2443 2522
rect 2559 2526 2563 2527
rect 2559 2521 2563 2522
rect 2631 2526 2635 2527
rect 2631 2521 2635 2522
rect 2783 2526 2787 2527
rect 2783 2521 2787 2522
rect 2823 2526 2827 2527
rect 2823 2521 2827 2522
rect 2999 2526 3003 2527
rect 2999 2521 3003 2522
rect 3007 2526 3011 2527
rect 3007 2521 3011 2522
rect 3175 2526 3179 2527
rect 3175 2521 3179 2522
rect 3199 2526 3203 2527
rect 3199 2521 3203 2522
rect 3335 2526 3339 2527
rect 3335 2521 3339 2522
rect 3383 2526 3387 2527
rect 3383 2521 3387 2522
rect 3487 2526 3491 2527
rect 3487 2521 3491 2522
rect 3559 2526 3563 2527
rect 3559 2521 3563 2522
rect 3631 2526 3635 2527
rect 3631 2521 3635 2522
rect 3735 2526 3739 2527
rect 3735 2521 3739 2522
rect 3775 2526 3779 2527
rect 3775 2521 3779 2522
rect 3895 2526 3899 2527
rect 3895 2521 3899 2522
rect 3991 2526 3995 2527
rect 3991 2521 3995 2522
rect 110 2518 116 2519
rect 278 2518 284 2519
rect 112 2487 114 2518
rect 278 2514 279 2518
rect 283 2514 284 2518
rect 278 2513 284 2514
rect 462 2518 468 2519
rect 462 2514 463 2518
rect 467 2514 468 2518
rect 462 2513 468 2514
rect 662 2518 668 2519
rect 662 2514 663 2518
rect 667 2514 668 2518
rect 662 2513 668 2514
rect 862 2518 868 2519
rect 862 2514 863 2518
rect 867 2514 868 2518
rect 862 2513 868 2514
rect 1062 2518 1068 2519
rect 1062 2514 1063 2518
rect 1067 2514 1068 2518
rect 1062 2513 1068 2514
rect 1254 2518 1260 2519
rect 1254 2514 1255 2518
rect 1259 2514 1260 2518
rect 1254 2513 1260 2514
rect 1430 2518 1436 2519
rect 1430 2514 1431 2518
rect 1435 2514 1436 2518
rect 1430 2513 1436 2514
rect 1606 2518 1612 2519
rect 1606 2514 1607 2518
rect 1611 2514 1612 2518
rect 1606 2513 1612 2514
rect 1782 2518 1788 2519
rect 1782 2514 1783 2518
rect 1787 2514 1788 2518
rect 1782 2513 1788 2514
rect 1934 2518 1940 2519
rect 2030 2518 2036 2519
rect 1934 2514 1935 2518
rect 1939 2514 1940 2518
rect 1934 2513 1940 2514
rect 280 2487 282 2513
rect 464 2487 466 2513
rect 664 2487 666 2513
rect 864 2487 866 2513
rect 1064 2487 1066 2513
rect 1256 2487 1258 2513
rect 1432 2487 1434 2513
rect 1608 2487 1610 2513
rect 1784 2487 1786 2513
rect 1936 2487 1938 2513
rect 2032 2487 2034 2518
rect 2072 2493 2074 2521
rect 2112 2512 2114 2521
rect 2256 2512 2258 2521
rect 2440 2512 2442 2521
rect 2632 2512 2634 2521
rect 2824 2512 2826 2521
rect 3008 2512 3010 2521
rect 3176 2512 3178 2521
rect 3336 2512 3338 2521
rect 3488 2512 3490 2521
rect 3632 2512 3634 2521
rect 3776 2512 3778 2521
rect 3896 2512 3898 2521
rect 2110 2511 2116 2512
rect 2110 2507 2111 2511
rect 2115 2507 2116 2511
rect 2110 2506 2116 2507
rect 2254 2511 2260 2512
rect 2254 2507 2255 2511
rect 2259 2507 2260 2511
rect 2254 2506 2260 2507
rect 2438 2511 2444 2512
rect 2438 2507 2439 2511
rect 2443 2507 2444 2511
rect 2438 2506 2444 2507
rect 2630 2511 2636 2512
rect 2630 2507 2631 2511
rect 2635 2507 2636 2511
rect 2630 2506 2636 2507
rect 2822 2511 2828 2512
rect 2822 2507 2823 2511
rect 2827 2507 2828 2511
rect 2822 2506 2828 2507
rect 3006 2511 3012 2512
rect 3006 2507 3007 2511
rect 3011 2507 3012 2511
rect 3006 2506 3012 2507
rect 3174 2511 3180 2512
rect 3174 2507 3175 2511
rect 3179 2507 3180 2511
rect 3174 2506 3180 2507
rect 3334 2511 3340 2512
rect 3334 2507 3335 2511
rect 3339 2507 3340 2511
rect 3334 2506 3340 2507
rect 3486 2511 3492 2512
rect 3486 2507 3487 2511
rect 3491 2507 3492 2511
rect 3486 2506 3492 2507
rect 3630 2511 3636 2512
rect 3630 2507 3631 2511
rect 3635 2507 3636 2511
rect 3630 2506 3636 2507
rect 3774 2511 3780 2512
rect 3774 2507 3775 2511
rect 3779 2507 3780 2511
rect 3774 2506 3780 2507
rect 3894 2511 3900 2512
rect 3894 2507 3895 2511
rect 3899 2507 3900 2511
rect 3894 2506 3900 2507
rect 3992 2493 3994 2521
rect 2070 2492 2076 2493
rect 2070 2488 2071 2492
rect 2075 2488 2076 2492
rect 2070 2487 2076 2488
rect 3990 2492 3996 2493
rect 3990 2488 3991 2492
rect 3995 2488 3996 2492
rect 3990 2487 3996 2488
rect 111 2486 115 2487
rect 111 2481 115 2482
rect 279 2486 283 2487
rect 279 2481 283 2482
rect 311 2486 315 2487
rect 311 2481 315 2482
rect 463 2486 467 2487
rect 463 2481 467 2482
rect 471 2486 475 2487
rect 471 2481 475 2482
rect 647 2486 651 2487
rect 647 2481 651 2482
rect 663 2486 667 2487
rect 663 2481 667 2482
rect 831 2486 835 2487
rect 831 2481 835 2482
rect 863 2486 867 2487
rect 863 2481 867 2482
rect 1015 2486 1019 2487
rect 1015 2481 1019 2482
rect 1063 2486 1067 2487
rect 1063 2481 1067 2482
rect 1191 2486 1195 2487
rect 1191 2481 1195 2482
rect 1255 2486 1259 2487
rect 1255 2481 1259 2482
rect 1367 2486 1371 2487
rect 1367 2481 1371 2482
rect 1431 2486 1435 2487
rect 1431 2481 1435 2482
rect 1535 2486 1539 2487
rect 1535 2481 1539 2482
rect 1607 2486 1611 2487
rect 1607 2481 1611 2482
rect 1703 2486 1707 2487
rect 1703 2481 1707 2482
rect 1783 2486 1787 2487
rect 1783 2481 1787 2482
rect 1871 2486 1875 2487
rect 1871 2481 1875 2482
rect 1935 2486 1939 2487
rect 1935 2481 1939 2482
rect 2031 2486 2035 2487
rect 2031 2481 2035 2482
rect 112 2466 114 2481
rect 312 2471 314 2481
rect 472 2471 474 2481
rect 648 2471 650 2481
rect 832 2471 834 2481
rect 1016 2471 1018 2481
rect 1192 2471 1194 2481
rect 1368 2471 1370 2481
rect 1536 2471 1538 2481
rect 1704 2471 1706 2481
rect 1872 2471 1874 2481
rect 310 2470 316 2471
rect 310 2466 311 2470
rect 315 2466 316 2470
rect 110 2465 116 2466
rect 310 2465 316 2466
rect 470 2470 476 2471
rect 470 2466 471 2470
rect 475 2466 476 2470
rect 470 2465 476 2466
rect 646 2470 652 2471
rect 646 2466 647 2470
rect 651 2466 652 2470
rect 646 2465 652 2466
rect 830 2470 836 2471
rect 830 2466 831 2470
rect 835 2466 836 2470
rect 830 2465 836 2466
rect 1014 2470 1020 2471
rect 1014 2466 1015 2470
rect 1019 2466 1020 2470
rect 1014 2465 1020 2466
rect 1190 2470 1196 2471
rect 1190 2466 1191 2470
rect 1195 2466 1196 2470
rect 1190 2465 1196 2466
rect 1366 2470 1372 2471
rect 1366 2466 1367 2470
rect 1371 2466 1372 2470
rect 1366 2465 1372 2466
rect 1534 2470 1540 2471
rect 1534 2466 1535 2470
rect 1539 2466 1540 2470
rect 1534 2465 1540 2466
rect 1702 2470 1708 2471
rect 1702 2466 1703 2470
rect 1707 2466 1708 2470
rect 1702 2465 1708 2466
rect 1870 2470 1876 2471
rect 1870 2466 1871 2470
rect 1875 2466 1876 2470
rect 2032 2466 2034 2481
rect 2070 2475 2076 2476
rect 2070 2471 2071 2475
rect 2075 2471 2076 2475
rect 3990 2475 3996 2476
rect 3990 2471 3991 2475
rect 3995 2471 3996 2475
rect 2070 2470 2076 2471
rect 2110 2470 2116 2471
rect 1870 2465 1876 2466
rect 2030 2465 2036 2466
rect 110 2461 111 2465
rect 115 2461 116 2465
rect 110 2460 116 2461
rect 2030 2461 2031 2465
rect 2035 2461 2036 2465
rect 2030 2460 2036 2461
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 110 2443 116 2444
rect 2030 2448 2036 2449
rect 2030 2444 2031 2448
rect 2035 2444 2036 2448
rect 2072 2447 2074 2470
rect 2110 2466 2111 2470
rect 2115 2466 2116 2470
rect 2110 2465 2116 2466
rect 2254 2470 2260 2471
rect 2254 2466 2255 2470
rect 2259 2466 2260 2470
rect 2254 2465 2260 2466
rect 2438 2470 2444 2471
rect 2438 2466 2439 2470
rect 2443 2466 2444 2470
rect 2438 2465 2444 2466
rect 2630 2470 2636 2471
rect 2630 2466 2631 2470
rect 2635 2466 2636 2470
rect 2630 2465 2636 2466
rect 2822 2470 2828 2471
rect 2822 2466 2823 2470
rect 2827 2466 2828 2470
rect 2822 2465 2828 2466
rect 3006 2470 3012 2471
rect 3006 2466 3007 2470
rect 3011 2466 3012 2470
rect 3006 2465 3012 2466
rect 3174 2470 3180 2471
rect 3174 2466 3175 2470
rect 3179 2466 3180 2470
rect 3174 2465 3180 2466
rect 3334 2470 3340 2471
rect 3334 2466 3335 2470
rect 3339 2466 3340 2470
rect 3334 2465 3340 2466
rect 3486 2470 3492 2471
rect 3486 2466 3487 2470
rect 3491 2466 3492 2470
rect 3486 2465 3492 2466
rect 3630 2470 3636 2471
rect 3630 2466 3631 2470
rect 3635 2466 3636 2470
rect 3630 2465 3636 2466
rect 3774 2470 3780 2471
rect 3774 2466 3775 2470
rect 3779 2466 3780 2470
rect 3774 2465 3780 2466
rect 3894 2470 3900 2471
rect 3990 2470 3996 2471
rect 3894 2466 3895 2470
rect 3899 2466 3900 2470
rect 3894 2465 3900 2466
rect 2112 2447 2114 2465
rect 2256 2447 2258 2465
rect 2440 2447 2442 2465
rect 2632 2447 2634 2465
rect 2824 2447 2826 2465
rect 3008 2447 3010 2465
rect 3176 2447 3178 2465
rect 3336 2447 3338 2465
rect 3488 2447 3490 2465
rect 3632 2447 3634 2465
rect 3776 2447 3778 2465
rect 3896 2447 3898 2465
rect 3992 2447 3994 2470
rect 2030 2443 2036 2444
rect 2071 2446 2075 2447
rect 112 2403 114 2443
rect 310 2429 316 2430
rect 310 2425 311 2429
rect 315 2425 316 2429
rect 310 2424 316 2425
rect 470 2429 476 2430
rect 470 2425 471 2429
rect 475 2425 476 2429
rect 470 2424 476 2425
rect 646 2429 652 2430
rect 646 2425 647 2429
rect 651 2425 652 2429
rect 646 2424 652 2425
rect 830 2429 836 2430
rect 830 2425 831 2429
rect 835 2425 836 2429
rect 830 2424 836 2425
rect 1014 2429 1020 2430
rect 1014 2425 1015 2429
rect 1019 2425 1020 2429
rect 1014 2424 1020 2425
rect 1190 2429 1196 2430
rect 1190 2425 1191 2429
rect 1195 2425 1196 2429
rect 1190 2424 1196 2425
rect 1366 2429 1372 2430
rect 1366 2425 1367 2429
rect 1371 2425 1372 2429
rect 1366 2424 1372 2425
rect 1534 2429 1540 2430
rect 1534 2425 1535 2429
rect 1539 2425 1540 2429
rect 1534 2424 1540 2425
rect 1702 2429 1708 2430
rect 1702 2425 1703 2429
rect 1707 2425 1708 2429
rect 1702 2424 1708 2425
rect 1870 2429 1876 2430
rect 1870 2425 1871 2429
rect 1875 2425 1876 2429
rect 1870 2424 1876 2425
rect 312 2403 314 2424
rect 472 2403 474 2424
rect 648 2403 650 2424
rect 832 2403 834 2424
rect 1016 2403 1018 2424
rect 1192 2403 1194 2424
rect 1368 2403 1370 2424
rect 1536 2403 1538 2424
rect 1704 2403 1706 2424
rect 1872 2403 1874 2424
rect 2032 2403 2034 2443
rect 2071 2441 2075 2442
rect 2111 2446 2115 2447
rect 2111 2441 2115 2442
rect 2255 2446 2259 2447
rect 2255 2441 2259 2442
rect 2311 2446 2315 2447
rect 2311 2441 2315 2442
rect 2439 2446 2443 2447
rect 2439 2441 2443 2442
rect 2535 2446 2539 2447
rect 2535 2441 2539 2442
rect 2631 2446 2635 2447
rect 2631 2441 2635 2442
rect 2751 2446 2755 2447
rect 2751 2441 2755 2442
rect 2823 2446 2827 2447
rect 2823 2441 2827 2442
rect 2951 2446 2955 2447
rect 2951 2441 2955 2442
rect 3007 2446 3011 2447
rect 3007 2441 3011 2442
rect 3135 2446 3139 2447
rect 3135 2441 3139 2442
rect 3175 2446 3179 2447
rect 3175 2441 3179 2442
rect 3311 2446 3315 2447
rect 3311 2441 3315 2442
rect 3335 2446 3339 2447
rect 3335 2441 3339 2442
rect 3471 2446 3475 2447
rect 3471 2441 3475 2442
rect 3487 2446 3491 2447
rect 3487 2441 3491 2442
rect 3623 2446 3627 2447
rect 3623 2441 3627 2442
rect 3631 2446 3635 2447
rect 3631 2441 3635 2442
rect 3767 2446 3771 2447
rect 3767 2441 3771 2442
rect 3775 2446 3779 2447
rect 3775 2441 3779 2442
rect 3895 2446 3899 2447
rect 3895 2441 3899 2442
rect 3991 2446 3995 2447
rect 3991 2441 3995 2442
rect 2072 2426 2074 2441
rect 2112 2431 2114 2441
rect 2312 2431 2314 2441
rect 2536 2431 2538 2441
rect 2752 2431 2754 2441
rect 2952 2431 2954 2441
rect 3136 2431 3138 2441
rect 3312 2431 3314 2441
rect 3472 2431 3474 2441
rect 3624 2431 3626 2441
rect 3768 2431 3770 2441
rect 3896 2431 3898 2441
rect 2110 2430 2116 2431
rect 2110 2426 2111 2430
rect 2115 2426 2116 2430
rect 2070 2425 2076 2426
rect 2110 2425 2116 2426
rect 2310 2430 2316 2431
rect 2310 2426 2311 2430
rect 2315 2426 2316 2430
rect 2310 2425 2316 2426
rect 2534 2430 2540 2431
rect 2534 2426 2535 2430
rect 2539 2426 2540 2430
rect 2534 2425 2540 2426
rect 2750 2430 2756 2431
rect 2750 2426 2751 2430
rect 2755 2426 2756 2430
rect 2750 2425 2756 2426
rect 2950 2430 2956 2431
rect 2950 2426 2951 2430
rect 2955 2426 2956 2430
rect 2950 2425 2956 2426
rect 3134 2430 3140 2431
rect 3134 2426 3135 2430
rect 3139 2426 3140 2430
rect 3134 2425 3140 2426
rect 3310 2430 3316 2431
rect 3310 2426 3311 2430
rect 3315 2426 3316 2430
rect 3310 2425 3316 2426
rect 3470 2430 3476 2431
rect 3470 2426 3471 2430
rect 3475 2426 3476 2430
rect 3470 2425 3476 2426
rect 3622 2430 3628 2431
rect 3622 2426 3623 2430
rect 3627 2426 3628 2430
rect 3622 2425 3628 2426
rect 3766 2430 3772 2431
rect 3766 2426 3767 2430
rect 3771 2426 3772 2430
rect 3766 2425 3772 2426
rect 3894 2430 3900 2431
rect 3894 2426 3895 2430
rect 3899 2426 3900 2430
rect 3992 2426 3994 2441
rect 3894 2425 3900 2426
rect 3990 2425 3996 2426
rect 2070 2421 2071 2425
rect 2075 2421 2076 2425
rect 2070 2420 2076 2421
rect 3990 2421 3991 2425
rect 3995 2421 3996 2425
rect 3990 2420 3996 2421
rect 2070 2408 2076 2409
rect 2070 2404 2071 2408
rect 2075 2404 2076 2408
rect 2070 2403 2076 2404
rect 3990 2408 3996 2409
rect 3990 2404 3991 2408
rect 3995 2404 3996 2408
rect 3990 2403 3996 2404
rect 111 2402 115 2403
rect 111 2397 115 2398
rect 207 2402 211 2403
rect 207 2397 211 2398
rect 311 2402 315 2403
rect 311 2397 315 2398
rect 351 2402 355 2403
rect 351 2397 355 2398
rect 471 2402 475 2403
rect 471 2397 475 2398
rect 503 2402 507 2403
rect 503 2397 507 2398
rect 647 2402 651 2403
rect 647 2397 651 2398
rect 655 2402 659 2403
rect 655 2397 659 2398
rect 815 2402 819 2403
rect 815 2397 819 2398
rect 831 2402 835 2403
rect 831 2397 835 2398
rect 967 2402 971 2403
rect 967 2397 971 2398
rect 1015 2402 1019 2403
rect 1015 2397 1019 2398
rect 1119 2402 1123 2403
rect 1119 2397 1123 2398
rect 1191 2402 1195 2403
rect 1191 2397 1195 2398
rect 1263 2402 1267 2403
rect 1263 2397 1267 2398
rect 1367 2402 1371 2403
rect 1367 2397 1371 2398
rect 1415 2402 1419 2403
rect 1415 2397 1419 2398
rect 1535 2402 1539 2403
rect 1535 2397 1539 2398
rect 1567 2402 1571 2403
rect 1567 2397 1571 2398
rect 1703 2402 1707 2403
rect 1703 2397 1707 2398
rect 1871 2402 1875 2403
rect 1871 2397 1875 2398
rect 2031 2402 2035 2403
rect 2031 2397 2035 2398
rect 112 2369 114 2397
rect 208 2388 210 2397
rect 352 2388 354 2397
rect 504 2388 506 2397
rect 656 2388 658 2397
rect 816 2388 818 2397
rect 968 2388 970 2397
rect 1120 2388 1122 2397
rect 1264 2388 1266 2397
rect 1416 2388 1418 2397
rect 1568 2388 1570 2397
rect 206 2387 212 2388
rect 206 2383 207 2387
rect 211 2383 212 2387
rect 206 2382 212 2383
rect 350 2387 356 2388
rect 350 2383 351 2387
rect 355 2383 356 2387
rect 350 2382 356 2383
rect 502 2387 508 2388
rect 502 2383 503 2387
rect 507 2383 508 2387
rect 502 2382 508 2383
rect 654 2387 660 2388
rect 654 2383 655 2387
rect 659 2383 660 2387
rect 654 2382 660 2383
rect 814 2387 820 2388
rect 814 2383 815 2387
rect 819 2383 820 2387
rect 814 2382 820 2383
rect 966 2387 972 2388
rect 966 2383 967 2387
rect 971 2383 972 2387
rect 966 2382 972 2383
rect 1118 2387 1124 2388
rect 1118 2383 1119 2387
rect 1123 2383 1124 2387
rect 1118 2382 1124 2383
rect 1262 2387 1268 2388
rect 1262 2383 1263 2387
rect 1267 2383 1268 2387
rect 1262 2382 1268 2383
rect 1414 2387 1420 2388
rect 1414 2383 1415 2387
rect 1419 2383 1420 2387
rect 1414 2382 1420 2383
rect 1566 2387 1572 2388
rect 1566 2383 1567 2387
rect 1571 2383 1572 2387
rect 1566 2382 1572 2383
rect 2032 2369 2034 2397
rect 2072 2375 2074 2403
rect 2110 2389 2116 2390
rect 2110 2385 2111 2389
rect 2115 2385 2116 2389
rect 2110 2384 2116 2385
rect 2310 2389 2316 2390
rect 2310 2385 2311 2389
rect 2315 2385 2316 2389
rect 2310 2384 2316 2385
rect 2534 2389 2540 2390
rect 2534 2385 2535 2389
rect 2539 2385 2540 2389
rect 2534 2384 2540 2385
rect 2750 2389 2756 2390
rect 2750 2385 2751 2389
rect 2755 2385 2756 2389
rect 2750 2384 2756 2385
rect 2950 2389 2956 2390
rect 2950 2385 2951 2389
rect 2955 2385 2956 2389
rect 2950 2384 2956 2385
rect 3134 2389 3140 2390
rect 3134 2385 3135 2389
rect 3139 2385 3140 2389
rect 3134 2384 3140 2385
rect 3310 2389 3316 2390
rect 3310 2385 3311 2389
rect 3315 2385 3316 2389
rect 3310 2384 3316 2385
rect 3470 2389 3476 2390
rect 3470 2385 3471 2389
rect 3475 2385 3476 2389
rect 3470 2384 3476 2385
rect 3622 2389 3628 2390
rect 3622 2385 3623 2389
rect 3627 2385 3628 2389
rect 3622 2384 3628 2385
rect 3766 2389 3772 2390
rect 3766 2385 3767 2389
rect 3771 2385 3772 2389
rect 3766 2384 3772 2385
rect 3894 2389 3900 2390
rect 3894 2385 3895 2389
rect 3899 2385 3900 2389
rect 3894 2384 3900 2385
rect 2112 2375 2114 2384
rect 2312 2375 2314 2384
rect 2536 2375 2538 2384
rect 2752 2375 2754 2384
rect 2952 2375 2954 2384
rect 3136 2375 3138 2384
rect 3312 2375 3314 2384
rect 3472 2375 3474 2384
rect 3624 2375 3626 2384
rect 3768 2375 3770 2384
rect 3896 2375 3898 2384
rect 3992 2375 3994 2403
rect 2071 2374 2075 2375
rect 2071 2369 2075 2370
rect 2111 2374 2115 2375
rect 2111 2369 2115 2370
rect 2311 2374 2315 2375
rect 2311 2369 2315 2370
rect 2327 2374 2331 2375
rect 2327 2369 2331 2370
rect 2535 2374 2539 2375
rect 2535 2369 2539 2370
rect 2559 2374 2563 2375
rect 2559 2369 2563 2370
rect 2751 2374 2755 2375
rect 2751 2369 2755 2370
rect 2783 2374 2787 2375
rect 2783 2369 2787 2370
rect 2951 2374 2955 2375
rect 2951 2369 2955 2370
rect 2999 2374 3003 2375
rect 2999 2369 3003 2370
rect 3135 2374 3139 2375
rect 3135 2369 3139 2370
rect 3191 2374 3195 2375
rect 3191 2369 3195 2370
rect 3311 2374 3315 2375
rect 3311 2369 3315 2370
rect 3375 2374 3379 2375
rect 3375 2369 3379 2370
rect 3471 2374 3475 2375
rect 3471 2369 3475 2370
rect 3543 2374 3547 2375
rect 3543 2369 3547 2370
rect 3623 2374 3627 2375
rect 3623 2369 3627 2370
rect 3711 2374 3715 2375
rect 3711 2369 3715 2370
rect 3767 2374 3771 2375
rect 3767 2369 3771 2370
rect 3887 2374 3891 2375
rect 3887 2369 3891 2370
rect 3895 2374 3899 2375
rect 3895 2369 3899 2370
rect 3991 2374 3995 2375
rect 3991 2369 3995 2370
rect 110 2368 116 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 2030 2368 2036 2369
rect 2030 2364 2031 2368
rect 2035 2364 2036 2368
rect 2030 2363 2036 2364
rect 110 2351 116 2352
rect 110 2347 111 2351
rect 115 2347 116 2351
rect 2030 2351 2036 2352
rect 2030 2347 2031 2351
rect 2035 2347 2036 2351
rect 110 2346 116 2347
rect 206 2346 212 2347
rect 112 2319 114 2346
rect 206 2342 207 2346
rect 211 2342 212 2346
rect 206 2341 212 2342
rect 350 2346 356 2347
rect 350 2342 351 2346
rect 355 2342 356 2346
rect 350 2341 356 2342
rect 502 2346 508 2347
rect 502 2342 503 2346
rect 507 2342 508 2346
rect 502 2341 508 2342
rect 654 2346 660 2347
rect 654 2342 655 2346
rect 659 2342 660 2346
rect 654 2341 660 2342
rect 814 2346 820 2347
rect 814 2342 815 2346
rect 819 2342 820 2346
rect 814 2341 820 2342
rect 966 2346 972 2347
rect 966 2342 967 2346
rect 971 2342 972 2346
rect 966 2341 972 2342
rect 1118 2346 1124 2347
rect 1118 2342 1119 2346
rect 1123 2342 1124 2346
rect 1118 2341 1124 2342
rect 1262 2346 1268 2347
rect 1262 2342 1263 2346
rect 1267 2342 1268 2346
rect 1262 2341 1268 2342
rect 1414 2346 1420 2347
rect 1414 2342 1415 2346
rect 1419 2342 1420 2346
rect 1414 2341 1420 2342
rect 1566 2346 1572 2347
rect 2030 2346 2036 2347
rect 1566 2342 1567 2346
rect 1571 2342 1572 2346
rect 1566 2341 1572 2342
rect 208 2319 210 2341
rect 352 2319 354 2341
rect 504 2319 506 2341
rect 656 2319 658 2341
rect 816 2319 818 2341
rect 968 2319 970 2341
rect 1120 2319 1122 2341
rect 1264 2319 1266 2341
rect 1416 2319 1418 2341
rect 1568 2319 1570 2341
rect 2032 2319 2034 2346
rect 2072 2341 2074 2369
rect 2112 2360 2114 2369
rect 2328 2360 2330 2369
rect 2560 2360 2562 2369
rect 2784 2360 2786 2369
rect 3000 2360 3002 2369
rect 3192 2360 3194 2369
rect 3376 2360 3378 2369
rect 3544 2360 3546 2369
rect 3712 2360 3714 2369
rect 3888 2360 3890 2369
rect 2110 2359 2116 2360
rect 2110 2355 2111 2359
rect 2115 2355 2116 2359
rect 2110 2354 2116 2355
rect 2326 2359 2332 2360
rect 2326 2355 2327 2359
rect 2331 2355 2332 2359
rect 2326 2354 2332 2355
rect 2558 2359 2564 2360
rect 2558 2355 2559 2359
rect 2563 2355 2564 2359
rect 2558 2354 2564 2355
rect 2782 2359 2788 2360
rect 2782 2355 2783 2359
rect 2787 2355 2788 2359
rect 2782 2354 2788 2355
rect 2998 2359 3004 2360
rect 2998 2355 2999 2359
rect 3003 2355 3004 2359
rect 2998 2354 3004 2355
rect 3190 2359 3196 2360
rect 3190 2355 3191 2359
rect 3195 2355 3196 2359
rect 3190 2354 3196 2355
rect 3374 2359 3380 2360
rect 3374 2355 3375 2359
rect 3379 2355 3380 2359
rect 3374 2354 3380 2355
rect 3542 2359 3548 2360
rect 3542 2355 3543 2359
rect 3547 2355 3548 2359
rect 3542 2354 3548 2355
rect 3710 2359 3716 2360
rect 3710 2355 3711 2359
rect 3715 2355 3716 2359
rect 3710 2354 3716 2355
rect 3886 2359 3892 2360
rect 3886 2355 3887 2359
rect 3891 2355 3892 2359
rect 3886 2354 3892 2355
rect 3992 2341 3994 2369
rect 2070 2340 2076 2341
rect 2070 2336 2071 2340
rect 2075 2336 2076 2340
rect 2070 2335 2076 2336
rect 3990 2340 3996 2341
rect 3990 2336 3991 2340
rect 3995 2336 3996 2340
rect 3990 2335 3996 2336
rect 2070 2323 2076 2324
rect 2070 2319 2071 2323
rect 2075 2319 2076 2323
rect 3990 2323 3996 2324
rect 3990 2319 3991 2323
rect 3995 2319 3996 2323
rect 111 2318 115 2319
rect 111 2313 115 2314
rect 207 2318 211 2319
rect 207 2313 211 2314
rect 255 2318 259 2319
rect 255 2313 259 2314
rect 351 2318 355 2319
rect 351 2313 355 2314
rect 359 2318 363 2319
rect 359 2313 363 2314
rect 471 2318 475 2319
rect 471 2313 475 2314
rect 503 2318 507 2319
rect 503 2313 507 2314
rect 583 2318 587 2319
rect 583 2313 587 2314
rect 655 2318 659 2319
rect 655 2313 659 2314
rect 695 2318 699 2319
rect 695 2313 699 2314
rect 807 2318 811 2319
rect 807 2313 811 2314
rect 815 2318 819 2319
rect 815 2313 819 2314
rect 919 2318 923 2319
rect 919 2313 923 2314
rect 967 2318 971 2319
rect 967 2313 971 2314
rect 1031 2318 1035 2319
rect 1031 2313 1035 2314
rect 1119 2318 1123 2319
rect 1119 2313 1123 2314
rect 1151 2318 1155 2319
rect 1151 2313 1155 2314
rect 1263 2318 1267 2319
rect 1263 2313 1267 2314
rect 1271 2318 1275 2319
rect 1271 2313 1275 2314
rect 1415 2318 1419 2319
rect 1415 2313 1419 2314
rect 1567 2318 1571 2319
rect 1567 2313 1571 2314
rect 2031 2318 2035 2319
rect 2070 2318 2076 2319
rect 2110 2318 2116 2319
rect 2031 2313 2035 2314
rect 112 2298 114 2313
rect 256 2303 258 2313
rect 360 2303 362 2313
rect 472 2303 474 2313
rect 584 2303 586 2313
rect 696 2303 698 2313
rect 808 2303 810 2313
rect 920 2303 922 2313
rect 1032 2303 1034 2313
rect 1152 2303 1154 2313
rect 1272 2303 1274 2313
rect 254 2302 260 2303
rect 254 2298 255 2302
rect 259 2298 260 2302
rect 110 2297 116 2298
rect 254 2297 260 2298
rect 358 2302 364 2303
rect 358 2298 359 2302
rect 363 2298 364 2302
rect 358 2297 364 2298
rect 470 2302 476 2303
rect 470 2298 471 2302
rect 475 2298 476 2302
rect 470 2297 476 2298
rect 582 2302 588 2303
rect 582 2298 583 2302
rect 587 2298 588 2302
rect 582 2297 588 2298
rect 694 2302 700 2303
rect 694 2298 695 2302
rect 699 2298 700 2302
rect 694 2297 700 2298
rect 806 2302 812 2303
rect 806 2298 807 2302
rect 811 2298 812 2302
rect 806 2297 812 2298
rect 918 2302 924 2303
rect 918 2298 919 2302
rect 923 2298 924 2302
rect 918 2297 924 2298
rect 1030 2302 1036 2303
rect 1030 2298 1031 2302
rect 1035 2298 1036 2302
rect 1030 2297 1036 2298
rect 1150 2302 1156 2303
rect 1150 2298 1151 2302
rect 1155 2298 1156 2302
rect 1150 2297 1156 2298
rect 1270 2302 1276 2303
rect 1270 2298 1271 2302
rect 1275 2298 1276 2302
rect 2032 2298 2034 2313
rect 2072 2303 2074 2318
rect 2110 2314 2111 2318
rect 2115 2314 2116 2318
rect 2110 2313 2116 2314
rect 2326 2318 2332 2319
rect 2326 2314 2327 2318
rect 2331 2314 2332 2318
rect 2326 2313 2332 2314
rect 2558 2318 2564 2319
rect 2558 2314 2559 2318
rect 2563 2314 2564 2318
rect 2558 2313 2564 2314
rect 2782 2318 2788 2319
rect 2782 2314 2783 2318
rect 2787 2314 2788 2318
rect 2782 2313 2788 2314
rect 2998 2318 3004 2319
rect 2998 2314 2999 2318
rect 3003 2314 3004 2318
rect 2998 2313 3004 2314
rect 3190 2318 3196 2319
rect 3190 2314 3191 2318
rect 3195 2314 3196 2318
rect 3190 2313 3196 2314
rect 3374 2318 3380 2319
rect 3374 2314 3375 2318
rect 3379 2314 3380 2318
rect 3374 2313 3380 2314
rect 3542 2318 3548 2319
rect 3542 2314 3543 2318
rect 3547 2314 3548 2318
rect 3542 2313 3548 2314
rect 3710 2318 3716 2319
rect 3710 2314 3711 2318
rect 3715 2314 3716 2318
rect 3710 2313 3716 2314
rect 3886 2318 3892 2319
rect 3990 2318 3996 2319
rect 3886 2314 3887 2318
rect 3891 2314 3892 2318
rect 3886 2313 3892 2314
rect 2112 2303 2114 2313
rect 2328 2303 2330 2313
rect 2560 2303 2562 2313
rect 2784 2303 2786 2313
rect 3000 2303 3002 2313
rect 3192 2303 3194 2313
rect 3376 2303 3378 2313
rect 3544 2303 3546 2313
rect 3712 2303 3714 2313
rect 3888 2303 3890 2313
rect 3992 2303 3994 2318
rect 2071 2302 2075 2303
rect 1270 2297 1276 2298
rect 2030 2297 2036 2298
rect 2071 2297 2075 2298
rect 2111 2302 2115 2303
rect 2111 2297 2115 2298
rect 2295 2302 2299 2303
rect 2295 2297 2299 2298
rect 2327 2302 2331 2303
rect 2327 2297 2331 2298
rect 2527 2302 2531 2303
rect 2527 2297 2531 2298
rect 2559 2302 2563 2303
rect 2559 2297 2563 2298
rect 2775 2302 2779 2303
rect 2775 2297 2779 2298
rect 2783 2302 2787 2303
rect 2783 2297 2787 2298
rect 2999 2302 3003 2303
rect 2999 2297 3003 2298
rect 3039 2302 3043 2303
rect 3039 2297 3043 2298
rect 3191 2302 3195 2303
rect 3191 2297 3195 2298
rect 3319 2302 3323 2303
rect 3319 2297 3323 2298
rect 3375 2302 3379 2303
rect 3375 2297 3379 2298
rect 3543 2302 3547 2303
rect 3543 2297 3547 2298
rect 3607 2302 3611 2303
rect 3607 2297 3611 2298
rect 3711 2302 3715 2303
rect 3711 2297 3715 2298
rect 3887 2302 3891 2303
rect 3887 2297 3891 2298
rect 3895 2302 3899 2303
rect 3895 2297 3899 2298
rect 3991 2302 3995 2303
rect 3991 2297 3995 2298
rect 110 2293 111 2297
rect 115 2293 116 2297
rect 110 2292 116 2293
rect 2030 2293 2031 2297
rect 2035 2293 2036 2297
rect 2030 2292 2036 2293
rect 2072 2282 2074 2297
rect 2112 2287 2114 2297
rect 2296 2287 2298 2297
rect 2528 2287 2530 2297
rect 2776 2287 2778 2297
rect 3040 2287 3042 2297
rect 3320 2287 3322 2297
rect 3608 2287 3610 2297
rect 3896 2287 3898 2297
rect 2110 2286 2116 2287
rect 2110 2282 2111 2286
rect 2115 2282 2116 2286
rect 2070 2281 2076 2282
rect 2110 2281 2116 2282
rect 2294 2286 2300 2287
rect 2294 2282 2295 2286
rect 2299 2282 2300 2286
rect 2294 2281 2300 2282
rect 2526 2286 2532 2287
rect 2526 2282 2527 2286
rect 2531 2282 2532 2286
rect 2526 2281 2532 2282
rect 2774 2286 2780 2287
rect 2774 2282 2775 2286
rect 2779 2282 2780 2286
rect 2774 2281 2780 2282
rect 3038 2286 3044 2287
rect 3038 2282 3039 2286
rect 3043 2282 3044 2286
rect 3038 2281 3044 2282
rect 3318 2286 3324 2287
rect 3318 2282 3319 2286
rect 3323 2282 3324 2286
rect 3318 2281 3324 2282
rect 3606 2286 3612 2287
rect 3606 2282 3607 2286
rect 3611 2282 3612 2286
rect 3606 2281 3612 2282
rect 3894 2286 3900 2287
rect 3894 2282 3895 2286
rect 3899 2282 3900 2286
rect 3992 2282 3994 2297
rect 3894 2281 3900 2282
rect 3990 2281 3996 2282
rect 110 2280 116 2281
rect 110 2276 111 2280
rect 115 2276 116 2280
rect 110 2275 116 2276
rect 2030 2280 2036 2281
rect 2030 2276 2031 2280
rect 2035 2276 2036 2280
rect 2070 2277 2071 2281
rect 2075 2277 2076 2281
rect 2070 2276 2076 2277
rect 3990 2277 3991 2281
rect 3995 2277 3996 2281
rect 3990 2276 3996 2277
rect 2030 2275 2036 2276
rect 112 2235 114 2275
rect 254 2261 260 2262
rect 254 2257 255 2261
rect 259 2257 260 2261
rect 254 2256 260 2257
rect 358 2261 364 2262
rect 358 2257 359 2261
rect 363 2257 364 2261
rect 358 2256 364 2257
rect 470 2261 476 2262
rect 470 2257 471 2261
rect 475 2257 476 2261
rect 470 2256 476 2257
rect 582 2261 588 2262
rect 582 2257 583 2261
rect 587 2257 588 2261
rect 582 2256 588 2257
rect 694 2261 700 2262
rect 694 2257 695 2261
rect 699 2257 700 2261
rect 694 2256 700 2257
rect 806 2261 812 2262
rect 806 2257 807 2261
rect 811 2257 812 2261
rect 806 2256 812 2257
rect 918 2261 924 2262
rect 918 2257 919 2261
rect 923 2257 924 2261
rect 918 2256 924 2257
rect 1030 2261 1036 2262
rect 1030 2257 1031 2261
rect 1035 2257 1036 2261
rect 1030 2256 1036 2257
rect 1150 2261 1156 2262
rect 1150 2257 1151 2261
rect 1155 2257 1156 2261
rect 1150 2256 1156 2257
rect 1270 2261 1276 2262
rect 1270 2257 1271 2261
rect 1275 2257 1276 2261
rect 1270 2256 1276 2257
rect 256 2235 258 2256
rect 360 2235 362 2256
rect 472 2235 474 2256
rect 584 2235 586 2256
rect 696 2235 698 2256
rect 808 2235 810 2256
rect 920 2235 922 2256
rect 1032 2235 1034 2256
rect 1152 2235 1154 2256
rect 1272 2235 1274 2256
rect 2032 2235 2034 2275
rect 2070 2264 2076 2265
rect 2070 2260 2071 2264
rect 2075 2260 2076 2264
rect 2070 2259 2076 2260
rect 3990 2264 3996 2265
rect 3990 2260 3991 2264
rect 3995 2260 3996 2264
rect 3990 2259 3996 2260
rect 111 2234 115 2235
rect 111 2229 115 2230
rect 183 2234 187 2235
rect 183 2229 187 2230
rect 255 2234 259 2235
rect 255 2229 259 2230
rect 343 2234 347 2235
rect 343 2229 347 2230
rect 359 2234 363 2235
rect 359 2229 363 2230
rect 471 2234 475 2235
rect 471 2229 475 2230
rect 495 2234 499 2235
rect 495 2229 499 2230
rect 583 2234 587 2235
rect 583 2229 587 2230
rect 647 2234 651 2235
rect 647 2229 651 2230
rect 695 2234 699 2235
rect 695 2229 699 2230
rect 791 2234 795 2235
rect 791 2229 795 2230
rect 807 2234 811 2235
rect 807 2229 811 2230
rect 919 2234 923 2235
rect 919 2229 923 2230
rect 935 2234 939 2235
rect 935 2229 939 2230
rect 1031 2234 1035 2235
rect 1031 2229 1035 2230
rect 1071 2234 1075 2235
rect 1071 2229 1075 2230
rect 1151 2234 1155 2235
rect 1151 2229 1155 2230
rect 1199 2234 1203 2235
rect 1199 2229 1203 2230
rect 1271 2234 1275 2235
rect 1271 2229 1275 2230
rect 1335 2234 1339 2235
rect 1335 2229 1339 2230
rect 1471 2234 1475 2235
rect 1471 2229 1475 2230
rect 2031 2234 2035 2235
rect 2031 2229 2035 2230
rect 112 2201 114 2229
rect 184 2220 186 2229
rect 344 2220 346 2229
rect 496 2220 498 2229
rect 648 2220 650 2229
rect 792 2220 794 2229
rect 936 2220 938 2229
rect 1072 2220 1074 2229
rect 1200 2220 1202 2229
rect 1336 2220 1338 2229
rect 1472 2220 1474 2229
rect 182 2219 188 2220
rect 182 2215 183 2219
rect 187 2215 188 2219
rect 182 2214 188 2215
rect 342 2219 348 2220
rect 342 2215 343 2219
rect 347 2215 348 2219
rect 342 2214 348 2215
rect 494 2219 500 2220
rect 494 2215 495 2219
rect 499 2215 500 2219
rect 494 2214 500 2215
rect 646 2219 652 2220
rect 646 2215 647 2219
rect 651 2215 652 2219
rect 646 2214 652 2215
rect 790 2219 796 2220
rect 790 2215 791 2219
rect 795 2215 796 2219
rect 790 2214 796 2215
rect 934 2219 940 2220
rect 934 2215 935 2219
rect 939 2215 940 2219
rect 934 2214 940 2215
rect 1070 2219 1076 2220
rect 1070 2215 1071 2219
rect 1075 2215 1076 2219
rect 1070 2214 1076 2215
rect 1198 2219 1204 2220
rect 1198 2215 1199 2219
rect 1203 2215 1204 2219
rect 1198 2214 1204 2215
rect 1334 2219 1340 2220
rect 1334 2215 1335 2219
rect 1339 2215 1340 2219
rect 1334 2214 1340 2215
rect 1470 2219 1476 2220
rect 1470 2215 1471 2219
rect 1475 2215 1476 2219
rect 1470 2214 1476 2215
rect 2032 2201 2034 2229
rect 2072 2223 2074 2259
rect 2110 2245 2116 2246
rect 2110 2241 2111 2245
rect 2115 2241 2116 2245
rect 2110 2240 2116 2241
rect 2294 2245 2300 2246
rect 2294 2241 2295 2245
rect 2299 2241 2300 2245
rect 2294 2240 2300 2241
rect 2526 2245 2532 2246
rect 2526 2241 2527 2245
rect 2531 2241 2532 2245
rect 2526 2240 2532 2241
rect 2774 2245 2780 2246
rect 2774 2241 2775 2245
rect 2779 2241 2780 2245
rect 2774 2240 2780 2241
rect 3038 2245 3044 2246
rect 3038 2241 3039 2245
rect 3043 2241 3044 2245
rect 3038 2240 3044 2241
rect 3318 2245 3324 2246
rect 3318 2241 3319 2245
rect 3323 2241 3324 2245
rect 3318 2240 3324 2241
rect 3606 2245 3612 2246
rect 3606 2241 3607 2245
rect 3611 2241 3612 2245
rect 3606 2240 3612 2241
rect 3894 2245 3900 2246
rect 3894 2241 3895 2245
rect 3899 2241 3900 2245
rect 3894 2240 3900 2241
rect 2112 2223 2114 2240
rect 2296 2223 2298 2240
rect 2528 2223 2530 2240
rect 2776 2223 2778 2240
rect 3040 2223 3042 2240
rect 3320 2223 3322 2240
rect 3608 2223 3610 2240
rect 3896 2223 3898 2240
rect 3992 2223 3994 2259
rect 2071 2222 2075 2223
rect 2071 2217 2075 2218
rect 2111 2222 2115 2223
rect 2111 2217 2115 2218
rect 2279 2222 2283 2223
rect 2279 2217 2283 2218
rect 2295 2222 2299 2223
rect 2295 2217 2299 2218
rect 2439 2222 2443 2223
rect 2439 2217 2443 2218
rect 2527 2222 2531 2223
rect 2527 2217 2531 2218
rect 2623 2222 2627 2223
rect 2623 2217 2627 2218
rect 2775 2222 2779 2223
rect 2775 2217 2779 2218
rect 2839 2222 2843 2223
rect 2839 2217 2843 2218
rect 3039 2222 3043 2223
rect 3039 2217 3043 2218
rect 3079 2222 3083 2223
rect 3079 2217 3083 2218
rect 3319 2222 3323 2223
rect 3319 2217 3323 2218
rect 3343 2222 3347 2223
rect 3343 2217 3347 2218
rect 3607 2222 3611 2223
rect 3607 2217 3611 2218
rect 3623 2222 3627 2223
rect 3623 2217 3627 2218
rect 3895 2222 3899 2223
rect 3895 2217 3899 2218
rect 3991 2222 3995 2223
rect 3991 2217 3995 2218
rect 110 2200 116 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 2030 2200 2036 2201
rect 2030 2196 2031 2200
rect 2035 2196 2036 2200
rect 2030 2195 2036 2196
rect 2072 2189 2074 2217
rect 2280 2208 2282 2217
rect 2440 2208 2442 2217
rect 2624 2208 2626 2217
rect 2840 2208 2842 2217
rect 3080 2208 3082 2217
rect 3344 2208 3346 2217
rect 3624 2208 3626 2217
rect 3896 2208 3898 2217
rect 2278 2207 2284 2208
rect 2278 2203 2279 2207
rect 2283 2203 2284 2207
rect 2278 2202 2284 2203
rect 2438 2207 2444 2208
rect 2438 2203 2439 2207
rect 2443 2203 2444 2207
rect 2438 2202 2444 2203
rect 2622 2207 2628 2208
rect 2622 2203 2623 2207
rect 2627 2203 2628 2207
rect 2622 2202 2628 2203
rect 2838 2207 2844 2208
rect 2838 2203 2839 2207
rect 2843 2203 2844 2207
rect 2838 2202 2844 2203
rect 3078 2207 3084 2208
rect 3078 2203 3079 2207
rect 3083 2203 3084 2207
rect 3078 2202 3084 2203
rect 3342 2207 3348 2208
rect 3342 2203 3343 2207
rect 3347 2203 3348 2207
rect 3342 2202 3348 2203
rect 3622 2207 3628 2208
rect 3622 2203 3623 2207
rect 3627 2203 3628 2207
rect 3622 2202 3628 2203
rect 3894 2207 3900 2208
rect 3894 2203 3895 2207
rect 3899 2203 3900 2207
rect 3894 2202 3900 2203
rect 3992 2189 3994 2217
rect 2070 2188 2076 2189
rect 2070 2184 2071 2188
rect 2075 2184 2076 2188
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 2030 2183 2036 2184
rect 2070 2183 2076 2184
rect 3990 2188 3996 2189
rect 3990 2184 3991 2188
rect 3995 2184 3996 2188
rect 3990 2183 3996 2184
rect 2030 2179 2031 2183
rect 2035 2179 2036 2183
rect 110 2178 116 2179
rect 182 2178 188 2179
rect 112 2147 114 2178
rect 182 2174 183 2178
rect 187 2174 188 2178
rect 182 2173 188 2174
rect 342 2178 348 2179
rect 342 2174 343 2178
rect 347 2174 348 2178
rect 342 2173 348 2174
rect 494 2178 500 2179
rect 494 2174 495 2178
rect 499 2174 500 2178
rect 494 2173 500 2174
rect 646 2178 652 2179
rect 646 2174 647 2178
rect 651 2174 652 2178
rect 646 2173 652 2174
rect 790 2178 796 2179
rect 790 2174 791 2178
rect 795 2174 796 2178
rect 790 2173 796 2174
rect 934 2178 940 2179
rect 934 2174 935 2178
rect 939 2174 940 2178
rect 934 2173 940 2174
rect 1070 2178 1076 2179
rect 1070 2174 1071 2178
rect 1075 2174 1076 2178
rect 1070 2173 1076 2174
rect 1198 2178 1204 2179
rect 1198 2174 1199 2178
rect 1203 2174 1204 2178
rect 1198 2173 1204 2174
rect 1334 2178 1340 2179
rect 1334 2174 1335 2178
rect 1339 2174 1340 2178
rect 1334 2173 1340 2174
rect 1470 2178 1476 2179
rect 2030 2178 2036 2179
rect 1470 2174 1471 2178
rect 1475 2174 1476 2178
rect 1470 2173 1476 2174
rect 184 2147 186 2173
rect 344 2147 346 2173
rect 496 2147 498 2173
rect 648 2147 650 2173
rect 792 2147 794 2173
rect 936 2147 938 2173
rect 1072 2147 1074 2173
rect 1200 2147 1202 2173
rect 1336 2147 1338 2173
rect 1472 2147 1474 2173
rect 2032 2147 2034 2178
rect 2070 2171 2076 2172
rect 2070 2167 2071 2171
rect 2075 2167 2076 2171
rect 3990 2171 3996 2172
rect 3990 2167 3991 2171
rect 3995 2167 3996 2171
rect 2070 2166 2076 2167
rect 2278 2166 2284 2167
rect 2072 2151 2074 2166
rect 2278 2162 2279 2166
rect 2283 2162 2284 2166
rect 2278 2161 2284 2162
rect 2438 2166 2444 2167
rect 2438 2162 2439 2166
rect 2443 2162 2444 2166
rect 2438 2161 2444 2162
rect 2622 2166 2628 2167
rect 2622 2162 2623 2166
rect 2627 2162 2628 2166
rect 2622 2161 2628 2162
rect 2838 2166 2844 2167
rect 2838 2162 2839 2166
rect 2843 2162 2844 2166
rect 2838 2161 2844 2162
rect 3078 2166 3084 2167
rect 3078 2162 3079 2166
rect 3083 2162 3084 2166
rect 3078 2161 3084 2162
rect 3342 2166 3348 2167
rect 3342 2162 3343 2166
rect 3347 2162 3348 2166
rect 3342 2161 3348 2162
rect 3622 2166 3628 2167
rect 3622 2162 3623 2166
rect 3627 2162 3628 2166
rect 3622 2161 3628 2162
rect 3894 2166 3900 2167
rect 3990 2166 3996 2167
rect 3894 2162 3895 2166
rect 3899 2162 3900 2166
rect 3894 2161 3900 2162
rect 2280 2151 2282 2161
rect 2440 2151 2442 2161
rect 2624 2151 2626 2161
rect 2840 2151 2842 2161
rect 3080 2151 3082 2161
rect 3344 2151 3346 2161
rect 3624 2151 3626 2161
rect 3896 2151 3898 2161
rect 3992 2151 3994 2166
rect 2071 2150 2075 2151
rect 111 2146 115 2147
rect 111 2141 115 2142
rect 151 2146 155 2147
rect 151 2141 155 2142
rect 183 2146 187 2147
rect 183 2141 187 2142
rect 327 2146 331 2147
rect 327 2141 331 2142
rect 343 2146 347 2147
rect 343 2141 347 2142
rect 495 2146 499 2147
rect 495 2141 499 2142
rect 535 2146 539 2147
rect 535 2141 539 2142
rect 647 2146 651 2147
rect 647 2141 651 2142
rect 735 2146 739 2147
rect 735 2141 739 2142
rect 791 2146 795 2147
rect 791 2141 795 2142
rect 927 2146 931 2147
rect 927 2141 931 2142
rect 935 2146 939 2147
rect 935 2141 939 2142
rect 1071 2146 1075 2147
rect 1071 2141 1075 2142
rect 1111 2146 1115 2147
rect 1111 2141 1115 2142
rect 1199 2146 1203 2147
rect 1199 2141 1203 2142
rect 1279 2146 1283 2147
rect 1279 2141 1283 2142
rect 1335 2146 1339 2147
rect 1335 2141 1339 2142
rect 1447 2146 1451 2147
rect 1447 2141 1451 2142
rect 1471 2146 1475 2147
rect 1471 2141 1475 2142
rect 1615 2146 1619 2147
rect 1615 2141 1619 2142
rect 1783 2146 1787 2147
rect 1783 2141 1787 2142
rect 2031 2146 2035 2147
rect 2071 2145 2075 2146
rect 2279 2150 2283 2151
rect 2279 2145 2283 2146
rect 2391 2150 2395 2151
rect 2391 2145 2395 2146
rect 2439 2150 2443 2151
rect 2439 2145 2443 2146
rect 2495 2150 2499 2151
rect 2495 2145 2499 2146
rect 2599 2150 2603 2151
rect 2599 2145 2603 2146
rect 2623 2150 2627 2151
rect 2623 2145 2627 2146
rect 2703 2150 2707 2151
rect 2703 2145 2707 2146
rect 2807 2150 2811 2151
rect 2807 2145 2811 2146
rect 2839 2150 2843 2151
rect 2839 2145 2843 2146
rect 2911 2150 2915 2151
rect 2911 2145 2915 2146
rect 3031 2150 3035 2151
rect 3031 2145 3035 2146
rect 3079 2150 3083 2151
rect 3079 2145 3083 2146
rect 3175 2150 3179 2151
rect 3175 2145 3179 2146
rect 3343 2150 3347 2151
rect 3343 2145 3347 2146
rect 3527 2150 3531 2151
rect 3527 2145 3531 2146
rect 3623 2150 3627 2151
rect 3623 2145 3627 2146
rect 3719 2150 3723 2151
rect 3719 2145 3723 2146
rect 3895 2150 3899 2151
rect 3895 2145 3899 2146
rect 3991 2150 3995 2151
rect 3991 2145 3995 2146
rect 2031 2141 2035 2142
rect 112 2126 114 2141
rect 152 2131 154 2141
rect 328 2131 330 2141
rect 536 2131 538 2141
rect 736 2131 738 2141
rect 928 2131 930 2141
rect 1112 2131 1114 2141
rect 1280 2131 1282 2141
rect 1448 2131 1450 2141
rect 1616 2131 1618 2141
rect 1784 2131 1786 2141
rect 150 2130 156 2131
rect 150 2126 151 2130
rect 155 2126 156 2130
rect 110 2125 116 2126
rect 150 2125 156 2126
rect 326 2130 332 2131
rect 326 2126 327 2130
rect 331 2126 332 2130
rect 326 2125 332 2126
rect 534 2130 540 2131
rect 534 2126 535 2130
rect 539 2126 540 2130
rect 534 2125 540 2126
rect 734 2130 740 2131
rect 734 2126 735 2130
rect 739 2126 740 2130
rect 734 2125 740 2126
rect 926 2130 932 2131
rect 926 2126 927 2130
rect 931 2126 932 2130
rect 926 2125 932 2126
rect 1110 2130 1116 2131
rect 1110 2126 1111 2130
rect 1115 2126 1116 2130
rect 1110 2125 1116 2126
rect 1278 2130 1284 2131
rect 1278 2126 1279 2130
rect 1283 2126 1284 2130
rect 1278 2125 1284 2126
rect 1446 2130 1452 2131
rect 1446 2126 1447 2130
rect 1451 2126 1452 2130
rect 1446 2125 1452 2126
rect 1614 2130 1620 2131
rect 1614 2126 1615 2130
rect 1619 2126 1620 2130
rect 1614 2125 1620 2126
rect 1782 2130 1788 2131
rect 1782 2126 1783 2130
rect 1787 2126 1788 2130
rect 2032 2126 2034 2141
rect 2072 2130 2074 2145
rect 2392 2135 2394 2145
rect 2496 2135 2498 2145
rect 2600 2135 2602 2145
rect 2704 2135 2706 2145
rect 2808 2135 2810 2145
rect 2912 2135 2914 2145
rect 3032 2135 3034 2145
rect 3176 2135 3178 2145
rect 3344 2135 3346 2145
rect 3528 2135 3530 2145
rect 3720 2135 3722 2145
rect 3896 2135 3898 2145
rect 2390 2134 2396 2135
rect 2390 2130 2391 2134
rect 2395 2130 2396 2134
rect 2070 2129 2076 2130
rect 2390 2129 2396 2130
rect 2494 2134 2500 2135
rect 2494 2130 2495 2134
rect 2499 2130 2500 2134
rect 2494 2129 2500 2130
rect 2598 2134 2604 2135
rect 2598 2130 2599 2134
rect 2603 2130 2604 2134
rect 2598 2129 2604 2130
rect 2702 2134 2708 2135
rect 2702 2130 2703 2134
rect 2707 2130 2708 2134
rect 2702 2129 2708 2130
rect 2806 2134 2812 2135
rect 2806 2130 2807 2134
rect 2811 2130 2812 2134
rect 2806 2129 2812 2130
rect 2910 2134 2916 2135
rect 2910 2130 2911 2134
rect 2915 2130 2916 2134
rect 2910 2129 2916 2130
rect 3030 2134 3036 2135
rect 3030 2130 3031 2134
rect 3035 2130 3036 2134
rect 3030 2129 3036 2130
rect 3174 2134 3180 2135
rect 3174 2130 3175 2134
rect 3179 2130 3180 2134
rect 3174 2129 3180 2130
rect 3342 2134 3348 2135
rect 3342 2130 3343 2134
rect 3347 2130 3348 2134
rect 3342 2129 3348 2130
rect 3526 2134 3532 2135
rect 3526 2130 3527 2134
rect 3531 2130 3532 2134
rect 3526 2129 3532 2130
rect 3718 2134 3724 2135
rect 3718 2130 3719 2134
rect 3723 2130 3724 2134
rect 3718 2129 3724 2130
rect 3894 2134 3900 2135
rect 3894 2130 3895 2134
rect 3899 2130 3900 2134
rect 3992 2130 3994 2145
rect 3894 2129 3900 2130
rect 3990 2129 3996 2130
rect 1782 2125 1788 2126
rect 2030 2125 2036 2126
rect 110 2121 111 2125
rect 115 2121 116 2125
rect 110 2120 116 2121
rect 2030 2121 2031 2125
rect 2035 2121 2036 2125
rect 2070 2125 2071 2129
rect 2075 2125 2076 2129
rect 2070 2124 2076 2125
rect 3990 2125 3991 2129
rect 3995 2125 3996 2129
rect 3990 2124 3996 2125
rect 2030 2120 2036 2121
rect 2070 2112 2076 2113
rect 110 2108 116 2109
rect 110 2104 111 2108
rect 115 2104 116 2108
rect 110 2103 116 2104
rect 2030 2108 2036 2109
rect 2030 2104 2031 2108
rect 2035 2104 2036 2108
rect 2070 2108 2071 2112
rect 2075 2108 2076 2112
rect 2070 2107 2076 2108
rect 3990 2112 3996 2113
rect 3990 2108 3991 2112
rect 3995 2108 3996 2112
rect 3990 2107 3996 2108
rect 2030 2103 2036 2104
rect 112 2063 114 2103
rect 150 2089 156 2090
rect 150 2085 151 2089
rect 155 2085 156 2089
rect 150 2084 156 2085
rect 326 2089 332 2090
rect 326 2085 327 2089
rect 331 2085 332 2089
rect 326 2084 332 2085
rect 534 2089 540 2090
rect 534 2085 535 2089
rect 539 2085 540 2089
rect 534 2084 540 2085
rect 734 2089 740 2090
rect 734 2085 735 2089
rect 739 2085 740 2089
rect 734 2084 740 2085
rect 926 2089 932 2090
rect 926 2085 927 2089
rect 931 2085 932 2089
rect 926 2084 932 2085
rect 1110 2089 1116 2090
rect 1110 2085 1111 2089
rect 1115 2085 1116 2089
rect 1110 2084 1116 2085
rect 1278 2089 1284 2090
rect 1278 2085 1279 2089
rect 1283 2085 1284 2089
rect 1278 2084 1284 2085
rect 1446 2089 1452 2090
rect 1446 2085 1447 2089
rect 1451 2085 1452 2089
rect 1446 2084 1452 2085
rect 1614 2089 1620 2090
rect 1614 2085 1615 2089
rect 1619 2085 1620 2089
rect 1614 2084 1620 2085
rect 1782 2089 1788 2090
rect 1782 2085 1783 2089
rect 1787 2085 1788 2089
rect 1782 2084 1788 2085
rect 152 2063 154 2084
rect 328 2063 330 2084
rect 536 2063 538 2084
rect 736 2063 738 2084
rect 928 2063 930 2084
rect 1112 2063 1114 2084
rect 1280 2063 1282 2084
rect 1448 2063 1450 2084
rect 1616 2063 1618 2084
rect 1784 2063 1786 2084
rect 2032 2063 2034 2103
rect 2072 2075 2074 2107
rect 2390 2093 2396 2094
rect 2390 2089 2391 2093
rect 2395 2089 2396 2093
rect 2390 2088 2396 2089
rect 2494 2093 2500 2094
rect 2494 2089 2495 2093
rect 2499 2089 2500 2093
rect 2494 2088 2500 2089
rect 2598 2093 2604 2094
rect 2598 2089 2599 2093
rect 2603 2089 2604 2093
rect 2598 2088 2604 2089
rect 2702 2093 2708 2094
rect 2702 2089 2703 2093
rect 2707 2089 2708 2093
rect 2702 2088 2708 2089
rect 2806 2093 2812 2094
rect 2806 2089 2807 2093
rect 2811 2089 2812 2093
rect 2806 2088 2812 2089
rect 2910 2093 2916 2094
rect 2910 2089 2911 2093
rect 2915 2089 2916 2093
rect 2910 2088 2916 2089
rect 3030 2093 3036 2094
rect 3030 2089 3031 2093
rect 3035 2089 3036 2093
rect 3030 2088 3036 2089
rect 3174 2093 3180 2094
rect 3174 2089 3175 2093
rect 3179 2089 3180 2093
rect 3174 2088 3180 2089
rect 3342 2093 3348 2094
rect 3342 2089 3343 2093
rect 3347 2089 3348 2093
rect 3342 2088 3348 2089
rect 3526 2093 3532 2094
rect 3526 2089 3527 2093
rect 3531 2089 3532 2093
rect 3526 2088 3532 2089
rect 3718 2093 3724 2094
rect 3718 2089 3719 2093
rect 3723 2089 3724 2093
rect 3718 2088 3724 2089
rect 3894 2093 3900 2094
rect 3894 2089 3895 2093
rect 3899 2089 3900 2093
rect 3894 2088 3900 2089
rect 2392 2075 2394 2088
rect 2496 2075 2498 2088
rect 2600 2075 2602 2088
rect 2704 2075 2706 2088
rect 2808 2075 2810 2088
rect 2912 2075 2914 2088
rect 3032 2075 3034 2088
rect 3176 2075 3178 2088
rect 3344 2075 3346 2088
rect 3528 2075 3530 2088
rect 3720 2075 3722 2088
rect 3896 2075 3898 2088
rect 3992 2075 3994 2107
rect 2071 2074 2075 2075
rect 2071 2069 2075 2070
rect 2391 2074 2395 2075
rect 2391 2069 2395 2070
rect 2487 2074 2491 2075
rect 2487 2069 2491 2070
rect 2495 2074 2499 2075
rect 2495 2069 2499 2070
rect 2591 2074 2595 2075
rect 2591 2069 2595 2070
rect 2599 2074 2603 2075
rect 2599 2069 2603 2070
rect 2695 2074 2699 2075
rect 2695 2069 2699 2070
rect 2703 2074 2707 2075
rect 2703 2069 2707 2070
rect 2807 2074 2811 2075
rect 2807 2069 2811 2070
rect 2911 2074 2915 2075
rect 2911 2069 2915 2070
rect 2935 2074 2939 2075
rect 2935 2069 2939 2070
rect 3031 2074 3035 2075
rect 3031 2069 3035 2070
rect 3095 2074 3099 2075
rect 3095 2069 3099 2070
rect 3175 2074 3179 2075
rect 3175 2069 3179 2070
rect 3279 2074 3283 2075
rect 3279 2069 3283 2070
rect 3343 2074 3347 2075
rect 3343 2069 3347 2070
rect 3479 2074 3483 2075
rect 3479 2069 3483 2070
rect 3527 2074 3531 2075
rect 3527 2069 3531 2070
rect 3695 2074 3699 2075
rect 3695 2069 3699 2070
rect 3719 2074 3723 2075
rect 3719 2069 3723 2070
rect 3895 2074 3899 2075
rect 3895 2069 3899 2070
rect 3991 2074 3995 2075
rect 3991 2069 3995 2070
rect 111 2062 115 2063
rect 111 2057 115 2058
rect 151 2062 155 2063
rect 151 2057 155 2058
rect 327 2062 331 2063
rect 327 2057 331 2058
rect 383 2062 387 2063
rect 383 2057 387 2058
rect 535 2062 539 2063
rect 535 2057 539 2058
rect 631 2062 635 2063
rect 631 2057 635 2058
rect 735 2062 739 2063
rect 735 2057 739 2058
rect 863 2062 867 2063
rect 863 2057 867 2058
rect 927 2062 931 2063
rect 927 2057 931 2058
rect 1071 2062 1075 2063
rect 1071 2057 1075 2058
rect 1111 2062 1115 2063
rect 1111 2057 1115 2058
rect 1263 2062 1267 2063
rect 1263 2057 1267 2058
rect 1279 2062 1283 2063
rect 1279 2057 1283 2058
rect 1447 2062 1451 2063
rect 1447 2057 1451 2058
rect 1615 2062 1619 2063
rect 1615 2057 1619 2058
rect 1783 2062 1787 2063
rect 1783 2057 1787 2058
rect 1935 2062 1939 2063
rect 1935 2057 1939 2058
rect 2031 2062 2035 2063
rect 2031 2057 2035 2058
rect 112 2029 114 2057
rect 152 2048 154 2057
rect 384 2048 386 2057
rect 632 2048 634 2057
rect 864 2048 866 2057
rect 1072 2048 1074 2057
rect 1264 2048 1266 2057
rect 1448 2048 1450 2057
rect 1616 2048 1618 2057
rect 1784 2048 1786 2057
rect 1936 2048 1938 2057
rect 150 2047 156 2048
rect 150 2043 151 2047
rect 155 2043 156 2047
rect 150 2042 156 2043
rect 382 2047 388 2048
rect 382 2043 383 2047
rect 387 2043 388 2047
rect 382 2042 388 2043
rect 630 2047 636 2048
rect 630 2043 631 2047
rect 635 2043 636 2047
rect 630 2042 636 2043
rect 862 2047 868 2048
rect 862 2043 863 2047
rect 867 2043 868 2047
rect 862 2042 868 2043
rect 1070 2047 1076 2048
rect 1070 2043 1071 2047
rect 1075 2043 1076 2047
rect 1070 2042 1076 2043
rect 1262 2047 1268 2048
rect 1262 2043 1263 2047
rect 1267 2043 1268 2047
rect 1262 2042 1268 2043
rect 1446 2047 1452 2048
rect 1446 2043 1447 2047
rect 1451 2043 1452 2047
rect 1446 2042 1452 2043
rect 1614 2047 1620 2048
rect 1614 2043 1615 2047
rect 1619 2043 1620 2047
rect 1614 2042 1620 2043
rect 1782 2047 1788 2048
rect 1782 2043 1783 2047
rect 1787 2043 1788 2047
rect 1782 2042 1788 2043
rect 1934 2047 1940 2048
rect 1934 2043 1935 2047
rect 1939 2043 1940 2047
rect 1934 2042 1940 2043
rect 2032 2029 2034 2057
rect 2072 2041 2074 2069
rect 2488 2060 2490 2069
rect 2592 2060 2594 2069
rect 2696 2060 2698 2069
rect 2808 2060 2810 2069
rect 2936 2060 2938 2069
rect 3096 2060 3098 2069
rect 3280 2060 3282 2069
rect 3480 2060 3482 2069
rect 3696 2060 3698 2069
rect 3896 2060 3898 2069
rect 2486 2059 2492 2060
rect 2486 2055 2487 2059
rect 2491 2055 2492 2059
rect 2486 2054 2492 2055
rect 2590 2059 2596 2060
rect 2590 2055 2591 2059
rect 2595 2055 2596 2059
rect 2590 2054 2596 2055
rect 2694 2059 2700 2060
rect 2694 2055 2695 2059
rect 2699 2055 2700 2059
rect 2694 2054 2700 2055
rect 2806 2059 2812 2060
rect 2806 2055 2807 2059
rect 2811 2055 2812 2059
rect 2806 2054 2812 2055
rect 2934 2059 2940 2060
rect 2934 2055 2935 2059
rect 2939 2055 2940 2059
rect 2934 2054 2940 2055
rect 3094 2059 3100 2060
rect 3094 2055 3095 2059
rect 3099 2055 3100 2059
rect 3094 2054 3100 2055
rect 3278 2059 3284 2060
rect 3278 2055 3279 2059
rect 3283 2055 3284 2059
rect 3278 2054 3284 2055
rect 3478 2059 3484 2060
rect 3478 2055 3479 2059
rect 3483 2055 3484 2059
rect 3478 2054 3484 2055
rect 3694 2059 3700 2060
rect 3694 2055 3695 2059
rect 3699 2055 3700 2059
rect 3694 2054 3700 2055
rect 3894 2059 3900 2060
rect 3894 2055 3895 2059
rect 3899 2055 3900 2059
rect 3894 2054 3900 2055
rect 3992 2041 3994 2069
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 3990 2040 3996 2041
rect 3990 2036 3991 2040
rect 3995 2036 3996 2040
rect 3990 2035 3996 2036
rect 110 2028 116 2029
rect 110 2024 111 2028
rect 115 2024 116 2028
rect 110 2023 116 2024
rect 2030 2028 2036 2029
rect 2030 2024 2031 2028
rect 2035 2024 2036 2028
rect 2030 2023 2036 2024
rect 2070 2023 2076 2024
rect 2070 2019 2071 2023
rect 2075 2019 2076 2023
rect 3990 2023 3996 2024
rect 3990 2019 3991 2023
rect 3995 2019 3996 2023
rect 2070 2018 2076 2019
rect 2486 2018 2492 2019
rect 110 2011 116 2012
rect 110 2007 111 2011
rect 115 2007 116 2011
rect 2030 2011 2036 2012
rect 2030 2007 2031 2011
rect 2035 2007 2036 2011
rect 110 2006 116 2007
rect 150 2006 156 2007
rect 112 1979 114 2006
rect 150 2002 151 2006
rect 155 2002 156 2006
rect 150 2001 156 2002
rect 382 2006 388 2007
rect 382 2002 383 2006
rect 387 2002 388 2006
rect 382 2001 388 2002
rect 630 2006 636 2007
rect 630 2002 631 2006
rect 635 2002 636 2006
rect 630 2001 636 2002
rect 862 2006 868 2007
rect 862 2002 863 2006
rect 867 2002 868 2006
rect 862 2001 868 2002
rect 1070 2006 1076 2007
rect 1070 2002 1071 2006
rect 1075 2002 1076 2006
rect 1070 2001 1076 2002
rect 1262 2006 1268 2007
rect 1262 2002 1263 2006
rect 1267 2002 1268 2006
rect 1262 2001 1268 2002
rect 1446 2006 1452 2007
rect 1446 2002 1447 2006
rect 1451 2002 1452 2006
rect 1446 2001 1452 2002
rect 1614 2006 1620 2007
rect 1614 2002 1615 2006
rect 1619 2002 1620 2006
rect 1614 2001 1620 2002
rect 1782 2006 1788 2007
rect 1782 2002 1783 2006
rect 1787 2002 1788 2006
rect 1782 2001 1788 2002
rect 1934 2006 1940 2007
rect 2030 2006 2036 2007
rect 1934 2002 1935 2006
rect 1939 2002 1940 2006
rect 1934 2001 1940 2002
rect 152 1979 154 2001
rect 384 1979 386 2001
rect 632 1979 634 2001
rect 864 1979 866 2001
rect 1072 1979 1074 2001
rect 1264 1979 1266 2001
rect 1448 1979 1450 2001
rect 1616 1979 1618 2001
rect 1784 1979 1786 2001
rect 1936 1979 1938 2001
rect 2032 1979 2034 2006
rect 2072 1995 2074 2018
rect 2486 2014 2487 2018
rect 2491 2014 2492 2018
rect 2486 2013 2492 2014
rect 2590 2018 2596 2019
rect 2590 2014 2591 2018
rect 2595 2014 2596 2018
rect 2590 2013 2596 2014
rect 2694 2018 2700 2019
rect 2694 2014 2695 2018
rect 2699 2014 2700 2018
rect 2694 2013 2700 2014
rect 2806 2018 2812 2019
rect 2806 2014 2807 2018
rect 2811 2014 2812 2018
rect 2806 2013 2812 2014
rect 2934 2018 2940 2019
rect 2934 2014 2935 2018
rect 2939 2014 2940 2018
rect 2934 2013 2940 2014
rect 3094 2018 3100 2019
rect 3094 2014 3095 2018
rect 3099 2014 3100 2018
rect 3094 2013 3100 2014
rect 3278 2018 3284 2019
rect 3278 2014 3279 2018
rect 3283 2014 3284 2018
rect 3278 2013 3284 2014
rect 3478 2018 3484 2019
rect 3478 2014 3479 2018
rect 3483 2014 3484 2018
rect 3478 2013 3484 2014
rect 3694 2018 3700 2019
rect 3694 2014 3695 2018
rect 3699 2014 3700 2018
rect 3694 2013 3700 2014
rect 3894 2018 3900 2019
rect 3990 2018 3996 2019
rect 3894 2014 3895 2018
rect 3899 2014 3900 2018
rect 3894 2013 3900 2014
rect 2488 1995 2490 2013
rect 2592 1995 2594 2013
rect 2696 1995 2698 2013
rect 2808 1995 2810 2013
rect 2936 1995 2938 2013
rect 3096 1995 3098 2013
rect 3280 1995 3282 2013
rect 3480 1995 3482 2013
rect 3696 1995 3698 2013
rect 3896 1995 3898 2013
rect 3992 1995 3994 2018
rect 2071 1994 2075 1995
rect 2071 1989 2075 1990
rect 2487 1994 2491 1995
rect 2487 1989 2491 1990
rect 2527 1994 2531 1995
rect 2527 1989 2531 1990
rect 2591 1994 2595 1995
rect 2591 1989 2595 1990
rect 2695 1994 2699 1995
rect 2695 1989 2699 1990
rect 2703 1994 2707 1995
rect 2703 1989 2707 1990
rect 2807 1994 2811 1995
rect 2807 1989 2811 1990
rect 2887 1994 2891 1995
rect 2887 1989 2891 1990
rect 2935 1994 2939 1995
rect 2935 1989 2939 1990
rect 3079 1994 3083 1995
rect 3079 1989 3083 1990
rect 3095 1994 3099 1995
rect 3095 1989 3099 1990
rect 3279 1994 3283 1995
rect 3279 1989 3283 1990
rect 3479 1994 3483 1995
rect 3479 1989 3483 1990
rect 3487 1994 3491 1995
rect 3487 1989 3491 1990
rect 3695 1994 3699 1995
rect 3695 1989 3699 1990
rect 3703 1994 3707 1995
rect 3703 1989 3707 1990
rect 3895 1994 3899 1995
rect 3895 1989 3899 1990
rect 3991 1994 3995 1995
rect 3991 1989 3995 1990
rect 111 1978 115 1979
rect 111 1973 115 1974
rect 151 1978 155 1979
rect 151 1973 155 1974
rect 327 1978 331 1979
rect 327 1973 331 1974
rect 383 1978 387 1979
rect 383 1973 387 1974
rect 535 1978 539 1979
rect 535 1973 539 1974
rect 631 1978 635 1979
rect 631 1973 635 1974
rect 735 1978 739 1979
rect 735 1973 739 1974
rect 863 1978 867 1979
rect 863 1973 867 1974
rect 935 1978 939 1979
rect 935 1973 939 1974
rect 1071 1978 1075 1979
rect 1071 1973 1075 1974
rect 1127 1978 1131 1979
rect 1127 1973 1131 1974
rect 1263 1978 1267 1979
rect 1263 1973 1267 1974
rect 1303 1978 1307 1979
rect 1303 1973 1307 1974
rect 1447 1978 1451 1979
rect 1447 1973 1451 1974
rect 1471 1978 1475 1979
rect 1471 1973 1475 1974
rect 1615 1978 1619 1979
rect 1615 1973 1619 1974
rect 1631 1978 1635 1979
rect 1631 1973 1635 1974
rect 1783 1978 1787 1979
rect 1783 1973 1787 1974
rect 1791 1978 1795 1979
rect 1791 1973 1795 1974
rect 1935 1978 1939 1979
rect 1935 1973 1939 1974
rect 2031 1978 2035 1979
rect 2072 1974 2074 1989
rect 2528 1979 2530 1989
rect 2704 1979 2706 1989
rect 2888 1979 2890 1989
rect 3080 1979 3082 1989
rect 3280 1979 3282 1989
rect 3488 1979 3490 1989
rect 3704 1979 3706 1989
rect 3896 1979 3898 1989
rect 2526 1978 2532 1979
rect 2526 1974 2527 1978
rect 2531 1974 2532 1978
rect 2031 1973 2035 1974
rect 2070 1973 2076 1974
rect 2526 1973 2532 1974
rect 2702 1978 2708 1979
rect 2702 1974 2703 1978
rect 2707 1974 2708 1978
rect 2702 1973 2708 1974
rect 2886 1978 2892 1979
rect 2886 1974 2887 1978
rect 2891 1974 2892 1978
rect 2886 1973 2892 1974
rect 3078 1978 3084 1979
rect 3078 1974 3079 1978
rect 3083 1974 3084 1978
rect 3078 1973 3084 1974
rect 3278 1978 3284 1979
rect 3278 1974 3279 1978
rect 3283 1974 3284 1978
rect 3278 1973 3284 1974
rect 3486 1978 3492 1979
rect 3486 1974 3487 1978
rect 3491 1974 3492 1978
rect 3486 1973 3492 1974
rect 3702 1978 3708 1979
rect 3702 1974 3703 1978
rect 3707 1974 3708 1978
rect 3702 1973 3708 1974
rect 3894 1978 3900 1979
rect 3894 1974 3895 1978
rect 3899 1974 3900 1978
rect 3992 1974 3994 1989
rect 3894 1973 3900 1974
rect 3990 1973 3996 1974
rect 112 1958 114 1973
rect 152 1963 154 1973
rect 328 1963 330 1973
rect 536 1963 538 1973
rect 736 1963 738 1973
rect 936 1963 938 1973
rect 1128 1963 1130 1973
rect 1304 1963 1306 1973
rect 1472 1963 1474 1973
rect 1632 1963 1634 1973
rect 1792 1963 1794 1973
rect 1936 1963 1938 1973
rect 150 1962 156 1963
rect 150 1958 151 1962
rect 155 1958 156 1962
rect 110 1957 116 1958
rect 150 1957 156 1958
rect 326 1962 332 1963
rect 326 1958 327 1962
rect 331 1958 332 1962
rect 326 1957 332 1958
rect 534 1962 540 1963
rect 534 1958 535 1962
rect 539 1958 540 1962
rect 534 1957 540 1958
rect 734 1962 740 1963
rect 734 1958 735 1962
rect 739 1958 740 1962
rect 734 1957 740 1958
rect 934 1962 940 1963
rect 934 1958 935 1962
rect 939 1958 940 1962
rect 934 1957 940 1958
rect 1126 1962 1132 1963
rect 1126 1958 1127 1962
rect 1131 1958 1132 1962
rect 1126 1957 1132 1958
rect 1302 1962 1308 1963
rect 1302 1958 1303 1962
rect 1307 1958 1308 1962
rect 1302 1957 1308 1958
rect 1470 1962 1476 1963
rect 1470 1958 1471 1962
rect 1475 1958 1476 1962
rect 1470 1957 1476 1958
rect 1630 1962 1636 1963
rect 1630 1958 1631 1962
rect 1635 1958 1636 1962
rect 1630 1957 1636 1958
rect 1790 1962 1796 1963
rect 1790 1958 1791 1962
rect 1795 1958 1796 1962
rect 1790 1957 1796 1958
rect 1934 1962 1940 1963
rect 1934 1958 1935 1962
rect 1939 1958 1940 1962
rect 2032 1958 2034 1973
rect 2070 1969 2071 1973
rect 2075 1969 2076 1973
rect 2070 1968 2076 1969
rect 3990 1969 3991 1973
rect 3995 1969 3996 1973
rect 3990 1968 3996 1969
rect 1934 1957 1940 1958
rect 2030 1957 2036 1958
rect 110 1953 111 1957
rect 115 1953 116 1957
rect 110 1952 116 1953
rect 2030 1953 2031 1957
rect 2035 1953 2036 1957
rect 2030 1952 2036 1953
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2070 1951 2076 1952
rect 3990 1956 3996 1957
rect 3990 1952 3991 1956
rect 3995 1952 3996 1956
rect 3990 1951 3996 1952
rect 110 1940 116 1941
rect 110 1936 111 1940
rect 115 1936 116 1940
rect 110 1935 116 1936
rect 2030 1940 2036 1941
rect 2030 1936 2031 1940
rect 2035 1936 2036 1940
rect 2030 1935 2036 1936
rect 112 1903 114 1935
rect 150 1921 156 1922
rect 150 1917 151 1921
rect 155 1917 156 1921
rect 150 1916 156 1917
rect 326 1921 332 1922
rect 326 1917 327 1921
rect 331 1917 332 1921
rect 326 1916 332 1917
rect 534 1921 540 1922
rect 534 1917 535 1921
rect 539 1917 540 1921
rect 534 1916 540 1917
rect 734 1921 740 1922
rect 734 1917 735 1921
rect 739 1917 740 1921
rect 734 1916 740 1917
rect 934 1921 940 1922
rect 934 1917 935 1921
rect 939 1917 940 1921
rect 934 1916 940 1917
rect 1126 1921 1132 1922
rect 1126 1917 1127 1921
rect 1131 1917 1132 1921
rect 1126 1916 1132 1917
rect 1302 1921 1308 1922
rect 1302 1917 1303 1921
rect 1307 1917 1308 1921
rect 1302 1916 1308 1917
rect 1470 1921 1476 1922
rect 1470 1917 1471 1921
rect 1475 1917 1476 1921
rect 1470 1916 1476 1917
rect 1630 1921 1636 1922
rect 1630 1917 1631 1921
rect 1635 1917 1636 1921
rect 1630 1916 1636 1917
rect 1790 1921 1796 1922
rect 1790 1917 1791 1921
rect 1795 1917 1796 1921
rect 1790 1916 1796 1917
rect 1934 1921 1940 1922
rect 1934 1917 1935 1921
rect 1939 1917 1940 1921
rect 1934 1916 1940 1917
rect 152 1903 154 1916
rect 328 1903 330 1916
rect 536 1903 538 1916
rect 736 1903 738 1916
rect 936 1903 938 1916
rect 1128 1903 1130 1916
rect 1304 1903 1306 1916
rect 1472 1903 1474 1916
rect 1632 1903 1634 1916
rect 1792 1903 1794 1916
rect 1936 1903 1938 1916
rect 2032 1903 2034 1935
rect 2072 1919 2074 1951
rect 2526 1937 2532 1938
rect 2526 1933 2527 1937
rect 2531 1933 2532 1937
rect 2526 1932 2532 1933
rect 2702 1937 2708 1938
rect 2702 1933 2703 1937
rect 2707 1933 2708 1937
rect 2702 1932 2708 1933
rect 2886 1937 2892 1938
rect 2886 1933 2887 1937
rect 2891 1933 2892 1937
rect 2886 1932 2892 1933
rect 3078 1937 3084 1938
rect 3078 1933 3079 1937
rect 3083 1933 3084 1937
rect 3078 1932 3084 1933
rect 3278 1937 3284 1938
rect 3278 1933 3279 1937
rect 3283 1933 3284 1937
rect 3278 1932 3284 1933
rect 3486 1937 3492 1938
rect 3486 1933 3487 1937
rect 3491 1933 3492 1937
rect 3486 1932 3492 1933
rect 3702 1937 3708 1938
rect 3702 1933 3703 1937
rect 3707 1933 3708 1937
rect 3702 1932 3708 1933
rect 3894 1937 3900 1938
rect 3894 1933 3895 1937
rect 3899 1933 3900 1937
rect 3894 1932 3900 1933
rect 2528 1919 2530 1932
rect 2704 1919 2706 1932
rect 2888 1919 2890 1932
rect 3080 1919 3082 1932
rect 3280 1919 3282 1932
rect 3488 1919 3490 1932
rect 3704 1919 3706 1932
rect 3896 1919 3898 1932
rect 3992 1919 3994 1951
rect 2071 1918 2075 1919
rect 2071 1913 2075 1914
rect 2111 1918 2115 1919
rect 2111 1913 2115 1914
rect 2303 1918 2307 1919
rect 2303 1913 2307 1914
rect 2519 1918 2523 1919
rect 2519 1913 2523 1914
rect 2527 1918 2531 1919
rect 2527 1913 2531 1914
rect 2703 1918 2707 1919
rect 2703 1913 2707 1914
rect 2735 1918 2739 1919
rect 2735 1913 2739 1914
rect 2887 1918 2891 1919
rect 2887 1913 2891 1914
rect 2959 1918 2963 1919
rect 2959 1913 2963 1914
rect 3079 1918 3083 1919
rect 3079 1913 3083 1914
rect 3191 1918 3195 1919
rect 3191 1913 3195 1914
rect 3279 1918 3283 1919
rect 3279 1913 3283 1914
rect 3431 1918 3435 1919
rect 3431 1913 3435 1914
rect 3487 1918 3491 1919
rect 3487 1913 3491 1914
rect 3671 1918 3675 1919
rect 3671 1913 3675 1914
rect 3703 1918 3707 1919
rect 3703 1913 3707 1914
rect 3895 1918 3899 1919
rect 3895 1913 3899 1914
rect 3991 1918 3995 1919
rect 3991 1913 3995 1914
rect 111 1902 115 1903
rect 111 1897 115 1898
rect 151 1902 155 1903
rect 151 1897 155 1898
rect 303 1902 307 1903
rect 303 1897 307 1898
rect 327 1902 331 1903
rect 327 1897 331 1898
rect 463 1902 467 1903
rect 463 1897 467 1898
rect 535 1902 539 1903
rect 535 1897 539 1898
rect 615 1902 619 1903
rect 615 1897 619 1898
rect 735 1902 739 1903
rect 735 1897 739 1898
rect 767 1902 771 1903
rect 767 1897 771 1898
rect 927 1902 931 1903
rect 927 1897 931 1898
rect 935 1902 939 1903
rect 935 1897 939 1898
rect 1103 1902 1107 1903
rect 1103 1897 1107 1898
rect 1127 1902 1131 1903
rect 1127 1897 1131 1898
rect 1295 1902 1299 1903
rect 1295 1897 1299 1898
rect 1303 1902 1307 1903
rect 1303 1897 1307 1898
rect 1471 1902 1475 1903
rect 1471 1897 1475 1898
rect 1511 1902 1515 1903
rect 1511 1897 1515 1898
rect 1631 1902 1635 1903
rect 1631 1897 1635 1898
rect 1735 1902 1739 1903
rect 1735 1897 1739 1898
rect 1791 1902 1795 1903
rect 1791 1897 1795 1898
rect 1935 1902 1939 1903
rect 1935 1897 1939 1898
rect 2031 1902 2035 1903
rect 2031 1897 2035 1898
rect 112 1869 114 1897
rect 152 1888 154 1897
rect 304 1888 306 1897
rect 464 1888 466 1897
rect 616 1888 618 1897
rect 768 1888 770 1897
rect 928 1888 930 1897
rect 1104 1888 1106 1897
rect 1296 1888 1298 1897
rect 1512 1888 1514 1897
rect 1736 1888 1738 1897
rect 1936 1888 1938 1897
rect 150 1887 156 1888
rect 150 1883 151 1887
rect 155 1883 156 1887
rect 150 1882 156 1883
rect 302 1887 308 1888
rect 302 1883 303 1887
rect 307 1883 308 1887
rect 302 1882 308 1883
rect 462 1887 468 1888
rect 462 1883 463 1887
rect 467 1883 468 1887
rect 462 1882 468 1883
rect 614 1887 620 1888
rect 614 1883 615 1887
rect 619 1883 620 1887
rect 614 1882 620 1883
rect 766 1887 772 1888
rect 766 1883 767 1887
rect 771 1883 772 1887
rect 766 1882 772 1883
rect 926 1887 932 1888
rect 926 1883 927 1887
rect 931 1883 932 1887
rect 926 1882 932 1883
rect 1102 1887 1108 1888
rect 1102 1883 1103 1887
rect 1107 1883 1108 1887
rect 1102 1882 1108 1883
rect 1294 1887 1300 1888
rect 1294 1883 1295 1887
rect 1299 1883 1300 1887
rect 1294 1882 1300 1883
rect 1510 1887 1516 1888
rect 1510 1883 1511 1887
rect 1515 1883 1516 1887
rect 1510 1882 1516 1883
rect 1734 1887 1740 1888
rect 1734 1883 1735 1887
rect 1739 1883 1740 1887
rect 1734 1882 1740 1883
rect 1934 1887 1940 1888
rect 1934 1883 1935 1887
rect 1939 1883 1940 1887
rect 1934 1882 1940 1883
rect 2032 1869 2034 1897
rect 2072 1885 2074 1913
rect 2112 1904 2114 1913
rect 2304 1904 2306 1913
rect 2520 1904 2522 1913
rect 2736 1904 2738 1913
rect 2960 1904 2962 1913
rect 3192 1904 3194 1913
rect 3432 1904 3434 1913
rect 3672 1904 3674 1913
rect 3896 1904 3898 1913
rect 2110 1903 2116 1904
rect 2110 1899 2111 1903
rect 2115 1899 2116 1903
rect 2110 1898 2116 1899
rect 2302 1903 2308 1904
rect 2302 1899 2303 1903
rect 2307 1899 2308 1903
rect 2302 1898 2308 1899
rect 2518 1903 2524 1904
rect 2518 1899 2519 1903
rect 2523 1899 2524 1903
rect 2518 1898 2524 1899
rect 2734 1903 2740 1904
rect 2734 1899 2735 1903
rect 2739 1899 2740 1903
rect 2734 1898 2740 1899
rect 2958 1903 2964 1904
rect 2958 1899 2959 1903
rect 2963 1899 2964 1903
rect 2958 1898 2964 1899
rect 3190 1903 3196 1904
rect 3190 1899 3191 1903
rect 3195 1899 3196 1903
rect 3190 1898 3196 1899
rect 3430 1903 3436 1904
rect 3430 1899 3431 1903
rect 3435 1899 3436 1903
rect 3430 1898 3436 1899
rect 3670 1903 3676 1904
rect 3670 1899 3671 1903
rect 3675 1899 3676 1903
rect 3670 1898 3676 1899
rect 3894 1903 3900 1904
rect 3894 1899 3895 1903
rect 3899 1899 3900 1903
rect 3894 1898 3900 1899
rect 3992 1885 3994 1913
rect 2070 1884 2076 1885
rect 2070 1880 2071 1884
rect 2075 1880 2076 1884
rect 2070 1879 2076 1880
rect 3990 1884 3996 1885
rect 3990 1880 3991 1884
rect 3995 1880 3996 1884
rect 3990 1879 3996 1880
rect 110 1868 116 1869
rect 110 1864 111 1868
rect 115 1864 116 1868
rect 110 1863 116 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2070 1867 2076 1868
rect 2070 1863 2071 1867
rect 2075 1863 2076 1867
rect 3990 1867 3996 1868
rect 3990 1863 3991 1867
rect 3995 1863 3996 1867
rect 2070 1862 2076 1863
rect 2110 1862 2116 1863
rect 110 1851 116 1852
rect 110 1847 111 1851
rect 115 1847 116 1851
rect 2030 1851 2036 1852
rect 2030 1847 2031 1851
rect 2035 1847 2036 1851
rect 2072 1847 2074 1862
rect 2110 1858 2111 1862
rect 2115 1858 2116 1862
rect 2110 1857 2116 1858
rect 2302 1862 2308 1863
rect 2302 1858 2303 1862
rect 2307 1858 2308 1862
rect 2302 1857 2308 1858
rect 2518 1862 2524 1863
rect 2518 1858 2519 1862
rect 2523 1858 2524 1862
rect 2518 1857 2524 1858
rect 2734 1862 2740 1863
rect 2734 1858 2735 1862
rect 2739 1858 2740 1862
rect 2734 1857 2740 1858
rect 2958 1862 2964 1863
rect 2958 1858 2959 1862
rect 2963 1858 2964 1862
rect 2958 1857 2964 1858
rect 3190 1862 3196 1863
rect 3190 1858 3191 1862
rect 3195 1858 3196 1862
rect 3190 1857 3196 1858
rect 3430 1862 3436 1863
rect 3430 1858 3431 1862
rect 3435 1858 3436 1862
rect 3430 1857 3436 1858
rect 3670 1862 3676 1863
rect 3670 1858 3671 1862
rect 3675 1858 3676 1862
rect 3670 1857 3676 1858
rect 3894 1862 3900 1863
rect 3990 1862 3996 1863
rect 3894 1858 3895 1862
rect 3899 1858 3900 1862
rect 3894 1857 3900 1858
rect 2112 1847 2114 1857
rect 2304 1847 2306 1857
rect 2520 1847 2522 1857
rect 2736 1847 2738 1857
rect 2960 1847 2962 1857
rect 3192 1847 3194 1857
rect 3432 1847 3434 1857
rect 3672 1847 3674 1857
rect 3896 1847 3898 1857
rect 3992 1847 3994 1862
rect 110 1846 116 1847
rect 150 1846 156 1847
rect 112 1819 114 1846
rect 150 1842 151 1846
rect 155 1842 156 1846
rect 150 1841 156 1842
rect 302 1846 308 1847
rect 302 1842 303 1846
rect 307 1842 308 1846
rect 302 1841 308 1842
rect 462 1846 468 1847
rect 462 1842 463 1846
rect 467 1842 468 1846
rect 462 1841 468 1842
rect 614 1846 620 1847
rect 614 1842 615 1846
rect 619 1842 620 1846
rect 614 1841 620 1842
rect 766 1846 772 1847
rect 766 1842 767 1846
rect 771 1842 772 1846
rect 766 1841 772 1842
rect 926 1846 932 1847
rect 926 1842 927 1846
rect 931 1842 932 1846
rect 926 1841 932 1842
rect 1102 1846 1108 1847
rect 1102 1842 1103 1846
rect 1107 1842 1108 1846
rect 1102 1841 1108 1842
rect 1294 1846 1300 1847
rect 1294 1842 1295 1846
rect 1299 1842 1300 1846
rect 1294 1841 1300 1842
rect 1510 1846 1516 1847
rect 1510 1842 1511 1846
rect 1515 1842 1516 1846
rect 1510 1841 1516 1842
rect 1734 1846 1740 1847
rect 1734 1842 1735 1846
rect 1739 1842 1740 1846
rect 1734 1841 1740 1842
rect 1934 1846 1940 1847
rect 2030 1846 2036 1847
rect 2071 1846 2075 1847
rect 1934 1842 1935 1846
rect 1939 1842 1940 1846
rect 1934 1841 1940 1842
rect 152 1819 154 1841
rect 304 1819 306 1841
rect 464 1819 466 1841
rect 616 1819 618 1841
rect 768 1819 770 1841
rect 928 1819 930 1841
rect 1104 1819 1106 1841
rect 1296 1819 1298 1841
rect 1512 1819 1514 1841
rect 1736 1819 1738 1841
rect 1936 1819 1938 1841
rect 2032 1819 2034 1846
rect 2071 1841 2075 1842
rect 2111 1846 2115 1847
rect 2111 1841 2115 1842
rect 2231 1846 2235 1847
rect 2231 1841 2235 1842
rect 2303 1846 2307 1847
rect 2303 1841 2307 1842
rect 2399 1846 2403 1847
rect 2399 1841 2403 1842
rect 2519 1846 2523 1847
rect 2519 1841 2523 1842
rect 2599 1846 2603 1847
rect 2599 1841 2603 1842
rect 2735 1846 2739 1847
rect 2735 1841 2739 1842
rect 2831 1846 2835 1847
rect 2831 1841 2835 1842
rect 2959 1846 2963 1847
rect 2959 1841 2963 1842
rect 3079 1846 3083 1847
rect 3079 1841 3083 1842
rect 3191 1846 3195 1847
rect 3191 1841 3195 1842
rect 3351 1846 3355 1847
rect 3351 1841 3355 1842
rect 3431 1846 3435 1847
rect 3431 1841 3435 1842
rect 3631 1846 3635 1847
rect 3631 1841 3635 1842
rect 3671 1846 3675 1847
rect 3671 1841 3675 1842
rect 3895 1846 3899 1847
rect 3895 1841 3899 1842
rect 3991 1846 3995 1847
rect 3991 1841 3995 1842
rect 2072 1826 2074 1841
rect 2112 1831 2114 1841
rect 2232 1831 2234 1841
rect 2400 1831 2402 1841
rect 2600 1831 2602 1841
rect 2832 1831 2834 1841
rect 3080 1831 3082 1841
rect 3352 1831 3354 1841
rect 3632 1831 3634 1841
rect 3896 1831 3898 1841
rect 2110 1830 2116 1831
rect 2110 1826 2111 1830
rect 2115 1826 2116 1830
rect 2070 1825 2076 1826
rect 2110 1825 2116 1826
rect 2230 1830 2236 1831
rect 2230 1826 2231 1830
rect 2235 1826 2236 1830
rect 2230 1825 2236 1826
rect 2398 1830 2404 1831
rect 2398 1826 2399 1830
rect 2403 1826 2404 1830
rect 2398 1825 2404 1826
rect 2598 1830 2604 1831
rect 2598 1826 2599 1830
rect 2603 1826 2604 1830
rect 2598 1825 2604 1826
rect 2830 1830 2836 1831
rect 2830 1826 2831 1830
rect 2835 1826 2836 1830
rect 2830 1825 2836 1826
rect 3078 1830 3084 1831
rect 3078 1826 3079 1830
rect 3083 1826 3084 1830
rect 3078 1825 3084 1826
rect 3350 1830 3356 1831
rect 3350 1826 3351 1830
rect 3355 1826 3356 1830
rect 3350 1825 3356 1826
rect 3630 1830 3636 1831
rect 3630 1826 3631 1830
rect 3635 1826 3636 1830
rect 3630 1825 3636 1826
rect 3894 1830 3900 1831
rect 3894 1826 3895 1830
rect 3899 1826 3900 1830
rect 3992 1826 3994 1841
rect 3894 1825 3900 1826
rect 3990 1825 3996 1826
rect 2070 1821 2071 1825
rect 2075 1821 2076 1825
rect 2070 1820 2076 1821
rect 3990 1821 3991 1825
rect 3995 1821 3996 1825
rect 3990 1820 3996 1821
rect 111 1818 115 1819
rect 111 1813 115 1814
rect 151 1818 155 1819
rect 151 1813 155 1814
rect 303 1818 307 1819
rect 303 1813 307 1814
rect 343 1818 347 1819
rect 343 1813 347 1814
rect 463 1818 467 1819
rect 463 1813 467 1814
rect 543 1818 547 1819
rect 543 1813 547 1814
rect 615 1818 619 1819
rect 615 1813 619 1814
rect 735 1818 739 1819
rect 735 1813 739 1814
rect 767 1818 771 1819
rect 767 1813 771 1814
rect 919 1818 923 1819
rect 919 1813 923 1814
rect 927 1818 931 1819
rect 927 1813 931 1814
rect 1095 1818 1099 1819
rect 1095 1813 1099 1814
rect 1103 1818 1107 1819
rect 1103 1813 1107 1814
rect 1271 1818 1275 1819
rect 1271 1813 1275 1814
rect 1295 1818 1299 1819
rect 1295 1813 1299 1814
rect 1447 1818 1451 1819
rect 1447 1813 1451 1814
rect 1511 1818 1515 1819
rect 1511 1813 1515 1814
rect 1623 1818 1627 1819
rect 1623 1813 1627 1814
rect 1735 1818 1739 1819
rect 1735 1813 1739 1814
rect 1807 1818 1811 1819
rect 1807 1813 1811 1814
rect 1935 1818 1939 1819
rect 1935 1813 1939 1814
rect 2031 1818 2035 1819
rect 2031 1813 2035 1814
rect 112 1798 114 1813
rect 152 1803 154 1813
rect 344 1803 346 1813
rect 544 1803 546 1813
rect 736 1803 738 1813
rect 920 1803 922 1813
rect 1096 1803 1098 1813
rect 1272 1803 1274 1813
rect 1448 1803 1450 1813
rect 1624 1803 1626 1813
rect 1808 1803 1810 1813
rect 150 1802 156 1803
rect 150 1798 151 1802
rect 155 1798 156 1802
rect 110 1797 116 1798
rect 150 1797 156 1798
rect 342 1802 348 1803
rect 342 1798 343 1802
rect 347 1798 348 1802
rect 342 1797 348 1798
rect 542 1802 548 1803
rect 542 1798 543 1802
rect 547 1798 548 1802
rect 542 1797 548 1798
rect 734 1802 740 1803
rect 734 1798 735 1802
rect 739 1798 740 1802
rect 734 1797 740 1798
rect 918 1802 924 1803
rect 918 1798 919 1802
rect 923 1798 924 1802
rect 918 1797 924 1798
rect 1094 1802 1100 1803
rect 1094 1798 1095 1802
rect 1099 1798 1100 1802
rect 1094 1797 1100 1798
rect 1270 1802 1276 1803
rect 1270 1798 1271 1802
rect 1275 1798 1276 1802
rect 1270 1797 1276 1798
rect 1446 1802 1452 1803
rect 1446 1798 1447 1802
rect 1451 1798 1452 1802
rect 1446 1797 1452 1798
rect 1622 1802 1628 1803
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1806 1802 1812 1803
rect 1806 1798 1807 1802
rect 1811 1798 1812 1802
rect 2032 1798 2034 1813
rect 2070 1808 2076 1809
rect 2070 1804 2071 1808
rect 2075 1804 2076 1808
rect 2070 1803 2076 1804
rect 3990 1808 3996 1809
rect 3990 1804 3991 1808
rect 3995 1804 3996 1808
rect 3990 1803 3996 1804
rect 1806 1797 1812 1798
rect 2030 1797 2036 1798
rect 110 1793 111 1797
rect 115 1793 116 1797
rect 110 1792 116 1793
rect 2030 1793 2031 1797
rect 2035 1793 2036 1797
rect 2030 1792 2036 1793
rect 110 1780 116 1781
rect 110 1776 111 1780
rect 115 1776 116 1780
rect 110 1775 116 1776
rect 2030 1780 2036 1781
rect 2030 1776 2031 1780
rect 2035 1776 2036 1780
rect 2030 1775 2036 1776
rect 112 1743 114 1775
rect 150 1761 156 1762
rect 150 1757 151 1761
rect 155 1757 156 1761
rect 150 1756 156 1757
rect 342 1761 348 1762
rect 342 1757 343 1761
rect 347 1757 348 1761
rect 342 1756 348 1757
rect 542 1761 548 1762
rect 542 1757 543 1761
rect 547 1757 548 1761
rect 542 1756 548 1757
rect 734 1761 740 1762
rect 734 1757 735 1761
rect 739 1757 740 1761
rect 734 1756 740 1757
rect 918 1761 924 1762
rect 918 1757 919 1761
rect 923 1757 924 1761
rect 918 1756 924 1757
rect 1094 1761 1100 1762
rect 1094 1757 1095 1761
rect 1099 1757 1100 1761
rect 1094 1756 1100 1757
rect 1270 1761 1276 1762
rect 1270 1757 1271 1761
rect 1275 1757 1276 1761
rect 1270 1756 1276 1757
rect 1446 1761 1452 1762
rect 1446 1757 1447 1761
rect 1451 1757 1452 1761
rect 1446 1756 1452 1757
rect 1622 1761 1628 1762
rect 1622 1757 1623 1761
rect 1627 1757 1628 1761
rect 1622 1756 1628 1757
rect 1806 1761 1812 1762
rect 1806 1757 1807 1761
rect 1811 1757 1812 1761
rect 1806 1756 1812 1757
rect 152 1743 154 1756
rect 344 1743 346 1756
rect 544 1743 546 1756
rect 736 1743 738 1756
rect 920 1743 922 1756
rect 1096 1743 1098 1756
rect 1272 1743 1274 1756
rect 1448 1743 1450 1756
rect 1624 1743 1626 1756
rect 1808 1743 1810 1756
rect 2032 1743 2034 1775
rect 2072 1771 2074 1803
rect 2110 1789 2116 1790
rect 2110 1785 2111 1789
rect 2115 1785 2116 1789
rect 2110 1784 2116 1785
rect 2230 1789 2236 1790
rect 2230 1785 2231 1789
rect 2235 1785 2236 1789
rect 2230 1784 2236 1785
rect 2398 1789 2404 1790
rect 2398 1785 2399 1789
rect 2403 1785 2404 1789
rect 2398 1784 2404 1785
rect 2598 1789 2604 1790
rect 2598 1785 2599 1789
rect 2603 1785 2604 1789
rect 2598 1784 2604 1785
rect 2830 1789 2836 1790
rect 2830 1785 2831 1789
rect 2835 1785 2836 1789
rect 2830 1784 2836 1785
rect 3078 1789 3084 1790
rect 3078 1785 3079 1789
rect 3083 1785 3084 1789
rect 3078 1784 3084 1785
rect 3350 1789 3356 1790
rect 3350 1785 3351 1789
rect 3355 1785 3356 1789
rect 3350 1784 3356 1785
rect 3630 1789 3636 1790
rect 3630 1785 3631 1789
rect 3635 1785 3636 1789
rect 3630 1784 3636 1785
rect 3894 1789 3900 1790
rect 3894 1785 3895 1789
rect 3899 1785 3900 1789
rect 3894 1784 3900 1785
rect 2112 1771 2114 1784
rect 2232 1771 2234 1784
rect 2400 1771 2402 1784
rect 2600 1771 2602 1784
rect 2832 1771 2834 1784
rect 3080 1771 3082 1784
rect 3352 1771 3354 1784
rect 3632 1771 3634 1784
rect 3896 1771 3898 1784
rect 3992 1771 3994 1803
rect 2071 1770 2075 1771
rect 2071 1765 2075 1766
rect 2111 1770 2115 1771
rect 2111 1765 2115 1766
rect 2231 1770 2235 1771
rect 2231 1765 2235 1766
rect 2239 1770 2243 1771
rect 2239 1765 2243 1766
rect 2399 1770 2403 1771
rect 2399 1765 2403 1766
rect 2575 1770 2579 1771
rect 2575 1765 2579 1766
rect 2599 1770 2603 1771
rect 2599 1765 2603 1766
rect 2751 1770 2755 1771
rect 2751 1765 2755 1766
rect 2831 1770 2835 1771
rect 2831 1765 2835 1766
rect 2935 1770 2939 1771
rect 2935 1765 2939 1766
rect 3079 1770 3083 1771
rect 3079 1765 3083 1766
rect 3127 1770 3131 1771
rect 3127 1765 3131 1766
rect 3319 1770 3323 1771
rect 3319 1765 3323 1766
rect 3351 1770 3355 1771
rect 3351 1765 3355 1766
rect 3511 1770 3515 1771
rect 3511 1765 3515 1766
rect 3631 1770 3635 1771
rect 3631 1765 3635 1766
rect 3711 1770 3715 1771
rect 3711 1765 3715 1766
rect 3895 1770 3899 1771
rect 3895 1765 3899 1766
rect 3991 1770 3995 1771
rect 3991 1765 3995 1766
rect 111 1742 115 1743
rect 111 1737 115 1738
rect 151 1742 155 1743
rect 151 1737 155 1738
rect 319 1742 323 1743
rect 319 1737 323 1738
rect 343 1742 347 1743
rect 343 1737 347 1738
rect 527 1742 531 1743
rect 527 1737 531 1738
rect 543 1742 547 1743
rect 543 1737 547 1738
rect 735 1742 739 1743
rect 735 1737 739 1738
rect 743 1742 747 1743
rect 743 1737 747 1738
rect 919 1742 923 1743
rect 919 1737 923 1738
rect 959 1742 963 1743
rect 959 1737 963 1738
rect 1095 1742 1099 1743
rect 1095 1737 1099 1738
rect 1167 1742 1171 1743
rect 1167 1737 1171 1738
rect 1271 1742 1275 1743
rect 1271 1737 1275 1738
rect 1367 1742 1371 1743
rect 1367 1737 1371 1738
rect 1447 1742 1451 1743
rect 1447 1737 1451 1738
rect 1559 1742 1563 1743
rect 1559 1737 1563 1738
rect 1623 1742 1627 1743
rect 1623 1737 1627 1738
rect 1759 1742 1763 1743
rect 1759 1737 1763 1738
rect 1807 1742 1811 1743
rect 1807 1737 1811 1738
rect 1935 1742 1939 1743
rect 1935 1737 1939 1738
rect 2031 1742 2035 1743
rect 2031 1737 2035 1738
rect 2072 1737 2074 1765
rect 2112 1756 2114 1765
rect 2240 1756 2242 1765
rect 2400 1756 2402 1765
rect 2576 1756 2578 1765
rect 2752 1756 2754 1765
rect 2936 1756 2938 1765
rect 3128 1756 3130 1765
rect 3320 1756 3322 1765
rect 3512 1756 3514 1765
rect 3712 1756 3714 1765
rect 3896 1756 3898 1765
rect 2110 1755 2116 1756
rect 2110 1751 2111 1755
rect 2115 1751 2116 1755
rect 2110 1750 2116 1751
rect 2238 1755 2244 1756
rect 2238 1751 2239 1755
rect 2243 1751 2244 1755
rect 2238 1750 2244 1751
rect 2398 1755 2404 1756
rect 2398 1751 2399 1755
rect 2403 1751 2404 1755
rect 2398 1750 2404 1751
rect 2574 1755 2580 1756
rect 2574 1751 2575 1755
rect 2579 1751 2580 1755
rect 2574 1750 2580 1751
rect 2750 1755 2756 1756
rect 2750 1751 2751 1755
rect 2755 1751 2756 1755
rect 2750 1750 2756 1751
rect 2934 1755 2940 1756
rect 2934 1751 2935 1755
rect 2939 1751 2940 1755
rect 2934 1750 2940 1751
rect 3126 1755 3132 1756
rect 3126 1751 3127 1755
rect 3131 1751 3132 1755
rect 3126 1750 3132 1751
rect 3318 1755 3324 1756
rect 3318 1751 3319 1755
rect 3323 1751 3324 1755
rect 3318 1750 3324 1751
rect 3510 1755 3516 1756
rect 3510 1751 3511 1755
rect 3515 1751 3516 1755
rect 3510 1750 3516 1751
rect 3710 1755 3716 1756
rect 3710 1751 3711 1755
rect 3715 1751 3716 1755
rect 3710 1750 3716 1751
rect 3894 1755 3900 1756
rect 3894 1751 3895 1755
rect 3899 1751 3900 1755
rect 3894 1750 3900 1751
rect 3992 1737 3994 1765
rect 112 1709 114 1737
rect 152 1728 154 1737
rect 320 1728 322 1737
rect 528 1728 530 1737
rect 744 1728 746 1737
rect 960 1728 962 1737
rect 1168 1728 1170 1737
rect 1368 1728 1370 1737
rect 1560 1728 1562 1737
rect 1760 1728 1762 1737
rect 1936 1728 1938 1737
rect 150 1727 156 1728
rect 150 1723 151 1727
rect 155 1723 156 1727
rect 150 1722 156 1723
rect 318 1727 324 1728
rect 318 1723 319 1727
rect 323 1723 324 1727
rect 318 1722 324 1723
rect 526 1727 532 1728
rect 526 1723 527 1727
rect 531 1723 532 1727
rect 526 1722 532 1723
rect 742 1727 748 1728
rect 742 1723 743 1727
rect 747 1723 748 1727
rect 742 1722 748 1723
rect 958 1727 964 1728
rect 958 1723 959 1727
rect 963 1723 964 1727
rect 958 1722 964 1723
rect 1166 1727 1172 1728
rect 1166 1723 1167 1727
rect 1171 1723 1172 1727
rect 1166 1722 1172 1723
rect 1366 1727 1372 1728
rect 1366 1723 1367 1727
rect 1371 1723 1372 1727
rect 1366 1722 1372 1723
rect 1558 1727 1564 1728
rect 1558 1723 1559 1727
rect 1563 1723 1564 1727
rect 1558 1722 1564 1723
rect 1758 1727 1764 1728
rect 1758 1723 1759 1727
rect 1763 1723 1764 1727
rect 1758 1722 1764 1723
rect 1934 1727 1940 1728
rect 1934 1723 1935 1727
rect 1939 1723 1940 1727
rect 1934 1722 1940 1723
rect 2032 1709 2034 1737
rect 2070 1736 2076 1737
rect 2070 1732 2071 1736
rect 2075 1732 2076 1736
rect 2070 1731 2076 1732
rect 3990 1736 3996 1737
rect 3990 1732 3991 1736
rect 3995 1732 3996 1736
rect 3990 1731 3996 1732
rect 2070 1719 2076 1720
rect 2070 1715 2071 1719
rect 2075 1715 2076 1719
rect 3990 1719 3996 1720
rect 3990 1715 3991 1719
rect 3995 1715 3996 1719
rect 2070 1714 2076 1715
rect 2110 1714 2116 1715
rect 110 1708 116 1709
rect 110 1704 111 1708
rect 115 1704 116 1708
rect 110 1703 116 1704
rect 2030 1708 2036 1709
rect 2030 1704 2031 1708
rect 2035 1704 2036 1708
rect 2030 1703 2036 1704
rect 110 1691 116 1692
rect 110 1687 111 1691
rect 115 1687 116 1691
rect 2030 1691 2036 1692
rect 2072 1691 2074 1714
rect 2110 1710 2111 1714
rect 2115 1710 2116 1714
rect 2110 1709 2116 1710
rect 2238 1714 2244 1715
rect 2238 1710 2239 1714
rect 2243 1710 2244 1714
rect 2238 1709 2244 1710
rect 2398 1714 2404 1715
rect 2398 1710 2399 1714
rect 2403 1710 2404 1714
rect 2398 1709 2404 1710
rect 2574 1714 2580 1715
rect 2574 1710 2575 1714
rect 2579 1710 2580 1714
rect 2574 1709 2580 1710
rect 2750 1714 2756 1715
rect 2750 1710 2751 1714
rect 2755 1710 2756 1714
rect 2750 1709 2756 1710
rect 2934 1714 2940 1715
rect 2934 1710 2935 1714
rect 2939 1710 2940 1714
rect 2934 1709 2940 1710
rect 3126 1714 3132 1715
rect 3126 1710 3127 1714
rect 3131 1710 3132 1714
rect 3126 1709 3132 1710
rect 3318 1714 3324 1715
rect 3318 1710 3319 1714
rect 3323 1710 3324 1714
rect 3318 1709 3324 1710
rect 3510 1714 3516 1715
rect 3510 1710 3511 1714
rect 3515 1710 3516 1714
rect 3510 1709 3516 1710
rect 3710 1714 3716 1715
rect 3710 1710 3711 1714
rect 3715 1710 3716 1714
rect 3710 1709 3716 1710
rect 3894 1714 3900 1715
rect 3990 1714 3996 1715
rect 3894 1710 3895 1714
rect 3899 1710 3900 1714
rect 3894 1709 3900 1710
rect 2112 1691 2114 1709
rect 2240 1691 2242 1709
rect 2400 1691 2402 1709
rect 2576 1691 2578 1709
rect 2752 1691 2754 1709
rect 2936 1691 2938 1709
rect 3128 1691 3130 1709
rect 3320 1691 3322 1709
rect 3512 1691 3514 1709
rect 3712 1691 3714 1709
rect 3896 1691 3898 1709
rect 3992 1691 3994 1714
rect 2030 1687 2031 1691
rect 2035 1687 2036 1691
rect 110 1686 116 1687
rect 150 1686 156 1687
rect 112 1671 114 1686
rect 150 1682 151 1686
rect 155 1682 156 1686
rect 150 1681 156 1682
rect 318 1686 324 1687
rect 318 1682 319 1686
rect 323 1682 324 1686
rect 318 1681 324 1682
rect 526 1686 532 1687
rect 526 1682 527 1686
rect 531 1682 532 1686
rect 526 1681 532 1682
rect 742 1686 748 1687
rect 742 1682 743 1686
rect 747 1682 748 1686
rect 742 1681 748 1682
rect 958 1686 964 1687
rect 958 1682 959 1686
rect 963 1682 964 1686
rect 958 1681 964 1682
rect 1166 1686 1172 1687
rect 1166 1682 1167 1686
rect 1171 1682 1172 1686
rect 1166 1681 1172 1682
rect 1366 1686 1372 1687
rect 1366 1682 1367 1686
rect 1371 1682 1372 1686
rect 1366 1681 1372 1682
rect 1558 1686 1564 1687
rect 1558 1682 1559 1686
rect 1563 1682 1564 1686
rect 1558 1681 1564 1682
rect 1758 1686 1764 1687
rect 1758 1682 1759 1686
rect 1763 1682 1764 1686
rect 1758 1681 1764 1682
rect 1934 1686 1940 1687
rect 2030 1686 2036 1687
rect 2071 1690 2075 1691
rect 1934 1682 1935 1686
rect 1939 1682 1940 1686
rect 1934 1681 1940 1682
rect 152 1671 154 1681
rect 320 1671 322 1681
rect 528 1671 530 1681
rect 744 1671 746 1681
rect 960 1671 962 1681
rect 1168 1671 1170 1681
rect 1368 1671 1370 1681
rect 1560 1671 1562 1681
rect 1760 1671 1762 1681
rect 1936 1671 1938 1681
rect 2032 1671 2034 1686
rect 2071 1685 2075 1686
rect 2111 1690 2115 1691
rect 2111 1685 2115 1686
rect 2239 1690 2243 1691
rect 2239 1685 2243 1686
rect 2311 1690 2315 1691
rect 2311 1685 2315 1686
rect 2399 1690 2403 1691
rect 2399 1685 2403 1686
rect 2527 1690 2531 1691
rect 2527 1685 2531 1686
rect 2575 1690 2579 1691
rect 2575 1685 2579 1686
rect 2743 1690 2747 1691
rect 2743 1685 2747 1686
rect 2751 1690 2755 1691
rect 2751 1685 2755 1686
rect 2935 1690 2939 1691
rect 2935 1685 2939 1686
rect 2951 1690 2955 1691
rect 2951 1685 2955 1686
rect 3127 1690 3131 1691
rect 3127 1685 3131 1686
rect 3151 1690 3155 1691
rect 3151 1685 3155 1686
rect 3319 1690 3323 1691
rect 3319 1685 3323 1686
rect 3343 1690 3347 1691
rect 3343 1685 3347 1686
rect 3511 1690 3515 1691
rect 3511 1685 3515 1686
rect 3527 1690 3531 1691
rect 3527 1685 3531 1686
rect 3711 1690 3715 1691
rect 3711 1685 3715 1686
rect 3719 1690 3723 1691
rect 3719 1685 3723 1686
rect 3895 1690 3899 1691
rect 3895 1685 3899 1686
rect 3991 1690 3995 1691
rect 3991 1685 3995 1686
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 151 1670 155 1671
rect 151 1665 155 1666
rect 319 1670 323 1671
rect 319 1665 323 1666
rect 503 1670 507 1671
rect 503 1665 507 1666
rect 527 1670 531 1671
rect 527 1665 531 1666
rect 695 1670 699 1671
rect 695 1665 699 1666
rect 743 1670 747 1671
rect 743 1665 747 1666
rect 887 1670 891 1671
rect 887 1665 891 1666
rect 959 1670 963 1671
rect 959 1665 963 1666
rect 1079 1670 1083 1671
rect 1079 1665 1083 1666
rect 1167 1670 1171 1671
rect 1167 1665 1171 1666
rect 1263 1670 1267 1671
rect 1263 1665 1267 1666
rect 1367 1670 1371 1671
rect 1367 1665 1371 1666
rect 1439 1670 1443 1671
rect 1439 1665 1443 1666
rect 1559 1670 1563 1671
rect 1559 1665 1563 1666
rect 1615 1670 1619 1671
rect 1615 1665 1619 1666
rect 1759 1670 1763 1671
rect 1759 1665 1763 1666
rect 1791 1670 1795 1671
rect 1791 1665 1795 1666
rect 1935 1670 1939 1671
rect 1935 1665 1939 1666
rect 2031 1670 2035 1671
rect 2072 1670 2074 1685
rect 2112 1675 2114 1685
rect 2312 1675 2314 1685
rect 2528 1675 2530 1685
rect 2744 1675 2746 1685
rect 2952 1675 2954 1685
rect 3152 1675 3154 1685
rect 3344 1675 3346 1685
rect 3528 1675 3530 1685
rect 3720 1675 3722 1685
rect 3896 1675 3898 1685
rect 2110 1674 2116 1675
rect 2110 1670 2111 1674
rect 2115 1670 2116 1674
rect 2031 1665 2035 1666
rect 2070 1669 2076 1670
rect 2110 1669 2116 1670
rect 2310 1674 2316 1675
rect 2310 1670 2311 1674
rect 2315 1670 2316 1674
rect 2310 1669 2316 1670
rect 2526 1674 2532 1675
rect 2526 1670 2527 1674
rect 2531 1670 2532 1674
rect 2526 1669 2532 1670
rect 2742 1674 2748 1675
rect 2742 1670 2743 1674
rect 2747 1670 2748 1674
rect 2742 1669 2748 1670
rect 2950 1674 2956 1675
rect 2950 1670 2951 1674
rect 2955 1670 2956 1674
rect 2950 1669 2956 1670
rect 3150 1674 3156 1675
rect 3150 1670 3151 1674
rect 3155 1670 3156 1674
rect 3150 1669 3156 1670
rect 3342 1674 3348 1675
rect 3342 1670 3343 1674
rect 3347 1670 3348 1674
rect 3342 1669 3348 1670
rect 3526 1674 3532 1675
rect 3526 1670 3527 1674
rect 3531 1670 3532 1674
rect 3526 1669 3532 1670
rect 3718 1674 3724 1675
rect 3718 1670 3719 1674
rect 3723 1670 3724 1674
rect 3718 1669 3724 1670
rect 3894 1674 3900 1675
rect 3894 1670 3895 1674
rect 3899 1670 3900 1674
rect 3992 1670 3994 1685
rect 3894 1669 3900 1670
rect 3990 1669 3996 1670
rect 2070 1665 2071 1669
rect 2075 1665 2076 1669
rect 112 1650 114 1665
rect 152 1655 154 1665
rect 320 1655 322 1665
rect 504 1655 506 1665
rect 696 1655 698 1665
rect 888 1655 890 1665
rect 1080 1655 1082 1665
rect 1264 1655 1266 1665
rect 1440 1655 1442 1665
rect 1616 1655 1618 1665
rect 1792 1655 1794 1665
rect 150 1654 156 1655
rect 150 1650 151 1654
rect 155 1650 156 1654
rect 110 1649 116 1650
rect 150 1649 156 1650
rect 318 1654 324 1655
rect 318 1650 319 1654
rect 323 1650 324 1654
rect 318 1649 324 1650
rect 502 1654 508 1655
rect 502 1650 503 1654
rect 507 1650 508 1654
rect 502 1649 508 1650
rect 694 1654 700 1655
rect 694 1650 695 1654
rect 699 1650 700 1654
rect 694 1649 700 1650
rect 886 1654 892 1655
rect 886 1650 887 1654
rect 891 1650 892 1654
rect 886 1649 892 1650
rect 1078 1654 1084 1655
rect 1078 1650 1079 1654
rect 1083 1650 1084 1654
rect 1078 1649 1084 1650
rect 1262 1654 1268 1655
rect 1262 1650 1263 1654
rect 1267 1650 1268 1654
rect 1262 1649 1268 1650
rect 1438 1654 1444 1655
rect 1438 1650 1439 1654
rect 1443 1650 1444 1654
rect 1438 1649 1444 1650
rect 1614 1654 1620 1655
rect 1614 1650 1615 1654
rect 1619 1650 1620 1654
rect 1614 1649 1620 1650
rect 1790 1654 1796 1655
rect 1790 1650 1791 1654
rect 1795 1650 1796 1654
rect 2032 1650 2034 1665
rect 2070 1664 2076 1665
rect 3990 1665 3991 1669
rect 3995 1665 3996 1669
rect 3990 1664 3996 1665
rect 2070 1652 2076 1653
rect 1790 1649 1796 1650
rect 2030 1649 2036 1650
rect 110 1645 111 1649
rect 115 1645 116 1649
rect 110 1644 116 1645
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2070 1648 2071 1652
rect 2075 1648 2076 1652
rect 2070 1647 2076 1648
rect 3990 1652 3996 1653
rect 3990 1648 3991 1652
rect 3995 1648 3996 1652
rect 3990 1647 3996 1648
rect 2030 1644 2036 1645
rect 110 1632 116 1633
rect 110 1628 111 1632
rect 115 1628 116 1632
rect 110 1627 116 1628
rect 2030 1632 2036 1633
rect 2030 1628 2031 1632
rect 2035 1628 2036 1632
rect 2030 1627 2036 1628
rect 112 1591 114 1627
rect 150 1613 156 1614
rect 150 1609 151 1613
rect 155 1609 156 1613
rect 150 1608 156 1609
rect 318 1613 324 1614
rect 318 1609 319 1613
rect 323 1609 324 1613
rect 318 1608 324 1609
rect 502 1613 508 1614
rect 502 1609 503 1613
rect 507 1609 508 1613
rect 502 1608 508 1609
rect 694 1613 700 1614
rect 694 1609 695 1613
rect 699 1609 700 1613
rect 694 1608 700 1609
rect 886 1613 892 1614
rect 886 1609 887 1613
rect 891 1609 892 1613
rect 886 1608 892 1609
rect 1078 1613 1084 1614
rect 1078 1609 1079 1613
rect 1083 1609 1084 1613
rect 1078 1608 1084 1609
rect 1262 1613 1268 1614
rect 1262 1609 1263 1613
rect 1267 1609 1268 1613
rect 1262 1608 1268 1609
rect 1438 1613 1444 1614
rect 1438 1609 1439 1613
rect 1443 1609 1444 1613
rect 1438 1608 1444 1609
rect 1614 1613 1620 1614
rect 1614 1609 1615 1613
rect 1619 1609 1620 1613
rect 1614 1608 1620 1609
rect 1790 1613 1796 1614
rect 1790 1609 1791 1613
rect 1795 1609 1796 1613
rect 1790 1608 1796 1609
rect 152 1591 154 1608
rect 320 1591 322 1608
rect 504 1591 506 1608
rect 696 1591 698 1608
rect 888 1591 890 1608
rect 1080 1591 1082 1608
rect 1264 1591 1266 1608
rect 1440 1591 1442 1608
rect 1616 1591 1618 1608
rect 1792 1591 1794 1608
rect 2032 1591 2034 1627
rect 2072 1607 2074 1647
rect 2110 1633 2116 1634
rect 2110 1629 2111 1633
rect 2115 1629 2116 1633
rect 2110 1628 2116 1629
rect 2310 1633 2316 1634
rect 2310 1629 2311 1633
rect 2315 1629 2316 1633
rect 2310 1628 2316 1629
rect 2526 1633 2532 1634
rect 2526 1629 2527 1633
rect 2531 1629 2532 1633
rect 2526 1628 2532 1629
rect 2742 1633 2748 1634
rect 2742 1629 2743 1633
rect 2747 1629 2748 1633
rect 2742 1628 2748 1629
rect 2950 1633 2956 1634
rect 2950 1629 2951 1633
rect 2955 1629 2956 1633
rect 2950 1628 2956 1629
rect 3150 1633 3156 1634
rect 3150 1629 3151 1633
rect 3155 1629 3156 1633
rect 3150 1628 3156 1629
rect 3342 1633 3348 1634
rect 3342 1629 3343 1633
rect 3347 1629 3348 1633
rect 3342 1628 3348 1629
rect 3526 1633 3532 1634
rect 3526 1629 3527 1633
rect 3531 1629 3532 1633
rect 3526 1628 3532 1629
rect 3718 1633 3724 1634
rect 3718 1629 3719 1633
rect 3723 1629 3724 1633
rect 3718 1628 3724 1629
rect 3894 1633 3900 1634
rect 3894 1629 3895 1633
rect 3899 1629 3900 1633
rect 3894 1628 3900 1629
rect 2112 1607 2114 1628
rect 2312 1607 2314 1628
rect 2528 1607 2530 1628
rect 2744 1607 2746 1628
rect 2952 1607 2954 1628
rect 3152 1607 3154 1628
rect 3344 1607 3346 1628
rect 3528 1607 3530 1628
rect 3720 1607 3722 1628
rect 3896 1607 3898 1628
rect 3992 1607 3994 1647
rect 2071 1606 2075 1607
rect 2071 1601 2075 1602
rect 2111 1606 2115 1607
rect 2111 1601 2115 1602
rect 2311 1606 2315 1607
rect 2311 1601 2315 1602
rect 2479 1606 2483 1607
rect 2479 1601 2483 1602
rect 2527 1606 2531 1607
rect 2527 1601 2531 1602
rect 2583 1606 2587 1607
rect 2583 1601 2587 1602
rect 2695 1606 2699 1607
rect 2695 1601 2699 1602
rect 2743 1606 2747 1607
rect 2743 1601 2747 1602
rect 2815 1606 2819 1607
rect 2815 1601 2819 1602
rect 2943 1606 2947 1607
rect 2943 1601 2947 1602
rect 2951 1606 2955 1607
rect 2951 1601 2955 1602
rect 3079 1606 3083 1607
rect 3079 1601 3083 1602
rect 3151 1606 3155 1607
rect 3151 1601 3155 1602
rect 3223 1606 3227 1607
rect 3223 1601 3227 1602
rect 3343 1606 3347 1607
rect 3343 1601 3347 1602
rect 3383 1606 3387 1607
rect 3383 1601 3387 1602
rect 3527 1606 3531 1607
rect 3527 1601 3531 1602
rect 3551 1606 3555 1607
rect 3551 1601 3555 1602
rect 3719 1606 3723 1607
rect 3719 1601 3723 1602
rect 3727 1606 3731 1607
rect 3727 1601 3731 1602
rect 3895 1606 3899 1607
rect 3895 1601 3899 1602
rect 3991 1606 3995 1607
rect 3991 1601 3995 1602
rect 111 1590 115 1591
rect 111 1585 115 1586
rect 151 1590 155 1591
rect 151 1585 155 1586
rect 319 1590 323 1591
rect 319 1585 323 1586
rect 455 1590 459 1591
rect 455 1585 459 1586
rect 503 1590 507 1591
rect 503 1585 507 1586
rect 599 1590 603 1591
rect 599 1585 603 1586
rect 695 1590 699 1591
rect 695 1585 699 1586
rect 743 1590 747 1591
rect 743 1585 747 1586
rect 887 1590 891 1591
rect 887 1585 891 1586
rect 1031 1590 1035 1591
rect 1031 1585 1035 1586
rect 1079 1590 1083 1591
rect 1079 1585 1083 1586
rect 1175 1590 1179 1591
rect 1175 1585 1179 1586
rect 1263 1590 1267 1591
rect 1263 1585 1267 1586
rect 1319 1590 1323 1591
rect 1319 1585 1323 1586
rect 1439 1590 1443 1591
rect 1439 1585 1443 1586
rect 1471 1590 1475 1591
rect 1471 1585 1475 1586
rect 1615 1590 1619 1591
rect 1615 1585 1619 1586
rect 1623 1590 1627 1591
rect 1623 1585 1627 1586
rect 1791 1590 1795 1591
rect 1791 1585 1795 1586
rect 2031 1590 2035 1591
rect 2031 1585 2035 1586
rect 112 1557 114 1585
rect 320 1576 322 1585
rect 456 1576 458 1585
rect 600 1576 602 1585
rect 744 1576 746 1585
rect 888 1576 890 1585
rect 1032 1576 1034 1585
rect 1176 1576 1178 1585
rect 1320 1576 1322 1585
rect 1472 1576 1474 1585
rect 1624 1576 1626 1585
rect 318 1575 324 1576
rect 318 1571 319 1575
rect 323 1571 324 1575
rect 318 1570 324 1571
rect 454 1575 460 1576
rect 454 1571 455 1575
rect 459 1571 460 1575
rect 454 1570 460 1571
rect 598 1575 604 1576
rect 598 1571 599 1575
rect 603 1571 604 1575
rect 598 1570 604 1571
rect 742 1575 748 1576
rect 742 1571 743 1575
rect 747 1571 748 1575
rect 742 1570 748 1571
rect 886 1575 892 1576
rect 886 1571 887 1575
rect 891 1571 892 1575
rect 886 1570 892 1571
rect 1030 1575 1036 1576
rect 1030 1571 1031 1575
rect 1035 1571 1036 1575
rect 1030 1570 1036 1571
rect 1174 1575 1180 1576
rect 1174 1571 1175 1575
rect 1179 1571 1180 1575
rect 1174 1570 1180 1571
rect 1318 1575 1324 1576
rect 1318 1571 1319 1575
rect 1323 1571 1324 1575
rect 1318 1570 1324 1571
rect 1470 1575 1476 1576
rect 1470 1571 1471 1575
rect 1475 1571 1476 1575
rect 1470 1570 1476 1571
rect 1622 1575 1628 1576
rect 1622 1571 1623 1575
rect 1627 1571 1628 1575
rect 1622 1570 1628 1571
rect 2032 1557 2034 1585
rect 2072 1573 2074 1601
rect 2480 1592 2482 1601
rect 2584 1592 2586 1601
rect 2696 1592 2698 1601
rect 2816 1592 2818 1601
rect 2944 1592 2946 1601
rect 3080 1592 3082 1601
rect 3224 1592 3226 1601
rect 3384 1592 3386 1601
rect 3552 1592 3554 1601
rect 3728 1592 3730 1601
rect 3896 1592 3898 1601
rect 2478 1591 2484 1592
rect 2478 1587 2479 1591
rect 2483 1587 2484 1591
rect 2478 1586 2484 1587
rect 2582 1591 2588 1592
rect 2582 1587 2583 1591
rect 2587 1587 2588 1591
rect 2582 1586 2588 1587
rect 2694 1591 2700 1592
rect 2694 1587 2695 1591
rect 2699 1587 2700 1591
rect 2694 1586 2700 1587
rect 2814 1591 2820 1592
rect 2814 1587 2815 1591
rect 2819 1587 2820 1591
rect 2814 1586 2820 1587
rect 2942 1591 2948 1592
rect 2942 1587 2943 1591
rect 2947 1587 2948 1591
rect 2942 1586 2948 1587
rect 3078 1591 3084 1592
rect 3078 1587 3079 1591
rect 3083 1587 3084 1591
rect 3078 1586 3084 1587
rect 3222 1591 3228 1592
rect 3222 1587 3223 1591
rect 3227 1587 3228 1591
rect 3222 1586 3228 1587
rect 3382 1591 3388 1592
rect 3382 1587 3383 1591
rect 3387 1587 3388 1591
rect 3382 1586 3388 1587
rect 3550 1591 3556 1592
rect 3550 1587 3551 1591
rect 3555 1587 3556 1591
rect 3550 1586 3556 1587
rect 3726 1591 3732 1592
rect 3726 1587 3727 1591
rect 3731 1587 3732 1591
rect 3726 1586 3732 1587
rect 3894 1591 3900 1592
rect 3894 1587 3895 1591
rect 3899 1587 3900 1591
rect 3894 1586 3900 1587
rect 3992 1573 3994 1601
rect 2070 1572 2076 1573
rect 2070 1568 2071 1572
rect 2075 1568 2076 1572
rect 2070 1567 2076 1568
rect 3990 1572 3996 1573
rect 3990 1568 3991 1572
rect 3995 1568 3996 1572
rect 3990 1567 3996 1568
rect 110 1556 116 1557
rect 110 1552 111 1556
rect 115 1552 116 1556
rect 110 1551 116 1552
rect 2030 1556 2036 1557
rect 2030 1552 2031 1556
rect 2035 1552 2036 1556
rect 2030 1551 2036 1552
rect 2070 1555 2076 1556
rect 2070 1551 2071 1555
rect 2075 1551 2076 1555
rect 3990 1555 3996 1556
rect 3990 1551 3991 1555
rect 3995 1551 3996 1555
rect 2070 1550 2076 1551
rect 2478 1550 2484 1551
rect 110 1539 116 1540
rect 110 1535 111 1539
rect 115 1535 116 1539
rect 2030 1539 2036 1540
rect 2030 1535 2031 1539
rect 2035 1535 2036 1539
rect 110 1534 116 1535
rect 318 1534 324 1535
rect 112 1511 114 1534
rect 318 1530 319 1534
rect 323 1530 324 1534
rect 318 1529 324 1530
rect 454 1534 460 1535
rect 454 1530 455 1534
rect 459 1530 460 1534
rect 454 1529 460 1530
rect 598 1534 604 1535
rect 598 1530 599 1534
rect 603 1530 604 1534
rect 598 1529 604 1530
rect 742 1534 748 1535
rect 742 1530 743 1534
rect 747 1530 748 1534
rect 742 1529 748 1530
rect 886 1534 892 1535
rect 886 1530 887 1534
rect 891 1530 892 1534
rect 886 1529 892 1530
rect 1030 1534 1036 1535
rect 1030 1530 1031 1534
rect 1035 1530 1036 1534
rect 1030 1529 1036 1530
rect 1174 1534 1180 1535
rect 1174 1530 1175 1534
rect 1179 1530 1180 1534
rect 1174 1529 1180 1530
rect 1318 1534 1324 1535
rect 1318 1530 1319 1534
rect 1323 1530 1324 1534
rect 1318 1529 1324 1530
rect 1470 1534 1476 1535
rect 1470 1530 1471 1534
rect 1475 1530 1476 1534
rect 1470 1529 1476 1530
rect 1622 1534 1628 1535
rect 2030 1534 2036 1535
rect 1622 1530 1623 1534
rect 1627 1530 1628 1534
rect 1622 1529 1628 1530
rect 320 1511 322 1529
rect 456 1511 458 1529
rect 600 1511 602 1529
rect 744 1511 746 1529
rect 888 1511 890 1529
rect 1032 1511 1034 1529
rect 1176 1511 1178 1529
rect 1320 1511 1322 1529
rect 1472 1511 1474 1529
rect 1624 1511 1626 1529
rect 2032 1511 2034 1534
rect 2072 1523 2074 1550
rect 2478 1546 2479 1550
rect 2483 1546 2484 1550
rect 2478 1545 2484 1546
rect 2582 1550 2588 1551
rect 2582 1546 2583 1550
rect 2587 1546 2588 1550
rect 2582 1545 2588 1546
rect 2694 1550 2700 1551
rect 2694 1546 2695 1550
rect 2699 1546 2700 1550
rect 2694 1545 2700 1546
rect 2814 1550 2820 1551
rect 2814 1546 2815 1550
rect 2819 1546 2820 1550
rect 2814 1545 2820 1546
rect 2942 1550 2948 1551
rect 2942 1546 2943 1550
rect 2947 1546 2948 1550
rect 2942 1545 2948 1546
rect 3078 1550 3084 1551
rect 3078 1546 3079 1550
rect 3083 1546 3084 1550
rect 3078 1545 3084 1546
rect 3222 1550 3228 1551
rect 3222 1546 3223 1550
rect 3227 1546 3228 1550
rect 3222 1545 3228 1546
rect 3382 1550 3388 1551
rect 3382 1546 3383 1550
rect 3387 1546 3388 1550
rect 3382 1545 3388 1546
rect 3550 1550 3556 1551
rect 3550 1546 3551 1550
rect 3555 1546 3556 1550
rect 3550 1545 3556 1546
rect 3726 1550 3732 1551
rect 3726 1546 3727 1550
rect 3731 1546 3732 1550
rect 3726 1545 3732 1546
rect 3894 1550 3900 1551
rect 3990 1550 3996 1551
rect 3894 1546 3895 1550
rect 3899 1546 3900 1550
rect 3894 1545 3900 1546
rect 2480 1523 2482 1545
rect 2584 1523 2586 1545
rect 2696 1523 2698 1545
rect 2816 1523 2818 1545
rect 2944 1523 2946 1545
rect 3080 1523 3082 1545
rect 3224 1523 3226 1545
rect 3384 1523 3386 1545
rect 3552 1523 3554 1545
rect 3728 1523 3730 1545
rect 3896 1523 3898 1545
rect 3992 1523 3994 1550
rect 2071 1522 2075 1523
rect 2071 1517 2075 1518
rect 2479 1522 2483 1523
rect 2479 1517 2483 1518
rect 2487 1522 2491 1523
rect 2487 1517 2491 1518
rect 2583 1522 2587 1523
rect 2583 1517 2587 1518
rect 2591 1522 2595 1523
rect 2591 1517 2595 1518
rect 2695 1522 2699 1523
rect 2695 1517 2699 1518
rect 2807 1522 2811 1523
rect 2807 1517 2811 1518
rect 2815 1522 2819 1523
rect 2815 1517 2819 1518
rect 2935 1522 2939 1523
rect 2935 1517 2939 1518
rect 2943 1522 2947 1523
rect 2943 1517 2947 1518
rect 3071 1522 3075 1523
rect 3071 1517 3075 1518
rect 3079 1522 3083 1523
rect 3079 1517 3083 1518
rect 3223 1522 3227 1523
rect 3223 1517 3227 1518
rect 3383 1522 3387 1523
rect 3383 1517 3387 1518
rect 3551 1522 3555 1523
rect 3551 1517 3555 1518
rect 3719 1522 3723 1523
rect 3719 1517 3723 1518
rect 3727 1522 3731 1523
rect 3727 1517 3731 1518
rect 3895 1522 3899 1523
rect 3895 1517 3899 1518
rect 3991 1522 3995 1523
rect 3991 1517 3995 1518
rect 111 1510 115 1511
rect 111 1505 115 1506
rect 319 1510 323 1511
rect 319 1505 323 1506
rect 359 1510 363 1511
rect 359 1505 363 1506
rect 455 1510 459 1511
rect 455 1505 459 1506
rect 487 1510 491 1511
rect 487 1505 491 1506
rect 599 1510 603 1511
rect 599 1505 603 1506
rect 623 1510 627 1511
rect 623 1505 627 1506
rect 743 1510 747 1511
rect 743 1505 747 1506
rect 775 1510 779 1511
rect 775 1505 779 1506
rect 887 1510 891 1511
rect 887 1505 891 1506
rect 927 1510 931 1511
rect 927 1505 931 1506
rect 1031 1510 1035 1511
rect 1031 1505 1035 1506
rect 1087 1510 1091 1511
rect 1087 1505 1091 1506
rect 1175 1510 1179 1511
rect 1175 1505 1179 1506
rect 1255 1510 1259 1511
rect 1255 1505 1259 1506
rect 1319 1510 1323 1511
rect 1319 1505 1323 1506
rect 1423 1510 1427 1511
rect 1423 1505 1427 1506
rect 1471 1510 1475 1511
rect 1471 1505 1475 1506
rect 1591 1510 1595 1511
rect 1591 1505 1595 1506
rect 1623 1510 1627 1511
rect 1623 1505 1627 1506
rect 1767 1510 1771 1511
rect 1767 1505 1771 1506
rect 2031 1510 2035 1511
rect 2031 1505 2035 1506
rect 112 1490 114 1505
rect 360 1495 362 1505
rect 488 1495 490 1505
rect 624 1495 626 1505
rect 776 1495 778 1505
rect 928 1495 930 1505
rect 1088 1495 1090 1505
rect 1256 1495 1258 1505
rect 1424 1495 1426 1505
rect 1592 1495 1594 1505
rect 1768 1495 1770 1505
rect 358 1494 364 1495
rect 358 1490 359 1494
rect 363 1490 364 1494
rect 110 1489 116 1490
rect 358 1489 364 1490
rect 486 1494 492 1495
rect 486 1490 487 1494
rect 491 1490 492 1494
rect 486 1489 492 1490
rect 622 1494 628 1495
rect 622 1490 623 1494
rect 627 1490 628 1494
rect 622 1489 628 1490
rect 774 1494 780 1495
rect 774 1490 775 1494
rect 779 1490 780 1494
rect 774 1489 780 1490
rect 926 1494 932 1495
rect 926 1490 927 1494
rect 931 1490 932 1494
rect 926 1489 932 1490
rect 1086 1494 1092 1495
rect 1086 1490 1087 1494
rect 1091 1490 1092 1494
rect 1086 1489 1092 1490
rect 1254 1494 1260 1495
rect 1254 1490 1255 1494
rect 1259 1490 1260 1494
rect 1254 1489 1260 1490
rect 1422 1494 1428 1495
rect 1422 1490 1423 1494
rect 1427 1490 1428 1494
rect 1422 1489 1428 1490
rect 1590 1494 1596 1495
rect 1590 1490 1591 1494
rect 1595 1490 1596 1494
rect 1590 1489 1596 1490
rect 1766 1494 1772 1495
rect 1766 1490 1767 1494
rect 1771 1490 1772 1494
rect 2032 1490 2034 1505
rect 2072 1502 2074 1517
rect 2488 1507 2490 1517
rect 2592 1507 2594 1517
rect 2696 1507 2698 1517
rect 2808 1507 2810 1517
rect 2936 1507 2938 1517
rect 3072 1507 3074 1517
rect 3224 1507 3226 1517
rect 3384 1507 3386 1517
rect 3552 1507 3554 1517
rect 3720 1507 3722 1517
rect 3896 1507 3898 1517
rect 2486 1506 2492 1507
rect 2486 1502 2487 1506
rect 2491 1502 2492 1506
rect 2070 1501 2076 1502
rect 2486 1501 2492 1502
rect 2590 1506 2596 1507
rect 2590 1502 2591 1506
rect 2595 1502 2596 1506
rect 2590 1501 2596 1502
rect 2694 1506 2700 1507
rect 2694 1502 2695 1506
rect 2699 1502 2700 1506
rect 2694 1501 2700 1502
rect 2806 1506 2812 1507
rect 2806 1502 2807 1506
rect 2811 1502 2812 1506
rect 2806 1501 2812 1502
rect 2934 1506 2940 1507
rect 2934 1502 2935 1506
rect 2939 1502 2940 1506
rect 2934 1501 2940 1502
rect 3070 1506 3076 1507
rect 3070 1502 3071 1506
rect 3075 1502 3076 1506
rect 3070 1501 3076 1502
rect 3222 1506 3228 1507
rect 3222 1502 3223 1506
rect 3227 1502 3228 1506
rect 3222 1501 3228 1502
rect 3382 1506 3388 1507
rect 3382 1502 3383 1506
rect 3387 1502 3388 1506
rect 3382 1501 3388 1502
rect 3550 1506 3556 1507
rect 3550 1502 3551 1506
rect 3555 1502 3556 1506
rect 3550 1501 3556 1502
rect 3718 1506 3724 1507
rect 3718 1502 3719 1506
rect 3723 1502 3724 1506
rect 3718 1501 3724 1502
rect 3894 1506 3900 1507
rect 3894 1502 3895 1506
rect 3899 1502 3900 1506
rect 3992 1502 3994 1517
rect 3894 1501 3900 1502
rect 3990 1501 3996 1502
rect 2070 1497 2071 1501
rect 2075 1497 2076 1501
rect 2070 1496 2076 1497
rect 3990 1497 3991 1501
rect 3995 1497 3996 1501
rect 3990 1496 3996 1497
rect 1766 1489 1772 1490
rect 2030 1489 2036 1490
rect 110 1485 111 1489
rect 115 1485 116 1489
rect 110 1484 116 1485
rect 2030 1485 2031 1489
rect 2035 1485 2036 1489
rect 2030 1484 2036 1485
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 3990 1484 3996 1485
rect 3990 1480 3991 1484
rect 3995 1480 3996 1484
rect 3990 1479 3996 1480
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 110 1467 116 1468
rect 2030 1472 2036 1473
rect 2030 1468 2031 1472
rect 2035 1468 2036 1472
rect 2030 1467 2036 1468
rect 112 1431 114 1467
rect 358 1453 364 1454
rect 358 1449 359 1453
rect 363 1449 364 1453
rect 358 1448 364 1449
rect 486 1453 492 1454
rect 486 1449 487 1453
rect 491 1449 492 1453
rect 486 1448 492 1449
rect 622 1453 628 1454
rect 622 1449 623 1453
rect 627 1449 628 1453
rect 622 1448 628 1449
rect 774 1453 780 1454
rect 774 1449 775 1453
rect 779 1449 780 1453
rect 774 1448 780 1449
rect 926 1453 932 1454
rect 926 1449 927 1453
rect 931 1449 932 1453
rect 926 1448 932 1449
rect 1086 1453 1092 1454
rect 1086 1449 1087 1453
rect 1091 1449 1092 1453
rect 1086 1448 1092 1449
rect 1254 1453 1260 1454
rect 1254 1449 1255 1453
rect 1259 1449 1260 1453
rect 1254 1448 1260 1449
rect 1422 1453 1428 1454
rect 1422 1449 1423 1453
rect 1427 1449 1428 1453
rect 1422 1448 1428 1449
rect 1590 1453 1596 1454
rect 1590 1449 1591 1453
rect 1595 1449 1596 1453
rect 1590 1448 1596 1449
rect 1766 1453 1772 1454
rect 1766 1449 1767 1453
rect 1771 1449 1772 1453
rect 1766 1448 1772 1449
rect 360 1431 362 1448
rect 488 1431 490 1448
rect 624 1431 626 1448
rect 776 1431 778 1448
rect 928 1431 930 1448
rect 1088 1431 1090 1448
rect 1256 1431 1258 1448
rect 1424 1431 1426 1448
rect 1592 1431 1594 1448
rect 1768 1431 1770 1448
rect 2032 1431 2034 1467
rect 2072 1447 2074 1479
rect 2486 1465 2492 1466
rect 2486 1461 2487 1465
rect 2491 1461 2492 1465
rect 2486 1460 2492 1461
rect 2590 1465 2596 1466
rect 2590 1461 2591 1465
rect 2595 1461 2596 1465
rect 2590 1460 2596 1461
rect 2694 1465 2700 1466
rect 2694 1461 2695 1465
rect 2699 1461 2700 1465
rect 2694 1460 2700 1461
rect 2806 1465 2812 1466
rect 2806 1461 2807 1465
rect 2811 1461 2812 1465
rect 2806 1460 2812 1461
rect 2934 1465 2940 1466
rect 2934 1461 2935 1465
rect 2939 1461 2940 1465
rect 2934 1460 2940 1461
rect 3070 1465 3076 1466
rect 3070 1461 3071 1465
rect 3075 1461 3076 1465
rect 3070 1460 3076 1461
rect 3222 1465 3228 1466
rect 3222 1461 3223 1465
rect 3227 1461 3228 1465
rect 3222 1460 3228 1461
rect 3382 1465 3388 1466
rect 3382 1461 3383 1465
rect 3387 1461 3388 1465
rect 3382 1460 3388 1461
rect 3550 1465 3556 1466
rect 3550 1461 3551 1465
rect 3555 1461 3556 1465
rect 3550 1460 3556 1461
rect 3718 1465 3724 1466
rect 3718 1461 3719 1465
rect 3723 1461 3724 1465
rect 3718 1460 3724 1461
rect 3894 1465 3900 1466
rect 3894 1461 3895 1465
rect 3899 1461 3900 1465
rect 3894 1460 3900 1461
rect 2488 1447 2490 1460
rect 2592 1447 2594 1460
rect 2696 1447 2698 1460
rect 2808 1447 2810 1460
rect 2936 1447 2938 1460
rect 3072 1447 3074 1460
rect 3224 1447 3226 1460
rect 3384 1447 3386 1460
rect 3552 1447 3554 1460
rect 3720 1447 3722 1460
rect 3896 1447 3898 1460
rect 3992 1447 3994 1479
rect 2071 1446 2075 1447
rect 2071 1441 2075 1442
rect 2239 1446 2243 1447
rect 2239 1441 2243 1442
rect 2351 1446 2355 1447
rect 2351 1441 2355 1442
rect 2471 1446 2475 1447
rect 2471 1441 2475 1442
rect 2487 1446 2491 1447
rect 2487 1441 2491 1442
rect 2591 1446 2595 1447
rect 2591 1441 2595 1442
rect 2695 1446 2699 1447
rect 2695 1441 2699 1442
rect 2727 1446 2731 1447
rect 2727 1441 2731 1442
rect 2807 1446 2811 1447
rect 2807 1441 2811 1442
rect 2879 1446 2883 1447
rect 2879 1441 2883 1442
rect 2935 1446 2939 1447
rect 2935 1441 2939 1442
rect 3055 1446 3059 1447
rect 3055 1441 3059 1442
rect 3071 1446 3075 1447
rect 3071 1441 3075 1442
rect 3223 1446 3227 1447
rect 3223 1441 3227 1442
rect 3247 1446 3251 1447
rect 3247 1441 3251 1442
rect 3383 1446 3387 1447
rect 3383 1441 3387 1442
rect 3455 1446 3459 1447
rect 3455 1441 3459 1442
rect 3551 1446 3555 1447
rect 3551 1441 3555 1442
rect 3671 1446 3675 1447
rect 3671 1441 3675 1442
rect 3719 1446 3723 1447
rect 3719 1441 3723 1442
rect 3887 1446 3891 1447
rect 3887 1441 3891 1442
rect 3895 1446 3899 1447
rect 3895 1441 3899 1442
rect 3991 1446 3995 1447
rect 3991 1441 3995 1442
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 151 1430 155 1431
rect 151 1425 155 1426
rect 271 1430 275 1431
rect 271 1425 275 1426
rect 359 1430 363 1431
rect 359 1425 363 1426
rect 431 1430 435 1431
rect 431 1425 435 1426
rect 487 1430 491 1431
rect 487 1425 491 1426
rect 615 1430 619 1431
rect 615 1425 619 1426
rect 623 1430 627 1431
rect 623 1425 627 1426
rect 775 1430 779 1431
rect 775 1425 779 1426
rect 807 1430 811 1431
rect 807 1425 811 1426
rect 927 1430 931 1431
rect 927 1425 931 1426
rect 1007 1430 1011 1431
rect 1007 1425 1011 1426
rect 1087 1430 1091 1431
rect 1087 1425 1091 1426
rect 1215 1430 1219 1431
rect 1215 1425 1219 1426
rect 1255 1430 1259 1431
rect 1255 1425 1259 1426
rect 1423 1430 1427 1431
rect 1423 1425 1427 1426
rect 1591 1430 1595 1431
rect 1591 1425 1595 1426
rect 1631 1430 1635 1431
rect 1631 1425 1635 1426
rect 1767 1430 1771 1431
rect 1767 1425 1771 1426
rect 1847 1430 1851 1431
rect 1847 1425 1851 1426
rect 2031 1430 2035 1431
rect 2031 1425 2035 1426
rect 112 1397 114 1425
rect 152 1416 154 1425
rect 272 1416 274 1425
rect 432 1416 434 1425
rect 616 1416 618 1425
rect 808 1416 810 1425
rect 1008 1416 1010 1425
rect 1216 1416 1218 1425
rect 1424 1416 1426 1425
rect 1632 1416 1634 1425
rect 1848 1416 1850 1425
rect 150 1415 156 1416
rect 150 1411 151 1415
rect 155 1411 156 1415
rect 150 1410 156 1411
rect 270 1415 276 1416
rect 270 1411 271 1415
rect 275 1411 276 1415
rect 270 1410 276 1411
rect 430 1415 436 1416
rect 430 1411 431 1415
rect 435 1411 436 1415
rect 430 1410 436 1411
rect 614 1415 620 1416
rect 614 1411 615 1415
rect 619 1411 620 1415
rect 614 1410 620 1411
rect 806 1415 812 1416
rect 806 1411 807 1415
rect 811 1411 812 1415
rect 806 1410 812 1411
rect 1006 1415 1012 1416
rect 1006 1411 1007 1415
rect 1011 1411 1012 1415
rect 1006 1410 1012 1411
rect 1214 1415 1220 1416
rect 1214 1411 1215 1415
rect 1219 1411 1220 1415
rect 1214 1410 1220 1411
rect 1422 1415 1428 1416
rect 1422 1411 1423 1415
rect 1427 1411 1428 1415
rect 1422 1410 1428 1411
rect 1630 1415 1636 1416
rect 1630 1411 1631 1415
rect 1635 1411 1636 1415
rect 1630 1410 1636 1411
rect 1846 1415 1852 1416
rect 1846 1411 1847 1415
rect 1851 1411 1852 1415
rect 1846 1410 1852 1411
rect 2032 1397 2034 1425
rect 2072 1413 2074 1441
rect 2240 1432 2242 1441
rect 2352 1432 2354 1441
rect 2472 1432 2474 1441
rect 2592 1432 2594 1441
rect 2728 1432 2730 1441
rect 2880 1432 2882 1441
rect 3056 1432 3058 1441
rect 3248 1432 3250 1441
rect 3456 1432 3458 1441
rect 3672 1432 3674 1441
rect 3888 1432 3890 1441
rect 2238 1431 2244 1432
rect 2238 1427 2239 1431
rect 2243 1427 2244 1431
rect 2238 1426 2244 1427
rect 2350 1431 2356 1432
rect 2350 1427 2351 1431
rect 2355 1427 2356 1431
rect 2350 1426 2356 1427
rect 2470 1431 2476 1432
rect 2470 1427 2471 1431
rect 2475 1427 2476 1431
rect 2470 1426 2476 1427
rect 2590 1431 2596 1432
rect 2590 1427 2591 1431
rect 2595 1427 2596 1431
rect 2590 1426 2596 1427
rect 2726 1431 2732 1432
rect 2726 1427 2727 1431
rect 2731 1427 2732 1431
rect 2726 1426 2732 1427
rect 2878 1431 2884 1432
rect 2878 1427 2879 1431
rect 2883 1427 2884 1431
rect 2878 1426 2884 1427
rect 3054 1431 3060 1432
rect 3054 1427 3055 1431
rect 3059 1427 3060 1431
rect 3054 1426 3060 1427
rect 3246 1431 3252 1432
rect 3246 1427 3247 1431
rect 3251 1427 3252 1431
rect 3246 1426 3252 1427
rect 3454 1431 3460 1432
rect 3454 1427 3455 1431
rect 3459 1427 3460 1431
rect 3454 1426 3460 1427
rect 3670 1431 3676 1432
rect 3670 1427 3671 1431
rect 3675 1427 3676 1431
rect 3670 1426 3676 1427
rect 3886 1431 3892 1432
rect 3886 1427 3887 1431
rect 3891 1427 3892 1431
rect 3886 1426 3892 1427
rect 3992 1413 3994 1441
rect 2070 1412 2076 1413
rect 2070 1408 2071 1412
rect 2075 1408 2076 1412
rect 2070 1407 2076 1408
rect 3990 1412 3996 1413
rect 3990 1408 3991 1412
rect 3995 1408 3996 1412
rect 3990 1407 3996 1408
rect 110 1396 116 1397
rect 110 1392 111 1396
rect 115 1392 116 1396
rect 110 1391 116 1392
rect 2030 1396 2036 1397
rect 2030 1392 2031 1396
rect 2035 1392 2036 1396
rect 2030 1391 2036 1392
rect 2070 1395 2076 1396
rect 2070 1391 2071 1395
rect 2075 1391 2076 1395
rect 3990 1395 3996 1396
rect 3990 1391 3991 1395
rect 3995 1391 3996 1395
rect 2070 1390 2076 1391
rect 2238 1390 2244 1391
rect 110 1379 116 1380
rect 110 1375 111 1379
rect 115 1375 116 1379
rect 2030 1379 2036 1380
rect 2030 1375 2031 1379
rect 2035 1375 2036 1379
rect 110 1374 116 1375
rect 150 1374 156 1375
rect 112 1347 114 1374
rect 150 1370 151 1374
rect 155 1370 156 1374
rect 150 1369 156 1370
rect 270 1374 276 1375
rect 270 1370 271 1374
rect 275 1370 276 1374
rect 270 1369 276 1370
rect 430 1374 436 1375
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 614 1374 620 1375
rect 614 1370 615 1374
rect 619 1370 620 1374
rect 614 1369 620 1370
rect 806 1374 812 1375
rect 806 1370 807 1374
rect 811 1370 812 1374
rect 806 1369 812 1370
rect 1006 1374 1012 1375
rect 1006 1370 1007 1374
rect 1011 1370 1012 1374
rect 1006 1369 1012 1370
rect 1214 1374 1220 1375
rect 1214 1370 1215 1374
rect 1219 1370 1220 1374
rect 1214 1369 1220 1370
rect 1422 1374 1428 1375
rect 1422 1370 1423 1374
rect 1427 1370 1428 1374
rect 1422 1369 1428 1370
rect 1630 1374 1636 1375
rect 1630 1370 1631 1374
rect 1635 1370 1636 1374
rect 1630 1369 1636 1370
rect 1846 1374 1852 1375
rect 2030 1374 2036 1375
rect 1846 1370 1847 1374
rect 1851 1370 1852 1374
rect 1846 1369 1852 1370
rect 152 1347 154 1369
rect 272 1347 274 1369
rect 432 1347 434 1369
rect 616 1347 618 1369
rect 808 1347 810 1369
rect 1008 1347 1010 1369
rect 1216 1347 1218 1369
rect 1424 1347 1426 1369
rect 1632 1347 1634 1369
rect 1848 1347 1850 1369
rect 2032 1347 2034 1374
rect 2072 1367 2074 1390
rect 2238 1386 2239 1390
rect 2243 1386 2244 1390
rect 2238 1385 2244 1386
rect 2350 1390 2356 1391
rect 2350 1386 2351 1390
rect 2355 1386 2356 1390
rect 2350 1385 2356 1386
rect 2470 1390 2476 1391
rect 2470 1386 2471 1390
rect 2475 1386 2476 1390
rect 2470 1385 2476 1386
rect 2590 1390 2596 1391
rect 2590 1386 2591 1390
rect 2595 1386 2596 1390
rect 2590 1385 2596 1386
rect 2726 1390 2732 1391
rect 2726 1386 2727 1390
rect 2731 1386 2732 1390
rect 2726 1385 2732 1386
rect 2878 1390 2884 1391
rect 2878 1386 2879 1390
rect 2883 1386 2884 1390
rect 2878 1385 2884 1386
rect 3054 1390 3060 1391
rect 3054 1386 3055 1390
rect 3059 1386 3060 1390
rect 3054 1385 3060 1386
rect 3246 1390 3252 1391
rect 3246 1386 3247 1390
rect 3251 1386 3252 1390
rect 3246 1385 3252 1386
rect 3454 1390 3460 1391
rect 3454 1386 3455 1390
rect 3459 1386 3460 1390
rect 3454 1385 3460 1386
rect 3670 1390 3676 1391
rect 3670 1386 3671 1390
rect 3675 1386 3676 1390
rect 3670 1385 3676 1386
rect 3886 1390 3892 1391
rect 3990 1390 3996 1391
rect 3886 1386 3887 1390
rect 3891 1386 3892 1390
rect 3886 1385 3892 1386
rect 2240 1367 2242 1385
rect 2352 1367 2354 1385
rect 2472 1367 2474 1385
rect 2592 1367 2594 1385
rect 2728 1367 2730 1385
rect 2880 1367 2882 1385
rect 3056 1367 3058 1385
rect 3248 1367 3250 1385
rect 3456 1367 3458 1385
rect 3672 1367 3674 1385
rect 3888 1367 3890 1385
rect 3992 1367 3994 1390
rect 2071 1366 2075 1367
rect 2071 1361 2075 1362
rect 2239 1366 2243 1367
rect 2239 1361 2243 1362
rect 2351 1366 2355 1367
rect 2351 1361 2355 1362
rect 2391 1366 2395 1367
rect 2391 1361 2395 1362
rect 2471 1366 2475 1367
rect 2471 1361 2475 1362
rect 2527 1366 2531 1367
rect 2527 1361 2531 1362
rect 2591 1366 2595 1367
rect 2591 1361 2595 1362
rect 2679 1366 2683 1367
rect 2679 1361 2683 1362
rect 2727 1366 2731 1367
rect 2727 1361 2731 1362
rect 2839 1366 2843 1367
rect 2839 1361 2843 1362
rect 2879 1366 2883 1367
rect 2879 1361 2883 1362
rect 2999 1366 3003 1367
rect 2999 1361 3003 1362
rect 3055 1366 3059 1367
rect 3055 1361 3059 1362
rect 3167 1366 3171 1367
rect 3167 1361 3171 1362
rect 3247 1366 3251 1367
rect 3247 1361 3251 1362
rect 3343 1366 3347 1367
rect 3343 1361 3347 1362
rect 3455 1366 3459 1367
rect 3455 1361 3459 1362
rect 3519 1366 3523 1367
rect 3519 1361 3523 1362
rect 3671 1366 3675 1367
rect 3671 1361 3675 1362
rect 3695 1366 3699 1367
rect 3695 1361 3699 1362
rect 3879 1366 3883 1367
rect 3879 1361 3883 1362
rect 3887 1366 3891 1367
rect 3887 1361 3891 1362
rect 3991 1366 3995 1367
rect 3991 1361 3995 1362
rect 111 1346 115 1347
rect 111 1341 115 1342
rect 151 1346 155 1347
rect 151 1341 155 1342
rect 271 1346 275 1347
rect 271 1341 275 1342
rect 287 1346 291 1347
rect 287 1341 291 1342
rect 431 1346 435 1347
rect 431 1341 435 1342
rect 463 1346 467 1347
rect 463 1341 467 1342
rect 615 1346 619 1347
rect 615 1341 619 1342
rect 663 1346 667 1347
rect 663 1341 667 1342
rect 807 1346 811 1347
rect 807 1341 811 1342
rect 863 1346 867 1347
rect 863 1341 867 1342
rect 1007 1346 1011 1347
rect 1007 1341 1011 1342
rect 1063 1346 1067 1347
rect 1063 1341 1067 1342
rect 1215 1346 1219 1347
rect 1215 1341 1219 1342
rect 1255 1346 1259 1347
rect 1255 1341 1259 1342
rect 1423 1346 1427 1347
rect 1423 1341 1427 1342
rect 1431 1346 1435 1347
rect 1431 1341 1435 1342
rect 1607 1346 1611 1347
rect 1607 1341 1611 1342
rect 1631 1346 1635 1347
rect 1631 1341 1635 1342
rect 1783 1346 1787 1347
rect 1783 1341 1787 1342
rect 1847 1346 1851 1347
rect 1847 1341 1851 1342
rect 1935 1346 1939 1347
rect 1935 1341 1939 1342
rect 2031 1346 2035 1347
rect 2072 1346 2074 1361
rect 2392 1351 2394 1361
rect 2528 1351 2530 1361
rect 2680 1351 2682 1361
rect 2840 1351 2842 1361
rect 3000 1351 3002 1361
rect 3168 1351 3170 1361
rect 3344 1351 3346 1361
rect 3520 1351 3522 1361
rect 3696 1351 3698 1361
rect 3880 1351 3882 1361
rect 2390 1350 2396 1351
rect 2390 1346 2391 1350
rect 2395 1346 2396 1350
rect 2031 1341 2035 1342
rect 2070 1345 2076 1346
rect 2390 1345 2396 1346
rect 2526 1350 2532 1351
rect 2526 1346 2527 1350
rect 2531 1346 2532 1350
rect 2526 1345 2532 1346
rect 2678 1350 2684 1351
rect 2678 1346 2679 1350
rect 2683 1346 2684 1350
rect 2678 1345 2684 1346
rect 2838 1350 2844 1351
rect 2838 1346 2839 1350
rect 2843 1346 2844 1350
rect 2838 1345 2844 1346
rect 2998 1350 3004 1351
rect 2998 1346 2999 1350
rect 3003 1346 3004 1350
rect 2998 1345 3004 1346
rect 3166 1350 3172 1351
rect 3166 1346 3167 1350
rect 3171 1346 3172 1350
rect 3166 1345 3172 1346
rect 3342 1350 3348 1351
rect 3342 1346 3343 1350
rect 3347 1346 3348 1350
rect 3342 1345 3348 1346
rect 3518 1350 3524 1351
rect 3518 1346 3519 1350
rect 3523 1346 3524 1350
rect 3518 1345 3524 1346
rect 3694 1350 3700 1351
rect 3694 1346 3695 1350
rect 3699 1346 3700 1350
rect 3694 1345 3700 1346
rect 3878 1350 3884 1351
rect 3878 1346 3879 1350
rect 3883 1346 3884 1350
rect 3992 1346 3994 1361
rect 3878 1345 3884 1346
rect 3990 1345 3996 1346
rect 2070 1341 2071 1345
rect 2075 1341 2076 1345
rect 112 1326 114 1341
rect 152 1331 154 1341
rect 288 1331 290 1341
rect 464 1331 466 1341
rect 664 1331 666 1341
rect 864 1331 866 1341
rect 1064 1331 1066 1341
rect 1256 1331 1258 1341
rect 1432 1331 1434 1341
rect 1608 1331 1610 1341
rect 1784 1331 1786 1341
rect 1936 1331 1938 1341
rect 150 1330 156 1331
rect 150 1326 151 1330
rect 155 1326 156 1330
rect 110 1325 116 1326
rect 150 1325 156 1326
rect 286 1330 292 1331
rect 286 1326 287 1330
rect 291 1326 292 1330
rect 286 1325 292 1326
rect 462 1330 468 1331
rect 462 1326 463 1330
rect 467 1326 468 1330
rect 462 1325 468 1326
rect 662 1330 668 1331
rect 662 1326 663 1330
rect 667 1326 668 1330
rect 662 1325 668 1326
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 862 1325 868 1326
rect 1062 1330 1068 1331
rect 1062 1326 1063 1330
rect 1067 1326 1068 1330
rect 1062 1325 1068 1326
rect 1254 1330 1260 1331
rect 1254 1326 1255 1330
rect 1259 1326 1260 1330
rect 1254 1325 1260 1326
rect 1430 1330 1436 1331
rect 1430 1326 1431 1330
rect 1435 1326 1436 1330
rect 1430 1325 1436 1326
rect 1606 1330 1612 1331
rect 1606 1326 1607 1330
rect 1611 1326 1612 1330
rect 1606 1325 1612 1326
rect 1782 1330 1788 1331
rect 1782 1326 1783 1330
rect 1787 1326 1788 1330
rect 1782 1325 1788 1326
rect 1934 1330 1940 1331
rect 1934 1326 1935 1330
rect 1939 1326 1940 1330
rect 2032 1326 2034 1341
rect 2070 1340 2076 1341
rect 3990 1341 3991 1345
rect 3995 1341 3996 1345
rect 3990 1340 3996 1341
rect 2070 1328 2076 1329
rect 1934 1325 1940 1326
rect 2030 1325 2036 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 110 1320 116 1321
rect 2030 1321 2031 1325
rect 2035 1321 2036 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 3990 1328 3996 1329
rect 3990 1324 3991 1328
rect 3995 1324 3996 1328
rect 3990 1323 3996 1324
rect 2030 1320 2036 1321
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 110 1303 116 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2030 1303 2036 1304
rect 112 1275 114 1303
rect 150 1289 156 1290
rect 150 1285 151 1289
rect 155 1285 156 1289
rect 150 1284 156 1285
rect 286 1289 292 1290
rect 286 1285 287 1289
rect 291 1285 292 1289
rect 286 1284 292 1285
rect 462 1289 468 1290
rect 462 1285 463 1289
rect 467 1285 468 1289
rect 462 1284 468 1285
rect 662 1289 668 1290
rect 662 1285 663 1289
rect 667 1285 668 1289
rect 662 1284 668 1285
rect 862 1289 868 1290
rect 862 1285 863 1289
rect 867 1285 868 1289
rect 862 1284 868 1285
rect 1062 1289 1068 1290
rect 1062 1285 1063 1289
rect 1067 1285 1068 1289
rect 1062 1284 1068 1285
rect 1254 1289 1260 1290
rect 1254 1285 1255 1289
rect 1259 1285 1260 1289
rect 1254 1284 1260 1285
rect 1430 1289 1436 1290
rect 1430 1285 1431 1289
rect 1435 1285 1436 1289
rect 1430 1284 1436 1285
rect 1606 1289 1612 1290
rect 1606 1285 1607 1289
rect 1611 1285 1612 1289
rect 1606 1284 1612 1285
rect 1782 1289 1788 1290
rect 1782 1285 1783 1289
rect 1787 1285 1788 1289
rect 1782 1284 1788 1285
rect 1934 1289 1940 1290
rect 1934 1285 1935 1289
rect 1939 1285 1940 1289
rect 1934 1284 1940 1285
rect 152 1275 154 1284
rect 288 1275 290 1284
rect 464 1275 466 1284
rect 664 1275 666 1284
rect 864 1275 866 1284
rect 1064 1275 1066 1284
rect 1256 1275 1258 1284
rect 1432 1275 1434 1284
rect 1608 1275 1610 1284
rect 1784 1275 1786 1284
rect 1936 1275 1938 1284
rect 2032 1275 2034 1303
rect 2072 1287 2074 1323
rect 2390 1309 2396 1310
rect 2390 1305 2391 1309
rect 2395 1305 2396 1309
rect 2390 1304 2396 1305
rect 2526 1309 2532 1310
rect 2526 1305 2527 1309
rect 2531 1305 2532 1309
rect 2526 1304 2532 1305
rect 2678 1309 2684 1310
rect 2678 1305 2679 1309
rect 2683 1305 2684 1309
rect 2678 1304 2684 1305
rect 2838 1309 2844 1310
rect 2838 1305 2839 1309
rect 2843 1305 2844 1309
rect 2838 1304 2844 1305
rect 2998 1309 3004 1310
rect 2998 1305 2999 1309
rect 3003 1305 3004 1309
rect 2998 1304 3004 1305
rect 3166 1309 3172 1310
rect 3166 1305 3167 1309
rect 3171 1305 3172 1309
rect 3166 1304 3172 1305
rect 3342 1309 3348 1310
rect 3342 1305 3343 1309
rect 3347 1305 3348 1309
rect 3342 1304 3348 1305
rect 3518 1309 3524 1310
rect 3518 1305 3519 1309
rect 3523 1305 3524 1309
rect 3518 1304 3524 1305
rect 3694 1309 3700 1310
rect 3694 1305 3695 1309
rect 3699 1305 3700 1309
rect 3694 1304 3700 1305
rect 3878 1309 3884 1310
rect 3878 1305 3879 1309
rect 3883 1305 3884 1309
rect 3878 1304 3884 1305
rect 2392 1287 2394 1304
rect 2528 1287 2530 1304
rect 2680 1287 2682 1304
rect 2840 1287 2842 1304
rect 3000 1287 3002 1304
rect 3168 1287 3170 1304
rect 3344 1287 3346 1304
rect 3520 1287 3522 1304
rect 3696 1287 3698 1304
rect 3880 1287 3882 1304
rect 3992 1287 3994 1323
rect 2071 1286 2075 1287
rect 2071 1281 2075 1282
rect 2111 1286 2115 1287
rect 2111 1281 2115 1282
rect 2343 1286 2347 1287
rect 2343 1281 2347 1282
rect 2391 1286 2395 1287
rect 2391 1281 2395 1282
rect 2527 1286 2531 1287
rect 2527 1281 2531 1282
rect 2583 1286 2587 1287
rect 2583 1281 2587 1282
rect 2679 1286 2683 1287
rect 2679 1281 2683 1282
rect 2799 1286 2803 1287
rect 2799 1281 2803 1282
rect 2839 1286 2843 1287
rect 2839 1281 2843 1282
rect 2999 1286 3003 1287
rect 2999 1281 3003 1282
rect 3167 1286 3171 1287
rect 3167 1281 3171 1282
rect 3183 1286 3187 1287
rect 3183 1281 3187 1282
rect 3343 1286 3347 1287
rect 3343 1281 3347 1282
rect 3495 1286 3499 1287
rect 3495 1281 3499 1282
rect 3519 1286 3523 1287
rect 3519 1281 3523 1282
rect 3639 1286 3643 1287
rect 3639 1281 3643 1282
rect 3695 1286 3699 1287
rect 3695 1281 3699 1282
rect 3775 1286 3779 1287
rect 3775 1281 3779 1282
rect 3879 1286 3883 1287
rect 3879 1281 3883 1282
rect 3895 1286 3899 1287
rect 3895 1281 3899 1282
rect 3991 1286 3995 1287
rect 3991 1281 3995 1282
rect 111 1274 115 1275
rect 111 1269 115 1270
rect 151 1274 155 1275
rect 151 1269 155 1270
rect 207 1274 211 1275
rect 207 1269 211 1270
rect 287 1274 291 1275
rect 287 1269 291 1270
rect 327 1274 331 1275
rect 327 1269 331 1270
rect 455 1274 459 1275
rect 455 1269 459 1270
rect 463 1274 467 1275
rect 463 1269 467 1270
rect 583 1274 587 1275
rect 583 1269 587 1270
rect 663 1274 667 1275
rect 663 1269 667 1270
rect 719 1274 723 1275
rect 719 1269 723 1270
rect 863 1274 867 1275
rect 863 1269 867 1270
rect 879 1274 883 1275
rect 879 1269 883 1270
rect 1055 1274 1059 1275
rect 1055 1269 1059 1270
rect 1063 1274 1067 1275
rect 1063 1269 1067 1270
rect 1255 1274 1259 1275
rect 1255 1269 1259 1270
rect 1263 1274 1267 1275
rect 1263 1269 1267 1270
rect 1431 1274 1435 1275
rect 1431 1269 1435 1270
rect 1487 1274 1491 1275
rect 1487 1269 1491 1270
rect 1607 1274 1611 1275
rect 1607 1269 1611 1270
rect 1719 1274 1723 1275
rect 1719 1269 1723 1270
rect 1783 1274 1787 1275
rect 1783 1269 1787 1270
rect 1935 1274 1939 1275
rect 1935 1269 1939 1270
rect 2031 1274 2035 1275
rect 2031 1269 2035 1270
rect 112 1241 114 1269
rect 208 1260 210 1269
rect 328 1260 330 1269
rect 456 1260 458 1269
rect 584 1260 586 1269
rect 720 1260 722 1269
rect 880 1260 882 1269
rect 1056 1260 1058 1269
rect 1264 1260 1266 1269
rect 1488 1260 1490 1269
rect 1720 1260 1722 1269
rect 1936 1260 1938 1269
rect 206 1259 212 1260
rect 206 1255 207 1259
rect 211 1255 212 1259
rect 206 1254 212 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 454 1259 460 1260
rect 454 1255 455 1259
rect 459 1255 460 1259
rect 454 1254 460 1255
rect 582 1259 588 1260
rect 582 1255 583 1259
rect 587 1255 588 1259
rect 582 1254 588 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 878 1259 884 1260
rect 878 1255 879 1259
rect 883 1255 884 1259
rect 878 1254 884 1255
rect 1054 1259 1060 1260
rect 1054 1255 1055 1259
rect 1059 1255 1060 1259
rect 1054 1254 1060 1255
rect 1262 1259 1268 1260
rect 1262 1255 1263 1259
rect 1267 1255 1268 1259
rect 1262 1254 1268 1255
rect 1486 1259 1492 1260
rect 1486 1255 1487 1259
rect 1491 1255 1492 1259
rect 1486 1254 1492 1255
rect 1718 1259 1724 1260
rect 1718 1255 1719 1259
rect 1723 1255 1724 1259
rect 1718 1254 1724 1255
rect 1934 1259 1940 1260
rect 1934 1255 1935 1259
rect 1939 1255 1940 1259
rect 1934 1254 1940 1255
rect 2032 1241 2034 1269
rect 2072 1253 2074 1281
rect 2112 1272 2114 1281
rect 2344 1272 2346 1281
rect 2584 1272 2586 1281
rect 2800 1272 2802 1281
rect 3000 1272 3002 1281
rect 3184 1272 3186 1281
rect 3344 1272 3346 1281
rect 3496 1272 3498 1281
rect 3640 1272 3642 1281
rect 3776 1272 3778 1281
rect 3896 1272 3898 1281
rect 2110 1271 2116 1272
rect 2110 1267 2111 1271
rect 2115 1267 2116 1271
rect 2110 1266 2116 1267
rect 2342 1271 2348 1272
rect 2342 1267 2343 1271
rect 2347 1267 2348 1271
rect 2342 1266 2348 1267
rect 2582 1271 2588 1272
rect 2582 1267 2583 1271
rect 2587 1267 2588 1271
rect 2582 1266 2588 1267
rect 2798 1271 2804 1272
rect 2798 1267 2799 1271
rect 2803 1267 2804 1271
rect 2798 1266 2804 1267
rect 2998 1271 3004 1272
rect 2998 1267 2999 1271
rect 3003 1267 3004 1271
rect 2998 1266 3004 1267
rect 3182 1271 3188 1272
rect 3182 1267 3183 1271
rect 3187 1267 3188 1271
rect 3182 1266 3188 1267
rect 3342 1271 3348 1272
rect 3342 1267 3343 1271
rect 3347 1267 3348 1271
rect 3342 1266 3348 1267
rect 3494 1271 3500 1272
rect 3494 1267 3495 1271
rect 3499 1267 3500 1271
rect 3494 1266 3500 1267
rect 3638 1271 3644 1272
rect 3638 1267 3639 1271
rect 3643 1267 3644 1271
rect 3638 1266 3644 1267
rect 3774 1271 3780 1272
rect 3774 1267 3775 1271
rect 3779 1267 3780 1271
rect 3774 1266 3780 1267
rect 3894 1271 3900 1272
rect 3894 1267 3895 1271
rect 3899 1267 3900 1271
rect 3894 1266 3900 1267
rect 3992 1253 3994 1281
rect 2070 1252 2076 1253
rect 2070 1248 2071 1252
rect 2075 1248 2076 1252
rect 2070 1247 2076 1248
rect 3990 1252 3996 1253
rect 3990 1248 3991 1252
rect 3995 1248 3996 1252
rect 3990 1247 3996 1248
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 110 1235 116 1236
rect 2030 1240 2036 1241
rect 2030 1236 2031 1240
rect 2035 1236 2036 1240
rect 2030 1235 2036 1236
rect 2070 1235 2076 1236
rect 2070 1231 2071 1235
rect 2075 1231 2076 1235
rect 3990 1235 3996 1236
rect 3990 1231 3991 1235
rect 3995 1231 3996 1235
rect 2070 1230 2076 1231
rect 2110 1230 2116 1231
rect 110 1223 116 1224
rect 110 1219 111 1223
rect 115 1219 116 1223
rect 2030 1223 2036 1224
rect 2030 1219 2031 1223
rect 2035 1219 2036 1223
rect 110 1218 116 1219
rect 206 1218 212 1219
rect 112 1195 114 1218
rect 206 1214 207 1218
rect 211 1214 212 1218
rect 206 1213 212 1214
rect 326 1218 332 1219
rect 326 1214 327 1218
rect 331 1214 332 1218
rect 326 1213 332 1214
rect 454 1218 460 1219
rect 454 1214 455 1218
rect 459 1214 460 1218
rect 454 1213 460 1214
rect 582 1218 588 1219
rect 582 1214 583 1218
rect 587 1214 588 1218
rect 582 1213 588 1214
rect 718 1218 724 1219
rect 718 1214 719 1218
rect 723 1214 724 1218
rect 718 1213 724 1214
rect 878 1218 884 1219
rect 878 1214 879 1218
rect 883 1214 884 1218
rect 878 1213 884 1214
rect 1054 1218 1060 1219
rect 1054 1214 1055 1218
rect 1059 1214 1060 1218
rect 1054 1213 1060 1214
rect 1262 1218 1268 1219
rect 1262 1214 1263 1218
rect 1267 1214 1268 1218
rect 1262 1213 1268 1214
rect 1486 1218 1492 1219
rect 1486 1214 1487 1218
rect 1491 1214 1492 1218
rect 1486 1213 1492 1214
rect 1718 1218 1724 1219
rect 1718 1214 1719 1218
rect 1723 1214 1724 1218
rect 1718 1213 1724 1214
rect 1934 1218 1940 1219
rect 2030 1218 2036 1219
rect 1934 1214 1935 1218
rect 1939 1214 1940 1218
rect 1934 1213 1940 1214
rect 208 1195 210 1213
rect 328 1195 330 1213
rect 456 1195 458 1213
rect 584 1195 586 1213
rect 720 1195 722 1213
rect 880 1195 882 1213
rect 1056 1195 1058 1213
rect 1264 1195 1266 1213
rect 1488 1195 1490 1213
rect 1720 1195 1722 1213
rect 1936 1195 1938 1213
rect 2032 1195 2034 1218
rect 2072 1211 2074 1230
rect 2110 1226 2111 1230
rect 2115 1226 2116 1230
rect 2110 1225 2116 1226
rect 2342 1230 2348 1231
rect 2342 1226 2343 1230
rect 2347 1226 2348 1230
rect 2342 1225 2348 1226
rect 2582 1230 2588 1231
rect 2582 1226 2583 1230
rect 2587 1226 2588 1230
rect 2582 1225 2588 1226
rect 2798 1230 2804 1231
rect 2798 1226 2799 1230
rect 2803 1226 2804 1230
rect 2798 1225 2804 1226
rect 2998 1230 3004 1231
rect 2998 1226 2999 1230
rect 3003 1226 3004 1230
rect 2998 1225 3004 1226
rect 3182 1230 3188 1231
rect 3182 1226 3183 1230
rect 3187 1226 3188 1230
rect 3182 1225 3188 1226
rect 3342 1230 3348 1231
rect 3342 1226 3343 1230
rect 3347 1226 3348 1230
rect 3342 1225 3348 1226
rect 3494 1230 3500 1231
rect 3494 1226 3495 1230
rect 3499 1226 3500 1230
rect 3494 1225 3500 1226
rect 3638 1230 3644 1231
rect 3638 1226 3639 1230
rect 3643 1226 3644 1230
rect 3638 1225 3644 1226
rect 3774 1230 3780 1231
rect 3774 1226 3775 1230
rect 3779 1226 3780 1230
rect 3774 1225 3780 1226
rect 3894 1230 3900 1231
rect 3990 1230 3996 1231
rect 3894 1226 3895 1230
rect 3899 1226 3900 1230
rect 3894 1225 3900 1226
rect 2112 1211 2114 1225
rect 2344 1211 2346 1225
rect 2584 1211 2586 1225
rect 2800 1211 2802 1225
rect 3000 1211 3002 1225
rect 3184 1211 3186 1225
rect 3344 1211 3346 1225
rect 3496 1211 3498 1225
rect 3640 1211 3642 1225
rect 3776 1211 3778 1225
rect 3896 1211 3898 1225
rect 3992 1211 3994 1230
rect 2071 1210 2075 1211
rect 2071 1205 2075 1206
rect 2111 1210 2115 1211
rect 2111 1205 2115 1206
rect 2279 1210 2283 1211
rect 2279 1205 2283 1206
rect 2343 1210 2347 1211
rect 2343 1205 2347 1206
rect 2471 1210 2475 1211
rect 2471 1205 2475 1206
rect 2583 1210 2587 1211
rect 2583 1205 2587 1206
rect 2655 1210 2659 1211
rect 2655 1205 2659 1206
rect 2799 1210 2803 1211
rect 2799 1205 2803 1206
rect 2831 1210 2835 1211
rect 2831 1205 2835 1206
rect 2999 1210 3003 1211
rect 2999 1205 3003 1206
rect 3159 1210 3163 1211
rect 3159 1205 3163 1206
rect 3183 1210 3187 1211
rect 3183 1205 3187 1206
rect 3327 1210 3331 1211
rect 3327 1205 3331 1206
rect 3343 1210 3347 1211
rect 3343 1205 3347 1206
rect 3495 1210 3499 1211
rect 3495 1205 3499 1206
rect 3639 1210 3643 1211
rect 3639 1205 3643 1206
rect 3775 1210 3779 1211
rect 3775 1205 3779 1206
rect 3895 1210 3899 1211
rect 3895 1205 3899 1206
rect 3991 1210 3995 1211
rect 3991 1205 3995 1206
rect 111 1194 115 1195
rect 111 1189 115 1190
rect 207 1194 211 1195
rect 207 1189 211 1190
rect 327 1194 331 1195
rect 327 1189 331 1190
rect 455 1194 459 1195
rect 455 1189 459 1190
rect 471 1194 475 1195
rect 471 1189 475 1190
rect 583 1194 587 1195
rect 583 1189 587 1190
rect 703 1194 707 1195
rect 703 1189 707 1190
rect 719 1194 723 1195
rect 719 1189 723 1190
rect 823 1194 827 1195
rect 823 1189 827 1190
rect 879 1194 883 1195
rect 879 1189 883 1190
rect 943 1194 947 1195
rect 943 1189 947 1190
rect 1055 1194 1059 1195
rect 1055 1189 1059 1190
rect 1063 1194 1067 1195
rect 1063 1189 1067 1190
rect 1183 1194 1187 1195
rect 1183 1189 1187 1190
rect 1263 1194 1267 1195
rect 1263 1189 1267 1190
rect 1303 1194 1307 1195
rect 1303 1189 1307 1190
rect 1423 1194 1427 1195
rect 1423 1189 1427 1190
rect 1487 1194 1491 1195
rect 1487 1189 1491 1190
rect 1543 1194 1547 1195
rect 1543 1189 1547 1190
rect 1719 1194 1723 1195
rect 1719 1189 1723 1190
rect 1935 1194 1939 1195
rect 1935 1189 1939 1190
rect 2031 1194 2035 1195
rect 2072 1190 2074 1205
rect 2112 1195 2114 1205
rect 2280 1195 2282 1205
rect 2472 1195 2474 1205
rect 2656 1195 2658 1205
rect 2832 1195 2834 1205
rect 3000 1195 3002 1205
rect 3160 1195 3162 1205
rect 3328 1195 3330 1205
rect 3496 1195 3498 1205
rect 2110 1194 2116 1195
rect 2110 1190 2111 1194
rect 2115 1190 2116 1194
rect 2031 1189 2035 1190
rect 2070 1189 2076 1190
rect 2110 1189 2116 1190
rect 2278 1194 2284 1195
rect 2278 1190 2279 1194
rect 2283 1190 2284 1194
rect 2278 1189 2284 1190
rect 2470 1194 2476 1195
rect 2470 1190 2471 1194
rect 2475 1190 2476 1194
rect 2470 1189 2476 1190
rect 2654 1194 2660 1195
rect 2654 1190 2655 1194
rect 2659 1190 2660 1194
rect 2654 1189 2660 1190
rect 2830 1194 2836 1195
rect 2830 1190 2831 1194
rect 2835 1190 2836 1194
rect 2830 1189 2836 1190
rect 2998 1194 3004 1195
rect 2998 1190 2999 1194
rect 3003 1190 3004 1194
rect 2998 1189 3004 1190
rect 3158 1194 3164 1195
rect 3158 1190 3159 1194
rect 3163 1190 3164 1194
rect 3158 1189 3164 1190
rect 3326 1194 3332 1195
rect 3326 1190 3327 1194
rect 3331 1190 3332 1194
rect 3326 1189 3332 1190
rect 3494 1194 3500 1195
rect 3494 1190 3495 1194
rect 3499 1190 3500 1194
rect 3992 1190 3994 1205
rect 3494 1189 3500 1190
rect 3990 1189 3996 1190
rect 112 1174 114 1189
rect 472 1179 474 1189
rect 584 1179 586 1189
rect 704 1179 706 1189
rect 824 1179 826 1189
rect 944 1179 946 1189
rect 1064 1179 1066 1189
rect 1184 1179 1186 1189
rect 1304 1179 1306 1189
rect 1424 1179 1426 1189
rect 1544 1179 1546 1189
rect 470 1178 476 1179
rect 470 1174 471 1178
rect 475 1174 476 1178
rect 110 1173 116 1174
rect 470 1173 476 1174
rect 582 1178 588 1179
rect 582 1174 583 1178
rect 587 1174 588 1178
rect 582 1173 588 1174
rect 702 1178 708 1179
rect 702 1174 703 1178
rect 707 1174 708 1178
rect 702 1173 708 1174
rect 822 1178 828 1179
rect 822 1174 823 1178
rect 827 1174 828 1178
rect 822 1173 828 1174
rect 942 1178 948 1179
rect 942 1174 943 1178
rect 947 1174 948 1178
rect 942 1173 948 1174
rect 1062 1178 1068 1179
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1182 1178 1188 1179
rect 1182 1174 1183 1178
rect 1187 1174 1188 1178
rect 1182 1173 1188 1174
rect 1302 1178 1308 1179
rect 1302 1174 1303 1178
rect 1307 1174 1308 1178
rect 1302 1173 1308 1174
rect 1422 1178 1428 1179
rect 1422 1174 1423 1178
rect 1427 1174 1428 1178
rect 1422 1173 1428 1174
rect 1542 1178 1548 1179
rect 1542 1174 1543 1178
rect 1547 1174 1548 1178
rect 2032 1174 2034 1189
rect 2070 1185 2071 1189
rect 2075 1185 2076 1189
rect 2070 1184 2076 1185
rect 3990 1185 3991 1189
rect 3995 1185 3996 1189
rect 3990 1184 3996 1185
rect 1542 1173 1548 1174
rect 2030 1173 2036 1174
rect 110 1169 111 1173
rect 115 1169 116 1173
rect 110 1168 116 1169
rect 2030 1169 2031 1173
rect 2035 1169 2036 1173
rect 2030 1168 2036 1169
rect 2070 1172 2076 1173
rect 2070 1168 2071 1172
rect 2075 1168 2076 1172
rect 2070 1167 2076 1168
rect 3990 1172 3996 1173
rect 3990 1168 3991 1172
rect 3995 1168 3996 1172
rect 3990 1167 3996 1168
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 110 1151 116 1152
rect 2030 1156 2036 1157
rect 2030 1152 2031 1156
rect 2035 1152 2036 1156
rect 2030 1151 2036 1152
rect 112 1115 114 1151
rect 470 1137 476 1138
rect 470 1133 471 1137
rect 475 1133 476 1137
rect 470 1132 476 1133
rect 582 1137 588 1138
rect 582 1133 583 1137
rect 587 1133 588 1137
rect 582 1132 588 1133
rect 702 1137 708 1138
rect 702 1133 703 1137
rect 707 1133 708 1137
rect 702 1132 708 1133
rect 822 1137 828 1138
rect 822 1133 823 1137
rect 827 1133 828 1137
rect 822 1132 828 1133
rect 942 1137 948 1138
rect 942 1133 943 1137
rect 947 1133 948 1137
rect 942 1132 948 1133
rect 1062 1137 1068 1138
rect 1062 1133 1063 1137
rect 1067 1133 1068 1137
rect 1062 1132 1068 1133
rect 1182 1137 1188 1138
rect 1182 1133 1183 1137
rect 1187 1133 1188 1137
rect 1182 1132 1188 1133
rect 1302 1137 1308 1138
rect 1302 1133 1303 1137
rect 1307 1133 1308 1137
rect 1302 1132 1308 1133
rect 1422 1137 1428 1138
rect 1422 1133 1423 1137
rect 1427 1133 1428 1137
rect 1422 1132 1428 1133
rect 1542 1137 1548 1138
rect 1542 1133 1543 1137
rect 1547 1133 1548 1137
rect 1542 1132 1548 1133
rect 472 1115 474 1132
rect 584 1115 586 1132
rect 704 1115 706 1132
rect 824 1115 826 1132
rect 944 1115 946 1132
rect 1064 1115 1066 1132
rect 1184 1115 1186 1132
rect 1304 1115 1306 1132
rect 1424 1115 1426 1132
rect 1544 1115 1546 1132
rect 2032 1115 2034 1151
rect 2072 1135 2074 1167
rect 2110 1153 2116 1154
rect 2110 1149 2111 1153
rect 2115 1149 2116 1153
rect 2110 1148 2116 1149
rect 2278 1153 2284 1154
rect 2278 1149 2279 1153
rect 2283 1149 2284 1153
rect 2278 1148 2284 1149
rect 2470 1153 2476 1154
rect 2470 1149 2471 1153
rect 2475 1149 2476 1153
rect 2470 1148 2476 1149
rect 2654 1153 2660 1154
rect 2654 1149 2655 1153
rect 2659 1149 2660 1153
rect 2654 1148 2660 1149
rect 2830 1153 2836 1154
rect 2830 1149 2831 1153
rect 2835 1149 2836 1153
rect 2830 1148 2836 1149
rect 2998 1153 3004 1154
rect 2998 1149 2999 1153
rect 3003 1149 3004 1153
rect 2998 1148 3004 1149
rect 3158 1153 3164 1154
rect 3158 1149 3159 1153
rect 3163 1149 3164 1153
rect 3158 1148 3164 1149
rect 3326 1153 3332 1154
rect 3326 1149 3327 1153
rect 3331 1149 3332 1153
rect 3326 1148 3332 1149
rect 3494 1153 3500 1154
rect 3494 1149 3495 1153
rect 3499 1149 3500 1153
rect 3494 1148 3500 1149
rect 2112 1135 2114 1148
rect 2280 1135 2282 1148
rect 2472 1135 2474 1148
rect 2656 1135 2658 1148
rect 2832 1135 2834 1148
rect 3000 1135 3002 1148
rect 3160 1135 3162 1148
rect 3328 1135 3330 1148
rect 3496 1135 3498 1148
rect 3992 1135 3994 1167
rect 2071 1134 2075 1135
rect 2071 1129 2075 1130
rect 2111 1134 2115 1135
rect 2111 1129 2115 1130
rect 2279 1134 2283 1135
rect 2279 1129 2283 1130
rect 2295 1134 2299 1135
rect 2295 1129 2299 1130
rect 2471 1134 2475 1135
rect 2471 1129 2475 1130
rect 2503 1134 2507 1135
rect 2503 1129 2507 1130
rect 2655 1134 2659 1135
rect 2655 1129 2659 1130
rect 2703 1134 2707 1135
rect 2703 1129 2707 1130
rect 2831 1134 2835 1135
rect 2831 1129 2835 1130
rect 2895 1134 2899 1135
rect 2895 1129 2899 1130
rect 2999 1134 3003 1135
rect 2999 1129 3003 1130
rect 3079 1134 3083 1135
rect 3079 1129 3083 1130
rect 3159 1134 3163 1135
rect 3159 1129 3163 1130
rect 3255 1134 3259 1135
rect 3255 1129 3259 1130
rect 3327 1134 3331 1135
rect 3327 1129 3331 1130
rect 3431 1134 3435 1135
rect 3431 1129 3435 1130
rect 3495 1134 3499 1135
rect 3495 1129 3499 1130
rect 3615 1134 3619 1135
rect 3615 1129 3619 1130
rect 3991 1134 3995 1135
rect 3991 1129 3995 1130
rect 111 1114 115 1115
rect 111 1109 115 1110
rect 471 1114 475 1115
rect 471 1109 475 1110
rect 583 1114 587 1115
rect 583 1109 587 1110
rect 623 1114 627 1115
rect 623 1109 627 1110
rect 703 1114 707 1115
rect 703 1109 707 1110
rect 735 1114 739 1115
rect 735 1109 739 1110
rect 823 1114 827 1115
rect 823 1109 827 1110
rect 855 1114 859 1115
rect 855 1109 859 1110
rect 943 1114 947 1115
rect 943 1109 947 1110
rect 975 1114 979 1115
rect 975 1109 979 1110
rect 1063 1114 1067 1115
rect 1063 1109 1067 1110
rect 1095 1114 1099 1115
rect 1095 1109 1099 1110
rect 1183 1114 1187 1115
rect 1183 1109 1187 1110
rect 1215 1114 1219 1115
rect 1215 1109 1219 1110
rect 1303 1114 1307 1115
rect 1303 1109 1307 1110
rect 1335 1114 1339 1115
rect 1335 1109 1339 1110
rect 1423 1114 1427 1115
rect 1423 1109 1427 1110
rect 1455 1114 1459 1115
rect 1455 1109 1459 1110
rect 1543 1114 1547 1115
rect 1543 1109 1547 1110
rect 1575 1114 1579 1115
rect 1575 1109 1579 1110
rect 1703 1114 1707 1115
rect 1703 1109 1707 1110
rect 2031 1114 2035 1115
rect 2031 1109 2035 1110
rect 112 1081 114 1109
rect 624 1100 626 1109
rect 736 1100 738 1109
rect 856 1100 858 1109
rect 976 1100 978 1109
rect 1096 1100 1098 1109
rect 1216 1100 1218 1109
rect 1336 1100 1338 1109
rect 1456 1100 1458 1109
rect 1576 1100 1578 1109
rect 1704 1100 1706 1109
rect 622 1099 628 1100
rect 622 1095 623 1099
rect 627 1095 628 1099
rect 622 1094 628 1095
rect 734 1099 740 1100
rect 734 1095 735 1099
rect 739 1095 740 1099
rect 734 1094 740 1095
rect 854 1099 860 1100
rect 854 1095 855 1099
rect 859 1095 860 1099
rect 854 1094 860 1095
rect 974 1099 980 1100
rect 974 1095 975 1099
rect 979 1095 980 1099
rect 974 1094 980 1095
rect 1094 1099 1100 1100
rect 1094 1095 1095 1099
rect 1099 1095 1100 1099
rect 1094 1094 1100 1095
rect 1214 1099 1220 1100
rect 1214 1095 1215 1099
rect 1219 1095 1220 1099
rect 1214 1094 1220 1095
rect 1334 1099 1340 1100
rect 1334 1095 1335 1099
rect 1339 1095 1340 1099
rect 1334 1094 1340 1095
rect 1454 1099 1460 1100
rect 1454 1095 1455 1099
rect 1459 1095 1460 1099
rect 1454 1094 1460 1095
rect 1574 1099 1580 1100
rect 1574 1095 1575 1099
rect 1579 1095 1580 1099
rect 1574 1094 1580 1095
rect 1702 1099 1708 1100
rect 1702 1095 1703 1099
rect 1707 1095 1708 1099
rect 1702 1094 1708 1095
rect 2032 1081 2034 1109
rect 2072 1101 2074 1129
rect 2112 1120 2114 1129
rect 2296 1120 2298 1129
rect 2504 1120 2506 1129
rect 2704 1120 2706 1129
rect 2896 1120 2898 1129
rect 3080 1120 3082 1129
rect 3256 1120 3258 1129
rect 3432 1120 3434 1129
rect 3616 1120 3618 1129
rect 2110 1119 2116 1120
rect 2110 1115 2111 1119
rect 2115 1115 2116 1119
rect 2110 1114 2116 1115
rect 2294 1119 2300 1120
rect 2294 1115 2295 1119
rect 2299 1115 2300 1119
rect 2294 1114 2300 1115
rect 2502 1119 2508 1120
rect 2502 1115 2503 1119
rect 2507 1115 2508 1119
rect 2502 1114 2508 1115
rect 2702 1119 2708 1120
rect 2702 1115 2703 1119
rect 2707 1115 2708 1119
rect 2702 1114 2708 1115
rect 2894 1119 2900 1120
rect 2894 1115 2895 1119
rect 2899 1115 2900 1119
rect 2894 1114 2900 1115
rect 3078 1119 3084 1120
rect 3078 1115 3079 1119
rect 3083 1115 3084 1119
rect 3078 1114 3084 1115
rect 3254 1119 3260 1120
rect 3254 1115 3255 1119
rect 3259 1115 3260 1119
rect 3254 1114 3260 1115
rect 3430 1119 3436 1120
rect 3430 1115 3431 1119
rect 3435 1115 3436 1119
rect 3430 1114 3436 1115
rect 3614 1119 3620 1120
rect 3614 1115 3615 1119
rect 3619 1115 3620 1119
rect 3614 1114 3620 1115
rect 3992 1101 3994 1129
rect 2070 1100 2076 1101
rect 2070 1096 2071 1100
rect 2075 1096 2076 1100
rect 2070 1095 2076 1096
rect 3990 1100 3996 1101
rect 3990 1096 3991 1100
rect 3995 1096 3996 1100
rect 3990 1095 3996 1096
rect 2070 1083 2076 1084
rect 110 1080 116 1081
rect 110 1076 111 1080
rect 115 1076 116 1080
rect 110 1075 116 1076
rect 2030 1080 2036 1081
rect 2030 1076 2031 1080
rect 2035 1076 2036 1080
rect 2070 1079 2071 1083
rect 2075 1079 2076 1083
rect 3990 1083 3996 1084
rect 3990 1079 3991 1083
rect 3995 1079 3996 1083
rect 2070 1078 2076 1079
rect 2110 1078 2116 1079
rect 2030 1075 2036 1076
rect 110 1063 116 1064
rect 110 1059 111 1063
rect 115 1059 116 1063
rect 2030 1063 2036 1064
rect 2030 1059 2031 1063
rect 2035 1059 2036 1063
rect 110 1058 116 1059
rect 622 1058 628 1059
rect 112 1035 114 1058
rect 622 1054 623 1058
rect 627 1054 628 1058
rect 622 1053 628 1054
rect 734 1058 740 1059
rect 734 1054 735 1058
rect 739 1054 740 1058
rect 734 1053 740 1054
rect 854 1058 860 1059
rect 854 1054 855 1058
rect 859 1054 860 1058
rect 854 1053 860 1054
rect 974 1058 980 1059
rect 974 1054 975 1058
rect 979 1054 980 1058
rect 974 1053 980 1054
rect 1094 1058 1100 1059
rect 1094 1054 1095 1058
rect 1099 1054 1100 1058
rect 1094 1053 1100 1054
rect 1214 1058 1220 1059
rect 1214 1054 1215 1058
rect 1219 1054 1220 1058
rect 1214 1053 1220 1054
rect 1334 1058 1340 1059
rect 1334 1054 1335 1058
rect 1339 1054 1340 1058
rect 1334 1053 1340 1054
rect 1454 1058 1460 1059
rect 1454 1054 1455 1058
rect 1459 1054 1460 1058
rect 1454 1053 1460 1054
rect 1574 1058 1580 1059
rect 1574 1054 1575 1058
rect 1579 1054 1580 1058
rect 1574 1053 1580 1054
rect 1702 1058 1708 1059
rect 2030 1058 2036 1059
rect 1702 1054 1703 1058
rect 1707 1054 1708 1058
rect 1702 1053 1708 1054
rect 624 1035 626 1053
rect 736 1035 738 1053
rect 856 1035 858 1053
rect 976 1035 978 1053
rect 1096 1035 1098 1053
rect 1216 1035 1218 1053
rect 1336 1035 1338 1053
rect 1456 1035 1458 1053
rect 1576 1035 1578 1053
rect 1704 1035 1706 1053
rect 2032 1035 2034 1058
rect 2072 1055 2074 1078
rect 2110 1074 2111 1078
rect 2115 1074 2116 1078
rect 2110 1073 2116 1074
rect 2294 1078 2300 1079
rect 2294 1074 2295 1078
rect 2299 1074 2300 1078
rect 2294 1073 2300 1074
rect 2502 1078 2508 1079
rect 2502 1074 2503 1078
rect 2507 1074 2508 1078
rect 2502 1073 2508 1074
rect 2702 1078 2708 1079
rect 2702 1074 2703 1078
rect 2707 1074 2708 1078
rect 2702 1073 2708 1074
rect 2894 1078 2900 1079
rect 2894 1074 2895 1078
rect 2899 1074 2900 1078
rect 2894 1073 2900 1074
rect 3078 1078 3084 1079
rect 3078 1074 3079 1078
rect 3083 1074 3084 1078
rect 3078 1073 3084 1074
rect 3254 1078 3260 1079
rect 3254 1074 3255 1078
rect 3259 1074 3260 1078
rect 3254 1073 3260 1074
rect 3430 1078 3436 1079
rect 3430 1074 3431 1078
rect 3435 1074 3436 1078
rect 3430 1073 3436 1074
rect 3614 1078 3620 1079
rect 3990 1078 3996 1079
rect 3614 1074 3615 1078
rect 3619 1074 3620 1078
rect 3614 1073 3620 1074
rect 2112 1055 2114 1073
rect 2296 1055 2298 1073
rect 2504 1055 2506 1073
rect 2704 1055 2706 1073
rect 2896 1055 2898 1073
rect 3080 1055 3082 1073
rect 3256 1055 3258 1073
rect 3432 1055 3434 1073
rect 3616 1055 3618 1073
rect 3992 1055 3994 1078
rect 2071 1054 2075 1055
rect 2071 1049 2075 1050
rect 2111 1054 2115 1055
rect 2111 1049 2115 1050
rect 2167 1054 2171 1055
rect 2167 1049 2171 1050
rect 2287 1054 2291 1055
rect 2287 1049 2291 1050
rect 2295 1054 2299 1055
rect 2295 1049 2299 1050
rect 2423 1054 2427 1055
rect 2423 1049 2427 1050
rect 2503 1054 2507 1055
rect 2503 1049 2507 1050
rect 2575 1054 2579 1055
rect 2575 1049 2579 1050
rect 2703 1054 2707 1055
rect 2703 1049 2707 1050
rect 2743 1054 2747 1055
rect 2743 1049 2747 1050
rect 2895 1054 2899 1055
rect 2895 1049 2899 1050
rect 2919 1054 2923 1055
rect 2919 1049 2923 1050
rect 3079 1054 3083 1055
rect 3079 1049 3083 1050
rect 3095 1054 3099 1055
rect 3095 1049 3099 1050
rect 3255 1054 3259 1055
rect 3255 1049 3259 1050
rect 3279 1054 3283 1055
rect 3279 1049 3283 1050
rect 3431 1054 3435 1055
rect 3431 1049 3435 1050
rect 3463 1054 3467 1055
rect 3463 1049 3467 1050
rect 3615 1054 3619 1055
rect 3615 1049 3619 1050
rect 3655 1054 3659 1055
rect 3655 1049 3659 1050
rect 3991 1054 3995 1055
rect 3991 1049 3995 1050
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 623 1034 627 1035
rect 623 1029 627 1030
rect 727 1034 731 1035
rect 727 1029 731 1030
rect 735 1034 739 1035
rect 735 1029 739 1030
rect 847 1034 851 1035
rect 847 1029 851 1030
rect 855 1034 859 1035
rect 855 1029 859 1030
rect 967 1034 971 1035
rect 967 1029 971 1030
rect 975 1034 979 1035
rect 975 1029 979 1030
rect 1095 1034 1099 1035
rect 1095 1029 1099 1030
rect 1215 1034 1219 1035
rect 1215 1029 1219 1030
rect 1223 1034 1227 1035
rect 1223 1029 1227 1030
rect 1335 1034 1339 1035
rect 1335 1029 1339 1030
rect 1351 1034 1355 1035
rect 1351 1029 1355 1030
rect 1455 1034 1459 1035
rect 1455 1029 1459 1030
rect 1479 1034 1483 1035
rect 1479 1029 1483 1030
rect 1575 1034 1579 1035
rect 1575 1029 1579 1030
rect 1607 1034 1611 1035
rect 1607 1029 1611 1030
rect 1703 1034 1707 1035
rect 1703 1029 1707 1030
rect 1735 1034 1739 1035
rect 1735 1029 1739 1030
rect 1863 1034 1867 1035
rect 1863 1029 1867 1030
rect 2031 1034 2035 1035
rect 2072 1034 2074 1049
rect 2168 1039 2170 1049
rect 2288 1039 2290 1049
rect 2424 1039 2426 1049
rect 2576 1039 2578 1049
rect 2744 1039 2746 1049
rect 2920 1039 2922 1049
rect 3096 1039 3098 1049
rect 3280 1039 3282 1049
rect 3464 1039 3466 1049
rect 3656 1039 3658 1049
rect 2166 1038 2172 1039
rect 2166 1034 2167 1038
rect 2171 1034 2172 1038
rect 2031 1029 2035 1030
rect 2070 1033 2076 1034
rect 2166 1033 2172 1034
rect 2286 1038 2292 1039
rect 2286 1034 2287 1038
rect 2291 1034 2292 1038
rect 2286 1033 2292 1034
rect 2422 1038 2428 1039
rect 2422 1034 2423 1038
rect 2427 1034 2428 1038
rect 2422 1033 2428 1034
rect 2574 1038 2580 1039
rect 2574 1034 2575 1038
rect 2579 1034 2580 1038
rect 2574 1033 2580 1034
rect 2742 1038 2748 1039
rect 2742 1034 2743 1038
rect 2747 1034 2748 1038
rect 2742 1033 2748 1034
rect 2918 1038 2924 1039
rect 2918 1034 2919 1038
rect 2923 1034 2924 1038
rect 2918 1033 2924 1034
rect 3094 1038 3100 1039
rect 3094 1034 3095 1038
rect 3099 1034 3100 1038
rect 3094 1033 3100 1034
rect 3278 1038 3284 1039
rect 3278 1034 3279 1038
rect 3283 1034 3284 1038
rect 3278 1033 3284 1034
rect 3462 1038 3468 1039
rect 3462 1034 3463 1038
rect 3467 1034 3468 1038
rect 3462 1033 3468 1034
rect 3654 1038 3660 1039
rect 3654 1034 3655 1038
rect 3659 1034 3660 1038
rect 3992 1034 3994 1049
rect 3654 1033 3660 1034
rect 3990 1033 3996 1034
rect 2070 1029 2071 1033
rect 2075 1029 2076 1033
rect 112 1014 114 1029
rect 728 1019 730 1029
rect 848 1019 850 1029
rect 968 1019 970 1029
rect 1096 1019 1098 1029
rect 1224 1019 1226 1029
rect 1352 1019 1354 1029
rect 1480 1019 1482 1029
rect 1608 1019 1610 1029
rect 1736 1019 1738 1029
rect 1864 1019 1866 1029
rect 726 1018 732 1019
rect 726 1014 727 1018
rect 731 1014 732 1018
rect 110 1013 116 1014
rect 726 1013 732 1014
rect 846 1018 852 1019
rect 846 1014 847 1018
rect 851 1014 852 1018
rect 846 1013 852 1014
rect 966 1018 972 1019
rect 966 1014 967 1018
rect 971 1014 972 1018
rect 966 1013 972 1014
rect 1094 1018 1100 1019
rect 1094 1014 1095 1018
rect 1099 1014 1100 1018
rect 1094 1013 1100 1014
rect 1222 1018 1228 1019
rect 1222 1014 1223 1018
rect 1227 1014 1228 1018
rect 1222 1013 1228 1014
rect 1350 1018 1356 1019
rect 1350 1014 1351 1018
rect 1355 1014 1356 1018
rect 1350 1013 1356 1014
rect 1478 1018 1484 1019
rect 1478 1014 1479 1018
rect 1483 1014 1484 1018
rect 1478 1013 1484 1014
rect 1606 1018 1612 1019
rect 1606 1014 1607 1018
rect 1611 1014 1612 1018
rect 1606 1013 1612 1014
rect 1734 1018 1740 1019
rect 1734 1014 1735 1018
rect 1739 1014 1740 1018
rect 1734 1013 1740 1014
rect 1862 1018 1868 1019
rect 1862 1014 1863 1018
rect 1867 1014 1868 1018
rect 2032 1014 2034 1029
rect 2070 1028 2076 1029
rect 3990 1029 3991 1033
rect 3995 1029 3996 1033
rect 3990 1028 3996 1029
rect 2070 1016 2076 1017
rect 1862 1013 1868 1014
rect 2030 1013 2036 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 110 1008 116 1009
rect 2030 1009 2031 1013
rect 2035 1009 2036 1013
rect 2070 1012 2071 1016
rect 2075 1012 2076 1016
rect 2070 1011 2076 1012
rect 3990 1016 3996 1017
rect 3990 1012 3991 1016
rect 3995 1012 3996 1016
rect 3990 1011 3996 1012
rect 2030 1008 2036 1009
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 110 991 116 992
rect 2030 996 2036 997
rect 2030 992 2031 996
rect 2035 992 2036 996
rect 2030 991 2036 992
rect 112 955 114 991
rect 726 977 732 978
rect 726 973 727 977
rect 731 973 732 977
rect 726 972 732 973
rect 846 977 852 978
rect 846 973 847 977
rect 851 973 852 977
rect 846 972 852 973
rect 966 977 972 978
rect 966 973 967 977
rect 971 973 972 977
rect 966 972 972 973
rect 1094 977 1100 978
rect 1094 973 1095 977
rect 1099 973 1100 977
rect 1094 972 1100 973
rect 1222 977 1228 978
rect 1222 973 1223 977
rect 1227 973 1228 977
rect 1222 972 1228 973
rect 1350 977 1356 978
rect 1350 973 1351 977
rect 1355 973 1356 977
rect 1350 972 1356 973
rect 1478 977 1484 978
rect 1478 973 1479 977
rect 1483 973 1484 977
rect 1478 972 1484 973
rect 1606 977 1612 978
rect 1606 973 1607 977
rect 1611 973 1612 977
rect 1606 972 1612 973
rect 1734 977 1740 978
rect 1734 973 1735 977
rect 1739 973 1740 977
rect 1734 972 1740 973
rect 1862 977 1868 978
rect 1862 973 1863 977
rect 1867 973 1868 977
rect 1862 972 1868 973
rect 728 955 730 972
rect 848 955 850 972
rect 968 955 970 972
rect 1096 955 1098 972
rect 1224 955 1226 972
rect 1352 955 1354 972
rect 1480 955 1482 972
rect 1608 955 1610 972
rect 1736 955 1738 972
rect 1864 955 1866 972
rect 2032 955 2034 991
rect 2072 975 2074 1011
rect 2166 997 2172 998
rect 2166 993 2167 997
rect 2171 993 2172 997
rect 2166 992 2172 993
rect 2286 997 2292 998
rect 2286 993 2287 997
rect 2291 993 2292 997
rect 2286 992 2292 993
rect 2422 997 2428 998
rect 2422 993 2423 997
rect 2427 993 2428 997
rect 2422 992 2428 993
rect 2574 997 2580 998
rect 2574 993 2575 997
rect 2579 993 2580 997
rect 2574 992 2580 993
rect 2742 997 2748 998
rect 2742 993 2743 997
rect 2747 993 2748 997
rect 2742 992 2748 993
rect 2918 997 2924 998
rect 2918 993 2919 997
rect 2923 993 2924 997
rect 2918 992 2924 993
rect 3094 997 3100 998
rect 3094 993 3095 997
rect 3099 993 3100 997
rect 3094 992 3100 993
rect 3278 997 3284 998
rect 3278 993 3279 997
rect 3283 993 3284 997
rect 3278 992 3284 993
rect 3462 997 3468 998
rect 3462 993 3463 997
rect 3467 993 3468 997
rect 3462 992 3468 993
rect 3654 997 3660 998
rect 3654 993 3655 997
rect 3659 993 3660 997
rect 3654 992 3660 993
rect 2168 975 2170 992
rect 2288 975 2290 992
rect 2424 975 2426 992
rect 2576 975 2578 992
rect 2744 975 2746 992
rect 2920 975 2922 992
rect 3096 975 3098 992
rect 3280 975 3282 992
rect 3464 975 3466 992
rect 3656 975 3658 992
rect 3992 975 3994 1011
rect 2071 974 2075 975
rect 2071 969 2075 970
rect 2167 974 2171 975
rect 2167 969 2171 970
rect 2287 974 2291 975
rect 2287 969 2291 970
rect 2423 974 2427 975
rect 2423 969 2427 970
rect 2527 974 2531 975
rect 2527 969 2531 970
rect 2575 974 2579 975
rect 2575 969 2579 970
rect 2647 974 2651 975
rect 2647 969 2651 970
rect 2743 974 2747 975
rect 2743 969 2747 970
rect 2775 974 2779 975
rect 2775 969 2779 970
rect 2919 974 2923 975
rect 2919 969 2923 970
rect 3071 974 3075 975
rect 3071 969 3075 970
rect 3095 974 3099 975
rect 3095 969 3099 970
rect 3231 974 3235 975
rect 3231 969 3235 970
rect 3279 974 3283 975
rect 3279 969 3283 970
rect 3399 974 3403 975
rect 3399 969 3403 970
rect 3463 974 3467 975
rect 3463 969 3467 970
rect 3567 974 3571 975
rect 3567 969 3571 970
rect 3655 974 3659 975
rect 3655 969 3659 970
rect 3735 974 3739 975
rect 3735 969 3739 970
rect 3991 974 3995 975
rect 3991 969 3995 970
rect 111 954 115 955
rect 111 949 115 950
rect 591 954 595 955
rect 591 949 595 950
rect 727 954 731 955
rect 727 949 731 950
rect 735 954 739 955
rect 735 949 739 950
rect 847 954 851 955
rect 847 949 851 950
rect 887 954 891 955
rect 887 949 891 950
rect 967 954 971 955
rect 967 949 971 950
rect 1039 954 1043 955
rect 1039 949 1043 950
rect 1095 954 1099 955
rect 1095 949 1099 950
rect 1199 954 1203 955
rect 1199 949 1203 950
rect 1223 954 1227 955
rect 1223 949 1227 950
rect 1351 954 1355 955
rect 1351 949 1355 950
rect 1479 954 1483 955
rect 1479 949 1483 950
rect 1503 954 1507 955
rect 1503 949 1507 950
rect 1607 954 1611 955
rect 1607 949 1611 950
rect 1655 954 1659 955
rect 1655 949 1659 950
rect 1735 954 1739 955
rect 1735 949 1739 950
rect 1807 954 1811 955
rect 1807 949 1811 950
rect 1863 954 1867 955
rect 1863 949 1867 950
rect 1935 954 1939 955
rect 1935 949 1939 950
rect 2031 954 2035 955
rect 2031 949 2035 950
rect 112 921 114 949
rect 592 940 594 949
rect 736 940 738 949
rect 888 940 890 949
rect 1040 940 1042 949
rect 1200 940 1202 949
rect 1352 940 1354 949
rect 1504 940 1506 949
rect 1656 940 1658 949
rect 1808 940 1810 949
rect 1936 940 1938 949
rect 590 939 596 940
rect 590 935 591 939
rect 595 935 596 939
rect 590 934 596 935
rect 734 939 740 940
rect 734 935 735 939
rect 739 935 740 939
rect 734 934 740 935
rect 886 939 892 940
rect 886 935 887 939
rect 891 935 892 939
rect 886 934 892 935
rect 1038 939 1044 940
rect 1038 935 1039 939
rect 1043 935 1044 939
rect 1038 934 1044 935
rect 1198 939 1204 940
rect 1198 935 1199 939
rect 1203 935 1204 939
rect 1198 934 1204 935
rect 1350 939 1356 940
rect 1350 935 1351 939
rect 1355 935 1356 939
rect 1350 934 1356 935
rect 1502 939 1508 940
rect 1502 935 1503 939
rect 1507 935 1508 939
rect 1502 934 1508 935
rect 1654 939 1660 940
rect 1654 935 1655 939
rect 1659 935 1660 939
rect 1654 934 1660 935
rect 1806 939 1812 940
rect 1806 935 1807 939
rect 1811 935 1812 939
rect 1806 934 1812 935
rect 1934 939 1940 940
rect 1934 935 1935 939
rect 1939 935 1940 939
rect 1934 934 1940 935
rect 2032 921 2034 949
rect 2072 941 2074 969
rect 2528 960 2530 969
rect 2648 960 2650 969
rect 2776 960 2778 969
rect 2920 960 2922 969
rect 3072 960 3074 969
rect 3232 960 3234 969
rect 3400 960 3402 969
rect 3568 960 3570 969
rect 3736 960 3738 969
rect 2526 959 2532 960
rect 2526 955 2527 959
rect 2531 955 2532 959
rect 2526 954 2532 955
rect 2646 959 2652 960
rect 2646 955 2647 959
rect 2651 955 2652 959
rect 2646 954 2652 955
rect 2774 959 2780 960
rect 2774 955 2775 959
rect 2779 955 2780 959
rect 2774 954 2780 955
rect 2918 959 2924 960
rect 2918 955 2919 959
rect 2923 955 2924 959
rect 2918 954 2924 955
rect 3070 959 3076 960
rect 3070 955 3071 959
rect 3075 955 3076 959
rect 3070 954 3076 955
rect 3230 959 3236 960
rect 3230 955 3231 959
rect 3235 955 3236 959
rect 3230 954 3236 955
rect 3398 959 3404 960
rect 3398 955 3399 959
rect 3403 955 3404 959
rect 3398 954 3404 955
rect 3566 959 3572 960
rect 3566 955 3567 959
rect 3571 955 3572 959
rect 3566 954 3572 955
rect 3734 959 3740 960
rect 3734 955 3735 959
rect 3739 955 3740 959
rect 3734 954 3740 955
rect 3992 941 3994 969
rect 2070 940 2076 941
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 3990 940 3996 941
rect 3990 936 3991 940
rect 3995 936 3996 940
rect 3990 935 3996 936
rect 2070 923 2076 924
rect 110 920 116 921
rect 110 916 111 920
rect 115 916 116 920
rect 110 915 116 916
rect 2030 920 2036 921
rect 2030 916 2031 920
rect 2035 916 2036 920
rect 2070 919 2071 923
rect 2075 919 2076 923
rect 3990 923 3996 924
rect 3990 919 3991 923
rect 3995 919 3996 923
rect 2070 918 2076 919
rect 2526 918 2532 919
rect 2030 915 2036 916
rect 110 903 116 904
rect 110 899 111 903
rect 115 899 116 903
rect 2030 903 2036 904
rect 2030 899 2031 903
rect 2035 899 2036 903
rect 110 898 116 899
rect 590 898 596 899
rect 112 875 114 898
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 734 898 740 899
rect 734 894 735 898
rect 739 894 740 898
rect 734 893 740 894
rect 886 898 892 899
rect 886 894 887 898
rect 891 894 892 898
rect 886 893 892 894
rect 1038 898 1044 899
rect 1038 894 1039 898
rect 1043 894 1044 898
rect 1038 893 1044 894
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1350 898 1356 899
rect 1350 894 1351 898
rect 1355 894 1356 898
rect 1350 893 1356 894
rect 1502 898 1508 899
rect 1502 894 1503 898
rect 1507 894 1508 898
rect 1502 893 1508 894
rect 1654 898 1660 899
rect 1654 894 1655 898
rect 1659 894 1660 898
rect 1654 893 1660 894
rect 1806 898 1812 899
rect 1806 894 1807 898
rect 1811 894 1812 898
rect 1806 893 1812 894
rect 1934 898 1940 899
rect 2030 898 2036 899
rect 1934 894 1935 898
rect 1939 894 1940 898
rect 1934 893 1940 894
rect 592 875 594 893
rect 736 875 738 893
rect 888 875 890 893
rect 1040 875 1042 893
rect 1200 875 1202 893
rect 1352 875 1354 893
rect 1504 875 1506 893
rect 1656 875 1658 893
rect 1808 875 1810 893
rect 1936 875 1938 893
rect 2032 875 2034 898
rect 2072 891 2074 918
rect 2526 914 2527 918
rect 2531 914 2532 918
rect 2526 913 2532 914
rect 2646 918 2652 919
rect 2646 914 2647 918
rect 2651 914 2652 918
rect 2646 913 2652 914
rect 2774 918 2780 919
rect 2774 914 2775 918
rect 2779 914 2780 918
rect 2774 913 2780 914
rect 2918 918 2924 919
rect 2918 914 2919 918
rect 2923 914 2924 918
rect 2918 913 2924 914
rect 3070 918 3076 919
rect 3070 914 3071 918
rect 3075 914 3076 918
rect 3070 913 3076 914
rect 3230 918 3236 919
rect 3230 914 3231 918
rect 3235 914 3236 918
rect 3230 913 3236 914
rect 3398 918 3404 919
rect 3398 914 3399 918
rect 3403 914 3404 918
rect 3398 913 3404 914
rect 3566 918 3572 919
rect 3566 914 3567 918
rect 3571 914 3572 918
rect 3566 913 3572 914
rect 3734 918 3740 919
rect 3990 918 3996 919
rect 3734 914 3735 918
rect 3739 914 3740 918
rect 3734 913 3740 914
rect 2528 891 2530 913
rect 2648 891 2650 913
rect 2776 891 2778 913
rect 2920 891 2922 913
rect 3072 891 3074 913
rect 3232 891 3234 913
rect 3400 891 3402 913
rect 3568 891 3570 913
rect 3736 891 3738 913
rect 3992 891 3994 918
rect 2071 890 2075 891
rect 2071 885 2075 886
rect 2455 890 2459 891
rect 2455 885 2459 886
rect 2527 890 2531 891
rect 2527 885 2531 886
rect 2575 890 2579 891
rect 2575 885 2579 886
rect 2647 890 2651 891
rect 2647 885 2651 886
rect 2711 890 2715 891
rect 2711 885 2715 886
rect 2775 890 2779 891
rect 2775 885 2779 886
rect 2863 890 2867 891
rect 2863 885 2867 886
rect 2919 890 2923 891
rect 2919 885 2923 886
rect 3015 890 3019 891
rect 3015 885 3019 886
rect 3071 890 3075 891
rect 3071 885 3075 886
rect 3167 890 3171 891
rect 3167 885 3171 886
rect 3231 890 3235 891
rect 3231 885 3235 886
rect 3319 890 3323 891
rect 3319 885 3323 886
rect 3399 890 3403 891
rect 3399 885 3403 886
rect 3471 890 3475 891
rect 3471 885 3475 886
rect 3567 890 3571 891
rect 3567 885 3571 886
rect 3615 890 3619 891
rect 3615 885 3619 886
rect 3735 890 3739 891
rect 3735 885 3739 886
rect 3767 890 3771 891
rect 3767 885 3771 886
rect 3895 890 3899 891
rect 3895 885 3899 886
rect 3991 890 3995 891
rect 3991 885 3995 886
rect 111 874 115 875
rect 111 869 115 870
rect 439 874 443 875
rect 439 869 443 870
rect 583 874 587 875
rect 583 869 587 870
rect 591 874 595 875
rect 591 869 595 870
rect 735 874 739 875
rect 735 869 739 870
rect 887 874 891 875
rect 887 869 891 870
rect 1039 874 1043 875
rect 1039 869 1043 870
rect 1047 874 1051 875
rect 1047 869 1051 870
rect 1199 874 1203 875
rect 1199 869 1203 870
rect 1351 874 1355 875
rect 1351 869 1355 870
rect 1495 874 1499 875
rect 1495 869 1499 870
rect 1503 874 1507 875
rect 1503 869 1507 870
rect 1647 874 1651 875
rect 1647 869 1651 870
rect 1655 874 1659 875
rect 1655 869 1659 870
rect 1799 874 1803 875
rect 1799 869 1803 870
rect 1807 874 1811 875
rect 1807 869 1811 870
rect 1935 874 1939 875
rect 1935 869 1939 870
rect 2031 874 2035 875
rect 2072 870 2074 885
rect 2456 875 2458 885
rect 2576 875 2578 885
rect 2712 875 2714 885
rect 2864 875 2866 885
rect 3016 875 3018 885
rect 3168 875 3170 885
rect 3320 875 3322 885
rect 3472 875 3474 885
rect 3616 875 3618 885
rect 3768 875 3770 885
rect 3896 875 3898 885
rect 2454 874 2460 875
rect 2454 870 2455 874
rect 2459 870 2460 874
rect 2031 869 2035 870
rect 2070 869 2076 870
rect 2454 869 2460 870
rect 2574 874 2580 875
rect 2574 870 2575 874
rect 2579 870 2580 874
rect 2574 869 2580 870
rect 2710 874 2716 875
rect 2710 870 2711 874
rect 2715 870 2716 874
rect 2710 869 2716 870
rect 2862 874 2868 875
rect 2862 870 2863 874
rect 2867 870 2868 874
rect 2862 869 2868 870
rect 3014 874 3020 875
rect 3014 870 3015 874
rect 3019 870 3020 874
rect 3014 869 3020 870
rect 3166 874 3172 875
rect 3166 870 3167 874
rect 3171 870 3172 874
rect 3166 869 3172 870
rect 3318 874 3324 875
rect 3318 870 3319 874
rect 3323 870 3324 874
rect 3318 869 3324 870
rect 3470 874 3476 875
rect 3470 870 3471 874
rect 3475 870 3476 874
rect 3470 869 3476 870
rect 3614 874 3620 875
rect 3614 870 3615 874
rect 3619 870 3620 874
rect 3614 869 3620 870
rect 3766 874 3772 875
rect 3766 870 3767 874
rect 3771 870 3772 874
rect 3766 869 3772 870
rect 3894 874 3900 875
rect 3894 870 3895 874
rect 3899 870 3900 874
rect 3992 870 3994 885
rect 3894 869 3900 870
rect 3990 869 3996 870
rect 112 854 114 869
rect 440 859 442 869
rect 584 859 586 869
rect 736 859 738 869
rect 888 859 890 869
rect 1048 859 1050 869
rect 1200 859 1202 869
rect 1352 859 1354 869
rect 1496 859 1498 869
rect 1648 859 1650 869
rect 1800 859 1802 869
rect 438 858 444 859
rect 438 854 439 858
rect 443 854 444 858
rect 110 853 116 854
rect 438 853 444 854
rect 582 858 588 859
rect 582 854 583 858
rect 587 854 588 858
rect 582 853 588 854
rect 734 858 740 859
rect 734 854 735 858
rect 739 854 740 858
rect 734 853 740 854
rect 886 858 892 859
rect 886 854 887 858
rect 891 854 892 858
rect 886 853 892 854
rect 1046 858 1052 859
rect 1046 854 1047 858
rect 1051 854 1052 858
rect 1046 853 1052 854
rect 1198 858 1204 859
rect 1198 854 1199 858
rect 1203 854 1204 858
rect 1198 853 1204 854
rect 1350 858 1356 859
rect 1350 854 1351 858
rect 1355 854 1356 858
rect 1350 853 1356 854
rect 1494 858 1500 859
rect 1494 854 1495 858
rect 1499 854 1500 858
rect 1494 853 1500 854
rect 1646 858 1652 859
rect 1646 854 1647 858
rect 1651 854 1652 858
rect 1646 853 1652 854
rect 1798 858 1804 859
rect 1798 854 1799 858
rect 1803 854 1804 858
rect 2032 854 2034 869
rect 2070 865 2071 869
rect 2075 865 2076 869
rect 2070 864 2076 865
rect 3990 865 3991 869
rect 3995 865 3996 869
rect 3990 864 3996 865
rect 1798 853 1804 854
rect 2030 853 2036 854
rect 110 849 111 853
rect 115 849 116 853
rect 110 848 116 849
rect 2030 849 2031 853
rect 2035 849 2036 853
rect 2030 848 2036 849
rect 2070 852 2076 853
rect 2070 848 2071 852
rect 2075 848 2076 852
rect 2070 847 2076 848
rect 3990 852 3996 853
rect 3990 848 3991 852
rect 3995 848 3996 852
rect 3990 847 3996 848
rect 110 836 116 837
rect 110 832 111 836
rect 115 832 116 836
rect 110 831 116 832
rect 2030 836 2036 837
rect 2030 832 2031 836
rect 2035 832 2036 836
rect 2030 831 2036 832
rect 112 803 114 831
rect 438 817 444 818
rect 438 813 439 817
rect 443 813 444 817
rect 438 812 444 813
rect 582 817 588 818
rect 582 813 583 817
rect 587 813 588 817
rect 582 812 588 813
rect 734 817 740 818
rect 734 813 735 817
rect 739 813 740 817
rect 734 812 740 813
rect 886 817 892 818
rect 886 813 887 817
rect 891 813 892 817
rect 886 812 892 813
rect 1046 817 1052 818
rect 1046 813 1047 817
rect 1051 813 1052 817
rect 1046 812 1052 813
rect 1198 817 1204 818
rect 1198 813 1199 817
rect 1203 813 1204 817
rect 1198 812 1204 813
rect 1350 817 1356 818
rect 1350 813 1351 817
rect 1355 813 1356 817
rect 1350 812 1356 813
rect 1494 817 1500 818
rect 1494 813 1495 817
rect 1499 813 1500 817
rect 1494 812 1500 813
rect 1646 817 1652 818
rect 1646 813 1647 817
rect 1651 813 1652 817
rect 1646 812 1652 813
rect 1798 817 1804 818
rect 1798 813 1799 817
rect 1803 813 1804 817
rect 1798 812 1804 813
rect 440 803 442 812
rect 584 803 586 812
rect 736 803 738 812
rect 888 803 890 812
rect 1048 803 1050 812
rect 1200 803 1202 812
rect 1352 803 1354 812
rect 1496 803 1498 812
rect 1648 803 1650 812
rect 1800 803 1802 812
rect 2032 803 2034 831
rect 2072 819 2074 847
rect 2454 833 2460 834
rect 2454 829 2455 833
rect 2459 829 2460 833
rect 2454 828 2460 829
rect 2574 833 2580 834
rect 2574 829 2575 833
rect 2579 829 2580 833
rect 2574 828 2580 829
rect 2710 833 2716 834
rect 2710 829 2711 833
rect 2715 829 2716 833
rect 2710 828 2716 829
rect 2862 833 2868 834
rect 2862 829 2863 833
rect 2867 829 2868 833
rect 2862 828 2868 829
rect 3014 833 3020 834
rect 3014 829 3015 833
rect 3019 829 3020 833
rect 3014 828 3020 829
rect 3166 833 3172 834
rect 3166 829 3167 833
rect 3171 829 3172 833
rect 3166 828 3172 829
rect 3318 833 3324 834
rect 3318 829 3319 833
rect 3323 829 3324 833
rect 3318 828 3324 829
rect 3470 833 3476 834
rect 3470 829 3471 833
rect 3475 829 3476 833
rect 3470 828 3476 829
rect 3614 833 3620 834
rect 3614 829 3615 833
rect 3619 829 3620 833
rect 3614 828 3620 829
rect 3766 833 3772 834
rect 3766 829 3767 833
rect 3771 829 3772 833
rect 3766 828 3772 829
rect 3894 833 3900 834
rect 3894 829 3895 833
rect 3899 829 3900 833
rect 3894 828 3900 829
rect 2456 819 2458 828
rect 2576 819 2578 828
rect 2712 819 2714 828
rect 2864 819 2866 828
rect 3016 819 3018 828
rect 3168 819 3170 828
rect 3320 819 3322 828
rect 3472 819 3474 828
rect 3616 819 3618 828
rect 3768 819 3770 828
rect 3896 819 3898 828
rect 3992 819 3994 847
rect 2071 818 2075 819
rect 2071 813 2075 814
rect 2215 818 2219 819
rect 2215 813 2219 814
rect 2343 818 2347 819
rect 2343 813 2347 814
rect 2455 818 2459 819
rect 2455 813 2459 814
rect 2479 818 2483 819
rect 2479 813 2483 814
rect 2575 818 2579 819
rect 2575 813 2579 814
rect 2623 818 2627 819
rect 2623 813 2627 814
rect 2711 818 2715 819
rect 2711 813 2715 814
rect 2783 818 2787 819
rect 2783 813 2787 814
rect 2863 818 2867 819
rect 2863 813 2867 814
rect 2959 818 2963 819
rect 2959 813 2963 814
rect 3015 818 3019 819
rect 3015 813 3019 814
rect 3167 818 3171 819
rect 3167 813 3171 814
rect 3319 818 3323 819
rect 3319 813 3323 814
rect 3391 818 3395 819
rect 3391 813 3395 814
rect 3471 818 3475 819
rect 3471 813 3475 814
rect 3615 818 3619 819
rect 3615 813 3619 814
rect 3623 818 3627 819
rect 3623 813 3627 814
rect 3767 818 3771 819
rect 3767 813 3771 814
rect 3863 818 3867 819
rect 3863 813 3867 814
rect 3895 818 3899 819
rect 3895 813 3899 814
rect 3991 818 3995 819
rect 3991 813 3995 814
rect 111 802 115 803
rect 111 797 115 798
rect 279 802 283 803
rect 279 797 283 798
rect 431 802 435 803
rect 431 797 435 798
rect 439 802 443 803
rect 439 797 443 798
rect 583 802 587 803
rect 583 797 587 798
rect 591 802 595 803
rect 591 797 595 798
rect 735 802 739 803
rect 735 797 739 798
rect 751 802 755 803
rect 751 797 755 798
rect 887 802 891 803
rect 887 797 891 798
rect 919 802 923 803
rect 919 797 923 798
rect 1047 802 1051 803
rect 1047 797 1051 798
rect 1087 802 1091 803
rect 1087 797 1091 798
rect 1199 802 1203 803
rect 1199 797 1203 798
rect 1255 802 1259 803
rect 1255 797 1259 798
rect 1351 802 1355 803
rect 1351 797 1355 798
rect 1423 802 1427 803
rect 1423 797 1427 798
rect 1495 802 1499 803
rect 1495 797 1499 798
rect 1591 802 1595 803
rect 1591 797 1595 798
rect 1647 802 1651 803
rect 1647 797 1651 798
rect 1799 802 1803 803
rect 1799 797 1803 798
rect 2031 802 2035 803
rect 2031 797 2035 798
rect 112 769 114 797
rect 280 788 282 797
rect 432 788 434 797
rect 592 788 594 797
rect 752 788 754 797
rect 920 788 922 797
rect 1088 788 1090 797
rect 1256 788 1258 797
rect 1424 788 1426 797
rect 1592 788 1594 797
rect 278 787 284 788
rect 278 783 279 787
rect 283 783 284 787
rect 278 782 284 783
rect 430 787 436 788
rect 430 783 431 787
rect 435 783 436 787
rect 430 782 436 783
rect 590 787 596 788
rect 590 783 591 787
rect 595 783 596 787
rect 590 782 596 783
rect 750 787 756 788
rect 750 783 751 787
rect 755 783 756 787
rect 750 782 756 783
rect 918 787 924 788
rect 918 783 919 787
rect 923 783 924 787
rect 918 782 924 783
rect 1086 787 1092 788
rect 1086 783 1087 787
rect 1091 783 1092 787
rect 1086 782 1092 783
rect 1254 787 1260 788
rect 1254 783 1255 787
rect 1259 783 1260 787
rect 1254 782 1260 783
rect 1422 787 1428 788
rect 1422 783 1423 787
rect 1427 783 1428 787
rect 1422 782 1428 783
rect 1590 787 1596 788
rect 1590 783 1591 787
rect 1595 783 1596 787
rect 1590 782 1596 783
rect 2032 769 2034 797
rect 2072 785 2074 813
rect 2216 804 2218 813
rect 2344 804 2346 813
rect 2480 804 2482 813
rect 2624 804 2626 813
rect 2784 804 2786 813
rect 2960 804 2962 813
rect 3168 804 3170 813
rect 3392 804 3394 813
rect 3624 804 3626 813
rect 3864 804 3866 813
rect 2214 803 2220 804
rect 2214 799 2215 803
rect 2219 799 2220 803
rect 2214 798 2220 799
rect 2342 803 2348 804
rect 2342 799 2343 803
rect 2347 799 2348 803
rect 2342 798 2348 799
rect 2478 803 2484 804
rect 2478 799 2479 803
rect 2483 799 2484 803
rect 2478 798 2484 799
rect 2622 803 2628 804
rect 2622 799 2623 803
rect 2627 799 2628 803
rect 2622 798 2628 799
rect 2782 803 2788 804
rect 2782 799 2783 803
rect 2787 799 2788 803
rect 2782 798 2788 799
rect 2958 803 2964 804
rect 2958 799 2959 803
rect 2963 799 2964 803
rect 2958 798 2964 799
rect 3166 803 3172 804
rect 3166 799 3167 803
rect 3171 799 3172 803
rect 3166 798 3172 799
rect 3390 803 3396 804
rect 3390 799 3391 803
rect 3395 799 3396 803
rect 3390 798 3396 799
rect 3622 803 3628 804
rect 3622 799 3623 803
rect 3627 799 3628 803
rect 3622 798 3628 799
rect 3862 803 3868 804
rect 3862 799 3863 803
rect 3867 799 3868 803
rect 3862 798 3868 799
rect 3992 785 3994 813
rect 2070 784 2076 785
rect 2070 780 2071 784
rect 2075 780 2076 784
rect 2070 779 2076 780
rect 3990 784 3996 785
rect 3990 780 3991 784
rect 3995 780 3996 784
rect 3990 779 3996 780
rect 110 768 116 769
rect 110 764 111 768
rect 115 764 116 768
rect 110 763 116 764
rect 2030 768 2036 769
rect 2030 764 2031 768
rect 2035 764 2036 768
rect 2030 763 2036 764
rect 2070 767 2076 768
rect 2070 763 2071 767
rect 2075 763 2076 767
rect 3990 767 3996 768
rect 3990 763 3991 767
rect 3995 763 3996 767
rect 2070 762 2076 763
rect 2214 762 2220 763
rect 110 751 116 752
rect 110 747 111 751
rect 115 747 116 751
rect 2030 751 2036 752
rect 2030 747 2031 751
rect 2035 747 2036 751
rect 110 746 116 747
rect 278 746 284 747
rect 112 727 114 746
rect 278 742 279 746
rect 283 742 284 746
rect 278 741 284 742
rect 430 746 436 747
rect 430 742 431 746
rect 435 742 436 746
rect 430 741 436 742
rect 590 746 596 747
rect 590 742 591 746
rect 595 742 596 746
rect 590 741 596 742
rect 750 746 756 747
rect 750 742 751 746
rect 755 742 756 746
rect 750 741 756 742
rect 918 746 924 747
rect 918 742 919 746
rect 923 742 924 746
rect 918 741 924 742
rect 1086 746 1092 747
rect 1086 742 1087 746
rect 1091 742 1092 746
rect 1086 741 1092 742
rect 1254 746 1260 747
rect 1254 742 1255 746
rect 1259 742 1260 746
rect 1254 741 1260 742
rect 1422 746 1428 747
rect 1422 742 1423 746
rect 1427 742 1428 746
rect 1422 741 1428 742
rect 1590 746 1596 747
rect 2030 746 2036 747
rect 1590 742 1591 746
rect 1595 742 1596 746
rect 1590 741 1596 742
rect 280 727 282 741
rect 432 727 434 741
rect 592 727 594 741
rect 752 727 754 741
rect 920 727 922 741
rect 1088 727 1090 741
rect 1256 727 1258 741
rect 1424 727 1426 741
rect 1592 727 1594 741
rect 2032 727 2034 746
rect 2072 739 2074 762
rect 2214 758 2215 762
rect 2219 758 2220 762
rect 2214 757 2220 758
rect 2342 762 2348 763
rect 2342 758 2343 762
rect 2347 758 2348 762
rect 2342 757 2348 758
rect 2478 762 2484 763
rect 2478 758 2479 762
rect 2483 758 2484 762
rect 2478 757 2484 758
rect 2622 762 2628 763
rect 2622 758 2623 762
rect 2627 758 2628 762
rect 2622 757 2628 758
rect 2782 762 2788 763
rect 2782 758 2783 762
rect 2787 758 2788 762
rect 2782 757 2788 758
rect 2958 762 2964 763
rect 2958 758 2959 762
rect 2963 758 2964 762
rect 2958 757 2964 758
rect 3166 762 3172 763
rect 3166 758 3167 762
rect 3171 758 3172 762
rect 3166 757 3172 758
rect 3390 762 3396 763
rect 3390 758 3391 762
rect 3395 758 3396 762
rect 3390 757 3396 758
rect 3622 762 3628 763
rect 3622 758 3623 762
rect 3627 758 3628 762
rect 3622 757 3628 758
rect 3862 762 3868 763
rect 3990 762 3996 763
rect 3862 758 3863 762
rect 3867 758 3868 762
rect 3862 757 3868 758
rect 2216 739 2218 757
rect 2344 739 2346 757
rect 2480 739 2482 757
rect 2624 739 2626 757
rect 2784 739 2786 757
rect 2960 739 2962 757
rect 3168 739 3170 757
rect 3392 739 3394 757
rect 3624 739 3626 757
rect 3864 739 3866 757
rect 3992 739 3994 762
rect 2071 738 2075 739
rect 2071 733 2075 734
rect 2111 738 2115 739
rect 2111 733 2115 734
rect 2215 738 2219 739
rect 2215 733 2219 734
rect 2247 738 2251 739
rect 2247 733 2251 734
rect 2343 738 2347 739
rect 2343 733 2347 734
rect 2423 738 2427 739
rect 2423 733 2427 734
rect 2479 738 2483 739
rect 2479 733 2483 734
rect 2599 738 2603 739
rect 2599 733 2603 734
rect 2623 738 2627 739
rect 2623 733 2627 734
rect 2783 738 2787 739
rect 2783 733 2787 734
rect 2959 738 2963 739
rect 2959 733 2963 734
rect 2967 738 2971 739
rect 2967 733 2971 734
rect 3151 738 3155 739
rect 3151 733 3155 734
rect 3167 738 3171 739
rect 3167 733 3171 734
rect 3335 738 3339 739
rect 3335 733 3339 734
rect 3391 738 3395 739
rect 3391 733 3395 734
rect 3519 738 3523 739
rect 3519 733 3523 734
rect 3623 738 3627 739
rect 3623 733 3627 734
rect 3703 738 3707 739
rect 3703 733 3707 734
rect 3863 738 3867 739
rect 3863 733 3867 734
rect 3895 738 3899 739
rect 3895 733 3899 734
rect 3991 738 3995 739
rect 3991 733 3995 734
rect 111 726 115 727
rect 111 721 115 722
rect 151 726 155 727
rect 151 721 155 722
rect 271 726 275 727
rect 271 721 275 722
rect 279 726 283 727
rect 279 721 283 722
rect 423 726 427 727
rect 423 721 427 722
rect 431 726 435 727
rect 431 721 435 722
rect 575 726 579 727
rect 575 721 579 722
rect 591 726 595 727
rect 591 721 595 722
rect 735 726 739 727
rect 735 721 739 722
rect 751 726 755 727
rect 751 721 755 722
rect 887 726 891 727
rect 887 721 891 722
rect 919 726 923 727
rect 919 721 923 722
rect 1039 726 1043 727
rect 1039 721 1043 722
rect 1087 726 1091 727
rect 1087 721 1091 722
rect 1191 726 1195 727
rect 1191 721 1195 722
rect 1255 726 1259 727
rect 1255 721 1259 722
rect 1343 726 1347 727
rect 1343 721 1347 722
rect 1423 726 1427 727
rect 1423 721 1427 722
rect 1495 726 1499 727
rect 1495 721 1499 722
rect 1591 726 1595 727
rect 1591 721 1595 722
rect 2031 726 2035 727
rect 2031 721 2035 722
rect 112 706 114 721
rect 152 711 154 721
rect 272 711 274 721
rect 424 711 426 721
rect 576 711 578 721
rect 736 711 738 721
rect 888 711 890 721
rect 1040 711 1042 721
rect 1192 711 1194 721
rect 1344 711 1346 721
rect 1496 711 1498 721
rect 150 710 156 711
rect 150 706 151 710
rect 155 706 156 710
rect 110 705 116 706
rect 150 705 156 706
rect 270 710 276 711
rect 270 706 271 710
rect 275 706 276 710
rect 270 705 276 706
rect 422 710 428 711
rect 422 706 423 710
rect 427 706 428 710
rect 422 705 428 706
rect 574 710 580 711
rect 574 706 575 710
rect 579 706 580 710
rect 574 705 580 706
rect 734 710 740 711
rect 734 706 735 710
rect 739 706 740 710
rect 734 705 740 706
rect 886 710 892 711
rect 886 706 887 710
rect 891 706 892 710
rect 886 705 892 706
rect 1038 710 1044 711
rect 1038 706 1039 710
rect 1043 706 1044 710
rect 1038 705 1044 706
rect 1190 710 1196 711
rect 1190 706 1191 710
rect 1195 706 1196 710
rect 1190 705 1196 706
rect 1342 710 1348 711
rect 1342 706 1343 710
rect 1347 706 1348 710
rect 1342 705 1348 706
rect 1494 710 1500 711
rect 1494 706 1495 710
rect 1499 706 1500 710
rect 2032 706 2034 721
rect 2072 718 2074 733
rect 2112 723 2114 733
rect 2248 723 2250 733
rect 2424 723 2426 733
rect 2600 723 2602 733
rect 2784 723 2786 733
rect 2968 723 2970 733
rect 3152 723 3154 733
rect 3336 723 3338 733
rect 3520 723 3522 733
rect 3704 723 3706 733
rect 3896 723 3898 733
rect 2110 722 2116 723
rect 2110 718 2111 722
rect 2115 718 2116 722
rect 2070 717 2076 718
rect 2110 717 2116 718
rect 2246 722 2252 723
rect 2246 718 2247 722
rect 2251 718 2252 722
rect 2246 717 2252 718
rect 2422 722 2428 723
rect 2422 718 2423 722
rect 2427 718 2428 722
rect 2422 717 2428 718
rect 2598 722 2604 723
rect 2598 718 2599 722
rect 2603 718 2604 722
rect 2598 717 2604 718
rect 2782 722 2788 723
rect 2782 718 2783 722
rect 2787 718 2788 722
rect 2782 717 2788 718
rect 2966 722 2972 723
rect 2966 718 2967 722
rect 2971 718 2972 722
rect 2966 717 2972 718
rect 3150 722 3156 723
rect 3150 718 3151 722
rect 3155 718 3156 722
rect 3150 717 3156 718
rect 3334 722 3340 723
rect 3334 718 3335 722
rect 3339 718 3340 722
rect 3334 717 3340 718
rect 3518 722 3524 723
rect 3518 718 3519 722
rect 3523 718 3524 722
rect 3518 717 3524 718
rect 3702 722 3708 723
rect 3702 718 3703 722
rect 3707 718 3708 722
rect 3702 717 3708 718
rect 3894 722 3900 723
rect 3894 718 3895 722
rect 3899 718 3900 722
rect 3992 718 3994 733
rect 3894 717 3900 718
rect 3990 717 3996 718
rect 2070 713 2071 717
rect 2075 713 2076 717
rect 2070 712 2076 713
rect 3990 713 3991 717
rect 3995 713 3996 717
rect 3990 712 3996 713
rect 1494 705 1500 706
rect 2030 705 2036 706
rect 110 701 111 705
rect 115 701 116 705
rect 110 700 116 701
rect 2030 701 2031 705
rect 2035 701 2036 705
rect 2030 700 2036 701
rect 2070 700 2076 701
rect 2070 696 2071 700
rect 2075 696 2076 700
rect 2070 695 2076 696
rect 3990 700 3996 701
rect 3990 696 3991 700
rect 3995 696 3996 700
rect 3990 695 3996 696
rect 110 688 116 689
rect 110 684 111 688
rect 115 684 116 688
rect 110 683 116 684
rect 2030 688 2036 689
rect 2030 684 2031 688
rect 2035 684 2036 688
rect 2030 683 2036 684
rect 112 647 114 683
rect 150 669 156 670
rect 150 665 151 669
rect 155 665 156 669
rect 150 664 156 665
rect 270 669 276 670
rect 270 665 271 669
rect 275 665 276 669
rect 270 664 276 665
rect 422 669 428 670
rect 422 665 423 669
rect 427 665 428 669
rect 422 664 428 665
rect 574 669 580 670
rect 574 665 575 669
rect 579 665 580 669
rect 574 664 580 665
rect 734 669 740 670
rect 734 665 735 669
rect 739 665 740 669
rect 734 664 740 665
rect 886 669 892 670
rect 886 665 887 669
rect 891 665 892 669
rect 886 664 892 665
rect 1038 669 1044 670
rect 1038 665 1039 669
rect 1043 665 1044 669
rect 1038 664 1044 665
rect 1190 669 1196 670
rect 1190 665 1191 669
rect 1195 665 1196 669
rect 1190 664 1196 665
rect 1342 669 1348 670
rect 1342 665 1343 669
rect 1347 665 1348 669
rect 1342 664 1348 665
rect 1494 669 1500 670
rect 1494 665 1495 669
rect 1499 665 1500 669
rect 1494 664 1500 665
rect 152 647 154 664
rect 272 647 274 664
rect 424 647 426 664
rect 576 647 578 664
rect 736 647 738 664
rect 888 647 890 664
rect 1040 647 1042 664
rect 1192 647 1194 664
rect 1344 647 1346 664
rect 1496 647 1498 664
rect 2032 647 2034 683
rect 2072 663 2074 695
rect 2110 681 2116 682
rect 2110 677 2111 681
rect 2115 677 2116 681
rect 2110 676 2116 677
rect 2246 681 2252 682
rect 2246 677 2247 681
rect 2251 677 2252 681
rect 2246 676 2252 677
rect 2422 681 2428 682
rect 2422 677 2423 681
rect 2427 677 2428 681
rect 2422 676 2428 677
rect 2598 681 2604 682
rect 2598 677 2599 681
rect 2603 677 2604 681
rect 2598 676 2604 677
rect 2782 681 2788 682
rect 2782 677 2783 681
rect 2787 677 2788 681
rect 2782 676 2788 677
rect 2966 681 2972 682
rect 2966 677 2967 681
rect 2971 677 2972 681
rect 2966 676 2972 677
rect 3150 681 3156 682
rect 3150 677 3151 681
rect 3155 677 3156 681
rect 3150 676 3156 677
rect 3334 681 3340 682
rect 3334 677 3335 681
rect 3339 677 3340 681
rect 3334 676 3340 677
rect 3518 681 3524 682
rect 3518 677 3519 681
rect 3523 677 3524 681
rect 3518 676 3524 677
rect 3702 681 3708 682
rect 3702 677 3703 681
rect 3707 677 3708 681
rect 3702 676 3708 677
rect 3894 681 3900 682
rect 3894 677 3895 681
rect 3899 677 3900 681
rect 3894 676 3900 677
rect 2112 663 2114 676
rect 2248 663 2250 676
rect 2424 663 2426 676
rect 2600 663 2602 676
rect 2784 663 2786 676
rect 2968 663 2970 676
rect 3152 663 3154 676
rect 3336 663 3338 676
rect 3520 663 3522 676
rect 3704 663 3706 676
rect 3896 663 3898 676
rect 3992 663 3994 695
rect 2071 662 2075 663
rect 2071 657 2075 658
rect 2111 662 2115 663
rect 2111 657 2115 658
rect 2247 662 2251 663
rect 2247 657 2251 658
rect 2375 662 2379 663
rect 2375 657 2379 658
rect 2423 662 2427 663
rect 2423 657 2427 658
rect 2599 662 2603 663
rect 2599 657 2603 658
rect 2655 662 2659 663
rect 2655 657 2659 658
rect 2783 662 2787 663
rect 2783 657 2787 658
rect 2919 662 2923 663
rect 2919 657 2923 658
rect 2967 662 2971 663
rect 2967 657 2971 658
rect 3151 662 3155 663
rect 3151 657 3155 658
rect 3175 662 3179 663
rect 3175 657 3179 658
rect 3335 662 3339 663
rect 3335 657 3339 658
rect 3423 662 3427 663
rect 3423 657 3427 658
rect 3519 662 3523 663
rect 3519 657 3523 658
rect 3671 662 3675 663
rect 3671 657 3675 658
rect 3703 662 3707 663
rect 3703 657 3707 658
rect 3895 662 3899 663
rect 3895 657 3899 658
rect 3991 662 3995 663
rect 3991 657 3995 658
rect 111 646 115 647
rect 111 641 115 642
rect 151 646 155 647
rect 151 641 155 642
rect 255 646 259 647
rect 255 641 259 642
rect 271 646 275 647
rect 271 641 275 642
rect 391 646 395 647
rect 391 641 395 642
rect 423 646 427 647
rect 423 641 427 642
rect 527 646 531 647
rect 527 641 531 642
rect 575 646 579 647
rect 575 641 579 642
rect 663 646 667 647
rect 663 641 667 642
rect 735 646 739 647
rect 735 641 739 642
rect 807 646 811 647
rect 807 641 811 642
rect 887 646 891 647
rect 887 641 891 642
rect 959 646 963 647
rect 959 641 963 642
rect 1039 646 1043 647
rect 1039 641 1043 642
rect 1119 646 1123 647
rect 1119 641 1123 642
rect 1191 646 1195 647
rect 1191 641 1195 642
rect 1287 646 1291 647
rect 1287 641 1291 642
rect 1343 646 1347 647
rect 1343 641 1347 642
rect 1455 646 1459 647
rect 1455 641 1459 642
rect 1495 646 1499 647
rect 1495 641 1499 642
rect 1623 646 1627 647
rect 1623 641 1627 642
rect 1791 646 1795 647
rect 1791 641 1795 642
rect 1935 646 1939 647
rect 1935 641 1939 642
rect 2031 646 2035 647
rect 2031 641 2035 642
rect 112 613 114 641
rect 152 632 154 641
rect 256 632 258 641
rect 392 632 394 641
rect 528 632 530 641
rect 664 632 666 641
rect 808 632 810 641
rect 960 632 962 641
rect 1120 632 1122 641
rect 1288 632 1290 641
rect 1456 632 1458 641
rect 1624 632 1626 641
rect 1792 632 1794 641
rect 1936 632 1938 641
rect 150 631 156 632
rect 150 627 151 631
rect 155 627 156 631
rect 150 626 156 627
rect 254 631 260 632
rect 254 627 255 631
rect 259 627 260 631
rect 254 626 260 627
rect 390 631 396 632
rect 390 627 391 631
rect 395 627 396 631
rect 390 626 396 627
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 662 631 668 632
rect 662 627 663 631
rect 667 627 668 631
rect 662 626 668 627
rect 806 631 812 632
rect 806 627 807 631
rect 811 627 812 631
rect 806 626 812 627
rect 958 631 964 632
rect 958 627 959 631
rect 963 627 964 631
rect 958 626 964 627
rect 1118 631 1124 632
rect 1118 627 1119 631
rect 1123 627 1124 631
rect 1118 626 1124 627
rect 1286 631 1292 632
rect 1286 627 1287 631
rect 1291 627 1292 631
rect 1286 626 1292 627
rect 1454 631 1460 632
rect 1454 627 1455 631
rect 1459 627 1460 631
rect 1454 626 1460 627
rect 1622 631 1628 632
rect 1622 627 1623 631
rect 1627 627 1628 631
rect 1622 626 1628 627
rect 1790 631 1796 632
rect 1790 627 1791 631
rect 1795 627 1796 631
rect 1790 626 1796 627
rect 1934 631 1940 632
rect 1934 627 1935 631
rect 1939 627 1940 631
rect 1934 626 1940 627
rect 2032 613 2034 641
rect 2072 629 2074 657
rect 2112 648 2114 657
rect 2376 648 2378 657
rect 2656 648 2658 657
rect 2920 648 2922 657
rect 3176 648 3178 657
rect 3424 648 3426 657
rect 3672 648 3674 657
rect 3896 648 3898 657
rect 2110 647 2116 648
rect 2110 643 2111 647
rect 2115 643 2116 647
rect 2110 642 2116 643
rect 2374 647 2380 648
rect 2374 643 2375 647
rect 2379 643 2380 647
rect 2374 642 2380 643
rect 2654 647 2660 648
rect 2654 643 2655 647
rect 2659 643 2660 647
rect 2654 642 2660 643
rect 2918 647 2924 648
rect 2918 643 2919 647
rect 2923 643 2924 647
rect 2918 642 2924 643
rect 3174 647 3180 648
rect 3174 643 3175 647
rect 3179 643 3180 647
rect 3174 642 3180 643
rect 3422 647 3428 648
rect 3422 643 3423 647
rect 3427 643 3428 647
rect 3422 642 3428 643
rect 3670 647 3676 648
rect 3670 643 3671 647
rect 3675 643 3676 647
rect 3670 642 3676 643
rect 3894 647 3900 648
rect 3894 643 3895 647
rect 3899 643 3900 647
rect 3894 642 3900 643
rect 3992 629 3994 657
rect 2070 628 2076 629
rect 2070 624 2071 628
rect 2075 624 2076 628
rect 2070 623 2076 624
rect 3990 628 3996 629
rect 3990 624 3991 628
rect 3995 624 3996 628
rect 3990 623 3996 624
rect 110 612 116 613
rect 110 608 111 612
rect 115 608 116 612
rect 110 607 116 608
rect 2030 612 2036 613
rect 2030 608 2031 612
rect 2035 608 2036 612
rect 2030 607 2036 608
rect 2070 611 2076 612
rect 2070 607 2071 611
rect 2075 607 2076 611
rect 3990 611 3996 612
rect 3990 607 3991 611
rect 3995 607 3996 611
rect 2070 606 2076 607
rect 2110 606 2116 607
rect 110 595 116 596
rect 110 591 111 595
rect 115 591 116 595
rect 2030 595 2036 596
rect 2030 591 2031 595
rect 2035 591 2036 595
rect 110 590 116 591
rect 150 590 156 591
rect 112 563 114 590
rect 150 586 151 590
rect 155 586 156 590
rect 150 585 156 586
rect 254 590 260 591
rect 254 586 255 590
rect 259 586 260 590
rect 254 585 260 586
rect 390 590 396 591
rect 390 586 391 590
rect 395 586 396 590
rect 390 585 396 586
rect 526 590 532 591
rect 526 586 527 590
rect 531 586 532 590
rect 526 585 532 586
rect 662 590 668 591
rect 662 586 663 590
rect 667 586 668 590
rect 662 585 668 586
rect 806 590 812 591
rect 806 586 807 590
rect 811 586 812 590
rect 806 585 812 586
rect 958 590 964 591
rect 958 586 959 590
rect 963 586 964 590
rect 958 585 964 586
rect 1118 590 1124 591
rect 1118 586 1119 590
rect 1123 586 1124 590
rect 1118 585 1124 586
rect 1286 590 1292 591
rect 1286 586 1287 590
rect 1291 586 1292 590
rect 1286 585 1292 586
rect 1454 590 1460 591
rect 1454 586 1455 590
rect 1459 586 1460 590
rect 1454 585 1460 586
rect 1622 590 1628 591
rect 1622 586 1623 590
rect 1627 586 1628 590
rect 1622 585 1628 586
rect 1790 590 1796 591
rect 1790 586 1791 590
rect 1795 586 1796 590
rect 1790 585 1796 586
rect 1934 590 1940 591
rect 2030 590 2036 591
rect 1934 586 1935 590
rect 1939 586 1940 590
rect 1934 585 1940 586
rect 152 563 154 585
rect 256 563 258 585
rect 392 563 394 585
rect 528 563 530 585
rect 664 563 666 585
rect 808 563 810 585
rect 960 563 962 585
rect 1120 563 1122 585
rect 1288 563 1290 585
rect 1456 563 1458 585
rect 1624 563 1626 585
rect 1792 563 1794 585
rect 1936 563 1938 585
rect 2032 563 2034 590
rect 2072 579 2074 606
rect 2110 602 2111 606
rect 2115 602 2116 606
rect 2110 601 2116 602
rect 2374 606 2380 607
rect 2374 602 2375 606
rect 2379 602 2380 606
rect 2374 601 2380 602
rect 2654 606 2660 607
rect 2654 602 2655 606
rect 2659 602 2660 606
rect 2654 601 2660 602
rect 2918 606 2924 607
rect 2918 602 2919 606
rect 2923 602 2924 606
rect 2918 601 2924 602
rect 3174 606 3180 607
rect 3174 602 3175 606
rect 3179 602 3180 606
rect 3174 601 3180 602
rect 3422 606 3428 607
rect 3422 602 3423 606
rect 3427 602 3428 606
rect 3422 601 3428 602
rect 3670 606 3676 607
rect 3670 602 3671 606
rect 3675 602 3676 606
rect 3670 601 3676 602
rect 3894 606 3900 607
rect 3990 606 3996 607
rect 3894 602 3895 606
rect 3899 602 3900 606
rect 3894 601 3900 602
rect 2112 579 2114 601
rect 2376 579 2378 601
rect 2656 579 2658 601
rect 2920 579 2922 601
rect 3176 579 3178 601
rect 3424 579 3426 601
rect 3672 579 3674 601
rect 3896 579 3898 601
rect 3992 579 3994 606
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2111 578 2115 579
rect 2111 573 2115 574
rect 2215 578 2219 579
rect 2215 573 2219 574
rect 2351 578 2355 579
rect 2351 573 2355 574
rect 2375 578 2379 579
rect 2375 573 2379 574
rect 2487 578 2491 579
rect 2487 573 2491 574
rect 2631 578 2635 579
rect 2631 573 2635 574
rect 2655 578 2659 579
rect 2655 573 2659 574
rect 2791 578 2795 579
rect 2791 573 2795 574
rect 2919 578 2923 579
rect 2919 573 2923 574
rect 2975 578 2979 579
rect 2975 573 2979 574
rect 3175 578 3179 579
rect 3175 573 3179 574
rect 3191 578 3195 579
rect 3191 573 3195 574
rect 3423 578 3427 579
rect 3423 573 3427 574
rect 3671 578 3675 579
rect 3671 573 3675 574
rect 3895 578 3899 579
rect 3895 573 3899 574
rect 3991 578 3995 579
rect 3991 573 3995 574
rect 111 562 115 563
rect 111 557 115 558
rect 151 562 155 563
rect 151 557 155 558
rect 207 562 211 563
rect 207 557 211 558
rect 255 562 259 563
rect 255 557 259 558
rect 327 562 331 563
rect 327 557 331 558
rect 391 562 395 563
rect 391 557 395 558
rect 447 562 451 563
rect 447 557 451 558
rect 527 562 531 563
rect 527 557 531 558
rect 567 562 571 563
rect 567 557 571 558
rect 663 562 667 563
rect 663 557 667 558
rect 687 562 691 563
rect 687 557 691 558
rect 799 562 803 563
rect 799 557 803 558
rect 807 562 811 563
rect 807 557 811 558
rect 911 562 915 563
rect 911 557 915 558
rect 959 562 963 563
rect 959 557 963 558
rect 1031 562 1035 563
rect 1031 557 1035 558
rect 1119 562 1123 563
rect 1119 557 1123 558
rect 1151 562 1155 563
rect 1151 557 1155 558
rect 1271 562 1275 563
rect 1271 557 1275 558
rect 1287 562 1291 563
rect 1287 557 1291 558
rect 1455 562 1459 563
rect 1455 557 1459 558
rect 1623 562 1627 563
rect 1623 557 1627 558
rect 1791 562 1795 563
rect 1791 557 1795 558
rect 1935 562 1939 563
rect 1935 557 1939 558
rect 2031 562 2035 563
rect 2072 558 2074 573
rect 2112 563 2114 573
rect 2216 563 2218 573
rect 2352 563 2354 573
rect 2488 563 2490 573
rect 2632 563 2634 573
rect 2792 563 2794 573
rect 2976 563 2978 573
rect 3192 563 3194 573
rect 3424 563 3426 573
rect 3672 563 3674 573
rect 3896 563 3898 573
rect 2110 562 2116 563
rect 2110 558 2111 562
rect 2115 558 2116 562
rect 2031 557 2035 558
rect 2070 557 2076 558
rect 2110 557 2116 558
rect 2214 562 2220 563
rect 2214 558 2215 562
rect 2219 558 2220 562
rect 2214 557 2220 558
rect 2350 562 2356 563
rect 2350 558 2351 562
rect 2355 558 2356 562
rect 2350 557 2356 558
rect 2486 562 2492 563
rect 2486 558 2487 562
rect 2491 558 2492 562
rect 2486 557 2492 558
rect 2630 562 2636 563
rect 2630 558 2631 562
rect 2635 558 2636 562
rect 2630 557 2636 558
rect 2790 562 2796 563
rect 2790 558 2791 562
rect 2795 558 2796 562
rect 2790 557 2796 558
rect 2974 562 2980 563
rect 2974 558 2975 562
rect 2979 558 2980 562
rect 2974 557 2980 558
rect 3190 562 3196 563
rect 3190 558 3191 562
rect 3195 558 3196 562
rect 3190 557 3196 558
rect 3422 562 3428 563
rect 3422 558 3423 562
rect 3427 558 3428 562
rect 3422 557 3428 558
rect 3670 562 3676 563
rect 3670 558 3671 562
rect 3675 558 3676 562
rect 3670 557 3676 558
rect 3894 562 3900 563
rect 3894 558 3895 562
rect 3899 558 3900 562
rect 3992 558 3994 573
rect 3894 557 3900 558
rect 3990 557 3996 558
rect 112 542 114 557
rect 208 547 210 557
rect 328 547 330 557
rect 448 547 450 557
rect 568 547 570 557
rect 688 547 690 557
rect 800 547 802 557
rect 912 547 914 557
rect 1032 547 1034 557
rect 1152 547 1154 557
rect 1272 547 1274 557
rect 206 546 212 547
rect 206 542 207 546
rect 211 542 212 546
rect 110 541 116 542
rect 206 541 212 542
rect 326 546 332 547
rect 326 542 327 546
rect 331 542 332 546
rect 326 541 332 542
rect 446 546 452 547
rect 446 542 447 546
rect 451 542 452 546
rect 446 541 452 542
rect 566 546 572 547
rect 566 542 567 546
rect 571 542 572 546
rect 566 541 572 542
rect 686 546 692 547
rect 686 542 687 546
rect 691 542 692 546
rect 686 541 692 542
rect 798 546 804 547
rect 798 542 799 546
rect 803 542 804 546
rect 798 541 804 542
rect 910 546 916 547
rect 910 542 911 546
rect 915 542 916 546
rect 910 541 916 542
rect 1030 546 1036 547
rect 1030 542 1031 546
rect 1035 542 1036 546
rect 1030 541 1036 542
rect 1150 546 1156 547
rect 1150 542 1151 546
rect 1155 542 1156 546
rect 1150 541 1156 542
rect 1270 546 1276 547
rect 1270 542 1271 546
rect 1275 542 1276 546
rect 2032 542 2034 557
rect 2070 553 2071 557
rect 2075 553 2076 557
rect 2070 552 2076 553
rect 3990 553 3991 557
rect 3995 553 3996 557
rect 3990 552 3996 553
rect 1270 541 1276 542
rect 2030 541 2036 542
rect 110 537 111 541
rect 115 537 116 541
rect 110 536 116 537
rect 2030 537 2031 541
rect 2035 537 2036 541
rect 2030 536 2036 537
rect 2070 540 2076 541
rect 2070 536 2071 540
rect 2075 536 2076 540
rect 2070 535 2076 536
rect 3990 540 3996 541
rect 3990 536 3991 540
rect 3995 536 3996 540
rect 3990 535 3996 536
rect 110 524 116 525
rect 110 520 111 524
rect 115 520 116 524
rect 110 519 116 520
rect 2030 524 2036 525
rect 2030 520 2031 524
rect 2035 520 2036 524
rect 2030 519 2036 520
rect 112 483 114 519
rect 206 505 212 506
rect 206 501 207 505
rect 211 501 212 505
rect 206 500 212 501
rect 326 505 332 506
rect 326 501 327 505
rect 331 501 332 505
rect 326 500 332 501
rect 446 505 452 506
rect 446 501 447 505
rect 451 501 452 505
rect 446 500 452 501
rect 566 505 572 506
rect 566 501 567 505
rect 571 501 572 505
rect 566 500 572 501
rect 686 505 692 506
rect 686 501 687 505
rect 691 501 692 505
rect 686 500 692 501
rect 798 505 804 506
rect 798 501 799 505
rect 803 501 804 505
rect 798 500 804 501
rect 910 505 916 506
rect 910 501 911 505
rect 915 501 916 505
rect 910 500 916 501
rect 1030 505 1036 506
rect 1030 501 1031 505
rect 1035 501 1036 505
rect 1030 500 1036 501
rect 1150 505 1156 506
rect 1150 501 1151 505
rect 1155 501 1156 505
rect 1150 500 1156 501
rect 1270 505 1276 506
rect 1270 501 1271 505
rect 1275 501 1276 505
rect 1270 500 1276 501
rect 208 483 210 500
rect 328 483 330 500
rect 448 483 450 500
rect 568 483 570 500
rect 688 483 690 500
rect 800 483 802 500
rect 912 483 914 500
rect 1032 483 1034 500
rect 1152 483 1154 500
rect 1272 483 1274 500
rect 2032 483 2034 519
rect 2072 503 2074 535
rect 2110 521 2116 522
rect 2110 517 2111 521
rect 2115 517 2116 521
rect 2110 516 2116 517
rect 2214 521 2220 522
rect 2214 517 2215 521
rect 2219 517 2220 521
rect 2214 516 2220 517
rect 2350 521 2356 522
rect 2350 517 2351 521
rect 2355 517 2356 521
rect 2350 516 2356 517
rect 2486 521 2492 522
rect 2486 517 2487 521
rect 2491 517 2492 521
rect 2486 516 2492 517
rect 2630 521 2636 522
rect 2630 517 2631 521
rect 2635 517 2636 521
rect 2630 516 2636 517
rect 2790 521 2796 522
rect 2790 517 2791 521
rect 2795 517 2796 521
rect 2790 516 2796 517
rect 2974 521 2980 522
rect 2974 517 2975 521
rect 2979 517 2980 521
rect 2974 516 2980 517
rect 3190 521 3196 522
rect 3190 517 3191 521
rect 3195 517 3196 521
rect 3190 516 3196 517
rect 3422 521 3428 522
rect 3422 517 3423 521
rect 3427 517 3428 521
rect 3422 516 3428 517
rect 3670 521 3676 522
rect 3670 517 3671 521
rect 3675 517 3676 521
rect 3670 516 3676 517
rect 3894 521 3900 522
rect 3894 517 3895 521
rect 3899 517 3900 521
rect 3894 516 3900 517
rect 2112 503 2114 516
rect 2216 503 2218 516
rect 2352 503 2354 516
rect 2488 503 2490 516
rect 2632 503 2634 516
rect 2792 503 2794 516
rect 2976 503 2978 516
rect 3192 503 3194 516
rect 3424 503 3426 516
rect 3672 503 3674 516
rect 3896 503 3898 516
rect 3992 503 3994 535
rect 2071 502 2075 503
rect 2071 497 2075 498
rect 2111 502 2115 503
rect 2111 497 2115 498
rect 2215 502 2219 503
rect 2215 497 2219 498
rect 2351 502 2355 503
rect 2351 497 2355 498
rect 2423 502 2427 503
rect 2423 497 2427 498
rect 2487 502 2491 503
rect 2487 497 2491 498
rect 2527 502 2531 503
rect 2527 497 2531 498
rect 2631 502 2635 503
rect 2631 497 2635 498
rect 2743 502 2747 503
rect 2743 497 2747 498
rect 2791 502 2795 503
rect 2791 497 2795 498
rect 2871 502 2875 503
rect 2871 497 2875 498
rect 2975 502 2979 503
rect 2975 497 2979 498
rect 3031 502 3035 503
rect 3031 497 3035 498
rect 3191 502 3195 503
rect 3191 497 3195 498
rect 3223 502 3227 503
rect 3223 497 3227 498
rect 3423 502 3427 503
rect 3423 497 3427 498
rect 3447 502 3451 503
rect 3447 497 3451 498
rect 3671 502 3675 503
rect 3671 497 3675 498
rect 3679 502 3683 503
rect 3679 497 3683 498
rect 3895 502 3899 503
rect 3895 497 3899 498
rect 3991 502 3995 503
rect 3991 497 3995 498
rect 111 482 115 483
rect 111 477 115 478
rect 207 482 211 483
rect 207 477 211 478
rect 327 482 331 483
rect 327 477 331 478
rect 439 482 443 483
rect 439 477 443 478
rect 447 482 451 483
rect 447 477 451 478
rect 543 482 547 483
rect 543 477 547 478
rect 567 482 571 483
rect 567 477 571 478
rect 647 482 651 483
rect 647 477 651 478
rect 687 482 691 483
rect 687 477 691 478
rect 751 482 755 483
rect 751 477 755 478
rect 799 482 803 483
rect 799 477 803 478
rect 855 482 859 483
rect 855 477 859 478
rect 911 482 915 483
rect 911 477 915 478
rect 959 482 963 483
rect 959 477 963 478
rect 1031 482 1035 483
rect 1031 477 1035 478
rect 1063 482 1067 483
rect 1063 477 1067 478
rect 1151 482 1155 483
rect 1151 477 1155 478
rect 1167 482 1171 483
rect 1167 477 1171 478
rect 1271 482 1275 483
rect 1271 477 1275 478
rect 1375 482 1379 483
rect 1375 477 1379 478
rect 2031 482 2035 483
rect 2031 477 2035 478
rect 112 449 114 477
rect 440 468 442 477
rect 544 468 546 477
rect 648 468 650 477
rect 752 468 754 477
rect 856 468 858 477
rect 960 468 962 477
rect 1064 468 1066 477
rect 1168 468 1170 477
rect 1272 468 1274 477
rect 1376 468 1378 477
rect 438 467 444 468
rect 438 463 439 467
rect 443 463 444 467
rect 438 462 444 463
rect 542 467 548 468
rect 542 463 543 467
rect 547 463 548 467
rect 542 462 548 463
rect 646 467 652 468
rect 646 463 647 467
rect 651 463 652 467
rect 646 462 652 463
rect 750 467 756 468
rect 750 463 751 467
rect 755 463 756 467
rect 750 462 756 463
rect 854 467 860 468
rect 854 463 855 467
rect 859 463 860 467
rect 854 462 860 463
rect 958 467 964 468
rect 958 463 959 467
rect 963 463 964 467
rect 958 462 964 463
rect 1062 467 1068 468
rect 1062 463 1063 467
rect 1067 463 1068 467
rect 1062 462 1068 463
rect 1166 467 1172 468
rect 1166 463 1167 467
rect 1171 463 1172 467
rect 1166 462 1172 463
rect 1270 467 1276 468
rect 1270 463 1271 467
rect 1275 463 1276 467
rect 1270 462 1276 463
rect 1374 467 1380 468
rect 1374 463 1375 467
rect 1379 463 1380 467
rect 1374 462 1380 463
rect 2032 449 2034 477
rect 2072 469 2074 497
rect 2424 488 2426 497
rect 2528 488 2530 497
rect 2632 488 2634 497
rect 2744 488 2746 497
rect 2872 488 2874 497
rect 3032 488 3034 497
rect 3224 488 3226 497
rect 3448 488 3450 497
rect 3680 488 3682 497
rect 3896 488 3898 497
rect 2422 487 2428 488
rect 2422 483 2423 487
rect 2427 483 2428 487
rect 2422 482 2428 483
rect 2526 487 2532 488
rect 2526 483 2527 487
rect 2531 483 2532 487
rect 2526 482 2532 483
rect 2630 487 2636 488
rect 2630 483 2631 487
rect 2635 483 2636 487
rect 2630 482 2636 483
rect 2742 487 2748 488
rect 2742 483 2743 487
rect 2747 483 2748 487
rect 2742 482 2748 483
rect 2870 487 2876 488
rect 2870 483 2871 487
rect 2875 483 2876 487
rect 2870 482 2876 483
rect 3030 487 3036 488
rect 3030 483 3031 487
rect 3035 483 3036 487
rect 3030 482 3036 483
rect 3222 487 3228 488
rect 3222 483 3223 487
rect 3227 483 3228 487
rect 3222 482 3228 483
rect 3446 487 3452 488
rect 3446 483 3447 487
rect 3451 483 3452 487
rect 3446 482 3452 483
rect 3678 487 3684 488
rect 3678 483 3679 487
rect 3683 483 3684 487
rect 3678 482 3684 483
rect 3894 487 3900 488
rect 3894 483 3895 487
rect 3899 483 3900 487
rect 3894 482 3900 483
rect 3992 469 3994 497
rect 2070 468 2076 469
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 3990 468 3996 469
rect 3990 464 3991 468
rect 3995 464 3996 468
rect 3990 463 3996 464
rect 2070 451 2076 452
rect 110 448 116 449
rect 110 444 111 448
rect 115 444 116 448
rect 110 443 116 444
rect 2030 448 2036 449
rect 2030 444 2031 448
rect 2035 444 2036 448
rect 2070 447 2071 451
rect 2075 447 2076 451
rect 3990 451 3996 452
rect 3990 447 3991 451
rect 3995 447 3996 451
rect 2070 446 2076 447
rect 2422 446 2428 447
rect 2030 443 2036 444
rect 110 431 116 432
rect 110 427 111 431
rect 115 427 116 431
rect 2030 431 2036 432
rect 2030 427 2031 431
rect 2035 427 2036 431
rect 2072 427 2074 446
rect 2422 442 2423 446
rect 2427 442 2428 446
rect 2422 441 2428 442
rect 2526 446 2532 447
rect 2526 442 2527 446
rect 2531 442 2532 446
rect 2526 441 2532 442
rect 2630 446 2636 447
rect 2630 442 2631 446
rect 2635 442 2636 446
rect 2630 441 2636 442
rect 2742 446 2748 447
rect 2742 442 2743 446
rect 2747 442 2748 446
rect 2742 441 2748 442
rect 2870 446 2876 447
rect 2870 442 2871 446
rect 2875 442 2876 446
rect 2870 441 2876 442
rect 3030 446 3036 447
rect 3030 442 3031 446
rect 3035 442 3036 446
rect 3030 441 3036 442
rect 3222 446 3228 447
rect 3222 442 3223 446
rect 3227 442 3228 446
rect 3222 441 3228 442
rect 3446 446 3452 447
rect 3446 442 3447 446
rect 3451 442 3452 446
rect 3446 441 3452 442
rect 3678 446 3684 447
rect 3678 442 3679 446
rect 3683 442 3684 446
rect 3678 441 3684 442
rect 3894 446 3900 447
rect 3990 446 3996 447
rect 3894 442 3895 446
rect 3899 442 3900 446
rect 3894 441 3900 442
rect 2424 427 2426 441
rect 2528 427 2530 441
rect 2632 427 2634 441
rect 2744 427 2746 441
rect 2872 427 2874 441
rect 3032 427 3034 441
rect 3224 427 3226 441
rect 3448 427 3450 441
rect 3680 427 3682 441
rect 3896 427 3898 441
rect 3992 427 3994 446
rect 110 426 116 427
rect 438 426 444 427
rect 112 403 114 426
rect 438 422 439 426
rect 443 422 444 426
rect 438 421 444 422
rect 542 426 548 427
rect 542 422 543 426
rect 547 422 548 426
rect 542 421 548 422
rect 646 426 652 427
rect 646 422 647 426
rect 651 422 652 426
rect 646 421 652 422
rect 750 426 756 427
rect 750 422 751 426
rect 755 422 756 426
rect 750 421 756 422
rect 854 426 860 427
rect 854 422 855 426
rect 859 422 860 426
rect 854 421 860 422
rect 958 426 964 427
rect 958 422 959 426
rect 963 422 964 426
rect 958 421 964 422
rect 1062 426 1068 427
rect 1062 422 1063 426
rect 1067 422 1068 426
rect 1062 421 1068 422
rect 1166 426 1172 427
rect 1166 422 1167 426
rect 1171 422 1172 426
rect 1166 421 1172 422
rect 1270 426 1276 427
rect 1270 422 1271 426
rect 1275 422 1276 426
rect 1270 421 1276 422
rect 1374 426 1380 427
rect 2030 426 2036 427
rect 2071 426 2075 427
rect 1374 422 1375 426
rect 1379 422 1380 426
rect 1374 421 1380 422
rect 440 403 442 421
rect 544 403 546 421
rect 648 403 650 421
rect 752 403 754 421
rect 856 403 858 421
rect 960 403 962 421
rect 1064 403 1066 421
rect 1168 403 1170 421
rect 1272 403 1274 421
rect 1376 403 1378 421
rect 2032 403 2034 426
rect 2071 421 2075 422
rect 2423 426 2427 427
rect 2423 421 2427 422
rect 2527 426 2531 427
rect 2527 421 2531 422
rect 2631 426 2635 427
rect 2631 421 2635 422
rect 2639 426 2643 427
rect 2639 421 2643 422
rect 2743 426 2747 427
rect 2743 421 2747 422
rect 2775 426 2779 427
rect 2775 421 2779 422
rect 2871 426 2875 427
rect 2871 421 2875 422
rect 2951 426 2955 427
rect 2951 421 2955 422
rect 3031 426 3035 427
rect 3031 421 3035 422
rect 3159 426 3163 427
rect 3159 421 3163 422
rect 3223 426 3227 427
rect 3223 421 3227 422
rect 3399 426 3403 427
rect 3399 421 3403 422
rect 3447 426 3451 427
rect 3447 421 3451 422
rect 3655 426 3659 427
rect 3655 421 3659 422
rect 3679 426 3683 427
rect 3679 421 3683 422
rect 3895 426 3899 427
rect 3895 421 3899 422
rect 3991 426 3995 427
rect 3991 421 3995 422
rect 2072 406 2074 421
rect 2528 411 2530 421
rect 2640 411 2642 421
rect 2776 411 2778 421
rect 2952 411 2954 421
rect 3160 411 3162 421
rect 3400 411 3402 421
rect 3656 411 3658 421
rect 3896 411 3898 421
rect 2526 410 2532 411
rect 2526 406 2527 410
rect 2531 406 2532 410
rect 2070 405 2076 406
rect 2526 405 2532 406
rect 2638 410 2644 411
rect 2638 406 2639 410
rect 2643 406 2644 410
rect 2638 405 2644 406
rect 2774 410 2780 411
rect 2774 406 2775 410
rect 2779 406 2780 410
rect 2774 405 2780 406
rect 2950 410 2956 411
rect 2950 406 2951 410
rect 2955 406 2956 410
rect 2950 405 2956 406
rect 3158 410 3164 411
rect 3158 406 3159 410
rect 3163 406 3164 410
rect 3158 405 3164 406
rect 3398 410 3404 411
rect 3398 406 3399 410
rect 3403 406 3404 410
rect 3398 405 3404 406
rect 3654 410 3660 411
rect 3654 406 3655 410
rect 3659 406 3660 410
rect 3654 405 3660 406
rect 3894 410 3900 411
rect 3894 406 3895 410
rect 3899 406 3900 410
rect 3992 406 3994 421
rect 3894 405 3900 406
rect 3990 405 3996 406
rect 111 402 115 403
rect 111 397 115 398
rect 439 402 443 403
rect 439 397 443 398
rect 543 402 547 403
rect 543 397 547 398
rect 623 402 627 403
rect 623 397 627 398
rect 647 402 651 403
rect 647 397 651 398
rect 727 402 731 403
rect 727 397 731 398
rect 751 402 755 403
rect 751 397 755 398
rect 831 402 835 403
rect 831 397 835 398
rect 855 402 859 403
rect 855 397 859 398
rect 935 402 939 403
rect 935 397 939 398
rect 959 402 963 403
rect 959 397 963 398
rect 1039 402 1043 403
rect 1039 397 1043 398
rect 1063 402 1067 403
rect 1063 397 1067 398
rect 1143 402 1147 403
rect 1143 397 1147 398
rect 1167 402 1171 403
rect 1167 397 1171 398
rect 1247 402 1251 403
rect 1247 397 1251 398
rect 1271 402 1275 403
rect 1271 397 1275 398
rect 1351 402 1355 403
rect 1351 397 1355 398
rect 1375 402 1379 403
rect 1375 397 1379 398
rect 1455 402 1459 403
rect 1455 397 1459 398
rect 1559 402 1563 403
rect 1559 397 1563 398
rect 2031 402 2035 403
rect 2070 401 2071 405
rect 2075 401 2076 405
rect 2070 400 2076 401
rect 3990 401 3991 405
rect 3995 401 3996 405
rect 3990 400 3996 401
rect 2031 397 2035 398
rect 112 382 114 397
rect 624 387 626 397
rect 728 387 730 397
rect 832 387 834 397
rect 936 387 938 397
rect 1040 387 1042 397
rect 1144 387 1146 397
rect 1248 387 1250 397
rect 1352 387 1354 397
rect 1456 387 1458 397
rect 1560 387 1562 397
rect 622 386 628 387
rect 622 382 623 386
rect 627 382 628 386
rect 110 381 116 382
rect 622 381 628 382
rect 726 386 732 387
rect 726 382 727 386
rect 731 382 732 386
rect 726 381 732 382
rect 830 386 836 387
rect 830 382 831 386
rect 835 382 836 386
rect 830 381 836 382
rect 934 386 940 387
rect 934 382 935 386
rect 939 382 940 386
rect 934 381 940 382
rect 1038 386 1044 387
rect 1038 382 1039 386
rect 1043 382 1044 386
rect 1038 381 1044 382
rect 1142 386 1148 387
rect 1142 382 1143 386
rect 1147 382 1148 386
rect 1142 381 1148 382
rect 1246 386 1252 387
rect 1246 382 1247 386
rect 1251 382 1252 386
rect 1246 381 1252 382
rect 1350 386 1356 387
rect 1350 382 1351 386
rect 1355 382 1356 386
rect 1350 381 1356 382
rect 1454 386 1460 387
rect 1454 382 1455 386
rect 1459 382 1460 386
rect 1454 381 1460 382
rect 1558 386 1564 387
rect 1558 382 1559 386
rect 1563 382 1564 386
rect 2032 382 2034 397
rect 2070 388 2076 389
rect 2070 384 2071 388
rect 2075 384 2076 388
rect 2070 383 2076 384
rect 3990 388 3996 389
rect 3990 384 3991 388
rect 3995 384 3996 388
rect 3990 383 3996 384
rect 1558 381 1564 382
rect 2030 381 2036 382
rect 110 377 111 381
rect 115 377 116 381
rect 110 376 116 377
rect 2030 377 2031 381
rect 2035 377 2036 381
rect 2030 376 2036 377
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 110 359 116 360
rect 2030 364 2036 365
rect 2030 360 2031 364
rect 2035 360 2036 364
rect 2030 359 2036 360
rect 112 331 114 359
rect 622 345 628 346
rect 622 341 623 345
rect 627 341 628 345
rect 622 340 628 341
rect 726 345 732 346
rect 726 341 727 345
rect 731 341 732 345
rect 726 340 732 341
rect 830 345 836 346
rect 830 341 831 345
rect 835 341 836 345
rect 830 340 836 341
rect 934 345 940 346
rect 934 341 935 345
rect 939 341 940 345
rect 934 340 940 341
rect 1038 345 1044 346
rect 1038 341 1039 345
rect 1043 341 1044 345
rect 1038 340 1044 341
rect 1142 345 1148 346
rect 1142 341 1143 345
rect 1147 341 1148 345
rect 1142 340 1148 341
rect 1246 345 1252 346
rect 1246 341 1247 345
rect 1251 341 1252 345
rect 1246 340 1252 341
rect 1350 345 1356 346
rect 1350 341 1351 345
rect 1355 341 1356 345
rect 1350 340 1356 341
rect 1454 345 1460 346
rect 1454 341 1455 345
rect 1459 341 1460 345
rect 1454 340 1460 341
rect 1558 345 1564 346
rect 1558 341 1559 345
rect 1563 341 1564 345
rect 1558 340 1564 341
rect 624 331 626 340
rect 728 331 730 340
rect 832 331 834 340
rect 936 331 938 340
rect 1040 331 1042 340
rect 1144 331 1146 340
rect 1248 331 1250 340
rect 1352 331 1354 340
rect 1456 331 1458 340
rect 1560 331 1562 340
rect 2032 331 2034 359
rect 2072 343 2074 383
rect 2526 369 2532 370
rect 2526 365 2527 369
rect 2531 365 2532 369
rect 2526 364 2532 365
rect 2638 369 2644 370
rect 2638 365 2639 369
rect 2643 365 2644 369
rect 2638 364 2644 365
rect 2774 369 2780 370
rect 2774 365 2775 369
rect 2779 365 2780 369
rect 2774 364 2780 365
rect 2950 369 2956 370
rect 2950 365 2951 369
rect 2955 365 2956 369
rect 2950 364 2956 365
rect 3158 369 3164 370
rect 3158 365 3159 369
rect 3163 365 3164 369
rect 3158 364 3164 365
rect 3398 369 3404 370
rect 3398 365 3399 369
rect 3403 365 3404 369
rect 3398 364 3404 365
rect 3654 369 3660 370
rect 3654 365 3655 369
rect 3659 365 3660 369
rect 3654 364 3660 365
rect 3894 369 3900 370
rect 3894 365 3895 369
rect 3899 365 3900 369
rect 3894 364 3900 365
rect 2528 343 2530 364
rect 2640 343 2642 364
rect 2776 343 2778 364
rect 2952 343 2954 364
rect 3160 343 3162 364
rect 3400 343 3402 364
rect 3656 343 3658 364
rect 3896 343 3898 364
rect 3992 343 3994 383
rect 2071 342 2075 343
rect 2071 337 2075 338
rect 2271 342 2275 343
rect 2271 337 2275 338
rect 2423 342 2427 343
rect 2423 337 2427 338
rect 2527 342 2531 343
rect 2527 337 2531 338
rect 2583 342 2587 343
rect 2583 337 2587 338
rect 2639 342 2643 343
rect 2639 337 2643 338
rect 2743 342 2747 343
rect 2743 337 2747 338
rect 2775 342 2779 343
rect 2775 337 2779 338
rect 2911 342 2915 343
rect 2911 337 2915 338
rect 2951 342 2955 343
rect 2951 337 2955 338
rect 3071 342 3075 343
rect 3071 337 3075 338
rect 3159 342 3163 343
rect 3159 337 3163 338
rect 3223 342 3227 343
rect 3223 337 3227 338
rect 3367 342 3371 343
rect 3367 337 3371 338
rect 3399 342 3403 343
rect 3399 337 3403 338
rect 3503 342 3507 343
rect 3503 337 3507 338
rect 3639 342 3643 343
rect 3639 337 3643 338
rect 3655 342 3659 343
rect 3655 337 3659 338
rect 3775 342 3779 343
rect 3775 337 3779 338
rect 3895 342 3899 343
rect 3895 337 3899 338
rect 3991 342 3995 343
rect 3991 337 3995 338
rect 111 330 115 331
rect 111 325 115 326
rect 399 330 403 331
rect 399 325 403 326
rect 543 330 547 331
rect 543 325 547 326
rect 623 330 627 331
rect 623 325 627 326
rect 687 330 691 331
rect 687 325 691 326
rect 727 330 731 331
rect 727 325 731 326
rect 831 330 835 331
rect 831 325 835 326
rect 839 330 843 331
rect 839 325 843 326
rect 935 330 939 331
rect 935 325 939 326
rect 991 330 995 331
rect 991 325 995 326
rect 1039 330 1043 331
rect 1039 325 1043 326
rect 1143 330 1147 331
rect 1143 325 1147 326
rect 1247 330 1251 331
rect 1247 325 1251 326
rect 1303 330 1307 331
rect 1303 325 1307 326
rect 1351 330 1355 331
rect 1351 325 1355 326
rect 1455 330 1459 331
rect 1455 325 1459 326
rect 1463 330 1467 331
rect 1463 325 1467 326
rect 1559 330 1563 331
rect 1559 325 1563 326
rect 1623 330 1627 331
rect 1623 325 1627 326
rect 2031 330 2035 331
rect 2031 325 2035 326
rect 112 297 114 325
rect 400 316 402 325
rect 544 316 546 325
rect 688 316 690 325
rect 840 316 842 325
rect 992 316 994 325
rect 1144 316 1146 325
rect 1304 316 1306 325
rect 1464 316 1466 325
rect 1624 316 1626 325
rect 398 315 404 316
rect 398 311 399 315
rect 403 311 404 315
rect 398 310 404 311
rect 542 315 548 316
rect 542 311 543 315
rect 547 311 548 315
rect 542 310 548 311
rect 686 315 692 316
rect 686 311 687 315
rect 691 311 692 315
rect 686 310 692 311
rect 838 315 844 316
rect 838 311 839 315
rect 843 311 844 315
rect 838 310 844 311
rect 990 315 996 316
rect 990 311 991 315
rect 995 311 996 315
rect 990 310 996 311
rect 1142 315 1148 316
rect 1142 311 1143 315
rect 1147 311 1148 315
rect 1142 310 1148 311
rect 1302 315 1308 316
rect 1302 311 1303 315
rect 1307 311 1308 315
rect 1302 310 1308 311
rect 1462 315 1468 316
rect 1462 311 1463 315
rect 1467 311 1468 315
rect 1462 310 1468 311
rect 1622 315 1628 316
rect 1622 311 1623 315
rect 1627 311 1628 315
rect 1622 310 1628 311
rect 2032 297 2034 325
rect 2072 309 2074 337
rect 2272 328 2274 337
rect 2424 328 2426 337
rect 2584 328 2586 337
rect 2744 328 2746 337
rect 2912 328 2914 337
rect 3072 328 3074 337
rect 3224 328 3226 337
rect 3368 328 3370 337
rect 3504 328 3506 337
rect 3640 328 3642 337
rect 3776 328 3778 337
rect 3896 328 3898 337
rect 2270 327 2276 328
rect 2270 323 2271 327
rect 2275 323 2276 327
rect 2270 322 2276 323
rect 2422 327 2428 328
rect 2422 323 2423 327
rect 2427 323 2428 327
rect 2422 322 2428 323
rect 2582 327 2588 328
rect 2582 323 2583 327
rect 2587 323 2588 327
rect 2582 322 2588 323
rect 2742 327 2748 328
rect 2742 323 2743 327
rect 2747 323 2748 327
rect 2742 322 2748 323
rect 2910 327 2916 328
rect 2910 323 2911 327
rect 2915 323 2916 327
rect 2910 322 2916 323
rect 3070 327 3076 328
rect 3070 323 3071 327
rect 3075 323 3076 327
rect 3070 322 3076 323
rect 3222 327 3228 328
rect 3222 323 3223 327
rect 3227 323 3228 327
rect 3222 322 3228 323
rect 3366 327 3372 328
rect 3366 323 3367 327
rect 3371 323 3372 327
rect 3366 322 3372 323
rect 3502 327 3508 328
rect 3502 323 3503 327
rect 3507 323 3508 327
rect 3502 322 3508 323
rect 3638 327 3644 328
rect 3638 323 3639 327
rect 3643 323 3644 327
rect 3638 322 3644 323
rect 3774 327 3780 328
rect 3774 323 3775 327
rect 3779 323 3780 327
rect 3774 322 3780 323
rect 3894 327 3900 328
rect 3894 323 3895 327
rect 3899 323 3900 327
rect 3894 322 3900 323
rect 3992 309 3994 337
rect 2070 308 2076 309
rect 2070 304 2071 308
rect 2075 304 2076 308
rect 2070 303 2076 304
rect 3990 308 3996 309
rect 3990 304 3991 308
rect 3995 304 3996 308
rect 3990 303 3996 304
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 2030 296 2036 297
rect 2030 292 2031 296
rect 2035 292 2036 296
rect 2030 291 2036 292
rect 2070 291 2076 292
rect 2070 287 2071 291
rect 2075 287 2076 291
rect 3990 291 3996 292
rect 3990 287 3991 291
rect 3995 287 3996 291
rect 2070 286 2076 287
rect 2270 286 2276 287
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 2030 279 2036 280
rect 2030 275 2031 279
rect 2035 275 2036 279
rect 110 274 116 275
rect 398 274 404 275
rect 112 255 114 274
rect 398 270 399 274
rect 403 270 404 274
rect 398 269 404 270
rect 542 274 548 275
rect 542 270 543 274
rect 547 270 548 274
rect 542 269 548 270
rect 686 274 692 275
rect 686 270 687 274
rect 691 270 692 274
rect 686 269 692 270
rect 838 274 844 275
rect 838 270 839 274
rect 843 270 844 274
rect 838 269 844 270
rect 990 274 996 275
rect 990 270 991 274
rect 995 270 996 274
rect 990 269 996 270
rect 1142 274 1148 275
rect 1142 270 1143 274
rect 1147 270 1148 274
rect 1142 269 1148 270
rect 1302 274 1308 275
rect 1302 270 1303 274
rect 1307 270 1308 274
rect 1302 269 1308 270
rect 1462 274 1468 275
rect 1462 270 1463 274
rect 1467 270 1468 274
rect 1462 269 1468 270
rect 1622 274 1628 275
rect 2030 274 2036 275
rect 1622 270 1623 274
rect 1627 270 1628 274
rect 1622 269 1628 270
rect 400 255 402 269
rect 544 255 546 269
rect 688 255 690 269
rect 840 255 842 269
rect 992 255 994 269
rect 1144 255 1146 269
rect 1304 255 1306 269
rect 1464 255 1466 269
rect 1624 255 1626 269
rect 2032 255 2034 274
rect 2072 263 2074 286
rect 2270 282 2271 286
rect 2275 282 2276 286
rect 2270 281 2276 282
rect 2422 286 2428 287
rect 2422 282 2423 286
rect 2427 282 2428 286
rect 2422 281 2428 282
rect 2582 286 2588 287
rect 2582 282 2583 286
rect 2587 282 2588 286
rect 2582 281 2588 282
rect 2742 286 2748 287
rect 2742 282 2743 286
rect 2747 282 2748 286
rect 2742 281 2748 282
rect 2910 286 2916 287
rect 2910 282 2911 286
rect 2915 282 2916 286
rect 2910 281 2916 282
rect 3070 286 3076 287
rect 3070 282 3071 286
rect 3075 282 3076 286
rect 3070 281 3076 282
rect 3222 286 3228 287
rect 3222 282 3223 286
rect 3227 282 3228 286
rect 3222 281 3228 282
rect 3366 286 3372 287
rect 3366 282 3367 286
rect 3371 282 3372 286
rect 3366 281 3372 282
rect 3502 286 3508 287
rect 3502 282 3503 286
rect 3507 282 3508 286
rect 3502 281 3508 282
rect 3638 286 3644 287
rect 3638 282 3639 286
rect 3643 282 3644 286
rect 3638 281 3644 282
rect 3774 286 3780 287
rect 3774 282 3775 286
rect 3779 282 3780 286
rect 3774 281 3780 282
rect 3894 286 3900 287
rect 3990 286 3996 287
rect 3894 282 3895 286
rect 3899 282 3900 286
rect 3894 281 3900 282
rect 2272 263 2274 281
rect 2424 263 2426 281
rect 2584 263 2586 281
rect 2744 263 2746 281
rect 2912 263 2914 281
rect 3072 263 3074 281
rect 3224 263 3226 281
rect 3368 263 3370 281
rect 3504 263 3506 281
rect 3640 263 3642 281
rect 3776 263 3778 281
rect 3896 263 3898 281
rect 3992 263 3994 286
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 2111 262 2115 263
rect 2111 257 2115 258
rect 2247 262 2251 263
rect 2247 257 2251 258
rect 2271 262 2275 263
rect 2271 257 2275 258
rect 2423 262 2427 263
rect 2423 257 2427 258
rect 2583 262 2587 263
rect 2583 257 2587 258
rect 2599 262 2603 263
rect 2599 257 2603 258
rect 2743 262 2747 263
rect 2743 257 2747 258
rect 2775 262 2779 263
rect 2775 257 2779 258
rect 2911 262 2915 263
rect 2911 257 2915 258
rect 2943 262 2947 263
rect 2943 257 2947 258
rect 3071 262 3075 263
rect 3071 257 3075 258
rect 3103 262 3107 263
rect 3103 257 3107 258
rect 3223 262 3227 263
rect 3223 257 3227 258
rect 3255 262 3259 263
rect 3255 257 3259 258
rect 3367 262 3371 263
rect 3367 257 3371 258
rect 3391 262 3395 263
rect 3391 257 3395 258
rect 3503 262 3507 263
rect 3503 257 3507 258
rect 3527 262 3531 263
rect 3527 257 3531 258
rect 3639 262 3643 263
rect 3639 257 3643 258
rect 3655 262 3659 263
rect 3655 257 3659 258
rect 3775 262 3779 263
rect 3775 257 3779 258
rect 3783 262 3787 263
rect 3783 257 3787 258
rect 3895 262 3899 263
rect 3895 257 3899 258
rect 3991 262 3995 263
rect 3991 257 3995 258
rect 111 254 115 255
rect 111 249 115 250
rect 207 254 211 255
rect 207 249 211 250
rect 399 254 403 255
rect 399 249 403 250
rect 431 254 435 255
rect 431 249 435 250
rect 543 254 547 255
rect 543 249 547 250
rect 655 254 659 255
rect 655 249 659 250
rect 687 254 691 255
rect 687 249 691 250
rect 839 254 843 255
rect 839 249 843 250
rect 871 254 875 255
rect 871 249 875 250
rect 991 254 995 255
rect 991 249 995 250
rect 1071 254 1075 255
rect 1071 249 1075 250
rect 1143 254 1147 255
rect 1143 249 1147 250
rect 1263 254 1267 255
rect 1263 249 1267 250
rect 1303 254 1307 255
rect 1303 249 1307 250
rect 1447 254 1451 255
rect 1447 249 1451 250
rect 1463 254 1467 255
rect 1463 249 1467 250
rect 1623 254 1627 255
rect 1623 249 1627 250
rect 1631 254 1635 255
rect 1631 249 1635 250
rect 1815 254 1819 255
rect 1815 249 1819 250
rect 2031 254 2035 255
rect 2031 249 2035 250
rect 112 234 114 249
rect 208 239 210 249
rect 432 239 434 249
rect 656 239 658 249
rect 872 239 874 249
rect 1072 239 1074 249
rect 1264 239 1266 249
rect 1448 239 1450 249
rect 1632 239 1634 249
rect 1816 239 1818 249
rect 206 238 212 239
rect 206 234 207 238
rect 211 234 212 238
rect 110 233 116 234
rect 206 233 212 234
rect 430 238 436 239
rect 430 234 431 238
rect 435 234 436 238
rect 430 233 436 234
rect 654 238 660 239
rect 654 234 655 238
rect 659 234 660 238
rect 654 233 660 234
rect 870 238 876 239
rect 870 234 871 238
rect 875 234 876 238
rect 870 233 876 234
rect 1070 238 1076 239
rect 1070 234 1071 238
rect 1075 234 1076 238
rect 1070 233 1076 234
rect 1262 238 1268 239
rect 1262 234 1263 238
rect 1267 234 1268 238
rect 1262 233 1268 234
rect 1446 238 1452 239
rect 1446 234 1447 238
rect 1451 234 1452 238
rect 1446 233 1452 234
rect 1630 238 1636 239
rect 1630 234 1631 238
rect 1635 234 1636 238
rect 1630 233 1636 234
rect 1814 238 1820 239
rect 1814 234 1815 238
rect 1819 234 1820 238
rect 2032 234 2034 249
rect 2072 242 2074 257
rect 2112 247 2114 257
rect 2248 247 2250 257
rect 2424 247 2426 257
rect 2600 247 2602 257
rect 2776 247 2778 257
rect 2944 247 2946 257
rect 3104 247 3106 257
rect 3256 247 3258 257
rect 3392 247 3394 257
rect 3528 247 3530 257
rect 3656 247 3658 257
rect 3784 247 3786 257
rect 3896 247 3898 257
rect 2110 246 2116 247
rect 2110 242 2111 246
rect 2115 242 2116 246
rect 2070 241 2076 242
rect 2110 241 2116 242
rect 2246 246 2252 247
rect 2246 242 2247 246
rect 2251 242 2252 246
rect 2246 241 2252 242
rect 2422 246 2428 247
rect 2422 242 2423 246
rect 2427 242 2428 246
rect 2422 241 2428 242
rect 2598 246 2604 247
rect 2598 242 2599 246
rect 2603 242 2604 246
rect 2598 241 2604 242
rect 2774 246 2780 247
rect 2774 242 2775 246
rect 2779 242 2780 246
rect 2774 241 2780 242
rect 2942 246 2948 247
rect 2942 242 2943 246
rect 2947 242 2948 246
rect 2942 241 2948 242
rect 3102 246 3108 247
rect 3102 242 3103 246
rect 3107 242 3108 246
rect 3102 241 3108 242
rect 3254 246 3260 247
rect 3254 242 3255 246
rect 3259 242 3260 246
rect 3254 241 3260 242
rect 3390 246 3396 247
rect 3390 242 3391 246
rect 3395 242 3396 246
rect 3390 241 3396 242
rect 3526 246 3532 247
rect 3526 242 3527 246
rect 3531 242 3532 246
rect 3526 241 3532 242
rect 3654 246 3660 247
rect 3654 242 3655 246
rect 3659 242 3660 246
rect 3654 241 3660 242
rect 3782 246 3788 247
rect 3782 242 3783 246
rect 3787 242 3788 246
rect 3782 241 3788 242
rect 3894 246 3900 247
rect 3894 242 3895 246
rect 3899 242 3900 246
rect 3992 242 3994 257
rect 3894 241 3900 242
rect 3990 241 3996 242
rect 2070 237 2071 241
rect 2075 237 2076 241
rect 2070 236 2076 237
rect 3990 237 3991 241
rect 3995 237 3996 241
rect 3990 236 3996 237
rect 1814 233 1820 234
rect 2030 233 2036 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 2030 229 2031 233
rect 2035 229 2036 233
rect 2030 228 2036 229
rect 2070 224 2076 225
rect 2070 220 2071 224
rect 2075 220 2076 224
rect 2070 219 2076 220
rect 3990 224 3996 225
rect 3990 220 3991 224
rect 3995 220 3996 224
rect 3990 219 3996 220
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 110 211 116 212
rect 2030 216 2036 217
rect 2030 212 2031 216
rect 2035 212 2036 216
rect 2030 211 2036 212
rect 112 155 114 211
rect 206 197 212 198
rect 206 193 207 197
rect 211 193 212 197
rect 206 192 212 193
rect 430 197 436 198
rect 430 193 431 197
rect 435 193 436 197
rect 430 192 436 193
rect 654 197 660 198
rect 654 193 655 197
rect 659 193 660 197
rect 654 192 660 193
rect 870 197 876 198
rect 870 193 871 197
rect 875 193 876 197
rect 870 192 876 193
rect 1070 197 1076 198
rect 1070 193 1071 197
rect 1075 193 1076 197
rect 1070 192 1076 193
rect 1262 197 1268 198
rect 1262 193 1263 197
rect 1267 193 1268 197
rect 1262 192 1268 193
rect 1446 197 1452 198
rect 1446 193 1447 197
rect 1451 193 1452 197
rect 1446 192 1452 193
rect 1630 197 1636 198
rect 1630 193 1631 197
rect 1635 193 1636 197
rect 1630 192 1636 193
rect 1814 197 1820 198
rect 1814 193 1815 197
rect 1819 193 1820 197
rect 1814 192 1820 193
rect 208 155 210 192
rect 432 155 434 192
rect 656 155 658 192
rect 872 155 874 192
rect 1072 155 1074 192
rect 1264 155 1266 192
rect 1448 155 1450 192
rect 1632 155 1634 192
rect 1816 155 1818 192
rect 2032 155 2034 211
rect 2072 179 2074 219
rect 2110 205 2116 206
rect 2110 201 2111 205
rect 2115 201 2116 205
rect 2110 200 2116 201
rect 2246 205 2252 206
rect 2246 201 2247 205
rect 2251 201 2252 205
rect 2246 200 2252 201
rect 2422 205 2428 206
rect 2422 201 2423 205
rect 2427 201 2428 205
rect 2422 200 2428 201
rect 2598 205 2604 206
rect 2598 201 2599 205
rect 2603 201 2604 205
rect 2598 200 2604 201
rect 2774 205 2780 206
rect 2774 201 2775 205
rect 2779 201 2780 205
rect 2774 200 2780 201
rect 2942 205 2948 206
rect 2942 201 2943 205
rect 2947 201 2948 205
rect 2942 200 2948 201
rect 3102 205 3108 206
rect 3102 201 3103 205
rect 3107 201 3108 205
rect 3102 200 3108 201
rect 3254 205 3260 206
rect 3254 201 3255 205
rect 3259 201 3260 205
rect 3254 200 3260 201
rect 3390 205 3396 206
rect 3390 201 3391 205
rect 3395 201 3396 205
rect 3390 200 3396 201
rect 3526 205 3532 206
rect 3526 201 3527 205
rect 3531 201 3532 205
rect 3526 200 3532 201
rect 3654 205 3660 206
rect 3654 201 3655 205
rect 3659 201 3660 205
rect 3654 200 3660 201
rect 3782 205 3788 206
rect 3782 201 3783 205
rect 3787 201 3788 205
rect 3782 200 3788 201
rect 3894 205 3900 206
rect 3894 201 3895 205
rect 3899 201 3900 205
rect 3894 200 3900 201
rect 2112 179 2114 200
rect 2248 179 2250 200
rect 2424 179 2426 200
rect 2600 179 2602 200
rect 2776 179 2778 200
rect 2944 179 2946 200
rect 3104 179 3106 200
rect 3256 179 3258 200
rect 3392 179 3394 200
rect 3528 179 3530 200
rect 3656 179 3658 200
rect 3784 179 3786 200
rect 3896 179 3898 200
rect 3992 179 3994 219
rect 2071 178 2075 179
rect 2071 173 2075 174
rect 2111 178 2115 179
rect 2111 173 2115 174
rect 2239 178 2243 179
rect 2239 173 2243 174
rect 2247 178 2251 179
rect 2247 173 2251 174
rect 2399 178 2403 179
rect 2399 173 2403 174
rect 2423 178 2427 179
rect 2423 173 2427 174
rect 2567 178 2571 179
rect 2567 173 2571 174
rect 2599 178 2603 179
rect 2599 173 2603 174
rect 2735 178 2739 179
rect 2735 173 2739 174
rect 2775 178 2779 179
rect 2775 173 2779 174
rect 2895 178 2899 179
rect 2895 173 2899 174
rect 2943 178 2947 179
rect 2943 173 2947 174
rect 3047 178 3051 179
rect 3047 173 3051 174
rect 3103 178 3107 179
rect 3103 173 3107 174
rect 3191 178 3195 179
rect 3191 173 3195 174
rect 3255 178 3259 179
rect 3255 173 3259 174
rect 3327 178 3331 179
rect 3327 173 3331 174
rect 3391 178 3395 179
rect 3391 173 3395 174
rect 3455 178 3459 179
rect 3455 173 3459 174
rect 3527 178 3531 179
rect 3527 173 3531 174
rect 3591 178 3595 179
rect 3591 173 3595 174
rect 3655 178 3659 179
rect 3655 173 3659 174
rect 3727 178 3731 179
rect 3727 173 3731 174
rect 3783 178 3787 179
rect 3783 173 3787 174
rect 3895 178 3899 179
rect 3895 173 3899 174
rect 3991 178 3995 179
rect 3991 173 3995 174
rect 111 154 115 155
rect 111 149 115 150
rect 151 154 155 155
rect 151 149 155 150
rect 207 154 211 155
rect 207 149 211 150
rect 255 154 259 155
rect 255 149 259 150
rect 359 154 363 155
rect 359 149 363 150
rect 431 154 435 155
rect 431 149 435 150
rect 463 154 467 155
rect 463 149 467 150
rect 567 154 571 155
rect 567 149 571 150
rect 655 154 659 155
rect 655 149 659 150
rect 671 154 675 155
rect 671 149 675 150
rect 775 154 779 155
rect 775 149 779 150
rect 871 154 875 155
rect 871 149 875 150
rect 879 154 883 155
rect 879 149 883 150
rect 983 154 987 155
rect 983 149 987 150
rect 1071 154 1075 155
rect 1071 149 1075 150
rect 1087 154 1091 155
rect 1087 149 1091 150
rect 1191 154 1195 155
rect 1191 149 1195 150
rect 1263 154 1267 155
rect 1263 149 1267 150
rect 1295 154 1299 155
rect 1295 149 1299 150
rect 1399 154 1403 155
rect 1399 149 1403 150
rect 1447 154 1451 155
rect 1447 149 1451 150
rect 1511 154 1515 155
rect 1511 149 1515 150
rect 1623 154 1627 155
rect 1623 149 1627 150
rect 1631 154 1635 155
rect 1631 149 1635 150
rect 1727 154 1731 155
rect 1727 149 1731 150
rect 1815 154 1819 155
rect 1815 149 1819 150
rect 1831 154 1835 155
rect 1831 149 1835 150
rect 1935 154 1939 155
rect 1935 149 1939 150
rect 2031 154 2035 155
rect 2031 149 2035 150
rect 112 121 114 149
rect 152 140 154 149
rect 256 140 258 149
rect 360 140 362 149
rect 464 140 466 149
rect 568 140 570 149
rect 672 140 674 149
rect 776 140 778 149
rect 880 140 882 149
rect 984 140 986 149
rect 1088 140 1090 149
rect 1192 140 1194 149
rect 1296 140 1298 149
rect 1400 140 1402 149
rect 1512 140 1514 149
rect 1624 140 1626 149
rect 1728 140 1730 149
rect 1832 140 1834 149
rect 1936 140 1938 149
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 150 134 156 135
rect 254 139 260 140
rect 254 135 255 139
rect 259 135 260 139
rect 254 134 260 135
rect 358 139 364 140
rect 358 135 359 139
rect 363 135 364 139
rect 358 134 364 135
rect 462 139 468 140
rect 462 135 463 139
rect 467 135 468 139
rect 462 134 468 135
rect 566 139 572 140
rect 566 135 567 139
rect 571 135 572 139
rect 566 134 572 135
rect 670 139 676 140
rect 670 135 671 139
rect 675 135 676 139
rect 670 134 676 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 878 139 884 140
rect 878 135 879 139
rect 883 135 884 139
rect 878 134 884 135
rect 982 139 988 140
rect 982 135 983 139
rect 987 135 988 139
rect 982 134 988 135
rect 1086 139 1092 140
rect 1086 135 1087 139
rect 1091 135 1092 139
rect 1086 134 1092 135
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1294 139 1300 140
rect 1294 135 1295 139
rect 1299 135 1300 139
rect 1294 134 1300 135
rect 1398 139 1404 140
rect 1398 135 1399 139
rect 1403 135 1404 139
rect 1398 134 1404 135
rect 1510 139 1516 140
rect 1510 135 1511 139
rect 1515 135 1516 139
rect 1510 134 1516 135
rect 1622 139 1628 140
rect 1622 135 1623 139
rect 1627 135 1628 139
rect 1622 134 1628 135
rect 1726 139 1732 140
rect 1726 135 1727 139
rect 1731 135 1732 139
rect 1726 134 1732 135
rect 1830 139 1836 140
rect 1830 135 1831 139
rect 1835 135 1836 139
rect 1830 134 1836 135
rect 1934 139 1940 140
rect 1934 135 1935 139
rect 1939 135 1940 139
rect 1934 134 1940 135
rect 2032 121 2034 149
rect 2072 145 2074 173
rect 2112 164 2114 173
rect 2240 164 2242 173
rect 2400 164 2402 173
rect 2568 164 2570 173
rect 2736 164 2738 173
rect 2896 164 2898 173
rect 3048 164 3050 173
rect 3192 164 3194 173
rect 3328 164 3330 173
rect 3456 164 3458 173
rect 3592 164 3594 173
rect 3728 164 3730 173
rect 2110 163 2116 164
rect 2110 159 2111 163
rect 2115 159 2116 163
rect 2110 158 2116 159
rect 2238 163 2244 164
rect 2238 159 2239 163
rect 2243 159 2244 163
rect 2238 158 2244 159
rect 2398 163 2404 164
rect 2398 159 2399 163
rect 2403 159 2404 163
rect 2398 158 2404 159
rect 2566 163 2572 164
rect 2566 159 2567 163
rect 2571 159 2572 163
rect 2566 158 2572 159
rect 2734 163 2740 164
rect 2734 159 2735 163
rect 2739 159 2740 163
rect 2734 158 2740 159
rect 2894 163 2900 164
rect 2894 159 2895 163
rect 2899 159 2900 163
rect 2894 158 2900 159
rect 3046 163 3052 164
rect 3046 159 3047 163
rect 3051 159 3052 163
rect 3046 158 3052 159
rect 3190 163 3196 164
rect 3190 159 3191 163
rect 3195 159 3196 163
rect 3190 158 3196 159
rect 3326 163 3332 164
rect 3326 159 3327 163
rect 3331 159 3332 163
rect 3326 158 3332 159
rect 3454 163 3460 164
rect 3454 159 3455 163
rect 3459 159 3460 163
rect 3454 158 3460 159
rect 3590 163 3596 164
rect 3590 159 3591 163
rect 3595 159 3596 163
rect 3590 158 3596 159
rect 3726 163 3732 164
rect 3726 159 3727 163
rect 3731 159 3732 163
rect 3726 158 3732 159
rect 3992 145 3994 173
rect 2070 144 2076 145
rect 2070 140 2071 144
rect 2075 140 2076 144
rect 2070 139 2076 140
rect 3990 144 3996 145
rect 3990 140 3991 144
rect 3995 140 3996 144
rect 3990 139 3996 140
rect 2070 127 2076 128
rect 2070 123 2071 127
rect 2075 123 2076 127
rect 3990 127 3996 128
rect 3990 123 3991 127
rect 3995 123 3996 127
rect 2070 122 2076 123
rect 2110 122 2116 123
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2030 115 2036 116
rect 2072 107 2074 122
rect 2110 118 2111 122
rect 2115 118 2116 122
rect 2110 117 2116 118
rect 2238 122 2244 123
rect 2238 118 2239 122
rect 2243 118 2244 122
rect 2238 117 2244 118
rect 2398 122 2404 123
rect 2398 118 2399 122
rect 2403 118 2404 122
rect 2398 117 2404 118
rect 2566 122 2572 123
rect 2566 118 2567 122
rect 2571 118 2572 122
rect 2566 117 2572 118
rect 2734 122 2740 123
rect 2734 118 2735 122
rect 2739 118 2740 122
rect 2734 117 2740 118
rect 2894 122 2900 123
rect 2894 118 2895 122
rect 2899 118 2900 122
rect 2894 117 2900 118
rect 3046 122 3052 123
rect 3046 118 3047 122
rect 3051 118 3052 122
rect 3046 117 3052 118
rect 3190 122 3196 123
rect 3190 118 3191 122
rect 3195 118 3196 122
rect 3190 117 3196 118
rect 3326 122 3332 123
rect 3326 118 3327 122
rect 3331 118 3332 122
rect 3326 117 3332 118
rect 3454 122 3460 123
rect 3454 118 3455 122
rect 3459 118 3460 122
rect 3454 117 3460 118
rect 3590 122 3596 123
rect 3590 118 3591 122
rect 3595 118 3596 122
rect 3590 117 3596 118
rect 3726 122 3732 123
rect 3990 122 3996 123
rect 3726 118 3727 122
rect 3731 118 3732 122
rect 3726 117 3732 118
rect 2112 107 2114 117
rect 2240 107 2242 117
rect 2400 107 2402 117
rect 2568 107 2570 117
rect 2736 107 2738 117
rect 2896 107 2898 117
rect 3048 107 3050 117
rect 3192 107 3194 117
rect 3328 107 3330 117
rect 3456 107 3458 117
rect 3592 107 3594 117
rect 3728 107 3730 117
rect 3992 107 3994 122
rect 2071 106 2075 107
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 2030 103 2036 104
rect 2030 99 2031 103
rect 2035 99 2036 103
rect 2071 101 2075 102
rect 2111 106 2115 107
rect 2111 101 2115 102
rect 2239 106 2243 107
rect 2239 101 2243 102
rect 2399 106 2403 107
rect 2399 101 2403 102
rect 2567 106 2571 107
rect 2567 101 2571 102
rect 2735 106 2739 107
rect 2735 101 2739 102
rect 2895 106 2899 107
rect 2895 101 2899 102
rect 3047 106 3051 107
rect 3047 101 3051 102
rect 3191 106 3195 107
rect 3191 101 3195 102
rect 3327 106 3331 107
rect 3327 101 3331 102
rect 3455 106 3459 107
rect 3455 101 3459 102
rect 3591 106 3595 107
rect 3591 101 3595 102
rect 3727 106 3731 107
rect 3727 101 3731 102
rect 3991 106 3995 107
rect 3991 101 3995 102
rect 110 98 116 99
rect 150 98 156 99
rect 112 83 114 98
rect 150 94 151 98
rect 155 94 156 98
rect 150 93 156 94
rect 254 98 260 99
rect 254 94 255 98
rect 259 94 260 98
rect 254 93 260 94
rect 358 98 364 99
rect 358 94 359 98
rect 363 94 364 98
rect 358 93 364 94
rect 462 98 468 99
rect 462 94 463 98
rect 467 94 468 98
rect 462 93 468 94
rect 566 98 572 99
rect 566 94 567 98
rect 571 94 572 98
rect 566 93 572 94
rect 670 98 676 99
rect 670 94 671 98
rect 675 94 676 98
rect 670 93 676 94
rect 774 98 780 99
rect 774 94 775 98
rect 779 94 780 98
rect 774 93 780 94
rect 878 98 884 99
rect 878 94 879 98
rect 883 94 884 98
rect 878 93 884 94
rect 982 98 988 99
rect 982 94 983 98
rect 987 94 988 98
rect 982 93 988 94
rect 1086 98 1092 99
rect 1086 94 1087 98
rect 1091 94 1092 98
rect 1086 93 1092 94
rect 1190 98 1196 99
rect 1190 94 1191 98
rect 1195 94 1196 98
rect 1190 93 1196 94
rect 1294 98 1300 99
rect 1294 94 1295 98
rect 1299 94 1300 98
rect 1294 93 1300 94
rect 1398 98 1404 99
rect 1398 94 1399 98
rect 1403 94 1404 98
rect 1398 93 1404 94
rect 1510 98 1516 99
rect 1510 94 1511 98
rect 1515 94 1516 98
rect 1510 93 1516 94
rect 1622 98 1628 99
rect 1622 94 1623 98
rect 1627 94 1628 98
rect 1622 93 1628 94
rect 1726 98 1732 99
rect 1726 94 1727 98
rect 1731 94 1732 98
rect 1726 93 1732 94
rect 1830 98 1836 99
rect 1830 94 1831 98
rect 1835 94 1836 98
rect 1830 93 1836 94
rect 1934 98 1940 99
rect 2030 98 2036 99
rect 1934 94 1935 98
rect 1939 94 1940 98
rect 1934 93 1940 94
rect 152 83 154 93
rect 256 83 258 93
rect 360 83 362 93
rect 464 83 466 93
rect 568 83 570 93
rect 672 83 674 93
rect 776 83 778 93
rect 880 83 882 93
rect 984 83 986 93
rect 1088 83 1090 93
rect 1192 83 1194 93
rect 1296 83 1298 93
rect 1400 83 1402 93
rect 1512 83 1514 93
rect 1624 83 1626 93
rect 1728 83 1730 93
rect 1832 83 1834 93
rect 1936 83 1938 93
rect 2032 83 2034 98
rect 111 82 115 83
rect 111 77 115 78
rect 151 82 155 83
rect 151 77 155 78
rect 255 82 259 83
rect 255 77 259 78
rect 359 82 363 83
rect 359 77 363 78
rect 463 82 467 83
rect 463 77 467 78
rect 567 82 571 83
rect 567 77 571 78
rect 671 82 675 83
rect 671 77 675 78
rect 775 82 779 83
rect 775 77 779 78
rect 879 82 883 83
rect 879 77 883 78
rect 983 82 987 83
rect 983 77 987 78
rect 1087 82 1091 83
rect 1087 77 1091 78
rect 1191 82 1195 83
rect 1191 77 1195 78
rect 1295 82 1299 83
rect 1295 77 1299 78
rect 1399 82 1403 83
rect 1399 77 1403 78
rect 1511 82 1515 83
rect 1511 77 1515 78
rect 1623 82 1627 83
rect 1623 77 1627 78
rect 1727 82 1731 83
rect 1727 77 1731 78
rect 1831 82 1835 83
rect 1831 77 1835 78
rect 1935 82 1939 83
rect 1935 77 1939 78
rect 2031 82 2035 83
rect 2031 77 2035 78
<< m4c >>
rect 2071 4078 2075 4082
rect 3399 4078 3403 4082
rect 3503 4078 3507 4082
rect 3607 4078 3611 4082
rect 3711 4078 3715 4082
rect 3991 4078 3995 4082
rect 111 4042 115 4046
rect 495 4042 499 4046
rect 599 4042 603 4046
rect 703 4042 707 4046
rect 807 4042 811 4046
rect 911 4042 915 4046
rect 1015 4042 1019 4046
rect 1119 4042 1123 4046
rect 1223 4042 1227 4046
rect 1327 4042 1331 4046
rect 1431 4042 1435 4046
rect 2031 4042 2035 4046
rect 2071 4006 2075 4010
rect 2111 4006 2115 4010
rect 2215 4006 2219 4010
rect 2319 4006 2323 4010
rect 2423 4006 2427 4010
rect 2527 4006 2531 4010
rect 2647 4006 2651 4010
rect 2775 4006 2779 4010
rect 2903 4006 2907 4010
rect 3031 4006 3035 4010
rect 3159 4006 3163 4010
rect 3287 4006 3291 4010
rect 3399 4006 3403 4010
rect 3415 4006 3419 4010
rect 3503 4006 3507 4010
rect 3551 4006 3555 4010
rect 3607 4006 3611 4010
rect 3711 4006 3715 4010
rect 3991 4006 3995 4010
rect 111 3970 115 3974
rect 391 3970 395 3974
rect 495 3970 499 3974
rect 599 3970 603 3974
rect 703 3970 707 3974
rect 807 3970 811 3974
rect 911 3970 915 3974
rect 1015 3970 1019 3974
rect 1119 3970 1123 3974
rect 1223 3970 1227 3974
rect 1327 3970 1331 3974
rect 1431 3970 1435 3974
rect 1535 3970 1539 3974
rect 2031 3970 2035 3974
rect 2071 3930 2075 3934
rect 2111 3930 2115 3934
rect 2143 3930 2147 3934
rect 2215 3930 2219 3934
rect 2319 3930 2323 3934
rect 2423 3930 2427 3934
rect 2487 3930 2491 3934
rect 2527 3930 2531 3934
rect 2647 3930 2651 3934
rect 2775 3930 2779 3934
rect 2799 3930 2803 3934
rect 2903 3930 2907 3934
rect 2951 3930 2955 3934
rect 3031 3930 3035 3934
rect 3103 3930 3107 3934
rect 3159 3930 3163 3934
rect 3255 3930 3259 3934
rect 3287 3930 3291 3934
rect 3415 3930 3419 3934
rect 3551 3930 3555 3934
rect 3991 3930 3995 3934
rect 111 3894 115 3898
rect 375 3894 379 3898
rect 391 3894 395 3898
rect 495 3894 499 3898
rect 599 3894 603 3898
rect 623 3894 627 3898
rect 703 3894 707 3898
rect 759 3894 763 3898
rect 807 3894 811 3898
rect 895 3894 899 3898
rect 911 3894 915 3898
rect 1015 3894 1019 3898
rect 1023 3894 1027 3898
rect 1119 3894 1123 3898
rect 1151 3894 1155 3898
rect 1223 3894 1227 3898
rect 1279 3894 1283 3898
rect 1327 3894 1331 3898
rect 1415 3894 1419 3898
rect 1431 3894 1435 3898
rect 1535 3894 1539 3898
rect 1551 3894 1555 3898
rect 2031 3894 2035 3898
rect 2071 3858 2075 3862
rect 2119 3858 2123 3862
rect 2143 3858 2147 3862
rect 2287 3858 2291 3862
rect 2319 3858 2323 3862
rect 2447 3858 2451 3862
rect 2487 3858 2491 3862
rect 2599 3858 2603 3862
rect 2647 3858 2651 3862
rect 2743 3858 2747 3862
rect 2799 3858 2803 3862
rect 2879 3858 2883 3862
rect 2951 3858 2955 3862
rect 3023 3858 3027 3862
rect 3103 3858 3107 3862
rect 3167 3858 3171 3862
rect 3255 3858 3259 3862
rect 3991 3858 3995 3862
rect 111 3814 115 3818
rect 375 3814 379 3818
rect 431 3814 435 3818
rect 495 3814 499 3818
rect 575 3814 579 3818
rect 623 3814 627 3818
rect 719 3814 723 3818
rect 759 3814 763 3818
rect 863 3814 867 3818
rect 895 3814 899 3818
rect 999 3814 1003 3818
rect 1023 3814 1027 3818
rect 1135 3814 1139 3818
rect 1151 3814 1155 3818
rect 1271 3814 1275 3818
rect 1279 3814 1283 3818
rect 1407 3814 1411 3818
rect 1415 3814 1419 3818
rect 1551 3814 1555 3818
rect 2031 3814 2035 3818
rect 2071 3782 2075 3786
rect 2111 3782 2115 3786
rect 2119 3782 2123 3786
rect 2239 3782 2243 3786
rect 2287 3782 2291 3786
rect 2391 3782 2395 3786
rect 2447 3782 2451 3786
rect 2543 3782 2547 3786
rect 2599 3782 2603 3786
rect 2687 3782 2691 3786
rect 2743 3782 2747 3786
rect 2823 3782 2827 3786
rect 2879 3782 2883 3786
rect 2951 3782 2955 3786
rect 3023 3782 3027 3786
rect 3087 3782 3091 3786
rect 3167 3782 3171 3786
rect 3223 3782 3227 3786
rect 3991 3782 3995 3786
rect 111 3734 115 3738
rect 359 3734 363 3738
rect 431 3734 435 3738
rect 495 3734 499 3738
rect 575 3734 579 3738
rect 631 3734 635 3738
rect 719 3734 723 3738
rect 775 3734 779 3738
rect 863 3734 867 3738
rect 919 3734 923 3738
rect 999 3734 1003 3738
rect 1071 3734 1075 3738
rect 1135 3734 1139 3738
rect 1223 3734 1227 3738
rect 1271 3734 1275 3738
rect 1375 3734 1379 3738
rect 1407 3734 1411 3738
rect 1527 3734 1531 3738
rect 1551 3734 1555 3738
rect 2031 3734 2035 3738
rect 2071 3702 2075 3706
rect 2111 3702 2115 3706
rect 2239 3702 2243 3706
rect 2295 3702 2299 3706
rect 2391 3702 2395 3706
rect 2487 3702 2491 3706
rect 2543 3702 2547 3706
rect 2671 3702 2675 3706
rect 2687 3702 2691 3706
rect 2823 3702 2827 3706
rect 2847 3702 2851 3706
rect 2951 3702 2955 3706
rect 3015 3702 3019 3706
rect 3087 3702 3091 3706
rect 3183 3702 3187 3706
rect 3223 3702 3227 3706
rect 3359 3702 3363 3706
rect 3991 3702 3995 3706
rect 111 3662 115 3666
rect 343 3662 347 3666
rect 359 3662 363 3666
rect 495 3662 499 3666
rect 519 3662 523 3666
rect 631 3662 635 3666
rect 695 3662 699 3666
rect 775 3662 779 3666
rect 863 3662 867 3666
rect 919 3662 923 3666
rect 1031 3662 1035 3666
rect 1071 3662 1075 3666
rect 1191 3662 1195 3666
rect 1223 3662 1227 3666
rect 1343 3662 1347 3666
rect 1375 3662 1379 3666
rect 1495 3662 1499 3666
rect 1527 3662 1531 3666
rect 1655 3662 1659 3666
rect 2031 3662 2035 3666
rect 2071 3622 2075 3626
rect 2111 3622 2115 3626
rect 2295 3622 2299 3626
rect 2487 3622 2491 3626
rect 2495 3622 2499 3626
rect 2671 3622 2675 3626
rect 2687 3622 2691 3626
rect 2847 3622 2851 3626
rect 2863 3622 2867 3626
rect 3015 3622 3019 3626
rect 3023 3622 3027 3626
rect 3167 3622 3171 3626
rect 3183 3622 3187 3626
rect 3303 3622 3307 3626
rect 3359 3622 3363 3626
rect 3431 3622 3435 3626
rect 3551 3622 3555 3626
rect 3671 3622 3675 3626
rect 3791 3622 3795 3626
rect 3895 3622 3899 3626
rect 3991 3622 3995 3626
rect 111 3590 115 3594
rect 239 3590 243 3594
rect 343 3590 347 3594
rect 399 3590 403 3594
rect 519 3590 523 3594
rect 551 3590 555 3594
rect 695 3590 699 3594
rect 703 3590 707 3594
rect 855 3590 859 3594
rect 863 3590 867 3594
rect 999 3590 1003 3594
rect 1031 3590 1035 3594
rect 1135 3590 1139 3594
rect 1191 3590 1195 3594
rect 1263 3590 1267 3594
rect 1343 3590 1347 3594
rect 1383 3590 1387 3594
rect 1495 3590 1499 3594
rect 1607 3590 1611 3594
rect 1655 3590 1659 3594
rect 1719 3590 1723 3594
rect 1831 3590 1835 3594
rect 1935 3590 1939 3594
rect 2031 3590 2035 3594
rect 2071 3538 2075 3542
rect 2111 3538 2115 3542
rect 2295 3538 2299 3542
rect 2447 3538 2451 3542
rect 2495 3538 2499 3542
rect 2591 3538 2595 3542
rect 2687 3538 2691 3542
rect 2727 3538 2731 3542
rect 2863 3538 2867 3542
rect 2991 3538 2995 3542
rect 3023 3538 3027 3542
rect 3119 3538 3123 3542
rect 3167 3538 3171 3542
rect 3239 3538 3243 3542
rect 3303 3538 3307 3542
rect 3351 3538 3355 3542
rect 3431 3538 3435 3542
rect 3463 3538 3467 3542
rect 3551 3538 3555 3542
rect 3575 3538 3579 3542
rect 3671 3538 3675 3542
rect 3687 3538 3691 3542
rect 3791 3538 3795 3542
rect 3895 3538 3899 3542
rect 3991 3538 3995 3542
rect 111 3518 115 3522
rect 151 3518 155 3522
rect 239 3518 243 3522
rect 375 3518 379 3522
rect 399 3518 403 3522
rect 551 3518 555 3522
rect 615 3518 619 3522
rect 703 3518 707 3522
rect 847 3518 851 3522
rect 855 3518 859 3522
rect 999 3518 1003 3522
rect 1063 3518 1067 3522
rect 1135 3518 1139 3522
rect 1255 3518 1259 3522
rect 1263 3518 1267 3522
rect 1383 3518 1387 3522
rect 1439 3518 1443 3522
rect 1495 3518 1499 3522
rect 1607 3518 1611 3522
rect 1615 3518 1619 3522
rect 1719 3518 1723 3522
rect 1783 3518 1787 3522
rect 1831 3518 1835 3522
rect 1935 3518 1939 3522
rect 2031 3518 2035 3522
rect 2071 3466 2075 3470
rect 2343 3466 2347 3470
rect 2447 3466 2451 3470
rect 2591 3466 2595 3470
rect 2727 3466 2731 3470
rect 2855 3466 2859 3470
rect 2863 3466 2867 3470
rect 2991 3466 2995 3470
rect 3119 3466 3123 3470
rect 3239 3466 3243 3470
rect 3351 3466 3355 3470
rect 3375 3466 3379 3470
rect 3463 3466 3467 3470
rect 3575 3466 3579 3470
rect 3687 3466 3691 3470
rect 3791 3466 3795 3470
rect 3895 3466 3899 3470
rect 3991 3466 3995 3470
rect 111 3422 115 3426
rect 151 3422 155 3426
rect 335 3422 339 3426
rect 375 3422 379 3426
rect 583 3422 587 3426
rect 615 3422 619 3426
rect 847 3422 851 3426
rect 863 3422 867 3426
rect 1063 3422 1067 3426
rect 1159 3422 1163 3426
rect 1255 3422 1259 3426
rect 1439 3422 1443 3426
rect 1463 3422 1467 3426
rect 1615 3422 1619 3426
rect 1783 3422 1787 3426
rect 1935 3422 1939 3426
rect 2031 3422 2035 3426
rect 2071 3390 2075 3394
rect 2183 3390 2187 3394
rect 2343 3390 2347 3394
rect 2583 3390 2587 3394
rect 2855 3390 2859 3394
rect 3007 3390 3011 3394
rect 3375 3390 3379 3394
rect 3447 3390 3451 3394
rect 3895 3390 3899 3394
rect 3991 3390 3995 3394
rect 111 3342 115 3346
rect 151 3342 155 3346
rect 287 3342 291 3346
rect 335 3342 339 3346
rect 463 3342 467 3346
rect 583 3342 587 3346
rect 639 3342 643 3346
rect 815 3342 819 3346
rect 863 3342 867 3346
rect 991 3342 995 3346
rect 1159 3342 1163 3346
rect 1319 3342 1323 3346
rect 1463 3342 1467 3346
rect 1487 3342 1491 3346
rect 1655 3342 1659 3346
rect 2031 3342 2035 3346
rect 2071 3302 2075 3306
rect 2111 3302 2115 3306
rect 2183 3302 2187 3306
rect 2295 3302 2299 3306
rect 2503 3302 2507 3306
rect 2583 3302 2587 3306
rect 2703 3302 2707 3306
rect 2895 3302 2899 3306
rect 3007 3302 3011 3306
rect 3071 3302 3075 3306
rect 3231 3302 3235 3306
rect 3375 3302 3379 3306
rect 3447 3302 3451 3306
rect 3511 3302 3515 3306
rect 3647 3302 3651 3306
rect 3783 3302 3787 3306
rect 3895 3302 3899 3306
rect 3991 3302 3995 3306
rect 111 3258 115 3262
rect 151 3258 155 3262
rect 287 3258 291 3262
rect 295 3258 299 3262
rect 463 3258 467 3262
rect 479 3258 483 3262
rect 639 3258 643 3262
rect 671 3258 675 3262
rect 815 3258 819 3262
rect 863 3258 867 3262
rect 991 3258 995 3262
rect 1055 3258 1059 3262
rect 1159 3258 1163 3262
rect 1247 3258 1251 3262
rect 1319 3258 1323 3262
rect 1431 3258 1435 3262
rect 1487 3258 1491 3262
rect 1615 3258 1619 3262
rect 1655 3258 1659 3262
rect 1807 3258 1811 3262
rect 2031 3258 2035 3262
rect 2071 3230 2075 3234
rect 2111 3230 2115 3234
rect 2239 3230 2243 3234
rect 2295 3230 2299 3234
rect 2399 3230 2403 3234
rect 2503 3230 2507 3234
rect 2559 3230 2563 3234
rect 2703 3230 2707 3234
rect 2719 3230 2723 3234
rect 2879 3230 2883 3234
rect 2895 3230 2899 3234
rect 3031 3230 3035 3234
rect 3071 3230 3075 3234
rect 3167 3230 3171 3234
rect 3231 3230 3235 3234
rect 3303 3230 3307 3234
rect 3375 3230 3379 3234
rect 3431 3230 3435 3234
rect 3511 3230 3515 3234
rect 3551 3230 3555 3234
rect 3647 3230 3651 3234
rect 3671 3230 3675 3234
rect 3783 3230 3787 3234
rect 3791 3230 3795 3234
rect 3895 3230 3899 3234
rect 3991 3230 3995 3234
rect 111 3174 115 3178
rect 151 3174 155 3178
rect 287 3174 291 3178
rect 295 3174 299 3178
rect 423 3174 427 3178
rect 479 3174 483 3178
rect 567 3174 571 3178
rect 671 3174 675 3178
rect 727 3174 731 3178
rect 863 3174 867 3178
rect 903 3174 907 3178
rect 1055 3174 1059 3178
rect 1095 3174 1099 3178
rect 1247 3174 1251 3178
rect 1295 3174 1299 3178
rect 1431 3174 1435 3178
rect 1495 3174 1499 3178
rect 1615 3174 1619 3178
rect 1703 3174 1707 3178
rect 1807 3174 1811 3178
rect 1919 3174 1923 3178
rect 2031 3174 2035 3178
rect 2071 3142 2075 3146
rect 2111 3142 2115 3146
rect 2183 3142 2187 3146
rect 2239 3142 2243 3146
rect 2367 3142 2371 3146
rect 2399 3142 2403 3146
rect 2551 3142 2555 3146
rect 2559 3142 2563 3146
rect 2719 3142 2723 3146
rect 2735 3142 2739 3146
rect 2879 3142 2883 3146
rect 2911 3142 2915 3146
rect 3031 3142 3035 3146
rect 3087 3142 3091 3146
rect 3167 3142 3171 3146
rect 3263 3142 3267 3146
rect 3303 3142 3307 3146
rect 3431 3142 3435 3146
rect 3447 3142 3451 3146
rect 3551 3142 3555 3146
rect 3671 3142 3675 3146
rect 3791 3142 3795 3146
rect 3895 3142 3899 3146
rect 3991 3142 3995 3146
rect 111 3086 115 3090
rect 287 3086 291 3090
rect 423 3086 427 3090
rect 567 3086 571 3090
rect 575 3086 579 3090
rect 679 3086 683 3090
rect 727 3086 731 3090
rect 799 3086 803 3090
rect 903 3086 907 3090
rect 935 3086 939 3090
rect 1079 3086 1083 3090
rect 1095 3086 1099 3090
rect 1231 3086 1235 3090
rect 1295 3086 1299 3090
rect 1391 3086 1395 3090
rect 1495 3086 1499 3090
rect 1559 3086 1563 3090
rect 1703 3086 1707 3090
rect 1727 3086 1731 3090
rect 1903 3086 1907 3090
rect 1919 3086 1923 3090
rect 2031 3086 2035 3090
rect 2071 3062 2075 3066
rect 2183 3062 2187 3066
rect 2351 3062 2355 3066
rect 2367 3062 2371 3066
rect 2455 3062 2459 3066
rect 2551 3062 2555 3066
rect 2567 3062 2571 3066
rect 2687 3062 2691 3066
rect 2735 3062 2739 3066
rect 2807 3062 2811 3066
rect 2911 3062 2915 3066
rect 2927 3062 2931 3066
rect 3047 3062 3051 3066
rect 3087 3062 3091 3066
rect 3167 3062 3171 3066
rect 3263 3062 3267 3066
rect 3295 3062 3299 3066
rect 3447 3062 3451 3066
rect 3991 3062 3995 3066
rect 111 3002 115 3006
rect 551 3002 555 3006
rect 575 3002 579 3006
rect 655 3002 659 3006
rect 679 3002 683 3006
rect 759 3002 763 3006
rect 799 3002 803 3006
rect 871 3002 875 3006
rect 935 3002 939 3006
rect 991 3002 995 3006
rect 1079 3002 1083 3006
rect 1119 3002 1123 3006
rect 1231 3002 1235 3006
rect 1255 3002 1259 3006
rect 1391 3002 1395 3006
rect 1535 3002 1539 3006
rect 1559 3002 1563 3006
rect 1687 3002 1691 3006
rect 1727 3002 1731 3006
rect 1903 3002 1907 3006
rect 2031 3002 2035 3006
rect 2071 2990 2075 2994
rect 2351 2990 2355 2994
rect 2455 2990 2459 2994
rect 2495 2990 2499 2994
rect 2567 2990 2571 2994
rect 2599 2990 2603 2994
rect 2687 2990 2691 2994
rect 2703 2990 2707 2994
rect 2807 2990 2811 2994
rect 2911 2990 2915 2994
rect 2927 2990 2931 2994
rect 3015 2990 3019 2994
rect 3047 2990 3051 2994
rect 3119 2990 3123 2994
rect 3167 2990 3171 2994
rect 3223 2990 3227 2994
rect 3295 2990 3299 2994
rect 3991 2990 3995 2994
rect 111 2918 115 2922
rect 311 2918 315 2922
rect 431 2918 435 2922
rect 551 2918 555 2922
rect 559 2918 563 2922
rect 655 2918 659 2922
rect 695 2918 699 2922
rect 759 2918 763 2922
rect 831 2918 835 2922
rect 871 2918 875 2922
rect 975 2918 979 2922
rect 991 2918 995 2922
rect 1119 2918 1123 2922
rect 1255 2918 1259 2922
rect 1271 2918 1275 2922
rect 1391 2918 1395 2922
rect 1423 2918 1427 2922
rect 1535 2918 1539 2922
rect 1575 2918 1579 2922
rect 1687 2918 1691 2922
rect 2031 2918 2035 2922
rect 2071 2918 2075 2922
rect 2415 2918 2419 2922
rect 2495 2918 2499 2922
rect 2519 2918 2523 2922
rect 2599 2918 2603 2922
rect 2623 2918 2627 2922
rect 2703 2918 2707 2922
rect 2727 2918 2731 2922
rect 2807 2918 2811 2922
rect 2831 2918 2835 2922
rect 2911 2918 2915 2922
rect 2935 2918 2939 2922
rect 3015 2918 3019 2922
rect 3039 2918 3043 2922
rect 3119 2918 3123 2922
rect 3143 2918 3147 2922
rect 3223 2918 3227 2922
rect 3247 2918 3251 2922
rect 3991 2918 3995 2922
rect 2071 2842 2075 2846
rect 2407 2842 2411 2846
rect 2415 2842 2419 2846
rect 2511 2842 2515 2846
rect 2519 2842 2523 2846
rect 2615 2842 2619 2846
rect 2623 2842 2627 2846
rect 2719 2842 2723 2846
rect 2727 2842 2731 2846
rect 2823 2842 2827 2846
rect 2831 2842 2835 2846
rect 2927 2842 2931 2846
rect 2935 2842 2939 2846
rect 3031 2842 3035 2846
rect 3039 2842 3043 2846
rect 3135 2842 3139 2846
rect 3143 2842 3147 2846
rect 3239 2842 3243 2846
rect 3247 2842 3251 2846
rect 3991 2842 3995 2846
rect 111 2830 115 2834
rect 151 2830 155 2834
rect 311 2830 315 2834
rect 431 2830 435 2834
rect 471 2830 475 2834
rect 559 2830 563 2834
rect 623 2830 627 2834
rect 695 2830 699 2834
rect 767 2830 771 2834
rect 831 2830 835 2834
rect 903 2830 907 2834
rect 975 2830 979 2834
rect 1031 2830 1035 2834
rect 1119 2830 1123 2834
rect 1159 2830 1163 2834
rect 1271 2830 1275 2834
rect 1287 2830 1291 2834
rect 1415 2830 1419 2834
rect 1423 2830 1427 2834
rect 1575 2830 1579 2834
rect 2031 2830 2035 2834
rect 2071 2762 2075 2766
rect 2303 2762 2307 2766
rect 2407 2762 2411 2766
rect 2415 2762 2419 2766
rect 2511 2762 2515 2766
rect 2535 2762 2539 2766
rect 2615 2762 2619 2766
rect 2655 2762 2659 2766
rect 2719 2762 2723 2766
rect 2775 2762 2779 2766
rect 2823 2762 2827 2766
rect 2895 2762 2899 2766
rect 2927 2762 2931 2766
rect 3015 2762 3019 2766
rect 3031 2762 3035 2766
rect 3135 2762 3139 2766
rect 3143 2762 3147 2766
rect 3239 2762 3243 2766
rect 3271 2762 3275 2766
rect 3399 2762 3403 2766
rect 3991 2762 3995 2766
rect 111 2742 115 2746
rect 151 2742 155 2746
rect 303 2742 307 2746
rect 311 2742 315 2746
rect 471 2742 475 2746
rect 623 2742 627 2746
rect 767 2742 771 2746
rect 903 2742 907 2746
rect 1031 2742 1035 2746
rect 1039 2742 1043 2746
rect 1159 2742 1163 2746
rect 1167 2742 1171 2746
rect 1287 2742 1291 2746
rect 1295 2742 1299 2746
rect 1415 2742 1419 2746
rect 1423 2742 1427 2746
rect 2031 2742 2035 2746
rect 2071 2674 2075 2678
rect 2151 2674 2155 2678
rect 2303 2674 2307 2678
rect 2415 2674 2419 2678
rect 2463 2674 2467 2678
rect 2535 2674 2539 2678
rect 2623 2674 2627 2678
rect 2655 2674 2659 2678
rect 2775 2674 2779 2678
rect 2791 2674 2795 2678
rect 2895 2674 2899 2678
rect 2951 2674 2955 2678
rect 3015 2674 3019 2678
rect 3111 2674 3115 2678
rect 3143 2674 3147 2678
rect 3263 2674 3267 2678
rect 3271 2674 3275 2678
rect 3399 2674 3403 2678
rect 3415 2674 3419 2678
rect 3575 2674 3579 2678
rect 3991 2674 3995 2678
rect 111 2658 115 2662
rect 151 2658 155 2662
rect 303 2658 307 2662
rect 319 2658 323 2662
rect 471 2658 475 2662
rect 511 2658 515 2662
rect 623 2658 627 2662
rect 703 2658 707 2662
rect 767 2658 771 2662
rect 887 2658 891 2662
rect 903 2658 907 2662
rect 1039 2658 1043 2662
rect 1063 2658 1067 2662
rect 1167 2658 1171 2662
rect 1231 2658 1235 2662
rect 1295 2658 1299 2662
rect 1391 2658 1395 2662
rect 1423 2658 1427 2662
rect 1551 2658 1555 2662
rect 1711 2658 1715 2662
rect 2031 2658 2035 2662
rect 2071 2594 2075 2598
rect 2111 2594 2115 2598
rect 2151 2594 2155 2598
rect 2303 2594 2307 2598
rect 2327 2594 2331 2598
rect 2463 2594 2467 2598
rect 2559 2594 2563 2598
rect 2623 2594 2627 2598
rect 2783 2594 2787 2598
rect 2791 2594 2795 2598
rect 2951 2594 2955 2598
rect 2999 2594 3003 2598
rect 3111 2594 3115 2598
rect 3199 2594 3203 2598
rect 3263 2594 3267 2598
rect 3383 2594 3387 2598
rect 3415 2594 3419 2598
rect 3559 2594 3563 2598
rect 3575 2594 3579 2598
rect 3735 2594 3739 2598
rect 3895 2594 3899 2598
rect 3991 2594 3995 2598
rect 111 2570 115 2574
rect 151 2570 155 2574
rect 279 2570 283 2574
rect 319 2570 323 2574
rect 463 2570 467 2574
rect 511 2570 515 2574
rect 663 2570 667 2574
rect 703 2570 707 2574
rect 863 2570 867 2574
rect 887 2570 891 2574
rect 1063 2570 1067 2574
rect 1231 2570 1235 2574
rect 1255 2570 1259 2574
rect 1391 2570 1395 2574
rect 1431 2570 1435 2574
rect 1551 2570 1555 2574
rect 1607 2570 1611 2574
rect 1711 2570 1715 2574
rect 1783 2570 1787 2574
rect 1935 2570 1939 2574
rect 2031 2570 2035 2574
rect 2071 2522 2075 2526
rect 2111 2522 2115 2526
rect 2255 2522 2259 2526
rect 2327 2522 2331 2526
rect 2439 2522 2443 2526
rect 2559 2522 2563 2526
rect 2631 2522 2635 2526
rect 2783 2522 2787 2526
rect 2823 2522 2827 2526
rect 2999 2522 3003 2526
rect 3007 2522 3011 2526
rect 3175 2522 3179 2526
rect 3199 2522 3203 2526
rect 3335 2522 3339 2526
rect 3383 2522 3387 2526
rect 3487 2522 3491 2526
rect 3559 2522 3563 2526
rect 3631 2522 3635 2526
rect 3735 2522 3739 2526
rect 3775 2522 3779 2526
rect 3895 2522 3899 2526
rect 3991 2522 3995 2526
rect 111 2482 115 2486
rect 279 2482 283 2486
rect 311 2482 315 2486
rect 463 2482 467 2486
rect 471 2482 475 2486
rect 647 2482 651 2486
rect 663 2482 667 2486
rect 831 2482 835 2486
rect 863 2482 867 2486
rect 1015 2482 1019 2486
rect 1063 2482 1067 2486
rect 1191 2482 1195 2486
rect 1255 2482 1259 2486
rect 1367 2482 1371 2486
rect 1431 2482 1435 2486
rect 1535 2482 1539 2486
rect 1607 2482 1611 2486
rect 1703 2482 1707 2486
rect 1783 2482 1787 2486
rect 1871 2482 1875 2486
rect 1935 2482 1939 2486
rect 2031 2482 2035 2486
rect 2071 2442 2075 2446
rect 2111 2442 2115 2446
rect 2255 2442 2259 2446
rect 2311 2442 2315 2446
rect 2439 2442 2443 2446
rect 2535 2442 2539 2446
rect 2631 2442 2635 2446
rect 2751 2442 2755 2446
rect 2823 2442 2827 2446
rect 2951 2442 2955 2446
rect 3007 2442 3011 2446
rect 3135 2442 3139 2446
rect 3175 2442 3179 2446
rect 3311 2442 3315 2446
rect 3335 2442 3339 2446
rect 3471 2442 3475 2446
rect 3487 2442 3491 2446
rect 3623 2442 3627 2446
rect 3631 2442 3635 2446
rect 3767 2442 3771 2446
rect 3775 2442 3779 2446
rect 3895 2442 3899 2446
rect 3991 2442 3995 2446
rect 111 2398 115 2402
rect 207 2398 211 2402
rect 311 2398 315 2402
rect 351 2398 355 2402
rect 471 2398 475 2402
rect 503 2398 507 2402
rect 647 2398 651 2402
rect 655 2398 659 2402
rect 815 2398 819 2402
rect 831 2398 835 2402
rect 967 2398 971 2402
rect 1015 2398 1019 2402
rect 1119 2398 1123 2402
rect 1191 2398 1195 2402
rect 1263 2398 1267 2402
rect 1367 2398 1371 2402
rect 1415 2398 1419 2402
rect 1535 2398 1539 2402
rect 1567 2398 1571 2402
rect 1703 2398 1707 2402
rect 1871 2398 1875 2402
rect 2031 2398 2035 2402
rect 2071 2370 2075 2374
rect 2111 2370 2115 2374
rect 2311 2370 2315 2374
rect 2327 2370 2331 2374
rect 2535 2370 2539 2374
rect 2559 2370 2563 2374
rect 2751 2370 2755 2374
rect 2783 2370 2787 2374
rect 2951 2370 2955 2374
rect 2999 2370 3003 2374
rect 3135 2370 3139 2374
rect 3191 2370 3195 2374
rect 3311 2370 3315 2374
rect 3375 2370 3379 2374
rect 3471 2370 3475 2374
rect 3543 2370 3547 2374
rect 3623 2370 3627 2374
rect 3711 2370 3715 2374
rect 3767 2370 3771 2374
rect 3887 2370 3891 2374
rect 3895 2370 3899 2374
rect 3991 2370 3995 2374
rect 111 2314 115 2318
rect 207 2314 211 2318
rect 255 2314 259 2318
rect 351 2314 355 2318
rect 359 2314 363 2318
rect 471 2314 475 2318
rect 503 2314 507 2318
rect 583 2314 587 2318
rect 655 2314 659 2318
rect 695 2314 699 2318
rect 807 2314 811 2318
rect 815 2314 819 2318
rect 919 2314 923 2318
rect 967 2314 971 2318
rect 1031 2314 1035 2318
rect 1119 2314 1123 2318
rect 1151 2314 1155 2318
rect 1263 2314 1267 2318
rect 1271 2314 1275 2318
rect 1415 2314 1419 2318
rect 1567 2314 1571 2318
rect 2031 2314 2035 2318
rect 2071 2298 2075 2302
rect 2111 2298 2115 2302
rect 2295 2298 2299 2302
rect 2327 2298 2331 2302
rect 2527 2298 2531 2302
rect 2559 2298 2563 2302
rect 2775 2298 2779 2302
rect 2783 2298 2787 2302
rect 2999 2298 3003 2302
rect 3039 2298 3043 2302
rect 3191 2298 3195 2302
rect 3319 2298 3323 2302
rect 3375 2298 3379 2302
rect 3543 2298 3547 2302
rect 3607 2298 3611 2302
rect 3711 2298 3715 2302
rect 3887 2298 3891 2302
rect 3895 2298 3899 2302
rect 3991 2298 3995 2302
rect 111 2230 115 2234
rect 183 2230 187 2234
rect 255 2230 259 2234
rect 343 2230 347 2234
rect 359 2230 363 2234
rect 471 2230 475 2234
rect 495 2230 499 2234
rect 583 2230 587 2234
rect 647 2230 651 2234
rect 695 2230 699 2234
rect 791 2230 795 2234
rect 807 2230 811 2234
rect 919 2230 923 2234
rect 935 2230 939 2234
rect 1031 2230 1035 2234
rect 1071 2230 1075 2234
rect 1151 2230 1155 2234
rect 1199 2230 1203 2234
rect 1271 2230 1275 2234
rect 1335 2230 1339 2234
rect 1471 2230 1475 2234
rect 2031 2230 2035 2234
rect 2071 2218 2075 2222
rect 2111 2218 2115 2222
rect 2279 2218 2283 2222
rect 2295 2218 2299 2222
rect 2439 2218 2443 2222
rect 2527 2218 2531 2222
rect 2623 2218 2627 2222
rect 2775 2218 2779 2222
rect 2839 2218 2843 2222
rect 3039 2218 3043 2222
rect 3079 2218 3083 2222
rect 3319 2218 3323 2222
rect 3343 2218 3347 2222
rect 3607 2218 3611 2222
rect 3623 2218 3627 2222
rect 3895 2218 3899 2222
rect 3991 2218 3995 2222
rect 111 2142 115 2146
rect 151 2142 155 2146
rect 183 2142 187 2146
rect 327 2142 331 2146
rect 343 2142 347 2146
rect 495 2142 499 2146
rect 535 2142 539 2146
rect 647 2142 651 2146
rect 735 2142 739 2146
rect 791 2142 795 2146
rect 927 2142 931 2146
rect 935 2142 939 2146
rect 1071 2142 1075 2146
rect 1111 2142 1115 2146
rect 1199 2142 1203 2146
rect 1279 2142 1283 2146
rect 1335 2142 1339 2146
rect 1447 2142 1451 2146
rect 1471 2142 1475 2146
rect 1615 2142 1619 2146
rect 1783 2142 1787 2146
rect 2031 2142 2035 2146
rect 2071 2146 2075 2150
rect 2279 2146 2283 2150
rect 2391 2146 2395 2150
rect 2439 2146 2443 2150
rect 2495 2146 2499 2150
rect 2599 2146 2603 2150
rect 2623 2146 2627 2150
rect 2703 2146 2707 2150
rect 2807 2146 2811 2150
rect 2839 2146 2843 2150
rect 2911 2146 2915 2150
rect 3031 2146 3035 2150
rect 3079 2146 3083 2150
rect 3175 2146 3179 2150
rect 3343 2146 3347 2150
rect 3527 2146 3531 2150
rect 3623 2146 3627 2150
rect 3719 2146 3723 2150
rect 3895 2146 3899 2150
rect 3991 2146 3995 2150
rect 2071 2070 2075 2074
rect 2391 2070 2395 2074
rect 2487 2070 2491 2074
rect 2495 2070 2499 2074
rect 2591 2070 2595 2074
rect 2599 2070 2603 2074
rect 2695 2070 2699 2074
rect 2703 2070 2707 2074
rect 2807 2070 2811 2074
rect 2911 2070 2915 2074
rect 2935 2070 2939 2074
rect 3031 2070 3035 2074
rect 3095 2070 3099 2074
rect 3175 2070 3179 2074
rect 3279 2070 3283 2074
rect 3343 2070 3347 2074
rect 3479 2070 3483 2074
rect 3527 2070 3531 2074
rect 3695 2070 3699 2074
rect 3719 2070 3723 2074
rect 3895 2070 3899 2074
rect 3991 2070 3995 2074
rect 111 2058 115 2062
rect 151 2058 155 2062
rect 327 2058 331 2062
rect 383 2058 387 2062
rect 535 2058 539 2062
rect 631 2058 635 2062
rect 735 2058 739 2062
rect 863 2058 867 2062
rect 927 2058 931 2062
rect 1071 2058 1075 2062
rect 1111 2058 1115 2062
rect 1263 2058 1267 2062
rect 1279 2058 1283 2062
rect 1447 2058 1451 2062
rect 1615 2058 1619 2062
rect 1783 2058 1787 2062
rect 1935 2058 1939 2062
rect 2031 2058 2035 2062
rect 2071 1990 2075 1994
rect 2487 1990 2491 1994
rect 2527 1990 2531 1994
rect 2591 1990 2595 1994
rect 2695 1990 2699 1994
rect 2703 1990 2707 1994
rect 2807 1990 2811 1994
rect 2887 1990 2891 1994
rect 2935 1990 2939 1994
rect 3079 1990 3083 1994
rect 3095 1990 3099 1994
rect 3279 1990 3283 1994
rect 3479 1990 3483 1994
rect 3487 1990 3491 1994
rect 3695 1990 3699 1994
rect 3703 1990 3707 1994
rect 3895 1990 3899 1994
rect 3991 1990 3995 1994
rect 111 1974 115 1978
rect 151 1974 155 1978
rect 327 1974 331 1978
rect 383 1974 387 1978
rect 535 1974 539 1978
rect 631 1974 635 1978
rect 735 1974 739 1978
rect 863 1974 867 1978
rect 935 1974 939 1978
rect 1071 1974 1075 1978
rect 1127 1974 1131 1978
rect 1263 1974 1267 1978
rect 1303 1974 1307 1978
rect 1447 1974 1451 1978
rect 1471 1974 1475 1978
rect 1615 1974 1619 1978
rect 1631 1974 1635 1978
rect 1783 1974 1787 1978
rect 1791 1974 1795 1978
rect 1935 1974 1939 1978
rect 2031 1974 2035 1978
rect 2071 1914 2075 1918
rect 2111 1914 2115 1918
rect 2303 1914 2307 1918
rect 2519 1914 2523 1918
rect 2527 1914 2531 1918
rect 2703 1914 2707 1918
rect 2735 1914 2739 1918
rect 2887 1914 2891 1918
rect 2959 1914 2963 1918
rect 3079 1914 3083 1918
rect 3191 1914 3195 1918
rect 3279 1914 3283 1918
rect 3431 1914 3435 1918
rect 3487 1914 3491 1918
rect 3671 1914 3675 1918
rect 3703 1914 3707 1918
rect 3895 1914 3899 1918
rect 3991 1914 3995 1918
rect 111 1898 115 1902
rect 151 1898 155 1902
rect 303 1898 307 1902
rect 327 1898 331 1902
rect 463 1898 467 1902
rect 535 1898 539 1902
rect 615 1898 619 1902
rect 735 1898 739 1902
rect 767 1898 771 1902
rect 927 1898 931 1902
rect 935 1898 939 1902
rect 1103 1898 1107 1902
rect 1127 1898 1131 1902
rect 1295 1898 1299 1902
rect 1303 1898 1307 1902
rect 1471 1898 1475 1902
rect 1511 1898 1515 1902
rect 1631 1898 1635 1902
rect 1735 1898 1739 1902
rect 1791 1898 1795 1902
rect 1935 1898 1939 1902
rect 2031 1898 2035 1902
rect 2071 1842 2075 1846
rect 2111 1842 2115 1846
rect 2231 1842 2235 1846
rect 2303 1842 2307 1846
rect 2399 1842 2403 1846
rect 2519 1842 2523 1846
rect 2599 1842 2603 1846
rect 2735 1842 2739 1846
rect 2831 1842 2835 1846
rect 2959 1842 2963 1846
rect 3079 1842 3083 1846
rect 3191 1842 3195 1846
rect 3351 1842 3355 1846
rect 3431 1842 3435 1846
rect 3631 1842 3635 1846
rect 3671 1842 3675 1846
rect 3895 1842 3899 1846
rect 3991 1842 3995 1846
rect 111 1814 115 1818
rect 151 1814 155 1818
rect 303 1814 307 1818
rect 343 1814 347 1818
rect 463 1814 467 1818
rect 543 1814 547 1818
rect 615 1814 619 1818
rect 735 1814 739 1818
rect 767 1814 771 1818
rect 919 1814 923 1818
rect 927 1814 931 1818
rect 1095 1814 1099 1818
rect 1103 1814 1107 1818
rect 1271 1814 1275 1818
rect 1295 1814 1299 1818
rect 1447 1814 1451 1818
rect 1511 1814 1515 1818
rect 1623 1814 1627 1818
rect 1735 1814 1739 1818
rect 1807 1814 1811 1818
rect 1935 1814 1939 1818
rect 2031 1814 2035 1818
rect 2071 1766 2075 1770
rect 2111 1766 2115 1770
rect 2231 1766 2235 1770
rect 2239 1766 2243 1770
rect 2399 1766 2403 1770
rect 2575 1766 2579 1770
rect 2599 1766 2603 1770
rect 2751 1766 2755 1770
rect 2831 1766 2835 1770
rect 2935 1766 2939 1770
rect 3079 1766 3083 1770
rect 3127 1766 3131 1770
rect 3319 1766 3323 1770
rect 3351 1766 3355 1770
rect 3511 1766 3515 1770
rect 3631 1766 3635 1770
rect 3711 1766 3715 1770
rect 3895 1766 3899 1770
rect 3991 1766 3995 1770
rect 111 1738 115 1742
rect 151 1738 155 1742
rect 319 1738 323 1742
rect 343 1738 347 1742
rect 527 1738 531 1742
rect 543 1738 547 1742
rect 735 1738 739 1742
rect 743 1738 747 1742
rect 919 1738 923 1742
rect 959 1738 963 1742
rect 1095 1738 1099 1742
rect 1167 1738 1171 1742
rect 1271 1738 1275 1742
rect 1367 1738 1371 1742
rect 1447 1738 1451 1742
rect 1559 1738 1563 1742
rect 1623 1738 1627 1742
rect 1759 1738 1763 1742
rect 1807 1738 1811 1742
rect 1935 1738 1939 1742
rect 2031 1738 2035 1742
rect 2071 1686 2075 1690
rect 2111 1686 2115 1690
rect 2239 1686 2243 1690
rect 2311 1686 2315 1690
rect 2399 1686 2403 1690
rect 2527 1686 2531 1690
rect 2575 1686 2579 1690
rect 2743 1686 2747 1690
rect 2751 1686 2755 1690
rect 2935 1686 2939 1690
rect 2951 1686 2955 1690
rect 3127 1686 3131 1690
rect 3151 1686 3155 1690
rect 3319 1686 3323 1690
rect 3343 1686 3347 1690
rect 3511 1686 3515 1690
rect 3527 1686 3531 1690
rect 3711 1686 3715 1690
rect 3719 1686 3723 1690
rect 3895 1686 3899 1690
rect 3991 1686 3995 1690
rect 111 1666 115 1670
rect 151 1666 155 1670
rect 319 1666 323 1670
rect 503 1666 507 1670
rect 527 1666 531 1670
rect 695 1666 699 1670
rect 743 1666 747 1670
rect 887 1666 891 1670
rect 959 1666 963 1670
rect 1079 1666 1083 1670
rect 1167 1666 1171 1670
rect 1263 1666 1267 1670
rect 1367 1666 1371 1670
rect 1439 1666 1443 1670
rect 1559 1666 1563 1670
rect 1615 1666 1619 1670
rect 1759 1666 1763 1670
rect 1791 1666 1795 1670
rect 1935 1666 1939 1670
rect 2031 1666 2035 1670
rect 2071 1602 2075 1606
rect 2111 1602 2115 1606
rect 2311 1602 2315 1606
rect 2479 1602 2483 1606
rect 2527 1602 2531 1606
rect 2583 1602 2587 1606
rect 2695 1602 2699 1606
rect 2743 1602 2747 1606
rect 2815 1602 2819 1606
rect 2943 1602 2947 1606
rect 2951 1602 2955 1606
rect 3079 1602 3083 1606
rect 3151 1602 3155 1606
rect 3223 1602 3227 1606
rect 3343 1602 3347 1606
rect 3383 1602 3387 1606
rect 3527 1602 3531 1606
rect 3551 1602 3555 1606
rect 3719 1602 3723 1606
rect 3727 1602 3731 1606
rect 3895 1602 3899 1606
rect 3991 1602 3995 1606
rect 111 1586 115 1590
rect 151 1586 155 1590
rect 319 1586 323 1590
rect 455 1586 459 1590
rect 503 1586 507 1590
rect 599 1586 603 1590
rect 695 1586 699 1590
rect 743 1586 747 1590
rect 887 1586 891 1590
rect 1031 1586 1035 1590
rect 1079 1586 1083 1590
rect 1175 1586 1179 1590
rect 1263 1586 1267 1590
rect 1319 1586 1323 1590
rect 1439 1586 1443 1590
rect 1471 1586 1475 1590
rect 1615 1586 1619 1590
rect 1623 1586 1627 1590
rect 1791 1586 1795 1590
rect 2031 1586 2035 1590
rect 2071 1518 2075 1522
rect 2479 1518 2483 1522
rect 2487 1518 2491 1522
rect 2583 1518 2587 1522
rect 2591 1518 2595 1522
rect 2695 1518 2699 1522
rect 2807 1518 2811 1522
rect 2815 1518 2819 1522
rect 2935 1518 2939 1522
rect 2943 1518 2947 1522
rect 3071 1518 3075 1522
rect 3079 1518 3083 1522
rect 3223 1518 3227 1522
rect 3383 1518 3387 1522
rect 3551 1518 3555 1522
rect 3719 1518 3723 1522
rect 3727 1518 3731 1522
rect 3895 1518 3899 1522
rect 3991 1518 3995 1522
rect 111 1506 115 1510
rect 319 1506 323 1510
rect 359 1506 363 1510
rect 455 1506 459 1510
rect 487 1506 491 1510
rect 599 1506 603 1510
rect 623 1506 627 1510
rect 743 1506 747 1510
rect 775 1506 779 1510
rect 887 1506 891 1510
rect 927 1506 931 1510
rect 1031 1506 1035 1510
rect 1087 1506 1091 1510
rect 1175 1506 1179 1510
rect 1255 1506 1259 1510
rect 1319 1506 1323 1510
rect 1423 1506 1427 1510
rect 1471 1506 1475 1510
rect 1591 1506 1595 1510
rect 1623 1506 1627 1510
rect 1767 1506 1771 1510
rect 2031 1506 2035 1510
rect 2071 1442 2075 1446
rect 2239 1442 2243 1446
rect 2351 1442 2355 1446
rect 2471 1442 2475 1446
rect 2487 1442 2491 1446
rect 2591 1442 2595 1446
rect 2695 1442 2699 1446
rect 2727 1442 2731 1446
rect 2807 1442 2811 1446
rect 2879 1442 2883 1446
rect 2935 1442 2939 1446
rect 3055 1442 3059 1446
rect 3071 1442 3075 1446
rect 3223 1442 3227 1446
rect 3247 1442 3251 1446
rect 3383 1442 3387 1446
rect 3455 1442 3459 1446
rect 3551 1442 3555 1446
rect 3671 1442 3675 1446
rect 3719 1442 3723 1446
rect 3887 1442 3891 1446
rect 3895 1442 3899 1446
rect 3991 1442 3995 1446
rect 111 1426 115 1430
rect 151 1426 155 1430
rect 271 1426 275 1430
rect 359 1426 363 1430
rect 431 1426 435 1430
rect 487 1426 491 1430
rect 615 1426 619 1430
rect 623 1426 627 1430
rect 775 1426 779 1430
rect 807 1426 811 1430
rect 927 1426 931 1430
rect 1007 1426 1011 1430
rect 1087 1426 1091 1430
rect 1215 1426 1219 1430
rect 1255 1426 1259 1430
rect 1423 1426 1427 1430
rect 1591 1426 1595 1430
rect 1631 1426 1635 1430
rect 1767 1426 1771 1430
rect 1847 1426 1851 1430
rect 2031 1426 2035 1430
rect 2071 1362 2075 1366
rect 2239 1362 2243 1366
rect 2351 1362 2355 1366
rect 2391 1362 2395 1366
rect 2471 1362 2475 1366
rect 2527 1362 2531 1366
rect 2591 1362 2595 1366
rect 2679 1362 2683 1366
rect 2727 1362 2731 1366
rect 2839 1362 2843 1366
rect 2879 1362 2883 1366
rect 2999 1362 3003 1366
rect 3055 1362 3059 1366
rect 3167 1362 3171 1366
rect 3247 1362 3251 1366
rect 3343 1362 3347 1366
rect 3455 1362 3459 1366
rect 3519 1362 3523 1366
rect 3671 1362 3675 1366
rect 3695 1362 3699 1366
rect 3879 1362 3883 1366
rect 3887 1362 3891 1366
rect 3991 1362 3995 1366
rect 111 1342 115 1346
rect 151 1342 155 1346
rect 271 1342 275 1346
rect 287 1342 291 1346
rect 431 1342 435 1346
rect 463 1342 467 1346
rect 615 1342 619 1346
rect 663 1342 667 1346
rect 807 1342 811 1346
rect 863 1342 867 1346
rect 1007 1342 1011 1346
rect 1063 1342 1067 1346
rect 1215 1342 1219 1346
rect 1255 1342 1259 1346
rect 1423 1342 1427 1346
rect 1431 1342 1435 1346
rect 1607 1342 1611 1346
rect 1631 1342 1635 1346
rect 1783 1342 1787 1346
rect 1847 1342 1851 1346
rect 1935 1342 1939 1346
rect 2031 1342 2035 1346
rect 2071 1282 2075 1286
rect 2111 1282 2115 1286
rect 2343 1282 2347 1286
rect 2391 1282 2395 1286
rect 2527 1282 2531 1286
rect 2583 1282 2587 1286
rect 2679 1282 2683 1286
rect 2799 1282 2803 1286
rect 2839 1282 2843 1286
rect 2999 1282 3003 1286
rect 3167 1282 3171 1286
rect 3183 1282 3187 1286
rect 3343 1282 3347 1286
rect 3495 1282 3499 1286
rect 3519 1282 3523 1286
rect 3639 1282 3643 1286
rect 3695 1282 3699 1286
rect 3775 1282 3779 1286
rect 3879 1282 3883 1286
rect 3895 1282 3899 1286
rect 3991 1282 3995 1286
rect 111 1270 115 1274
rect 151 1270 155 1274
rect 207 1270 211 1274
rect 287 1270 291 1274
rect 327 1270 331 1274
rect 455 1270 459 1274
rect 463 1270 467 1274
rect 583 1270 587 1274
rect 663 1270 667 1274
rect 719 1270 723 1274
rect 863 1270 867 1274
rect 879 1270 883 1274
rect 1055 1270 1059 1274
rect 1063 1270 1067 1274
rect 1255 1270 1259 1274
rect 1263 1270 1267 1274
rect 1431 1270 1435 1274
rect 1487 1270 1491 1274
rect 1607 1270 1611 1274
rect 1719 1270 1723 1274
rect 1783 1270 1787 1274
rect 1935 1270 1939 1274
rect 2031 1270 2035 1274
rect 2071 1206 2075 1210
rect 2111 1206 2115 1210
rect 2279 1206 2283 1210
rect 2343 1206 2347 1210
rect 2471 1206 2475 1210
rect 2583 1206 2587 1210
rect 2655 1206 2659 1210
rect 2799 1206 2803 1210
rect 2831 1206 2835 1210
rect 2999 1206 3003 1210
rect 3159 1206 3163 1210
rect 3183 1206 3187 1210
rect 3327 1206 3331 1210
rect 3343 1206 3347 1210
rect 3495 1206 3499 1210
rect 3639 1206 3643 1210
rect 3775 1206 3779 1210
rect 3895 1206 3899 1210
rect 3991 1206 3995 1210
rect 111 1190 115 1194
rect 207 1190 211 1194
rect 327 1190 331 1194
rect 455 1190 459 1194
rect 471 1190 475 1194
rect 583 1190 587 1194
rect 703 1190 707 1194
rect 719 1190 723 1194
rect 823 1190 827 1194
rect 879 1190 883 1194
rect 943 1190 947 1194
rect 1055 1190 1059 1194
rect 1063 1190 1067 1194
rect 1183 1190 1187 1194
rect 1263 1190 1267 1194
rect 1303 1190 1307 1194
rect 1423 1190 1427 1194
rect 1487 1190 1491 1194
rect 1543 1190 1547 1194
rect 1719 1190 1723 1194
rect 1935 1190 1939 1194
rect 2031 1190 2035 1194
rect 2071 1130 2075 1134
rect 2111 1130 2115 1134
rect 2279 1130 2283 1134
rect 2295 1130 2299 1134
rect 2471 1130 2475 1134
rect 2503 1130 2507 1134
rect 2655 1130 2659 1134
rect 2703 1130 2707 1134
rect 2831 1130 2835 1134
rect 2895 1130 2899 1134
rect 2999 1130 3003 1134
rect 3079 1130 3083 1134
rect 3159 1130 3163 1134
rect 3255 1130 3259 1134
rect 3327 1130 3331 1134
rect 3431 1130 3435 1134
rect 3495 1130 3499 1134
rect 3615 1130 3619 1134
rect 3991 1130 3995 1134
rect 111 1110 115 1114
rect 471 1110 475 1114
rect 583 1110 587 1114
rect 623 1110 627 1114
rect 703 1110 707 1114
rect 735 1110 739 1114
rect 823 1110 827 1114
rect 855 1110 859 1114
rect 943 1110 947 1114
rect 975 1110 979 1114
rect 1063 1110 1067 1114
rect 1095 1110 1099 1114
rect 1183 1110 1187 1114
rect 1215 1110 1219 1114
rect 1303 1110 1307 1114
rect 1335 1110 1339 1114
rect 1423 1110 1427 1114
rect 1455 1110 1459 1114
rect 1543 1110 1547 1114
rect 1575 1110 1579 1114
rect 1703 1110 1707 1114
rect 2031 1110 2035 1114
rect 2071 1050 2075 1054
rect 2111 1050 2115 1054
rect 2167 1050 2171 1054
rect 2287 1050 2291 1054
rect 2295 1050 2299 1054
rect 2423 1050 2427 1054
rect 2503 1050 2507 1054
rect 2575 1050 2579 1054
rect 2703 1050 2707 1054
rect 2743 1050 2747 1054
rect 2895 1050 2899 1054
rect 2919 1050 2923 1054
rect 3079 1050 3083 1054
rect 3095 1050 3099 1054
rect 3255 1050 3259 1054
rect 3279 1050 3283 1054
rect 3431 1050 3435 1054
rect 3463 1050 3467 1054
rect 3615 1050 3619 1054
rect 3655 1050 3659 1054
rect 3991 1050 3995 1054
rect 111 1030 115 1034
rect 623 1030 627 1034
rect 727 1030 731 1034
rect 735 1030 739 1034
rect 847 1030 851 1034
rect 855 1030 859 1034
rect 967 1030 971 1034
rect 975 1030 979 1034
rect 1095 1030 1099 1034
rect 1215 1030 1219 1034
rect 1223 1030 1227 1034
rect 1335 1030 1339 1034
rect 1351 1030 1355 1034
rect 1455 1030 1459 1034
rect 1479 1030 1483 1034
rect 1575 1030 1579 1034
rect 1607 1030 1611 1034
rect 1703 1030 1707 1034
rect 1735 1030 1739 1034
rect 1863 1030 1867 1034
rect 2031 1030 2035 1034
rect 2071 970 2075 974
rect 2167 970 2171 974
rect 2287 970 2291 974
rect 2423 970 2427 974
rect 2527 970 2531 974
rect 2575 970 2579 974
rect 2647 970 2651 974
rect 2743 970 2747 974
rect 2775 970 2779 974
rect 2919 970 2923 974
rect 3071 970 3075 974
rect 3095 970 3099 974
rect 3231 970 3235 974
rect 3279 970 3283 974
rect 3399 970 3403 974
rect 3463 970 3467 974
rect 3567 970 3571 974
rect 3655 970 3659 974
rect 3735 970 3739 974
rect 3991 970 3995 974
rect 111 950 115 954
rect 591 950 595 954
rect 727 950 731 954
rect 735 950 739 954
rect 847 950 851 954
rect 887 950 891 954
rect 967 950 971 954
rect 1039 950 1043 954
rect 1095 950 1099 954
rect 1199 950 1203 954
rect 1223 950 1227 954
rect 1351 950 1355 954
rect 1479 950 1483 954
rect 1503 950 1507 954
rect 1607 950 1611 954
rect 1655 950 1659 954
rect 1735 950 1739 954
rect 1807 950 1811 954
rect 1863 950 1867 954
rect 1935 950 1939 954
rect 2031 950 2035 954
rect 2071 886 2075 890
rect 2455 886 2459 890
rect 2527 886 2531 890
rect 2575 886 2579 890
rect 2647 886 2651 890
rect 2711 886 2715 890
rect 2775 886 2779 890
rect 2863 886 2867 890
rect 2919 886 2923 890
rect 3015 886 3019 890
rect 3071 886 3075 890
rect 3167 886 3171 890
rect 3231 886 3235 890
rect 3319 886 3323 890
rect 3399 886 3403 890
rect 3471 886 3475 890
rect 3567 886 3571 890
rect 3615 886 3619 890
rect 3735 886 3739 890
rect 3767 886 3771 890
rect 3895 886 3899 890
rect 3991 886 3995 890
rect 111 870 115 874
rect 439 870 443 874
rect 583 870 587 874
rect 591 870 595 874
rect 735 870 739 874
rect 887 870 891 874
rect 1039 870 1043 874
rect 1047 870 1051 874
rect 1199 870 1203 874
rect 1351 870 1355 874
rect 1495 870 1499 874
rect 1503 870 1507 874
rect 1647 870 1651 874
rect 1655 870 1659 874
rect 1799 870 1803 874
rect 1807 870 1811 874
rect 1935 870 1939 874
rect 2031 870 2035 874
rect 2071 814 2075 818
rect 2215 814 2219 818
rect 2343 814 2347 818
rect 2455 814 2459 818
rect 2479 814 2483 818
rect 2575 814 2579 818
rect 2623 814 2627 818
rect 2711 814 2715 818
rect 2783 814 2787 818
rect 2863 814 2867 818
rect 2959 814 2963 818
rect 3015 814 3019 818
rect 3167 814 3171 818
rect 3319 814 3323 818
rect 3391 814 3395 818
rect 3471 814 3475 818
rect 3615 814 3619 818
rect 3623 814 3627 818
rect 3767 814 3771 818
rect 3863 814 3867 818
rect 3895 814 3899 818
rect 3991 814 3995 818
rect 111 798 115 802
rect 279 798 283 802
rect 431 798 435 802
rect 439 798 443 802
rect 583 798 587 802
rect 591 798 595 802
rect 735 798 739 802
rect 751 798 755 802
rect 887 798 891 802
rect 919 798 923 802
rect 1047 798 1051 802
rect 1087 798 1091 802
rect 1199 798 1203 802
rect 1255 798 1259 802
rect 1351 798 1355 802
rect 1423 798 1427 802
rect 1495 798 1499 802
rect 1591 798 1595 802
rect 1647 798 1651 802
rect 1799 798 1803 802
rect 2031 798 2035 802
rect 2071 734 2075 738
rect 2111 734 2115 738
rect 2215 734 2219 738
rect 2247 734 2251 738
rect 2343 734 2347 738
rect 2423 734 2427 738
rect 2479 734 2483 738
rect 2599 734 2603 738
rect 2623 734 2627 738
rect 2783 734 2787 738
rect 2959 734 2963 738
rect 2967 734 2971 738
rect 3151 734 3155 738
rect 3167 734 3171 738
rect 3335 734 3339 738
rect 3391 734 3395 738
rect 3519 734 3523 738
rect 3623 734 3627 738
rect 3703 734 3707 738
rect 3863 734 3867 738
rect 3895 734 3899 738
rect 3991 734 3995 738
rect 111 722 115 726
rect 151 722 155 726
rect 271 722 275 726
rect 279 722 283 726
rect 423 722 427 726
rect 431 722 435 726
rect 575 722 579 726
rect 591 722 595 726
rect 735 722 739 726
rect 751 722 755 726
rect 887 722 891 726
rect 919 722 923 726
rect 1039 722 1043 726
rect 1087 722 1091 726
rect 1191 722 1195 726
rect 1255 722 1259 726
rect 1343 722 1347 726
rect 1423 722 1427 726
rect 1495 722 1499 726
rect 1591 722 1595 726
rect 2031 722 2035 726
rect 2071 658 2075 662
rect 2111 658 2115 662
rect 2247 658 2251 662
rect 2375 658 2379 662
rect 2423 658 2427 662
rect 2599 658 2603 662
rect 2655 658 2659 662
rect 2783 658 2787 662
rect 2919 658 2923 662
rect 2967 658 2971 662
rect 3151 658 3155 662
rect 3175 658 3179 662
rect 3335 658 3339 662
rect 3423 658 3427 662
rect 3519 658 3523 662
rect 3671 658 3675 662
rect 3703 658 3707 662
rect 3895 658 3899 662
rect 3991 658 3995 662
rect 111 642 115 646
rect 151 642 155 646
rect 255 642 259 646
rect 271 642 275 646
rect 391 642 395 646
rect 423 642 427 646
rect 527 642 531 646
rect 575 642 579 646
rect 663 642 667 646
rect 735 642 739 646
rect 807 642 811 646
rect 887 642 891 646
rect 959 642 963 646
rect 1039 642 1043 646
rect 1119 642 1123 646
rect 1191 642 1195 646
rect 1287 642 1291 646
rect 1343 642 1347 646
rect 1455 642 1459 646
rect 1495 642 1499 646
rect 1623 642 1627 646
rect 1791 642 1795 646
rect 1935 642 1939 646
rect 2031 642 2035 646
rect 2071 574 2075 578
rect 2111 574 2115 578
rect 2215 574 2219 578
rect 2351 574 2355 578
rect 2375 574 2379 578
rect 2487 574 2491 578
rect 2631 574 2635 578
rect 2655 574 2659 578
rect 2791 574 2795 578
rect 2919 574 2923 578
rect 2975 574 2979 578
rect 3175 574 3179 578
rect 3191 574 3195 578
rect 3423 574 3427 578
rect 3671 574 3675 578
rect 3895 574 3899 578
rect 3991 574 3995 578
rect 111 558 115 562
rect 151 558 155 562
rect 207 558 211 562
rect 255 558 259 562
rect 327 558 331 562
rect 391 558 395 562
rect 447 558 451 562
rect 527 558 531 562
rect 567 558 571 562
rect 663 558 667 562
rect 687 558 691 562
rect 799 558 803 562
rect 807 558 811 562
rect 911 558 915 562
rect 959 558 963 562
rect 1031 558 1035 562
rect 1119 558 1123 562
rect 1151 558 1155 562
rect 1271 558 1275 562
rect 1287 558 1291 562
rect 1455 558 1459 562
rect 1623 558 1627 562
rect 1791 558 1795 562
rect 1935 558 1939 562
rect 2031 558 2035 562
rect 2071 498 2075 502
rect 2111 498 2115 502
rect 2215 498 2219 502
rect 2351 498 2355 502
rect 2423 498 2427 502
rect 2487 498 2491 502
rect 2527 498 2531 502
rect 2631 498 2635 502
rect 2743 498 2747 502
rect 2791 498 2795 502
rect 2871 498 2875 502
rect 2975 498 2979 502
rect 3031 498 3035 502
rect 3191 498 3195 502
rect 3223 498 3227 502
rect 3423 498 3427 502
rect 3447 498 3451 502
rect 3671 498 3675 502
rect 3679 498 3683 502
rect 3895 498 3899 502
rect 3991 498 3995 502
rect 111 478 115 482
rect 207 478 211 482
rect 327 478 331 482
rect 439 478 443 482
rect 447 478 451 482
rect 543 478 547 482
rect 567 478 571 482
rect 647 478 651 482
rect 687 478 691 482
rect 751 478 755 482
rect 799 478 803 482
rect 855 478 859 482
rect 911 478 915 482
rect 959 478 963 482
rect 1031 478 1035 482
rect 1063 478 1067 482
rect 1151 478 1155 482
rect 1167 478 1171 482
rect 1271 478 1275 482
rect 1375 478 1379 482
rect 2031 478 2035 482
rect 2071 422 2075 426
rect 2423 422 2427 426
rect 2527 422 2531 426
rect 2631 422 2635 426
rect 2639 422 2643 426
rect 2743 422 2747 426
rect 2775 422 2779 426
rect 2871 422 2875 426
rect 2951 422 2955 426
rect 3031 422 3035 426
rect 3159 422 3163 426
rect 3223 422 3227 426
rect 3399 422 3403 426
rect 3447 422 3451 426
rect 3655 422 3659 426
rect 3679 422 3683 426
rect 3895 422 3899 426
rect 3991 422 3995 426
rect 111 398 115 402
rect 439 398 443 402
rect 543 398 547 402
rect 623 398 627 402
rect 647 398 651 402
rect 727 398 731 402
rect 751 398 755 402
rect 831 398 835 402
rect 855 398 859 402
rect 935 398 939 402
rect 959 398 963 402
rect 1039 398 1043 402
rect 1063 398 1067 402
rect 1143 398 1147 402
rect 1167 398 1171 402
rect 1247 398 1251 402
rect 1271 398 1275 402
rect 1351 398 1355 402
rect 1375 398 1379 402
rect 1455 398 1459 402
rect 1559 398 1563 402
rect 2031 398 2035 402
rect 2071 338 2075 342
rect 2271 338 2275 342
rect 2423 338 2427 342
rect 2527 338 2531 342
rect 2583 338 2587 342
rect 2639 338 2643 342
rect 2743 338 2747 342
rect 2775 338 2779 342
rect 2911 338 2915 342
rect 2951 338 2955 342
rect 3071 338 3075 342
rect 3159 338 3163 342
rect 3223 338 3227 342
rect 3367 338 3371 342
rect 3399 338 3403 342
rect 3503 338 3507 342
rect 3639 338 3643 342
rect 3655 338 3659 342
rect 3775 338 3779 342
rect 3895 338 3899 342
rect 3991 338 3995 342
rect 111 326 115 330
rect 399 326 403 330
rect 543 326 547 330
rect 623 326 627 330
rect 687 326 691 330
rect 727 326 731 330
rect 831 326 835 330
rect 839 326 843 330
rect 935 326 939 330
rect 991 326 995 330
rect 1039 326 1043 330
rect 1143 326 1147 330
rect 1247 326 1251 330
rect 1303 326 1307 330
rect 1351 326 1355 330
rect 1455 326 1459 330
rect 1463 326 1467 330
rect 1559 326 1563 330
rect 1623 326 1627 330
rect 2031 326 2035 330
rect 2071 258 2075 262
rect 2111 258 2115 262
rect 2247 258 2251 262
rect 2271 258 2275 262
rect 2423 258 2427 262
rect 2583 258 2587 262
rect 2599 258 2603 262
rect 2743 258 2747 262
rect 2775 258 2779 262
rect 2911 258 2915 262
rect 2943 258 2947 262
rect 3071 258 3075 262
rect 3103 258 3107 262
rect 3223 258 3227 262
rect 3255 258 3259 262
rect 3367 258 3371 262
rect 3391 258 3395 262
rect 3503 258 3507 262
rect 3527 258 3531 262
rect 3639 258 3643 262
rect 3655 258 3659 262
rect 3775 258 3779 262
rect 3783 258 3787 262
rect 3895 258 3899 262
rect 3991 258 3995 262
rect 111 250 115 254
rect 207 250 211 254
rect 399 250 403 254
rect 431 250 435 254
rect 543 250 547 254
rect 655 250 659 254
rect 687 250 691 254
rect 839 250 843 254
rect 871 250 875 254
rect 991 250 995 254
rect 1071 250 1075 254
rect 1143 250 1147 254
rect 1263 250 1267 254
rect 1303 250 1307 254
rect 1447 250 1451 254
rect 1463 250 1467 254
rect 1623 250 1627 254
rect 1631 250 1635 254
rect 1815 250 1819 254
rect 2031 250 2035 254
rect 2071 174 2075 178
rect 2111 174 2115 178
rect 2239 174 2243 178
rect 2247 174 2251 178
rect 2399 174 2403 178
rect 2423 174 2427 178
rect 2567 174 2571 178
rect 2599 174 2603 178
rect 2735 174 2739 178
rect 2775 174 2779 178
rect 2895 174 2899 178
rect 2943 174 2947 178
rect 3047 174 3051 178
rect 3103 174 3107 178
rect 3191 174 3195 178
rect 3255 174 3259 178
rect 3327 174 3331 178
rect 3391 174 3395 178
rect 3455 174 3459 178
rect 3527 174 3531 178
rect 3591 174 3595 178
rect 3655 174 3659 178
rect 3727 174 3731 178
rect 3783 174 3787 178
rect 3895 174 3899 178
rect 3991 174 3995 178
rect 111 150 115 154
rect 151 150 155 154
rect 207 150 211 154
rect 255 150 259 154
rect 359 150 363 154
rect 431 150 435 154
rect 463 150 467 154
rect 567 150 571 154
rect 655 150 659 154
rect 671 150 675 154
rect 775 150 779 154
rect 871 150 875 154
rect 879 150 883 154
rect 983 150 987 154
rect 1071 150 1075 154
rect 1087 150 1091 154
rect 1191 150 1195 154
rect 1263 150 1267 154
rect 1295 150 1299 154
rect 1399 150 1403 154
rect 1447 150 1451 154
rect 1511 150 1515 154
rect 1623 150 1627 154
rect 1631 150 1635 154
rect 1727 150 1731 154
rect 1815 150 1819 154
rect 1831 150 1835 154
rect 1935 150 1939 154
rect 2031 150 2035 154
rect 2071 102 2075 106
rect 2111 102 2115 106
rect 2239 102 2243 106
rect 2399 102 2403 106
rect 2567 102 2571 106
rect 2735 102 2739 106
rect 2895 102 2899 106
rect 3047 102 3051 106
rect 3191 102 3195 106
rect 3327 102 3331 106
rect 3455 102 3459 106
rect 3591 102 3595 106
rect 3727 102 3731 106
rect 3991 102 3995 106
rect 111 78 115 82
rect 151 78 155 82
rect 255 78 259 82
rect 359 78 363 82
rect 463 78 467 82
rect 567 78 571 82
rect 671 78 675 82
rect 775 78 779 82
rect 879 78 883 82
rect 983 78 987 82
rect 1087 78 1091 82
rect 1191 78 1195 82
rect 1295 78 1299 82
rect 1399 78 1403 82
rect 1511 78 1515 82
rect 1623 78 1627 82
rect 1727 78 1731 82
rect 1831 78 1835 82
rect 1935 78 1939 82
rect 2031 78 2035 82
<< m4 >>
rect 2054 4077 2055 4083
rect 2061 4082 4027 4083
rect 2061 4078 2071 4082
rect 2075 4078 3399 4082
rect 3403 4078 3503 4082
rect 3507 4078 3607 4082
rect 3611 4078 3711 4082
rect 3715 4078 3991 4082
rect 3995 4078 4027 4082
rect 2061 4077 4027 4078
rect 4033 4077 4034 4083
rect 96 4041 97 4047
rect 103 4046 2055 4047
rect 103 4042 111 4046
rect 115 4042 495 4046
rect 499 4042 599 4046
rect 603 4042 703 4046
rect 707 4042 807 4046
rect 811 4042 911 4046
rect 915 4042 1015 4046
rect 1019 4042 1119 4046
rect 1123 4042 1223 4046
rect 1227 4042 1327 4046
rect 1331 4042 1431 4046
rect 1435 4042 2031 4046
rect 2035 4042 2055 4046
rect 103 4041 2055 4042
rect 2061 4041 2062 4047
rect 2042 4005 2043 4011
rect 2049 4010 4015 4011
rect 2049 4006 2071 4010
rect 2075 4006 2111 4010
rect 2115 4006 2215 4010
rect 2219 4006 2319 4010
rect 2323 4006 2423 4010
rect 2427 4006 2527 4010
rect 2531 4006 2647 4010
rect 2651 4006 2775 4010
rect 2779 4006 2903 4010
rect 2907 4006 3031 4010
rect 3035 4006 3159 4010
rect 3163 4006 3287 4010
rect 3291 4006 3399 4010
rect 3403 4006 3415 4010
rect 3419 4006 3503 4010
rect 3507 4006 3551 4010
rect 3555 4006 3607 4010
rect 3611 4006 3711 4010
rect 3715 4006 3991 4010
rect 3995 4006 4015 4010
rect 2049 4005 4015 4006
rect 4021 4005 4022 4011
rect 84 3969 85 3975
rect 91 3974 2043 3975
rect 91 3970 111 3974
rect 115 3970 391 3974
rect 395 3970 495 3974
rect 499 3970 599 3974
rect 603 3970 703 3974
rect 707 3970 807 3974
rect 811 3970 911 3974
rect 915 3970 1015 3974
rect 1019 3970 1119 3974
rect 1123 3970 1223 3974
rect 1227 3970 1327 3974
rect 1331 3970 1431 3974
rect 1435 3970 1535 3974
rect 1539 3970 2031 3974
rect 2035 3970 2043 3974
rect 91 3969 2043 3970
rect 2049 3969 2050 3975
rect 2054 3929 2055 3935
rect 2061 3934 4027 3935
rect 2061 3930 2071 3934
rect 2075 3930 2111 3934
rect 2115 3930 2143 3934
rect 2147 3930 2215 3934
rect 2219 3930 2319 3934
rect 2323 3930 2423 3934
rect 2427 3930 2487 3934
rect 2491 3930 2527 3934
rect 2531 3930 2647 3934
rect 2651 3930 2775 3934
rect 2779 3930 2799 3934
rect 2803 3930 2903 3934
rect 2907 3930 2951 3934
rect 2955 3930 3031 3934
rect 3035 3930 3103 3934
rect 3107 3930 3159 3934
rect 3163 3930 3255 3934
rect 3259 3930 3287 3934
rect 3291 3930 3415 3934
rect 3419 3930 3551 3934
rect 3555 3930 3991 3934
rect 3995 3930 4027 3934
rect 2061 3929 4027 3930
rect 4033 3929 4034 3935
rect 96 3893 97 3899
rect 103 3898 2055 3899
rect 103 3894 111 3898
rect 115 3894 375 3898
rect 379 3894 391 3898
rect 395 3894 495 3898
rect 499 3894 599 3898
rect 603 3894 623 3898
rect 627 3894 703 3898
rect 707 3894 759 3898
rect 763 3894 807 3898
rect 811 3894 895 3898
rect 899 3894 911 3898
rect 915 3894 1015 3898
rect 1019 3894 1023 3898
rect 1027 3894 1119 3898
rect 1123 3894 1151 3898
rect 1155 3894 1223 3898
rect 1227 3894 1279 3898
rect 1283 3894 1327 3898
rect 1331 3894 1415 3898
rect 1419 3894 1431 3898
rect 1435 3894 1535 3898
rect 1539 3894 1551 3898
rect 1555 3894 2031 3898
rect 2035 3894 2055 3898
rect 103 3893 2055 3894
rect 2061 3893 2062 3899
rect 2042 3857 2043 3863
rect 2049 3862 4015 3863
rect 2049 3858 2071 3862
rect 2075 3858 2119 3862
rect 2123 3858 2143 3862
rect 2147 3858 2287 3862
rect 2291 3858 2319 3862
rect 2323 3858 2447 3862
rect 2451 3858 2487 3862
rect 2491 3858 2599 3862
rect 2603 3858 2647 3862
rect 2651 3858 2743 3862
rect 2747 3858 2799 3862
rect 2803 3858 2879 3862
rect 2883 3858 2951 3862
rect 2955 3858 3023 3862
rect 3027 3858 3103 3862
rect 3107 3858 3167 3862
rect 3171 3858 3255 3862
rect 3259 3858 3991 3862
rect 3995 3858 4015 3862
rect 2049 3857 4015 3858
rect 4021 3857 4022 3863
rect 84 3813 85 3819
rect 91 3818 2043 3819
rect 91 3814 111 3818
rect 115 3814 375 3818
rect 379 3814 431 3818
rect 435 3814 495 3818
rect 499 3814 575 3818
rect 579 3814 623 3818
rect 627 3814 719 3818
rect 723 3814 759 3818
rect 763 3814 863 3818
rect 867 3814 895 3818
rect 899 3814 999 3818
rect 1003 3814 1023 3818
rect 1027 3814 1135 3818
rect 1139 3814 1151 3818
rect 1155 3814 1271 3818
rect 1275 3814 1279 3818
rect 1283 3814 1407 3818
rect 1411 3814 1415 3818
rect 1419 3814 1551 3818
rect 1555 3814 2031 3818
rect 2035 3814 2043 3818
rect 91 3813 2043 3814
rect 2049 3813 2050 3819
rect 2054 3781 2055 3787
rect 2061 3786 4027 3787
rect 2061 3782 2071 3786
rect 2075 3782 2111 3786
rect 2115 3782 2119 3786
rect 2123 3782 2239 3786
rect 2243 3782 2287 3786
rect 2291 3782 2391 3786
rect 2395 3782 2447 3786
rect 2451 3782 2543 3786
rect 2547 3782 2599 3786
rect 2603 3782 2687 3786
rect 2691 3782 2743 3786
rect 2747 3782 2823 3786
rect 2827 3782 2879 3786
rect 2883 3782 2951 3786
rect 2955 3782 3023 3786
rect 3027 3782 3087 3786
rect 3091 3782 3167 3786
rect 3171 3782 3223 3786
rect 3227 3782 3991 3786
rect 3995 3782 4027 3786
rect 2061 3781 4027 3782
rect 4033 3781 4034 3787
rect 96 3733 97 3739
rect 103 3738 2055 3739
rect 103 3734 111 3738
rect 115 3734 359 3738
rect 363 3734 431 3738
rect 435 3734 495 3738
rect 499 3734 575 3738
rect 579 3734 631 3738
rect 635 3734 719 3738
rect 723 3734 775 3738
rect 779 3734 863 3738
rect 867 3734 919 3738
rect 923 3734 999 3738
rect 1003 3734 1071 3738
rect 1075 3734 1135 3738
rect 1139 3734 1223 3738
rect 1227 3734 1271 3738
rect 1275 3734 1375 3738
rect 1379 3734 1407 3738
rect 1411 3734 1527 3738
rect 1531 3734 1551 3738
rect 1555 3734 2031 3738
rect 2035 3734 2055 3738
rect 103 3733 2055 3734
rect 2061 3733 2062 3739
rect 2042 3701 2043 3707
rect 2049 3706 4015 3707
rect 2049 3702 2071 3706
rect 2075 3702 2111 3706
rect 2115 3702 2239 3706
rect 2243 3702 2295 3706
rect 2299 3702 2391 3706
rect 2395 3702 2487 3706
rect 2491 3702 2543 3706
rect 2547 3702 2671 3706
rect 2675 3702 2687 3706
rect 2691 3702 2823 3706
rect 2827 3702 2847 3706
rect 2851 3702 2951 3706
rect 2955 3702 3015 3706
rect 3019 3702 3087 3706
rect 3091 3702 3183 3706
rect 3187 3702 3223 3706
rect 3227 3702 3359 3706
rect 3363 3702 3991 3706
rect 3995 3702 4015 3706
rect 2049 3701 4015 3702
rect 4021 3701 4022 3707
rect 84 3661 85 3667
rect 91 3666 2043 3667
rect 91 3662 111 3666
rect 115 3662 343 3666
rect 347 3662 359 3666
rect 363 3662 495 3666
rect 499 3662 519 3666
rect 523 3662 631 3666
rect 635 3662 695 3666
rect 699 3662 775 3666
rect 779 3662 863 3666
rect 867 3662 919 3666
rect 923 3662 1031 3666
rect 1035 3662 1071 3666
rect 1075 3662 1191 3666
rect 1195 3662 1223 3666
rect 1227 3662 1343 3666
rect 1347 3662 1375 3666
rect 1379 3662 1495 3666
rect 1499 3662 1527 3666
rect 1531 3662 1655 3666
rect 1659 3662 2031 3666
rect 2035 3662 2043 3666
rect 91 3661 2043 3662
rect 2049 3661 2050 3667
rect 2054 3621 2055 3627
rect 2061 3626 4027 3627
rect 2061 3622 2071 3626
rect 2075 3622 2111 3626
rect 2115 3622 2295 3626
rect 2299 3622 2487 3626
rect 2491 3622 2495 3626
rect 2499 3622 2671 3626
rect 2675 3622 2687 3626
rect 2691 3622 2847 3626
rect 2851 3622 2863 3626
rect 2867 3622 3015 3626
rect 3019 3622 3023 3626
rect 3027 3622 3167 3626
rect 3171 3622 3183 3626
rect 3187 3622 3303 3626
rect 3307 3622 3359 3626
rect 3363 3622 3431 3626
rect 3435 3622 3551 3626
rect 3555 3622 3671 3626
rect 3675 3622 3791 3626
rect 3795 3622 3895 3626
rect 3899 3622 3991 3626
rect 3995 3622 4027 3626
rect 2061 3621 4027 3622
rect 4033 3621 4034 3627
rect 96 3589 97 3595
rect 103 3594 2055 3595
rect 103 3590 111 3594
rect 115 3590 239 3594
rect 243 3590 343 3594
rect 347 3590 399 3594
rect 403 3590 519 3594
rect 523 3590 551 3594
rect 555 3590 695 3594
rect 699 3590 703 3594
rect 707 3590 855 3594
rect 859 3590 863 3594
rect 867 3590 999 3594
rect 1003 3590 1031 3594
rect 1035 3590 1135 3594
rect 1139 3590 1191 3594
rect 1195 3590 1263 3594
rect 1267 3590 1343 3594
rect 1347 3590 1383 3594
rect 1387 3590 1495 3594
rect 1499 3590 1607 3594
rect 1611 3590 1655 3594
rect 1659 3590 1719 3594
rect 1723 3590 1831 3594
rect 1835 3590 1935 3594
rect 1939 3590 2031 3594
rect 2035 3590 2055 3594
rect 103 3589 2055 3590
rect 2061 3589 2062 3595
rect 2042 3537 2043 3543
rect 2049 3542 4015 3543
rect 2049 3538 2071 3542
rect 2075 3538 2111 3542
rect 2115 3538 2295 3542
rect 2299 3538 2447 3542
rect 2451 3538 2495 3542
rect 2499 3538 2591 3542
rect 2595 3538 2687 3542
rect 2691 3538 2727 3542
rect 2731 3538 2863 3542
rect 2867 3538 2991 3542
rect 2995 3538 3023 3542
rect 3027 3538 3119 3542
rect 3123 3538 3167 3542
rect 3171 3538 3239 3542
rect 3243 3538 3303 3542
rect 3307 3538 3351 3542
rect 3355 3538 3431 3542
rect 3435 3538 3463 3542
rect 3467 3538 3551 3542
rect 3555 3538 3575 3542
rect 3579 3538 3671 3542
rect 3675 3538 3687 3542
rect 3691 3538 3791 3542
rect 3795 3538 3895 3542
rect 3899 3538 3991 3542
rect 3995 3538 4015 3542
rect 2049 3537 4015 3538
rect 4021 3537 4022 3543
rect 84 3517 85 3523
rect 91 3522 2043 3523
rect 91 3518 111 3522
rect 115 3518 151 3522
rect 155 3518 239 3522
rect 243 3518 375 3522
rect 379 3518 399 3522
rect 403 3518 551 3522
rect 555 3518 615 3522
rect 619 3518 703 3522
rect 707 3518 847 3522
rect 851 3518 855 3522
rect 859 3518 999 3522
rect 1003 3518 1063 3522
rect 1067 3518 1135 3522
rect 1139 3518 1255 3522
rect 1259 3518 1263 3522
rect 1267 3518 1383 3522
rect 1387 3518 1439 3522
rect 1443 3518 1495 3522
rect 1499 3518 1607 3522
rect 1611 3518 1615 3522
rect 1619 3518 1719 3522
rect 1723 3518 1783 3522
rect 1787 3518 1831 3522
rect 1835 3518 1935 3522
rect 1939 3518 2031 3522
rect 2035 3518 2043 3522
rect 91 3517 2043 3518
rect 2049 3517 2050 3523
rect 2054 3465 2055 3471
rect 2061 3470 4027 3471
rect 2061 3466 2071 3470
rect 2075 3466 2343 3470
rect 2347 3466 2447 3470
rect 2451 3466 2591 3470
rect 2595 3466 2727 3470
rect 2731 3466 2855 3470
rect 2859 3466 2863 3470
rect 2867 3466 2991 3470
rect 2995 3466 3119 3470
rect 3123 3466 3239 3470
rect 3243 3466 3351 3470
rect 3355 3466 3375 3470
rect 3379 3466 3463 3470
rect 3467 3466 3575 3470
rect 3579 3466 3687 3470
rect 3691 3466 3791 3470
rect 3795 3466 3895 3470
rect 3899 3466 3991 3470
rect 3995 3466 4027 3470
rect 2061 3465 4027 3466
rect 4033 3465 4034 3471
rect 96 3421 97 3427
rect 103 3426 2055 3427
rect 103 3422 111 3426
rect 115 3422 151 3426
rect 155 3422 335 3426
rect 339 3422 375 3426
rect 379 3422 583 3426
rect 587 3422 615 3426
rect 619 3422 847 3426
rect 851 3422 863 3426
rect 867 3422 1063 3426
rect 1067 3422 1159 3426
rect 1163 3422 1255 3426
rect 1259 3422 1439 3426
rect 1443 3422 1463 3426
rect 1467 3422 1615 3426
rect 1619 3422 1783 3426
rect 1787 3422 1935 3426
rect 1939 3422 2031 3426
rect 2035 3422 2055 3426
rect 103 3421 2055 3422
rect 2061 3421 2062 3427
rect 2042 3389 2043 3395
rect 2049 3394 4015 3395
rect 2049 3390 2071 3394
rect 2075 3390 2183 3394
rect 2187 3390 2343 3394
rect 2347 3390 2583 3394
rect 2587 3390 2855 3394
rect 2859 3390 3007 3394
rect 3011 3390 3375 3394
rect 3379 3390 3447 3394
rect 3451 3390 3895 3394
rect 3899 3390 3991 3394
rect 3995 3390 4015 3394
rect 2049 3389 4015 3390
rect 4021 3389 4022 3395
rect 84 3341 85 3347
rect 91 3346 2043 3347
rect 91 3342 111 3346
rect 115 3342 151 3346
rect 155 3342 287 3346
rect 291 3342 335 3346
rect 339 3342 463 3346
rect 467 3342 583 3346
rect 587 3342 639 3346
rect 643 3342 815 3346
rect 819 3342 863 3346
rect 867 3342 991 3346
rect 995 3342 1159 3346
rect 1163 3342 1319 3346
rect 1323 3342 1463 3346
rect 1467 3342 1487 3346
rect 1491 3342 1655 3346
rect 1659 3342 2031 3346
rect 2035 3342 2043 3346
rect 91 3341 2043 3342
rect 2049 3341 2050 3347
rect 2054 3301 2055 3307
rect 2061 3306 4027 3307
rect 2061 3302 2071 3306
rect 2075 3302 2111 3306
rect 2115 3302 2183 3306
rect 2187 3302 2295 3306
rect 2299 3302 2503 3306
rect 2507 3302 2583 3306
rect 2587 3302 2703 3306
rect 2707 3302 2895 3306
rect 2899 3302 3007 3306
rect 3011 3302 3071 3306
rect 3075 3302 3231 3306
rect 3235 3302 3375 3306
rect 3379 3302 3447 3306
rect 3451 3302 3511 3306
rect 3515 3302 3647 3306
rect 3651 3302 3783 3306
rect 3787 3302 3895 3306
rect 3899 3302 3991 3306
rect 3995 3302 4027 3306
rect 2061 3301 4027 3302
rect 4033 3301 4034 3307
rect 96 3257 97 3263
rect 103 3262 2055 3263
rect 103 3258 111 3262
rect 115 3258 151 3262
rect 155 3258 287 3262
rect 291 3258 295 3262
rect 299 3258 463 3262
rect 467 3258 479 3262
rect 483 3258 639 3262
rect 643 3258 671 3262
rect 675 3258 815 3262
rect 819 3258 863 3262
rect 867 3258 991 3262
rect 995 3258 1055 3262
rect 1059 3258 1159 3262
rect 1163 3258 1247 3262
rect 1251 3258 1319 3262
rect 1323 3258 1431 3262
rect 1435 3258 1487 3262
rect 1491 3258 1615 3262
rect 1619 3258 1655 3262
rect 1659 3258 1807 3262
rect 1811 3258 2031 3262
rect 2035 3258 2055 3262
rect 103 3257 2055 3258
rect 2061 3257 2062 3263
rect 2042 3229 2043 3235
rect 2049 3234 4015 3235
rect 2049 3230 2071 3234
rect 2075 3230 2111 3234
rect 2115 3230 2239 3234
rect 2243 3230 2295 3234
rect 2299 3230 2399 3234
rect 2403 3230 2503 3234
rect 2507 3230 2559 3234
rect 2563 3230 2703 3234
rect 2707 3230 2719 3234
rect 2723 3230 2879 3234
rect 2883 3230 2895 3234
rect 2899 3230 3031 3234
rect 3035 3230 3071 3234
rect 3075 3230 3167 3234
rect 3171 3230 3231 3234
rect 3235 3230 3303 3234
rect 3307 3230 3375 3234
rect 3379 3230 3431 3234
rect 3435 3230 3511 3234
rect 3515 3230 3551 3234
rect 3555 3230 3647 3234
rect 3651 3230 3671 3234
rect 3675 3230 3783 3234
rect 3787 3230 3791 3234
rect 3795 3230 3895 3234
rect 3899 3230 3991 3234
rect 3995 3230 4015 3234
rect 2049 3229 4015 3230
rect 4021 3229 4022 3235
rect 84 3173 85 3179
rect 91 3178 2043 3179
rect 91 3174 111 3178
rect 115 3174 151 3178
rect 155 3174 287 3178
rect 291 3174 295 3178
rect 299 3174 423 3178
rect 427 3174 479 3178
rect 483 3174 567 3178
rect 571 3174 671 3178
rect 675 3174 727 3178
rect 731 3174 863 3178
rect 867 3174 903 3178
rect 907 3174 1055 3178
rect 1059 3174 1095 3178
rect 1099 3174 1247 3178
rect 1251 3174 1295 3178
rect 1299 3174 1431 3178
rect 1435 3174 1495 3178
rect 1499 3174 1615 3178
rect 1619 3174 1703 3178
rect 1707 3174 1807 3178
rect 1811 3174 1919 3178
rect 1923 3174 2031 3178
rect 2035 3174 2043 3178
rect 91 3173 2043 3174
rect 2049 3173 2050 3179
rect 2054 3141 2055 3147
rect 2061 3146 4027 3147
rect 2061 3142 2071 3146
rect 2075 3142 2111 3146
rect 2115 3142 2183 3146
rect 2187 3142 2239 3146
rect 2243 3142 2367 3146
rect 2371 3142 2399 3146
rect 2403 3142 2551 3146
rect 2555 3142 2559 3146
rect 2563 3142 2719 3146
rect 2723 3142 2735 3146
rect 2739 3142 2879 3146
rect 2883 3142 2911 3146
rect 2915 3142 3031 3146
rect 3035 3142 3087 3146
rect 3091 3142 3167 3146
rect 3171 3142 3263 3146
rect 3267 3142 3303 3146
rect 3307 3142 3431 3146
rect 3435 3142 3447 3146
rect 3451 3142 3551 3146
rect 3555 3142 3671 3146
rect 3675 3142 3791 3146
rect 3795 3142 3895 3146
rect 3899 3142 3991 3146
rect 3995 3142 4027 3146
rect 2061 3141 4027 3142
rect 4033 3141 4034 3147
rect 96 3085 97 3091
rect 103 3090 2055 3091
rect 103 3086 111 3090
rect 115 3086 287 3090
rect 291 3086 423 3090
rect 427 3086 567 3090
rect 571 3086 575 3090
rect 579 3086 679 3090
rect 683 3086 727 3090
rect 731 3086 799 3090
rect 803 3086 903 3090
rect 907 3086 935 3090
rect 939 3086 1079 3090
rect 1083 3086 1095 3090
rect 1099 3086 1231 3090
rect 1235 3086 1295 3090
rect 1299 3086 1391 3090
rect 1395 3086 1495 3090
rect 1499 3086 1559 3090
rect 1563 3086 1703 3090
rect 1707 3086 1727 3090
rect 1731 3086 1903 3090
rect 1907 3086 1919 3090
rect 1923 3086 2031 3090
rect 2035 3086 2055 3090
rect 103 3085 2055 3086
rect 2061 3085 2062 3091
rect 2042 3061 2043 3067
rect 2049 3066 4015 3067
rect 2049 3062 2071 3066
rect 2075 3062 2183 3066
rect 2187 3062 2351 3066
rect 2355 3062 2367 3066
rect 2371 3062 2455 3066
rect 2459 3062 2551 3066
rect 2555 3062 2567 3066
rect 2571 3062 2687 3066
rect 2691 3062 2735 3066
rect 2739 3062 2807 3066
rect 2811 3062 2911 3066
rect 2915 3062 2927 3066
rect 2931 3062 3047 3066
rect 3051 3062 3087 3066
rect 3091 3062 3167 3066
rect 3171 3062 3263 3066
rect 3267 3062 3295 3066
rect 3299 3062 3447 3066
rect 3451 3062 3991 3066
rect 3995 3062 4015 3066
rect 2049 3061 4015 3062
rect 4021 3061 4022 3067
rect 84 3001 85 3007
rect 91 3006 2043 3007
rect 91 3002 111 3006
rect 115 3002 551 3006
rect 555 3002 575 3006
rect 579 3002 655 3006
rect 659 3002 679 3006
rect 683 3002 759 3006
rect 763 3002 799 3006
rect 803 3002 871 3006
rect 875 3002 935 3006
rect 939 3002 991 3006
rect 995 3002 1079 3006
rect 1083 3002 1119 3006
rect 1123 3002 1231 3006
rect 1235 3002 1255 3006
rect 1259 3002 1391 3006
rect 1395 3002 1535 3006
rect 1539 3002 1559 3006
rect 1563 3002 1687 3006
rect 1691 3002 1727 3006
rect 1731 3002 1903 3006
rect 1907 3002 2031 3006
rect 2035 3002 2043 3006
rect 91 3001 2043 3002
rect 2049 3001 2050 3007
rect 2054 2989 2055 2995
rect 2061 2994 4027 2995
rect 2061 2990 2071 2994
rect 2075 2990 2351 2994
rect 2355 2990 2455 2994
rect 2459 2990 2495 2994
rect 2499 2990 2567 2994
rect 2571 2990 2599 2994
rect 2603 2990 2687 2994
rect 2691 2990 2703 2994
rect 2707 2990 2807 2994
rect 2811 2990 2911 2994
rect 2915 2990 2927 2994
rect 2931 2990 3015 2994
rect 3019 2990 3047 2994
rect 3051 2990 3119 2994
rect 3123 2990 3167 2994
rect 3171 2990 3223 2994
rect 3227 2990 3295 2994
rect 3299 2990 3991 2994
rect 3995 2990 4027 2994
rect 2061 2989 4027 2990
rect 4033 2989 4034 2995
rect 2042 2927 2043 2933
rect 2049 2927 2074 2933
rect 2068 2923 2074 2927
rect 96 2917 97 2923
rect 103 2922 2055 2923
rect 103 2918 111 2922
rect 115 2918 311 2922
rect 315 2918 431 2922
rect 435 2918 551 2922
rect 555 2918 559 2922
rect 563 2918 655 2922
rect 659 2918 695 2922
rect 699 2918 759 2922
rect 763 2918 831 2922
rect 835 2918 871 2922
rect 875 2918 975 2922
rect 979 2918 991 2922
rect 995 2918 1119 2922
rect 1123 2918 1255 2922
rect 1259 2918 1271 2922
rect 1275 2918 1391 2922
rect 1395 2918 1423 2922
rect 1427 2918 1535 2922
rect 1539 2918 1575 2922
rect 1579 2918 1687 2922
rect 1691 2918 2031 2922
rect 2035 2918 2055 2922
rect 103 2917 2055 2918
rect 2061 2917 2062 2923
rect 2068 2922 4015 2923
rect 2068 2918 2071 2922
rect 2075 2918 2415 2922
rect 2419 2918 2495 2922
rect 2499 2918 2519 2922
rect 2523 2918 2599 2922
rect 2603 2918 2623 2922
rect 2627 2918 2703 2922
rect 2707 2918 2727 2922
rect 2731 2918 2807 2922
rect 2811 2918 2831 2922
rect 2835 2918 2911 2922
rect 2915 2918 2935 2922
rect 2939 2918 3015 2922
rect 3019 2918 3039 2922
rect 3043 2918 3119 2922
rect 3123 2918 3143 2922
rect 3147 2918 3223 2922
rect 3227 2918 3247 2922
rect 3251 2918 3991 2922
rect 3995 2918 4015 2922
rect 2068 2917 4015 2918
rect 4021 2917 4022 2923
rect 2054 2841 2055 2847
rect 2061 2846 4027 2847
rect 2061 2842 2071 2846
rect 2075 2842 2407 2846
rect 2411 2842 2415 2846
rect 2419 2842 2511 2846
rect 2515 2842 2519 2846
rect 2523 2842 2615 2846
rect 2619 2842 2623 2846
rect 2627 2842 2719 2846
rect 2723 2842 2727 2846
rect 2731 2842 2823 2846
rect 2827 2842 2831 2846
rect 2835 2842 2927 2846
rect 2931 2842 2935 2846
rect 2939 2842 3031 2846
rect 3035 2842 3039 2846
rect 3043 2842 3135 2846
rect 3139 2842 3143 2846
rect 3147 2842 3239 2846
rect 3243 2842 3247 2846
rect 3251 2842 3991 2846
rect 3995 2842 4027 2846
rect 2061 2841 4027 2842
rect 4033 2841 4034 2847
rect 84 2829 85 2835
rect 91 2834 2043 2835
rect 91 2830 111 2834
rect 115 2830 151 2834
rect 155 2830 311 2834
rect 315 2830 431 2834
rect 435 2830 471 2834
rect 475 2830 559 2834
rect 563 2830 623 2834
rect 627 2830 695 2834
rect 699 2830 767 2834
rect 771 2830 831 2834
rect 835 2830 903 2834
rect 907 2830 975 2834
rect 979 2830 1031 2834
rect 1035 2830 1119 2834
rect 1123 2830 1159 2834
rect 1163 2830 1271 2834
rect 1275 2830 1287 2834
rect 1291 2830 1415 2834
rect 1419 2830 1423 2834
rect 1427 2830 1575 2834
rect 1579 2830 2031 2834
rect 2035 2830 2043 2834
rect 91 2829 2043 2830
rect 2049 2829 2050 2835
rect 2042 2761 2043 2767
rect 2049 2766 4015 2767
rect 2049 2762 2071 2766
rect 2075 2762 2303 2766
rect 2307 2762 2407 2766
rect 2411 2762 2415 2766
rect 2419 2762 2511 2766
rect 2515 2762 2535 2766
rect 2539 2762 2615 2766
rect 2619 2762 2655 2766
rect 2659 2762 2719 2766
rect 2723 2762 2775 2766
rect 2779 2762 2823 2766
rect 2827 2762 2895 2766
rect 2899 2762 2927 2766
rect 2931 2762 3015 2766
rect 3019 2762 3031 2766
rect 3035 2762 3135 2766
rect 3139 2762 3143 2766
rect 3147 2762 3239 2766
rect 3243 2762 3271 2766
rect 3275 2762 3399 2766
rect 3403 2762 3991 2766
rect 3995 2762 4015 2766
rect 2049 2761 4015 2762
rect 4021 2761 4022 2767
rect 96 2741 97 2747
rect 103 2746 2055 2747
rect 103 2742 111 2746
rect 115 2742 151 2746
rect 155 2742 303 2746
rect 307 2742 311 2746
rect 315 2742 471 2746
rect 475 2742 623 2746
rect 627 2742 767 2746
rect 771 2742 903 2746
rect 907 2742 1031 2746
rect 1035 2742 1039 2746
rect 1043 2742 1159 2746
rect 1163 2742 1167 2746
rect 1171 2742 1287 2746
rect 1291 2742 1295 2746
rect 1299 2742 1415 2746
rect 1419 2742 1423 2746
rect 1427 2742 2031 2746
rect 2035 2742 2055 2746
rect 103 2741 2055 2742
rect 2061 2741 2062 2747
rect 2054 2673 2055 2679
rect 2061 2678 4027 2679
rect 2061 2674 2071 2678
rect 2075 2674 2151 2678
rect 2155 2674 2303 2678
rect 2307 2674 2415 2678
rect 2419 2674 2463 2678
rect 2467 2674 2535 2678
rect 2539 2674 2623 2678
rect 2627 2674 2655 2678
rect 2659 2674 2775 2678
rect 2779 2674 2791 2678
rect 2795 2674 2895 2678
rect 2899 2674 2951 2678
rect 2955 2674 3015 2678
rect 3019 2674 3111 2678
rect 3115 2674 3143 2678
rect 3147 2674 3263 2678
rect 3267 2674 3271 2678
rect 3275 2674 3399 2678
rect 3403 2674 3415 2678
rect 3419 2674 3575 2678
rect 3579 2674 3991 2678
rect 3995 2674 4027 2678
rect 2061 2673 4027 2674
rect 4033 2673 4034 2679
rect 84 2657 85 2663
rect 91 2662 2043 2663
rect 91 2658 111 2662
rect 115 2658 151 2662
rect 155 2658 303 2662
rect 307 2658 319 2662
rect 323 2658 471 2662
rect 475 2658 511 2662
rect 515 2658 623 2662
rect 627 2658 703 2662
rect 707 2658 767 2662
rect 771 2658 887 2662
rect 891 2658 903 2662
rect 907 2658 1039 2662
rect 1043 2658 1063 2662
rect 1067 2658 1167 2662
rect 1171 2658 1231 2662
rect 1235 2658 1295 2662
rect 1299 2658 1391 2662
rect 1395 2658 1423 2662
rect 1427 2658 1551 2662
rect 1555 2658 1711 2662
rect 1715 2658 2031 2662
rect 2035 2658 2043 2662
rect 91 2657 2043 2658
rect 2049 2657 2050 2663
rect 2042 2593 2043 2599
rect 2049 2598 4015 2599
rect 2049 2594 2071 2598
rect 2075 2594 2111 2598
rect 2115 2594 2151 2598
rect 2155 2594 2303 2598
rect 2307 2594 2327 2598
rect 2331 2594 2463 2598
rect 2467 2594 2559 2598
rect 2563 2594 2623 2598
rect 2627 2594 2783 2598
rect 2787 2594 2791 2598
rect 2795 2594 2951 2598
rect 2955 2594 2999 2598
rect 3003 2594 3111 2598
rect 3115 2594 3199 2598
rect 3203 2594 3263 2598
rect 3267 2594 3383 2598
rect 3387 2594 3415 2598
rect 3419 2594 3559 2598
rect 3563 2594 3575 2598
rect 3579 2594 3735 2598
rect 3739 2594 3895 2598
rect 3899 2594 3991 2598
rect 3995 2594 4015 2598
rect 2049 2593 4015 2594
rect 4021 2593 4022 2599
rect 96 2569 97 2575
rect 103 2574 2055 2575
rect 103 2570 111 2574
rect 115 2570 151 2574
rect 155 2570 279 2574
rect 283 2570 319 2574
rect 323 2570 463 2574
rect 467 2570 511 2574
rect 515 2570 663 2574
rect 667 2570 703 2574
rect 707 2570 863 2574
rect 867 2570 887 2574
rect 891 2570 1063 2574
rect 1067 2570 1231 2574
rect 1235 2570 1255 2574
rect 1259 2570 1391 2574
rect 1395 2570 1431 2574
rect 1435 2570 1551 2574
rect 1555 2570 1607 2574
rect 1611 2570 1711 2574
rect 1715 2570 1783 2574
rect 1787 2570 1935 2574
rect 1939 2570 2031 2574
rect 2035 2570 2055 2574
rect 103 2569 2055 2570
rect 2061 2569 2062 2575
rect 2054 2521 2055 2527
rect 2061 2526 4027 2527
rect 2061 2522 2071 2526
rect 2075 2522 2111 2526
rect 2115 2522 2255 2526
rect 2259 2522 2327 2526
rect 2331 2522 2439 2526
rect 2443 2522 2559 2526
rect 2563 2522 2631 2526
rect 2635 2522 2783 2526
rect 2787 2522 2823 2526
rect 2827 2522 2999 2526
rect 3003 2522 3007 2526
rect 3011 2522 3175 2526
rect 3179 2522 3199 2526
rect 3203 2522 3335 2526
rect 3339 2522 3383 2526
rect 3387 2522 3487 2526
rect 3491 2522 3559 2526
rect 3563 2522 3631 2526
rect 3635 2522 3735 2526
rect 3739 2522 3775 2526
rect 3779 2522 3895 2526
rect 3899 2522 3991 2526
rect 3995 2522 4027 2526
rect 2061 2521 4027 2522
rect 4033 2521 4034 2527
rect 84 2481 85 2487
rect 91 2486 2043 2487
rect 91 2482 111 2486
rect 115 2482 279 2486
rect 283 2482 311 2486
rect 315 2482 463 2486
rect 467 2482 471 2486
rect 475 2482 647 2486
rect 651 2482 663 2486
rect 667 2482 831 2486
rect 835 2482 863 2486
rect 867 2482 1015 2486
rect 1019 2482 1063 2486
rect 1067 2482 1191 2486
rect 1195 2482 1255 2486
rect 1259 2482 1367 2486
rect 1371 2482 1431 2486
rect 1435 2482 1535 2486
rect 1539 2482 1607 2486
rect 1611 2482 1703 2486
rect 1707 2482 1783 2486
rect 1787 2482 1871 2486
rect 1875 2482 1935 2486
rect 1939 2482 2031 2486
rect 2035 2482 2043 2486
rect 91 2481 2043 2482
rect 2049 2481 2050 2487
rect 2042 2441 2043 2447
rect 2049 2446 4015 2447
rect 2049 2442 2071 2446
rect 2075 2442 2111 2446
rect 2115 2442 2255 2446
rect 2259 2442 2311 2446
rect 2315 2442 2439 2446
rect 2443 2442 2535 2446
rect 2539 2442 2631 2446
rect 2635 2442 2751 2446
rect 2755 2442 2823 2446
rect 2827 2442 2951 2446
rect 2955 2442 3007 2446
rect 3011 2442 3135 2446
rect 3139 2442 3175 2446
rect 3179 2442 3311 2446
rect 3315 2442 3335 2446
rect 3339 2442 3471 2446
rect 3475 2442 3487 2446
rect 3491 2442 3623 2446
rect 3627 2442 3631 2446
rect 3635 2442 3767 2446
rect 3771 2442 3775 2446
rect 3779 2442 3895 2446
rect 3899 2442 3991 2446
rect 3995 2442 4015 2446
rect 2049 2441 4015 2442
rect 4021 2441 4022 2447
rect 96 2397 97 2403
rect 103 2402 2055 2403
rect 103 2398 111 2402
rect 115 2398 207 2402
rect 211 2398 311 2402
rect 315 2398 351 2402
rect 355 2398 471 2402
rect 475 2398 503 2402
rect 507 2398 647 2402
rect 651 2398 655 2402
rect 659 2398 815 2402
rect 819 2398 831 2402
rect 835 2398 967 2402
rect 971 2398 1015 2402
rect 1019 2398 1119 2402
rect 1123 2398 1191 2402
rect 1195 2398 1263 2402
rect 1267 2398 1367 2402
rect 1371 2398 1415 2402
rect 1419 2398 1535 2402
rect 1539 2398 1567 2402
rect 1571 2398 1703 2402
rect 1707 2398 1871 2402
rect 1875 2398 2031 2402
rect 2035 2398 2055 2402
rect 103 2397 2055 2398
rect 2061 2397 2062 2403
rect 2054 2369 2055 2375
rect 2061 2374 4027 2375
rect 2061 2370 2071 2374
rect 2075 2370 2111 2374
rect 2115 2370 2311 2374
rect 2315 2370 2327 2374
rect 2331 2370 2535 2374
rect 2539 2370 2559 2374
rect 2563 2370 2751 2374
rect 2755 2370 2783 2374
rect 2787 2370 2951 2374
rect 2955 2370 2999 2374
rect 3003 2370 3135 2374
rect 3139 2370 3191 2374
rect 3195 2370 3311 2374
rect 3315 2370 3375 2374
rect 3379 2370 3471 2374
rect 3475 2370 3543 2374
rect 3547 2370 3623 2374
rect 3627 2370 3711 2374
rect 3715 2370 3767 2374
rect 3771 2370 3887 2374
rect 3891 2370 3895 2374
rect 3899 2370 3991 2374
rect 3995 2370 4027 2374
rect 2061 2369 4027 2370
rect 4033 2369 4034 2375
rect 84 2313 85 2319
rect 91 2318 2043 2319
rect 91 2314 111 2318
rect 115 2314 207 2318
rect 211 2314 255 2318
rect 259 2314 351 2318
rect 355 2314 359 2318
rect 363 2314 471 2318
rect 475 2314 503 2318
rect 507 2314 583 2318
rect 587 2314 655 2318
rect 659 2314 695 2318
rect 699 2314 807 2318
rect 811 2314 815 2318
rect 819 2314 919 2318
rect 923 2314 967 2318
rect 971 2314 1031 2318
rect 1035 2314 1119 2318
rect 1123 2314 1151 2318
rect 1155 2314 1263 2318
rect 1267 2314 1271 2318
rect 1275 2314 1415 2318
rect 1419 2314 1567 2318
rect 1571 2314 2031 2318
rect 2035 2314 2043 2318
rect 91 2313 2043 2314
rect 2049 2313 2050 2319
rect 2042 2297 2043 2303
rect 2049 2302 4015 2303
rect 2049 2298 2071 2302
rect 2075 2298 2111 2302
rect 2115 2298 2295 2302
rect 2299 2298 2327 2302
rect 2331 2298 2527 2302
rect 2531 2298 2559 2302
rect 2563 2298 2775 2302
rect 2779 2298 2783 2302
rect 2787 2298 2999 2302
rect 3003 2298 3039 2302
rect 3043 2298 3191 2302
rect 3195 2298 3319 2302
rect 3323 2298 3375 2302
rect 3379 2298 3543 2302
rect 3547 2298 3607 2302
rect 3611 2298 3711 2302
rect 3715 2298 3887 2302
rect 3891 2298 3895 2302
rect 3899 2298 3991 2302
rect 3995 2298 4015 2302
rect 2049 2297 4015 2298
rect 4021 2297 4022 2303
rect 96 2229 97 2235
rect 103 2234 2055 2235
rect 103 2230 111 2234
rect 115 2230 183 2234
rect 187 2230 255 2234
rect 259 2230 343 2234
rect 347 2230 359 2234
rect 363 2230 471 2234
rect 475 2230 495 2234
rect 499 2230 583 2234
rect 587 2230 647 2234
rect 651 2230 695 2234
rect 699 2230 791 2234
rect 795 2230 807 2234
rect 811 2230 919 2234
rect 923 2230 935 2234
rect 939 2230 1031 2234
rect 1035 2230 1071 2234
rect 1075 2230 1151 2234
rect 1155 2230 1199 2234
rect 1203 2230 1271 2234
rect 1275 2230 1335 2234
rect 1339 2230 1471 2234
rect 1475 2230 2031 2234
rect 2035 2230 2055 2234
rect 103 2229 2055 2230
rect 2061 2229 2062 2235
rect 2054 2217 2055 2223
rect 2061 2222 4027 2223
rect 2061 2218 2071 2222
rect 2075 2218 2111 2222
rect 2115 2218 2279 2222
rect 2283 2218 2295 2222
rect 2299 2218 2439 2222
rect 2443 2218 2527 2222
rect 2531 2218 2623 2222
rect 2627 2218 2775 2222
rect 2779 2218 2839 2222
rect 2843 2218 3039 2222
rect 3043 2218 3079 2222
rect 3083 2218 3319 2222
rect 3323 2218 3343 2222
rect 3347 2218 3607 2222
rect 3611 2218 3623 2222
rect 3627 2218 3895 2222
rect 3899 2218 3991 2222
rect 3995 2218 4027 2222
rect 2061 2217 4027 2218
rect 4033 2217 4034 2223
rect 2042 2150 4022 2151
rect 2042 2147 2071 2150
rect 84 2141 85 2147
rect 91 2146 2043 2147
rect 91 2142 111 2146
rect 115 2142 151 2146
rect 155 2142 183 2146
rect 187 2142 327 2146
rect 331 2142 343 2146
rect 347 2142 495 2146
rect 499 2142 535 2146
rect 539 2142 647 2146
rect 651 2142 735 2146
rect 739 2142 791 2146
rect 795 2142 927 2146
rect 931 2142 935 2146
rect 939 2142 1071 2146
rect 1075 2142 1111 2146
rect 1115 2142 1199 2146
rect 1203 2142 1279 2146
rect 1283 2142 1335 2146
rect 1339 2142 1447 2146
rect 1451 2142 1471 2146
rect 1475 2142 1615 2146
rect 1619 2142 1783 2146
rect 1787 2142 2031 2146
rect 2035 2142 2043 2146
rect 91 2141 2043 2142
rect 2049 2146 2071 2147
rect 2075 2146 2279 2150
rect 2283 2146 2391 2150
rect 2395 2146 2439 2150
rect 2443 2146 2495 2150
rect 2499 2146 2599 2150
rect 2603 2146 2623 2150
rect 2627 2146 2703 2150
rect 2707 2146 2807 2150
rect 2811 2146 2839 2150
rect 2843 2146 2911 2150
rect 2915 2146 3031 2150
rect 3035 2146 3079 2150
rect 3083 2146 3175 2150
rect 3179 2146 3343 2150
rect 3347 2146 3527 2150
rect 3531 2146 3623 2150
rect 3627 2146 3719 2150
rect 3723 2146 3895 2150
rect 3899 2146 3991 2150
rect 3995 2146 4022 2150
rect 2049 2145 4022 2146
rect 2049 2141 2050 2145
rect 2054 2069 2055 2075
rect 2061 2074 4027 2075
rect 2061 2070 2071 2074
rect 2075 2070 2391 2074
rect 2395 2070 2487 2074
rect 2491 2070 2495 2074
rect 2499 2070 2591 2074
rect 2595 2070 2599 2074
rect 2603 2070 2695 2074
rect 2699 2070 2703 2074
rect 2707 2070 2807 2074
rect 2811 2070 2911 2074
rect 2915 2070 2935 2074
rect 2939 2070 3031 2074
rect 3035 2070 3095 2074
rect 3099 2070 3175 2074
rect 3179 2070 3279 2074
rect 3283 2070 3343 2074
rect 3347 2070 3479 2074
rect 3483 2070 3527 2074
rect 3531 2070 3695 2074
rect 3699 2070 3719 2074
rect 3723 2070 3895 2074
rect 3899 2070 3991 2074
rect 3995 2070 4027 2074
rect 2061 2069 4027 2070
rect 4033 2069 4034 2075
rect 96 2057 97 2063
rect 103 2062 2055 2063
rect 103 2058 111 2062
rect 115 2058 151 2062
rect 155 2058 327 2062
rect 331 2058 383 2062
rect 387 2058 535 2062
rect 539 2058 631 2062
rect 635 2058 735 2062
rect 739 2058 863 2062
rect 867 2058 927 2062
rect 931 2058 1071 2062
rect 1075 2058 1111 2062
rect 1115 2058 1263 2062
rect 1267 2058 1279 2062
rect 1283 2058 1447 2062
rect 1451 2058 1615 2062
rect 1619 2058 1783 2062
rect 1787 2058 1935 2062
rect 1939 2058 2031 2062
rect 2035 2058 2055 2062
rect 103 2057 2055 2058
rect 2061 2057 2062 2063
rect 2042 1989 2043 1995
rect 2049 1994 4015 1995
rect 2049 1990 2071 1994
rect 2075 1990 2487 1994
rect 2491 1990 2527 1994
rect 2531 1990 2591 1994
rect 2595 1990 2695 1994
rect 2699 1990 2703 1994
rect 2707 1990 2807 1994
rect 2811 1990 2887 1994
rect 2891 1990 2935 1994
rect 2939 1990 3079 1994
rect 3083 1990 3095 1994
rect 3099 1990 3279 1994
rect 3283 1990 3479 1994
rect 3483 1990 3487 1994
rect 3491 1990 3695 1994
rect 3699 1990 3703 1994
rect 3707 1990 3895 1994
rect 3899 1990 3991 1994
rect 3995 1990 4015 1994
rect 2049 1989 4015 1990
rect 4021 1989 4022 1995
rect 84 1973 85 1979
rect 91 1978 2043 1979
rect 91 1974 111 1978
rect 115 1974 151 1978
rect 155 1974 327 1978
rect 331 1974 383 1978
rect 387 1974 535 1978
rect 539 1974 631 1978
rect 635 1974 735 1978
rect 739 1974 863 1978
rect 867 1974 935 1978
rect 939 1974 1071 1978
rect 1075 1974 1127 1978
rect 1131 1974 1263 1978
rect 1267 1974 1303 1978
rect 1307 1974 1447 1978
rect 1451 1974 1471 1978
rect 1475 1974 1615 1978
rect 1619 1974 1631 1978
rect 1635 1974 1783 1978
rect 1787 1974 1791 1978
rect 1795 1974 1935 1978
rect 1939 1974 2031 1978
rect 2035 1974 2043 1978
rect 91 1973 2043 1974
rect 2049 1973 2050 1979
rect 2054 1913 2055 1919
rect 2061 1918 4027 1919
rect 2061 1914 2071 1918
rect 2075 1914 2111 1918
rect 2115 1914 2303 1918
rect 2307 1914 2519 1918
rect 2523 1914 2527 1918
rect 2531 1914 2703 1918
rect 2707 1914 2735 1918
rect 2739 1914 2887 1918
rect 2891 1914 2959 1918
rect 2963 1914 3079 1918
rect 3083 1914 3191 1918
rect 3195 1914 3279 1918
rect 3283 1914 3431 1918
rect 3435 1914 3487 1918
rect 3491 1914 3671 1918
rect 3675 1914 3703 1918
rect 3707 1914 3895 1918
rect 3899 1914 3991 1918
rect 3995 1914 4027 1918
rect 2061 1913 4027 1914
rect 4033 1913 4034 1919
rect 96 1897 97 1903
rect 103 1902 2055 1903
rect 103 1898 111 1902
rect 115 1898 151 1902
rect 155 1898 303 1902
rect 307 1898 327 1902
rect 331 1898 463 1902
rect 467 1898 535 1902
rect 539 1898 615 1902
rect 619 1898 735 1902
rect 739 1898 767 1902
rect 771 1898 927 1902
rect 931 1898 935 1902
rect 939 1898 1103 1902
rect 1107 1898 1127 1902
rect 1131 1898 1295 1902
rect 1299 1898 1303 1902
rect 1307 1898 1471 1902
rect 1475 1898 1511 1902
rect 1515 1898 1631 1902
rect 1635 1898 1735 1902
rect 1739 1898 1791 1902
rect 1795 1898 1935 1902
rect 1939 1898 2031 1902
rect 2035 1898 2055 1902
rect 103 1897 2055 1898
rect 2061 1897 2062 1903
rect 2042 1841 2043 1847
rect 2049 1846 4015 1847
rect 2049 1842 2071 1846
rect 2075 1842 2111 1846
rect 2115 1842 2231 1846
rect 2235 1842 2303 1846
rect 2307 1842 2399 1846
rect 2403 1842 2519 1846
rect 2523 1842 2599 1846
rect 2603 1842 2735 1846
rect 2739 1842 2831 1846
rect 2835 1842 2959 1846
rect 2963 1842 3079 1846
rect 3083 1842 3191 1846
rect 3195 1842 3351 1846
rect 3355 1842 3431 1846
rect 3435 1842 3631 1846
rect 3635 1842 3671 1846
rect 3675 1842 3895 1846
rect 3899 1842 3991 1846
rect 3995 1842 4015 1846
rect 2049 1841 4015 1842
rect 4021 1841 4022 1847
rect 84 1813 85 1819
rect 91 1818 2043 1819
rect 91 1814 111 1818
rect 115 1814 151 1818
rect 155 1814 303 1818
rect 307 1814 343 1818
rect 347 1814 463 1818
rect 467 1814 543 1818
rect 547 1814 615 1818
rect 619 1814 735 1818
rect 739 1814 767 1818
rect 771 1814 919 1818
rect 923 1814 927 1818
rect 931 1814 1095 1818
rect 1099 1814 1103 1818
rect 1107 1814 1271 1818
rect 1275 1814 1295 1818
rect 1299 1814 1447 1818
rect 1451 1814 1511 1818
rect 1515 1814 1623 1818
rect 1627 1814 1735 1818
rect 1739 1814 1807 1818
rect 1811 1814 1935 1818
rect 1939 1814 2031 1818
rect 2035 1814 2043 1818
rect 91 1813 2043 1814
rect 2049 1813 2050 1819
rect 2054 1765 2055 1771
rect 2061 1770 4027 1771
rect 2061 1766 2071 1770
rect 2075 1766 2111 1770
rect 2115 1766 2231 1770
rect 2235 1766 2239 1770
rect 2243 1766 2399 1770
rect 2403 1766 2575 1770
rect 2579 1766 2599 1770
rect 2603 1766 2751 1770
rect 2755 1766 2831 1770
rect 2835 1766 2935 1770
rect 2939 1766 3079 1770
rect 3083 1766 3127 1770
rect 3131 1766 3319 1770
rect 3323 1766 3351 1770
rect 3355 1766 3511 1770
rect 3515 1766 3631 1770
rect 3635 1766 3711 1770
rect 3715 1766 3895 1770
rect 3899 1766 3991 1770
rect 3995 1766 4027 1770
rect 2061 1765 4027 1766
rect 4033 1765 4034 1771
rect 96 1737 97 1743
rect 103 1742 2055 1743
rect 103 1738 111 1742
rect 115 1738 151 1742
rect 155 1738 319 1742
rect 323 1738 343 1742
rect 347 1738 527 1742
rect 531 1738 543 1742
rect 547 1738 735 1742
rect 739 1738 743 1742
rect 747 1738 919 1742
rect 923 1738 959 1742
rect 963 1738 1095 1742
rect 1099 1738 1167 1742
rect 1171 1738 1271 1742
rect 1275 1738 1367 1742
rect 1371 1738 1447 1742
rect 1451 1738 1559 1742
rect 1563 1738 1623 1742
rect 1627 1738 1759 1742
rect 1763 1738 1807 1742
rect 1811 1738 1935 1742
rect 1939 1738 2031 1742
rect 2035 1738 2055 1742
rect 103 1737 2055 1738
rect 2061 1737 2062 1743
rect 2042 1685 2043 1691
rect 2049 1690 4015 1691
rect 2049 1686 2071 1690
rect 2075 1686 2111 1690
rect 2115 1686 2239 1690
rect 2243 1686 2311 1690
rect 2315 1686 2399 1690
rect 2403 1686 2527 1690
rect 2531 1686 2575 1690
rect 2579 1686 2743 1690
rect 2747 1686 2751 1690
rect 2755 1686 2935 1690
rect 2939 1686 2951 1690
rect 2955 1686 3127 1690
rect 3131 1686 3151 1690
rect 3155 1686 3319 1690
rect 3323 1686 3343 1690
rect 3347 1686 3511 1690
rect 3515 1686 3527 1690
rect 3531 1686 3711 1690
rect 3715 1686 3719 1690
rect 3723 1686 3895 1690
rect 3899 1686 3991 1690
rect 3995 1686 4015 1690
rect 2049 1685 4015 1686
rect 4021 1685 4022 1691
rect 84 1665 85 1671
rect 91 1670 2043 1671
rect 91 1666 111 1670
rect 115 1666 151 1670
rect 155 1666 319 1670
rect 323 1666 503 1670
rect 507 1666 527 1670
rect 531 1666 695 1670
rect 699 1666 743 1670
rect 747 1666 887 1670
rect 891 1666 959 1670
rect 963 1666 1079 1670
rect 1083 1666 1167 1670
rect 1171 1666 1263 1670
rect 1267 1666 1367 1670
rect 1371 1666 1439 1670
rect 1443 1666 1559 1670
rect 1563 1666 1615 1670
rect 1619 1666 1759 1670
rect 1763 1666 1791 1670
rect 1795 1666 1935 1670
rect 1939 1666 2031 1670
rect 2035 1666 2043 1670
rect 91 1665 2043 1666
rect 2049 1665 2050 1671
rect 2054 1601 2055 1607
rect 2061 1606 4027 1607
rect 2061 1602 2071 1606
rect 2075 1602 2111 1606
rect 2115 1602 2311 1606
rect 2315 1602 2479 1606
rect 2483 1602 2527 1606
rect 2531 1602 2583 1606
rect 2587 1602 2695 1606
rect 2699 1602 2743 1606
rect 2747 1602 2815 1606
rect 2819 1602 2943 1606
rect 2947 1602 2951 1606
rect 2955 1602 3079 1606
rect 3083 1602 3151 1606
rect 3155 1602 3223 1606
rect 3227 1602 3343 1606
rect 3347 1602 3383 1606
rect 3387 1602 3527 1606
rect 3531 1602 3551 1606
rect 3555 1602 3719 1606
rect 3723 1602 3727 1606
rect 3731 1602 3895 1606
rect 3899 1602 3991 1606
rect 3995 1602 4027 1606
rect 2061 1601 4027 1602
rect 4033 1601 4034 1607
rect 96 1585 97 1591
rect 103 1590 2055 1591
rect 103 1586 111 1590
rect 115 1586 151 1590
rect 155 1586 319 1590
rect 323 1586 455 1590
rect 459 1586 503 1590
rect 507 1586 599 1590
rect 603 1586 695 1590
rect 699 1586 743 1590
rect 747 1586 887 1590
rect 891 1586 1031 1590
rect 1035 1586 1079 1590
rect 1083 1586 1175 1590
rect 1179 1586 1263 1590
rect 1267 1586 1319 1590
rect 1323 1586 1439 1590
rect 1443 1586 1471 1590
rect 1475 1586 1615 1590
rect 1619 1586 1623 1590
rect 1627 1586 1791 1590
rect 1795 1586 2031 1590
rect 2035 1586 2055 1590
rect 103 1585 2055 1586
rect 2061 1585 2062 1591
rect 2042 1517 2043 1523
rect 2049 1522 4015 1523
rect 2049 1518 2071 1522
rect 2075 1518 2479 1522
rect 2483 1518 2487 1522
rect 2491 1518 2583 1522
rect 2587 1518 2591 1522
rect 2595 1518 2695 1522
rect 2699 1518 2807 1522
rect 2811 1518 2815 1522
rect 2819 1518 2935 1522
rect 2939 1518 2943 1522
rect 2947 1518 3071 1522
rect 3075 1518 3079 1522
rect 3083 1518 3223 1522
rect 3227 1518 3383 1522
rect 3387 1518 3551 1522
rect 3555 1518 3719 1522
rect 3723 1518 3727 1522
rect 3731 1518 3895 1522
rect 3899 1518 3991 1522
rect 3995 1518 4015 1522
rect 2049 1517 4015 1518
rect 4021 1517 4022 1523
rect 84 1505 85 1511
rect 91 1510 2043 1511
rect 91 1506 111 1510
rect 115 1506 319 1510
rect 323 1506 359 1510
rect 363 1506 455 1510
rect 459 1506 487 1510
rect 491 1506 599 1510
rect 603 1506 623 1510
rect 627 1506 743 1510
rect 747 1506 775 1510
rect 779 1506 887 1510
rect 891 1506 927 1510
rect 931 1506 1031 1510
rect 1035 1506 1087 1510
rect 1091 1506 1175 1510
rect 1179 1506 1255 1510
rect 1259 1506 1319 1510
rect 1323 1506 1423 1510
rect 1427 1506 1471 1510
rect 1475 1506 1591 1510
rect 1595 1506 1623 1510
rect 1627 1506 1767 1510
rect 1771 1506 2031 1510
rect 2035 1506 2043 1510
rect 91 1505 2043 1506
rect 2049 1505 2050 1511
rect 2054 1441 2055 1447
rect 2061 1446 4027 1447
rect 2061 1442 2071 1446
rect 2075 1442 2239 1446
rect 2243 1442 2351 1446
rect 2355 1442 2471 1446
rect 2475 1442 2487 1446
rect 2491 1442 2591 1446
rect 2595 1442 2695 1446
rect 2699 1442 2727 1446
rect 2731 1442 2807 1446
rect 2811 1442 2879 1446
rect 2883 1442 2935 1446
rect 2939 1442 3055 1446
rect 3059 1442 3071 1446
rect 3075 1442 3223 1446
rect 3227 1442 3247 1446
rect 3251 1442 3383 1446
rect 3387 1442 3455 1446
rect 3459 1442 3551 1446
rect 3555 1442 3671 1446
rect 3675 1442 3719 1446
rect 3723 1442 3887 1446
rect 3891 1442 3895 1446
rect 3899 1442 3991 1446
rect 3995 1442 4027 1446
rect 2061 1441 4027 1442
rect 4033 1441 4034 1447
rect 96 1425 97 1431
rect 103 1430 2055 1431
rect 103 1426 111 1430
rect 115 1426 151 1430
rect 155 1426 271 1430
rect 275 1426 359 1430
rect 363 1426 431 1430
rect 435 1426 487 1430
rect 491 1426 615 1430
rect 619 1426 623 1430
rect 627 1426 775 1430
rect 779 1426 807 1430
rect 811 1426 927 1430
rect 931 1426 1007 1430
rect 1011 1426 1087 1430
rect 1091 1426 1215 1430
rect 1219 1426 1255 1430
rect 1259 1426 1423 1430
rect 1427 1426 1591 1430
rect 1595 1426 1631 1430
rect 1635 1426 1767 1430
rect 1771 1426 1847 1430
rect 1851 1426 2031 1430
rect 2035 1426 2055 1430
rect 103 1425 2055 1426
rect 2061 1425 2062 1431
rect 2042 1361 2043 1367
rect 2049 1366 4015 1367
rect 2049 1362 2071 1366
rect 2075 1362 2239 1366
rect 2243 1362 2351 1366
rect 2355 1362 2391 1366
rect 2395 1362 2471 1366
rect 2475 1362 2527 1366
rect 2531 1362 2591 1366
rect 2595 1362 2679 1366
rect 2683 1362 2727 1366
rect 2731 1362 2839 1366
rect 2843 1362 2879 1366
rect 2883 1362 2999 1366
rect 3003 1362 3055 1366
rect 3059 1362 3167 1366
rect 3171 1362 3247 1366
rect 3251 1362 3343 1366
rect 3347 1362 3455 1366
rect 3459 1362 3519 1366
rect 3523 1362 3671 1366
rect 3675 1362 3695 1366
rect 3699 1362 3879 1366
rect 3883 1362 3887 1366
rect 3891 1362 3991 1366
rect 3995 1362 4015 1366
rect 2049 1361 4015 1362
rect 4021 1361 4022 1367
rect 84 1341 85 1347
rect 91 1346 2043 1347
rect 91 1342 111 1346
rect 115 1342 151 1346
rect 155 1342 271 1346
rect 275 1342 287 1346
rect 291 1342 431 1346
rect 435 1342 463 1346
rect 467 1342 615 1346
rect 619 1342 663 1346
rect 667 1342 807 1346
rect 811 1342 863 1346
rect 867 1342 1007 1346
rect 1011 1342 1063 1346
rect 1067 1342 1215 1346
rect 1219 1342 1255 1346
rect 1259 1342 1423 1346
rect 1427 1342 1431 1346
rect 1435 1342 1607 1346
rect 1611 1342 1631 1346
rect 1635 1342 1783 1346
rect 1787 1342 1847 1346
rect 1851 1342 1935 1346
rect 1939 1342 2031 1346
rect 2035 1342 2043 1346
rect 91 1341 2043 1342
rect 2049 1341 2050 1347
rect 2054 1281 2055 1287
rect 2061 1286 4027 1287
rect 2061 1282 2071 1286
rect 2075 1282 2111 1286
rect 2115 1282 2343 1286
rect 2347 1282 2391 1286
rect 2395 1282 2527 1286
rect 2531 1282 2583 1286
rect 2587 1282 2679 1286
rect 2683 1282 2799 1286
rect 2803 1282 2839 1286
rect 2843 1282 2999 1286
rect 3003 1282 3167 1286
rect 3171 1282 3183 1286
rect 3187 1282 3343 1286
rect 3347 1282 3495 1286
rect 3499 1282 3519 1286
rect 3523 1282 3639 1286
rect 3643 1282 3695 1286
rect 3699 1282 3775 1286
rect 3779 1282 3879 1286
rect 3883 1282 3895 1286
rect 3899 1282 3991 1286
rect 3995 1282 4027 1286
rect 2061 1281 4027 1282
rect 4033 1281 4034 1287
rect 96 1269 97 1275
rect 103 1274 2055 1275
rect 103 1270 111 1274
rect 115 1270 151 1274
rect 155 1270 207 1274
rect 211 1270 287 1274
rect 291 1270 327 1274
rect 331 1270 455 1274
rect 459 1270 463 1274
rect 467 1270 583 1274
rect 587 1270 663 1274
rect 667 1270 719 1274
rect 723 1270 863 1274
rect 867 1270 879 1274
rect 883 1270 1055 1274
rect 1059 1270 1063 1274
rect 1067 1270 1255 1274
rect 1259 1270 1263 1274
rect 1267 1270 1431 1274
rect 1435 1270 1487 1274
rect 1491 1270 1607 1274
rect 1611 1270 1719 1274
rect 1723 1270 1783 1274
rect 1787 1270 1935 1274
rect 1939 1270 2031 1274
rect 2035 1270 2055 1274
rect 103 1269 2055 1270
rect 2061 1269 2062 1275
rect 2042 1205 2043 1211
rect 2049 1210 4015 1211
rect 2049 1206 2071 1210
rect 2075 1206 2111 1210
rect 2115 1206 2279 1210
rect 2283 1206 2343 1210
rect 2347 1206 2471 1210
rect 2475 1206 2583 1210
rect 2587 1206 2655 1210
rect 2659 1206 2799 1210
rect 2803 1206 2831 1210
rect 2835 1206 2999 1210
rect 3003 1206 3159 1210
rect 3163 1206 3183 1210
rect 3187 1206 3327 1210
rect 3331 1206 3343 1210
rect 3347 1206 3495 1210
rect 3499 1206 3639 1210
rect 3643 1206 3775 1210
rect 3779 1206 3895 1210
rect 3899 1206 3991 1210
rect 3995 1206 4015 1210
rect 2049 1205 4015 1206
rect 4021 1205 4022 1211
rect 84 1189 85 1195
rect 91 1194 2043 1195
rect 91 1190 111 1194
rect 115 1190 207 1194
rect 211 1190 327 1194
rect 331 1190 455 1194
rect 459 1190 471 1194
rect 475 1190 583 1194
rect 587 1190 703 1194
rect 707 1190 719 1194
rect 723 1190 823 1194
rect 827 1190 879 1194
rect 883 1190 943 1194
rect 947 1190 1055 1194
rect 1059 1190 1063 1194
rect 1067 1190 1183 1194
rect 1187 1190 1263 1194
rect 1267 1190 1303 1194
rect 1307 1190 1423 1194
rect 1427 1190 1487 1194
rect 1491 1190 1543 1194
rect 1547 1190 1719 1194
rect 1723 1190 1935 1194
rect 1939 1190 2031 1194
rect 2035 1190 2043 1194
rect 91 1189 2043 1190
rect 2049 1189 2050 1195
rect 2054 1129 2055 1135
rect 2061 1134 4027 1135
rect 2061 1130 2071 1134
rect 2075 1130 2111 1134
rect 2115 1130 2279 1134
rect 2283 1130 2295 1134
rect 2299 1130 2471 1134
rect 2475 1130 2503 1134
rect 2507 1130 2655 1134
rect 2659 1130 2703 1134
rect 2707 1130 2831 1134
rect 2835 1130 2895 1134
rect 2899 1130 2999 1134
rect 3003 1130 3079 1134
rect 3083 1130 3159 1134
rect 3163 1130 3255 1134
rect 3259 1130 3327 1134
rect 3331 1130 3431 1134
rect 3435 1130 3495 1134
rect 3499 1130 3615 1134
rect 3619 1130 3991 1134
rect 3995 1130 4027 1134
rect 2061 1129 4027 1130
rect 4033 1129 4034 1135
rect 96 1109 97 1115
rect 103 1114 2055 1115
rect 103 1110 111 1114
rect 115 1110 471 1114
rect 475 1110 583 1114
rect 587 1110 623 1114
rect 627 1110 703 1114
rect 707 1110 735 1114
rect 739 1110 823 1114
rect 827 1110 855 1114
rect 859 1110 943 1114
rect 947 1110 975 1114
rect 979 1110 1063 1114
rect 1067 1110 1095 1114
rect 1099 1110 1183 1114
rect 1187 1110 1215 1114
rect 1219 1110 1303 1114
rect 1307 1110 1335 1114
rect 1339 1110 1423 1114
rect 1427 1110 1455 1114
rect 1459 1110 1543 1114
rect 1547 1110 1575 1114
rect 1579 1110 1703 1114
rect 1707 1110 2031 1114
rect 2035 1110 2055 1114
rect 103 1109 2055 1110
rect 2061 1109 2062 1115
rect 2042 1049 2043 1055
rect 2049 1054 4015 1055
rect 2049 1050 2071 1054
rect 2075 1050 2111 1054
rect 2115 1050 2167 1054
rect 2171 1050 2287 1054
rect 2291 1050 2295 1054
rect 2299 1050 2423 1054
rect 2427 1050 2503 1054
rect 2507 1050 2575 1054
rect 2579 1050 2703 1054
rect 2707 1050 2743 1054
rect 2747 1050 2895 1054
rect 2899 1050 2919 1054
rect 2923 1050 3079 1054
rect 3083 1050 3095 1054
rect 3099 1050 3255 1054
rect 3259 1050 3279 1054
rect 3283 1050 3431 1054
rect 3435 1050 3463 1054
rect 3467 1050 3615 1054
rect 3619 1050 3655 1054
rect 3659 1050 3991 1054
rect 3995 1050 4015 1054
rect 2049 1049 4015 1050
rect 4021 1049 4022 1055
rect 84 1029 85 1035
rect 91 1034 2043 1035
rect 91 1030 111 1034
rect 115 1030 623 1034
rect 627 1030 727 1034
rect 731 1030 735 1034
rect 739 1030 847 1034
rect 851 1030 855 1034
rect 859 1030 967 1034
rect 971 1030 975 1034
rect 979 1030 1095 1034
rect 1099 1030 1215 1034
rect 1219 1030 1223 1034
rect 1227 1030 1335 1034
rect 1339 1030 1351 1034
rect 1355 1030 1455 1034
rect 1459 1030 1479 1034
rect 1483 1030 1575 1034
rect 1579 1030 1607 1034
rect 1611 1030 1703 1034
rect 1707 1030 1735 1034
rect 1739 1030 1863 1034
rect 1867 1030 2031 1034
rect 2035 1030 2043 1034
rect 91 1029 2043 1030
rect 2049 1029 2050 1035
rect 2054 969 2055 975
rect 2061 974 4027 975
rect 2061 970 2071 974
rect 2075 970 2167 974
rect 2171 970 2287 974
rect 2291 970 2423 974
rect 2427 970 2527 974
rect 2531 970 2575 974
rect 2579 970 2647 974
rect 2651 970 2743 974
rect 2747 970 2775 974
rect 2779 970 2919 974
rect 2923 970 3071 974
rect 3075 970 3095 974
rect 3099 970 3231 974
rect 3235 970 3279 974
rect 3283 970 3399 974
rect 3403 970 3463 974
rect 3467 970 3567 974
rect 3571 970 3655 974
rect 3659 970 3735 974
rect 3739 970 3991 974
rect 3995 970 4027 974
rect 2061 969 4027 970
rect 4033 969 4034 975
rect 96 949 97 955
rect 103 954 2055 955
rect 103 950 111 954
rect 115 950 591 954
rect 595 950 727 954
rect 731 950 735 954
rect 739 950 847 954
rect 851 950 887 954
rect 891 950 967 954
rect 971 950 1039 954
rect 1043 950 1095 954
rect 1099 950 1199 954
rect 1203 950 1223 954
rect 1227 950 1351 954
rect 1355 950 1479 954
rect 1483 950 1503 954
rect 1507 950 1607 954
rect 1611 950 1655 954
rect 1659 950 1735 954
rect 1739 950 1807 954
rect 1811 950 1863 954
rect 1867 950 1935 954
rect 1939 950 2031 954
rect 2035 950 2055 954
rect 103 949 2055 950
rect 2061 949 2062 955
rect 2042 885 2043 891
rect 2049 890 4015 891
rect 2049 886 2071 890
rect 2075 886 2455 890
rect 2459 886 2527 890
rect 2531 886 2575 890
rect 2579 886 2647 890
rect 2651 886 2711 890
rect 2715 886 2775 890
rect 2779 886 2863 890
rect 2867 886 2919 890
rect 2923 886 3015 890
rect 3019 886 3071 890
rect 3075 886 3167 890
rect 3171 886 3231 890
rect 3235 886 3319 890
rect 3323 886 3399 890
rect 3403 886 3471 890
rect 3475 886 3567 890
rect 3571 886 3615 890
rect 3619 886 3735 890
rect 3739 886 3767 890
rect 3771 886 3895 890
rect 3899 886 3991 890
rect 3995 886 4015 890
rect 2049 885 4015 886
rect 4021 885 4022 891
rect 84 869 85 875
rect 91 874 2043 875
rect 91 870 111 874
rect 115 870 439 874
rect 443 870 583 874
rect 587 870 591 874
rect 595 870 735 874
rect 739 870 887 874
rect 891 870 1039 874
rect 1043 870 1047 874
rect 1051 870 1199 874
rect 1203 870 1351 874
rect 1355 870 1495 874
rect 1499 870 1503 874
rect 1507 870 1647 874
rect 1651 870 1655 874
rect 1659 870 1799 874
rect 1803 870 1807 874
rect 1811 870 1935 874
rect 1939 870 2031 874
rect 2035 870 2043 874
rect 91 869 2043 870
rect 2049 869 2050 875
rect 2054 813 2055 819
rect 2061 818 4027 819
rect 2061 814 2071 818
rect 2075 814 2215 818
rect 2219 814 2343 818
rect 2347 814 2455 818
rect 2459 814 2479 818
rect 2483 814 2575 818
rect 2579 814 2623 818
rect 2627 814 2711 818
rect 2715 814 2783 818
rect 2787 814 2863 818
rect 2867 814 2959 818
rect 2963 814 3015 818
rect 3019 814 3167 818
rect 3171 814 3319 818
rect 3323 814 3391 818
rect 3395 814 3471 818
rect 3475 814 3615 818
rect 3619 814 3623 818
rect 3627 814 3767 818
rect 3771 814 3863 818
rect 3867 814 3895 818
rect 3899 814 3991 818
rect 3995 814 4027 818
rect 2061 813 4027 814
rect 4033 813 4034 819
rect 96 797 97 803
rect 103 802 2055 803
rect 103 798 111 802
rect 115 798 279 802
rect 283 798 431 802
rect 435 798 439 802
rect 443 798 583 802
rect 587 798 591 802
rect 595 798 735 802
rect 739 798 751 802
rect 755 798 887 802
rect 891 798 919 802
rect 923 798 1047 802
rect 1051 798 1087 802
rect 1091 798 1199 802
rect 1203 798 1255 802
rect 1259 798 1351 802
rect 1355 798 1423 802
rect 1427 798 1495 802
rect 1499 798 1591 802
rect 1595 798 1647 802
rect 1651 798 1799 802
rect 1803 798 2031 802
rect 2035 798 2055 802
rect 103 797 2055 798
rect 2061 797 2062 803
rect 2042 733 2043 739
rect 2049 738 4015 739
rect 2049 734 2071 738
rect 2075 734 2111 738
rect 2115 734 2215 738
rect 2219 734 2247 738
rect 2251 734 2343 738
rect 2347 734 2423 738
rect 2427 734 2479 738
rect 2483 734 2599 738
rect 2603 734 2623 738
rect 2627 734 2783 738
rect 2787 734 2959 738
rect 2963 734 2967 738
rect 2971 734 3151 738
rect 3155 734 3167 738
rect 3171 734 3335 738
rect 3339 734 3391 738
rect 3395 734 3519 738
rect 3523 734 3623 738
rect 3627 734 3703 738
rect 3707 734 3863 738
rect 3867 734 3895 738
rect 3899 734 3991 738
rect 3995 734 4015 738
rect 2049 733 4015 734
rect 4021 733 4022 739
rect 84 721 85 727
rect 91 726 2043 727
rect 91 722 111 726
rect 115 722 151 726
rect 155 722 271 726
rect 275 722 279 726
rect 283 722 423 726
rect 427 722 431 726
rect 435 722 575 726
rect 579 722 591 726
rect 595 722 735 726
rect 739 722 751 726
rect 755 722 887 726
rect 891 722 919 726
rect 923 722 1039 726
rect 1043 722 1087 726
rect 1091 722 1191 726
rect 1195 722 1255 726
rect 1259 722 1343 726
rect 1347 722 1423 726
rect 1427 722 1495 726
rect 1499 722 1591 726
rect 1595 722 2031 726
rect 2035 722 2043 726
rect 91 721 2043 722
rect 2049 721 2050 727
rect 2054 657 2055 663
rect 2061 662 4027 663
rect 2061 658 2071 662
rect 2075 658 2111 662
rect 2115 658 2247 662
rect 2251 658 2375 662
rect 2379 658 2423 662
rect 2427 658 2599 662
rect 2603 658 2655 662
rect 2659 658 2783 662
rect 2787 658 2919 662
rect 2923 658 2967 662
rect 2971 658 3151 662
rect 3155 658 3175 662
rect 3179 658 3335 662
rect 3339 658 3423 662
rect 3427 658 3519 662
rect 3523 658 3671 662
rect 3675 658 3703 662
rect 3707 658 3895 662
rect 3899 658 3991 662
rect 3995 658 4027 662
rect 2061 657 4027 658
rect 4033 657 4034 663
rect 96 641 97 647
rect 103 646 2055 647
rect 103 642 111 646
rect 115 642 151 646
rect 155 642 255 646
rect 259 642 271 646
rect 275 642 391 646
rect 395 642 423 646
rect 427 642 527 646
rect 531 642 575 646
rect 579 642 663 646
rect 667 642 735 646
rect 739 642 807 646
rect 811 642 887 646
rect 891 642 959 646
rect 963 642 1039 646
rect 1043 642 1119 646
rect 1123 642 1191 646
rect 1195 642 1287 646
rect 1291 642 1343 646
rect 1347 642 1455 646
rect 1459 642 1495 646
rect 1499 642 1623 646
rect 1627 642 1791 646
rect 1795 642 1935 646
rect 1939 642 2031 646
rect 2035 642 2055 646
rect 103 641 2055 642
rect 2061 641 2062 647
rect 2042 573 2043 579
rect 2049 578 4015 579
rect 2049 574 2071 578
rect 2075 574 2111 578
rect 2115 574 2215 578
rect 2219 574 2351 578
rect 2355 574 2375 578
rect 2379 574 2487 578
rect 2491 574 2631 578
rect 2635 574 2655 578
rect 2659 574 2791 578
rect 2795 574 2919 578
rect 2923 574 2975 578
rect 2979 574 3175 578
rect 3179 574 3191 578
rect 3195 574 3423 578
rect 3427 574 3671 578
rect 3675 574 3895 578
rect 3899 574 3991 578
rect 3995 574 4015 578
rect 2049 573 4015 574
rect 4021 573 4022 579
rect 84 557 85 563
rect 91 562 2043 563
rect 91 558 111 562
rect 115 558 151 562
rect 155 558 207 562
rect 211 558 255 562
rect 259 558 327 562
rect 331 558 391 562
rect 395 558 447 562
rect 451 558 527 562
rect 531 558 567 562
rect 571 558 663 562
rect 667 558 687 562
rect 691 558 799 562
rect 803 558 807 562
rect 811 558 911 562
rect 915 558 959 562
rect 963 558 1031 562
rect 1035 558 1119 562
rect 1123 558 1151 562
rect 1155 558 1271 562
rect 1275 558 1287 562
rect 1291 558 1455 562
rect 1459 558 1623 562
rect 1627 558 1791 562
rect 1795 558 1935 562
rect 1939 558 2031 562
rect 2035 558 2043 562
rect 91 557 2043 558
rect 2049 557 2050 563
rect 2054 497 2055 503
rect 2061 502 4027 503
rect 2061 498 2071 502
rect 2075 498 2111 502
rect 2115 498 2215 502
rect 2219 498 2351 502
rect 2355 498 2423 502
rect 2427 498 2487 502
rect 2491 498 2527 502
rect 2531 498 2631 502
rect 2635 498 2743 502
rect 2747 498 2791 502
rect 2795 498 2871 502
rect 2875 498 2975 502
rect 2979 498 3031 502
rect 3035 498 3191 502
rect 3195 498 3223 502
rect 3227 498 3423 502
rect 3427 498 3447 502
rect 3451 498 3671 502
rect 3675 498 3679 502
rect 3683 498 3895 502
rect 3899 498 3991 502
rect 3995 498 4027 502
rect 2061 497 4027 498
rect 4033 497 4034 503
rect 96 477 97 483
rect 103 482 2055 483
rect 103 478 111 482
rect 115 478 207 482
rect 211 478 327 482
rect 331 478 439 482
rect 443 478 447 482
rect 451 478 543 482
rect 547 478 567 482
rect 571 478 647 482
rect 651 478 687 482
rect 691 478 751 482
rect 755 478 799 482
rect 803 478 855 482
rect 859 478 911 482
rect 915 478 959 482
rect 963 478 1031 482
rect 1035 478 1063 482
rect 1067 478 1151 482
rect 1155 478 1167 482
rect 1171 478 1271 482
rect 1275 478 1375 482
rect 1379 478 2031 482
rect 2035 478 2055 482
rect 103 477 2055 478
rect 2061 477 2062 483
rect 2042 421 2043 427
rect 2049 426 4015 427
rect 2049 422 2071 426
rect 2075 422 2423 426
rect 2427 422 2527 426
rect 2531 422 2631 426
rect 2635 422 2639 426
rect 2643 422 2743 426
rect 2747 422 2775 426
rect 2779 422 2871 426
rect 2875 422 2951 426
rect 2955 422 3031 426
rect 3035 422 3159 426
rect 3163 422 3223 426
rect 3227 422 3399 426
rect 3403 422 3447 426
rect 3451 422 3655 426
rect 3659 422 3679 426
rect 3683 422 3895 426
rect 3899 422 3991 426
rect 3995 422 4015 426
rect 2049 421 4015 422
rect 4021 421 4022 427
rect 84 397 85 403
rect 91 402 2043 403
rect 91 398 111 402
rect 115 398 439 402
rect 443 398 543 402
rect 547 398 623 402
rect 627 398 647 402
rect 651 398 727 402
rect 731 398 751 402
rect 755 398 831 402
rect 835 398 855 402
rect 859 398 935 402
rect 939 398 959 402
rect 963 398 1039 402
rect 1043 398 1063 402
rect 1067 398 1143 402
rect 1147 398 1167 402
rect 1171 398 1247 402
rect 1251 398 1271 402
rect 1275 398 1351 402
rect 1355 398 1375 402
rect 1379 398 1455 402
rect 1459 398 1559 402
rect 1563 398 2031 402
rect 2035 398 2043 402
rect 91 397 2043 398
rect 2049 397 2050 403
rect 2054 337 2055 343
rect 2061 342 4027 343
rect 2061 338 2071 342
rect 2075 338 2271 342
rect 2275 338 2423 342
rect 2427 338 2527 342
rect 2531 338 2583 342
rect 2587 338 2639 342
rect 2643 338 2743 342
rect 2747 338 2775 342
rect 2779 338 2911 342
rect 2915 338 2951 342
rect 2955 338 3071 342
rect 3075 338 3159 342
rect 3163 338 3223 342
rect 3227 338 3367 342
rect 3371 338 3399 342
rect 3403 338 3503 342
rect 3507 338 3639 342
rect 3643 338 3655 342
rect 3659 338 3775 342
rect 3779 338 3895 342
rect 3899 338 3991 342
rect 3995 338 4027 342
rect 2061 337 4027 338
rect 4033 337 4034 343
rect 96 325 97 331
rect 103 330 2055 331
rect 103 326 111 330
rect 115 326 399 330
rect 403 326 543 330
rect 547 326 623 330
rect 627 326 687 330
rect 691 326 727 330
rect 731 326 831 330
rect 835 326 839 330
rect 843 326 935 330
rect 939 326 991 330
rect 995 326 1039 330
rect 1043 326 1143 330
rect 1147 326 1247 330
rect 1251 326 1303 330
rect 1307 326 1351 330
rect 1355 326 1455 330
rect 1459 326 1463 330
rect 1467 326 1559 330
rect 1563 326 1623 330
rect 1627 326 2031 330
rect 2035 326 2055 330
rect 103 325 2055 326
rect 2061 325 2062 331
rect 2042 257 2043 263
rect 2049 262 4015 263
rect 2049 258 2071 262
rect 2075 258 2111 262
rect 2115 258 2247 262
rect 2251 258 2271 262
rect 2275 258 2423 262
rect 2427 258 2583 262
rect 2587 258 2599 262
rect 2603 258 2743 262
rect 2747 258 2775 262
rect 2779 258 2911 262
rect 2915 258 2943 262
rect 2947 258 3071 262
rect 3075 258 3103 262
rect 3107 258 3223 262
rect 3227 258 3255 262
rect 3259 258 3367 262
rect 3371 258 3391 262
rect 3395 258 3503 262
rect 3507 258 3527 262
rect 3531 258 3639 262
rect 3643 258 3655 262
rect 3659 258 3775 262
rect 3779 258 3783 262
rect 3787 258 3895 262
rect 3899 258 3991 262
rect 3995 258 4015 262
rect 2049 257 4015 258
rect 4021 257 4022 263
rect 2042 255 2050 257
rect 84 249 85 255
rect 91 254 2043 255
rect 91 250 111 254
rect 115 250 207 254
rect 211 250 399 254
rect 403 250 431 254
rect 435 250 543 254
rect 547 250 655 254
rect 659 250 687 254
rect 691 250 839 254
rect 843 250 871 254
rect 875 250 991 254
rect 995 250 1071 254
rect 1075 250 1143 254
rect 1147 250 1263 254
rect 1267 250 1303 254
rect 1307 250 1447 254
rect 1451 250 1463 254
rect 1467 250 1623 254
rect 1627 250 1631 254
rect 1635 250 1815 254
rect 1819 250 2031 254
rect 2035 250 2043 254
rect 91 249 2043 250
rect 2049 249 2050 255
rect 2054 173 2055 179
rect 2061 178 4027 179
rect 2061 174 2071 178
rect 2075 174 2111 178
rect 2115 174 2239 178
rect 2243 174 2247 178
rect 2251 174 2399 178
rect 2403 174 2423 178
rect 2427 174 2567 178
rect 2571 174 2599 178
rect 2603 174 2735 178
rect 2739 174 2775 178
rect 2779 174 2895 178
rect 2899 174 2943 178
rect 2947 174 3047 178
rect 3051 174 3103 178
rect 3107 174 3191 178
rect 3195 174 3255 178
rect 3259 174 3327 178
rect 3331 174 3391 178
rect 3395 174 3455 178
rect 3459 174 3527 178
rect 3531 174 3591 178
rect 3595 174 3655 178
rect 3659 174 3727 178
rect 3731 174 3783 178
rect 3787 174 3895 178
rect 3899 174 3991 178
rect 3995 174 4027 178
rect 2061 173 4027 174
rect 4033 173 4034 179
rect 96 149 97 155
rect 103 154 2055 155
rect 103 150 111 154
rect 115 150 151 154
rect 155 150 207 154
rect 211 150 255 154
rect 259 150 359 154
rect 363 150 431 154
rect 435 150 463 154
rect 467 150 567 154
rect 571 150 655 154
rect 659 150 671 154
rect 675 150 775 154
rect 779 150 871 154
rect 875 150 879 154
rect 883 150 983 154
rect 987 150 1071 154
rect 1075 150 1087 154
rect 1091 150 1191 154
rect 1195 150 1263 154
rect 1267 150 1295 154
rect 1299 150 1399 154
rect 1403 150 1447 154
rect 1451 150 1511 154
rect 1515 150 1623 154
rect 1627 150 1631 154
rect 1635 150 1727 154
rect 1731 150 1815 154
rect 1819 150 1831 154
rect 1835 150 1935 154
rect 1939 150 2031 154
rect 2035 150 2055 154
rect 103 149 2055 150
rect 2061 149 2062 155
rect 2042 101 2043 107
rect 2049 106 4015 107
rect 2049 102 2071 106
rect 2075 102 2111 106
rect 2115 102 2239 106
rect 2243 102 2399 106
rect 2403 102 2567 106
rect 2571 102 2735 106
rect 2739 102 2895 106
rect 2899 102 3047 106
rect 3051 102 3191 106
rect 3195 102 3327 106
rect 3331 102 3455 106
rect 3459 102 3591 106
rect 3595 102 3727 106
rect 3731 102 3991 106
rect 3995 102 4015 106
rect 2049 101 4015 102
rect 4021 101 4022 107
rect 84 77 85 83
rect 91 82 2043 83
rect 91 78 111 82
rect 115 78 151 82
rect 155 78 255 82
rect 259 78 359 82
rect 363 78 463 82
rect 467 78 567 82
rect 571 78 671 82
rect 675 78 775 82
rect 779 78 879 82
rect 883 78 983 82
rect 987 78 1087 82
rect 1091 78 1191 82
rect 1195 78 1295 82
rect 1299 78 1399 82
rect 1403 78 1511 82
rect 1515 78 1623 82
rect 1627 78 1727 82
rect 1731 78 1831 82
rect 1835 78 1935 82
rect 1939 78 2031 82
rect 2035 78 2043 82
rect 91 77 2043 78
rect 2049 77 2050 83
<< m5c >>
rect 2055 4077 2061 4083
rect 4027 4077 4033 4083
rect 97 4041 103 4047
rect 2055 4041 2061 4047
rect 2043 4005 2049 4011
rect 4015 4005 4021 4011
rect 85 3969 91 3975
rect 2043 3969 2049 3975
rect 2055 3929 2061 3935
rect 4027 3929 4033 3935
rect 97 3893 103 3899
rect 2055 3893 2061 3899
rect 2043 3857 2049 3863
rect 4015 3857 4021 3863
rect 85 3813 91 3819
rect 2043 3813 2049 3819
rect 2055 3781 2061 3787
rect 4027 3781 4033 3787
rect 97 3733 103 3739
rect 2055 3733 2061 3739
rect 2043 3701 2049 3707
rect 4015 3701 4021 3707
rect 85 3661 91 3667
rect 2043 3661 2049 3667
rect 2055 3621 2061 3627
rect 4027 3621 4033 3627
rect 97 3589 103 3595
rect 2055 3589 2061 3595
rect 2043 3537 2049 3543
rect 4015 3537 4021 3543
rect 85 3517 91 3523
rect 2043 3517 2049 3523
rect 2055 3465 2061 3471
rect 4027 3465 4033 3471
rect 97 3421 103 3427
rect 2055 3421 2061 3427
rect 2043 3389 2049 3395
rect 4015 3389 4021 3395
rect 85 3341 91 3347
rect 2043 3341 2049 3347
rect 2055 3301 2061 3307
rect 4027 3301 4033 3307
rect 97 3257 103 3263
rect 2055 3257 2061 3263
rect 2043 3229 2049 3235
rect 4015 3229 4021 3235
rect 85 3173 91 3179
rect 2043 3173 2049 3179
rect 2055 3141 2061 3147
rect 4027 3141 4033 3147
rect 97 3085 103 3091
rect 2055 3085 2061 3091
rect 2043 3061 2049 3067
rect 4015 3061 4021 3067
rect 85 3001 91 3007
rect 2043 3001 2049 3007
rect 2055 2989 2061 2995
rect 4027 2989 4033 2995
rect 2043 2927 2049 2933
rect 97 2917 103 2923
rect 2055 2917 2061 2923
rect 4015 2917 4021 2923
rect 2055 2841 2061 2847
rect 4027 2841 4033 2847
rect 85 2829 91 2835
rect 2043 2829 2049 2835
rect 2043 2761 2049 2767
rect 4015 2761 4021 2767
rect 97 2741 103 2747
rect 2055 2741 2061 2747
rect 2055 2673 2061 2679
rect 4027 2673 4033 2679
rect 85 2657 91 2663
rect 2043 2657 2049 2663
rect 2043 2593 2049 2599
rect 4015 2593 4021 2599
rect 97 2569 103 2575
rect 2055 2569 2061 2575
rect 2055 2521 2061 2527
rect 4027 2521 4033 2527
rect 85 2481 91 2487
rect 2043 2481 2049 2487
rect 2043 2441 2049 2447
rect 4015 2441 4021 2447
rect 97 2397 103 2403
rect 2055 2397 2061 2403
rect 2055 2369 2061 2375
rect 4027 2369 4033 2375
rect 85 2313 91 2319
rect 2043 2313 2049 2319
rect 2043 2297 2049 2303
rect 4015 2297 4021 2303
rect 97 2229 103 2235
rect 2055 2229 2061 2235
rect 2055 2217 2061 2223
rect 4027 2217 4033 2223
rect 85 2141 91 2147
rect 2043 2141 2049 2147
rect 2055 2069 2061 2075
rect 4027 2069 4033 2075
rect 97 2057 103 2063
rect 2055 2057 2061 2063
rect 2043 1989 2049 1995
rect 4015 1989 4021 1995
rect 85 1973 91 1979
rect 2043 1973 2049 1979
rect 2055 1913 2061 1919
rect 4027 1913 4033 1919
rect 97 1897 103 1903
rect 2055 1897 2061 1903
rect 2043 1841 2049 1847
rect 4015 1841 4021 1847
rect 85 1813 91 1819
rect 2043 1813 2049 1819
rect 2055 1765 2061 1771
rect 4027 1765 4033 1771
rect 97 1737 103 1743
rect 2055 1737 2061 1743
rect 2043 1685 2049 1691
rect 4015 1685 4021 1691
rect 85 1665 91 1671
rect 2043 1665 2049 1671
rect 2055 1601 2061 1607
rect 4027 1601 4033 1607
rect 97 1585 103 1591
rect 2055 1585 2061 1591
rect 2043 1517 2049 1523
rect 4015 1517 4021 1523
rect 85 1505 91 1511
rect 2043 1505 2049 1511
rect 2055 1441 2061 1447
rect 4027 1441 4033 1447
rect 97 1425 103 1431
rect 2055 1425 2061 1431
rect 2043 1361 2049 1367
rect 4015 1361 4021 1367
rect 85 1341 91 1347
rect 2043 1341 2049 1347
rect 2055 1281 2061 1287
rect 4027 1281 4033 1287
rect 97 1269 103 1275
rect 2055 1269 2061 1275
rect 2043 1205 2049 1211
rect 4015 1205 4021 1211
rect 85 1189 91 1195
rect 2043 1189 2049 1195
rect 2055 1129 2061 1135
rect 4027 1129 4033 1135
rect 97 1109 103 1115
rect 2055 1109 2061 1115
rect 2043 1049 2049 1055
rect 4015 1049 4021 1055
rect 85 1029 91 1035
rect 2043 1029 2049 1035
rect 2055 969 2061 975
rect 4027 969 4033 975
rect 97 949 103 955
rect 2055 949 2061 955
rect 2043 885 2049 891
rect 4015 885 4021 891
rect 85 869 91 875
rect 2043 869 2049 875
rect 2055 813 2061 819
rect 4027 813 4033 819
rect 97 797 103 803
rect 2055 797 2061 803
rect 2043 733 2049 739
rect 4015 733 4021 739
rect 85 721 91 727
rect 2043 721 2049 727
rect 2055 657 2061 663
rect 4027 657 4033 663
rect 97 641 103 647
rect 2055 641 2061 647
rect 2043 573 2049 579
rect 4015 573 4021 579
rect 85 557 91 563
rect 2043 557 2049 563
rect 2055 497 2061 503
rect 4027 497 4033 503
rect 97 477 103 483
rect 2055 477 2061 483
rect 2043 421 2049 427
rect 4015 421 4021 427
rect 85 397 91 403
rect 2043 397 2049 403
rect 2055 337 2061 343
rect 4027 337 4033 343
rect 97 325 103 331
rect 2055 325 2061 331
rect 2043 257 2049 263
rect 4015 257 4021 263
rect 85 249 91 255
rect 2043 249 2049 255
rect 2055 173 2061 179
rect 4027 173 4033 179
rect 97 149 103 155
rect 2055 149 2061 155
rect 2043 101 2049 107
rect 4015 101 4021 107
rect 85 77 91 83
rect 2043 77 2049 83
<< m5 >>
rect 84 3975 92 4104
rect 84 3969 85 3975
rect 91 3969 92 3975
rect 84 3819 92 3969
rect 84 3813 85 3819
rect 91 3813 92 3819
rect 84 3667 92 3813
rect 84 3661 85 3667
rect 91 3661 92 3667
rect 84 3523 92 3661
rect 84 3517 85 3523
rect 91 3517 92 3523
rect 84 3347 92 3517
rect 84 3341 85 3347
rect 91 3341 92 3347
rect 84 3179 92 3341
rect 84 3173 85 3179
rect 91 3173 92 3179
rect 84 3007 92 3173
rect 84 3001 85 3007
rect 91 3001 92 3007
rect 84 2835 92 3001
rect 84 2829 85 2835
rect 91 2829 92 2835
rect 84 2663 92 2829
rect 84 2657 85 2663
rect 91 2657 92 2663
rect 84 2487 92 2657
rect 84 2481 85 2487
rect 91 2481 92 2487
rect 84 2319 92 2481
rect 84 2313 85 2319
rect 91 2313 92 2319
rect 84 2147 92 2313
rect 84 2141 85 2147
rect 91 2141 92 2147
rect 84 1979 92 2141
rect 84 1973 85 1979
rect 91 1973 92 1979
rect 84 1819 92 1973
rect 84 1813 85 1819
rect 91 1813 92 1819
rect 84 1671 92 1813
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1511 92 1665
rect 84 1505 85 1511
rect 91 1505 92 1511
rect 84 1347 92 1505
rect 84 1341 85 1347
rect 91 1341 92 1347
rect 84 1195 92 1341
rect 84 1189 85 1195
rect 91 1189 92 1195
rect 84 1035 92 1189
rect 84 1029 85 1035
rect 91 1029 92 1035
rect 84 875 92 1029
rect 84 869 85 875
rect 91 869 92 875
rect 84 727 92 869
rect 84 721 85 727
rect 91 721 92 727
rect 84 563 92 721
rect 84 557 85 563
rect 91 557 92 563
rect 84 403 92 557
rect 84 397 85 403
rect 91 397 92 403
rect 84 255 92 397
rect 84 249 85 255
rect 91 249 92 255
rect 84 83 92 249
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 4047 104 4104
rect 96 4041 97 4047
rect 103 4041 104 4047
rect 96 3899 104 4041
rect 96 3893 97 3899
rect 103 3893 104 3899
rect 96 3739 104 3893
rect 96 3733 97 3739
rect 103 3733 104 3739
rect 96 3595 104 3733
rect 96 3589 97 3595
rect 103 3589 104 3595
rect 96 3427 104 3589
rect 96 3421 97 3427
rect 103 3421 104 3427
rect 96 3263 104 3421
rect 96 3257 97 3263
rect 103 3257 104 3263
rect 96 3091 104 3257
rect 96 3085 97 3091
rect 103 3085 104 3091
rect 96 2923 104 3085
rect 96 2917 97 2923
rect 103 2917 104 2923
rect 96 2747 104 2917
rect 96 2741 97 2747
rect 103 2741 104 2747
rect 96 2575 104 2741
rect 96 2569 97 2575
rect 103 2569 104 2575
rect 96 2403 104 2569
rect 96 2397 97 2403
rect 103 2397 104 2403
rect 96 2235 104 2397
rect 96 2229 97 2235
rect 103 2229 104 2235
rect 96 2063 104 2229
rect 96 2057 97 2063
rect 103 2057 104 2063
rect 96 1903 104 2057
rect 96 1897 97 1903
rect 103 1897 104 1903
rect 96 1743 104 1897
rect 96 1737 97 1743
rect 103 1737 104 1743
rect 96 1591 104 1737
rect 96 1585 97 1591
rect 103 1585 104 1591
rect 96 1431 104 1585
rect 96 1425 97 1431
rect 103 1425 104 1431
rect 96 1275 104 1425
rect 96 1269 97 1275
rect 103 1269 104 1275
rect 96 1115 104 1269
rect 96 1109 97 1115
rect 103 1109 104 1115
rect 96 955 104 1109
rect 96 949 97 955
rect 103 949 104 955
rect 96 803 104 949
rect 96 797 97 803
rect 103 797 104 803
rect 96 647 104 797
rect 96 641 97 647
rect 103 641 104 647
rect 96 483 104 641
rect 96 477 97 483
rect 103 477 104 483
rect 96 331 104 477
rect 96 325 97 331
rect 103 325 104 331
rect 96 155 104 325
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 2042 4011 2050 4104
rect 2042 4005 2043 4011
rect 2049 4005 2050 4011
rect 2042 3975 2050 4005
rect 2042 3969 2043 3975
rect 2049 3969 2050 3975
rect 2042 3863 2050 3969
rect 2042 3857 2043 3863
rect 2049 3857 2050 3863
rect 2042 3819 2050 3857
rect 2042 3813 2043 3819
rect 2049 3813 2050 3819
rect 2042 3707 2050 3813
rect 2042 3701 2043 3707
rect 2049 3701 2050 3707
rect 2042 3667 2050 3701
rect 2042 3661 2043 3667
rect 2049 3661 2050 3667
rect 2042 3543 2050 3661
rect 2042 3537 2043 3543
rect 2049 3537 2050 3543
rect 2042 3523 2050 3537
rect 2042 3517 2043 3523
rect 2049 3517 2050 3523
rect 2042 3395 2050 3517
rect 2042 3389 2043 3395
rect 2049 3389 2050 3395
rect 2042 3347 2050 3389
rect 2042 3341 2043 3347
rect 2049 3341 2050 3347
rect 2042 3235 2050 3341
rect 2042 3229 2043 3235
rect 2049 3229 2050 3235
rect 2042 3179 2050 3229
rect 2042 3173 2043 3179
rect 2049 3173 2050 3179
rect 2042 3067 2050 3173
rect 2042 3061 2043 3067
rect 2049 3061 2050 3067
rect 2042 3007 2050 3061
rect 2042 3001 2043 3007
rect 2049 3001 2050 3007
rect 2042 2933 2050 3001
rect 2042 2927 2043 2933
rect 2049 2927 2050 2933
rect 2042 2835 2050 2927
rect 2042 2829 2043 2835
rect 2049 2829 2050 2835
rect 2042 2767 2050 2829
rect 2042 2761 2043 2767
rect 2049 2761 2050 2767
rect 2042 2663 2050 2761
rect 2042 2657 2043 2663
rect 2049 2657 2050 2663
rect 2042 2599 2050 2657
rect 2042 2593 2043 2599
rect 2049 2593 2050 2599
rect 2042 2487 2050 2593
rect 2042 2481 2043 2487
rect 2049 2481 2050 2487
rect 2042 2447 2050 2481
rect 2042 2441 2043 2447
rect 2049 2441 2050 2447
rect 2042 2319 2050 2441
rect 2042 2313 2043 2319
rect 2049 2313 2050 2319
rect 2042 2303 2050 2313
rect 2042 2297 2043 2303
rect 2049 2297 2050 2303
rect 2042 2147 2050 2297
rect 2042 2141 2043 2147
rect 2049 2141 2050 2147
rect 2042 1995 2050 2141
rect 2042 1989 2043 1995
rect 2049 1989 2050 1995
rect 2042 1979 2050 1989
rect 2042 1973 2043 1979
rect 2049 1973 2050 1979
rect 2042 1847 2050 1973
rect 2042 1841 2043 1847
rect 2049 1841 2050 1847
rect 2042 1819 2050 1841
rect 2042 1813 2043 1819
rect 2049 1813 2050 1819
rect 2042 1691 2050 1813
rect 2042 1685 2043 1691
rect 2049 1685 2050 1691
rect 2042 1671 2050 1685
rect 2042 1665 2043 1671
rect 2049 1665 2050 1671
rect 2042 1523 2050 1665
rect 2042 1517 2043 1523
rect 2049 1517 2050 1523
rect 2042 1511 2050 1517
rect 2042 1505 2043 1511
rect 2049 1505 2050 1511
rect 2042 1367 2050 1505
rect 2042 1361 2043 1367
rect 2049 1361 2050 1367
rect 2042 1347 2050 1361
rect 2042 1341 2043 1347
rect 2049 1341 2050 1347
rect 2042 1211 2050 1341
rect 2042 1205 2043 1211
rect 2049 1205 2050 1211
rect 2042 1195 2050 1205
rect 2042 1189 2043 1195
rect 2049 1189 2050 1195
rect 2042 1055 2050 1189
rect 2042 1049 2043 1055
rect 2049 1049 2050 1055
rect 2042 1035 2050 1049
rect 2042 1029 2043 1035
rect 2049 1029 2050 1035
rect 2042 891 2050 1029
rect 2042 885 2043 891
rect 2049 885 2050 891
rect 2042 875 2050 885
rect 2042 869 2043 875
rect 2049 869 2050 875
rect 2042 739 2050 869
rect 2042 733 2043 739
rect 2049 733 2050 739
rect 2042 727 2050 733
rect 2042 721 2043 727
rect 2049 721 2050 727
rect 2042 579 2050 721
rect 2042 573 2043 579
rect 2049 573 2050 579
rect 2042 563 2050 573
rect 2042 557 2043 563
rect 2049 557 2050 563
rect 2042 427 2050 557
rect 2042 421 2043 427
rect 2049 421 2050 427
rect 2042 403 2050 421
rect 2042 397 2043 403
rect 2049 397 2050 403
rect 2042 263 2050 397
rect 2042 257 2043 263
rect 2049 257 2050 263
rect 2042 255 2050 257
rect 2042 249 2043 255
rect 2049 249 2050 255
rect 2042 107 2050 249
rect 2042 101 2043 107
rect 2049 101 2050 107
rect 2042 83 2050 101
rect 2042 77 2043 83
rect 2049 77 2050 83
rect 2042 72 2050 77
rect 2054 4083 2062 4104
rect 2054 4077 2055 4083
rect 2061 4077 2062 4083
rect 2054 4047 2062 4077
rect 2054 4041 2055 4047
rect 2061 4041 2062 4047
rect 2054 3935 2062 4041
rect 2054 3929 2055 3935
rect 2061 3929 2062 3935
rect 2054 3899 2062 3929
rect 2054 3893 2055 3899
rect 2061 3893 2062 3899
rect 2054 3787 2062 3893
rect 2054 3781 2055 3787
rect 2061 3781 2062 3787
rect 2054 3739 2062 3781
rect 2054 3733 2055 3739
rect 2061 3733 2062 3739
rect 2054 3627 2062 3733
rect 2054 3621 2055 3627
rect 2061 3621 2062 3627
rect 2054 3595 2062 3621
rect 2054 3589 2055 3595
rect 2061 3589 2062 3595
rect 2054 3471 2062 3589
rect 2054 3465 2055 3471
rect 2061 3465 2062 3471
rect 2054 3427 2062 3465
rect 2054 3421 2055 3427
rect 2061 3421 2062 3427
rect 2054 3307 2062 3421
rect 2054 3301 2055 3307
rect 2061 3301 2062 3307
rect 2054 3263 2062 3301
rect 2054 3257 2055 3263
rect 2061 3257 2062 3263
rect 2054 3147 2062 3257
rect 2054 3141 2055 3147
rect 2061 3141 2062 3147
rect 2054 3091 2062 3141
rect 2054 3085 2055 3091
rect 2061 3085 2062 3091
rect 2054 2995 2062 3085
rect 2054 2989 2055 2995
rect 2061 2989 2062 2995
rect 2054 2923 2062 2989
rect 2054 2917 2055 2923
rect 2061 2917 2062 2923
rect 2054 2847 2062 2917
rect 2054 2841 2055 2847
rect 2061 2841 2062 2847
rect 2054 2747 2062 2841
rect 2054 2741 2055 2747
rect 2061 2741 2062 2747
rect 2054 2679 2062 2741
rect 2054 2673 2055 2679
rect 2061 2673 2062 2679
rect 2054 2575 2062 2673
rect 2054 2569 2055 2575
rect 2061 2569 2062 2575
rect 2054 2527 2062 2569
rect 2054 2521 2055 2527
rect 2061 2521 2062 2527
rect 2054 2403 2062 2521
rect 2054 2397 2055 2403
rect 2061 2397 2062 2403
rect 2054 2375 2062 2397
rect 2054 2369 2055 2375
rect 2061 2369 2062 2375
rect 2054 2235 2062 2369
rect 2054 2229 2055 2235
rect 2061 2229 2062 2235
rect 2054 2223 2062 2229
rect 2054 2217 2055 2223
rect 2061 2217 2062 2223
rect 2054 2075 2062 2217
rect 2054 2069 2055 2075
rect 2061 2069 2062 2075
rect 2054 2063 2062 2069
rect 2054 2057 2055 2063
rect 2061 2057 2062 2063
rect 2054 1919 2062 2057
rect 2054 1913 2055 1919
rect 2061 1913 2062 1919
rect 2054 1903 2062 1913
rect 2054 1897 2055 1903
rect 2061 1897 2062 1903
rect 2054 1771 2062 1897
rect 2054 1765 2055 1771
rect 2061 1765 2062 1771
rect 2054 1743 2062 1765
rect 2054 1737 2055 1743
rect 2061 1737 2062 1743
rect 2054 1607 2062 1737
rect 2054 1601 2055 1607
rect 2061 1601 2062 1607
rect 2054 1591 2062 1601
rect 2054 1585 2055 1591
rect 2061 1585 2062 1591
rect 2054 1447 2062 1585
rect 2054 1441 2055 1447
rect 2061 1441 2062 1447
rect 2054 1431 2062 1441
rect 2054 1425 2055 1431
rect 2061 1425 2062 1431
rect 2054 1287 2062 1425
rect 2054 1281 2055 1287
rect 2061 1281 2062 1287
rect 2054 1275 2062 1281
rect 2054 1269 2055 1275
rect 2061 1269 2062 1275
rect 2054 1135 2062 1269
rect 2054 1129 2055 1135
rect 2061 1129 2062 1135
rect 2054 1115 2062 1129
rect 2054 1109 2055 1115
rect 2061 1109 2062 1115
rect 2054 975 2062 1109
rect 2054 969 2055 975
rect 2061 969 2062 975
rect 2054 955 2062 969
rect 2054 949 2055 955
rect 2061 949 2062 955
rect 2054 819 2062 949
rect 2054 813 2055 819
rect 2061 813 2062 819
rect 2054 803 2062 813
rect 2054 797 2055 803
rect 2061 797 2062 803
rect 2054 663 2062 797
rect 2054 657 2055 663
rect 2061 657 2062 663
rect 2054 647 2062 657
rect 2054 641 2055 647
rect 2061 641 2062 647
rect 2054 503 2062 641
rect 2054 497 2055 503
rect 2061 497 2062 503
rect 2054 483 2062 497
rect 2054 477 2055 483
rect 2061 477 2062 483
rect 2054 343 2062 477
rect 2054 337 2055 343
rect 2061 337 2062 343
rect 2054 331 2062 337
rect 2054 325 2055 331
rect 2061 325 2062 331
rect 2054 179 2062 325
rect 2054 173 2055 179
rect 2061 173 2062 179
rect 2054 155 2062 173
rect 2054 149 2055 155
rect 2061 149 2062 155
rect 2054 72 2062 149
rect 4014 4011 4022 4104
rect 4014 4005 4015 4011
rect 4021 4005 4022 4011
rect 4014 3863 4022 4005
rect 4014 3857 4015 3863
rect 4021 3857 4022 3863
rect 4014 3707 4022 3857
rect 4014 3701 4015 3707
rect 4021 3701 4022 3707
rect 4014 3543 4022 3701
rect 4014 3537 4015 3543
rect 4021 3537 4022 3543
rect 4014 3395 4022 3537
rect 4014 3389 4015 3395
rect 4021 3389 4022 3395
rect 4014 3235 4022 3389
rect 4014 3229 4015 3235
rect 4021 3229 4022 3235
rect 4014 3067 4022 3229
rect 4014 3061 4015 3067
rect 4021 3061 4022 3067
rect 4014 2923 4022 3061
rect 4014 2917 4015 2923
rect 4021 2917 4022 2923
rect 4014 2767 4022 2917
rect 4014 2761 4015 2767
rect 4021 2761 4022 2767
rect 4014 2599 4022 2761
rect 4014 2593 4015 2599
rect 4021 2593 4022 2599
rect 4014 2447 4022 2593
rect 4014 2441 4015 2447
rect 4021 2441 4022 2447
rect 4014 2303 4022 2441
rect 4014 2297 4015 2303
rect 4021 2297 4022 2303
rect 4014 1995 4022 2297
rect 4014 1989 4015 1995
rect 4021 1989 4022 1995
rect 4014 1847 4022 1989
rect 4014 1841 4015 1847
rect 4021 1841 4022 1847
rect 4014 1691 4022 1841
rect 4014 1685 4015 1691
rect 4021 1685 4022 1691
rect 4014 1523 4022 1685
rect 4014 1517 4015 1523
rect 4021 1517 4022 1523
rect 4014 1367 4022 1517
rect 4014 1361 4015 1367
rect 4021 1361 4022 1367
rect 4014 1211 4022 1361
rect 4014 1205 4015 1211
rect 4021 1205 4022 1211
rect 4014 1055 4022 1205
rect 4014 1049 4015 1055
rect 4021 1049 4022 1055
rect 4014 891 4022 1049
rect 4014 885 4015 891
rect 4021 885 4022 891
rect 4014 739 4022 885
rect 4014 733 4015 739
rect 4021 733 4022 739
rect 4014 579 4022 733
rect 4014 573 4015 579
rect 4021 573 4022 579
rect 4014 427 4022 573
rect 4014 421 4015 427
rect 4021 421 4022 427
rect 4014 263 4022 421
rect 4014 257 4015 263
rect 4021 257 4022 263
rect 4014 107 4022 257
rect 4014 101 4015 107
rect 4021 101 4022 107
rect 4014 72 4022 101
rect 4026 4083 4034 4104
rect 4026 4077 4027 4083
rect 4033 4077 4034 4083
rect 4026 3935 4034 4077
rect 4026 3929 4027 3935
rect 4033 3929 4034 3935
rect 4026 3787 4034 3929
rect 4026 3781 4027 3787
rect 4033 3781 4034 3787
rect 4026 3627 4034 3781
rect 4026 3621 4027 3627
rect 4033 3621 4034 3627
rect 4026 3471 4034 3621
rect 4026 3465 4027 3471
rect 4033 3465 4034 3471
rect 4026 3307 4034 3465
rect 4026 3301 4027 3307
rect 4033 3301 4034 3307
rect 4026 3147 4034 3301
rect 4026 3141 4027 3147
rect 4033 3141 4034 3147
rect 4026 2995 4034 3141
rect 4026 2989 4027 2995
rect 4033 2989 4034 2995
rect 4026 2847 4034 2989
rect 4026 2841 4027 2847
rect 4033 2841 4034 2847
rect 4026 2679 4034 2841
rect 4026 2673 4027 2679
rect 4033 2673 4034 2679
rect 4026 2527 4034 2673
rect 4026 2521 4027 2527
rect 4033 2521 4034 2527
rect 4026 2375 4034 2521
rect 4026 2369 4027 2375
rect 4033 2369 4034 2375
rect 4026 2223 4034 2369
rect 4026 2217 4027 2223
rect 4033 2217 4034 2223
rect 4026 2075 4034 2217
rect 4026 2069 4027 2075
rect 4033 2069 4034 2075
rect 4026 1919 4034 2069
rect 4026 1913 4027 1919
rect 4033 1913 4034 1919
rect 4026 1771 4034 1913
rect 4026 1765 4027 1771
rect 4033 1765 4034 1771
rect 4026 1607 4034 1765
rect 4026 1601 4027 1607
rect 4033 1601 4034 1607
rect 4026 1447 4034 1601
rect 4026 1441 4027 1447
rect 4033 1441 4034 1447
rect 4026 1287 4034 1441
rect 4026 1281 4027 1287
rect 4033 1281 4034 1287
rect 4026 1135 4034 1281
rect 4026 1129 4027 1135
rect 4033 1129 4034 1135
rect 4026 975 4034 1129
rect 4026 969 4027 975
rect 4033 969 4034 975
rect 4026 819 4034 969
rect 4026 813 4027 819
rect 4033 813 4034 819
rect 4026 663 4034 813
rect 4026 657 4027 663
rect 4033 657 4034 663
rect 4026 503 4034 657
rect 4026 497 4027 503
rect 4033 497 4034 503
rect 4026 343 4034 497
rect 4026 337 4027 343
rect 4033 337 4034 343
rect 4026 179 4034 337
rect 4026 173 4027 179
rect 4033 173 4034 179
rect 4026 72 4034 173
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__199
timestamp 1731220536
transform 1 0 3984 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220536
transform 1 0 2064 0 1 4024
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220536
transform 1 0 3984 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220536
transform 1 0 2064 0 -1 3992
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220536
transform 1 0 3984 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220536
transform 1 0 2064 0 1 3876
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220536
transform 1 0 3984 0 -1 3844
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220536
transform 1 0 2064 0 -1 3844
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220536
transform 1 0 3984 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220536
transform 1 0 2064 0 1 3728
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220536
transform 1 0 3984 0 -1 3688
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220536
transform 1 0 2064 0 -1 3688
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220536
transform 1 0 3984 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220536
transform 1 0 2064 0 1 3568
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220536
transform 1 0 3984 0 -1 3524
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220536
transform 1 0 2064 0 -1 3524
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220536
transform 1 0 3984 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220536
transform 1 0 2064 0 1 3412
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220536
transform 1 0 3984 0 -1 3376
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220536
transform 1 0 2064 0 -1 3376
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220536
transform 1 0 3984 0 1 3248
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220536
transform 1 0 2064 0 1 3248
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220536
transform 1 0 3984 0 -1 3216
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220536
transform 1 0 2064 0 -1 3216
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220536
transform 1 0 3984 0 1 3088
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220536
transform 1 0 2064 0 1 3088
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220536
transform 1 0 3984 0 -1 3048
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220536
transform 1 0 2064 0 -1 3048
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220536
transform 1 0 3984 0 1 2936
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220536
transform 1 0 2064 0 1 2936
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220536
transform 1 0 3984 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220536
transform 1 0 2064 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220536
transform 1 0 3984 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220536
transform 1 0 2064 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220536
transform 1 0 3984 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220536
transform 1 0 2064 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220536
transform 1 0 3984 0 1 2620
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220536
transform 1 0 2064 0 1 2620
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220536
transform 1 0 3984 0 -1 2580
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220536
transform 1 0 2064 0 -1 2580
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220536
transform 1 0 3984 0 1 2468
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220536
transform 1 0 2064 0 1 2468
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220536
transform 1 0 3984 0 -1 2428
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220536
transform 1 0 2064 0 -1 2428
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220536
transform 1 0 3984 0 1 2316
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220536
transform 1 0 2064 0 1 2316
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220536
transform 1 0 3984 0 -1 2284
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220536
transform 1 0 2064 0 -1 2284
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220536
transform 1 0 3984 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220536
transform 1 0 2064 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220536
transform 1 0 3984 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220536
transform 1 0 2064 0 -1 2132
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220536
transform 1 0 3984 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220536
transform 1 0 2064 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220536
transform 1 0 3984 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220536
transform 1 0 2064 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220536
transform 1 0 3984 0 1 1860
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220536
transform 1 0 2064 0 1 1860
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220536
transform 1 0 3984 0 -1 1828
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220536
transform 1 0 2064 0 -1 1828
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220536
transform 1 0 3984 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220536
transform 1 0 2064 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220536
transform 1 0 3984 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220536
transform 1 0 2064 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220536
transform 1 0 3984 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220536
transform 1 0 2064 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220536
transform 1 0 3984 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220536
transform 1 0 2064 0 -1 1504
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220536
transform 1 0 3984 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220536
transform 1 0 2064 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220536
transform 1 0 3984 0 -1 1348
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220536
transform 1 0 2064 0 -1 1348
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220536
transform 1 0 3984 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220536
transform 1 0 2064 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220536
transform 1 0 3984 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220536
transform 1 0 2064 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220536
transform 1 0 3984 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220536
transform 1 0 2064 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220536
transform 1 0 3984 0 -1 1036
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220536
transform 1 0 2064 0 -1 1036
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220536
transform 1 0 3984 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220536
transform 1 0 2064 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220536
transform 1 0 3984 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220536
transform 1 0 2064 0 -1 872
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220536
transform 1 0 3984 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220536
transform 1 0 2064 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220536
transform 1 0 3984 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220536
transform 1 0 2064 0 -1 720
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220536
transform 1 0 3984 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220536
transform 1 0 2064 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220536
transform 1 0 3984 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220536
transform 1 0 2064 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220536
transform 1 0 3984 0 1 444
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220536
transform 1 0 2064 0 1 444
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220536
transform 1 0 3984 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220536
transform 1 0 2064 0 -1 408
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220536
transform 1 0 3984 0 1 284
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220536
transform 1 0 2064 0 1 284
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220536
transform 1 0 3984 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220536
transform 1 0 2064 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220536
transform 1 0 3984 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220536
transform 1 0 2064 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220536
transform 1 0 2024 0 1 3988
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220536
transform 1 0 104 0 1 3988
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220536
transform 1 0 2024 0 -1 3956
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220536
transform 1 0 104 0 -1 3956
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220536
transform 1 0 2024 0 1 3840
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220536
transform 1 0 104 0 1 3840
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220536
transform 1 0 2024 0 -1 3800
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220536
transform 1 0 104 0 -1 3800
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220536
transform 1 0 2024 0 1 3680
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220536
transform 1 0 104 0 1 3680
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220536
transform 1 0 2024 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220536
transform 1 0 104 0 -1 3648
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220536
transform 1 0 2024 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220536
transform 1 0 104 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220536
transform 1 0 2024 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220536
transform 1 0 104 0 -1 3504
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220536
transform 1 0 2024 0 1 3368
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220536
transform 1 0 104 0 1 3368
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220536
transform 1 0 2024 0 -1 3328
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220536
transform 1 0 104 0 -1 3328
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220536
transform 1 0 2024 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220536
transform 1 0 104 0 1 3204
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220536
transform 1 0 2024 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220536
transform 1 0 104 0 -1 3160
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220536
transform 1 0 2024 0 1 3032
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220536
transform 1 0 104 0 1 3032
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220536
transform 1 0 2024 0 -1 2988
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220536
transform 1 0 104 0 -1 2988
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220536
transform 1 0 2024 0 1 2864
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220536
transform 1 0 104 0 1 2864
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220536
transform 1 0 2024 0 -1 2816
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220536
transform 1 0 104 0 -1 2816
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220536
transform 1 0 2024 0 1 2688
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220536
transform 1 0 104 0 1 2688
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220536
transform 1 0 2024 0 -1 2644
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220536
transform 1 0 104 0 -1 2644
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220536
transform 1 0 2024 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220536
transform 1 0 104 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220536
transform 1 0 2024 0 -1 2468
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220536
transform 1 0 104 0 -1 2468
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220536
transform 1 0 2024 0 1 2344
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220536
transform 1 0 104 0 1 2344
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220536
transform 1 0 2024 0 -1 2300
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220536
transform 1 0 104 0 -1 2300
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220536
transform 1 0 2024 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220536
transform 1 0 104 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220536
transform 1 0 2024 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220536
transform 1 0 104 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220536
transform 1 0 2024 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220536
transform 1 0 104 0 1 2004
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220536
transform 1 0 2024 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220536
transform 1 0 104 0 -1 1960
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220536
transform 1 0 2024 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220536
transform 1 0 104 0 1 1844
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220536
transform 1 0 2024 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220536
transform 1 0 104 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220536
transform 1 0 2024 0 1 1684
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220536
transform 1 0 104 0 1 1684
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220536
transform 1 0 2024 0 -1 1652
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220536
transform 1 0 104 0 -1 1652
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220536
transform 1 0 2024 0 1 1532
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220536
transform 1 0 104 0 1 1532
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220536
transform 1 0 2024 0 -1 1492
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220536
transform 1 0 104 0 -1 1492
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220536
transform 1 0 2024 0 1 1372
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220536
transform 1 0 104 0 1 1372
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220536
transform 1 0 2024 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220536
transform 1 0 104 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220536
transform 1 0 2024 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220536
transform 1 0 104 0 1 1216
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220536
transform 1 0 2024 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220536
transform 1 0 104 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220536
transform 1 0 2024 0 1 1056
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220536
transform 1 0 104 0 1 1056
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220536
transform 1 0 2024 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220536
transform 1 0 104 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220536
transform 1 0 2024 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220536
transform 1 0 104 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220536
transform 1 0 2024 0 -1 856
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220536
transform 1 0 104 0 -1 856
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220536
transform 1 0 2024 0 1 744
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220536
transform 1 0 104 0 1 744
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220536
transform 1 0 2024 0 -1 708
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220536
transform 1 0 104 0 -1 708
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220536
transform 1 0 2024 0 1 588
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220536
transform 1 0 104 0 1 588
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220536
transform 1 0 2024 0 -1 544
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220536
transform 1 0 104 0 -1 544
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220536
transform 1 0 2024 0 1 424
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220536
transform 1 0 104 0 1 424
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220536
transform 1 0 2024 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220536
transform 1 0 104 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220536
transform 1 0 2024 0 1 272
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220536
transform 1 0 104 0 1 272
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220536
transform 1 0 2024 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220536
transform 1 0 104 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220536
transform 1 0 2024 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220536
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCH  tst_5999_6
timestamp 1731220536
transform 1 0 3688 0 1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5998_6
timestamp 1731220536
transform 1 0 3584 0 1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5997_6
timestamp 1731220536
transform 1 0 3480 0 1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5996_6
timestamp 1731220536
transform 1 0 3376 0 1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5995_6
timestamp 1731220536
transform 1 0 3528 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5994_6
timestamp 1731220536
transform 1 0 3392 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5993_6
timestamp 1731220536
transform 1 0 3264 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5992_6
timestamp 1731220536
transform 1 0 3136 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5991_6
timestamp 1731220536
transform 1 0 3008 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5990_6
timestamp 1731220536
transform 1 0 3232 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5989_6
timestamp 1731220536
transform 1 0 3080 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5988_6
timestamp 1731220536
transform 1 0 2928 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5987_6
timestamp 1731220536
transform 1 0 2776 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5986_6
timestamp 1731220536
transform 1 0 3144 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5985_6
timestamp 1731220536
transform 1 0 3000 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5984_6
timestamp 1731220536
transform 1 0 2856 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5983_6
timestamp 1731220536
transform 1 0 2720 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5982_6
timestamp 1731220536
transform 1 0 2800 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5981_6
timestamp 1731220536
transform 1 0 2928 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5980_6
timestamp 1731220536
transform 1 0 3200 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5979_6
timestamp 1731220536
transform 1 0 3064 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5978_6
timestamp 1731220536
transform 1 0 2992 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5977_6
timestamp 1731220536
transform 1 0 2824 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5976_6
timestamp 1731220536
transform 1 0 3160 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5975_6
timestamp 1731220536
transform 1 0 3336 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5974_6
timestamp 1731220536
transform 1 0 3280 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5973_6
timestamp 1731220536
transform 1 0 3144 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5972_6
timestamp 1731220536
transform 1 0 3000 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5971_6
timestamp 1731220536
transform 1 0 2840 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5970_6
timestamp 1731220536
transform 1 0 2840 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5969_6
timestamp 1731220536
transform 1 0 2968 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5968_6
timestamp 1731220536
transform 1 0 3096 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5967_6
timestamp 1731220536
transform 1 0 3216 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5966_6
timestamp 1731220536
transform 1 0 3328 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5965_6
timestamp 1731220536
transform 1 0 3440 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5964_6
timestamp 1731220536
transform 1 0 3768 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5963_6
timestamp 1731220536
transform 1 0 3664 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5962_6
timestamp 1731220536
transform 1 0 3552 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5961_6
timestamp 1731220536
transform 1 0 3528 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5960_6
timestamp 1731220536
transform 1 0 3408 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5959_6
timestamp 1731220536
transform 1 0 3648 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5958_6
timestamp 1731220536
transform 1 0 3768 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5957_6
timestamp 1731220536
transform 1 0 3872 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5956_6
timestamp 1731220536
transform 1 0 3872 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5955_6
timestamp 1731220536
transform 1 0 3872 0 1 3396
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5954_6
timestamp 1731220536
transform 1 0 3872 0 -1 3392
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5953_6
timestamp 1731220536
transform 1 0 3760 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5952_6
timestamp 1731220536
transform 1 0 3872 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5951_6
timestamp 1731220536
transform 1 0 3872 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5950_6
timestamp 1731220536
transform 1 0 3768 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5949_6
timestamp 1731220536
transform 1 0 3648 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5948_6
timestamp 1731220536
transform 1 0 3528 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5947_6
timestamp 1731220536
transform 1 0 3624 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5946_6
timestamp 1731220536
transform 1 0 3488 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5945_6
timestamp 1731220536
transform 1 0 3352 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5944_6
timestamp 1731220536
transform 1 0 3208 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5943_6
timestamp 1731220536
transform 1 0 3048 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5942_6
timestamp 1731220536
transform 1 0 2872 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5941_6
timestamp 1731220536
transform 1 0 3408 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5940_6
timestamp 1731220536
transform 1 0 3280 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5939_6
timestamp 1731220536
transform 1 0 3144 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5938_6
timestamp 1731220536
transform 1 0 3008 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5937_6
timestamp 1731220536
transform 1 0 2856 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5936_6
timestamp 1731220536
transform 1 0 3424 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5935_6
timestamp 1731220536
transform 1 0 3240 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5934_6
timestamp 1731220536
transform 1 0 3064 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5933_6
timestamp 1731220536
transform 1 0 2888 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5932_6
timestamp 1731220536
transform 1 0 3272 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5931_6
timestamp 1731220536
transform 1 0 3144 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5930_6
timestamp 1731220536
transform 1 0 3024 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5929_6
timestamp 1731220536
transform 1 0 2904 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5928_6
timestamp 1731220536
transform 1 0 3200 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5927_6
timestamp 1731220536
transform 1 0 3096 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5926_6
timestamp 1731220536
transform 1 0 2992 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5925_6
timestamp 1731220536
transform 1 0 2888 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5924_6
timestamp 1731220536
transform 1 0 2912 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5923_6
timestamp 1731220536
transform 1 0 3016 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5922_6
timestamp 1731220536
transform 1 0 3120 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5921_6
timestamp 1731220536
transform 1 0 3224 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5920_6
timestamp 1731220536
transform 1 0 3216 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5919_6
timestamp 1731220536
transform 1 0 3112 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5918_6
timestamp 1731220536
transform 1 0 3008 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5917_6
timestamp 1731220536
transform 1 0 2904 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5916_6
timestamp 1731220536
transform 1 0 2872 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5915_6
timestamp 1731220536
transform 1 0 2992 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5914_6
timestamp 1731220536
transform 1 0 3120 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5913_6
timestamp 1731220536
transform 1 0 3376 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5912_6
timestamp 1731220536
transform 1 0 3248 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5911_6
timestamp 1731220536
transform 1 0 3240 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5910_6
timestamp 1731220536
transform 1 0 3088 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5909_6
timestamp 1731220536
transform 1 0 2928 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5908_6
timestamp 1731220536
transform 1 0 3552 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5907_6
timestamp 1731220536
transform 1 0 3392 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5906_6
timestamp 1731220536
transform 1 0 3360 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5905_6
timestamp 1731220536
transform 1 0 3176 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5904_6
timestamp 1731220536
transform 1 0 2976 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5903_6
timestamp 1731220536
transform 1 0 3536 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5902_6
timestamp 1731220536
transform 1 0 3464 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5901_6
timestamp 1731220536
transform 1 0 3312 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5900_6
timestamp 1731220536
transform 1 0 3152 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5899_6
timestamp 1731220536
transform 1 0 2984 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5898_6
timestamp 1731220536
transform 1 0 3448 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5897_6
timestamp 1731220536
transform 1 0 3288 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5896_6
timestamp 1731220536
transform 1 0 3112 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5895_6
timestamp 1731220536
transform 1 0 2928 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5894_6
timestamp 1731220536
transform 1 0 2976 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5893_6
timestamp 1731220536
transform 1 0 3168 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5892_6
timestamp 1731220536
transform 1 0 3520 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5891_6
timestamp 1731220536
transform 1 0 3352 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5890_6
timestamp 1731220536
transform 1 0 3296 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5889_6
timestamp 1731220536
transform 1 0 3584 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5888_6
timestamp 1731220536
transform 1 0 3688 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5887_6
timestamp 1731220536
transform 1 0 3864 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5886_6
timestamp 1731220536
transform 1 0 3744 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5885_6
timestamp 1731220536
transform 1 0 3600 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5884_6
timestamp 1731220536
transform 1 0 3608 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5883_6
timestamp 1731220536
transform 1 0 3712 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5882_6
timestamp 1731220536
transform 1 0 3872 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5881_6
timestamp 1731220536
transform 1 0 3752 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5880_6
timestamp 1731220536
transform 1 0 3872 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5879_6
timestamp 1731220536
transform 1 0 3872 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5878_6
timestamp 1731220536
transform 1 0 3872 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5877_6
timestamp 1731220536
transform 1 0 3872 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5876_6
timestamp 1731220536
transform 1 0 3872 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5875_6
timestamp 1731220536
transform 1 0 3872 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5874_6
timestamp 1731220536
transform 1 0 3872 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5873_6
timestamp 1731220536
transform 1 0 3872 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5872_6
timestamp 1731220536
transform 1 0 3872 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5871_6
timestamp 1731220536
transform 1 0 3872 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5870_6
timestamp 1731220536
transform 1 0 3872 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5869_6
timestamp 1731220536
transform 1 0 3872 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5868_6
timestamp 1731220536
transform 1 0 3872 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5867_6
timestamp 1731220536
transform 1 0 3864 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5866_6
timestamp 1731220536
transform 1 0 3856 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5865_6
timestamp 1731220536
transform 1 0 3872 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5864_6
timestamp 1731220536
transform 1 0 3752 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5863_6
timestamp 1731220536
transform 1 0 3616 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5862_6
timestamp 1731220536
transform 1 0 3472 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5861_6
timestamp 1731220536
transform 1 0 3320 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5860_6
timestamp 1731220536
transform 1 0 3496 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5859_6
timestamp 1731220536
transform 1 0 3672 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5858_6
timestamp 1731220536
transform 1 0 3648 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5857_6
timestamp 1731220536
transform 1 0 3528 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5856_6
timestamp 1731220536
transform 1 0 3696 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5855_6
timestamp 1731220536
transform 1 0 3704 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5854_6
timestamp 1731220536
transform 1 0 3696 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5853_6
timestamp 1731220536
transform 1 0 3504 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5852_6
timestamp 1731220536
transform 1 0 3488 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5851_6
timestamp 1731220536
transform 1 0 3688 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5850_6
timestamp 1731220536
transform 1 0 3608 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5849_6
timestamp 1731220536
transform 1 0 3408 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5848_6
timestamp 1731220536
transform 1 0 3648 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5847_6
timestamp 1731220536
transform 1 0 3680 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5846_6
timestamp 1731220536
transform 1 0 3464 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5845_6
timestamp 1731220536
transform 1 0 3256 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5844_6
timestamp 1731220536
transform 1 0 3456 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5843_6
timestamp 1731220536
transform 1 0 3672 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5842_6
timestamp 1731220536
transform 1 0 3696 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5841_6
timestamp 1731220536
transform 1 0 3504 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5840_6
timestamp 1731220536
transform 1 0 3320 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5839_6
timestamp 1731220536
transform 1 0 3600 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5838_6
timestamp 1731220536
transform 1 0 3320 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5837_6
timestamp 1731220536
transform 1 0 3056 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5836_6
timestamp 1731220536
transform 1 0 3008 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5835_6
timestamp 1731220536
transform 1 0 2888 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5834_6
timestamp 1731220536
transform 1 0 3152 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5833_6
timestamp 1731220536
transform 1 0 3256 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5832_6
timestamp 1731220536
transform 1 0 3072 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5831_6
timestamp 1731220536
transform 1 0 2912 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5830_6
timestamp 1731220536
transform 1 0 2864 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5829_6
timestamp 1731220536
transform 1 0 3056 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5828_6
timestamp 1731220536
transform 1 0 2936 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5827_6
timestamp 1731220536
transform 1 0 2712 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5826_6
timestamp 1731220536
transform 1 0 3168 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5825_6
timestamp 1731220536
transform 1 0 3328 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5824_6
timestamp 1731220536
transform 1 0 3056 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5823_6
timestamp 1731220536
transform 1 0 2912 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5822_6
timestamp 1731220536
transform 1 0 3104 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5821_6
timestamp 1731220536
transform 1 0 3296 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5820_6
timestamp 1731220536
transform 1 0 3128 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5819_6
timestamp 1731220536
transform 1 0 2928 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5818_6
timestamp 1731220536
transform 1 0 3320 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5817_6
timestamp 1731220536
transform 1 0 3528 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5816_6
timestamp 1731220536
transform 1 0 3360 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5815_6
timestamp 1731220536
transform 1 0 3200 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5814_6
timestamp 1731220536
transform 1 0 3056 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5813_6
timestamp 1731220536
transform 1 0 3360 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5812_6
timestamp 1731220536
transform 1 0 3200 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5811_6
timestamp 1731220536
transform 1 0 3048 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5810_6
timestamp 1731220536
transform 1 0 3032 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5809_6
timestamp 1731220536
transform 1 0 2856 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5808_6
timestamp 1731220536
transform 1 0 3224 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5807_6
timestamp 1731220536
transform 1 0 3432 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5806_6
timestamp 1731220536
transform 1 0 3320 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5805_6
timestamp 1731220536
transform 1 0 3144 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5804_6
timestamp 1731220536
transform 1 0 2976 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5803_6
timestamp 1731220536
transform 1 0 2776 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5802_6
timestamp 1731220536
transform 1 0 2976 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5801_6
timestamp 1731220536
transform 1 0 3160 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5800_6
timestamp 1731220536
transform 1 0 3136 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5799_6
timestamp 1731220536
transform 1 0 2976 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5798_6
timestamp 1731220536
transform 1 0 3472 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5797_6
timestamp 1731220536
transform 1 0 3304 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5796_6
timestamp 1731220536
transform 1 0 3232 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5795_6
timestamp 1731220536
transform 1 0 3056 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5794_6
timestamp 1731220536
transform 1 0 3408 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5793_6
timestamp 1731220536
transform 1 0 3592 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5792_6
timestamp 1731220536
transform 1 0 3632 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5791_6
timestamp 1731220536
transform 1 0 3440 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5790_6
timestamp 1731220536
transform 1 0 3256 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5789_6
timestamp 1731220536
transform 1 0 3376 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5788_6
timestamp 1731220536
transform 1 0 3544 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5787_6
timestamp 1731220536
transform 1 0 3712 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5786_6
timestamp 1731220536
transform 1 0 3592 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5785_6
timestamp 1731220536
transform 1 0 3448 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5784_6
timestamp 1731220536
transform 1 0 3296 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5783_6
timestamp 1731220536
transform 1 0 3744 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5782_6
timestamp 1731220536
transform 1 0 3872 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5781_6
timestamp 1731220536
transform 1 0 3840 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5780_6
timestamp 1731220536
transform 1 0 3872 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5779_6
timestamp 1731220536
transform 1 0 3872 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5778_6
timestamp 1731220536
transform 1 0 3872 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5777_6
timestamp 1731220536
transform 1 0 3872 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5776_6
timestamp 1731220536
transform 1 0 3872 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5775_6
timestamp 1731220536
transform 1 0 3872 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5774_6
timestamp 1731220536
transform 1 0 3872 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5773_6
timestamp 1731220536
transform 1 0 3760 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5772_6
timestamp 1731220536
transform 1 0 3632 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5771_6
timestamp 1731220536
transform 1 0 3752 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5770_6
timestamp 1731220536
transform 1 0 3616 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5769_6
timestamp 1731220536
transform 1 0 3480 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5768_6
timestamp 1731220536
transform 1 0 3344 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5767_6
timestamp 1731220536
transform 1 0 3200 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5766_6
timestamp 1731220536
transform 1 0 3232 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5765_6
timestamp 1731220536
transform 1 0 3368 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5764_6
timestamp 1731220536
transform 1 0 3504 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5763_6
timestamp 1731220536
transform 1 0 3704 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5762_6
timestamp 1731220536
transform 1 0 3568 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5761_6
timestamp 1731220536
transform 1 0 3432 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5760_6
timestamp 1731220536
transform 1 0 3304 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5759_6
timestamp 1731220536
transform 1 0 3168 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5758_6
timestamp 1731220536
transform 1 0 3024 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5757_6
timestamp 1731220536
transform 1 0 2872 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5756_6
timestamp 1731220536
transform 1 0 2920 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5755_6
timestamp 1731220536
transform 1 0 3080 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5754_6
timestamp 1731220536
transform 1 0 3048 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5753_6
timestamp 1731220536
transform 1 0 3632 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5752_6
timestamp 1731220536
transform 1 0 3656 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5751_6
timestamp 1731220536
transform 1 0 3424 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5750_6
timestamp 1731220536
transform 1 0 3200 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5749_6
timestamp 1731220536
transform 1 0 3008 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5748_6
timestamp 1731220536
transform 1 0 2952 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5747_6
timestamp 1731220536
transform 1 0 2768 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5746_6
timestamp 1731220536
transform 1 0 3648 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5745_6
timestamp 1731220536
transform 1 0 3400 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5744_6
timestamp 1731220536
transform 1 0 3168 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5743_6
timestamp 1731220536
transform 1 0 3152 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5742_6
timestamp 1731220536
transform 1 0 2896 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5741_6
timestamp 1731220536
transform 1 0 2632 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5740_6
timestamp 1731220536
transform 1 0 3400 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5739_6
timestamp 1731220536
transform 1 0 3648 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5738_6
timestamp 1731220536
transform 1 0 3680 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5737_6
timestamp 1731220536
transform 1 0 3496 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5736_6
timestamp 1731220536
transform 1 0 3312 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5735_6
timestamp 1731220536
transform 1 0 3128 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5734_6
timestamp 1731220536
transform 1 0 2944 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5733_6
timestamp 1731220536
transform 1 0 3600 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5732_6
timestamp 1731220536
transform 1 0 3368 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5731_6
timestamp 1731220536
transform 1 0 3144 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5730_6
timestamp 1731220536
transform 1 0 2936 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5729_6
timestamp 1731220536
transform 1 0 3144 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5728_6
timestamp 1731220536
transform 1 0 3208 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5727_6
timestamp 1731220536
transform 1 0 3072 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5726_6
timestamp 1731220536
transform 1 0 2896 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5725_6
timestamp 1731220536
transform 1 0 2872 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5724_6
timestamp 1731220536
transform 1 0 2680 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5723_6
timestamp 1731220536
transform 1 0 2808 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5722_6
timestamp 1731220536
transform 1 0 2632 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5721_6
timestamp 1731220536
transform 1 0 2560 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5720_6
timestamp 1731220536
transform 1 0 2320 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5719_6
timestamp 1731220536
transform 1 0 2816 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5718_6
timestamp 1731220536
transform 1 0 2656 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5717_6
timestamp 1731220536
transform 1 0 2504 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5716_6
timestamp 1731220536
transform 1 0 2368 0 -1 1364
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5715_6
timestamp 1731220536
transform 1 0 2328 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5714_6
timestamp 1731220536
transform 1 0 2216 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5713_6
timestamp 1731220536
transform 1 0 2448 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5712_6
timestamp 1731220536
transform 1 0 2704 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5711_6
timestamp 1731220536
transform 1 0 2568 0 1 1372
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5710_6
timestamp 1731220536
transform 1 0 2464 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5709_6
timestamp 1731220536
transform 1 0 2568 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5708_6
timestamp 1731220536
transform 1 0 2672 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5707_6
timestamp 1731220536
transform 1 0 2784 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5706_6
timestamp 1731220536
transform 1 0 2912 0 -1 1520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5705_6
timestamp 1731220536
transform 1 0 2920 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5704_6
timestamp 1731220536
transform 1 0 2792 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5703_6
timestamp 1731220536
transform 1 0 2672 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5702_6
timestamp 1731220536
transform 1 0 2560 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5701_6
timestamp 1731220536
transform 1 0 2456 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5700_6
timestamp 1731220536
transform 1 0 2288 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5699_6
timestamp 1731220536
transform 1 0 2504 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5698_6
timestamp 1731220536
transform 1 0 2720 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5697_6
timestamp 1731220536
transform 1 0 2728 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5696_6
timestamp 1731220536
transform 1 0 2552 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5695_6
timestamp 1731220536
transform 1 0 2208 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5694_6
timestamp 1731220536
transform 1 0 2088 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5693_6
timestamp 1731220536
transform 1 0 2088 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5692_6
timestamp 1731220536
transform 1 0 1912 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5691_6
timestamp 1731220536
transform 1 0 1768 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5690_6
timestamp 1731220536
transform 1 0 1608 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5689_6
timestamp 1731220536
transform 1 0 1448 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5688_6
timestamp 1731220536
transform 1 0 1280 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5687_6
timestamp 1731220536
transform 1 0 1912 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5686_6
timestamp 1731220536
transform 1 0 1912 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5685_6
timestamp 1731220536
transform 1 0 1760 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5684_6
timestamp 1731220536
transform 1 0 1592 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5683_6
timestamp 1731220536
transform 1 0 1424 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5682_6
timestamp 1731220536
transform 1 0 1240 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5681_6
timestamp 1731220536
transform 1 0 1760 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5680_6
timestamp 1731220536
transform 1 0 1592 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5679_6
timestamp 1731220536
transform 1 0 1424 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5678_6
timestamp 1731220536
transform 1 0 1256 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5677_6
timestamp 1731220536
transform 1 0 1088 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5676_6
timestamp 1731220536
transform 1 0 1448 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5675_6
timestamp 1731220536
transform 1 0 1312 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5674_6
timestamp 1731220536
transform 1 0 1176 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5673_6
timestamp 1731220536
transform 1 0 1048 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5672_6
timestamp 1731220536
transform 1 0 912 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5671_6
timestamp 1731220536
transform 1 0 896 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5670_6
timestamp 1731220536
transform 1 0 784 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5669_6
timestamp 1731220536
transform 1 0 1248 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5668_6
timestamp 1731220536
transform 1 0 1128 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5667_6
timestamp 1731220536
transform 1 0 1008 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5666_6
timestamp 1731220536
transform 1 0 944 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5665_6
timestamp 1731220536
transform 1 0 1096 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5664_6
timestamp 1731220536
transform 1 0 1240 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5663_6
timestamp 1731220536
transform 1 0 1544 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5662_6
timestamp 1731220536
transform 1 0 1392 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5661_6
timestamp 1731220536
transform 1 0 1344 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5660_6
timestamp 1731220536
transform 1 0 1168 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5659_6
timestamp 1731220536
transform 1 0 1512 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5658_6
timestamp 1731220536
transform 1 0 1680 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5657_6
timestamp 1731220536
transform 1 0 1848 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5656_6
timestamp 1731220536
transform 1 0 1912 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5655_6
timestamp 1731220536
transform 1 0 1760 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5654_6
timestamp 1731220536
transform 1 0 1584 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5653_6
timestamp 1731220536
transform 1 0 1408 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5652_6
timestamp 1731220536
transform 1 0 1232 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5651_6
timestamp 1731220536
transform 1 0 1688 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5650_6
timestamp 1731220536
transform 1 0 1528 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5649_6
timestamp 1731220536
transform 1 0 1368 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5648_6
timestamp 1731220536
transform 1 0 1208 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5647_6
timestamp 1731220536
transform 1 0 1040 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5646_6
timestamp 1731220536
transform 1 0 1400 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5645_6
timestamp 1731220536
transform 1 0 1272 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5644_6
timestamp 1731220536
transform 1 0 1144 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5643_6
timestamp 1731220536
transform 1 0 1016 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5642_6
timestamp 1731220536
transform 1 0 880 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5641_6
timestamp 1731220536
transform 1 0 1136 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5640_6
timestamp 1731220536
transform 1 0 1392 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5639_6
timestamp 1731220536
transform 1 0 1264 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5638_6
timestamp 1731220536
transform 1 0 1248 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5637_6
timestamp 1731220536
transform 1 0 1400 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5636_6
timestamp 1731220536
transform 1 0 1552 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5635_6
timestamp 1731220536
transform 1 0 1664 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5634_6
timestamp 1731220536
transform 1 0 1512 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5633_6
timestamp 1731220536
transform 1 0 1536 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5632_6
timestamp 1731220536
transform 1 0 1704 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5631_6
timestamp 1731220536
transform 1 0 1880 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5630_6
timestamp 1731220536
transform 1 0 1896 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5629_6
timestamp 1731220536
transform 1 0 1680 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5628_6
timestamp 1731220536
transform 1 0 1784 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5627_6
timestamp 1731220536
transform 1 0 1592 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5626_6
timestamp 1731220536
transform 1 0 1408 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5625_6
timestamp 1731220536
transform 1 0 1632 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5624_6
timestamp 1731220536
transform 1 0 1464 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5623_6
timestamp 1731220536
transform 1 0 1440 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5622_6
timestamp 1731220536
transform 1 0 1296 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5621_6
timestamp 1731220536
transform 1 0 1136 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5620_6
timestamp 1731220536
transform 1 0 968 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5619_6
timestamp 1731220536
transform 1 0 1032 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5618_6
timestamp 1731220536
transform 1 0 1224 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5617_6
timestamp 1731220536
transform 1 0 1472 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5616_6
timestamp 1731220536
transform 1 0 1272 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5615_6
timestamp 1731220536
transform 1 0 1072 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5614_6
timestamp 1731220536
transform 1 0 1208 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5613_6
timestamp 1731220536
transform 1 0 1368 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5612_6
timestamp 1731220536
transform 1 0 1368 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5611_6
timestamp 1731220536
transform 1 0 1232 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5610_6
timestamp 1731220536
transform 1 0 1096 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5609_6
timestamp 1731220536
transform 1 0 1096 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5608_6
timestamp 1731220536
transform 1 0 952 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5607_6
timestamp 1731220536
transform 1 0 1008 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5606_6
timestamp 1731220536
transform 1 0 880 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5605_6
timestamp 1731220536
transform 1 0 744 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5604_6
timestamp 1731220536
transform 1 0 600 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5603_6
timestamp 1731220536
transform 1 0 600 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5602_6
timestamp 1731220536
transform 1 0 448 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5601_6
timestamp 1731220536
transform 1 0 744 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5600_6
timestamp 1731220536
transform 1 0 864 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5599_6
timestamp 1731220536
transform 1 0 680 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5598_6
timestamp 1731220536
transform 1 0 640 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5597_6
timestamp 1731220536
transform 1 0 840 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5596_6
timestamp 1731220536
transform 1 0 1040 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5595_6
timestamp 1731220536
transform 1 0 992 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5594_6
timestamp 1731220536
transform 1 0 808 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5593_6
timestamp 1731220536
transform 1 0 624 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5592_6
timestamp 1731220536
transform 1 0 448 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5591_6
timestamp 1731220536
transform 1 0 288 0 -1 2484
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5590_6
timestamp 1731220536
transform 1 0 256 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5589_6
timestamp 1731220536
transform 1 0 440 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5588_6
timestamp 1731220536
transform 1 0 488 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5587_6
timestamp 1731220536
transform 1 0 296 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5586_6
timestamp 1731220536
transform 1 0 128 0 -1 2660
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5585_6
timestamp 1731220536
transform 1 0 128 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5584_6
timestamp 1731220536
transform 1 0 280 0 1 2672
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5583_6
timestamp 1731220536
transform 1 0 128 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5582_6
timestamp 1731220536
transform 1 0 448 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5581_6
timestamp 1731220536
transform 1 0 288 0 -1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5580_6
timestamp 1731220536
transform 1 0 288 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5579_6
timestamp 1731220536
transform 1 0 408 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5578_6
timestamp 1731220536
transform 1 0 536 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5577_6
timestamp 1731220536
transform 1 0 808 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5576_6
timestamp 1731220536
transform 1 0 672 0 1 2848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5575_6
timestamp 1731220536
transform 1 0 632 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5574_6
timestamp 1731220536
transform 1 0 528 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5573_6
timestamp 1731220536
transform 1 0 736 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5572_6
timestamp 1731220536
transform 1 0 848 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5571_6
timestamp 1731220536
transform 1 0 968 0 -1 3004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5570_6
timestamp 1731220536
transform 1 0 1056 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5569_6
timestamp 1731220536
transform 1 0 912 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5568_6
timestamp 1731220536
transform 1 0 776 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5567_6
timestamp 1731220536
transform 1 0 656 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5566_6
timestamp 1731220536
transform 1 0 552 0 1 3016
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5565_6
timestamp 1731220536
transform 1 0 880 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5564_6
timestamp 1731220536
transform 1 0 704 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5563_6
timestamp 1731220536
transform 1 0 544 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5562_6
timestamp 1731220536
transform 1 0 400 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5561_6
timestamp 1731220536
transform 1 0 264 0 -1 3176
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5560_6
timestamp 1731220536
transform 1 0 840 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5559_6
timestamp 1731220536
transform 1 0 648 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5558_6
timestamp 1731220536
transform 1 0 456 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5557_6
timestamp 1731220536
transform 1 0 272 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5556_6
timestamp 1731220536
transform 1 0 128 0 1 3188
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5555_6
timestamp 1731220536
transform 1 0 792 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5554_6
timestamp 1731220536
transform 1 0 616 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5553_6
timestamp 1731220536
transform 1 0 440 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5552_6
timestamp 1731220536
transform 1 0 264 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5551_6
timestamp 1731220536
transform 1 0 128 0 -1 3344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5550_6
timestamp 1731220536
transform 1 0 128 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5549_6
timestamp 1731220536
transform 1 0 312 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5548_6
timestamp 1731220536
transform 1 0 1136 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5547_6
timestamp 1731220536
transform 1 0 840 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5546_6
timestamp 1731220536
transform 1 0 560 0 1 3352
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5545_6
timestamp 1731220536
transform 1 0 352 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5544_6
timestamp 1731220536
transform 1 0 128 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5543_6
timestamp 1731220536
transform 1 0 592 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5542_6
timestamp 1731220536
transform 1 0 824 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5541_6
timestamp 1731220536
transform 1 0 680 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5540_6
timestamp 1731220536
transform 1 0 528 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5539_6
timestamp 1731220536
transform 1 0 376 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5538_6
timestamp 1731220536
transform 1 0 216 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5537_6
timestamp 1731220536
transform 1 0 320 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5536_6
timestamp 1731220536
transform 1 0 840 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5535_6
timestamp 1731220536
transform 1 0 672 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5534_6
timestamp 1731220536
transform 1 0 496 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5533_6
timestamp 1731220536
transform 1 0 472 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5532_6
timestamp 1731220536
transform 1 0 336 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5531_6
timestamp 1731220536
transform 1 0 608 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5530_6
timestamp 1731220536
transform 1 0 752 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5529_6
timestamp 1731220536
transform 1 0 896 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5528_6
timestamp 1731220536
transform 1 0 840 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5527_6
timestamp 1731220536
transform 1 0 696 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5526_6
timestamp 1731220536
transform 1 0 552 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5525_6
timestamp 1731220536
transform 1 0 408 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5524_6
timestamp 1731220536
transform 1 0 352 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5523_6
timestamp 1731220536
transform 1 0 472 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5522_6
timestamp 1731220536
transform 1 0 872 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5521_6
timestamp 1731220536
transform 1 0 736 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5520_6
timestamp 1731220536
transform 1 0 600 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5519_6
timestamp 1731220536
transform 1 0 576 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5518_6
timestamp 1731220536
transform 1 0 472 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5517_6
timestamp 1731220536
transform 1 0 368 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5516_6
timestamp 1731220536
transform 1 0 888 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5515_6
timestamp 1731220536
transform 1 0 784 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5514_6
timestamp 1731220536
transform 1 0 680 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5513_6
timestamp 1731220536
transform 1 0 576 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5512_6
timestamp 1731220536
transform 1 0 472 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5511_6
timestamp 1731220536
transform 1 0 680 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5510_6
timestamp 1731220536
transform 1 0 784 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5509_6
timestamp 1731220536
transform 1 0 888 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5508_6
timestamp 1731220536
transform 1 0 992 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5507_6
timestamp 1731220536
transform 1 0 1096 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5506_6
timestamp 1731220536
transform 1 0 1200 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5505_6
timestamp 1731220536
transform 1 0 1408 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5504_6
timestamp 1731220536
transform 1 0 1304 0 1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5503_6
timestamp 1731220536
transform 1 0 1200 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5502_6
timestamp 1731220536
transform 1 0 1096 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5501_6
timestamp 1731220536
transform 1 0 992 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5500_6
timestamp 1731220536
transform 1 0 1304 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5499_6
timestamp 1731220536
transform 1 0 1408 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5498_6
timestamp 1731220536
transform 1 0 1512 0 -1 3972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5497_6
timestamp 1731220536
transform 1 0 1528 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5496_6
timestamp 1731220536
transform 1 0 1392 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5495_6
timestamp 1731220536
transform 1 0 1256 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5494_6
timestamp 1731220536
transform 1 0 1128 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5493_6
timestamp 1731220536
transform 1 0 1000 0 1 3824
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5492_6
timestamp 1731220536
transform 1 0 976 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5491_6
timestamp 1731220536
transform 1 0 1112 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5490_6
timestamp 1731220536
transform 1 0 1248 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5489_6
timestamp 1731220536
transform 1 0 1384 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5488_6
timestamp 1731220536
transform 1 0 1528 0 -1 3816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5487_6
timestamp 1731220536
transform 1 0 1504 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5486_6
timestamp 1731220536
transform 1 0 1352 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5485_6
timestamp 1731220536
transform 1 0 1200 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5484_6
timestamp 1731220536
transform 1 0 1048 0 1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5483_6
timestamp 1731220536
transform 1 0 1008 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5482_6
timestamp 1731220536
transform 1 0 1168 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5481_6
timestamp 1731220536
transform 1 0 1632 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5480_6
timestamp 1731220536
transform 1 0 1472 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5479_6
timestamp 1731220536
transform 1 0 1320 0 -1 3664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5478_6
timestamp 1731220536
transform 1 0 1112 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5477_6
timestamp 1731220536
transform 1 0 976 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5476_6
timestamp 1731220536
transform 1 0 832 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5475_6
timestamp 1731220536
transform 1 0 1472 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5474_6
timestamp 1731220536
transform 1 0 1360 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5473_6
timestamp 1731220536
transform 1 0 1240 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5472_6
timestamp 1731220536
transform 1 0 1232 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5471_6
timestamp 1731220536
transform 1 0 1040 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5470_6
timestamp 1731220536
transform 1 0 1416 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5469_6
timestamp 1731220536
transform 1 0 1912 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5468_6
timestamp 1731220536
transform 1 0 1760 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5467_6
timestamp 1731220536
transform 1 0 1592 0 -1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5466_6
timestamp 1731220536
transform 1 0 1584 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5465_6
timestamp 1731220536
transform 1 0 1696 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5464_6
timestamp 1731220536
transform 1 0 1808 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5463_6
timestamp 1731220536
transform 1 0 1912 0 1 3520
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5462_6
timestamp 1731220536
transform 1 0 2088 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5461_6
timestamp 1731220536
transform 1 0 2272 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5460_6
timestamp 1731220536
transform 1 0 2272 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5459_6
timestamp 1731220536
transform 1 0 2088 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5458_6
timestamp 1731220536
transform 1 0 2088 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5457_6
timestamp 1731220536
transform 1 0 2216 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5456_6
timestamp 1731220536
transform 1 0 2368 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5455_6
timestamp 1731220536
transform 1 0 2264 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5454_6
timestamp 1731220536
transform 1 0 2096 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5453_6
timestamp 1731220536
transform 1 0 2296 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5452_6
timestamp 1731220536
transform 1 0 2120 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5451_6
timestamp 1731220536
transform 1 0 2088 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5450_6
timestamp 1731220536
transform 1 0 2192 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5449_6
timestamp 1731220536
transform 1 0 2296 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5448_6
timestamp 1731220536
transform 1 0 2400 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5447_6
timestamp 1731220536
transform 1 0 2504 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5446_6
timestamp 1731220536
transform 1 0 2624 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5445_6
timestamp 1731220536
transform 1 0 2880 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5444_6
timestamp 1731220536
transform 1 0 2752 0 -1 4008
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5443_6
timestamp 1731220536
transform 1 0 2624 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5442_6
timestamp 1731220536
transform 1 0 2464 0 1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5441_6
timestamp 1731220536
transform 1 0 2424 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5440_6
timestamp 1731220536
transform 1 0 2576 0 -1 3860
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5439_6
timestamp 1731220536
transform 1 0 2520 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5438_6
timestamp 1731220536
transform 1 0 2664 0 1 3712
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5437_6
timestamp 1731220536
transform 1 0 2648 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5436_6
timestamp 1731220536
transform 1 0 2464 0 -1 3704
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5435_6
timestamp 1731220536
transform 1 0 2472 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5434_6
timestamp 1731220536
transform 1 0 2664 0 1 3552
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5433_6
timestamp 1731220536
transform 1 0 2704 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5432_6
timestamp 1731220536
transform 1 0 2568 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5431_6
timestamp 1731220536
transform 1 0 2424 0 -1 3540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5430_6
timestamp 1731220536
transform 1 0 2320 0 1 3396
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5429_6
timestamp 1731220536
transform 1 0 2832 0 1 3396
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5428_6
timestamp 1731220536
transform 1 0 3352 0 1 3396
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5427_6
timestamp 1731220536
transform 1 0 3424 0 -1 3392
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5426_6
timestamp 1731220536
transform 1 0 2984 0 -1 3392
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5425_6
timestamp 1731220536
transform 1 0 2560 0 -1 3392
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5424_6
timestamp 1731220536
transform 1 0 2160 0 -1 3392
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5423_6
timestamp 1731220536
transform 1 0 2680 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5422_6
timestamp 1731220536
transform 1 0 2480 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5421_6
timestamp 1731220536
transform 1 0 2272 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5420_6
timestamp 1731220536
transform 1 0 2088 0 1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5419_6
timestamp 1731220536
transform 1 0 2088 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5418_6
timestamp 1731220536
transform 1 0 2216 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5417_6
timestamp 1731220536
transform 1 0 2376 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5416_6
timestamp 1731220536
transform 1 0 2536 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5415_6
timestamp 1731220536
transform 1 0 2696 0 -1 3232
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5414_6
timestamp 1731220536
transform 1 0 2712 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5413_6
timestamp 1731220536
transform 1 0 2528 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5412_6
timestamp 1731220536
transform 1 0 2344 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5411_6
timestamp 1731220536
transform 1 0 2160 0 1 3072
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5410_6
timestamp 1731220536
transform 1 0 2328 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5409_6
timestamp 1731220536
transform 1 0 2432 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5408_6
timestamp 1731220536
transform 1 0 2544 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5407_6
timestamp 1731220536
transform 1 0 2664 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5406_6
timestamp 1731220536
transform 1 0 2784 0 -1 3064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5405_6
timestamp 1731220536
transform 1 0 2680 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5404_6
timestamp 1731220536
transform 1 0 2576 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5403_6
timestamp 1731220536
transform 1 0 2472 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5402_6
timestamp 1731220536
transform 1 0 2784 0 1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5401_6
timestamp 1731220536
transform 1 0 2808 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5400_6
timestamp 1731220536
transform 1 0 2704 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5399_6
timestamp 1731220536
transform 1 0 2600 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5398_6
timestamp 1731220536
transform 1 0 2496 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5397_6
timestamp 1731220536
transform 1 0 2392 0 -1 2920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5396_6
timestamp 1731220536
transform 1 0 2800 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5395_6
timestamp 1731220536
transform 1 0 2696 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5394_6
timestamp 1731220536
transform 1 0 2592 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5393_6
timestamp 1731220536
transform 1 0 2488 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5392_6
timestamp 1731220536
transform 1 0 2384 0 1 2772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5391_6
timestamp 1731220536
transform 1 0 2752 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5390_6
timestamp 1731220536
transform 1 0 2632 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5389_6
timestamp 1731220536
transform 1 0 2512 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5388_6
timestamp 1731220536
transform 1 0 2392 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5387_6
timestamp 1731220536
transform 1 0 2280 0 -1 2764
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5386_6
timestamp 1731220536
transform 1 0 2768 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5385_6
timestamp 1731220536
transform 1 0 2600 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5384_6
timestamp 1731220536
transform 1 0 2440 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5383_6
timestamp 1731220536
transform 1 0 2280 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5382_6
timestamp 1731220536
transform 1 0 2128 0 1 2604
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5381_6
timestamp 1731220536
transform 1 0 2760 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5380_6
timestamp 1731220536
transform 1 0 2536 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5379_6
timestamp 1731220536
transform 1 0 2304 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5378_6
timestamp 1731220536
transform 1 0 2088 0 -1 2596
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5377_6
timestamp 1731220536
transform 1 0 2800 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5376_6
timestamp 1731220536
transform 1 0 2608 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5375_6
timestamp 1731220536
transform 1 0 2416 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5374_6
timestamp 1731220536
transform 1 0 2232 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5373_6
timestamp 1731220536
transform 1 0 2088 0 1 2452
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5372_6
timestamp 1731220536
transform 1 0 2088 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5371_6
timestamp 1731220536
transform 1 0 2288 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5370_6
timestamp 1731220536
transform 1 0 2512 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5369_6
timestamp 1731220536
transform 1 0 2728 0 -1 2444
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5368_6
timestamp 1731220536
transform 1 0 2760 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5367_6
timestamp 1731220536
transform 1 0 2536 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5366_6
timestamp 1731220536
transform 1 0 2304 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5365_6
timestamp 1731220536
transform 1 0 2088 0 1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5364_6
timestamp 1731220536
transform 1 0 2088 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5363_6
timestamp 1731220536
transform 1 0 2272 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5362_6
timestamp 1731220536
transform 1 0 2504 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5361_6
timestamp 1731220536
transform 1 0 2752 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5360_6
timestamp 1731220536
transform 1 0 3016 0 -1 2300
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5359_6
timestamp 1731220536
transform 1 0 2816 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5358_6
timestamp 1731220536
transform 1 0 2600 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5357_6
timestamp 1731220536
transform 1 0 2416 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5356_6
timestamp 1731220536
transform 1 0 2256 0 1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5355_6
timestamp 1731220536
transform 1 0 2368 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5354_6
timestamp 1731220536
transform 1 0 2472 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5353_6
timestamp 1731220536
transform 1 0 2576 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5352_6
timestamp 1731220536
transform 1 0 2680 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5351_6
timestamp 1731220536
transform 1 0 2784 0 -1 2148
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5350_6
timestamp 1731220536
transform 1 0 2784 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5349_6
timestamp 1731220536
transform 1 0 2672 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5348_6
timestamp 1731220536
transform 1 0 2568 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5347_6
timestamp 1731220536
transform 1 0 2464 0 1 2000
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5346_6
timestamp 1731220536
transform 1 0 2680 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5345_6
timestamp 1731220536
transform 1 0 2504 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5344_6
timestamp 1731220536
transform 1 0 2496 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5343_6
timestamp 1731220536
transform 1 0 2280 0 1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5342_6
timestamp 1731220536
transform 1 0 2376 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5341_6
timestamp 1731220536
transform 1 0 2808 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5340_6
timestamp 1731220536
transform 1 0 2576 0 -1 1844
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5339_6
timestamp 1731220536
transform 1 0 2376 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5338_6
timestamp 1731220536
transform 1 0 2216 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5337_6
timestamp 1731220536
transform 1 0 2088 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5336_6
timestamp 1731220536
transform 1 0 2088 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5335_6
timestamp 1731220536
transform 1 0 1912 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5334_6
timestamp 1731220536
transform 1 0 1736 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5333_6
timestamp 1731220536
transform 1 0 1784 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5332_6
timestamp 1731220536
transform 1 0 1536 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5331_6
timestamp 1731220536
transform 1 0 1344 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5330_6
timestamp 1731220536
transform 1 0 1768 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5329_6
timestamp 1731220536
transform 1 0 1592 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5328_6
timestamp 1731220536
transform 1 0 1416 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5327_6
timestamp 1731220536
transform 1 0 1240 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5326_6
timestamp 1731220536
transform 1 0 1296 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5325_6
timestamp 1731220536
transform 1 0 1600 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5324_6
timestamp 1731220536
transform 1 0 1448 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5323_6
timestamp 1731220536
transform 1 0 1400 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5322_6
timestamp 1731220536
transform 1 0 1568 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5321_6
timestamp 1731220536
transform 1 0 1744 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5320_6
timestamp 1731220536
transform 1 0 1824 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5319_6
timestamp 1731220536
transform 1 0 1608 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5318_6
timestamp 1731220536
transform 1 0 1400 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5317_6
timestamp 1731220536
transform 1 0 1232 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5316_6
timestamp 1731220536
transform 1 0 1408 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5315_6
timestamp 1731220536
transform 1 0 1584 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5314_6
timestamp 1731220536
transform 1 0 1760 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5313_6
timestamp 1731220536
transform 1 0 1912 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5312_6
timestamp 1731220536
transform 1 0 1912 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5311_6
timestamp 1731220536
transform 1 0 2088 0 1 1212
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5310_6
timestamp 1731220536
transform 1 0 2088 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5309_6
timestamp 1731220536
transform 1 0 2256 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5308_6
timestamp 1731220536
transform 1 0 2448 0 -1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5307_6
timestamp 1731220536
transform 1 0 2480 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5306_6
timestamp 1731220536
transform 1 0 2272 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5305_6
timestamp 1731220536
transform 1 0 2088 0 1 1060
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5304_6
timestamp 1731220536
transform 1 0 2144 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5303_6
timestamp 1731220536
transform 1 0 2264 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5302_6
timestamp 1731220536
transform 1 0 2400 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5301_6
timestamp 1731220536
transform 1 0 2552 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5300_6
timestamp 1731220536
transform 1 0 2720 0 -1 1052
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5299_6
timestamp 1731220536
transform 1 0 2624 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5298_6
timestamp 1731220536
transform 1 0 2504 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5297_6
timestamp 1731220536
transform 1 0 2752 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5296_6
timestamp 1731220536
transform 1 0 2896 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5295_6
timestamp 1731220536
transform 1 0 3048 0 1 900
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5294_6
timestamp 1731220536
transform 1 0 2992 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5293_6
timestamp 1731220536
transform 1 0 2840 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5292_6
timestamp 1731220536
transform 1 0 2688 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5291_6
timestamp 1731220536
transform 1 0 2552 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5290_6
timestamp 1731220536
transform 1 0 2432 0 -1 888
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5289_6
timestamp 1731220536
transform 1 0 2760 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5288_6
timestamp 1731220536
transform 1 0 2600 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5287_6
timestamp 1731220536
transform 1 0 2456 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5286_6
timestamp 1731220536
transform 1 0 2320 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5285_6
timestamp 1731220536
transform 1 0 2192 0 1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5284_6
timestamp 1731220536
transform 1 0 2760 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5283_6
timestamp 1731220536
transform 1 0 2576 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5282_6
timestamp 1731220536
transform 1 0 2400 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5281_6
timestamp 1731220536
transform 1 0 2224 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5280_6
timestamp 1731220536
transform 1 0 2088 0 -1 736
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5279_6
timestamp 1731220536
transform 1 0 2088 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5278_6
timestamp 1731220536
transform 1 0 1912 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5277_6
timestamp 1731220536
transform 1 0 1768 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5276_6
timestamp 1731220536
transform 1 0 1600 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5275_6
timestamp 1731220536
transform 1 0 2352 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5274_6
timestamp 1731220536
transform 1 0 2328 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5273_6
timestamp 1731220536
transform 1 0 2192 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5272_6
timestamp 1731220536
transform 1 0 2088 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5271_6
timestamp 1731220536
transform 1 0 2464 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5270_6
timestamp 1731220536
transform 1 0 2608 0 -1 576
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5269_6
timestamp 1731220536
transform 1 0 2504 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5268_6
timestamp 1731220536
transform 1 0 2400 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5267_6
timestamp 1731220536
transform 1 0 2608 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5266_6
timestamp 1731220536
transform 1 0 2720 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5265_6
timestamp 1731220536
transform 1 0 2848 0 1 428
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5264_6
timestamp 1731220536
transform 1 0 3376 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5263_6
timestamp 1731220536
transform 1 0 3136 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5262_6
timestamp 1731220536
transform 1 0 2928 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5261_6
timestamp 1731220536
transform 1 0 2752 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5260_6
timestamp 1731220536
transform 1 0 2616 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5259_6
timestamp 1731220536
transform 1 0 2504 0 -1 424
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5258_6
timestamp 1731220536
transform 1 0 2888 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5257_6
timestamp 1731220536
transform 1 0 2720 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5256_6
timestamp 1731220536
transform 1 0 2560 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5255_6
timestamp 1731220536
transform 1 0 2400 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5254_6
timestamp 1731220536
transform 1 0 2248 0 1 268
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5253_6
timestamp 1731220536
transform 1 0 2752 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5252_6
timestamp 1731220536
transform 1 0 2576 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5251_6
timestamp 1731220536
transform 1 0 2400 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5250_6
timestamp 1731220536
transform 1 0 2224 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5249_6
timestamp 1731220536
transform 1 0 2088 0 -1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5248_6
timestamp 1731220536
transform 1 0 2712 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5247_6
timestamp 1731220536
transform 1 0 2544 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5246_6
timestamp 1731220536
transform 1 0 2376 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5245_6
timestamp 1731220536
transform 1 0 2216 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5244_6
timestamp 1731220536
transform 1 0 2088 0 1 104
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5243_6
timestamp 1731220536
transform 1 0 1912 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5242_6
timestamp 1731220536
transform 1 0 1808 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5241_6
timestamp 1731220536
transform 1 0 1704 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5240_6
timestamp 1731220536
transform 1 0 1600 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5239_6
timestamp 1731220536
transform 1 0 1488 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5238_6
timestamp 1731220536
transform 1 0 1376 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5237_6
timestamp 1731220536
transform 1 0 1272 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5236_6
timestamp 1731220536
transform 1 0 1168 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5235_6
timestamp 1731220536
transform 1 0 1064 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5234_6
timestamp 1731220536
transform 1 0 960 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5233_6
timestamp 1731220536
transform 1 0 1792 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5232_6
timestamp 1731220536
transform 1 0 1608 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5231_6
timestamp 1731220536
transform 1 0 1424 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5230_6
timestamp 1731220536
transform 1 0 1240 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5229_6
timestamp 1731220536
transform 1 0 1048 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5228_6
timestamp 1731220536
transform 1 0 1600 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5227_6
timestamp 1731220536
transform 1 0 1440 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5226_6
timestamp 1731220536
transform 1 0 1280 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5225_6
timestamp 1731220536
transform 1 0 1120 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5224_6
timestamp 1731220536
transform 1 0 1536 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5223_6
timestamp 1731220536
transform 1 0 1432 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5222_6
timestamp 1731220536
transform 1 0 1328 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5221_6
timestamp 1731220536
transform 1 0 1224 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5220_6
timestamp 1731220536
transform 1 0 1120 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5219_6
timestamp 1731220536
transform 1 0 1352 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5218_6
timestamp 1731220536
transform 1 0 1248 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5217_6
timestamp 1731220536
transform 1 0 1144 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5216_6
timestamp 1731220536
transform 1 0 1040 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5215_6
timestamp 1731220536
transform 1 0 936 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5214_6
timestamp 1731220536
transform 1 0 1248 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5213_6
timestamp 1731220536
transform 1 0 1128 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5212_6
timestamp 1731220536
transform 1 0 1008 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5211_6
timestamp 1731220536
transform 1 0 888 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5210_6
timestamp 1731220536
transform 1 0 776 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5209_6
timestamp 1731220536
transform 1 0 664 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5208_6
timestamp 1731220536
transform 1 0 784 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5207_6
timestamp 1731220536
transform 1 0 936 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5206_6
timestamp 1731220536
transform 1 0 1432 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5205_6
timestamp 1731220536
transform 1 0 1264 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5204_6
timestamp 1731220536
transform 1 0 1096 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5203_6
timestamp 1731220536
transform 1 0 1016 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5202_6
timestamp 1731220536
transform 1 0 864 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5201_6
timestamp 1731220536
transform 1 0 1168 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5200_6
timestamp 1731220536
transform 1 0 1472 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5199_6
timestamp 1731220536
transform 1 0 1320 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5198_6
timestamp 1731220536
transform 1 0 1232 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5197_6
timestamp 1731220536
transform 1 0 1064 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5196_6
timestamp 1731220536
transform 1 0 1568 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5195_6
timestamp 1731220536
transform 1 0 1400 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5194_6
timestamp 1731220536
transform 1 0 1328 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5193_6
timestamp 1731220536
transform 1 0 1176 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5192_6
timestamp 1731220536
transform 1 0 1472 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5191_6
timestamp 1731220536
transform 1 0 1624 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5190_6
timestamp 1731220536
transform 1 0 1776 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5189_6
timestamp 1731220536
transform 1 0 1912 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5188_6
timestamp 1731220536
transform 1 0 1784 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5187_6
timestamp 1731220536
transform 1 0 1632 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5186_6
timestamp 1731220536
transform 1 0 1480 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5185_6
timestamp 1731220536
transform 1 0 1328 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5184_6
timestamp 1731220536
transform 1 0 1840 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5183_6
timestamp 1731220536
transform 1 0 1712 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5182_6
timestamp 1731220536
transform 1 0 1584 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5181_6
timestamp 1731220536
transform 1 0 1456 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5180_6
timestamp 1731220536
transform 1 0 1328 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5179_6
timestamp 1731220536
transform 1 0 1680 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5178_6
timestamp 1731220536
transform 1 0 1552 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5177_6
timestamp 1731220536
transform 1 0 1432 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5176_6
timestamp 1731220536
transform 1 0 1312 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5175_6
timestamp 1731220536
transform 1 0 1192 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5174_6
timestamp 1731220536
transform 1 0 1520 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5173_6
timestamp 1731220536
transform 1 0 1400 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5172_6
timestamp 1731220536
transform 1 0 1280 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5171_6
timestamp 1731220536
transform 1 0 1160 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5170_6
timestamp 1731220536
transform 1 0 1040 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5169_6
timestamp 1731220536
transform 1 0 1696 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5168_6
timestamp 1731220536
transform 1 0 1464 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5167_6
timestamp 1731220536
transform 1 0 1240 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5166_6
timestamp 1731220536
transform 1 0 1032 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5165_6
timestamp 1731220536
transform 1 0 856 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5164_6
timestamp 1731220536
transform 1 0 1040 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5163_6
timestamp 1731220536
transform 1 0 984 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5162_6
timestamp 1731220536
transform 1 0 1192 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5161_6
timestamp 1731220536
transform 1 0 1232 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5160_6
timestamp 1731220536
transform 1 0 1064 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5159_6
timestamp 1731220536
transform 1 0 1008 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5158_6
timestamp 1731220536
transform 1 0 1152 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5157_6
timestamp 1731220536
transform 1 0 1056 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5156_6
timestamp 1731220536
transform 1 0 1144 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5155_6
timestamp 1731220536
transform 1 0 1600 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5154_6
timestamp 1731220536
transform 1 0 1424 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5153_6
timestamp 1731220536
transform 1 0 1248 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5152_6
timestamp 1731220536
transform 1 0 1072 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5151_6
timestamp 1731220536
transform 1 0 1712 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5150_6
timestamp 1731220536
transform 1 0 1488 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5149_6
timestamp 1731220536
transform 1 0 1272 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5148_6
timestamp 1731220536
transform 1 0 1080 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5147_6
timestamp 1731220536
transform 1 0 904 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5146_6
timestamp 1731220536
transform 1 0 912 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5145_6
timestamp 1731220536
transform 1 0 744 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5144_6
timestamp 1731220536
transform 1 0 592 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5143_6
timestamp 1731220536
transform 1 0 896 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5142_6
timestamp 1731220536
transform 1 0 712 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5141_6
timestamp 1731220536
transform 1 0 520 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5140_6
timestamp 1731220536
transform 1 0 320 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5139_6
timestamp 1731220536
transform 1 0 280 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5138_6
timestamp 1731220536
transform 1 0 440 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5137_6
timestamp 1731220536
transform 1 0 512 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5136_6
timestamp 1731220536
transform 1 0 712 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5135_6
timestamp 1731220536
transform 1 0 1104 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5134_6
timestamp 1731220536
transform 1 0 1048 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5133_6
timestamp 1731220536
transform 1 0 840 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5132_6
timestamp 1731220536
transform 1 0 608 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5131_6
timestamp 1731220536
transform 1 0 360 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5130_6
timestamp 1731220536
transform 1 0 712 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5129_6
timestamp 1731220536
transform 1 0 904 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5128_6
timestamp 1731220536
transform 1 0 768 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5127_6
timestamp 1731220536
transform 1 0 624 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5126_6
timestamp 1731220536
transform 1 0 472 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5125_6
timestamp 1731220536
transform 1 0 448 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5124_6
timestamp 1731220536
transform 1 0 560 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5123_6
timestamp 1731220536
transform 1 0 672 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5122_6
timestamp 1731220536
transform 1 0 792 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5121_6
timestamp 1731220536
transform 1 0 632 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5120_6
timestamp 1731220536
transform 1 0 480 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5119_6
timestamp 1731220536
transform 1 0 328 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5118_6
timestamp 1731220536
transform 1 0 184 0 1 2328
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5117_6
timestamp 1731220536
transform 1 0 336 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5116_6
timestamp 1731220536
transform 1 0 232 0 -1 2316
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5115_6
timestamp 1731220536
transform 1 0 160 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5114_6
timestamp 1731220536
transform 1 0 320 0 1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5113_6
timestamp 1731220536
transform 1 0 512 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5112_6
timestamp 1731220536
transform 1 0 304 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5111_6
timestamp 1731220536
transform 1 0 128 0 -1 2144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5110_6
timestamp 1731220536
transform 1 0 128 0 1 1988
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5109_6
timestamp 1731220536
transform 1 0 304 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5108_6
timestamp 1731220536
transform 1 0 128 0 -1 1976
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5107_6
timestamp 1731220536
transform 1 0 128 0 1 1828
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5106_6
timestamp 1731220536
transform 1 0 128 0 -1 1816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5105_6
timestamp 1731220536
transform 1 0 128 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5104_6
timestamp 1731220536
transform 1 0 296 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5103_6
timestamp 1731220536
transform 1 0 504 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5102_6
timestamp 1731220536
transform 1 0 720 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5101_6
timestamp 1731220536
transform 1 0 936 0 1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5100_6
timestamp 1731220536
transform 1 0 864 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_599_6
timestamp 1731220536
transform 1 0 672 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_598_6
timestamp 1731220536
transform 1 0 480 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_597_6
timestamp 1731220536
transform 1 0 296 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_596_6
timestamp 1731220536
transform 1 0 128 0 -1 1668
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_595_6
timestamp 1731220536
transform 1 0 296 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_594_6
timestamp 1731220536
transform 1 0 432 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_593_6
timestamp 1731220536
transform 1 0 576 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_592_6
timestamp 1731220536
transform 1 0 720 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_591_6
timestamp 1731220536
transform 1 0 864 0 1 1516
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_590_6
timestamp 1731220536
transform 1 0 904 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_589_6
timestamp 1731220536
transform 1 0 752 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_588_6
timestamp 1731220536
transform 1 0 600 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_587_6
timestamp 1731220536
transform 1 0 464 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_586_6
timestamp 1731220536
transform 1 0 336 0 -1 1508
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_585_6
timestamp 1731220536
transform 1 0 784 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_584_6
timestamp 1731220536
transform 1 0 592 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_583_6
timestamp 1731220536
transform 1 0 408 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_582_6
timestamp 1731220536
transform 1 0 248 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_581_6
timestamp 1731220536
transform 1 0 128 0 1 1356
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_580_6
timestamp 1731220536
transform 1 0 128 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_579_6
timestamp 1731220536
transform 1 0 264 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_578_6
timestamp 1731220536
transform 1 0 840 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_577_6
timestamp 1731220536
transform 1 0 640 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_576_6
timestamp 1731220536
transform 1 0 440 0 -1 1344
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_575_6
timestamp 1731220536
transform 1 0 432 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_574_6
timestamp 1731220536
transform 1 0 304 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_573_6
timestamp 1731220536
transform 1 0 184 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_572_6
timestamp 1731220536
transform 1 0 560 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_571_6
timestamp 1731220536
transform 1 0 696 0 1 1200
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_570_6
timestamp 1731220536
transform 1 0 680 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_569_6
timestamp 1731220536
transform 1 0 560 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_568_6
timestamp 1731220536
transform 1 0 448 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_567_6
timestamp 1731220536
transform 1 0 800 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_566_6
timestamp 1731220536
transform 1 0 920 0 -1 1192
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_565_6
timestamp 1731220536
transform 1 0 832 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_564_6
timestamp 1731220536
transform 1 0 712 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_563_6
timestamp 1731220536
transform 1 0 600 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_562_6
timestamp 1731220536
transform 1 0 952 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_561_6
timestamp 1731220536
transform 1 0 1072 0 1 1040
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_560_6
timestamp 1731220536
transform 1 0 1200 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_559_6
timestamp 1731220536
transform 1 0 1072 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_558_6
timestamp 1731220536
transform 1 0 944 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_557_6
timestamp 1731220536
transform 1 0 824 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_556_6
timestamp 1731220536
transform 1 0 704 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_555_6
timestamp 1731220536
transform 1 0 1176 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_554_6
timestamp 1731220536
transform 1 0 1016 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_553_6
timestamp 1731220536
transform 1 0 864 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_552_6
timestamp 1731220536
transform 1 0 712 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_551_6
timestamp 1731220536
transform 1 0 568 0 1 880
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_550_6
timestamp 1731220536
transform 1 0 1024 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_549_6
timestamp 1731220536
transform 1 0 864 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_548_6
timestamp 1731220536
transform 1 0 712 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_547_6
timestamp 1731220536
transform 1 0 560 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_546_6
timestamp 1731220536
transform 1 0 416 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_545_6
timestamp 1731220536
transform 1 0 896 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_544_6
timestamp 1731220536
transform 1 0 728 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_543_6
timestamp 1731220536
transform 1 0 568 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_542_6
timestamp 1731220536
transform 1 0 408 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_541_6
timestamp 1731220536
transform 1 0 256 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_540_6
timestamp 1731220536
transform 1 0 712 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_539_6
timestamp 1731220536
transform 1 0 552 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_538_6
timestamp 1731220536
transform 1 0 400 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_537_6
timestamp 1731220536
transform 1 0 248 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_536_6
timestamp 1731220536
transform 1 0 128 0 -1 724
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_535_6
timestamp 1731220536
transform 1 0 128 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_534_6
timestamp 1731220536
transform 1 0 232 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_533_6
timestamp 1731220536
transform 1 0 368 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_532_6
timestamp 1731220536
transform 1 0 504 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_531_6
timestamp 1731220536
transform 1 0 640 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_530_6
timestamp 1731220536
transform 1 0 544 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_529_6
timestamp 1731220536
transform 1 0 424 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_528_6
timestamp 1731220536
transform 1 0 304 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_527_6
timestamp 1731220536
transform 1 0 184 0 -1 560
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_526_6
timestamp 1731220536
transform 1 0 416 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_525_6
timestamp 1731220536
transform 1 0 520 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_524_6
timestamp 1731220536
transform 1 0 624 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_523_6
timestamp 1731220536
transform 1 0 728 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_522_6
timestamp 1731220536
transform 1 0 832 0 1 408
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_521_6
timestamp 1731220536
transform 1 0 1016 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_520_6
timestamp 1731220536
transform 1 0 912 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_519_6
timestamp 1731220536
transform 1 0 808 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_518_6
timestamp 1731220536
transform 1 0 704 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_517_6
timestamp 1731220536
transform 1 0 600 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_516_6
timestamp 1731220536
transform 1 0 968 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_515_6
timestamp 1731220536
transform 1 0 816 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_514_6
timestamp 1731220536
transform 1 0 664 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_513_6
timestamp 1731220536
transform 1 0 520 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_512_6
timestamp 1731220536
transform 1 0 376 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_511_6
timestamp 1731220536
transform 1 0 848 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_510_6
timestamp 1731220536
transform 1 0 632 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_59_6
timestamp 1731220536
transform 1 0 408 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_58_6
timestamp 1731220536
transform 1 0 184 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_57_6
timestamp 1731220536
transform 1 0 856 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_56_6
timestamp 1731220536
transform 1 0 752 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_55_6
timestamp 1731220536
transform 1 0 648 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_54_6
timestamp 1731220536
transform 1 0 544 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_53_6
timestamp 1731220536
transform 1 0 440 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_52_6
timestamp 1731220536
transform 1 0 336 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_51_6
timestamp 1731220536
transform 1 0 232 0 1 80
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_50_6
timestamp 1731220536
transform 1 0 128 0 1 80
box 8 5 100 68
<< end >>
