magic
tech sky130l
timestamp 1731220534
<< m1 >>
rect 576 1691 580 1707
rect 632 1691 636 1707
rect 688 1691 692 1707
rect 752 1691 756 1707
rect 920 1691 924 1707
rect 976 1691 980 1707
rect 1032 1691 1036 1707
rect 1312 1691 1316 1707
rect 1360 1691 1364 1707
rect 1400 1691 1404 1707
rect 1496 1691 1500 1707
rect 208 1611 212 1627
rect 272 1611 276 1627
rect 328 1611 332 1627
rect 384 1611 388 1627
rect 560 1611 564 1627
rect 688 1611 692 1627
rect 824 1611 828 1627
rect 896 1611 900 1627
rect 656 1547 660 1579
rect 384 1531 388 1547
rect 432 1531 436 1547
rect 480 1531 484 1547
rect 536 1531 540 1547
rect 1648 1547 1652 1579
rect 664 1531 668 1547
rect 720 1531 724 1547
rect 1432 1531 1436 1547
rect 1496 1531 1500 1547
rect 1552 1531 1556 1547
rect 1648 1463 1652 1495
rect 552 1447 556 1463
rect 624 1447 628 1463
rect 688 1447 692 1463
rect 744 1447 748 1463
rect 1184 1447 1188 1463
rect 1232 1447 1236 1463
rect 1288 1447 1292 1463
rect 1352 1447 1356 1463
rect 1424 1447 1428 1463
rect 1488 1383 1492 1411
rect 1496 1391 1500 1411
rect 528 1363 532 1379
rect 608 1363 612 1379
rect 768 1363 772 1379
rect 912 1363 916 1379
rect 984 1363 988 1379
rect 1056 1363 1060 1379
rect 1128 1363 1132 1379
rect 1200 1363 1204 1379
rect 1328 1363 1332 1379
rect 1392 1363 1396 1379
rect 1520 1363 1524 1379
rect 1648 1319 1652 1411
rect 160 1279 164 1295
rect 208 1279 212 1295
rect 304 1279 308 1295
rect 352 1279 356 1295
rect 632 1279 636 1295
rect 800 1279 804 1295
rect 856 1279 860 1295
rect 920 1279 924 1295
rect 984 1279 988 1295
rect 1048 1279 1052 1295
rect 1384 1279 1388 1295
rect 1472 1279 1476 1295
rect 792 1227 796 1247
rect 192 1195 196 1211
rect 360 1195 364 1211
rect 456 1195 460 1211
rect 512 1195 516 1211
rect 568 1195 572 1211
rect 624 1195 628 1211
rect 680 1195 684 1211
rect 792 1195 796 1211
rect 848 1195 852 1211
rect 1040 1195 1044 1211
rect 1168 1195 1172 1211
rect 1232 1195 1236 1211
rect 1304 1195 1308 1211
rect 1384 1195 1388 1211
rect 1472 1195 1476 1211
rect 1648 1163 1652 1291
rect 1544 1135 1548 1159
rect 200 1107 204 1123
rect 240 1107 244 1123
rect 360 1107 364 1123
rect 424 1107 428 1123
rect 552 1107 556 1123
rect 624 1107 628 1123
rect 688 1107 692 1123
rect 752 1107 756 1123
rect 816 1107 820 1123
rect 936 1107 940 1123
rect 992 1107 996 1123
rect 1176 1107 1180 1123
rect 1240 1107 1244 1123
rect 1360 1107 1364 1123
rect 1416 1107 1420 1123
rect 1472 1107 1476 1123
rect 1568 1107 1572 1123
rect 528 1019 532 1035
rect 584 1019 588 1035
rect 656 1019 660 1035
rect 824 1019 828 1035
rect 984 1019 988 1035
rect 1056 1019 1060 1035
rect 1120 1019 1124 1035
rect 1184 1019 1188 1035
rect 1248 1019 1252 1035
rect 1360 1019 1364 1035
rect 224 939 228 955
rect 264 939 268 955
rect 312 939 316 955
rect 368 939 372 955
rect 496 939 500 955
rect 560 939 564 955
rect 624 939 628 955
rect 872 939 876 955
rect 936 939 940 955
rect 1000 939 1004 955
rect 1064 939 1068 955
rect 1128 939 1132 955
rect 1416 939 1420 955
rect 192 851 196 867
rect 232 851 236 867
rect 296 851 300 867
rect 360 851 364 867
rect 496 851 500 867
rect 728 851 732 867
rect 1064 851 1068 867
rect 1192 851 1196 867
rect 1256 851 1260 867
rect 1312 851 1316 867
rect 1368 851 1372 867
rect 1424 851 1428 867
rect 1064 799 1068 819
rect 160 767 164 783
rect 200 767 204 783
rect 392 767 396 783
rect 552 767 556 783
rect 728 767 732 783
rect 816 767 820 783
rect 976 767 980 783
rect 1048 767 1052 783
rect 1120 767 1124 783
rect 1192 767 1196 783
rect 1256 767 1260 783
rect 1384 767 1388 783
rect 1440 767 1444 783
rect 464 703 468 735
rect 528 683 532 699
rect 568 683 572 699
rect 616 683 620 699
rect 672 683 676 699
rect 784 683 788 699
rect 848 683 852 699
rect 1048 683 1052 699
rect 1184 683 1188 699
rect 1208 695 1212 735
rect 1248 683 1252 699
rect 1312 683 1316 699
rect 1376 683 1380 699
rect 1496 683 1500 699
rect 1608 683 1612 699
rect 1648 619 1652 651
rect 304 603 308 619
rect 352 603 356 619
rect 392 603 396 619
rect 448 603 452 619
rect 544 603 548 619
rect 592 603 596 619
rect 640 603 644 619
rect 688 603 692 619
rect 744 603 748 619
rect 856 603 860 619
rect 920 603 924 619
rect 1072 603 1076 619
rect 1384 603 1388 619
rect 1456 603 1460 619
rect 1528 603 1532 619
rect 904 551 908 571
rect 1648 535 1652 571
rect 256 519 260 535
rect 304 519 308 535
rect 400 519 404 535
rect 712 519 716 535
rect 904 519 908 535
rect 968 519 972 535
rect 1256 519 1260 535
rect 1304 519 1308 535
rect 1360 519 1364 535
rect 1416 519 1420 535
rect 1472 519 1476 535
rect 264 467 268 487
rect 360 459 364 487
rect 640 467 644 487
rect 232 439 236 455
rect 352 427 356 451
rect 392 439 396 455
rect 512 411 516 455
rect 544 439 548 455
rect 624 439 628 455
rect 864 439 868 455
rect 1288 439 1292 455
rect 1192 375 1196 407
rect 1408 387 1412 407
rect 488 355 492 371
rect 544 355 548 371
rect 600 355 604 371
rect 768 355 772 371
rect 944 355 948 371
rect 1008 355 1012 371
rect 1280 355 1284 371
rect 1328 355 1332 371
rect 1376 355 1380 371
rect 1520 355 1524 371
rect 1568 355 1572 371
rect 656 303 660 323
rect 776 291 780 323
rect 1368 311 1372 339
rect 1648 291 1652 323
rect 784 275 788 291
rect 832 275 836 291
rect 904 275 908 291
rect 976 275 980 291
rect 1136 275 1140 291
rect 1216 275 1220 291
rect 1352 275 1356 291
rect 400 191 404 207
rect 440 191 444 207
rect 640 191 644 207
rect 720 191 724 207
rect 880 191 884 207
rect 952 191 956 207
rect 1024 191 1028 207
rect 1096 191 1100 207
rect 1168 191 1172 207
rect 1552 191 1556 207
rect 1608 191 1612 207
rect 1648 111 1652 159
rect 488 95 492 111
rect 528 95 532 111
rect 920 95 924 111
rect 960 95 964 111
rect 1000 95 1004 111
rect 1040 95 1044 111
rect 1088 95 1092 111
rect 1128 95 1132 111
rect 1208 95 1212 111
rect 1248 95 1252 111
rect 1320 95 1324 111
rect 1360 95 1364 111
rect 1400 95 1404 111
rect 1440 95 1444 111
rect 1480 95 1484 111
rect 1528 95 1532 111
<< m2c >>
rect 576 1707 580 1711
rect 632 1707 636 1711
rect 688 1707 692 1711
rect 752 1707 756 1711
rect 920 1707 924 1711
rect 976 1707 980 1711
rect 1032 1707 1036 1711
rect 272 1703 276 1707
rect 304 1703 308 1707
rect 336 1703 340 1707
rect 376 1703 380 1707
rect 424 1703 428 1707
rect 520 1703 524 1707
rect 568 1703 572 1707
rect 624 1703 628 1707
rect 680 1703 684 1707
rect 744 1703 748 1707
rect 800 1703 804 1707
rect 856 1703 860 1707
rect 912 1703 916 1707
rect 968 1703 972 1707
rect 1024 1703 1028 1707
rect 1080 1703 1084 1707
rect 1136 1703 1140 1707
rect 1192 1705 1196 1709
rect 1312 1707 1316 1711
rect 1360 1707 1364 1711
rect 1400 1707 1404 1711
rect 1496 1707 1500 1711
rect 1248 1703 1252 1707
rect 1304 1703 1308 1707
rect 1352 1703 1356 1707
rect 1392 1703 1396 1707
rect 1440 1703 1444 1707
rect 1488 1703 1492 1707
rect 1536 1703 1540 1707
rect 272 1687 276 1691
rect 304 1687 308 1691
rect 336 1687 340 1691
rect 376 1687 380 1691
rect 424 1687 428 1691
rect 472 1687 476 1691
rect 520 1687 524 1691
rect 568 1687 572 1691
rect 576 1687 580 1691
rect 624 1687 628 1691
rect 632 1687 636 1691
rect 680 1687 684 1691
rect 688 1687 692 1691
rect 744 1687 748 1691
rect 752 1687 756 1691
rect 800 1687 804 1691
rect 856 1687 860 1691
rect 912 1687 916 1691
rect 920 1687 924 1691
rect 968 1687 972 1691
rect 976 1687 980 1691
rect 1024 1687 1028 1691
rect 1032 1687 1036 1691
rect 1080 1687 1084 1691
rect 1136 1687 1140 1691
rect 1192 1687 1196 1691
rect 1248 1687 1252 1691
rect 1304 1687 1308 1691
rect 1312 1687 1316 1691
rect 1352 1687 1356 1691
rect 1360 1687 1364 1691
rect 1392 1687 1396 1691
rect 1400 1687 1404 1691
rect 1440 1687 1444 1691
rect 1488 1687 1492 1691
rect 1496 1687 1500 1691
rect 1536 1687 1540 1691
rect 152 1659 156 1663
rect 184 1659 188 1663
rect 232 1659 236 1663
rect 296 1659 300 1663
rect 360 1659 364 1663
rect 432 1659 436 1663
rect 504 1661 508 1665
rect 576 1659 580 1663
rect 648 1659 652 1663
rect 728 1659 732 1663
rect 808 1659 812 1663
rect 888 1659 892 1663
rect 968 1659 972 1663
rect 1048 1659 1052 1663
rect 1120 1659 1124 1663
rect 1192 1659 1196 1663
rect 1264 1659 1268 1663
rect 1336 1659 1340 1663
rect 1408 1659 1412 1663
rect 1472 1659 1476 1663
rect 1536 1659 1540 1663
rect 1600 1659 1604 1663
rect 1640 1659 1644 1663
rect 152 1643 156 1647
rect 184 1643 188 1647
rect 232 1643 236 1647
rect 296 1643 300 1647
rect 360 1643 364 1647
rect 432 1643 436 1647
rect 504 1643 508 1647
rect 576 1643 580 1647
rect 648 1643 652 1647
rect 728 1643 732 1647
rect 808 1643 812 1647
rect 888 1643 892 1647
rect 968 1643 972 1647
rect 1048 1643 1052 1647
rect 1120 1643 1124 1647
rect 1192 1643 1196 1647
rect 1264 1643 1268 1647
rect 1336 1643 1340 1647
rect 1408 1643 1412 1647
rect 1472 1643 1476 1647
rect 1536 1643 1540 1647
rect 1600 1643 1604 1647
rect 1640 1643 1644 1647
rect 208 1627 212 1631
rect 272 1627 276 1631
rect 328 1627 332 1631
rect 384 1627 388 1631
rect 560 1627 564 1631
rect 688 1627 692 1631
rect 824 1627 828 1631
rect 896 1627 900 1631
rect 152 1623 156 1627
rect 200 1623 204 1627
rect 264 1623 268 1627
rect 320 1623 324 1627
rect 376 1623 380 1627
rect 432 1623 436 1627
rect 488 1623 492 1627
rect 552 1623 556 1627
rect 616 1623 620 1627
rect 680 1623 684 1627
rect 744 1623 748 1627
rect 816 1623 820 1627
rect 888 1623 892 1627
rect 960 1623 964 1627
rect 1040 1623 1044 1627
rect 1120 1623 1124 1627
rect 1192 1623 1196 1627
rect 1264 1623 1268 1627
rect 1336 1623 1340 1627
rect 1416 1623 1420 1627
rect 1496 1623 1500 1627
rect 1576 1623 1580 1627
rect 1640 1623 1644 1627
rect 152 1607 156 1611
rect 200 1607 204 1611
rect 208 1607 212 1611
rect 264 1607 268 1611
rect 272 1607 276 1611
rect 320 1607 324 1611
rect 328 1607 332 1611
rect 376 1607 380 1611
rect 384 1607 388 1611
rect 432 1607 436 1611
rect 488 1607 492 1611
rect 552 1607 556 1611
rect 560 1607 564 1611
rect 616 1607 620 1611
rect 680 1607 684 1611
rect 688 1607 692 1611
rect 744 1607 748 1611
rect 816 1607 820 1611
rect 824 1607 828 1611
rect 888 1607 892 1611
rect 896 1607 900 1611
rect 960 1607 964 1611
rect 1040 1607 1044 1611
rect 1120 1607 1124 1611
rect 1192 1607 1196 1611
rect 1264 1607 1268 1611
rect 1336 1607 1340 1611
rect 1416 1607 1420 1611
rect 1496 1607 1500 1611
rect 1576 1607 1580 1611
rect 1640 1607 1644 1611
rect 152 1579 156 1583
rect 184 1579 188 1583
rect 240 1579 244 1583
rect 296 1581 300 1585
rect 352 1579 356 1583
rect 400 1579 404 1583
rect 448 1579 452 1583
rect 496 1579 500 1583
rect 552 1579 556 1583
rect 616 1579 620 1583
rect 656 1579 660 1583
rect 680 1579 684 1583
rect 744 1579 748 1583
rect 816 1579 820 1583
rect 888 1579 892 1583
rect 968 1579 972 1583
rect 1056 1579 1060 1583
rect 1136 1579 1140 1583
rect 1216 1579 1220 1583
rect 1296 1579 1300 1583
rect 1368 1579 1372 1583
rect 1432 1579 1436 1583
rect 1488 1579 1492 1583
rect 1544 1579 1548 1583
rect 1600 1579 1604 1583
rect 1640 1579 1644 1583
rect 1648 1579 1652 1583
rect 152 1563 156 1567
rect 184 1563 188 1567
rect 240 1563 244 1567
rect 296 1563 300 1567
rect 352 1563 356 1567
rect 400 1563 404 1567
rect 448 1563 452 1567
rect 496 1563 500 1567
rect 552 1563 556 1567
rect 616 1563 620 1567
rect 384 1547 388 1551
rect 432 1547 436 1551
rect 480 1547 484 1551
rect 536 1547 540 1551
rect 680 1563 684 1567
rect 744 1563 748 1567
rect 816 1563 820 1567
rect 888 1563 892 1567
rect 968 1563 972 1567
rect 1056 1563 1060 1567
rect 1136 1563 1140 1567
rect 1216 1563 1220 1567
rect 1296 1563 1300 1567
rect 1368 1563 1372 1567
rect 1432 1563 1436 1567
rect 1488 1563 1492 1567
rect 1544 1563 1548 1567
rect 1600 1563 1604 1567
rect 1640 1563 1644 1567
rect 152 1543 156 1547
rect 184 1543 188 1547
rect 232 1543 236 1547
rect 280 1543 284 1547
rect 328 1543 332 1547
rect 376 1543 380 1547
rect 424 1543 428 1547
rect 472 1543 476 1547
rect 528 1543 532 1547
rect 584 1543 588 1547
rect 648 1543 652 1547
rect 656 1543 660 1547
rect 664 1547 668 1551
rect 720 1547 724 1551
rect 1432 1547 1436 1551
rect 1496 1547 1500 1551
rect 1552 1547 1556 1551
rect 712 1543 716 1547
rect 776 1543 780 1547
rect 848 1543 852 1547
rect 936 1543 940 1547
rect 1024 1543 1028 1547
rect 1112 1543 1116 1547
rect 1200 1543 1204 1547
rect 1280 1543 1284 1547
rect 1352 1543 1356 1547
rect 1424 1543 1428 1547
rect 1488 1543 1492 1547
rect 1544 1543 1548 1547
rect 1600 1543 1604 1547
rect 1640 1543 1644 1547
rect 1648 1543 1652 1547
rect 152 1527 156 1531
rect 184 1527 188 1531
rect 232 1527 236 1531
rect 280 1527 284 1531
rect 328 1527 332 1531
rect 376 1527 380 1531
rect 384 1527 388 1531
rect 424 1527 428 1531
rect 432 1527 436 1531
rect 472 1527 476 1531
rect 480 1527 484 1531
rect 528 1527 532 1531
rect 536 1527 540 1531
rect 584 1527 588 1531
rect 648 1527 652 1531
rect 664 1527 668 1531
rect 712 1527 716 1531
rect 720 1527 724 1531
rect 776 1527 780 1531
rect 848 1527 852 1531
rect 936 1527 940 1531
rect 1024 1527 1028 1531
rect 1112 1527 1116 1531
rect 1200 1527 1204 1531
rect 1280 1527 1284 1531
rect 1352 1527 1356 1531
rect 1424 1527 1428 1531
rect 1432 1527 1436 1531
rect 1488 1527 1492 1531
rect 1496 1527 1500 1531
rect 1544 1527 1548 1531
rect 1552 1527 1556 1531
rect 1600 1527 1604 1531
rect 1640 1527 1644 1531
rect 152 1495 156 1499
rect 184 1495 188 1499
rect 240 1495 244 1499
rect 312 1495 316 1499
rect 392 1495 396 1499
rect 472 1495 476 1499
rect 544 1495 548 1499
rect 616 1495 620 1499
rect 688 1495 692 1499
rect 760 1495 764 1499
rect 832 1495 836 1499
rect 896 1495 900 1499
rect 960 1495 964 1499
rect 1024 1495 1028 1499
rect 1080 1495 1084 1499
rect 1128 1495 1132 1499
rect 1168 1495 1172 1499
rect 1200 1495 1204 1499
rect 1232 1495 1236 1499
rect 1272 1495 1276 1499
rect 1312 1495 1316 1499
rect 1368 1495 1372 1499
rect 1432 1495 1436 1499
rect 1504 1495 1508 1499
rect 1584 1495 1588 1499
rect 1640 1495 1644 1499
rect 1648 1495 1652 1499
rect 152 1479 156 1483
rect 184 1479 188 1483
rect 240 1479 244 1483
rect 312 1479 316 1483
rect 392 1479 396 1483
rect 472 1479 476 1483
rect 544 1479 548 1483
rect 616 1479 620 1483
rect 688 1479 692 1483
rect 760 1479 764 1483
rect 832 1479 836 1483
rect 896 1479 900 1483
rect 960 1479 964 1483
rect 1024 1479 1028 1483
rect 1080 1479 1084 1483
rect 1128 1479 1132 1483
rect 1168 1479 1172 1483
rect 1200 1479 1204 1483
rect 1232 1479 1236 1483
rect 1272 1479 1276 1483
rect 1312 1479 1316 1483
rect 1368 1479 1372 1483
rect 1432 1479 1436 1483
rect 1504 1479 1508 1483
rect 1584 1479 1588 1483
rect 1640 1479 1644 1483
rect 552 1463 556 1467
rect 624 1463 628 1467
rect 688 1463 692 1467
rect 744 1463 748 1467
rect 1184 1463 1188 1467
rect 1232 1463 1236 1467
rect 1288 1463 1292 1467
rect 1352 1463 1356 1467
rect 1424 1463 1428 1467
rect 152 1459 156 1463
rect 184 1459 188 1463
rect 240 1459 244 1463
rect 312 1459 316 1463
rect 392 1459 396 1463
rect 472 1459 476 1463
rect 544 1459 548 1463
rect 616 1459 620 1463
rect 680 1459 684 1463
rect 736 1459 740 1463
rect 800 1459 804 1463
rect 864 1459 868 1463
rect 920 1459 924 1463
rect 976 1459 980 1463
rect 1032 1459 1036 1463
rect 1088 1459 1092 1463
rect 1136 1459 1140 1463
rect 1176 1459 1180 1463
rect 1224 1459 1228 1463
rect 1280 1459 1284 1463
rect 1344 1459 1348 1463
rect 1416 1459 1420 1463
rect 1496 1459 1500 1463
rect 1576 1459 1580 1463
rect 1640 1459 1644 1463
rect 1648 1459 1652 1463
rect 152 1443 156 1447
rect 184 1443 188 1447
rect 240 1443 244 1447
rect 312 1443 316 1447
rect 392 1443 396 1447
rect 472 1443 476 1447
rect 544 1443 548 1447
rect 552 1443 556 1447
rect 616 1443 620 1447
rect 624 1443 628 1447
rect 680 1443 684 1447
rect 688 1443 692 1447
rect 736 1443 740 1447
rect 744 1443 748 1447
rect 800 1443 804 1447
rect 864 1443 868 1447
rect 920 1443 924 1447
rect 976 1443 980 1447
rect 1032 1443 1036 1447
rect 1088 1443 1092 1447
rect 1136 1443 1140 1447
rect 1176 1443 1180 1447
rect 1184 1443 1188 1447
rect 1224 1443 1228 1447
rect 1232 1443 1236 1447
rect 1280 1443 1284 1447
rect 1288 1443 1292 1447
rect 1344 1443 1348 1447
rect 1352 1443 1356 1447
rect 1416 1443 1420 1447
rect 1424 1443 1428 1447
rect 1496 1443 1500 1447
rect 1576 1443 1580 1447
rect 1640 1443 1644 1447
rect 152 1411 156 1415
rect 184 1411 188 1415
rect 232 1411 236 1415
rect 304 1411 308 1415
rect 376 1411 380 1415
rect 456 1411 460 1415
rect 536 1411 540 1415
rect 616 1411 620 1415
rect 696 1411 700 1415
rect 776 1411 780 1415
rect 848 1411 852 1415
rect 920 1411 924 1415
rect 984 1411 988 1415
rect 1048 1411 1052 1415
rect 1120 1411 1124 1415
rect 1184 1411 1188 1415
rect 1248 1411 1252 1415
rect 1312 1411 1316 1415
rect 1376 1411 1380 1415
rect 1432 1411 1436 1415
rect 1480 1411 1484 1415
rect 1488 1411 1492 1415
rect 152 1395 156 1399
rect 184 1395 188 1399
rect 232 1395 236 1399
rect 304 1395 308 1399
rect 376 1395 380 1399
rect 456 1395 460 1399
rect 536 1395 540 1399
rect 616 1395 620 1399
rect 696 1395 700 1399
rect 776 1395 780 1399
rect 848 1395 852 1399
rect 920 1395 924 1399
rect 984 1395 988 1399
rect 1048 1395 1052 1399
rect 1120 1395 1124 1399
rect 1184 1395 1188 1399
rect 1248 1395 1252 1399
rect 1312 1395 1316 1399
rect 1376 1395 1380 1399
rect 1432 1395 1436 1399
rect 1480 1395 1484 1399
rect 1496 1411 1500 1415
rect 1520 1411 1524 1415
rect 1568 1411 1572 1415
rect 1608 1411 1612 1415
rect 1640 1411 1644 1415
rect 1648 1411 1652 1415
rect 1520 1395 1524 1399
rect 1568 1395 1572 1399
rect 1608 1395 1612 1399
rect 1640 1395 1644 1399
rect 1496 1387 1500 1391
rect 528 1379 532 1383
rect 608 1379 612 1383
rect 768 1379 772 1383
rect 912 1379 916 1383
rect 984 1379 988 1383
rect 1056 1379 1060 1383
rect 1128 1379 1132 1383
rect 1200 1379 1204 1383
rect 1328 1379 1332 1383
rect 1392 1379 1396 1383
rect 1488 1379 1492 1383
rect 1520 1379 1524 1383
rect 152 1375 156 1379
rect 184 1375 188 1379
rect 240 1375 244 1379
rect 304 1375 308 1379
rect 376 1375 380 1379
rect 448 1375 452 1379
rect 520 1375 524 1379
rect 600 1375 604 1379
rect 680 1375 684 1379
rect 760 1375 764 1379
rect 832 1375 836 1379
rect 904 1375 908 1379
rect 976 1375 980 1379
rect 1048 1375 1052 1379
rect 1120 1375 1124 1379
rect 1192 1375 1196 1379
rect 1256 1375 1260 1379
rect 1320 1375 1324 1379
rect 1384 1375 1388 1379
rect 1448 1375 1452 1379
rect 1512 1375 1516 1379
rect 1584 1375 1588 1379
rect 1640 1375 1644 1379
rect 152 1359 156 1363
rect 184 1359 188 1363
rect 240 1359 244 1363
rect 304 1359 308 1363
rect 376 1359 380 1363
rect 448 1359 452 1363
rect 520 1359 524 1363
rect 528 1359 532 1363
rect 600 1359 604 1363
rect 608 1359 612 1363
rect 680 1359 684 1363
rect 760 1359 764 1363
rect 768 1359 772 1363
rect 832 1359 836 1363
rect 904 1359 908 1363
rect 912 1359 916 1363
rect 976 1359 980 1363
rect 984 1359 988 1363
rect 1048 1359 1052 1363
rect 1056 1359 1060 1363
rect 1120 1359 1124 1363
rect 1128 1359 1132 1363
rect 1192 1359 1196 1363
rect 1200 1359 1204 1363
rect 1256 1359 1260 1363
rect 1320 1359 1324 1363
rect 1328 1359 1332 1363
rect 1384 1359 1388 1363
rect 1392 1359 1396 1363
rect 1448 1359 1452 1363
rect 1512 1359 1516 1363
rect 1520 1359 1524 1363
rect 1584 1359 1588 1363
rect 1640 1359 1644 1363
rect 152 1331 156 1335
rect 200 1331 204 1335
rect 256 1331 260 1335
rect 312 1331 316 1335
rect 368 1331 372 1335
rect 416 1331 420 1335
rect 472 1331 476 1335
rect 528 1331 532 1335
rect 584 1331 588 1335
rect 648 1331 652 1335
rect 712 1331 716 1335
rect 776 1331 780 1335
rect 840 1331 844 1335
rect 904 1331 908 1335
rect 976 1331 980 1335
rect 1040 1331 1044 1335
rect 1104 1331 1108 1335
rect 1168 1331 1172 1335
rect 1232 1331 1236 1335
rect 1296 1331 1300 1335
rect 1360 1331 1364 1335
rect 1424 1331 1428 1335
rect 1496 1331 1500 1335
rect 1576 1331 1580 1335
rect 1640 1331 1644 1335
rect 152 1315 156 1319
rect 200 1315 204 1319
rect 256 1315 260 1319
rect 312 1315 316 1319
rect 368 1315 372 1319
rect 416 1315 420 1319
rect 472 1315 476 1319
rect 528 1315 532 1319
rect 584 1315 588 1319
rect 648 1315 652 1319
rect 712 1315 716 1319
rect 776 1315 780 1319
rect 840 1315 844 1319
rect 904 1315 908 1319
rect 976 1315 980 1319
rect 1040 1315 1044 1319
rect 1104 1315 1108 1319
rect 1168 1315 1172 1319
rect 1232 1315 1236 1319
rect 1296 1315 1300 1319
rect 1360 1315 1364 1319
rect 1424 1315 1428 1319
rect 1496 1315 1500 1319
rect 1576 1315 1580 1319
rect 1640 1315 1644 1319
rect 1648 1315 1652 1319
rect 160 1295 164 1299
rect 208 1295 212 1299
rect 304 1295 308 1299
rect 352 1295 356 1299
rect 632 1295 636 1299
rect 800 1295 804 1299
rect 856 1295 860 1299
rect 920 1295 924 1299
rect 984 1295 988 1299
rect 1048 1295 1052 1299
rect 1384 1295 1388 1299
rect 1472 1295 1476 1299
rect 152 1291 156 1295
rect 200 1291 204 1295
rect 248 1291 252 1295
rect 296 1291 300 1295
rect 344 1291 348 1295
rect 392 1291 396 1295
rect 448 1291 452 1295
rect 504 1291 508 1295
rect 560 1291 564 1295
rect 624 1291 628 1295
rect 680 1291 684 1295
rect 736 1291 740 1295
rect 792 1291 796 1295
rect 848 1291 852 1295
rect 912 1291 916 1295
rect 976 1291 980 1295
rect 1040 1291 1044 1295
rect 1096 1291 1100 1295
rect 1160 1291 1164 1295
rect 1224 1291 1228 1295
rect 1296 1291 1300 1295
rect 1376 1291 1380 1295
rect 1464 1291 1468 1295
rect 1560 1291 1564 1295
rect 1640 1291 1644 1295
rect 1648 1291 1652 1295
rect 152 1275 156 1279
rect 160 1275 164 1279
rect 200 1275 204 1279
rect 208 1275 212 1279
rect 248 1275 252 1279
rect 296 1275 300 1279
rect 304 1275 308 1279
rect 344 1275 348 1279
rect 352 1275 356 1279
rect 392 1275 396 1279
rect 448 1275 452 1279
rect 504 1275 508 1279
rect 560 1275 564 1279
rect 624 1275 628 1279
rect 632 1275 636 1279
rect 680 1275 684 1279
rect 736 1275 740 1279
rect 792 1275 796 1279
rect 800 1275 804 1279
rect 848 1275 852 1279
rect 856 1275 860 1279
rect 912 1275 916 1279
rect 920 1275 924 1279
rect 976 1275 980 1279
rect 984 1275 988 1279
rect 1040 1275 1044 1279
rect 1048 1275 1052 1279
rect 1096 1275 1100 1279
rect 1160 1275 1164 1279
rect 1224 1275 1228 1279
rect 1296 1275 1300 1279
rect 1376 1275 1380 1279
rect 1384 1275 1388 1279
rect 1464 1275 1468 1279
rect 1472 1275 1476 1279
rect 1560 1275 1564 1279
rect 1640 1275 1644 1279
rect 152 1247 156 1251
rect 184 1247 188 1251
rect 240 1247 244 1251
rect 296 1247 300 1251
rect 344 1247 348 1251
rect 400 1247 404 1251
rect 456 1247 460 1251
rect 512 1247 516 1251
rect 568 1247 572 1251
rect 624 1247 628 1251
rect 680 1247 684 1251
rect 736 1247 740 1251
rect 784 1247 788 1251
rect 792 1247 796 1251
rect 832 1247 836 1251
rect 888 1247 892 1251
rect 944 1247 948 1251
rect 1000 1247 1004 1251
rect 1056 1247 1060 1251
rect 1112 1247 1116 1251
rect 1176 1247 1180 1251
rect 1248 1247 1252 1251
rect 1336 1247 1340 1251
rect 1440 1247 1444 1251
rect 1552 1247 1556 1251
rect 1640 1247 1644 1251
rect 152 1231 156 1235
rect 184 1231 188 1235
rect 240 1231 244 1235
rect 296 1231 300 1235
rect 344 1231 348 1235
rect 400 1231 404 1235
rect 456 1231 460 1235
rect 512 1231 516 1235
rect 568 1231 572 1235
rect 624 1231 628 1235
rect 680 1231 684 1235
rect 736 1231 740 1235
rect 784 1231 788 1235
rect 832 1231 836 1235
rect 888 1231 892 1235
rect 944 1231 948 1235
rect 1000 1231 1004 1235
rect 1056 1231 1060 1235
rect 1112 1231 1116 1235
rect 1176 1231 1180 1235
rect 1248 1231 1252 1235
rect 1336 1231 1340 1235
rect 1440 1231 1444 1235
rect 1552 1231 1556 1235
rect 1640 1231 1644 1235
rect 792 1223 796 1227
rect 192 1211 196 1215
rect 360 1211 364 1215
rect 456 1211 460 1215
rect 512 1211 516 1215
rect 568 1211 572 1215
rect 624 1211 628 1215
rect 680 1211 684 1215
rect 792 1211 796 1215
rect 848 1211 852 1215
rect 1040 1211 1044 1215
rect 1168 1211 1172 1215
rect 1232 1211 1236 1215
rect 1304 1211 1308 1215
rect 1384 1211 1388 1215
rect 1472 1211 1476 1215
rect 152 1207 156 1211
rect 184 1207 188 1211
rect 240 1207 244 1211
rect 296 1207 300 1211
rect 352 1207 356 1211
rect 400 1207 404 1211
rect 448 1207 452 1211
rect 504 1207 508 1211
rect 560 1207 564 1211
rect 616 1207 620 1211
rect 672 1207 676 1211
rect 728 1207 732 1211
rect 784 1207 788 1211
rect 840 1207 844 1211
rect 904 1207 908 1211
rect 968 1207 972 1211
rect 1032 1207 1036 1211
rect 1096 1207 1100 1211
rect 1160 1207 1164 1211
rect 1224 1207 1228 1211
rect 1296 1207 1300 1211
rect 1376 1207 1380 1211
rect 1464 1207 1468 1211
rect 1560 1207 1564 1211
rect 1640 1207 1644 1211
rect 152 1191 156 1195
rect 184 1191 188 1195
rect 192 1191 196 1195
rect 240 1191 244 1195
rect 296 1191 300 1195
rect 352 1191 356 1195
rect 360 1191 364 1195
rect 400 1191 404 1195
rect 448 1191 452 1195
rect 456 1191 460 1195
rect 504 1191 508 1195
rect 512 1191 516 1195
rect 560 1191 564 1195
rect 568 1191 572 1195
rect 616 1191 620 1195
rect 624 1191 628 1195
rect 672 1191 676 1195
rect 680 1191 684 1195
rect 728 1191 732 1195
rect 784 1191 788 1195
rect 792 1191 796 1195
rect 840 1191 844 1195
rect 848 1191 852 1195
rect 904 1191 908 1195
rect 968 1191 972 1195
rect 1032 1191 1036 1195
rect 1040 1191 1044 1195
rect 1096 1191 1100 1195
rect 1160 1191 1164 1195
rect 1168 1191 1172 1195
rect 1224 1191 1228 1195
rect 1232 1191 1236 1195
rect 1296 1191 1300 1195
rect 1304 1191 1308 1195
rect 1376 1191 1380 1195
rect 1384 1191 1388 1195
rect 1464 1191 1468 1195
rect 1472 1191 1476 1195
rect 1560 1191 1564 1195
rect 1640 1191 1644 1195
rect 152 1159 156 1163
rect 184 1159 188 1163
rect 240 1159 244 1163
rect 304 1159 308 1163
rect 368 1159 372 1163
rect 432 1159 436 1163
rect 488 1159 492 1163
rect 552 1159 556 1163
rect 616 1159 620 1163
rect 680 1159 684 1163
rect 744 1159 748 1163
rect 800 1159 804 1163
rect 856 1159 860 1163
rect 920 1159 924 1163
rect 984 1159 988 1163
rect 1048 1159 1052 1163
rect 1112 1159 1116 1163
rect 1176 1159 1180 1163
rect 1232 1159 1236 1163
rect 1296 1159 1300 1163
rect 1360 1159 1364 1163
rect 1424 1159 1428 1163
rect 1496 1159 1500 1163
rect 1544 1159 1548 1163
rect 1576 1159 1580 1163
rect 1640 1159 1644 1163
rect 1648 1159 1652 1163
rect 152 1143 156 1147
rect 184 1143 188 1147
rect 240 1143 244 1147
rect 304 1143 308 1147
rect 368 1143 372 1147
rect 432 1143 436 1147
rect 488 1143 492 1147
rect 552 1143 556 1147
rect 616 1143 620 1147
rect 680 1143 684 1147
rect 744 1143 748 1147
rect 800 1143 804 1147
rect 856 1143 860 1147
rect 920 1143 924 1147
rect 984 1143 988 1147
rect 1048 1143 1052 1147
rect 1112 1143 1116 1147
rect 1176 1143 1180 1147
rect 1232 1143 1236 1147
rect 1296 1143 1300 1147
rect 1360 1143 1364 1147
rect 1424 1143 1428 1147
rect 1496 1143 1500 1147
rect 1576 1143 1580 1147
rect 1640 1143 1644 1147
rect 1544 1131 1548 1135
rect 200 1123 204 1127
rect 240 1123 244 1127
rect 360 1123 364 1127
rect 424 1123 428 1127
rect 552 1123 556 1127
rect 624 1123 628 1127
rect 688 1123 692 1127
rect 752 1123 756 1127
rect 816 1123 820 1127
rect 936 1123 940 1127
rect 992 1123 996 1127
rect 1176 1123 1180 1127
rect 1240 1123 1244 1127
rect 1360 1123 1364 1127
rect 1416 1123 1420 1127
rect 1472 1123 1476 1127
rect 1568 1123 1572 1127
rect 160 1119 164 1123
rect 192 1119 196 1123
rect 232 1119 236 1123
rect 288 1119 292 1123
rect 352 1119 356 1123
rect 416 1119 420 1123
rect 480 1119 484 1123
rect 544 1119 548 1123
rect 616 1119 620 1123
rect 680 1119 684 1123
rect 744 1119 748 1123
rect 808 1119 812 1123
rect 872 1119 876 1123
rect 928 1119 932 1123
rect 984 1119 988 1123
rect 1040 1119 1044 1123
rect 1104 1119 1108 1123
rect 1168 1119 1172 1123
rect 1232 1119 1236 1123
rect 1296 1119 1300 1123
rect 1352 1119 1356 1123
rect 1408 1119 1412 1123
rect 1464 1119 1468 1123
rect 1512 1119 1516 1123
rect 1560 1119 1564 1123
rect 1608 1119 1612 1123
rect 1640 1119 1644 1123
rect 160 1103 164 1107
rect 192 1103 196 1107
rect 200 1103 204 1107
rect 232 1103 236 1107
rect 240 1103 244 1107
rect 288 1103 292 1107
rect 352 1103 356 1107
rect 360 1103 364 1107
rect 416 1103 420 1107
rect 424 1103 428 1107
rect 480 1103 484 1107
rect 544 1103 548 1107
rect 552 1103 556 1107
rect 616 1103 620 1107
rect 624 1103 628 1107
rect 680 1103 684 1107
rect 688 1103 692 1107
rect 744 1103 748 1107
rect 752 1103 756 1107
rect 808 1103 812 1107
rect 816 1103 820 1107
rect 872 1103 876 1107
rect 928 1103 932 1107
rect 936 1103 940 1107
rect 984 1103 988 1107
rect 992 1103 996 1107
rect 1040 1103 1044 1107
rect 1104 1103 1108 1107
rect 1168 1103 1172 1107
rect 1176 1103 1180 1107
rect 1232 1103 1236 1107
rect 1240 1103 1244 1107
rect 1296 1103 1300 1107
rect 1352 1103 1356 1107
rect 1360 1103 1364 1107
rect 1408 1103 1412 1107
rect 1416 1103 1420 1107
rect 1464 1103 1468 1107
rect 1472 1103 1476 1107
rect 1512 1103 1516 1107
rect 1560 1103 1564 1107
rect 1568 1103 1572 1107
rect 1608 1103 1612 1107
rect 1640 1103 1644 1107
rect 232 1071 236 1075
rect 264 1071 268 1075
rect 296 1071 300 1075
rect 328 1071 332 1075
rect 368 1071 372 1075
rect 408 1071 412 1075
rect 456 1071 460 1075
rect 520 1071 524 1075
rect 592 1071 596 1075
rect 672 1071 676 1075
rect 752 1071 756 1075
rect 832 1071 836 1075
rect 912 1071 916 1075
rect 984 1071 988 1075
rect 1056 1071 1060 1075
rect 1128 1071 1132 1075
rect 1192 1071 1196 1075
rect 1256 1071 1260 1075
rect 1320 1071 1324 1075
rect 1376 1071 1380 1075
rect 1432 1071 1436 1075
rect 1480 1071 1484 1075
rect 1520 1071 1524 1075
rect 1568 1071 1572 1075
rect 1608 1071 1612 1075
rect 1640 1071 1644 1075
rect 232 1055 236 1059
rect 264 1055 268 1059
rect 296 1055 300 1059
rect 328 1055 332 1059
rect 368 1055 372 1059
rect 408 1055 412 1059
rect 456 1055 460 1059
rect 520 1055 524 1059
rect 592 1055 596 1059
rect 672 1055 676 1059
rect 752 1055 756 1059
rect 832 1055 836 1059
rect 912 1055 916 1059
rect 984 1055 988 1059
rect 1056 1055 1060 1059
rect 1128 1055 1132 1059
rect 1192 1055 1196 1059
rect 1256 1055 1260 1059
rect 1320 1055 1324 1059
rect 1376 1055 1380 1059
rect 1432 1055 1436 1059
rect 1480 1055 1484 1059
rect 1520 1055 1524 1059
rect 1568 1055 1572 1059
rect 1608 1055 1612 1059
rect 1640 1055 1644 1059
rect 528 1035 532 1039
rect 584 1035 588 1039
rect 656 1035 660 1039
rect 824 1035 828 1039
rect 984 1035 988 1039
rect 1056 1035 1060 1039
rect 1120 1035 1124 1039
rect 1184 1035 1188 1039
rect 1248 1035 1252 1039
rect 1360 1035 1364 1039
rect 312 1031 316 1035
rect 344 1031 348 1035
rect 376 1031 380 1035
rect 408 1031 412 1035
rect 440 1031 444 1035
rect 472 1031 476 1035
rect 520 1031 524 1035
rect 576 1031 580 1035
rect 648 1031 652 1035
rect 728 1031 732 1035
rect 816 1031 820 1035
rect 896 1031 900 1035
rect 976 1031 980 1035
rect 1048 1031 1052 1035
rect 1112 1031 1116 1035
rect 1176 1031 1180 1035
rect 1240 1031 1244 1035
rect 1296 1031 1300 1035
rect 1352 1031 1356 1035
rect 1400 1031 1404 1035
rect 1448 1031 1452 1035
rect 1496 1031 1500 1035
rect 1552 1031 1556 1035
rect 1608 1031 1612 1035
rect 1640 1031 1644 1035
rect 312 1015 316 1019
rect 344 1015 348 1019
rect 376 1015 380 1019
rect 408 1015 412 1019
rect 440 1015 444 1019
rect 472 1015 476 1019
rect 520 1015 524 1019
rect 528 1015 532 1019
rect 576 1015 580 1019
rect 584 1015 588 1019
rect 648 1015 652 1019
rect 656 1015 660 1019
rect 728 1015 732 1019
rect 816 1015 820 1019
rect 824 1015 828 1019
rect 896 1015 900 1019
rect 976 1015 980 1019
rect 984 1015 988 1019
rect 1048 1015 1052 1019
rect 1056 1015 1060 1019
rect 1112 1015 1116 1019
rect 1120 1015 1124 1019
rect 1176 1015 1180 1019
rect 1184 1015 1188 1019
rect 1240 1015 1244 1019
rect 1248 1015 1252 1019
rect 1296 1015 1300 1019
rect 1352 1015 1356 1019
rect 1360 1015 1364 1019
rect 1400 1015 1404 1019
rect 1448 1015 1452 1019
rect 1496 1015 1500 1019
rect 1552 1015 1556 1019
rect 1608 1015 1612 1019
rect 1640 1015 1644 1019
rect 264 987 268 991
rect 296 987 300 991
rect 328 987 332 991
rect 360 987 364 991
rect 400 987 404 991
rect 440 987 444 991
rect 496 987 500 991
rect 560 987 564 991
rect 632 987 636 991
rect 704 987 708 991
rect 776 987 780 991
rect 848 987 852 991
rect 920 987 924 991
rect 984 987 988 991
rect 1048 987 1052 991
rect 1112 987 1116 991
rect 1176 987 1180 991
rect 1240 987 1244 991
rect 1304 987 1308 991
rect 1360 987 1364 991
rect 1416 987 1420 991
rect 1464 987 1468 991
rect 1512 987 1516 991
rect 1560 987 1564 991
rect 1608 987 1612 991
rect 1640 987 1644 991
rect 264 971 268 975
rect 296 973 300 977
rect 328 971 332 975
rect 360 971 364 975
rect 400 971 404 975
rect 440 971 444 975
rect 496 971 500 975
rect 560 971 564 975
rect 632 971 636 975
rect 704 971 708 975
rect 776 971 780 975
rect 848 971 852 975
rect 920 971 924 975
rect 984 971 988 975
rect 1048 971 1052 975
rect 1112 971 1116 975
rect 1176 971 1180 975
rect 1240 971 1244 975
rect 1304 971 1308 975
rect 1360 971 1364 975
rect 1416 971 1420 975
rect 1464 971 1468 975
rect 1512 971 1516 975
rect 1560 971 1564 975
rect 1608 971 1612 975
rect 1640 971 1644 975
rect 224 955 228 959
rect 264 955 268 959
rect 312 955 316 959
rect 368 955 372 959
rect 496 955 500 959
rect 560 955 564 959
rect 624 955 628 959
rect 872 955 876 959
rect 936 955 940 959
rect 1000 955 1004 959
rect 1064 955 1068 959
rect 1128 955 1132 959
rect 1416 955 1420 959
rect 184 951 188 955
rect 216 951 220 955
rect 256 951 260 955
rect 304 951 308 955
rect 360 951 364 955
rect 424 951 428 955
rect 488 951 492 955
rect 552 951 556 955
rect 616 951 620 955
rect 680 951 684 955
rect 744 951 748 955
rect 808 951 812 955
rect 864 951 868 955
rect 928 951 932 955
rect 992 951 996 955
rect 1056 951 1060 955
rect 1120 951 1124 955
rect 1184 951 1188 955
rect 1248 951 1252 955
rect 1304 951 1308 955
rect 1360 951 1364 955
rect 1408 951 1412 955
rect 1448 951 1452 955
rect 1488 951 1492 955
rect 1528 951 1532 955
rect 1568 951 1572 955
rect 1608 951 1612 955
rect 1640 951 1644 955
rect 184 935 188 939
rect 216 935 220 939
rect 224 935 228 939
rect 256 935 260 939
rect 264 935 268 939
rect 304 935 308 939
rect 312 935 316 939
rect 360 935 364 939
rect 368 935 372 939
rect 424 935 428 939
rect 488 935 492 939
rect 496 935 500 939
rect 552 935 556 939
rect 560 935 564 939
rect 616 935 620 939
rect 624 935 628 939
rect 680 935 684 939
rect 744 935 748 939
rect 808 935 812 939
rect 864 935 868 939
rect 872 935 876 939
rect 928 935 932 939
rect 936 935 940 939
rect 992 935 996 939
rect 1000 935 1004 939
rect 1056 935 1060 939
rect 1064 935 1068 939
rect 1120 935 1124 939
rect 1128 935 1132 939
rect 1184 935 1188 939
rect 1248 935 1252 939
rect 1304 935 1308 939
rect 1360 935 1364 939
rect 1408 935 1412 939
rect 1416 935 1420 939
rect 1448 937 1452 941
rect 1488 935 1492 939
rect 1528 935 1532 939
rect 1568 935 1572 939
rect 1608 935 1612 939
rect 1640 935 1644 939
rect 152 903 156 907
rect 184 903 188 907
rect 224 903 228 907
rect 288 903 292 907
rect 352 903 356 907
rect 424 903 428 907
rect 488 903 492 907
rect 552 903 556 907
rect 608 903 612 907
rect 664 903 668 907
rect 720 903 724 907
rect 768 903 772 907
rect 816 903 820 907
rect 864 903 868 907
rect 920 903 924 907
rect 976 903 980 907
rect 1040 903 1044 907
rect 1104 903 1108 907
rect 1160 903 1164 907
rect 1216 903 1220 907
rect 1272 903 1276 907
rect 1336 903 1340 907
rect 1400 903 1404 907
rect 152 887 156 891
rect 184 887 188 891
rect 224 887 228 891
rect 288 887 292 891
rect 352 887 356 891
rect 424 887 428 891
rect 488 887 492 891
rect 552 887 556 891
rect 608 887 612 891
rect 664 887 668 891
rect 720 887 724 891
rect 768 887 772 891
rect 816 887 820 891
rect 864 887 868 891
rect 920 887 924 891
rect 976 887 980 891
rect 1040 887 1044 891
rect 1104 887 1108 891
rect 1160 887 1164 891
rect 1216 887 1220 891
rect 1272 887 1276 891
rect 1336 887 1340 891
rect 1400 887 1404 891
rect 192 867 196 871
rect 232 867 236 871
rect 296 867 300 871
rect 360 867 364 871
rect 496 867 500 871
rect 728 867 732 871
rect 1064 867 1068 871
rect 1192 867 1196 871
rect 1256 867 1260 871
rect 1312 867 1316 871
rect 1368 867 1372 871
rect 1424 867 1428 871
rect 152 863 156 867
rect 184 863 188 867
rect 224 863 228 867
rect 288 863 292 867
rect 352 863 356 867
rect 424 863 428 867
rect 488 863 492 867
rect 552 863 556 867
rect 616 863 620 867
rect 672 863 676 867
rect 720 863 724 867
rect 768 863 772 867
rect 816 863 820 867
rect 864 863 868 867
rect 920 863 924 867
rect 984 863 988 867
rect 1056 863 1060 867
rect 1120 863 1124 867
rect 1184 863 1188 867
rect 1248 863 1252 867
rect 1304 863 1308 867
rect 1360 863 1364 867
rect 1416 863 1420 867
rect 1480 863 1484 867
rect 152 847 156 851
rect 184 847 188 851
rect 192 847 196 851
rect 224 847 228 851
rect 232 847 236 851
rect 288 847 292 851
rect 296 847 300 851
rect 352 847 356 851
rect 360 847 364 851
rect 424 847 428 851
rect 488 847 492 851
rect 496 847 500 851
rect 552 847 556 851
rect 616 847 620 851
rect 672 847 676 851
rect 720 847 724 851
rect 728 847 732 851
rect 768 847 772 851
rect 816 847 820 851
rect 864 847 868 851
rect 920 847 924 851
rect 984 847 988 851
rect 1056 847 1060 851
rect 1064 847 1068 851
rect 1120 847 1124 851
rect 1184 847 1188 851
rect 1192 847 1196 851
rect 1248 847 1252 851
rect 1256 847 1260 851
rect 1304 847 1308 851
rect 1312 847 1316 851
rect 1360 847 1364 851
rect 1368 847 1372 851
rect 1416 847 1420 851
rect 1424 847 1428 851
rect 1480 847 1484 851
rect 152 819 156 823
rect 184 819 188 823
rect 232 819 236 823
rect 296 819 300 823
rect 360 819 364 823
rect 432 819 436 823
rect 496 819 500 823
rect 560 819 564 823
rect 624 819 628 823
rect 688 819 692 823
rect 752 819 756 823
rect 808 819 812 823
rect 864 819 868 823
rect 928 819 932 823
rect 992 819 996 823
rect 1056 819 1060 823
rect 1064 819 1068 823
rect 1128 819 1132 823
rect 1200 819 1204 823
rect 1264 819 1268 823
rect 1328 819 1332 823
rect 1384 819 1388 823
rect 1440 819 1444 823
rect 1496 819 1500 823
rect 1552 819 1556 823
rect 1608 819 1612 823
rect 152 803 156 807
rect 184 803 188 807
rect 232 803 236 807
rect 296 803 300 807
rect 360 803 364 807
rect 432 803 436 807
rect 496 803 500 807
rect 560 803 564 807
rect 624 803 628 807
rect 688 803 692 807
rect 752 803 756 807
rect 808 803 812 807
rect 864 803 868 807
rect 928 803 932 807
rect 992 803 996 807
rect 1056 803 1060 807
rect 1128 803 1132 807
rect 1200 803 1204 807
rect 1264 803 1268 807
rect 1328 803 1332 807
rect 1384 803 1388 807
rect 1440 803 1444 807
rect 1496 803 1500 807
rect 1552 803 1556 807
rect 1608 803 1612 807
rect 1064 795 1068 799
rect 160 783 164 787
rect 200 783 204 787
rect 392 783 396 787
rect 552 783 556 787
rect 728 783 732 787
rect 816 783 820 787
rect 976 783 980 787
rect 1048 783 1052 787
rect 1120 783 1124 787
rect 1192 783 1196 787
rect 1256 783 1260 787
rect 1384 783 1388 787
rect 1440 783 1444 787
rect 152 779 156 783
rect 192 779 196 783
rect 248 779 252 783
rect 312 779 316 783
rect 384 779 388 783
rect 464 779 468 783
rect 544 779 548 783
rect 632 779 636 783
rect 720 779 724 783
rect 808 779 812 783
rect 888 779 892 783
rect 968 779 972 783
rect 1040 779 1044 783
rect 1112 779 1116 783
rect 1184 779 1188 783
rect 1248 779 1252 783
rect 1312 779 1316 783
rect 1376 779 1380 783
rect 1432 779 1436 783
rect 1488 779 1492 783
rect 1544 779 1548 783
rect 1608 779 1612 783
rect 152 763 156 767
rect 160 763 164 767
rect 192 763 196 767
rect 200 763 204 767
rect 248 763 252 767
rect 312 763 316 767
rect 384 763 388 767
rect 392 763 396 767
rect 464 763 468 767
rect 544 763 548 767
rect 552 763 556 767
rect 632 763 636 767
rect 720 763 724 767
rect 728 763 732 767
rect 808 763 812 767
rect 816 763 820 767
rect 888 763 892 767
rect 968 763 972 767
rect 976 763 980 767
rect 1040 763 1044 767
rect 1048 763 1052 767
rect 1112 763 1116 767
rect 1120 763 1124 767
rect 1184 763 1188 767
rect 1192 763 1196 767
rect 1248 763 1252 767
rect 1256 763 1260 767
rect 1312 763 1316 767
rect 1376 763 1380 767
rect 1384 763 1388 767
rect 1432 763 1436 767
rect 1440 763 1444 767
rect 1488 763 1492 767
rect 1544 763 1548 767
rect 1608 763 1612 767
rect 232 735 236 739
rect 264 735 268 739
rect 296 737 300 741
rect 336 735 340 739
rect 376 735 380 739
rect 416 735 420 739
rect 456 735 460 739
rect 464 735 468 739
rect 504 735 508 739
rect 560 735 564 739
rect 624 735 628 739
rect 688 735 692 739
rect 752 735 756 739
rect 816 735 820 739
rect 880 735 884 739
rect 944 735 948 739
rect 1008 735 1012 739
rect 1072 735 1076 739
rect 1136 735 1140 739
rect 1200 735 1204 739
rect 1208 735 1212 739
rect 1256 735 1260 739
rect 1312 735 1316 739
rect 1368 735 1372 739
rect 1424 735 1428 739
rect 1480 735 1484 739
rect 1536 735 1540 739
rect 1600 735 1604 739
rect 1640 735 1644 739
rect 232 719 236 723
rect 264 719 268 723
rect 296 719 300 723
rect 336 719 340 723
rect 376 719 380 723
rect 416 719 420 723
rect 456 719 460 723
rect 504 719 508 723
rect 560 719 564 723
rect 624 719 628 723
rect 688 719 692 723
rect 752 719 756 723
rect 816 719 820 723
rect 880 719 884 723
rect 944 719 948 723
rect 1008 719 1012 723
rect 1072 719 1076 723
rect 1136 719 1140 723
rect 1200 719 1204 723
rect 464 699 468 703
rect 528 699 532 703
rect 568 699 572 703
rect 616 699 620 703
rect 672 699 676 703
rect 784 699 788 703
rect 848 699 852 703
rect 1048 699 1052 703
rect 1184 699 1188 703
rect 296 695 300 699
rect 328 695 332 699
rect 360 695 364 699
rect 392 695 396 699
rect 424 695 428 699
rect 456 695 460 699
rect 488 695 492 699
rect 520 695 524 699
rect 560 695 564 699
rect 608 695 612 699
rect 664 695 668 699
rect 720 695 724 699
rect 776 695 780 699
rect 840 695 844 699
rect 904 695 908 699
rect 976 695 980 699
rect 1040 695 1044 699
rect 1104 695 1108 699
rect 1176 695 1180 699
rect 1256 719 1260 723
rect 1312 719 1316 723
rect 1368 719 1372 723
rect 1424 719 1428 723
rect 1480 719 1484 723
rect 1536 719 1540 723
rect 1600 719 1604 723
rect 1640 719 1644 723
rect 1248 699 1252 703
rect 1312 699 1316 703
rect 1376 699 1380 703
rect 1496 699 1500 703
rect 1608 699 1612 703
rect 1240 695 1244 699
rect 1208 691 1212 695
rect 1304 695 1308 699
rect 1368 695 1372 699
rect 1432 695 1436 699
rect 1488 695 1492 699
rect 1544 695 1548 699
rect 1600 695 1604 699
rect 1640 695 1644 699
rect 296 679 300 683
rect 328 679 332 683
rect 360 679 364 683
rect 392 679 396 683
rect 424 679 428 683
rect 456 679 460 683
rect 488 679 492 683
rect 520 679 524 683
rect 528 679 532 683
rect 560 679 564 683
rect 568 679 572 683
rect 608 679 612 683
rect 616 679 620 683
rect 664 679 668 683
rect 672 679 676 683
rect 720 679 724 683
rect 776 679 780 683
rect 784 679 788 683
rect 840 679 844 683
rect 848 679 852 683
rect 904 679 908 683
rect 976 679 980 683
rect 1040 679 1044 683
rect 1048 679 1052 683
rect 1104 679 1108 683
rect 1176 679 1180 683
rect 1184 679 1188 683
rect 1240 679 1244 683
rect 1248 679 1252 683
rect 1304 679 1308 683
rect 1312 679 1316 683
rect 1368 679 1372 683
rect 1376 679 1380 683
rect 1432 679 1436 683
rect 1488 679 1492 683
rect 1496 679 1500 683
rect 1544 679 1548 683
rect 1600 679 1604 683
rect 1608 679 1612 683
rect 1640 679 1644 683
rect 312 651 316 655
rect 344 651 348 655
rect 376 651 380 655
rect 408 651 412 655
rect 440 651 444 655
rect 472 651 476 655
rect 504 651 508 655
rect 536 651 540 655
rect 568 651 572 655
rect 608 651 612 655
rect 656 651 660 655
rect 704 651 708 655
rect 752 651 756 655
rect 808 651 812 655
rect 864 651 868 655
rect 928 651 932 655
rect 992 651 996 655
rect 1064 651 1068 655
rect 1144 651 1148 655
rect 1232 651 1236 655
rect 1312 651 1316 655
rect 1400 651 1404 655
rect 1488 651 1492 655
rect 1576 651 1580 655
rect 1640 651 1644 655
rect 1648 651 1652 655
rect 312 635 316 639
rect 344 635 348 639
rect 376 635 380 639
rect 408 635 412 639
rect 440 635 444 639
rect 472 635 476 639
rect 504 635 508 639
rect 536 635 540 639
rect 568 635 572 639
rect 608 635 612 639
rect 656 635 660 639
rect 704 635 708 639
rect 752 635 756 639
rect 808 635 812 639
rect 864 635 868 639
rect 928 635 932 639
rect 992 635 996 639
rect 1064 635 1068 639
rect 1144 635 1148 639
rect 1232 635 1236 639
rect 1312 635 1316 639
rect 1400 635 1404 639
rect 1488 635 1492 639
rect 1576 635 1580 639
rect 1640 635 1644 639
rect 304 619 308 623
rect 352 619 356 623
rect 392 619 396 623
rect 448 619 452 623
rect 544 619 548 623
rect 592 619 596 623
rect 640 619 644 623
rect 688 619 692 623
rect 744 619 748 623
rect 856 619 860 623
rect 920 619 924 623
rect 1072 619 1076 623
rect 1384 619 1388 623
rect 1456 619 1460 623
rect 1528 619 1532 623
rect 264 615 268 619
rect 296 615 300 619
rect 336 615 340 619
rect 384 615 388 619
rect 440 615 444 619
rect 488 615 492 619
rect 536 615 540 619
rect 584 615 588 619
rect 632 615 636 619
rect 680 615 684 619
rect 736 615 740 619
rect 792 615 796 619
rect 848 615 852 619
rect 912 615 916 619
rect 984 615 988 619
rect 1064 615 1068 619
rect 1144 615 1148 619
rect 1224 615 1228 619
rect 1304 615 1308 619
rect 1376 615 1380 619
rect 1448 615 1452 619
rect 1520 615 1524 619
rect 1592 615 1596 619
rect 1640 615 1644 619
rect 1648 615 1652 619
rect 264 599 268 603
rect 296 599 300 603
rect 304 599 308 603
rect 336 599 340 603
rect 352 599 356 603
rect 384 599 388 603
rect 392 599 396 603
rect 440 599 444 603
rect 448 599 452 603
rect 488 599 492 603
rect 536 599 540 603
rect 544 599 548 603
rect 584 599 588 603
rect 592 599 596 603
rect 632 599 636 603
rect 640 599 644 603
rect 680 599 684 603
rect 688 599 692 603
rect 736 599 740 603
rect 744 599 748 603
rect 792 599 796 603
rect 848 599 852 603
rect 856 599 860 603
rect 912 599 916 603
rect 920 599 924 603
rect 984 599 988 603
rect 1064 599 1068 603
rect 1072 599 1076 603
rect 1144 599 1148 603
rect 1224 599 1228 603
rect 1304 599 1308 603
rect 1376 599 1380 603
rect 1384 599 1388 603
rect 1448 599 1452 603
rect 1456 599 1460 603
rect 1520 599 1524 603
rect 1528 599 1532 603
rect 1592 599 1596 603
rect 1640 599 1644 603
rect 184 571 188 575
rect 232 571 236 575
rect 288 571 292 575
rect 352 571 356 575
rect 424 571 428 575
rect 504 571 508 575
rect 576 571 580 575
rect 648 571 652 575
rect 720 571 724 575
rect 784 571 788 575
rect 840 571 844 575
rect 896 571 900 575
rect 904 571 908 575
rect 952 571 956 575
rect 1008 571 1012 575
rect 1064 571 1068 575
rect 1120 571 1124 575
rect 1176 571 1180 575
rect 1232 571 1236 575
rect 1288 571 1292 575
rect 1344 571 1348 575
rect 1400 571 1404 575
rect 1464 571 1468 575
rect 1528 571 1532 575
rect 1592 571 1596 575
rect 1640 571 1644 575
rect 1648 571 1652 575
rect 184 555 188 559
rect 232 555 236 559
rect 288 555 292 559
rect 352 555 356 559
rect 424 555 428 559
rect 504 555 508 559
rect 576 555 580 559
rect 648 555 652 559
rect 720 555 724 559
rect 784 555 788 559
rect 840 555 844 559
rect 896 555 900 559
rect 952 555 956 559
rect 1008 555 1012 559
rect 1064 555 1068 559
rect 1120 555 1124 559
rect 1176 555 1180 559
rect 1232 555 1236 559
rect 1288 555 1292 559
rect 1344 555 1348 559
rect 1400 555 1404 559
rect 1464 555 1468 559
rect 1528 555 1532 559
rect 1592 555 1596 559
rect 1640 555 1644 559
rect 904 547 908 551
rect 256 535 260 539
rect 304 535 308 539
rect 400 535 404 539
rect 712 535 716 539
rect 904 535 908 539
rect 968 535 972 539
rect 1256 535 1260 539
rect 1304 535 1308 539
rect 1360 535 1364 539
rect 1416 535 1420 539
rect 1472 535 1476 539
rect 152 531 156 535
rect 184 531 188 535
rect 216 531 220 535
rect 248 531 252 535
rect 296 531 300 535
rect 344 531 348 535
rect 392 531 396 535
rect 448 531 452 535
rect 512 531 516 535
rect 576 531 580 535
rect 640 531 644 535
rect 704 531 708 535
rect 768 531 772 535
rect 832 531 836 535
rect 896 531 900 535
rect 960 531 964 535
rect 1024 531 1028 535
rect 1088 531 1092 535
rect 1144 531 1148 535
rect 1200 531 1204 535
rect 1248 531 1252 535
rect 1296 531 1300 535
rect 1352 531 1356 535
rect 1408 531 1412 535
rect 1464 531 1468 535
rect 1528 531 1532 535
rect 1592 531 1596 535
rect 1640 531 1644 535
rect 1648 531 1652 535
rect 152 515 156 519
rect 184 515 188 519
rect 216 515 220 519
rect 248 515 252 519
rect 256 515 260 519
rect 296 515 300 519
rect 304 515 308 519
rect 344 515 348 519
rect 392 515 396 519
rect 400 515 404 519
rect 448 515 452 519
rect 512 515 516 519
rect 576 515 580 519
rect 640 515 644 519
rect 704 515 708 519
rect 712 515 716 519
rect 768 515 772 519
rect 832 515 836 519
rect 896 515 900 519
rect 904 515 908 519
rect 960 515 964 519
rect 968 515 972 519
rect 1024 515 1028 519
rect 1088 515 1092 519
rect 1144 515 1148 519
rect 1200 515 1204 519
rect 1248 515 1252 519
rect 1256 515 1260 519
rect 1296 515 1300 519
rect 1304 515 1308 519
rect 1352 515 1356 519
rect 1360 515 1364 519
rect 1408 515 1412 519
rect 1416 515 1420 519
rect 1464 515 1468 519
rect 1472 515 1476 519
rect 1528 515 1532 519
rect 1592 515 1596 519
rect 1640 515 1644 519
rect 152 487 156 491
rect 184 487 188 491
rect 216 487 220 491
rect 256 487 260 491
rect 264 487 268 491
rect 304 487 308 491
rect 344 487 348 491
rect 360 487 364 491
rect 392 487 396 491
rect 440 487 444 491
rect 496 487 500 491
rect 560 487 564 491
rect 632 487 636 491
rect 640 487 644 491
rect 712 487 716 491
rect 792 487 796 491
rect 864 487 868 491
rect 936 487 940 491
rect 1000 487 1004 491
rect 1056 487 1060 491
rect 1112 487 1116 491
rect 1160 487 1164 491
rect 1208 487 1212 491
rect 1256 487 1260 491
rect 1304 487 1308 491
rect 1352 487 1356 491
rect 1400 489 1404 493
rect 1448 487 1452 491
rect 1496 487 1500 491
rect 1552 487 1556 491
rect 1608 487 1612 491
rect 1640 487 1644 491
rect 152 471 156 475
rect 184 471 188 475
rect 216 471 220 475
rect 256 471 260 475
rect 304 471 308 475
rect 344 471 348 475
rect 264 463 268 467
rect 392 471 396 475
rect 440 471 444 475
rect 496 471 500 475
rect 560 471 564 475
rect 632 471 636 475
rect 712 471 716 475
rect 792 471 796 475
rect 864 471 868 475
rect 936 471 940 475
rect 1000 471 1004 475
rect 1056 471 1060 475
rect 1112 471 1116 475
rect 1160 471 1164 475
rect 1208 471 1212 475
rect 1256 471 1260 475
rect 1304 471 1308 475
rect 1352 471 1356 475
rect 1400 471 1404 475
rect 1448 471 1452 475
rect 1496 471 1500 475
rect 1552 471 1556 475
rect 1608 471 1612 475
rect 1640 471 1644 475
rect 640 463 644 467
rect 232 455 236 459
rect 360 455 364 459
rect 392 455 396 459
rect 512 455 516 459
rect 544 455 548 459
rect 624 455 628 459
rect 864 455 868 459
rect 1288 455 1292 459
rect 168 451 172 455
rect 224 451 228 455
rect 272 451 276 455
rect 328 451 332 455
rect 352 451 356 455
rect 384 451 388 455
rect 168 435 172 439
rect 224 435 228 439
rect 232 435 236 439
rect 272 435 276 439
rect 328 435 332 439
rect 456 451 460 455
rect 384 435 388 439
rect 392 435 396 439
rect 456 435 460 439
rect 352 423 356 427
rect 536 451 540 455
rect 616 451 620 455
rect 696 451 700 455
rect 776 451 780 455
rect 856 451 860 455
rect 928 451 932 455
rect 1000 451 1004 455
rect 1072 451 1076 455
rect 1144 451 1148 455
rect 1216 451 1220 455
rect 1280 451 1284 455
rect 1336 451 1340 455
rect 1392 451 1396 455
rect 1448 451 1452 455
rect 1512 451 1516 455
rect 536 435 540 439
rect 544 435 548 439
rect 616 435 620 439
rect 624 435 628 439
rect 696 435 700 439
rect 776 435 780 439
rect 856 435 860 439
rect 864 435 868 439
rect 928 435 932 439
rect 1000 435 1004 439
rect 1072 435 1076 439
rect 1144 435 1148 439
rect 1216 435 1220 439
rect 1280 435 1284 439
rect 1288 435 1292 439
rect 1336 435 1340 439
rect 1392 435 1396 439
rect 1448 435 1452 439
rect 1512 435 1516 439
rect 192 407 196 411
rect 240 407 244 411
rect 288 407 292 411
rect 336 407 340 411
rect 384 407 388 411
rect 432 407 436 411
rect 488 407 492 411
rect 512 407 516 411
rect 544 407 548 411
rect 608 407 612 411
rect 680 407 684 411
rect 752 407 756 411
rect 824 407 828 411
rect 888 407 892 411
rect 952 407 956 411
rect 1008 407 1012 411
rect 1056 407 1060 411
rect 1104 407 1108 411
rect 1144 407 1148 411
rect 1184 407 1188 411
rect 1192 407 1196 411
rect 1224 407 1228 411
rect 1264 407 1268 411
rect 1304 407 1308 411
rect 1352 407 1356 411
rect 1400 407 1404 411
rect 1408 407 1412 411
rect 192 391 196 395
rect 240 391 244 395
rect 288 391 292 395
rect 336 391 340 395
rect 384 391 388 395
rect 432 391 436 395
rect 488 391 492 395
rect 544 391 548 395
rect 608 391 612 395
rect 680 391 684 395
rect 752 391 756 395
rect 824 391 828 395
rect 888 391 892 395
rect 952 391 956 395
rect 1008 391 1012 395
rect 1056 391 1060 395
rect 1104 391 1108 395
rect 1144 391 1148 395
rect 1184 391 1188 395
rect 1224 391 1228 395
rect 1264 391 1268 395
rect 1304 391 1308 395
rect 1352 391 1356 395
rect 1400 391 1404 395
rect 1408 383 1412 387
rect 488 371 492 375
rect 544 371 548 375
rect 600 371 604 375
rect 768 371 772 375
rect 944 371 948 375
rect 1008 371 1012 375
rect 1192 371 1196 375
rect 1280 371 1284 375
rect 1328 371 1332 375
rect 1376 371 1380 375
rect 1520 371 1524 375
rect 1568 371 1572 375
rect 152 367 156 371
rect 184 367 188 371
rect 216 367 220 371
rect 256 367 260 371
rect 312 367 316 371
rect 368 367 372 371
rect 424 367 428 371
rect 480 367 484 371
rect 536 367 540 371
rect 592 367 596 371
rect 648 367 652 371
rect 704 367 708 371
rect 760 367 764 371
rect 816 367 820 371
rect 872 367 876 371
rect 936 367 940 371
rect 1000 367 1004 371
rect 1056 367 1060 371
rect 1112 367 1116 371
rect 1168 367 1172 371
rect 1224 367 1228 371
rect 1272 367 1276 371
rect 1320 367 1324 371
rect 1368 367 1372 371
rect 1416 367 1420 371
rect 1464 367 1468 371
rect 1512 367 1516 371
rect 1560 367 1564 371
rect 1608 367 1612 371
rect 1640 367 1644 371
rect 152 351 156 355
rect 184 351 188 355
rect 216 351 220 355
rect 256 351 260 355
rect 312 351 316 355
rect 368 351 372 355
rect 424 351 428 355
rect 480 351 484 355
rect 488 351 492 355
rect 536 351 540 355
rect 544 351 548 355
rect 592 351 596 355
rect 600 351 604 355
rect 648 351 652 355
rect 704 351 708 355
rect 760 351 764 355
rect 768 351 772 355
rect 816 351 820 355
rect 872 351 876 355
rect 936 351 940 355
rect 944 351 948 355
rect 1000 351 1004 355
rect 1008 351 1012 355
rect 1056 351 1060 355
rect 1112 351 1116 355
rect 1168 351 1172 355
rect 1224 351 1228 355
rect 1272 351 1276 355
rect 1280 351 1284 355
rect 1320 351 1324 355
rect 1328 351 1332 355
rect 1368 351 1372 355
rect 1376 351 1380 355
rect 1416 351 1420 355
rect 1464 351 1468 355
rect 1512 351 1516 355
rect 1520 351 1524 355
rect 1560 351 1564 355
rect 1568 351 1572 355
rect 1608 351 1612 355
rect 1640 351 1644 355
rect 1368 339 1372 343
rect 152 323 156 327
rect 184 323 188 327
rect 224 323 228 327
rect 280 323 284 327
rect 344 323 348 327
rect 408 323 412 327
rect 472 323 476 327
rect 536 323 540 327
rect 592 323 596 327
rect 648 323 652 327
rect 656 323 660 327
rect 704 323 708 327
rect 768 323 772 327
rect 776 323 780 327
rect 832 323 836 327
rect 896 323 900 327
rect 968 323 972 327
rect 1048 323 1052 327
rect 1128 323 1132 327
rect 1208 323 1212 327
rect 1288 323 1292 327
rect 1360 323 1364 327
rect 152 307 156 311
rect 184 307 188 311
rect 224 307 228 311
rect 280 307 284 311
rect 344 307 348 311
rect 408 307 412 311
rect 472 307 476 311
rect 536 307 540 311
rect 592 307 596 311
rect 648 307 652 311
rect 704 307 708 311
rect 768 307 772 311
rect 656 299 660 303
rect 1424 323 1428 327
rect 1480 323 1484 327
rect 1536 323 1540 327
rect 1600 323 1604 327
rect 1640 323 1644 327
rect 1648 323 1652 327
rect 832 307 836 311
rect 896 307 900 311
rect 968 307 972 311
rect 1048 307 1052 311
rect 1128 307 1132 311
rect 1208 307 1212 311
rect 1288 307 1292 311
rect 1360 307 1364 311
rect 1368 307 1372 311
rect 1424 307 1428 311
rect 1480 307 1484 311
rect 1536 307 1540 311
rect 1600 307 1604 311
rect 1640 307 1644 311
rect 152 287 156 291
rect 184 287 188 291
rect 248 287 252 291
rect 312 287 316 291
rect 384 287 388 291
rect 456 287 460 291
rect 520 287 524 291
rect 584 287 588 291
rect 648 287 652 291
rect 704 287 708 291
rect 760 287 764 291
rect 776 287 780 291
rect 784 291 788 295
rect 832 291 836 295
rect 904 291 908 295
rect 976 291 980 295
rect 1136 291 1140 295
rect 1216 291 1220 295
rect 1352 291 1356 295
rect 824 287 828 291
rect 896 287 900 291
rect 968 287 972 291
rect 1048 287 1052 291
rect 1128 287 1132 291
rect 1208 287 1212 291
rect 1280 287 1284 291
rect 1344 287 1348 291
rect 1408 287 1412 291
rect 1464 287 1468 291
rect 1512 287 1516 291
rect 1560 287 1564 291
rect 1608 287 1612 291
rect 1640 287 1644 291
rect 1648 287 1652 291
rect 152 271 156 275
rect 184 271 188 275
rect 248 271 252 275
rect 312 271 316 275
rect 384 271 388 275
rect 456 271 460 275
rect 520 271 524 275
rect 584 271 588 275
rect 648 271 652 275
rect 704 271 708 275
rect 760 271 764 275
rect 784 271 788 275
rect 824 271 828 275
rect 832 271 836 275
rect 896 271 900 275
rect 904 271 908 275
rect 968 271 972 275
rect 976 271 980 275
rect 1048 271 1052 275
rect 1128 271 1132 275
rect 1136 271 1140 275
rect 1208 271 1212 275
rect 1216 271 1220 275
rect 1280 271 1284 275
rect 1344 271 1348 275
rect 1352 271 1356 275
rect 1408 271 1412 275
rect 1464 271 1468 275
rect 1512 271 1516 275
rect 1560 271 1564 275
rect 1608 271 1612 275
rect 1640 271 1644 275
rect 152 239 156 243
rect 192 239 196 243
rect 264 239 268 243
rect 336 239 340 243
rect 400 239 404 243
rect 464 239 468 243
rect 536 239 540 243
rect 608 239 612 243
rect 680 239 684 243
rect 760 239 764 243
rect 840 239 844 243
rect 912 239 916 243
rect 984 239 988 243
rect 1048 239 1052 243
rect 1104 239 1108 243
rect 1160 239 1164 243
rect 1216 239 1220 243
rect 1272 239 1276 243
rect 1328 239 1332 243
rect 1384 239 1388 243
rect 1432 239 1436 243
rect 1480 239 1484 243
rect 1536 239 1540 243
rect 1592 239 1596 243
rect 1640 239 1644 243
rect 152 223 156 227
rect 192 223 196 227
rect 264 223 268 227
rect 336 223 340 227
rect 400 223 404 227
rect 464 223 468 227
rect 536 223 540 227
rect 608 223 612 227
rect 680 223 684 227
rect 760 223 764 227
rect 840 223 844 227
rect 912 223 916 227
rect 984 223 988 227
rect 1048 223 1052 227
rect 1104 223 1108 227
rect 1160 223 1164 227
rect 1216 223 1220 227
rect 1272 223 1276 227
rect 1328 223 1332 227
rect 1384 223 1388 227
rect 1432 223 1436 227
rect 1480 223 1484 227
rect 1536 223 1540 227
rect 1592 223 1596 227
rect 1640 223 1644 227
rect 400 207 404 211
rect 440 207 444 211
rect 640 207 644 211
rect 720 207 724 211
rect 880 207 884 211
rect 952 207 956 211
rect 1024 207 1028 211
rect 1096 207 1100 211
rect 1168 207 1172 211
rect 1552 207 1556 211
rect 1608 207 1612 211
rect 152 203 156 207
rect 184 203 188 207
rect 224 203 228 207
rect 272 203 276 207
rect 320 203 324 207
rect 360 203 364 207
rect 392 203 396 207
rect 432 203 436 207
rect 488 203 492 207
rect 552 203 556 207
rect 632 203 636 207
rect 712 203 716 207
rect 792 203 796 207
rect 872 203 876 207
rect 944 203 948 207
rect 1016 203 1020 207
rect 1088 203 1092 207
rect 1160 203 1164 207
rect 1232 203 1236 207
rect 1304 203 1308 207
rect 1368 203 1372 207
rect 1432 203 1436 207
rect 1488 203 1492 207
rect 1544 203 1548 207
rect 1600 203 1604 207
rect 1640 203 1644 207
rect 152 187 156 191
rect 184 187 188 191
rect 224 187 228 191
rect 272 187 276 191
rect 320 187 324 191
rect 360 187 364 191
rect 392 187 396 191
rect 400 187 404 191
rect 432 187 436 191
rect 440 187 444 191
rect 488 187 492 191
rect 552 187 556 191
rect 632 187 636 191
rect 640 187 644 191
rect 712 187 716 191
rect 720 187 724 191
rect 792 187 796 191
rect 872 187 876 191
rect 880 187 884 191
rect 944 187 948 191
rect 952 187 956 191
rect 1016 187 1020 191
rect 1024 187 1028 191
rect 1088 187 1092 191
rect 1096 187 1100 191
rect 1160 187 1164 191
rect 1168 187 1172 191
rect 1232 187 1236 191
rect 1304 187 1308 191
rect 1368 187 1372 191
rect 1432 187 1436 191
rect 1488 187 1492 191
rect 1544 187 1548 191
rect 1552 187 1556 191
rect 1600 187 1604 191
rect 1608 187 1612 191
rect 1640 187 1644 191
rect 152 159 156 163
rect 192 159 196 163
rect 248 159 252 163
rect 304 159 308 163
rect 360 159 364 163
rect 416 159 420 163
rect 472 159 476 163
rect 528 159 532 163
rect 592 159 596 163
rect 656 159 660 163
rect 720 159 724 163
rect 784 159 788 163
rect 848 159 852 163
rect 912 159 916 163
rect 968 159 972 163
rect 1032 159 1036 163
rect 1096 159 1100 163
rect 1160 159 1164 163
rect 1224 159 1228 163
rect 1296 159 1300 163
rect 1368 159 1372 163
rect 1440 159 1444 163
rect 1512 159 1516 163
rect 1584 159 1588 163
rect 1640 159 1644 163
rect 1648 159 1652 163
rect 152 143 156 147
rect 192 143 196 147
rect 248 143 252 147
rect 304 143 308 147
rect 360 143 364 147
rect 416 143 420 147
rect 472 143 476 147
rect 528 143 532 147
rect 592 143 596 147
rect 656 143 660 147
rect 720 143 724 147
rect 784 143 788 147
rect 848 143 852 147
rect 912 143 916 147
rect 968 143 972 147
rect 1032 143 1036 147
rect 1096 143 1100 147
rect 1160 143 1164 147
rect 1224 143 1228 147
rect 1296 143 1300 147
rect 1368 143 1372 147
rect 1440 143 1444 147
rect 1512 143 1516 147
rect 1584 143 1588 147
rect 1640 143 1644 147
rect 488 111 492 115
rect 528 111 532 115
rect 920 111 924 115
rect 960 111 964 115
rect 1000 111 1004 115
rect 1040 111 1044 115
rect 1088 111 1092 115
rect 1128 111 1132 115
rect 1208 111 1212 115
rect 1248 111 1252 115
rect 1320 111 1324 115
rect 1360 111 1364 115
rect 1400 111 1404 115
rect 1440 111 1444 115
rect 1480 111 1484 115
rect 1528 111 1532 115
rect 152 107 156 111
rect 184 107 188 111
rect 216 107 220 111
rect 248 107 252 111
rect 280 107 284 111
rect 312 107 316 111
rect 344 107 348 111
rect 376 107 380 111
rect 408 107 412 111
rect 440 107 444 111
rect 480 107 484 111
rect 520 107 524 111
rect 560 107 564 111
rect 592 107 596 111
rect 624 107 628 111
rect 656 107 660 111
rect 688 107 692 111
rect 720 107 724 111
rect 752 107 756 111
rect 784 107 788 111
rect 816 107 820 111
rect 848 107 852 111
rect 880 107 884 111
rect 912 107 916 111
rect 952 107 956 111
rect 992 107 996 111
rect 1032 107 1036 111
rect 1080 107 1084 111
rect 1120 107 1124 111
rect 1160 107 1164 111
rect 1200 107 1204 111
rect 1240 107 1244 111
rect 1280 107 1284 111
rect 1312 107 1316 111
rect 1352 107 1356 111
rect 1392 107 1396 111
rect 1432 107 1436 111
rect 1472 107 1476 111
rect 1520 107 1524 111
rect 1568 107 1572 111
rect 1608 107 1612 111
rect 1640 107 1644 111
rect 1648 107 1652 111
rect 152 91 156 95
rect 184 91 188 95
rect 216 91 220 95
rect 248 91 252 95
rect 280 91 284 95
rect 312 91 316 95
rect 344 91 348 95
rect 376 91 380 95
rect 408 91 412 95
rect 440 91 444 95
rect 480 91 484 95
rect 488 91 492 95
rect 520 91 524 95
rect 528 91 532 95
rect 560 91 564 95
rect 592 91 596 95
rect 624 91 628 95
rect 656 91 660 95
rect 688 91 692 95
rect 720 91 724 95
rect 752 91 756 95
rect 784 91 788 95
rect 816 91 820 95
rect 848 91 852 95
rect 880 91 884 95
rect 912 91 916 95
rect 920 91 924 95
rect 952 91 956 95
rect 960 91 964 95
rect 992 91 996 95
rect 1000 91 1004 95
rect 1032 91 1036 95
rect 1040 91 1044 95
rect 1080 91 1084 95
rect 1088 91 1092 95
rect 1120 91 1124 95
rect 1128 91 1132 95
rect 1160 91 1164 95
rect 1200 91 1204 95
rect 1208 91 1212 95
rect 1240 91 1244 95
rect 1248 91 1252 95
rect 1280 91 1284 95
rect 1312 91 1316 95
rect 1320 91 1324 95
rect 1352 91 1356 95
rect 1360 91 1364 95
rect 1392 91 1396 95
rect 1400 91 1404 95
rect 1432 91 1436 95
rect 1440 91 1444 95
rect 1472 91 1476 95
rect 1480 91 1484 95
rect 1520 91 1524 95
rect 1528 91 1532 95
rect 1568 91 1572 95
rect 1640 91 1644 95
<< m2 >>
rect 374 1715 380 1716
rect 374 1714 375 1715
rect 276 1712 375 1714
rect 276 1708 278 1712
rect 374 1711 375 1712
rect 379 1711 380 1715
rect 1138 1715 1144 1716
rect 374 1710 380 1711
rect 470 1711 476 1712
rect 470 1710 471 1711
rect 271 1707 278 1708
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 271 1703 272 1707
rect 276 1704 278 1707
rect 280 1708 307 1710
rect 400 1708 418 1710
rect 425 1708 471 1710
rect 276 1703 277 1704
rect 110 1699 116 1700
rect 254 1702 260 1703
rect 271 1702 277 1703
rect 254 1698 255 1702
rect 259 1698 260 1702
rect 254 1697 260 1698
rect 271 1691 277 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 271 1687 272 1691
rect 276 1690 277 1691
rect 280 1690 282 1708
rect 303 1707 309 1708
rect 303 1703 304 1707
rect 308 1703 309 1707
rect 335 1707 341 1708
rect 335 1706 336 1707
rect 328 1704 336 1706
rect 286 1702 292 1703
rect 303 1702 309 1703
rect 318 1702 324 1703
rect 286 1698 287 1702
rect 291 1698 292 1702
rect 286 1697 292 1698
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 328 1692 330 1704
rect 335 1703 336 1704
rect 340 1703 341 1707
rect 375 1707 381 1708
rect 375 1703 376 1707
rect 380 1706 381 1707
rect 400 1706 402 1708
rect 380 1704 402 1706
rect 380 1703 381 1704
rect 335 1702 341 1703
rect 358 1702 364 1703
rect 375 1702 381 1703
rect 406 1702 412 1703
rect 358 1698 359 1702
rect 363 1698 364 1702
rect 358 1697 364 1698
rect 406 1698 407 1702
rect 411 1698 412 1702
rect 406 1697 412 1698
rect 416 1694 418 1708
rect 423 1707 429 1708
rect 423 1703 424 1707
rect 428 1703 429 1707
rect 470 1707 471 1708
rect 475 1707 476 1711
rect 538 1711 544 1712
rect 470 1706 476 1707
rect 514 1707 525 1708
rect 514 1703 515 1707
rect 519 1703 520 1707
rect 524 1703 525 1707
rect 538 1707 539 1711
rect 543 1710 544 1711
rect 575 1711 581 1712
rect 543 1708 562 1710
rect 543 1707 544 1708
rect 538 1706 544 1707
rect 560 1706 562 1708
rect 567 1707 573 1708
rect 567 1706 568 1707
rect 560 1704 568 1706
rect 567 1703 568 1704
rect 572 1703 573 1707
rect 575 1707 576 1711
rect 580 1710 581 1711
rect 631 1711 637 1712
rect 580 1708 627 1710
rect 580 1707 581 1708
rect 575 1706 581 1707
rect 623 1707 629 1708
rect 623 1703 624 1707
rect 628 1703 629 1707
rect 631 1707 632 1711
rect 636 1710 637 1711
rect 687 1711 693 1712
rect 636 1708 683 1710
rect 636 1707 637 1708
rect 631 1706 637 1707
rect 679 1707 685 1708
rect 679 1703 680 1707
rect 684 1703 685 1707
rect 687 1707 688 1711
rect 692 1710 693 1711
rect 751 1711 757 1712
rect 692 1708 747 1710
rect 692 1707 693 1708
rect 687 1706 693 1707
rect 743 1707 749 1708
rect 743 1703 744 1707
rect 748 1703 749 1707
rect 751 1707 752 1711
rect 756 1710 757 1711
rect 919 1711 925 1712
rect 756 1708 803 1710
rect 756 1707 757 1708
rect 751 1706 757 1707
rect 799 1707 805 1708
rect 799 1703 800 1707
rect 804 1703 805 1707
rect 855 1707 861 1708
rect 855 1703 856 1707
rect 860 1706 861 1707
rect 886 1707 892 1708
rect 886 1706 887 1707
rect 860 1704 887 1706
rect 860 1703 861 1704
rect 423 1702 429 1703
rect 454 1702 460 1703
rect 454 1698 455 1702
rect 459 1698 460 1702
rect 454 1697 460 1698
rect 502 1702 508 1703
rect 514 1702 525 1703
rect 550 1702 556 1703
rect 567 1702 573 1703
rect 606 1702 612 1703
rect 623 1702 629 1703
rect 662 1702 668 1703
rect 679 1702 685 1703
rect 726 1702 732 1703
rect 743 1702 749 1703
rect 782 1702 788 1703
rect 799 1702 805 1703
rect 838 1702 844 1703
rect 855 1702 861 1703
rect 886 1703 887 1704
rect 891 1703 892 1707
rect 911 1707 917 1708
rect 911 1706 912 1707
rect 904 1704 912 1706
rect 886 1702 892 1703
rect 894 1702 900 1703
rect 502 1698 503 1702
rect 507 1698 508 1702
rect 502 1697 508 1698
rect 550 1698 551 1702
rect 555 1698 556 1702
rect 550 1697 556 1698
rect 606 1698 607 1702
rect 611 1698 612 1702
rect 606 1697 612 1698
rect 662 1698 663 1702
rect 667 1698 668 1702
rect 662 1697 668 1698
rect 726 1698 727 1702
rect 731 1698 732 1702
rect 726 1697 732 1698
rect 782 1698 783 1702
rect 787 1698 788 1702
rect 782 1697 788 1698
rect 838 1698 839 1702
rect 843 1698 844 1702
rect 838 1697 844 1698
rect 894 1698 895 1702
rect 899 1698 900 1702
rect 894 1697 900 1698
rect 416 1692 427 1694
rect 904 1692 906 1704
rect 911 1703 912 1704
rect 916 1703 917 1707
rect 919 1707 920 1711
rect 924 1710 925 1711
rect 975 1711 981 1712
rect 924 1708 962 1710
rect 924 1707 925 1708
rect 919 1706 925 1707
rect 960 1706 962 1708
rect 967 1707 973 1708
rect 967 1706 968 1707
rect 960 1704 968 1706
rect 967 1703 968 1704
rect 972 1703 973 1707
rect 975 1707 976 1711
rect 980 1710 981 1711
rect 1031 1711 1037 1712
rect 980 1708 1018 1710
rect 980 1707 981 1708
rect 975 1706 981 1707
rect 1016 1706 1018 1708
rect 1023 1707 1029 1708
rect 1023 1706 1024 1707
rect 1016 1704 1024 1706
rect 1023 1703 1024 1704
rect 1028 1703 1029 1707
rect 1031 1707 1032 1711
rect 1036 1710 1037 1711
rect 1106 1711 1112 1712
rect 1036 1708 1074 1710
rect 1036 1707 1037 1708
rect 1031 1706 1037 1707
rect 1072 1706 1074 1708
rect 1079 1707 1085 1708
rect 1079 1706 1080 1707
rect 1072 1704 1080 1706
rect 1079 1703 1080 1704
rect 1084 1703 1085 1707
rect 1106 1707 1107 1711
rect 1111 1710 1112 1711
rect 1138 1711 1139 1715
rect 1143 1714 1144 1715
rect 1143 1712 1194 1714
rect 1143 1711 1144 1712
rect 1138 1710 1144 1711
rect 1192 1710 1194 1712
rect 1270 1711 1276 1712
rect 1111 1708 1130 1710
rect 1191 1709 1197 1710
rect 1111 1707 1112 1708
rect 1106 1706 1112 1707
rect 1128 1706 1130 1708
rect 1135 1707 1141 1708
rect 1135 1706 1136 1707
rect 1128 1704 1136 1706
rect 1135 1703 1136 1704
rect 1140 1703 1141 1707
rect 1191 1705 1192 1709
rect 1196 1705 1197 1709
rect 1191 1704 1197 1705
rect 1247 1707 1253 1708
rect 1247 1703 1248 1707
rect 1252 1706 1253 1707
rect 1262 1707 1268 1708
rect 1262 1706 1263 1707
rect 1252 1704 1263 1706
rect 1252 1703 1253 1704
rect 911 1702 917 1703
rect 950 1702 956 1703
rect 967 1702 973 1703
rect 1006 1702 1012 1703
rect 1023 1702 1029 1703
rect 1062 1702 1068 1703
rect 1079 1702 1085 1703
rect 1118 1702 1124 1703
rect 1135 1702 1141 1703
rect 1174 1702 1180 1703
rect 950 1698 951 1702
rect 955 1698 956 1702
rect 950 1697 956 1698
rect 1006 1698 1007 1702
rect 1011 1698 1012 1702
rect 1006 1697 1012 1698
rect 1062 1698 1063 1702
rect 1067 1698 1068 1702
rect 1062 1697 1068 1698
rect 1118 1698 1119 1702
rect 1123 1698 1124 1702
rect 1118 1697 1124 1698
rect 1174 1698 1175 1702
rect 1179 1698 1180 1702
rect 1174 1697 1180 1698
rect 1230 1702 1236 1703
rect 1247 1702 1253 1703
rect 1262 1703 1263 1704
rect 1267 1703 1268 1707
rect 1270 1707 1271 1711
rect 1275 1710 1276 1711
rect 1311 1711 1317 1712
rect 1275 1708 1298 1710
rect 1275 1707 1276 1708
rect 1270 1706 1276 1707
rect 1296 1706 1298 1708
rect 1303 1707 1309 1708
rect 1303 1706 1304 1707
rect 1296 1704 1304 1706
rect 1303 1703 1304 1704
rect 1308 1703 1309 1707
rect 1311 1707 1312 1711
rect 1316 1710 1317 1711
rect 1359 1711 1365 1712
rect 1316 1708 1355 1710
rect 1316 1707 1317 1708
rect 1311 1706 1317 1707
rect 1351 1707 1357 1708
rect 1351 1703 1352 1707
rect 1356 1703 1357 1707
rect 1359 1707 1360 1711
rect 1364 1710 1365 1711
rect 1399 1711 1405 1712
rect 1364 1708 1386 1710
rect 1364 1707 1365 1708
rect 1359 1706 1365 1707
rect 1384 1706 1386 1708
rect 1391 1707 1397 1708
rect 1391 1706 1392 1707
rect 1384 1704 1392 1706
rect 1391 1703 1392 1704
rect 1396 1703 1397 1707
rect 1399 1707 1400 1711
rect 1404 1710 1405 1711
rect 1458 1711 1464 1712
rect 1404 1708 1434 1710
rect 1404 1707 1405 1708
rect 1399 1706 1405 1707
rect 1432 1706 1434 1708
rect 1439 1707 1445 1708
rect 1439 1706 1440 1707
rect 1432 1704 1440 1706
rect 1439 1703 1440 1704
rect 1444 1703 1445 1707
rect 1458 1707 1459 1711
rect 1463 1710 1464 1711
rect 1495 1711 1501 1712
rect 1463 1708 1482 1710
rect 1463 1707 1464 1708
rect 1458 1706 1464 1707
rect 1480 1706 1482 1708
rect 1487 1707 1493 1708
rect 1487 1706 1488 1707
rect 1480 1704 1488 1706
rect 1487 1703 1488 1704
rect 1492 1703 1493 1707
rect 1495 1707 1496 1711
rect 1500 1710 1501 1711
rect 1500 1708 1530 1710
rect 1500 1707 1501 1708
rect 1495 1706 1501 1707
rect 1528 1706 1530 1708
rect 1535 1707 1541 1708
rect 1535 1706 1536 1707
rect 1528 1704 1536 1706
rect 1535 1703 1536 1704
rect 1540 1703 1541 1707
rect 1262 1702 1268 1703
rect 1286 1702 1292 1703
rect 1303 1702 1309 1703
rect 1334 1702 1340 1703
rect 1351 1702 1357 1703
rect 1374 1702 1380 1703
rect 1391 1702 1397 1703
rect 1422 1702 1428 1703
rect 1439 1702 1445 1703
rect 1470 1702 1476 1703
rect 1487 1702 1493 1703
rect 1518 1702 1524 1703
rect 1535 1702 1541 1703
rect 1662 1704 1668 1705
rect 1230 1698 1231 1702
rect 1235 1698 1236 1702
rect 1230 1697 1236 1698
rect 1286 1698 1287 1702
rect 1291 1698 1292 1702
rect 1286 1697 1292 1698
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1374 1698 1375 1702
rect 1379 1698 1380 1702
rect 1374 1697 1380 1698
rect 1422 1698 1423 1702
rect 1427 1698 1428 1702
rect 1422 1697 1428 1698
rect 1470 1698 1471 1702
rect 1475 1698 1476 1702
rect 1470 1697 1476 1698
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1662 1700 1663 1704
rect 1667 1700 1668 1704
rect 1662 1699 1668 1700
rect 1518 1697 1524 1698
rect 276 1688 282 1690
rect 303 1691 309 1692
rect 276 1687 277 1688
rect 271 1686 277 1687
rect 303 1687 304 1691
rect 308 1690 309 1691
rect 316 1690 330 1692
rect 335 1691 341 1692
rect 308 1688 318 1690
rect 308 1687 309 1688
rect 303 1686 309 1687
rect 335 1687 336 1691
rect 340 1690 341 1691
rect 350 1691 356 1692
rect 350 1690 351 1691
rect 340 1688 351 1690
rect 340 1687 341 1688
rect 335 1686 341 1687
rect 350 1687 351 1688
rect 355 1687 356 1691
rect 350 1686 356 1687
rect 374 1691 381 1692
rect 374 1687 375 1691
rect 380 1687 381 1691
rect 374 1686 381 1687
rect 423 1691 429 1692
rect 423 1687 424 1691
rect 428 1687 429 1691
rect 423 1686 429 1687
rect 470 1691 477 1692
rect 470 1687 471 1691
rect 476 1687 477 1691
rect 470 1686 477 1687
rect 519 1691 525 1692
rect 519 1687 520 1691
rect 524 1690 525 1691
rect 538 1691 544 1692
rect 538 1690 539 1691
rect 524 1688 539 1690
rect 524 1687 525 1688
rect 519 1686 525 1687
rect 538 1687 539 1688
rect 543 1687 544 1691
rect 538 1686 544 1687
rect 567 1691 573 1692
rect 567 1687 568 1691
rect 572 1690 573 1691
rect 575 1691 581 1692
rect 575 1690 576 1691
rect 572 1688 576 1690
rect 572 1687 573 1688
rect 567 1686 573 1687
rect 575 1687 576 1688
rect 580 1687 581 1691
rect 575 1686 581 1687
rect 623 1691 629 1692
rect 623 1687 624 1691
rect 628 1690 629 1691
rect 631 1691 637 1692
rect 631 1690 632 1691
rect 628 1688 632 1690
rect 628 1687 629 1688
rect 623 1686 629 1687
rect 631 1687 632 1688
rect 636 1687 637 1691
rect 631 1686 637 1687
rect 679 1691 685 1692
rect 679 1687 680 1691
rect 684 1690 685 1691
rect 687 1691 693 1692
rect 687 1690 688 1691
rect 684 1688 688 1690
rect 684 1687 685 1688
rect 679 1686 685 1687
rect 687 1687 688 1688
rect 692 1687 693 1691
rect 687 1686 693 1687
rect 743 1691 749 1692
rect 743 1687 744 1691
rect 748 1690 749 1691
rect 751 1691 757 1692
rect 751 1690 752 1691
rect 748 1688 752 1690
rect 748 1687 749 1688
rect 743 1686 749 1687
rect 751 1687 752 1688
rect 756 1687 757 1691
rect 751 1686 757 1687
rect 799 1691 808 1692
rect 799 1687 800 1691
rect 807 1687 808 1691
rect 799 1686 808 1687
rect 855 1691 861 1692
rect 855 1687 856 1691
rect 860 1690 861 1691
rect 892 1690 906 1692
rect 911 1691 917 1692
rect 860 1688 894 1690
rect 860 1687 861 1688
rect 855 1686 861 1687
rect 911 1687 912 1691
rect 916 1690 917 1691
rect 919 1691 925 1692
rect 919 1690 920 1691
rect 916 1688 920 1690
rect 916 1687 917 1688
rect 911 1686 917 1687
rect 919 1687 920 1688
rect 924 1687 925 1691
rect 919 1686 925 1687
rect 967 1691 973 1692
rect 967 1687 968 1691
rect 972 1690 973 1691
rect 975 1691 981 1692
rect 975 1690 976 1691
rect 972 1688 976 1690
rect 972 1687 973 1688
rect 967 1686 973 1687
rect 975 1687 976 1688
rect 980 1687 981 1691
rect 975 1686 981 1687
rect 1023 1691 1029 1692
rect 1023 1687 1024 1691
rect 1028 1690 1029 1691
rect 1031 1691 1037 1692
rect 1031 1690 1032 1691
rect 1028 1688 1032 1690
rect 1028 1687 1029 1688
rect 1023 1686 1029 1687
rect 1031 1687 1032 1688
rect 1036 1687 1037 1691
rect 1031 1686 1037 1687
rect 1079 1691 1085 1692
rect 1079 1687 1080 1691
rect 1084 1690 1085 1691
rect 1106 1691 1112 1692
rect 1106 1690 1107 1691
rect 1084 1688 1107 1690
rect 1084 1687 1085 1688
rect 1079 1686 1085 1687
rect 1106 1687 1107 1688
rect 1111 1687 1112 1691
rect 1106 1686 1112 1687
rect 1135 1691 1144 1692
rect 1135 1687 1136 1691
rect 1143 1687 1144 1691
rect 1135 1686 1144 1687
rect 1190 1691 1197 1692
rect 1190 1687 1191 1691
rect 1196 1687 1197 1691
rect 1190 1686 1197 1687
rect 1247 1691 1253 1692
rect 1247 1687 1248 1691
rect 1252 1690 1253 1691
rect 1270 1691 1276 1692
rect 1270 1690 1271 1691
rect 1252 1688 1271 1690
rect 1252 1687 1253 1688
rect 1247 1686 1253 1687
rect 1270 1687 1271 1688
rect 1275 1687 1276 1691
rect 1270 1686 1276 1687
rect 1303 1691 1309 1692
rect 1303 1687 1304 1691
rect 1308 1690 1309 1691
rect 1311 1691 1317 1692
rect 1311 1690 1312 1691
rect 1308 1688 1312 1690
rect 1308 1687 1309 1688
rect 1303 1686 1309 1687
rect 1311 1687 1312 1688
rect 1316 1687 1317 1691
rect 1311 1686 1317 1687
rect 1351 1691 1357 1692
rect 1351 1687 1352 1691
rect 1356 1690 1357 1691
rect 1359 1691 1365 1692
rect 1359 1690 1360 1691
rect 1356 1688 1360 1690
rect 1356 1687 1357 1688
rect 1351 1686 1357 1687
rect 1359 1687 1360 1688
rect 1364 1687 1365 1691
rect 1359 1686 1365 1687
rect 1391 1691 1397 1692
rect 1391 1687 1392 1691
rect 1396 1690 1397 1691
rect 1399 1691 1405 1692
rect 1399 1690 1400 1691
rect 1396 1688 1400 1690
rect 1396 1687 1397 1688
rect 1391 1686 1397 1687
rect 1399 1687 1400 1688
rect 1404 1687 1405 1691
rect 1399 1686 1405 1687
rect 1439 1691 1445 1692
rect 1439 1687 1440 1691
rect 1444 1690 1445 1691
rect 1458 1691 1464 1692
rect 1458 1690 1459 1691
rect 1444 1688 1459 1690
rect 1444 1687 1445 1688
rect 1439 1686 1445 1687
rect 1458 1687 1459 1688
rect 1463 1687 1464 1691
rect 1458 1686 1464 1687
rect 1487 1691 1493 1692
rect 1487 1687 1488 1691
rect 1492 1690 1493 1691
rect 1495 1691 1501 1692
rect 1495 1690 1496 1691
rect 1492 1688 1496 1690
rect 1492 1687 1493 1688
rect 1487 1686 1493 1687
rect 1495 1687 1496 1688
rect 1500 1687 1501 1691
rect 1535 1691 1541 1692
rect 1535 1690 1536 1691
rect 1495 1686 1501 1687
rect 1528 1688 1536 1690
rect 110 1682 116 1683
rect 254 1685 260 1686
rect 254 1681 255 1685
rect 259 1681 260 1685
rect 254 1680 260 1681
rect 286 1685 292 1686
rect 286 1681 287 1685
rect 291 1681 292 1685
rect 286 1680 292 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 358 1685 364 1686
rect 358 1681 359 1685
rect 363 1681 364 1685
rect 358 1680 364 1681
rect 406 1685 412 1686
rect 406 1681 407 1685
rect 411 1681 412 1685
rect 406 1680 412 1681
rect 454 1685 460 1686
rect 454 1681 455 1685
rect 459 1681 460 1685
rect 454 1680 460 1681
rect 502 1685 508 1686
rect 502 1681 503 1685
rect 507 1681 508 1685
rect 502 1680 508 1681
rect 550 1685 556 1686
rect 550 1681 551 1685
rect 555 1681 556 1685
rect 550 1680 556 1681
rect 606 1685 612 1686
rect 606 1681 607 1685
rect 611 1681 612 1685
rect 606 1680 612 1681
rect 662 1685 668 1686
rect 662 1681 663 1685
rect 667 1681 668 1685
rect 662 1680 668 1681
rect 726 1685 732 1686
rect 726 1681 727 1685
rect 731 1681 732 1685
rect 726 1680 732 1681
rect 782 1685 788 1686
rect 782 1681 783 1685
rect 787 1681 788 1685
rect 782 1680 788 1681
rect 838 1685 844 1686
rect 838 1681 839 1685
rect 843 1681 844 1685
rect 838 1680 844 1681
rect 894 1685 900 1686
rect 894 1681 895 1685
rect 899 1681 900 1685
rect 894 1680 900 1681
rect 950 1685 956 1686
rect 950 1681 951 1685
rect 955 1681 956 1685
rect 950 1680 956 1681
rect 1006 1685 1012 1686
rect 1006 1681 1007 1685
rect 1011 1681 1012 1685
rect 1006 1680 1012 1681
rect 1062 1685 1068 1686
rect 1062 1681 1063 1685
rect 1067 1681 1068 1685
rect 1062 1680 1068 1681
rect 1118 1685 1124 1686
rect 1118 1681 1119 1685
rect 1123 1681 1124 1685
rect 1118 1680 1124 1681
rect 1174 1685 1180 1686
rect 1174 1681 1175 1685
rect 1179 1681 1180 1685
rect 1174 1680 1180 1681
rect 1230 1685 1236 1686
rect 1230 1681 1231 1685
rect 1235 1681 1236 1685
rect 1230 1680 1236 1681
rect 1286 1685 1292 1686
rect 1286 1681 1287 1685
rect 1291 1681 1292 1685
rect 1286 1680 1292 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1374 1685 1380 1686
rect 1374 1681 1375 1685
rect 1379 1681 1380 1685
rect 1374 1680 1380 1681
rect 1422 1685 1428 1686
rect 1422 1681 1423 1685
rect 1427 1681 1428 1685
rect 1422 1680 1428 1681
rect 1470 1685 1476 1686
rect 1470 1681 1471 1685
rect 1475 1681 1476 1685
rect 1470 1680 1476 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1518 1680 1524 1681
rect 1410 1679 1416 1680
rect 1410 1675 1411 1679
rect 1415 1678 1416 1679
rect 1528 1678 1530 1688
rect 1535 1687 1536 1688
rect 1540 1687 1541 1691
rect 1535 1686 1541 1687
rect 1662 1687 1668 1688
rect 1662 1683 1663 1687
rect 1667 1683 1668 1687
rect 1662 1682 1668 1683
rect 1415 1676 1530 1678
rect 1415 1675 1416 1676
rect 1410 1674 1416 1675
rect 134 1671 140 1672
rect 110 1669 116 1670
rect 110 1665 111 1669
rect 115 1665 116 1669
rect 134 1667 135 1671
rect 139 1667 140 1671
rect 134 1666 140 1667
rect 166 1671 172 1672
rect 166 1667 167 1671
rect 171 1667 172 1671
rect 166 1666 172 1667
rect 214 1671 220 1672
rect 214 1667 215 1671
rect 219 1667 220 1671
rect 214 1666 220 1667
rect 278 1671 284 1672
rect 278 1667 279 1671
rect 283 1667 284 1671
rect 278 1666 284 1667
rect 342 1671 348 1672
rect 342 1667 343 1671
rect 347 1667 348 1671
rect 342 1666 348 1667
rect 414 1671 420 1672
rect 414 1667 415 1671
rect 419 1667 420 1671
rect 414 1666 420 1667
rect 486 1671 492 1672
rect 486 1667 487 1671
rect 491 1667 492 1671
rect 558 1671 564 1672
rect 486 1666 492 1667
rect 514 1667 520 1668
rect 514 1666 515 1667
rect 110 1664 116 1665
rect 503 1665 515 1666
rect 150 1663 157 1664
rect 150 1659 151 1663
rect 156 1659 157 1663
rect 183 1663 189 1664
rect 183 1662 184 1663
rect 150 1658 157 1659
rect 176 1660 184 1662
rect 134 1654 140 1655
rect 110 1652 116 1653
rect 110 1648 111 1652
rect 115 1648 116 1652
rect 134 1650 135 1654
rect 139 1650 140 1654
rect 134 1649 140 1650
rect 166 1654 172 1655
rect 166 1650 167 1654
rect 171 1650 172 1654
rect 166 1649 172 1650
rect 110 1647 116 1648
rect 151 1647 157 1648
rect 151 1643 152 1647
rect 156 1646 157 1647
rect 176 1646 178 1660
rect 183 1659 184 1660
rect 188 1659 189 1663
rect 231 1663 237 1664
rect 231 1662 232 1663
rect 183 1658 189 1659
rect 208 1660 232 1662
rect 156 1644 178 1646
rect 183 1647 189 1648
rect 156 1643 157 1644
rect 151 1642 157 1643
rect 183 1643 184 1647
rect 188 1646 189 1647
rect 208 1646 210 1660
rect 231 1659 232 1660
rect 236 1659 237 1663
rect 295 1663 301 1664
rect 295 1662 296 1663
rect 231 1658 237 1659
rect 268 1660 296 1662
rect 214 1654 220 1655
rect 214 1650 215 1654
rect 219 1650 220 1654
rect 214 1649 220 1650
rect 188 1644 210 1646
rect 231 1647 237 1648
rect 188 1643 189 1644
rect 183 1642 189 1643
rect 231 1643 232 1647
rect 236 1646 237 1647
rect 268 1646 270 1660
rect 295 1659 296 1660
rect 300 1659 301 1663
rect 359 1663 365 1664
rect 359 1662 360 1663
rect 295 1658 301 1659
rect 319 1660 360 1662
rect 278 1654 284 1655
rect 278 1650 279 1654
rect 283 1650 284 1654
rect 278 1649 284 1650
rect 236 1644 270 1646
rect 295 1647 301 1648
rect 236 1643 237 1644
rect 231 1642 237 1643
rect 295 1643 296 1647
rect 300 1646 301 1647
rect 319 1646 321 1660
rect 359 1659 360 1660
rect 364 1659 365 1663
rect 359 1658 365 1659
rect 431 1663 437 1664
rect 431 1659 432 1663
rect 436 1662 437 1663
rect 436 1660 483 1662
rect 503 1661 504 1665
rect 508 1664 515 1665
rect 508 1661 509 1664
rect 514 1663 515 1664
rect 519 1663 520 1667
rect 558 1667 559 1671
rect 563 1667 564 1671
rect 558 1666 564 1667
rect 630 1671 636 1672
rect 630 1667 631 1671
rect 635 1667 636 1671
rect 630 1666 636 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 710 1666 716 1667
rect 790 1671 796 1672
rect 790 1667 791 1671
rect 795 1667 796 1671
rect 790 1666 796 1667
rect 870 1671 876 1672
rect 870 1667 871 1671
rect 875 1667 876 1671
rect 870 1666 876 1667
rect 950 1671 956 1672
rect 950 1667 951 1671
rect 955 1667 956 1671
rect 950 1666 956 1667
rect 1030 1671 1036 1672
rect 1030 1667 1031 1671
rect 1035 1667 1036 1671
rect 1030 1666 1036 1667
rect 1102 1671 1108 1672
rect 1102 1667 1103 1671
rect 1107 1667 1108 1671
rect 1102 1666 1108 1667
rect 1174 1671 1180 1672
rect 1174 1667 1175 1671
rect 1179 1667 1180 1671
rect 1174 1666 1180 1667
rect 1246 1671 1252 1672
rect 1246 1667 1247 1671
rect 1251 1667 1252 1671
rect 1246 1666 1252 1667
rect 1318 1671 1324 1672
rect 1318 1667 1319 1671
rect 1323 1667 1324 1671
rect 1318 1666 1324 1667
rect 1390 1671 1396 1672
rect 1390 1667 1391 1671
rect 1395 1667 1396 1671
rect 1390 1666 1396 1667
rect 1454 1671 1460 1672
rect 1454 1667 1455 1671
rect 1459 1667 1460 1671
rect 1454 1666 1460 1667
rect 1518 1671 1524 1672
rect 1518 1667 1519 1671
rect 1523 1667 1524 1671
rect 1518 1666 1524 1667
rect 1582 1671 1588 1672
rect 1582 1667 1583 1671
rect 1587 1667 1588 1671
rect 1582 1666 1588 1667
rect 1622 1671 1628 1672
rect 1622 1667 1623 1671
rect 1627 1667 1628 1671
rect 1622 1666 1628 1667
rect 1662 1669 1668 1670
rect 1662 1665 1663 1669
rect 1667 1665 1668 1669
rect 1662 1664 1668 1665
rect 514 1662 520 1663
rect 522 1663 528 1664
rect 503 1660 509 1661
rect 436 1659 437 1660
rect 431 1658 437 1659
rect 342 1654 348 1655
rect 342 1650 343 1654
rect 347 1650 348 1654
rect 342 1649 348 1650
rect 414 1654 420 1655
rect 414 1650 415 1654
rect 419 1650 420 1654
rect 414 1649 420 1650
rect 300 1644 321 1646
rect 350 1647 356 1648
rect 300 1643 301 1644
rect 295 1642 301 1643
rect 350 1643 351 1647
rect 355 1646 356 1647
rect 359 1647 365 1648
rect 359 1646 360 1647
rect 355 1644 360 1646
rect 355 1643 356 1644
rect 350 1642 356 1643
rect 359 1643 360 1644
rect 364 1643 365 1647
rect 359 1642 365 1643
rect 431 1647 437 1648
rect 431 1643 432 1647
rect 436 1643 437 1647
rect 481 1646 483 1660
rect 522 1659 523 1663
rect 527 1662 528 1663
rect 575 1663 581 1664
rect 575 1662 576 1663
rect 527 1660 576 1662
rect 527 1659 528 1660
rect 522 1658 528 1659
rect 575 1659 576 1660
rect 580 1659 581 1663
rect 575 1658 581 1659
rect 647 1663 653 1664
rect 647 1659 648 1663
rect 652 1662 653 1663
rect 678 1663 684 1664
rect 678 1662 679 1663
rect 652 1660 679 1662
rect 652 1659 653 1660
rect 647 1658 653 1659
rect 678 1659 679 1660
rect 683 1659 684 1663
rect 727 1663 733 1664
rect 727 1662 728 1663
rect 678 1658 684 1659
rect 689 1660 728 1662
rect 486 1654 492 1655
rect 486 1650 487 1654
rect 491 1650 492 1654
rect 486 1649 492 1650
rect 558 1654 564 1655
rect 558 1650 559 1654
rect 563 1650 564 1654
rect 558 1649 564 1650
rect 630 1654 636 1655
rect 630 1650 631 1654
rect 635 1650 636 1654
rect 630 1649 636 1650
rect 503 1647 509 1648
rect 503 1646 504 1647
rect 481 1644 504 1646
rect 431 1642 437 1643
rect 503 1643 504 1644
rect 508 1643 509 1647
rect 503 1642 509 1643
rect 575 1647 581 1648
rect 575 1643 576 1647
rect 580 1646 581 1647
rect 614 1647 620 1648
rect 614 1646 615 1647
rect 580 1644 615 1646
rect 580 1643 581 1644
rect 575 1642 581 1643
rect 614 1643 615 1644
rect 619 1643 620 1647
rect 614 1642 620 1643
rect 647 1647 653 1648
rect 647 1643 648 1647
rect 652 1646 653 1647
rect 689 1646 691 1660
rect 727 1659 728 1660
rect 732 1659 733 1663
rect 807 1663 813 1664
rect 807 1662 808 1663
rect 727 1658 733 1659
rect 772 1660 808 1662
rect 710 1654 716 1655
rect 710 1650 711 1654
rect 715 1650 716 1654
rect 710 1649 716 1650
rect 652 1644 691 1646
rect 727 1647 733 1648
rect 652 1643 653 1644
rect 647 1642 653 1643
rect 727 1643 728 1647
rect 732 1646 733 1647
rect 772 1646 774 1660
rect 807 1659 808 1660
rect 812 1659 813 1663
rect 807 1658 813 1659
rect 886 1663 893 1664
rect 886 1659 887 1663
rect 892 1659 893 1663
rect 967 1663 973 1664
rect 967 1662 968 1663
rect 886 1658 893 1659
rect 929 1660 968 1662
rect 790 1654 796 1655
rect 790 1650 791 1654
rect 795 1650 796 1654
rect 790 1649 796 1650
rect 870 1654 876 1655
rect 870 1650 871 1654
rect 875 1650 876 1654
rect 870 1649 876 1650
rect 732 1644 774 1646
rect 802 1647 813 1648
rect 732 1643 733 1644
rect 727 1642 733 1643
rect 802 1643 803 1647
rect 807 1643 808 1647
rect 812 1643 813 1647
rect 802 1642 813 1643
rect 887 1647 893 1648
rect 887 1643 888 1647
rect 892 1646 893 1647
rect 929 1646 931 1660
rect 967 1659 968 1660
rect 972 1659 973 1663
rect 967 1658 973 1659
rect 1047 1663 1053 1664
rect 1047 1659 1048 1663
rect 1052 1662 1053 1663
rect 1119 1663 1125 1664
rect 1052 1660 1114 1662
rect 1052 1659 1053 1660
rect 1047 1658 1053 1659
rect 950 1654 956 1655
rect 950 1650 951 1654
rect 955 1650 956 1654
rect 950 1649 956 1650
rect 1030 1654 1036 1655
rect 1030 1650 1031 1654
rect 1035 1650 1036 1654
rect 1030 1649 1036 1650
rect 1102 1654 1108 1655
rect 1102 1650 1103 1654
rect 1107 1650 1108 1654
rect 1102 1649 1108 1650
rect 892 1644 931 1646
rect 962 1647 973 1648
rect 892 1643 893 1644
rect 887 1642 893 1643
rect 962 1643 963 1647
rect 967 1643 968 1647
rect 972 1643 973 1647
rect 962 1642 973 1643
rect 1047 1647 1053 1648
rect 1047 1643 1048 1647
rect 1052 1643 1053 1647
rect 1112 1646 1114 1660
rect 1119 1659 1120 1663
rect 1124 1662 1125 1663
rect 1146 1663 1152 1664
rect 1124 1660 1142 1662
rect 1124 1659 1125 1660
rect 1119 1658 1125 1659
rect 1140 1654 1142 1660
rect 1146 1659 1147 1663
rect 1151 1662 1152 1663
rect 1191 1663 1197 1664
rect 1191 1662 1192 1663
rect 1151 1660 1192 1662
rect 1151 1659 1152 1660
rect 1146 1658 1152 1659
rect 1191 1659 1192 1660
rect 1196 1659 1197 1663
rect 1191 1658 1197 1659
rect 1262 1663 1269 1664
rect 1262 1659 1263 1663
rect 1268 1659 1269 1663
rect 1335 1663 1341 1664
rect 1335 1662 1336 1663
rect 1262 1658 1269 1659
rect 1300 1660 1336 1662
rect 1166 1655 1172 1656
rect 1166 1654 1167 1655
rect 1140 1652 1167 1654
rect 1166 1651 1167 1652
rect 1171 1651 1172 1655
rect 1166 1650 1172 1651
rect 1174 1654 1180 1655
rect 1174 1650 1175 1654
rect 1179 1650 1180 1654
rect 1174 1649 1180 1650
rect 1246 1654 1252 1655
rect 1246 1650 1247 1654
rect 1251 1650 1252 1654
rect 1246 1649 1252 1650
rect 1119 1647 1125 1648
rect 1119 1646 1120 1647
rect 1112 1644 1120 1646
rect 1047 1642 1053 1643
rect 1119 1643 1120 1644
rect 1124 1643 1125 1647
rect 1119 1642 1125 1643
rect 1190 1647 1197 1648
rect 1190 1643 1191 1647
rect 1196 1643 1197 1647
rect 1190 1642 1197 1643
rect 1263 1647 1269 1648
rect 1263 1643 1264 1647
rect 1268 1646 1269 1647
rect 1300 1646 1302 1660
rect 1335 1659 1336 1660
rect 1340 1659 1341 1663
rect 1335 1658 1341 1659
rect 1407 1663 1413 1664
rect 1407 1659 1408 1663
rect 1412 1662 1413 1663
rect 1471 1663 1477 1664
rect 1412 1660 1442 1662
rect 1412 1659 1413 1660
rect 1407 1658 1413 1659
rect 1318 1654 1324 1655
rect 1318 1650 1319 1654
rect 1323 1650 1324 1654
rect 1318 1649 1324 1650
rect 1390 1654 1396 1655
rect 1390 1650 1391 1654
rect 1395 1650 1396 1654
rect 1390 1649 1396 1650
rect 1268 1644 1302 1646
rect 1334 1647 1341 1648
rect 1268 1643 1269 1644
rect 1263 1642 1269 1643
rect 1334 1643 1335 1647
rect 1340 1643 1341 1647
rect 1334 1642 1341 1643
rect 1407 1647 1416 1648
rect 1407 1643 1408 1647
rect 1415 1643 1416 1647
rect 1440 1646 1442 1660
rect 1471 1659 1472 1663
rect 1476 1662 1477 1663
rect 1535 1663 1541 1664
rect 1476 1660 1530 1662
rect 1476 1659 1477 1660
rect 1471 1658 1477 1659
rect 1454 1654 1460 1655
rect 1454 1650 1455 1654
rect 1459 1650 1460 1654
rect 1454 1649 1460 1650
rect 1518 1654 1524 1655
rect 1518 1650 1519 1654
rect 1523 1650 1524 1654
rect 1518 1649 1524 1650
rect 1471 1647 1477 1648
rect 1471 1646 1472 1647
rect 1440 1644 1472 1646
rect 1407 1642 1416 1643
rect 1471 1643 1472 1644
rect 1476 1643 1477 1647
rect 1528 1646 1530 1660
rect 1535 1659 1536 1663
rect 1540 1662 1541 1663
rect 1574 1663 1580 1664
rect 1574 1662 1575 1663
rect 1540 1660 1575 1662
rect 1540 1659 1541 1660
rect 1535 1658 1541 1659
rect 1574 1659 1575 1660
rect 1579 1659 1580 1663
rect 1574 1658 1580 1659
rect 1599 1663 1605 1664
rect 1599 1659 1600 1663
rect 1604 1662 1605 1663
rect 1638 1663 1645 1664
rect 1604 1660 1618 1662
rect 1604 1659 1605 1660
rect 1599 1658 1605 1659
rect 1582 1654 1588 1655
rect 1582 1650 1583 1654
rect 1587 1650 1588 1654
rect 1582 1649 1588 1650
rect 1535 1647 1541 1648
rect 1535 1646 1536 1647
rect 1528 1644 1536 1646
rect 1471 1642 1477 1643
rect 1535 1643 1536 1644
rect 1540 1643 1541 1647
rect 1535 1642 1541 1643
rect 1546 1647 1552 1648
rect 1546 1643 1547 1647
rect 1551 1646 1552 1647
rect 1599 1647 1605 1648
rect 1599 1646 1600 1647
rect 1551 1644 1600 1646
rect 1551 1643 1552 1644
rect 1546 1642 1552 1643
rect 1599 1643 1600 1644
rect 1604 1643 1605 1647
rect 1616 1646 1618 1660
rect 1638 1659 1639 1663
rect 1644 1659 1645 1663
rect 1638 1658 1645 1659
rect 1622 1654 1628 1655
rect 1622 1650 1623 1654
rect 1627 1650 1628 1654
rect 1622 1649 1628 1650
rect 1662 1652 1668 1653
rect 1662 1648 1663 1652
rect 1667 1648 1668 1652
rect 1639 1647 1645 1648
rect 1662 1647 1668 1648
rect 1639 1646 1640 1647
rect 1616 1644 1640 1646
rect 1599 1642 1605 1643
rect 1639 1643 1640 1644
rect 1644 1643 1645 1647
rect 1639 1642 1645 1643
rect 433 1638 435 1642
rect 522 1639 528 1640
rect 522 1638 523 1639
rect 433 1636 523 1638
rect 522 1635 523 1636
rect 527 1635 528 1639
rect 1049 1638 1051 1642
rect 1146 1639 1152 1640
rect 1146 1638 1147 1639
rect 1049 1636 1147 1638
rect 522 1634 528 1635
rect 1146 1635 1147 1636
rect 1151 1635 1152 1639
rect 1146 1634 1152 1635
rect 207 1631 213 1632
rect 150 1627 157 1628
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 150 1623 151 1627
rect 156 1623 157 1627
rect 198 1627 205 1628
rect 198 1623 199 1627
rect 204 1623 205 1627
rect 207 1627 208 1631
rect 212 1630 213 1631
rect 271 1631 277 1632
rect 212 1628 258 1630
rect 212 1627 213 1628
rect 207 1626 213 1627
rect 256 1626 258 1628
rect 263 1627 269 1628
rect 263 1626 264 1627
rect 256 1624 264 1626
rect 263 1623 264 1624
rect 268 1623 269 1627
rect 271 1627 272 1631
rect 276 1630 277 1631
rect 327 1631 333 1632
rect 276 1628 321 1630
rect 276 1627 277 1628
rect 271 1626 277 1627
rect 319 1627 325 1628
rect 319 1623 320 1627
rect 324 1623 325 1627
rect 327 1627 328 1631
rect 332 1630 333 1631
rect 383 1631 389 1632
rect 332 1628 370 1630
rect 332 1627 333 1628
rect 327 1626 333 1627
rect 368 1626 370 1628
rect 375 1627 381 1628
rect 375 1626 376 1627
rect 368 1624 376 1626
rect 375 1623 376 1624
rect 380 1623 381 1627
rect 383 1627 384 1631
rect 388 1630 389 1631
rect 498 1631 504 1632
rect 388 1628 435 1630
rect 388 1627 389 1628
rect 383 1626 389 1627
rect 431 1627 437 1628
rect 431 1623 432 1627
rect 436 1623 437 1627
rect 487 1627 496 1628
rect 487 1623 488 1627
rect 495 1623 496 1627
rect 498 1627 499 1631
rect 503 1630 504 1631
rect 559 1631 565 1632
rect 503 1628 555 1630
rect 503 1627 504 1628
rect 498 1626 504 1627
rect 551 1627 557 1628
rect 551 1623 552 1627
rect 556 1623 557 1627
rect 559 1627 560 1631
rect 564 1630 565 1631
rect 687 1631 693 1632
rect 564 1628 619 1630
rect 564 1627 565 1628
rect 559 1626 565 1627
rect 615 1627 621 1628
rect 615 1623 616 1627
rect 620 1623 621 1627
rect 678 1627 685 1628
rect 678 1623 679 1627
rect 684 1623 685 1627
rect 687 1627 688 1631
rect 692 1630 693 1631
rect 823 1631 829 1632
rect 692 1628 747 1630
rect 692 1627 693 1628
rect 687 1626 693 1627
rect 743 1627 749 1628
rect 743 1623 744 1627
rect 748 1623 749 1627
rect 814 1627 821 1628
rect 814 1623 815 1627
rect 820 1623 821 1627
rect 823 1627 824 1631
rect 828 1630 829 1631
rect 895 1631 901 1632
rect 828 1628 882 1630
rect 828 1627 829 1628
rect 823 1626 829 1627
rect 880 1626 882 1628
rect 887 1627 893 1628
rect 887 1626 888 1627
rect 880 1624 888 1626
rect 887 1623 888 1624
rect 892 1623 893 1627
rect 895 1627 896 1631
rect 900 1630 901 1631
rect 1166 1631 1172 1632
rect 900 1628 954 1630
rect 1096 1628 1114 1630
rect 900 1627 901 1628
rect 895 1626 901 1627
rect 952 1626 954 1628
rect 959 1627 965 1628
rect 959 1626 960 1627
rect 952 1624 960 1626
rect 959 1623 960 1624
rect 964 1623 965 1627
rect 1039 1627 1045 1628
rect 1039 1623 1040 1627
rect 1044 1626 1045 1627
rect 1096 1626 1098 1628
rect 1044 1624 1098 1626
rect 1044 1623 1045 1624
rect 110 1619 116 1620
rect 134 1622 140 1623
rect 150 1622 157 1623
rect 182 1622 188 1623
rect 198 1622 205 1623
rect 246 1622 252 1623
rect 263 1622 269 1623
rect 302 1622 308 1623
rect 319 1622 325 1623
rect 358 1622 364 1623
rect 375 1622 381 1623
rect 414 1622 420 1623
rect 431 1622 437 1623
rect 470 1622 476 1623
rect 487 1622 496 1623
rect 534 1622 540 1623
rect 551 1622 557 1623
rect 598 1622 604 1623
rect 615 1622 621 1623
rect 662 1622 668 1623
rect 678 1622 685 1623
rect 726 1622 732 1623
rect 743 1622 749 1623
rect 798 1622 804 1623
rect 814 1622 821 1623
rect 870 1622 876 1623
rect 887 1622 893 1623
rect 942 1622 948 1623
rect 959 1622 965 1623
rect 1022 1622 1028 1623
rect 1039 1622 1045 1623
rect 1102 1622 1108 1623
rect 134 1618 135 1622
rect 139 1618 140 1622
rect 134 1617 140 1618
rect 182 1618 183 1622
rect 187 1618 188 1622
rect 182 1617 188 1618
rect 246 1618 247 1622
rect 251 1618 252 1622
rect 246 1617 252 1618
rect 302 1618 303 1622
rect 307 1618 308 1622
rect 302 1617 308 1618
rect 358 1618 359 1622
rect 363 1618 364 1622
rect 358 1617 364 1618
rect 414 1618 415 1622
rect 419 1618 420 1622
rect 414 1617 420 1618
rect 470 1618 471 1622
rect 475 1618 476 1622
rect 470 1617 476 1618
rect 534 1618 535 1622
rect 539 1618 540 1622
rect 534 1617 540 1618
rect 598 1618 599 1622
rect 603 1618 604 1622
rect 598 1617 604 1618
rect 662 1618 663 1622
rect 667 1618 668 1622
rect 662 1617 668 1618
rect 726 1618 727 1622
rect 731 1618 732 1622
rect 726 1617 732 1618
rect 798 1618 799 1622
rect 803 1618 804 1622
rect 798 1617 804 1618
rect 870 1618 871 1622
rect 875 1618 876 1622
rect 870 1617 876 1618
rect 942 1618 943 1622
rect 947 1618 948 1622
rect 942 1617 948 1618
rect 1022 1618 1023 1622
rect 1027 1618 1028 1622
rect 1022 1617 1028 1618
rect 1102 1618 1103 1622
rect 1107 1618 1108 1622
rect 1102 1617 1108 1618
rect 150 1611 157 1612
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 150 1607 151 1611
rect 156 1607 157 1611
rect 150 1606 157 1607
rect 199 1611 205 1612
rect 199 1607 200 1611
rect 204 1610 205 1611
rect 207 1611 213 1612
rect 207 1610 208 1611
rect 204 1608 208 1610
rect 204 1607 205 1608
rect 199 1606 205 1607
rect 207 1607 208 1608
rect 212 1607 213 1611
rect 207 1606 213 1607
rect 263 1611 269 1612
rect 263 1607 264 1611
rect 268 1610 269 1611
rect 271 1611 277 1612
rect 271 1610 272 1611
rect 268 1608 272 1610
rect 268 1607 269 1608
rect 263 1606 269 1607
rect 271 1607 272 1608
rect 276 1607 277 1611
rect 271 1606 277 1607
rect 319 1611 325 1612
rect 319 1607 320 1611
rect 324 1610 325 1611
rect 327 1611 333 1612
rect 327 1610 328 1611
rect 324 1608 328 1610
rect 324 1607 325 1608
rect 319 1606 325 1607
rect 327 1607 328 1608
rect 332 1607 333 1611
rect 327 1606 333 1607
rect 375 1611 381 1612
rect 375 1607 376 1611
rect 380 1610 381 1611
rect 383 1611 389 1612
rect 383 1610 384 1611
rect 380 1608 384 1610
rect 380 1607 381 1608
rect 375 1606 381 1607
rect 383 1607 384 1608
rect 388 1607 389 1611
rect 383 1606 389 1607
rect 431 1611 437 1612
rect 431 1607 432 1611
rect 436 1610 437 1611
rect 446 1611 452 1612
rect 446 1610 447 1611
rect 436 1608 447 1610
rect 436 1607 437 1608
rect 431 1606 437 1607
rect 446 1607 447 1608
rect 451 1607 452 1611
rect 446 1606 452 1607
rect 487 1611 493 1612
rect 487 1607 488 1611
rect 492 1610 493 1611
rect 498 1611 504 1612
rect 498 1610 499 1611
rect 492 1608 499 1610
rect 492 1607 493 1608
rect 487 1606 493 1607
rect 498 1607 499 1608
rect 503 1607 504 1611
rect 498 1606 504 1607
rect 551 1611 557 1612
rect 551 1607 552 1611
rect 556 1610 557 1611
rect 559 1611 565 1612
rect 559 1610 560 1611
rect 556 1608 560 1610
rect 556 1607 557 1608
rect 551 1606 557 1607
rect 559 1607 560 1608
rect 564 1607 565 1611
rect 559 1606 565 1607
rect 614 1611 621 1612
rect 614 1607 615 1611
rect 620 1607 621 1611
rect 614 1606 621 1607
rect 679 1611 685 1612
rect 679 1607 680 1611
rect 684 1610 685 1611
rect 687 1611 693 1612
rect 687 1610 688 1611
rect 684 1608 688 1610
rect 684 1607 685 1608
rect 679 1606 685 1607
rect 687 1607 688 1608
rect 692 1607 693 1611
rect 687 1606 693 1607
rect 742 1611 749 1612
rect 742 1607 743 1611
rect 748 1607 749 1611
rect 742 1606 749 1607
rect 815 1611 821 1612
rect 815 1607 816 1611
rect 820 1610 821 1611
rect 823 1611 829 1612
rect 823 1610 824 1611
rect 820 1608 824 1610
rect 820 1607 821 1608
rect 815 1606 821 1607
rect 823 1607 824 1608
rect 828 1607 829 1611
rect 823 1606 829 1607
rect 887 1611 893 1612
rect 887 1607 888 1611
rect 892 1610 893 1611
rect 895 1611 901 1612
rect 895 1610 896 1611
rect 892 1608 896 1610
rect 892 1607 893 1608
rect 887 1606 893 1607
rect 895 1607 896 1608
rect 900 1607 901 1611
rect 895 1606 901 1607
rect 959 1611 968 1612
rect 959 1607 960 1611
rect 967 1607 968 1611
rect 959 1606 968 1607
rect 1034 1611 1045 1612
rect 1034 1607 1035 1611
rect 1039 1607 1040 1611
rect 1044 1607 1045 1611
rect 1112 1610 1114 1628
rect 1119 1627 1125 1628
rect 1119 1623 1120 1627
rect 1124 1626 1125 1627
rect 1166 1627 1167 1631
rect 1171 1630 1172 1631
rect 1302 1631 1308 1632
rect 1171 1628 1186 1630
rect 1171 1627 1172 1628
rect 1166 1626 1172 1627
rect 1184 1626 1186 1628
rect 1191 1627 1197 1628
rect 1191 1626 1192 1627
rect 1124 1624 1161 1626
rect 1184 1624 1192 1626
rect 1124 1623 1125 1624
rect 1119 1622 1125 1623
rect 1159 1614 1161 1624
rect 1191 1623 1192 1624
rect 1196 1623 1197 1627
rect 1263 1627 1269 1628
rect 1263 1623 1264 1627
rect 1268 1626 1269 1627
rect 1294 1627 1300 1628
rect 1294 1626 1295 1627
rect 1268 1624 1295 1626
rect 1268 1623 1269 1624
rect 1174 1622 1180 1623
rect 1191 1622 1197 1623
rect 1246 1622 1252 1623
rect 1263 1622 1269 1623
rect 1294 1623 1295 1624
rect 1299 1623 1300 1627
rect 1302 1627 1303 1631
rect 1307 1630 1308 1631
rect 1307 1628 1330 1630
rect 1417 1628 1490 1630
rect 1497 1628 1570 1630
rect 1307 1627 1308 1628
rect 1302 1626 1308 1627
rect 1328 1626 1330 1628
rect 1335 1627 1341 1628
rect 1335 1626 1336 1627
rect 1328 1624 1336 1626
rect 1335 1623 1336 1624
rect 1340 1623 1341 1627
rect 1415 1627 1421 1628
rect 1415 1623 1416 1627
rect 1420 1623 1421 1627
rect 1294 1622 1300 1623
rect 1318 1622 1324 1623
rect 1335 1622 1341 1623
rect 1398 1622 1404 1623
rect 1415 1622 1421 1623
rect 1478 1622 1484 1623
rect 1174 1618 1175 1622
rect 1179 1618 1180 1622
rect 1174 1617 1180 1618
rect 1246 1618 1247 1622
rect 1251 1618 1252 1622
rect 1246 1617 1252 1618
rect 1318 1618 1319 1622
rect 1323 1618 1324 1622
rect 1318 1617 1324 1618
rect 1398 1618 1399 1622
rect 1403 1618 1404 1622
rect 1398 1617 1404 1618
rect 1478 1618 1479 1622
rect 1483 1618 1484 1622
rect 1478 1617 1484 1618
rect 1159 1612 1174 1614
rect 1119 1611 1125 1612
rect 1119 1610 1120 1611
rect 1112 1608 1120 1610
rect 1034 1606 1045 1607
rect 1119 1607 1120 1608
rect 1124 1607 1125 1611
rect 1172 1610 1186 1612
rect 1191 1611 1197 1612
rect 1191 1610 1192 1611
rect 1184 1608 1192 1610
rect 1119 1606 1125 1607
rect 1191 1607 1192 1608
rect 1196 1607 1197 1611
rect 1191 1606 1197 1607
rect 1263 1611 1269 1612
rect 1263 1607 1264 1611
rect 1268 1610 1269 1611
rect 1302 1611 1308 1612
rect 1302 1610 1303 1611
rect 1268 1608 1303 1610
rect 1268 1607 1269 1608
rect 1263 1606 1269 1607
rect 1302 1607 1303 1608
rect 1307 1607 1308 1611
rect 1302 1606 1308 1607
rect 1334 1611 1341 1612
rect 1334 1607 1335 1611
rect 1340 1607 1341 1611
rect 1334 1606 1341 1607
rect 1415 1611 1421 1612
rect 1415 1607 1416 1611
rect 1420 1610 1421 1611
rect 1430 1611 1436 1612
rect 1430 1610 1431 1611
rect 1420 1608 1431 1610
rect 1420 1607 1421 1608
rect 1415 1606 1421 1607
rect 1430 1607 1431 1608
rect 1435 1607 1436 1611
rect 1488 1610 1490 1628
rect 1495 1627 1501 1628
rect 1495 1623 1496 1627
rect 1500 1623 1501 1627
rect 1495 1622 1501 1623
rect 1558 1622 1564 1623
rect 1558 1618 1559 1622
rect 1563 1618 1564 1622
rect 1558 1617 1564 1618
rect 1495 1611 1501 1612
rect 1495 1610 1496 1611
rect 1488 1608 1496 1610
rect 1430 1606 1436 1607
rect 1495 1607 1496 1608
rect 1500 1607 1501 1611
rect 1568 1610 1570 1628
rect 1574 1627 1581 1628
rect 1574 1623 1575 1627
rect 1580 1623 1581 1627
rect 1638 1627 1645 1628
rect 1638 1623 1639 1627
rect 1644 1623 1645 1627
rect 1574 1622 1581 1623
rect 1622 1622 1628 1623
rect 1638 1622 1645 1623
rect 1662 1624 1668 1625
rect 1622 1618 1623 1622
rect 1627 1618 1628 1622
rect 1662 1620 1663 1624
rect 1667 1620 1668 1624
rect 1662 1619 1668 1620
rect 1622 1617 1628 1618
rect 1575 1611 1581 1612
rect 1575 1610 1576 1611
rect 1568 1608 1576 1610
rect 1495 1606 1501 1607
rect 1575 1607 1576 1608
rect 1580 1607 1581 1611
rect 1575 1606 1581 1607
rect 1638 1611 1645 1612
rect 1638 1607 1639 1611
rect 1644 1607 1645 1611
rect 1638 1606 1645 1607
rect 1662 1607 1668 1608
rect 110 1602 116 1603
rect 134 1605 140 1606
rect 134 1601 135 1605
rect 139 1601 140 1605
rect 134 1600 140 1601
rect 182 1605 188 1606
rect 182 1601 183 1605
rect 187 1601 188 1605
rect 182 1600 188 1601
rect 246 1605 252 1606
rect 246 1601 247 1605
rect 251 1601 252 1605
rect 246 1600 252 1601
rect 302 1605 308 1606
rect 302 1601 303 1605
rect 307 1601 308 1605
rect 302 1600 308 1601
rect 358 1605 364 1606
rect 358 1601 359 1605
rect 363 1601 364 1605
rect 358 1600 364 1601
rect 414 1605 420 1606
rect 414 1601 415 1605
rect 419 1601 420 1605
rect 414 1600 420 1601
rect 470 1605 476 1606
rect 470 1601 471 1605
rect 475 1601 476 1605
rect 470 1600 476 1601
rect 534 1605 540 1606
rect 534 1601 535 1605
rect 539 1601 540 1605
rect 534 1600 540 1601
rect 598 1605 604 1606
rect 598 1601 599 1605
rect 603 1601 604 1605
rect 598 1600 604 1601
rect 662 1605 668 1606
rect 662 1601 663 1605
rect 667 1601 668 1605
rect 662 1600 668 1601
rect 726 1605 732 1606
rect 726 1601 727 1605
rect 731 1601 732 1605
rect 726 1600 732 1601
rect 798 1605 804 1606
rect 798 1601 799 1605
rect 803 1601 804 1605
rect 798 1600 804 1601
rect 870 1605 876 1606
rect 870 1601 871 1605
rect 875 1601 876 1605
rect 870 1600 876 1601
rect 942 1605 948 1606
rect 942 1601 943 1605
rect 947 1601 948 1605
rect 942 1600 948 1601
rect 1022 1605 1028 1606
rect 1022 1601 1023 1605
rect 1027 1601 1028 1605
rect 1022 1600 1028 1601
rect 1102 1605 1108 1606
rect 1102 1601 1103 1605
rect 1107 1601 1108 1605
rect 1102 1600 1108 1601
rect 1174 1605 1180 1606
rect 1174 1601 1175 1605
rect 1179 1601 1180 1605
rect 1174 1600 1180 1601
rect 1246 1605 1252 1606
rect 1246 1601 1247 1605
rect 1251 1601 1252 1605
rect 1246 1600 1252 1601
rect 1318 1605 1324 1606
rect 1318 1601 1319 1605
rect 1323 1601 1324 1605
rect 1318 1600 1324 1601
rect 1398 1605 1404 1606
rect 1398 1601 1399 1605
rect 1403 1601 1404 1605
rect 1398 1600 1404 1601
rect 1478 1605 1484 1606
rect 1478 1601 1479 1605
rect 1483 1601 1484 1605
rect 1478 1600 1484 1601
rect 1558 1605 1564 1606
rect 1558 1601 1559 1605
rect 1563 1601 1564 1605
rect 1558 1600 1564 1601
rect 1622 1605 1628 1606
rect 1622 1601 1623 1605
rect 1627 1601 1628 1605
rect 1662 1603 1663 1607
rect 1667 1603 1668 1607
rect 1662 1602 1668 1603
rect 1622 1600 1628 1601
rect 198 1599 204 1600
rect 198 1595 199 1599
rect 203 1598 204 1599
rect 203 1596 298 1598
rect 203 1595 204 1596
rect 198 1594 204 1595
rect 134 1591 140 1592
rect 110 1589 116 1590
rect 110 1585 111 1589
rect 115 1585 116 1589
rect 134 1587 135 1591
rect 139 1587 140 1591
rect 134 1586 140 1587
rect 166 1591 172 1592
rect 166 1587 167 1591
rect 171 1587 172 1591
rect 166 1586 172 1587
rect 222 1591 228 1592
rect 222 1587 223 1591
rect 227 1587 228 1591
rect 222 1586 228 1587
rect 278 1591 284 1592
rect 278 1587 279 1591
rect 283 1587 284 1591
rect 278 1586 284 1587
rect 296 1586 298 1596
rect 334 1591 340 1592
rect 334 1587 335 1591
rect 339 1587 340 1591
rect 334 1586 340 1587
rect 382 1591 388 1592
rect 382 1587 383 1591
rect 387 1587 388 1591
rect 382 1586 388 1587
rect 430 1591 436 1592
rect 430 1587 431 1591
rect 435 1587 436 1591
rect 430 1586 436 1587
rect 478 1591 484 1592
rect 478 1587 479 1591
rect 483 1587 484 1591
rect 478 1586 484 1587
rect 534 1591 540 1592
rect 534 1587 535 1591
rect 539 1587 540 1591
rect 534 1586 540 1587
rect 598 1591 604 1592
rect 598 1587 599 1591
rect 603 1587 604 1591
rect 598 1586 604 1587
rect 662 1591 668 1592
rect 662 1587 663 1591
rect 667 1587 668 1591
rect 662 1586 668 1587
rect 726 1591 732 1592
rect 726 1587 727 1591
rect 731 1587 732 1591
rect 726 1586 732 1587
rect 798 1591 804 1592
rect 798 1587 799 1591
rect 803 1587 804 1591
rect 798 1586 804 1587
rect 870 1591 876 1592
rect 870 1587 871 1591
rect 875 1587 876 1591
rect 870 1586 876 1587
rect 950 1591 956 1592
rect 950 1587 951 1591
rect 955 1587 956 1591
rect 950 1586 956 1587
rect 1038 1591 1044 1592
rect 1038 1587 1039 1591
rect 1043 1587 1044 1591
rect 1038 1586 1044 1587
rect 1118 1591 1124 1592
rect 1118 1587 1119 1591
rect 1123 1587 1124 1591
rect 1118 1586 1124 1587
rect 1198 1591 1204 1592
rect 1198 1587 1199 1591
rect 1203 1587 1204 1591
rect 1198 1586 1204 1587
rect 1278 1591 1284 1592
rect 1278 1587 1279 1591
rect 1283 1587 1284 1591
rect 1278 1586 1284 1587
rect 1350 1591 1356 1592
rect 1350 1587 1351 1591
rect 1355 1587 1356 1591
rect 1350 1586 1356 1587
rect 1414 1591 1420 1592
rect 1414 1587 1415 1591
rect 1419 1587 1420 1591
rect 1414 1586 1420 1587
rect 1470 1591 1476 1592
rect 1470 1587 1471 1591
rect 1475 1587 1476 1591
rect 1470 1586 1476 1587
rect 1526 1591 1532 1592
rect 1526 1587 1527 1591
rect 1531 1587 1532 1591
rect 1526 1586 1532 1587
rect 1582 1591 1588 1592
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1622 1591 1628 1592
rect 1622 1587 1623 1591
rect 1627 1587 1628 1591
rect 1622 1586 1628 1587
rect 1662 1589 1668 1590
rect 110 1584 116 1585
rect 295 1585 301 1586
rect 151 1583 157 1584
rect 151 1579 152 1583
rect 156 1582 157 1583
rect 182 1583 189 1584
rect 156 1580 178 1582
rect 156 1579 157 1580
rect 151 1578 157 1579
rect 134 1574 140 1575
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 134 1570 135 1574
rect 139 1570 140 1574
rect 134 1569 140 1570
rect 166 1574 172 1575
rect 166 1570 167 1574
rect 171 1570 172 1574
rect 166 1569 172 1570
rect 110 1567 116 1568
rect 150 1567 157 1568
rect 150 1563 151 1567
rect 156 1563 157 1567
rect 176 1566 178 1580
rect 182 1579 183 1583
rect 188 1579 189 1583
rect 182 1578 189 1579
rect 239 1583 245 1584
rect 239 1579 240 1583
rect 244 1582 245 1583
rect 244 1580 290 1582
rect 295 1581 296 1585
rect 300 1581 301 1585
rect 1662 1585 1663 1589
rect 1667 1585 1668 1589
rect 1662 1584 1668 1585
rect 295 1580 301 1581
rect 351 1583 357 1584
rect 244 1579 245 1580
rect 239 1578 245 1579
rect 222 1574 228 1575
rect 222 1570 223 1574
rect 227 1570 228 1574
rect 222 1569 228 1570
rect 278 1574 284 1575
rect 278 1570 279 1574
rect 283 1570 284 1574
rect 278 1569 284 1570
rect 183 1567 189 1568
rect 183 1566 184 1567
rect 176 1564 184 1566
rect 150 1562 157 1563
rect 183 1563 184 1564
rect 188 1563 189 1567
rect 183 1562 189 1563
rect 234 1567 245 1568
rect 234 1563 235 1567
rect 239 1563 240 1567
rect 244 1563 245 1567
rect 288 1566 290 1580
rect 351 1579 352 1583
rect 356 1582 357 1583
rect 374 1583 380 1584
rect 374 1582 375 1583
rect 356 1580 375 1582
rect 356 1579 357 1580
rect 351 1578 357 1579
rect 374 1579 375 1580
rect 379 1579 380 1583
rect 399 1583 405 1584
rect 399 1582 400 1583
rect 374 1578 380 1579
rect 392 1580 400 1582
rect 334 1574 340 1575
rect 334 1570 335 1574
rect 339 1570 340 1574
rect 334 1569 340 1570
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 295 1567 301 1568
rect 295 1566 296 1567
rect 288 1564 296 1566
rect 234 1562 245 1563
rect 295 1563 296 1564
rect 300 1563 301 1567
rect 295 1562 301 1563
rect 351 1567 357 1568
rect 351 1563 352 1567
rect 356 1566 357 1567
rect 392 1566 394 1580
rect 399 1579 400 1580
rect 404 1579 405 1583
rect 447 1583 453 1584
rect 447 1582 448 1583
rect 399 1578 405 1579
rect 425 1580 448 1582
rect 356 1564 394 1566
rect 399 1567 405 1568
rect 356 1563 357 1564
rect 351 1562 357 1563
rect 399 1563 400 1567
rect 404 1566 405 1567
rect 425 1566 427 1580
rect 447 1579 448 1580
rect 452 1579 453 1583
rect 447 1578 453 1579
rect 490 1583 501 1584
rect 490 1579 491 1583
rect 495 1579 496 1583
rect 500 1579 501 1583
rect 551 1583 557 1584
rect 551 1582 552 1583
rect 490 1578 501 1579
rect 524 1580 552 1582
rect 430 1574 436 1575
rect 430 1570 431 1574
rect 435 1570 436 1574
rect 430 1569 436 1570
rect 478 1574 484 1575
rect 478 1570 479 1574
rect 483 1570 484 1574
rect 478 1569 484 1570
rect 404 1564 427 1566
rect 446 1567 453 1568
rect 404 1563 405 1564
rect 399 1562 405 1563
rect 446 1563 447 1567
rect 452 1563 453 1567
rect 446 1562 453 1563
rect 495 1567 501 1568
rect 495 1563 496 1567
rect 500 1566 501 1567
rect 524 1566 526 1580
rect 551 1579 552 1580
rect 556 1579 557 1583
rect 615 1583 621 1584
rect 615 1582 616 1583
rect 551 1578 557 1579
rect 560 1580 616 1582
rect 534 1574 540 1575
rect 534 1570 535 1574
rect 539 1570 540 1574
rect 534 1569 540 1570
rect 500 1564 526 1566
rect 551 1567 557 1568
rect 500 1563 501 1564
rect 495 1562 501 1563
rect 551 1563 552 1567
rect 556 1566 557 1567
rect 560 1566 562 1580
rect 615 1579 616 1580
rect 620 1579 621 1583
rect 615 1578 621 1579
rect 655 1583 661 1584
rect 655 1579 656 1583
rect 660 1582 661 1583
rect 679 1583 685 1584
rect 679 1582 680 1583
rect 660 1580 680 1582
rect 660 1579 661 1580
rect 655 1578 661 1579
rect 679 1579 680 1580
rect 684 1579 685 1583
rect 743 1583 749 1584
rect 743 1582 744 1583
rect 679 1578 685 1579
rect 716 1580 744 1582
rect 598 1574 604 1575
rect 598 1570 599 1574
rect 603 1570 604 1574
rect 598 1569 604 1570
rect 662 1574 668 1575
rect 662 1570 663 1574
rect 667 1570 668 1574
rect 662 1569 668 1570
rect 556 1564 562 1566
rect 586 1567 592 1568
rect 556 1563 557 1564
rect 551 1562 557 1563
rect 586 1563 587 1567
rect 591 1566 592 1567
rect 615 1567 621 1568
rect 615 1566 616 1567
rect 591 1564 616 1566
rect 591 1563 592 1564
rect 586 1562 592 1563
rect 615 1563 616 1564
rect 620 1563 621 1567
rect 615 1562 621 1563
rect 679 1567 685 1568
rect 679 1563 680 1567
rect 684 1566 685 1567
rect 716 1566 718 1580
rect 743 1579 744 1580
rect 748 1579 749 1583
rect 743 1578 749 1579
rect 814 1583 821 1584
rect 814 1579 815 1583
rect 820 1579 821 1583
rect 887 1583 893 1584
rect 887 1582 888 1583
rect 814 1578 821 1579
rect 856 1580 888 1582
rect 726 1574 732 1575
rect 726 1570 727 1574
rect 731 1570 732 1574
rect 726 1569 732 1570
rect 798 1574 804 1575
rect 856 1574 858 1580
rect 887 1579 888 1580
rect 892 1579 893 1583
rect 887 1578 893 1579
rect 967 1583 973 1584
rect 967 1579 968 1583
rect 972 1582 973 1583
rect 1055 1583 1061 1584
rect 972 1580 1050 1582
rect 972 1579 973 1580
rect 967 1578 973 1579
rect 798 1570 799 1574
rect 803 1570 804 1574
rect 798 1569 804 1570
rect 817 1572 858 1574
rect 870 1574 876 1575
rect 817 1568 819 1572
rect 870 1570 871 1574
rect 875 1570 876 1574
rect 870 1569 876 1570
rect 950 1574 956 1575
rect 950 1570 951 1574
rect 955 1570 956 1574
rect 950 1569 956 1570
rect 1038 1574 1044 1575
rect 1038 1570 1039 1574
rect 1043 1570 1044 1574
rect 1038 1569 1044 1570
rect 684 1564 718 1566
rect 742 1567 749 1568
rect 684 1563 685 1564
rect 679 1562 685 1563
rect 742 1563 743 1567
rect 748 1563 749 1567
rect 742 1562 749 1563
rect 815 1567 821 1568
rect 815 1563 816 1567
rect 820 1563 821 1567
rect 815 1562 821 1563
rect 850 1567 856 1568
rect 850 1563 851 1567
rect 855 1566 856 1567
rect 887 1567 893 1568
rect 887 1566 888 1567
rect 855 1564 888 1566
rect 855 1563 856 1564
rect 850 1562 856 1563
rect 887 1563 888 1564
rect 892 1563 893 1567
rect 887 1562 893 1563
rect 967 1567 973 1568
rect 967 1563 968 1567
rect 972 1566 973 1567
rect 1030 1567 1036 1568
rect 1030 1566 1031 1567
rect 972 1564 1031 1566
rect 972 1563 973 1564
rect 967 1562 973 1563
rect 1030 1563 1031 1564
rect 1035 1563 1036 1567
rect 1048 1566 1050 1580
rect 1055 1579 1056 1583
rect 1060 1582 1061 1583
rect 1135 1583 1141 1584
rect 1060 1580 1098 1582
rect 1060 1579 1061 1580
rect 1055 1578 1061 1579
rect 1055 1567 1061 1568
rect 1055 1566 1056 1567
rect 1048 1564 1056 1566
rect 1030 1562 1036 1563
rect 1055 1563 1056 1564
rect 1060 1563 1061 1567
rect 1096 1566 1098 1580
rect 1135 1579 1136 1583
rect 1140 1582 1141 1583
rect 1210 1583 1221 1584
rect 1140 1580 1161 1582
rect 1140 1579 1141 1580
rect 1135 1578 1141 1579
rect 1118 1574 1124 1575
rect 1118 1570 1119 1574
rect 1123 1570 1124 1574
rect 1118 1569 1124 1570
rect 1135 1567 1141 1568
rect 1135 1566 1136 1567
rect 1096 1564 1136 1566
rect 1055 1562 1061 1563
rect 1135 1563 1136 1564
rect 1140 1563 1141 1567
rect 1159 1566 1161 1580
rect 1210 1579 1211 1583
rect 1215 1579 1216 1583
rect 1220 1579 1221 1583
rect 1210 1578 1221 1579
rect 1294 1583 1301 1584
rect 1294 1579 1295 1583
rect 1300 1579 1301 1583
rect 1294 1578 1301 1579
rect 1362 1583 1373 1584
rect 1362 1579 1363 1583
rect 1367 1579 1368 1583
rect 1372 1579 1373 1583
rect 1362 1578 1373 1579
rect 1431 1583 1437 1584
rect 1431 1579 1432 1583
rect 1436 1582 1437 1583
rect 1482 1583 1493 1584
rect 1436 1580 1462 1582
rect 1436 1579 1437 1580
rect 1431 1578 1437 1579
rect 1198 1574 1204 1575
rect 1198 1570 1199 1574
rect 1203 1570 1204 1574
rect 1198 1569 1204 1570
rect 1278 1574 1284 1575
rect 1278 1570 1279 1574
rect 1283 1570 1284 1574
rect 1278 1569 1284 1570
rect 1350 1574 1356 1575
rect 1350 1570 1351 1574
rect 1355 1570 1356 1574
rect 1350 1569 1356 1570
rect 1414 1574 1420 1575
rect 1414 1570 1415 1574
rect 1419 1570 1420 1574
rect 1414 1569 1420 1570
rect 1215 1567 1221 1568
rect 1215 1566 1216 1567
rect 1159 1564 1216 1566
rect 1135 1562 1141 1563
rect 1215 1563 1216 1564
rect 1220 1563 1221 1567
rect 1215 1562 1221 1563
rect 1286 1567 1292 1568
rect 1286 1563 1287 1567
rect 1291 1566 1292 1567
rect 1295 1567 1301 1568
rect 1295 1566 1296 1567
rect 1291 1564 1296 1566
rect 1291 1563 1292 1564
rect 1286 1562 1292 1563
rect 1295 1563 1296 1564
rect 1300 1563 1301 1567
rect 1295 1562 1301 1563
rect 1367 1567 1373 1568
rect 1367 1563 1368 1567
rect 1372 1566 1373 1567
rect 1430 1567 1437 1568
rect 1372 1564 1427 1566
rect 1372 1563 1373 1564
rect 1367 1562 1373 1563
rect 1425 1558 1427 1564
rect 1430 1563 1431 1567
rect 1436 1563 1437 1567
rect 1460 1566 1462 1580
rect 1482 1579 1483 1583
rect 1487 1579 1488 1583
rect 1492 1579 1493 1583
rect 1482 1578 1493 1579
rect 1543 1583 1552 1584
rect 1543 1579 1544 1583
rect 1551 1579 1552 1583
rect 1599 1583 1605 1584
rect 1599 1582 1600 1583
rect 1543 1578 1552 1579
rect 1576 1580 1600 1582
rect 1470 1574 1476 1575
rect 1470 1570 1471 1574
rect 1475 1570 1476 1574
rect 1470 1569 1476 1570
rect 1526 1574 1532 1575
rect 1526 1570 1527 1574
rect 1531 1570 1532 1574
rect 1526 1569 1532 1570
rect 1487 1567 1493 1568
rect 1487 1566 1488 1567
rect 1460 1564 1488 1566
rect 1430 1562 1437 1563
rect 1487 1563 1488 1564
rect 1492 1563 1493 1567
rect 1487 1562 1493 1563
rect 1543 1567 1549 1568
rect 1543 1563 1544 1567
rect 1548 1566 1549 1567
rect 1576 1566 1578 1580
rect 1599 1579 1600 1580
rect 1604 1579 1605 1583
rect 1599 1578 1605 1579
rect 1639 1583 1645 1584
rect 1639 1579 1640 1583
rect 1644 1582 1645 1583
rect 1647 1583 1653 1584
rect 1647 1582 1648 1583
rect 1644 1580 1648 1582
rect 1644 1579 1645 1580
rect 1639 1578 1645 1579
rect 1647 1579 1648 1580
rect 1652 1579 1653 1583
rect 1647 1578 1653 1579
rect 1582 1574 1588 1575
rect 1582 1570 1583 1574
rect 1587 1570 1588 1574
rect 1582 1569 1588 1570
rect 1622 1574 1628 1575
rect 1622 1570 1623 1574
rect 1627 1570 1628 1574
rect 1622 1569 1628 1570
rect 1662 1572 1668 1573
rect 1662 1568 1663 1572
rect 1667 1568 1668 1572
rect 1548 1564 1578 1566
rect 1598 1567 1605 1568
rect 1548 1563 1549 1564
rect 1543 1562 1549 1563
rect 1598 1563 1599 1567
rect 1604 1563 1605 1567
rect 1598 1562 1605 1563
rect 1638 1567 1645 1568
rect 1662 1567 1668 1568
rect 1638 1563 1639 1567
rect 1644 1563 1645 1567
rect 1638 1562 1645 1563
rect 1482 1559 1488 1560
rect 1482 1558 1483 1559
rect 1425 1556 1483 1558
rect 1482 1555 1483 1556
rect 1487 1555 1488 1559
rect 1482 1554 1488 1555
rect 383 1551 389 1552
rect 153 1548 178 1550
rect 233 1548 274 1550
rect 300 1548 321 1550
rect 151 1547 157 1548
rect 110 1544 116 1545
rect 110 1540 111 1544
rect 115 1540 116 1544
rect 151 1543 152 1547
rect 156 1543 157 1547
rect 110 1539 116 1540
rect 134 1542 140 1543
rect 151 1542 157 1543
rect 166 1542 172 1543
rect 134 1538 135 1542
rect 139 1538 140 1542
rect 134 1537 140 1538
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 150 1531 157 1532
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 150 1527 151 1531
rect 156 1527 157 1531
rect 176 1530 178 1548
rect 182 1547 189 1548
rect 182 1543 183 1547
rect 188 1543 189 1547
rect 231 1547 237 1548
rect 231 1543 232 1547
rect 236 1543 237 1547
rect 182 1542 189 1543
rect 214 1542 220 1543
rect 231 1542 237 1543
rect 262 1542 268 1543
rect 214 1538 215 1542
rect 219 1538 220 1542
rect 214 1537 220 1538
rect 262 1538 263 1542
rect 267 1538 268 1542
rect 262 1537 268 1538
rect 183 1531 189 1532
rect 183 1530 184 1531
rect 176 1528 184 1530
rect 150 1526 157 1527
rect 183 1527 184 1528
rect 188 1527 189 1531
rect 183 1526 189 1527
rect 231 1531 240 1532
rect 231 1527 232 1531
rect 239 1527 240 1531
rect 272 1530 274 1548
rect 279 1547 285 1548
rect 279 1543 280 1547
rect 284 1546 285 1547
rect 300 1546 302 1548
rect 284 1544 302 1546
rect 284 1543 285 1544
rect 279 1542 285 1543
rect 310 1542 316 1543
rect 310 1538 311 1542
rect 315 1538 316 1542
rect 310 1537 316 1538
rect 279 1531 285 1532
rect 279 1530 280 1531
rect 272 1528 280 1530
rect 231 1526 240 1527
rect 279 1527 280 1528
rect 284 1527 285 1531
rect 319 1530 321 1548
rect 327 1547 333 1548
rect 327 1543 328 1547
rect 332 1546 333 1547
rect 350 1547 356 1548
rect 350 1546 351 1547
rect 332 1544 351 1546
rect 332 1543 333 1544
rect 327 1542 333 1543
rect 350 1543 351 1544
rect 355 1543 356 1547
rect 374 1547 381 1548
rect 374 1543 375 1547
rect 380 1543 381 1547
rect 383 1547 384 1551
rect 388 1550 389 1551
rect 431 1551 437 1552
rect 388 1548 427 1550
rect 388 1547 389 1548
rect 383 1546 389 1547
rect 423 1547 429 1548
rect 423 1543 424 1547
rect 428 1543 429 1547
rect 431 1547 432 1551
rect 436 1550 437 1551
rect 479 1551 485 1552
rect 436 1548 466 1550
rect 436 1547 437 1548
rect 431 1546 437 1547
rect 464 1546 466 1548
rect 471 1547 477 1548
rect 471 1546 472 1547
rect 464 1544 472 1546
rect 471 1543 472 1544
rect 476 1543 477 1547
rect 479 1547 480 1551
rect 484 1550 485 1551
rect 535 1551 541 1552
rect 484 1548 522 1550
rect 484 1547 485 1548
rect 479 1546 485 1547
rect 520 1546 522 1548
rect 527 1547 533 1548
rect 527 1546 528 1547
rect 520 1544 528 1546
rect 527 1543 528 1544
rect 532 1543 533 1547
rect 535 1547 536 1551
rect 540 1550 541 1551
rect 663 1551 669 1552
rect 540 1548 578 1550
rect 540 1547 541 1548
rect 535 1546 541 1547
rect 576 1546 578 1548
rect 583 1547 589 1548
rect 583 1546 584 1547
rect 576 1544 584 1546
rect 583 1543 584 1544
rect 588 1543 589 1547
rect 647 1547 653 1548
rect 647 1543 648 1547
rect 652 1546 653 1547
rect 655 1547 661 1548
rect 655 1546 656 1547
rect 652 1544 656 1546
rect 652 1543 653 1544
rect 350 1542 356 1543
rect 358 1542 364 1543
rect 374 1542 381 1543
rect 406 1542 412 1543
rect 423 1542 429 1543
rect 454 1542 460 1543
rect 471 1542 477 1543
rect 510 1542 516 1543
rect 527 1542 533 1543
rect 566 1542 572 1543
rect 583 1542 589 1543
rect 630 1542 636 1543
rect 647 1542 653 1543
rect 655 1543 656 1544
rect 660 1543 661 1547
rect 663 1547 664 1551
rect 668 1550 669 1551
rect 719 1551 725 1552
rect 668 1548 706 1550
rect 668 1547 669 1548
rect 663 1546 669 1547
rect 704 1546 706 1548
rect 711 1547 717 1548
rect 711 1546 712 1547
rect 704 1544 712 1546
rect 711 1543 712 1544
rect 716 1543 717 1547
rect 719 1547 720 1551
rect 724 1550 725 1551
rect 1370 1551 1376 1552
rect 724 1548 770 1550
rect 937 1548 1018 1550
rect 1088 1548 1106 1550
rect 1113 1548 1194 1550
rect 724 1547 725 1548
rect 719 1546 725 1547
rect 768 1546 770 1548
rect 775 1547 781 1548
rect 775 1546 776 1547
rect 768 1544 776 1546
rect 775 1543 776 1544
rect 780 1543 781 1547
rect 847 1547 853 1548
rect 847 1543 848 1547
rect 852 1546 853 1547
rect 894 1547 900 1548
rect 894 1546 895 1547
rect 852 1544 895 1546
rect 852 1543 853 1544
rect 655 1542 661 1543
rect 694 1542 700 1543
rect 711 1542 717 1543
rect 758 1542 764 1543
rect 775 1542 781 1543
rect 830 1542 836 1543
rect 847 1542 853 1543
rect 894 1543 895 1544
rect 899 1543 900 1547
rect 935 1547 941 1548
rect 935 1543 936 1547
rect 940 1543 941 1547
rect 894 1542 900 1543
rect 918 1542 924 1543
rect 935 1542 941 1543
rect 1006 1542 1012 1543
rect 358 1538 359 1542
rect 363 1538 364 1542
rect 358 1537 364 1538
rect 406 1538 407 1542
rect 411 1538 412 1542
rect 406 1537 412 1538
rect 454 1538 455 1542
rect 459 1538 460 1542
rect 454 1537 460 1538
rect 510 1538 511 1542
rect 515 1538 516 1542
rect 510 1537 516 1538
rect 566 1538 567 1542
rect 571 1538 572 1542
rect 566 1537 572 1538
rect 630 1538 631 1542
rect 635 1538 636 1542
rect 630 1537 636 1538
rect 694 1538 695 1542
rect 699 1538 700 1542
rect 694 1537 700 1538
rect 758 1538 759 1542
rect 763 1538 764 1542
rect 758 1537 764 1538
rect 830 1538 831 1542
rect 835 1538 836 1542
rect 830 1537 836 1538
rect 918 1538 919 1542
rect 923 1538 924 1542
rect 918 1537 924 1538
rect 1006 1538 1007 1542
rect 1011 1538 1012 1542
rect 1006 1537 1012 1538
rect 327 1531 333 1532
rect 327 1530 328 1531
rect 319 1528 328 1530
rect 279 1526 285 1527
rect 327 1527 328 1528
rect 332 1527 333 1531
rect 327 1526 333 1527
rect 375 1531 381 1532
rect 375 1527 376 1531
rect 380 1530 381 1531
rect 383 1531 389 1532
rect 383 1530 384 1531
rect 380 1528 384 1530
rect 380 1527 381 1528
rect 375 1526 381 1527
rect 383 1527 384 1528
rect 388 1527 389 1531
rect 383 1526 389 1527
rect 423 1531 429 1532
rect 423 1527 424 1531
rect 428 1530 429 1531
rect 431 1531 437 1532
rect 431 1530 432 1531
rect 428 1528 432 1530
rect 428 1527 429 1528
rect 423 1526 429 1527
rect 431 1527 432 1528
rect 436 1527 437 1531
rect 431 1526 437 1527
rect 471 1531 477 1532
rect 471 1527 472 1531
rect 476 1530 477 1531
rect 479 1531 485 1532
rect 479 1530 480 1531
rect 476 1528 480 1530
rect 476 1527 477 1528
rect 471 1526 477 1527
rect 479 1527 480 1528
rect 484 1527 485 1531
rect 479 1526 485 1527
rect 527 1531 533 1532
rect 527 1527 528 1531
rect 532 1530 533 1531
rect 535 1531 541 1532
rect 535 1530 536 1531
rect 532 1528 536 1530
rect 532 1527 533 1528
rect 527 1526 533 1527
rect 535 1527 536 1528
rect 540 1527 541 1531
rect 535 1526 541 1527
rect 583 1531 592 1532
rect 583 1527 584 1531
rect 591 1527 592 1531
rect 583 1526 592 1527
rect 647 1531 653 1532
rect 647 1527 648 1531
rect 652 1530 653 1531
rect 663 1531 669 1532
rect 663 1530 664 1531
rect 652 1528 664 1530
rect 652 1527 653 1528
rect 647 1526 653 1527
rect 663 1527 664 1528
rect 668 1527 669 1531
rect 663 1526 669 1527
rect 711 1531 717 1532
rect 711 1527 712 1531
rect 716 1530 717 1531
rect 719 1531 725 1532
rect 719 1530 720 1531
rect 716 1528 720 1530
rect 716 1527 717 1528
rect 711 1526 717 1527
rect 719 1527 720 1528
rect 724 1527 725 1531
rect 719 1526 725 1527
rect 770 1531 781 1532
rect 770 1527 771 1531
rect 775 1527 776 1531
rect 780 1527 781 1531
rect 770 1526 781 1527
rect 847 1531 856 1532
rect 847 1527 848 1531
rect 855 1527 856 1531
rect 847 1526 856 1527
rect 935 1531 941 1532
rect 935 1527 936 1531
rect 940 1530 941 1531
rect 958 1531 964 1532
rect 958 1530 959 1531
rect 940 1528 959 1530
rect 940 1527 941 1528
rect 935 1526 941 1527
rect 958 1527 959 1528
rect 963 1527 964 1531
rect 1016 1530 1018 1548
rect 1023 1547 1029 1548
rect 1023 1543 1024 1547
rect 1028 1546 1029 1547
rect 1088 1546 1090 1548
rect 1028 1544 1090 1546
rect 1028 1543 1029 1544
rect 1023 1542 1029 1543
rect 1094 1542 1100 1543
rect 1094 1538 1095 1542
rect 1099 1538 1100 1542
rect 1094 1537 1100 1538
rect 1023 1531 1029 1532
rect 1023 1530 1024 1531
rect 1016 1528 1024 1530
rect 958 1526 964 1527
rect 1023 1527 1024 1528
rect 1028 1527 1029 1531
rect 1104 1530 1106 1548
rect 1111 1547 1117 1548
rect 1111 1543 1112 1547
rect 1116 1543 1117 1547
rect 1111 1542 1117 1543
rect 1182 1542 1188 1543
rect 1182 1538 1183 1542
rect 1187 1538 1188 1542
rect 1182 1537 1188 1538
rect 1111 1531 1117 1532
rect 1111 1530 1112 1531
rect 1104 1528 1112 1530
rect 1023 1526 1029 1527
rect 1111 1527 1112 1528
rect 1116 1527 1117 1531
rect 1192 1530 1194 1548
rect 1199 1547 1205 1548
rect 1199 1543 1200 1547
rect 1204 1546 1205 1547
rect 1210 1547 1216 1548
rect 1210 1546 1211 1547
rect 1204 1544 1211 1546
rect 1204 1543 1205 1544
rect 1199 1542 1205 1543
rect 1210 1543 1211 1544
rect 1215 1543 1216 1547
rect 1279 1547 1285 1548
rect 1279 1543 1280 1547
rect 1284 1546 1285 1547
rect 1326 1547 1332 1548
rect 1326 1546 1327 1547
rect 1284 1544 1327 1546
rect 1284 1543 1285 1544
rect 1210 1542 1216 1543
rect 1262 1542 1268 1543
rect 1279 1542 1285 1543
rect 1326 1543 1327 1544
rect 1331 1543 1332 1547
rect 1351 1547 1357 1548
rect 1351 1543 1352 1547
rect 1356 1546 1357 1547
rect 1362 1547 1368 1548
rect 1362 1546 1363 1547
rect 1356 1544 1363 1546
rect 1356 1543 1357 1544
rect 1326 1542 1332 1543
rect 1334 1542 1340 1543
rect 1351 1542 1357 1543
rect 1362 1543 1363 1544
rect 1367 1543 1368 1547
rect 1370 1547 1371 1551
rect 1375 1550 1376 1551
rect 1431 1551 1437 1552
rect 1375 1548 1427 1550
rect 1375 1547 1376 1548
rect 1370 1546 1376 1547
rect 1423 1547 1429 1548
rect 1423 1543 1424 1547
rect 1428 1543 1429 1547
rect 1431 1547 1432 1551
rect 1436 1550 1437 1551
rect 1495 1551 1501 1552
rect 1436 1548 1482 1550
rect 1436 1547 1437 1548
rect 1431 1546 1437 1547
rect 1480 1546 1482 1548
rect 1487 1547 1493 1548
rect 1487 1546 1488 1547
rect 1480 1544 1488 1546
rect 1487 1543 1488 1544
rect 1492 1543 1493 1547
rect 1495 1547 1496 1551
rect 1500 1550 1501 1551
rect 1551 1551 1557 1552
rect 1500 1548 1547 1550
rect 1500 1547 1501 1548
rect 1495 1546 1501 1547
rect 1543 1547 1549 1548
rect 1543 1543 1544 1547
rect 1548 1543 1549 1547
rect 1551 1547 1552 1551
rect 1556 1550 1557 1551
rect 1556 1548 1594 1550
rect 1556 1547 1557 1548
rect 1551 1546 1557 1547
rect 1592 1546 1594 1548
rect 1599 1547 1605 1548
rect 1599 1546 1600 1547
rect 1592 1544 1600 1546
rect 1599 1543 1600 1544
rect 1604 1543 1605 1547
rect 1639 1547 1645 1548
rect 1639 1543 1640 1547
rect 1644 1546 1645 1547
rect 1647 1547 1653 1548
rect 1647 1546 1648 1547
rect 1644 1544 1648 1546
rect 1644 1543 1645 1544
rect 1362 1542 1368 1543
rect 1406 1542 1412 1543
rect 1423 1542 1429 1543
rect 1470 1542 1476 1543
rect 1487 1542 1493 1543
rect 1526 1542 1532 1543
rect 1543 1542 1549 1543
rect 1582 1542 1588 1543
rect 1599 1542 1605 1543
rect 1622 1542 1628 1543
rect 1639 1542 1645 1543
rect 1647 1543 1648 1544
rect 1652 1543 1653 1547
rect 1647 1542 1653 1543
rect 1662 1544 1668 1545
rect 1262 1538 1263 1542
rect 1267 1538 1268 1542
rect 1262 1537 1268 1538
rect 1334 1538 1335 1542
rect 1339 1538 1340 1542
rect 1334 1537 1340 1538
rect 1406 1538 1407 1542
rect 1411 1538 1412 1542
rect 1406 1537 1412 1538
rect 1470 1538 1471 1542
rect 1475 1538 1476 1542
rect 1470 1537 1476 1538
rect 1526 1538 1527 1542
rect 1531 1538 1532 1542
rect 1526 1537 1532 1538
rect 1582 1538 1583 1542
rect 1587 1538 1588 1542
rect 1582 1537 1588 1538
rect 1622 1538 1623 1542
rect 1627 1538 1628 1542
rect 1662 1540 1663 1544
rect 1667 1540 1668 1544
rect 1662 1539 1668 1540
rect 1622 1537 1628 1538
rect 1199 1531 1205 1532
rect 1199 1530 1200 1531
rect 1192 1528 1200 1530
rect 1111 1526 1117 1527
rect 1199 1527 1200 1528
rect 1204 1527 1205 1531
rect 1199 1526 1205 1527
rect 1279 1531 1285 1532
rect 1279 1527 1280 1531
rect 1284 1527 1285 1531
rect 1279 1526 1285 1527
rect 1351 1531 1357 1532
rect 1351 1527 1352 1531
rect 1356 1530 1357 1531
rect 1370 1531 1376 1532
rect 1370 1530 1371 1531
rect 1356 1528 1371 1530
rect 1356 1527 1357 1528
rect 1351 1526 1357 1527
rect 1370 1527 1371 1528
rect 1375 1527 1376 1531
rect 1370 1526 1376 1527
rect 1423 1531 1429 1532
rect 1423 1527 1424 1531
rect 1428 1530 1429 1531
rect 1431 1531 1437 1532
rect 1431 1530 1432 1531
rect 1428 1528 1432 1530
rect 1428 1527 1429 1528
rect 1423 1526 1429 1527
rect 1431 1527 1432 1528
rect 1436 1527 1437 1531
rect 1431 1526 1437 1527
rect 1487 1531 1493 1532
rect 1487 1527 1488 1531
rect 1492 1530 1493 1531
rect 1495 1531 1501 1532
rect 1495 1530 1496 1531
rect 1492 1528 1496 1530
rect 1492 1527 1493 1528
rect 1487 1526 1493 1527
rect 1495 1527 1496 1528
rect 1500 1527 1501 1531
rect 1495 1526 1501 1527
rect 1543 1531 1549 1532
rect 1543 1527 1544 1531
rect 1548 1530 1549 1531
rect 1551 1531 1557 1532
rect 1551 1530 1552 1531
rect 1548 1528 1552 1530
rect 1548 1527 1549 1528
rect 1543 1526 1549 1527
rect 1551 1527 1552 1528
rect 1556 1527 1557 1531
rect 1551 1526 1557 1527
rect 1598 1531 1605 1532
rect 1598 1527 1599 1531
rect 1604 1527 1605 1531
rect 1598 1526 1605 1527
rect 1638 1531 1645 1532
rect 1638 1527 1639 1531
rect 1644 1527 1645 1531
rect 1638 1526 1645 1527
rect 1662 1527 1668 1528
rect 110 1522 116 1523
rect 134 1525 140 1526
rect 134 1521 135 1525
rect 139 1521 140 1525
rect 134 1520 140 1521
rect 166 1525 172 1526
rect 166 1521 167 1525
rect 171 1521 172 1525
rect 166 1520 172 1521
rect 214 1525 220 1526
rect 214 1521 215 1525
rect 219 1521 220 1525
rect 214 1520 220 1521
rect 262 1525 268 1526
rect 262 1521 263 1525
rect 267 1521 268 1525
rect 262 1520 268 1521
rect 310 1525 316 1526
rect 310 1521 311 1525
rect 315 1521 316 1525
rect 310 1520 316 1521
rect 358 1525 364 1526
rect 358 1521 359 1525
rect 363 1521 364 1525
rect 358 1520 364 1521
rect 406 1525 412 1526
rect 406 1521 407 1525
rect 411 1521 412 1525
rect 406 1520 412 1521
rect 454 1525 460 1526
rect 454 1521 455 1525
rect 459 1521 460 1525
rect 454 1520 460 1521
rect 510 1525 516 1526
rect 510 1521 511 1525
rect 515 1521 516 1525
rect 510 1520 516 1521
rect 566 1525 572 1526
rect 566 1521 567 1525
rect 571 1521 572 1525
rect 566 1520 572 1521
rect 630 1525 636 1526
rect 630 1521 631 1525
rect 635 1521 636 1525
rect 630 1520 636 1521
rect 694 1525 700 1526
rect 694 1521 695 1525
rect 699 1521 700 1525
rect 694 1520 700 1521
rect 758 1525 764 1526
rect 758 1521 759 1525
rect 763 1521 764 1525
rect 758 1520 764 1521
rect 830 1525 836 1526
rect 830 1521 831 1525
rect 835 1521 836 1525
rect 830 1520 836 1521
rect 918 1525 924 1526
rect 918 1521 919 1525
rect 923 1521 924 1525
rect 918 1520 924 1521
rect 1006 1525 1012 1526
rect 1006 1521 1007 1525
rect 1011 1521 1012 1525
rect 1006 1520 1012 1521
rect 1094 1525 1100 1526
rect 1094 1521 1095 1525
rect 1099 1521 1100 1525
rect 1094 1520 1100 1521
rect 1182 1525 1188 1526
rect 1182 1521 1183 1525
rect 1187 1521 1188 1525
rect 1182 1520 1188 1521
rect 1262 1525 1268 1526
rect 1262 1521 1263 1525
rect 1267 1521 1268 1525
rect 1262 1520 1268 1521
rect 1334 1525 1340 1526
rect 1334 1521 1335 1525
rect 1339 1521 1340 1525
rect 1334 1520 1340 1521
rect 1406 1525 1412 1526
rect 1406 1521 1407 1525
rect 1411 1521 1412 1525
rect 1406 1520 1412 1521
rect 1470 1525 1476 1526
rect 1470 1521 1471 1525
rect 1475 1521 1476 1525
rect 1470 1520 1476 1521
rect 1526 1525 1532 1526
rect 1526 1521 1527 1525
rect 1531 1521 1532 1525
rect 1526 1520 1532 1521
rect 1582 1525 1588 1526
rect 1582 1521 1583 1525
rect 1587 1521 1588 1525
rect 1582 1520 1588 1521
rect 1622 1525 1628 1526
rect 1622 1521 1623 1525
rect 1627 1521 1628 1525
rect 1662 1523 1663 1527
rect 1667 1523 1668 1527
rect 1662 1522 1668 1523
rect 1622 1520 1628 1521
rect 350 1515 356 1516
rect 350 1511 351 1515
rect 355 1514 356 1515
rect 1326 1515 1332 1516
rect 355 1512 438 1514
rect 355 1511 356 1512
rect 350 1510 356 1511
rect 134 1507 140 1508
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 134 1503 135 1507
rect 139 1503 140 1507
rect 134 1502 140 1503
rect 166 1507 172 1508
rect 166 1503 167 1507
rect 171 1503 172 1507
rect 166 1502 172 1503
rect 222 1507 228 1508
rect 222 1503 223 1507
rect 227 1503 228 1507
rect 222 1502 228 1503
rect 294 1507 300 1508
rect 294 1503 295 1507
rect 299 1503 300 1507
rect 294 1502 300 1503
rect 374 1507 380 1508
rect 374 1503 375 1507
rect 379 1503 380 1507
rect 374 1502 380 1503
rect 110 1500 116 1501
rect 151 1499 157 1500
rect 151 1495 152 1499
rect 156 1498 157 1499
rect 183 1499 189 1500
rect 156 1496 178 1498
rect 156 1495 157 1496
rect 151 1494 157 1495
rect 134 1490 140 1491
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 134 1486 135 1490
rect 139 1486 140 1490
rect 134 1485 140 1486
rect 166 1490 172 1491
rect 166 1486 167 1490
rect 171 1486 172 1490
rect 176 1490 178 1496
rect 183 1495 184 1499
rect 188 1498 189 1499
rect 239 1499 245 1500
rect 188 1496 234 1498
rect 188 1495 189 1496
rect 183 1494 189 1495
rect 182 1491 188 1492
rect 182 1490 183 1491
rect 176 1488 183 1490
rect 182 1487 183 1488
rect 187 1487 188 1491
rect 182 1486 188 1487
rect 222 1490 228 1491
rect 222 1486 223 1490
rect 227 1486 228 1490
rect 166 1485 172 1486
rect 222 1485 228 1486
rect 110 1483 116 1484
rect 150 1483 157 1484
rect 150 1479 151 1483
rect 156 1479 157 1483
rect 150 1478 157 1479
rect 183 1483 189 1484
rect 183 1479 184 1483
rect 188 1479 189 1483
rect 232 1482 234 1496
rect 239 1495 240 1499
rect 244 1498 245 1499
rect 311 1499 317 1500
rect 244 1496 306 1498
rect 244 1495 245 1496
rect 239 1494 245 1495
rect 294 1490 300 1491
rect 294 1486 295 1490
rect 299 1486 300 1490
rect 294 1485 300 1486
rect 239 1483 245 1484
rect 239 1482 240 1483
rect 232 1480 240 1482
rect 183 1478 189 1479
rect 239 1479 240 1480
rect 244 1479 245 1483
rect 304 1482 306 1496
rect 311 1495 312 1499
rect 316 1498 317 1499
rect 391 1499 397 1500
rect 316 1496 321 1498
rect 316 1495 317 1496
rect 311 1494 317 1495
rect 311 1483 317 1484
rect 311 1482 312 1483
rect 304 1480 312 1482
rect 239 1478 245 1479
rect 311 1479 312 1480
rect 316 1479 317 1483
rect 319 1482 321 1496
rect 391 1495 392 1499
rect 396 1498 397 1499
rect 436 1498 438 1512
rect 1326 1511 1327 1515
rect 1331 1514 1332 1515
rect 1331 1512 1550 1514
rect 1331 1511 1332 1512
rect 1326 1510 1332 1511
rect 454 1507 460 1508
rect 454 1503 455 1507
rect 459 1503 460 1507
rect 454 1502 460 1503
rect 526 1507 532 1508
rect 526 1503 527 1507
rect 531 1503 532 1507
rect 526 1502 532 1503
rect 598 1507 604 1508
rect 598 1503 599 1507
rect 603 1503 604 1507
rect 598 1502 604 1503
rect 670 1507 676 1508
rect 670 1503 671 1507
rect 675 1503 676 1507
rect 670 1502 676 1503
rect 742 1507 748 1508
rect 742 1503 743 1507
rect 747 1503 748 1507
rect 742 1502 748 1503
rect 814 1507 820 1508
rect 814 1503 815 1507
rect 819 1503 820 1507
rect 814 1502 820 1503
rect 878 1507 884 1508
rect 878 1503 879 1507
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 942 1507 948 1508
rect 942 1503 943 1507
rect 947 1503 948 1507
rect 942 1502 948 1503
rect 1006 1507 1012 1508
rect 1006 1503 1007 1507
rect 1011 1503 1012 1507
rect 1006 1502 1012 1503
rect 1062 1507 1068 1508
rect 1062 1503 1063 1507
rect 1067 1503 1068 1507
rect 1062 1502 1068 1503
rect 1110 1507 1116 1508
rect 1110 1503 1111 1507
rect 1115 1503 1116 1507
rect 1110 1502 1116 1503
rect 1150 1507 1156 1508
rect 1150 1503 1151 1507
rect 1155 1503 1156 1507
rect 1150 1502 1156 1503
rect 1182 1507 1188 1508
rect 1182 1503 1183 1507
rect 1187 1503 1188 1507
rect 1182 1502 1188 1503
rect 1214 1507 1220 1508
rect 1214 1503 1215 1507
rect 1219 1503 1220 1507
rect 1214 1502 1220 1503
rect 1254 1507 1260 1508
rect 1254 1503 1255 1507
rect 1259 1503 1260 1507
rect 1254 1502 1260 1503
rect 1294 1507 1300 1508
rect 1294 1503 1295 1507
rect 1299 1503 1300 1507
rect 1294 1502 1300 1503
rect 1350 1507 1356 1508
rect 1350 1503 1351 1507
rect 1355 1503 1356 1507
rect 1350 1502 1356 1503
rect 1414 1507 1420 1508
rect 1414 1503 1415 1507
rect 1419 1503 1420 1507
rect 1414 1502 1420 1503
rect 1486 1507 1492 1508
rect 1486 1503 1487 1507
rect 1491 1503 1492 1507
rect 1486 1502 1492 1503
rect 471 1499 477 1500
rect 471 1498 472 1499
rect 396 1496 434 1498
rect 436 1496 472 1498
rect 396 1495 397 1496
rect 391 1494 397 1495
rect 374 1490 380 1491
rect 374 1486 375 1490
rect 379 1486 380 1490
rect 374 1485 380 1486
rect 391 1483 397 1484
rect 391 1482 392 1483
rect 319 1480 392 1482
rect 311 1478 317 1479
rect 391 1479 392 1480
rect 396 1479 397 1483
rect 432 1482 434 1496
rect 471 1495 472 1496
rect 476 1495 477 1499
rect 471 1494 477 1495
rect 542 1499 549 1500
rect 542 1495 543 1499
rect 548 1495 549 1499
rect 615 1499 621 1500
rect 615 1498 616 1499
rect 542 1494 549 1495
rect 580 1496 616 1498
rect 454 1490 460 1491
rect 454 1486 455 1490
rect 459 1486 460 1490
rect 454 1485 460 1486
rect 526 1490 532 1491
rect 526 1486 527 1490
rect 531 1486 532 1490
rect 526 1485 532 1486
rect 471 1483 477 1484
rect 471 1482 472 1483
rect 432 1480 472 1482
rect 391 1478 397 1479
rect 471 1479 472 1480
rect 476 1479 477 1483
rect 471 1478 477 1479
rect 543 1483 549 1484
rect 543 1479 544 1483
rect 548 1482 549 1483
rect 580 1482 582 1496
rect 615 1495 616 1496
rect 620 1495 621 1499
rect 687 1499 693 1500
rect 687 1498 688 1499
rect 615 1494 621 1495
rect 652 1496 688 1498
rect 598 1490 604 1491
rect 598 1486 599 1490
rect 603 1486 604 1490
rect 598 1485 604 1486
rect 548 1480 582 1482
rect 615 1483 621 1484
rect 548 1479 549 1480
rect 543 1478 549 1479
rect 615 1479 616 1483
rect 620 1482 621 1483
rect 652 1482 654 1496
rect 687 1495 688 1496
rect 692 1495 693 1499
rect 687 1494 693 1495
rect 759 1499 765 1500
rect 759 1495 760 1499
rect 764 1498 765 1499
rect 831 1499 837 1500
rect 764 1496 811 1498
rect 764 1495 765 1496
rect 759 1494 765 1495
rect 770 1491 776 1492
rect 670 1490 676 1491
rect 670 1486 671 1490
rect 675 1486 676 1490
rect 670 1485 676 1486
rect 742 1490 748 1491
rect 770 1490 771 1491
rect 742 1486 743 1490
rect 747 1486 748 1490
rect 742 1485 748 1486
rect 752 1488 771 1490
rect 620 1480 654 1482
rect 687 1483 693 1484
rect 620 1479 621 1480
rect 615 1478 621 1479
rect 687 1479 688 1483
rect 692 1482 693 1483
rect 752 1482 754 1488
rect 770 1487 771 1488
rect 775 1487 776 1491
rect 770 1486 776 1487
rect 692 1480 754 1482
rect 759 1483 765 1484
rect 692 1479 693 1480
rect 687 1478 693 1479
rect 759 1479 760 1483
rect 764 1482 765 1483
rect 798 1483 804 1484
rect 798 1482 799 1483
rect 764 1480 799 1482
rect 764 1479 765 1480
rect 759 1478 765 1479
rect 798 1479 799 1480
rect 803 1479 804 1483
rect 809 1482 811 1496
rect 831 1495 832 1499
rect 836 1498 837 1499
rect 894 1499 901 1500
rect 836 1496 866 1498
rect 836 1495 837 1496
rect 831 1494 837 1495
rect 814 1490 820 1491
rect 814 1486 815 1490
rect 819 1486 820 1490
rect 814 1485 820 1486
rect 831 1483 837 1484
rect 831 1482 832 1483
rect 809 1480 832 1482
rect 798 1478 804 1479
rect 831 1479 832 1480
rect 836 1479 837 1483
rect 864 1482 866 1496
rect 894 1495 895 1499
rect 900 1495 901 1499
rect 894 1494 901 1495
rect 959 1499 965 1500
rect 959 1495 960 1499
rect 964 1498 965 1499
rect 974 1499 980 1500
rect 974 1498 975 1499
rect 964 1496 975 1498
rect 964 1495 965 1496
rect 959 1494 965 1495
rect 974 1495 975 1496
rect 979 1495 980 1499
rect 974 1494 980 1495
rect 1023 1499 1029 1500
rect 1023 1495 1024 1499
rect 1028 1498 1029 1499
rect 1079 1499 1085 1500
rect 1028 1496 1054 1498
rect 1028 1495 1029 1496
rect 1023 1494 1029 1495
rect 878 1490 884 1491
rect 878 1486 879 1490
rect 883 1486 884 1490
rect 878 1485 884 1486
rect 942 1490 948 1491
rect 942 1486 943 1490
rect 947 1486 948 1490
rect 942 1485 948 1486
rect 1006 1490 1012 1491
rect 1006 1486 1007 1490
rect 1011 1486 1012 1490
rect 1006 1485 1012 1486
rect 895 1483 901 1484
rect 895 1482 896 1483
rect 864 1480 896 1482
rect 831 1478 837 1479
rect 895 1479 896 1480
rect 900 1479 901 1483
rect 895 1478 901 1479
rect 958 1483 965 1484
rect 958 1479 959 1483
rect 964 1479 965 1483
rect 958 1478 965 1479
rect 1023 1483 1032 1484
rect 1023 1479 1024 1483
rect 1031 1479 1032 1483
rect 1052 1482 1054 1496
rect 1079 1495 1080 1499
rect 1084 1498 1085 1499
rect 1127 1499 1133 1500
rect 1084 1496 1106 1498
rect 1084 1495 1085 1496
rect 1079 1494 1085 1495
rect 1062 1490 1068 1491
rect 1062 1486 1063 1490
rect 1067 1486 1068 1490
rect 1062 1485 1068 1486
rect 1079 1483 1085 1484
rect 1079 1482 1080 1483
rect 1052 1480 1080 1482
rect 1023 1478 1032 1479
rect 1079 1479 1080 1480
rect 1084 1479 1085 1483
rect 1104 1482 1106 1496
rect 1127 1495 1128 1499
rect 1132 1498 1133 1499
rect 1167 1499 1173 1500
rect 1132 1496 1161 1498
rect 1132 1495 1133 1496
rect 1127 1494 1133 1495
rect 1110 1490 1116 1491
rect 1110 1486 1111 1490
rect 1115 1486 1116 1490
rect 1110 1485 1116 1486
rect 1150 1490 1156 1491
rect 1150 1486 1151 1490
rect 1155 1486 1156 1490
rect 1150 1485 1156 1486
rect 1127 1483 1133 1484
rect 1127 1482 1128 1483
rect 1104 1480 1128 1482
rect 1079 1478 1085 1479
rect 1127 1479 1128 1480
rect 1132 1479 1133 1483
rect 1159 1482 1161 1496
rect 1167 1495 1168 1499
rect 1172 1498 1173 1499
rect 1199 1499 1205 1500
rect 1172 1496 1194 1498
rect 1172 1495 1173 1496
rect 1167 1494 1173 1495
rect 1182 1490 1188 1491
rect 1182 1486 1183 1490
rect 1187 1486 1188 1490
rect 1182 1485 1188 1486
rect 1167 1483 1173 1484
rect 1167 1482 1168 1483
rect 1159 1480 1168 1482
rect 1127 1478 1133 1479
rect 1167 1479 1168 1480
rect 1172 1479 1173 1483
rect 1192 1482 1194 1496
rect 1199 1495 1200 1499
rect 1204 1498 1205 1499
rect 1230 1499 1237 1500
rect 1204 1496 1226 1498
rect 1204 1495 1205 1496
rect 1199 1494 1205 1495
rect 1214 1490 1220 1491
rect 1214 1486 1215 1490
rect 1219 1486 1220 1490
rect 1214 1485 1220 1486
rect 1199 1483 1205 1484
rect 1199 1482 1200 1483
rect 1192 1480 1200 1482
rect 1167 1478 1173 1479
rect 1199 1479 1200 1480
rect 1204 1479 1205 1483
rect 1224 1482 1226 1496
rect 1230 1495 1231 1499
rect 1236 1495 1237 1499
rect 1230 1494 1237 1495
rect 1271 1499 1277 1500
rect 1271 1495 1272 1499
rect 1276 1498 1277 1499
rect 1311 1499 1317 1500
rect 1276 1496 1290 1498
rect 1276 1495 1277 1496
rect 1271 1494 1277 1495
rect 1254 1490 1260 1491
rect 1254 1486 1255 1490
rect 1259 1486 1260 1490
rect 1254 1485 1260 1486
rect 1231 1483 1237 1484
rect 1231 1482 1232 1483
rect 1224 1480 1232 1482
rect 1199 1478 1205 1479
rect 1231 1479 1232 1480
rect 1236 1479 1237 1483
rect 1231 1478 1237 1479
rect 1271 1483 1277 1484
rect 1271 1479 1272 1483
rect 1276 1482 1277 1483
rect 1288 1482 1290 1496
rect 1311 1495 1312 1499
rect 1316 1498 1317 1499
rect 1367 1499 1373 1500
rect 1316 1496 1342 1498
rect 1316 1495 1317 1496
rect 1311 1494 1317 1495
rect 1294 1490 1300 1491
rect 1294 1486 1295 1490
rect 1299 1486 1300 1490
rect 1294 1485 1300 1486
rect 1311 1483 1317 1484
rect 1311 1482 1312 1483
rect 1276 1480 1286 1482
rect 1288 1480 1312 1482
rect 1276 1479 1277 1480
rect 1271 1478 1277 1479
rect 185 1474 187 1478
rect 238 1475 244 1476
rect 238 1474 239 1475
rect 185 1472 239 1474
rect 238 1471 239 1472
rect 243 1471 244 1475
rect 1230 1475 1236 1476
rect 1230 1474 1231 1475
rect 238 1470 244 1471
rect 1177 1472 1231 1474
rect 551 1467 557 1468
rect 153 1464 178 1466
rect 241 1464 306 1466
rect 319 1464 386 1466
rect 151 1463 157 1464
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 151 1459 152 1463
rect 156 1459 157 1463
rect 110 1455 116 1456
rect 134 1458 140 1459
rect 151 1458 157 1459
rect 166 1458 172 1459
rect 134 1454 135 1458
rect 139 1454 140 1458
rect 134 1453 140 1454
rect 166 1454 167 1458
rect 171 1454 172 1458
rect 166 1453 172 1454
rect 150 1447 157 1448
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 150 1443 151 1447
rect 156 1443 157 1447
rect 176 1446 178 1464
rect 182 1463 189 1464
rect 182 1459 183 1463
rect 188 1459 189 1463
rect 239 1463 245 1464
rect 239 1459 240 1463
rect 244 1459 245 1463
rect 182 1458 189 1459
rect 222 1458 228 1459
rect 239 1458 245 1459
rect 294 1458 300 1459
rect 222 1454 223 1458
rect 227 1454 228 1458
rect 222 1453 228 1454
rect 294 1454 295 1458
rect 299 1454 300 1458
rect 294 1453 300 1454
rect 183 1447 189 1448
rect 183 1446 184 1447
rect 176 1444 184 1446
rect 150 1442 157 1443
rect 183 1443 184 1444
rect 188 1443 189 1447
rect 183 1442 189 1443
rect 238 1447 245 1448
rect 238 1443 239 1447
rect 244 1443 245 1447
rect 304 1446 306 1464
rect 311 1463 317 1464
rect 311 1459 312 1463
rect 316 1462 317 1463
rect 319 1462 321 1464
rect 316 1460 321 1462
rect 316 1459 317 1460
rect 311 1458 317 1459
rect 374 1458 380 1459
rect 374 1454 375 1458
rect 379 1454 380 1458
rect 374 1453 380 1454
rect 311 1447 317 1448
rect 311 1446 312 1447
rect 304 1444 312 1446
rect 238 1442 245 1443
rect 311 1443 312 1444
rect 316 1443 317 1447
rect 384 1446 386 1464
rect 391 1463 397 1464
rect 391 1459 392 1463
rect 396 1462 397 1463
rect 462 1463 468 1464
rect 396 1460 434 1462
rect 396 1459 397 1460
rect 391 1458 397 1459
rect 432 1450 434 1460
rect 462 1459 463 1463
rect 467 1462 468 1463
rect 471 1463 477 1464
rect 471 1462 472 1463
rect 467 1460 472 1462
rect 467 1459 468 1460
rect 454 1458 460 1459
rect 462 1458 468 1459
rect 471 1459 472 1460
rect 476 1459 477 1463
rect 542 1463 549 1464
rect 542 1459 543 1463
rect 548 1459 549 1463
rect 551 1463 552 1467
rect 556 1466 557 1467
rect 623 1467 629 1468
rect 556 1464 619 1466
rect 556 1463 557 1464
rect 551 1462 557 1463
rect 615 1463 621 1464
rect 615 1459 616 1463
rect 620 1459 621 1463
rect 623 1463 624 1467
rect 628 1466 629 1467
rect 687 1467 693 1468
rect 628 1464 683 1466
rect 628 1463 629 1464
rect 623 1462 629 1463
rect 679 1463 685 1464
rect 679 1459 680 1463
rect 684 1459 685 1463
rect 687 1463 688 1467
rect 692 1466 693 1467
rect 743 1467 749 1468
rect 692 1464 730 1466
rect 692 1463 693 1464
rect 687 1462 693 1463
rect 728 1462 730 1464
rect 735 1463 741 1464
rect 735 1462 736 1463
rect 728 1460 736 1462
rect 735 1459 736 1460
rect 740 1459 741 1463
rect 743 1463 744 1467
rect 748 1466 749 1467
rect 748 1464 803 1466
rect 896 1464 914 1466
rect 921 1464 970 1466
rect 1064 1464 1082 1466
rect 1113 1464 1130 1466
rect 1177 1464 1179 1472
rect 1230 1471 1231 1472
rect 1235 1471 1236 1475
rect 1284 1474 1286 1480
rect 1311 1479 1312 1480
rect 1316 1479 1317 1483
rect 1340 1482 1342 1496
rect 1367 1495 1368 1499
rect 1372 1498 1373 1499
rect 1431 1499 1437 1500
rect 1372 1496 1402 1498
rect 1372 1495 1373 1496
rect 1367 1494 1373 1495
rect 1350 1490 1356 1491
rect 1350 1486 1351 1490
rect 1355 1486 1356 1490
rect 1350 1485 1356 1486
rect 1367 1483 1373 1484
rect 1367 1482 1368 1483
rect 1340 1480 1368 1482
rect 1311 1478 1317 1479
rect 1367 1479 1368 1480
rect 1372 1479 1373 1483
rect 1400 1482 1402 1496
rect 1431 1495 1432 1499
rect 1436 1498 1437 1499
rect 1503 1499 1509 1500
rect 1436 1496 1470 1498
rect 1436 1495 1437 1496
rect 1431 1494 1437 1495
rect 1414 1490 1420 1491
rect 1414 1486 1415 1490
rect 1419 1486 1420 1490
rect 1414 1485 1420 1486
rect 1431 1483 1437 1484
rect 1431 1482 1432 1483
rect 1400 1480 1432 1482
rect 1367 1478 1373 1479
rect 1431 1479 1432 1480
rect 1436 1479 1437 1483
rect 1468 1482 1470 1496
rect 1503 1495 1504 1499
rect 1508 1498 1509 1499
rect 1548 1498 1550 1512
rect 1566 1507 1572 1508
rect 1566 1503 1567 1507
rect 1571 1503 1572 1507
rect 1566 1502 1572 1503
rect 1622 1507 1628 1508
rect 1622 1503 1623 1507
rect 1627 1503 1628 1507
rect 1622 1502 1628 1503
rect 1662 1505 1668 1506
rect 1662 1501 1663 1505
rect 1667 1501 1668 1505
rect 1662 1500 1668 1501
rect 1583 1499 1589 1500
rect 1583 1498 1584 1499
rect 1508 1496 1546 1498
rect 1548 1496 1584 1498
rect 1508 1495 1509 1496
rect 1503 1494 1509 1495
rect 1486 1490 1492 1491
rect 1486 1486 1487 1490
rect 1491 1486 1492 1490
rect 1486 1485 1492 1486
rect 1503 1483 1509 1484
rect 1503 1482 1504 1483
rect 1468 1480 1504 1482
rect 1431 1478 1437 1479
rect 1503 1479 1504 1480
rect 1508 1479 1509 1483
rect 1544 1482 1546 1496
rect 1583 1495 1584 1496
rect 1588 1495 1589 1499
rect 1583 1494 1589 1495
rect 1639 1499 1645 1500
rect 1639 1495 1640 1499
rect 1644 1498 1645 1499
rect 1647 1499 1653 1500
rect 1647 1498 1648 1499
rect 1644 1496 1648 1498
rect 1644 1495 1645 1496
rect 1639 1494 1645 1495
rect 1647 1495 1648 1496
rect 1652 1495 1653 1499
rect 1647 1494 1653 1495
rect 1566 1490 1572 1491
rect 1566 1486 1567 1490
rect 1571 1486 1572 1490
rect 1566 1485 1572 1486
rect 1622 1490 1628 1491
rect 1622 1486 1623 1490
rect 1627 1486 1628 1490
rect 1622 1485 1628 1486
rect 1662 1488 1668 1489
rect 1662 1484 1663 1488
rect 1667 1484 1668 1488
rect 1583 1483 1589 1484
rect 1583 1482 1584 1483
rect 1544 1480 1584 1482
rect 1503 1478 1509 1479
rect 1583 1479 1584 1480
rect 1588 1479 1589 1483
rect 1583 1478 1589 1479
rect 1638 1483 1645 1484
rect 1662 1483 1668 1484
rect 1638 1479 1639 1483
rect 1644 1479 1645 1483
rect 1638 1478 1645 1479
rect 1494 1475 1500 1476
rect 1494 1474 1495 1475
rect 1284 1472 1495 1474
rect 1230 1470 1236 1471
rect 1494 1471 1495 1472
rect 1499 1471 1500 1475
rect 1494 1470 1500 1471
rect 1183 1467 1189 1468
rect 748 1463 749 1464
rect 743 1462 749 1463
rect 799 1463 805 1464
rect 799 1459 800 1463
rect 804 1459 805 1463
rect 863 1463 869 1464
rect 863 1459 864 1463
rect 868 1462 869 1463
rect 896 1462 898 1464
rect 868 1460 898 1462
rect 868 1459 869 1460
rect 471 1458 477 1459
rect 526 1458 532 1459
rect 542 1458 549 1459
rect 598 1458 604 1459
rect 615 1458 621 1459
rect 662 1458 668 1459
rect 679 1458 685 1459
rect 718 1458 724 1459
rect 735 1458 741 1459
rect 782 1458 788 1459
rect 799 1458 805 1459
rect 846 1458 852 1459
rect 863 1458 869 1459
rect 902 1458 908 1459
rect 454 1454 455 1458
rect 459 1454 460 1458
rect 454 1453 460 1454
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 598 1454 599 1458
rect 603 1454 604 1458
rect 598 1453 604 1454
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 782 1454 783 1458
rect 787 1454 788 1458
rect 782 1453 788 1454
rect 846 1454 847 1458
rect 851 1454 852 1458
rect 846 1453 852 1454
rect 902 1454 903 1458
rect 907 1454 908 1458
rect 902 1453 908 1454
rect 912 1450 914 1464
rect 919 1463 925 1464
rect 919 1459 920 1463
rect 924 1459 925 1463
rect 919 1458 925 1459
rect 958 1458 964 1459
rect 958 1454 959 1458
rect 963 1454 964 1458
rect 958 1453 964 1454
rect 432 1448 454 1450
rect 912 1448 923 1450
rect 391 1447 397 1448
rect 391 1446 392 1447
rect 384 1444 392 1446
rect 311 1442 317 1443
rect 391 1443 392 1444
rect 396 1443 397 1447
rect 452 1446 466 1448
rect 471 1447 477 1448
rect 471 1446 472 1447
rect 464 1444 472 1446
rect 391 1442 397 1443
rect 471 1443 472 1444
rect 476 1443 477 1447
rect 471 1442 477 1443
rect 543 1447 549 1448
rect 543 1443 544 1447
rect 548 1446 549 1447
rect 551 1447 557 1448
rect 551 1446 552 1447
rect 548 1444 552 1446
rect 548 1443 549 1444
rect 543 1442 549 1443
rect 551 1443 552 1444
rect 556 1443 557 1447
rect 551 1442 557 1443
rect 615 1447 621 1448
rect 615 1443 616 1447
rect 620 1446 621 1447
rect 623 1447 629 1448
rect 623 1446 624 1447
rect 620 1444 624 1446
rect 620 1443 621 1444
rect 615 1442 621 1443
rect 623 1443 624 1444
rect 628 1443 629 1447
rect 623 1442 629 1443
rect 679 1447 685 1448
rect 679 1443 680 1447
rect 684 1446 685 1447
rect 687 1447 693 1448
rect 687 1446 688 1447
rect 684 1444 688 1446
rect 684 1443 685 1444
rect 679 1442 685 1443
rect 687 1443 688 1444
rect 692 1443 693 1447
rect 687 1442 693 1443
rect 735 1447 741 1448
rect 735 1443 736 1447
rect 740 1446 741 1447
rect 743 1447 749 1448
rect 743 1446 744 1447
rect 740 1444 744 1446
rect 740 1443 741 1444
rect 735 1442 741 1443
rect 743 1443 744 1444
rect 748 1443 749 1447
rect 743 1442 749 1443
rect 798 1447 805 1448
rect 798 1443 799 1447
rect 804 1443 805 1447
rect 798 1442 805 1443
rect 863 1447 869 1448
rect 863 1443 864 1447
rect 868 1446 869 1447
rect 894 1447 900 1448
rect 894 1446 895 1447
rect 868 1444 895 1446
rect 868 1443 869 1444
rect 863 1442 869 1443
rect 894 1443 895 1444
rect 899 1443 900 1447
rect 894 1442 900 1443
rect 919 1447 925 1448
rect 919 1443 920 1447
rect 924 1443 925 1447
rect 968 1446 970 1464
rect 974 1463 981 1464
rect 974 1459 975 1463
rect 980 1459 981 1463
rect 1031 1463 1037 1464
rect 1031 1459 1032 1463
rect 1036 1462 1037 1463
rect 1064 1462 1066 1464
rect 1036 1460 1066 1462
rect 1036 1459 1037 1460
rect 974 1458 981 1459
rect 1014 1458 1020 1459
rect 1031 1458 1037 1459
rect 1070 1458 1076 1459
rect 1014 1454 1015 1458
rect 1019 1454 1020 1458
rect 1014 1453 1020 1454
rect 1070 1454 1071 1458
rect 1075 1454 1076 1458
rect 1070 1453 1076 1454
rect 975 1447 981 1448
rect 975 1446 976 1447
rect 968 1444 976 1446
rect 919 1442 925 1443
rect 975 1443 976 1444
rect 980 1443 981 1447
rect 975 1442 981 1443
rect 1026 1447 1037 1448
rect 1026 1443 1027 1447
rect 1031 1443 1032 1447
rect 1036 1443 1037 1447
rect 1080 1446 1082 1464
rect 1087 1463 1093 1464
rect 1087 1459 1088 1463
rect 1092 1462 1093 1463
rect 1113 1462 1115 1464
rect 1092 1460 1115 1462
rect 1092 1459 1093 1460
rect 1087 1458 1093 1459
rect 1118 1458 1124 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 1087 1447 1093 1448
rect 1087 1446 1088 1447
rect 1080 1444 1088 1446
rect 1026 1442 1037 1443
rect 1087 1443 1088 1444
rect 1092 1443 1093 1447
rect 1128 1446 1130 1464
rect 1135 1463 1141 1464
rect 1135 1459 1136 1463
rect 1140 1462 1141 1463
rect 1146 1463 1152 1464
rect 1146 1462 1147 1463
rect 1140 1460 1147 1462
rect 1140 1459 1141 1460
rect 1135 1458 1141 1459
rect 1146 1459 1147 1460
rect 1151 1459 1152 1463
rect 1175 1463 1181 1464
rect 1175 1459 1176 1463
rect 1180 1459 1181 1463
rect 1183 1463 1184 1467
rect 1188 1466 1189 1467
rect 1231 1467 1237 1468
rect 1188 1464 1218 1466
rect 1188 1463 1189 1464
rect 1183 1462 1189 1463
rect 1216 1462 1218 1464
rect 1223 1463 1229 1464
rect 1223 1462 1224 1463
rect 1216 1460 1224 1462
rect 1223 1459 1224 1460
rect 1228 1459 1229 1463
rect 1231 1463 1232 1467
rect 1236 1466 1237 1467
rect 1287 1467 1293 1468
rect 1236 1464 1274 1466
rect 1236 1463 1237 1464
rect 1231 1462 1237 1463
rect 1272 1462 1274 1464
rect 1279 1463 1285 1464
rect 1279 1462 1280 1463
rect 1272 1460 1280 1462
rect 1279 1459 1280 1460
rect 1284 1459 1285 1463
rect 1287 1463 1288 1467
rect 1292 1466 1293 1467
rect 1351 1467 1357 1468
rect 1292 1464 1338 1466
rect 1292 1463 1293 1464
rect 1287 1462 1293 1463
rect 1336 1462 1338 1464
rect 1343 1463 1349 1464
rect 1343 1462 1344 1463
rect 1336 1460 1344 1462
rect 1343 1459 1344 1460
rect 1348 1459 1349 1463
rect 1351 1463 1352 1467
rect 1356 1466 1357 1467
rect 1423 1467 1429 1468
rect 1356 1464 1419 1466
rect 1356 1463 1357 1464
rect 1351 1462 1357 1463
rect 1415 1463 1421 1464
rect 1415 1459 1416 1463
rect 1420 1459 1421 1463
rect 1423 1463 1424 1467
rect 1428 1466 1429 1467
rect 1428 1464 1499 1466
rect 1428 1463 1429 1464
rect 1423 1462 1429 1463
rect 1495 1463 1501 1464
rect 1495 1459 1496 1463
rect 1500 1459 1501 1463
rect 1570 1463 1581 1464
rect 1570 1459 1571 1463
rect 1575 1459 1576 1463
rect 1580 1459 1581 1463
rect 1639 1463 1645 1464
rect 1639 1459 1640 1463
rect 1644 1462 1645 1463
rect 1647 1463 1653 1464
rect 1647 1462 1648 1463
rect 1644 1460 1648 1462
rect 1644 1459 1645 1460
rect 1146 1458 1152 1459
rect 1158 1458 1164 1459
rect 1175 1458 1181 1459
rect 1206 1458 1212 1459
rect 1223 1458 1229 1459
rect 1262 1458 1268 1459
rect 1279 1458 1285 1459
rect 1326 1458 1332 1459
rect 1343 1458 1349 1459
rect 1398 1458 1404 1459
rect 1415 1458 1421 1459
rect 1478 1458 1484 1459
rect 1495 1458 1501 1459
rect 1558 1458 1564 1459
rect 1570 1458 1581 1459
rect 1622 1458 1628 1459
rect 1639 1458 1645 1459
rect 1647 1459 1648 1460
rect 1652 1459 1653 1463
rect 1647 1458 1653 1459
rect 1662 1460 1668 1461
rect 1158 1454 1159 1458
rect 1163 1454 1164 1458
rect 1158 1453 1164 1454
rect 1206 1454 1207 1458
rect 1211 1454 1212 1458
rect 1206 1453 1212 1454
rect 1262 1454 1263 1458
rect 1267 1454 1268 1458
rect 1262 1453 1268 1454
rect 1326 1454 1327 1458
rect 1331 1454 1332 1458
rect 1326 1453 1332 1454
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1662 1456 1663 1460
rect 1667 1456 1668 1460
rect 1662 1455 1668 1456
rect 1622 1453 1628 1454
rect 1135 1447 1141 1448
rect 1135 1446 1136 1447
rect 1128 1444 1136 1446
rect 1087 1442 1093 1443
rect 1135 1443 1136 1444
rect 1140 1443 1141 1447
rect 1135 1442 1141 1443
rect 1175 1447 1181 1448
rect 1175 1443 1176 1447
rect 1180 1446 1181 1447
rect 1183 1447 1189 1448
rect 1183 1446 1184 1447
rect 1180 1444 1184 1446
rect 1180 1443 1181 1444
rect 1175 1442 1181 1443
rect 1183 1443 1184 1444
rect 1188 1443 1189 1447
rect 1183 1442 1189 1443
rect 1223 1447 1229 1448
rect 1223 1443 1224 1447
rect 1228 1446 1229 1447
rect 1231 1447 1237 1448
rect 1231 1446 1232 1447
rect 1228 1444 1232 1446
rect 1228 1443 1229 1444
rect 1223 1442 1229 1443
rect 1231 1443 1232 1444
rect 1236 1443 1237 1447
rect 1231 1442 1237 1443
rect 1279 1447 1285 1448
rect 1279 1443 1280 1447
rect 1284 1446 1285 1447
rect 1287 1447 1293 1448
rect 1287 1446 1288 1447
rect 1284 1444 1288 1446
rect 1284 1443 1285 1444
rect 1279 1442 1285 1443
rect 1287 1443 1288 1444
rect 1292 1443 1293 1447
rect 1287 1442 1293 1443
rect 1343 1447 1349 1448
rect 1343 1443 1344 1447
rect 1348 1446 1349 1447
rect 1351 1447 1357 1448
rect 1351 1446 1352 1447
rect 1348 1444 1352 1446
rect 1348 1443 1349 1444
rect 1343 1442 1349 1443
rect 1351 1443 1352 1444
rect 1356 1443 1357 1447
rect 1351 1442 1357 1443
rect 1415 1447 1421 1448
rect 1415 1443 1416 1447
rect 1420 1446 1421 1447
rect 1423 1447 1429 1448
rect 1423 1446 1424 1447
rect 1420 1444 1424 1446
rect 1420 1443 1421 1444
rect 1415 1442 1421 1443
rect 1423 1443 1424 1444
rect 1428 1443 1429 1447
rect 1423 1442 1429 1443
rect 1494 1447 1501 1448
rect 1494 1443 1495 1447
rect 1500 1443 1501 1447
rect 1494 1442 1501 1443
rect 1575 1447 1581 1448
rect 1575 1443 1576 1447
rect 1580 1443 1581 1447
rect 1575 1442 1581 1443
rect 1638 1447 1645 1448
rect 1638 1443 1639 1447
rect 1644 1443 1645 1447
rect 1638 1442 1645 1443
rect 1662 1443 1668 1444
rect 110 1438 116 1439
rect 134 1441 140 1442
rect 134 1437 135 1441
rect 139 1437 140 1441
rect 134 1436 140 1437
rect 166 1441 172 1442
rect 166 1437 167 1441
rect 171 1437 172 1441
rect 166 1436 172 1437
rect 222 1441 228 1442
rect 222 1437 223 1441
rect 227 1437 228 1441
rect 222 1436 228 1437
rect 294 1441 300 1442
rect 294 1437 295 1441
rect 299 1437 300 1441
rect 294 1436 300 1437
rect 374 1441 380 1442
rect 374 1437 375 1441
rect 379 1437 380 1441
rect 374 1436 380 1437
rect 454 1441 460 1442
rect 454 1437 455 1441
rect 459 1437 460 1441
rect 454 1436 460 1437
rect 526 1441 532 1442
rect 526 1437 527 1441
rect 531 1437 532 1441
rect 526 1436 532 1437
rect 598 1441 604 1442
rect 598 1437 599 1441
rect 603 1437 604 1441
rect 598 1436 604 1437
rect 662 1441 668 1442
rect 662 1437 663 1441
rect 667 1437 668 1441
rect 662 1436 668 1437
rect 718 1441 724 1442
rect 718 1437 719 1441
rect 723 1437 724 1441
rect 718 1436 724 1437
rect 782 1441 788 1442
rect 782 1437 783 1441
rect 787 1437 788 1441
rect 782 1436 788 1437
rect 846 1441 852 1442
rect 846 1437 847 1441
rect 851 1437 852 1441
rect 846 1436 852 1437
rect 902 1441 908 1442
rect 902 1437 903 1441
rect 907 1437 908 1441
rect 902 1436 908 1437
rect 958 1441 964 1442
rect 958 1437 959 1441
rect 963 1437 964 1441
rect 958 1436 964 1437
rect 1014 1441 1020 1442
rect 1014 1437 1015 1441
rect 1019 1437 1020 1441
rect 1014 1436 1020 1437
rect 1070 1441 1076 1442
rect 1070 1437 1071 1441
rect 1075 1437 1076 1441
rect 1070 1436 1076 1437
rect 1118 1441 1124 1442
rect 1118 1437 1119 1441
rect 1123 1437 1124 1441
rect 1118 1436 1124 1437
rect 1158 1441 1164 1442
rect 1158 1437 1159 1441
rect 1163 1437 1164 1441
rect 1158 1436 1164 1437
rect 1206 1441 1212 1442
rect 1206 1437 1207 1441
rect 1211 1437 1212 1441
rect 1206 1436 1212 1437
rect 1262 1441 1268 1442
rect 1262 1437 1263 1441
rect 1267 1437 1268 1441
rect 1262 1436 1268 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1326 1436 1332 1437
rect 1398 1441 1404 1442
rect 1398 1437 1399 1441
rect 1403 1437 1404 1441
rect 1398 1436 1404 1437
rect 1478 1441 1484 1442
rect 1478 1437 1479 1441
rect 1483 1437 1484 1441
rect 1478 1436 1484 1437
rect 1558 1441 1564 1442
rect 1558 1437 1559 1441
rect 1563 1437 1564 1441
rect 1558 1436 1564 1437
rect 1522 1435 1528 1436
rect 1146 1431 1152 1432
rect 1146 1427 1147 1431
rect 1151 1430 1152 1431
rect 1522 1431 1523 1435
rect 1527 1434 1528 1435
rect 1577 1434 1579 1442
rect 1622 1441 1628 1442
rect 1622 1437 1623 1441
rect 1627 1437 1628 1441
rect 1662 1439 1663 1443
rect 1667 1439 1668 1443
rect 1662 1438 1668 1439
rect 1622 1436 1628 1437
rect 1527 1432 1579 1434
rect 1527 1431 1528 1432
rect 1522 1430 1528 1431
rect 1151 1428 1306 1430
rect 1151 1427 1152 1428
rect 1146 1426 1152 1427
rect 134 1423 140 1424
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 134 1419 135 1423
rect 139 1419 140 1423
rect 134 1418 140 1419
rect 166 1423 172 1424
rect 166 1419 167 1423
rect 171 1419 172 1423
rect 166 1418 172 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1419 220 1423
rect 214 1418 220 1419
rect 286 1423 292 1424
rect 286 1419 287 1423
rect 291 1419 292 1423
rect 286 1418 292 1419
rect 358 1423 364 1424
rect 358 1419 359 1423
rect 363 1419 364 1423
rect 358 1418 364 1419
rect 438 1423 444 1424
rect 438 1419 439 1423
rect 443 1419 444 1423
rect 438 1418 444 1419
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 598 1423 604 1424
rect 598 1419 599 1423
rect 603 1419 604 1423
rect 598 1418 604 1419
rect 678 1423 684 1424
rect 678 1419 679 1423
rect 683 1419 684 1423
rect 678 1418 684 1419
rect 758 1423 764 1424
rect 758 1419 759 1423
rect 763 1419 764 1423
rect 758 1418 764 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 902 1423 908 1424
rect 902 1419 903 1423
rect 907 1419 908 1423
rect 902 1418 908 1419
rect 966 1423 972 1424
rect 966 1419 967 1423
rect 971 1419 972 1423
rect 966 1418 972 1419
rect 1030 1423 1036 1424
rect 1030 1419 1031 1423
rect 1035 1419 1036 1423
rect 1030 1418 1036 1419
rect 1102 1423 1108 1424
rect 1102 1419 1103 1423
rect 1107 1419 1108 1423
rect 1102 1418 1108 1419
rect 1166 1423 1172 1424
rect 1166 1419 1167 1423
rect 1171 1419 1172 1423
rect 1166 1418 1172 1419
rect 1230 1423 1236 1424
rect 1230 1419 1231 1423
rect 1235 1419 1236 1423
rect 1230 1418 1236 1419
rect 1294 1423 1300 1424
rect 1294 1419 1295 1423
rect 1299 1419 1300 1423
rect 1294 1418 1300 1419
rect 110 1416 116 1417
rect 151 1415 157 1416
rect 151 1411 152 1415
rect 156 1414 157 1415
rect 183 1415 189 1416
rect 156 1412 178 1414
rect 156 1411 157 1412
rect 151 1410 157 1411
rect 134 1406 140 1407
rect 110 1404 116 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 134 1402 135 1406
rect 139 1402 140 1406
rect 134 1401 140 1402
rect 166 1406 172 1407
rect 166 1402 167 1406
rect 171 1402 172 1406
rect 166 1401 172 1402
rect 110 1399 116 1400
rect 150 1399 157 1400
rect 150 1395 151 1399
rect 156 1395 157 1399
rect 176 1398 178 1412
rect 183 1411 184 1415
rect 188 1414 189 1415
rect 230 1415 237 1416
rect 188 1412 226 1414
rect 188 1411 189 1412
rect 183 1410 189 1411
rect 214 1406 220 1407
rect 214 1402 215 1406
rect 219 1402 220 1406
rect 214 1401 220 1402
rect 183 1399 189 1400
rect 183 1398 184 1399
rect 176 1396 184 1398
rect 150 1394 157 1395
rect 183 1395 184 1396
rect 188 1395 189 1399
rect 224 1398 226 1412
rect 230 1411 231 1415
rect 236 1411 237 1415
rect 230 1410 237 1411
rect 303 1415 309 1416
rect 303 1411 304 1415
rect 308 1414 309 1415
rect 375 1415 381 1416
rect 308 1412 321 1414
rect 308 1411 309 1412
rect 303 1410 309 1411
rect 286 1406 292 1407
rect 286 1402 287 1406
rect 291 1402 292 1406
rect 286 1401 292 1402
rect 231 1399 237 1400
rect 231 1398 232 1399
rect 224 1396 232 1398
rect 183 1394 189 1395
rect 231 1395 232 1396
rect 236 1395 237 1399
rect 231 1394 237 1395
rect 242 1399 248 1400
rect 242 1395 243 1399
rect 247 1398 248 1399
rect 303 1399 309 1400
rect 303 1398 304 1399
rect 247 1396 304 1398
rect 247 1395 248 1396
rect 242 1394 248 1395
rect 303 1395 304 1396
rect 308 1395 309 1399
rect 319 1398 321 1412
rect 375 1411 376 1415
rect 380 1414 381 1415
rect 455 1415 461 1416
rect 380 1412 418 1414
rect 380 1411 381 1412
rect 375 1410 381 1411
rect 358 1406 364 1407
rect 358 1402 359 1406
rect 363 1402 364 1406
rect 358 1401 364 1402
rect 375 1399 381 1400
rect 375 1398 376 1399
rect 319 1396 376 1398
rect 303 1394 309 1395
rect 375 1395 376 1396
rect 380 1395 381 1399
rect 416 1398 418 1412
rect 455 1411 456 1415
rect 460 1411 461 1415
rect 455 1410 461 1411
rect 535 1415 541 1416
rect 535 1411 536 1415
rect 540 1414 541 1415
rect 615 1415 621 1416
rect 540 1412 578 1414
rect 540 1411 541 1412
rect 535 1410 541 1411
rect 438 1406 444 1407
rect 438 1402 439 1406
rect 443 1402 444 1406
rect 438 1401 444 1402
rect 518 1406 524 1407
rect 518 1402 519 1406
rect 523 1402 524 1406
rect 518 1401 524 1402
rect 455 1399 461 1400
rect 455 1398 456 1399
rect 416 1396 456 1398
rect 375 1394 381 1395
rect 455 1395 456 1396
rect 460 1395 461 1399
rect 455 1394 461 1395
rect 535 1399 541 1400
rect 535 1395 536 1399
rect 540 1398 541 1399
rect 576 1398 578 1412
rect 615 1411 616 1415
rect 620 1414 621 1415
rect 695 1415 701 1416
rect 620 1412 690 1414
rect 620 1411 621 1412
rect 615 1410 621 1411
rect 598 1406 604 1407
rect 598 1402 599 1406
rect 603 1402 604 1406
rect 598 1401 604 1402
rect 678 1406 684 1407
rect 678 1402 679 1406
rect 683 1402 684 1406
rect 678 1401 684 1402
rect 615 1399 621 1400
rect 615 1398 616 1399
rect 540 1396 562 1398
rect 576 1396 616 1398
rect 540 1395 541 1396
rect 535 1394 541 1395
rect 560 1390 562 1396
rect 615 1395 616 1396
rect 620 1395 621 1399
rect 688 1398 690 1412
rect 695 1411 696 1415
rect 700 1414 701 1415
rect 750 1415 756 1416
rect 750 1414 751 1415
rect 700 1412 751 1414
rect 700 1411 701 1412
rect 695 1410 701 1411
rect 750 1411 751 1412
rect 755 1411 756 1415
rect 750 1410 756 1411
rect 770 1415 781 1416
rect 770 1411 771 1415
rect 775 1411 776 1415
rect 780 1411 781 1415
rect 847 1415 853 1416
rect 847 1414 848 1415
rect 770 1410 781 1411
rect 816 1412 848 1414
rect 758 1406 764 1407
rect 758 1402 759 1406
rect 763 1402 764 1406
rect 758 1401 764 1402
rect 695 1399 701 1400
rect 695 1398 696 1399
rect 688 1396 696 1398
rect 615 1394 621 1395
rect 695 1395 696 1396
rect 700 1395 701 1399
rect 695 1394 701 1395
rect 775 1399 781 1400
rect 775 1395 776 1399
rect 780 1398 781 1399
rect 816 1398 818 1412
rect 847 1411 848 1412
rect 852 1411 853 1415
rect 919 1415 925 1416
rect 919 1414 920 1415
rect 847 1410 853 1411
rect 884 1412 920 1414
rect 830 1406 836 1407
rect 830 1402 831 1406
rect 835 1402 836 1406
rect 830 1401 836 1402
rect 780 1396 818 1398
rect 847 1399 853 1400
rect 780 1395 781 1396
rect 775 1394 781 1395
rect 847 1395 848 1399
rect 852 1398 853 1399
rect 884 1398 886 1412
rect 919 1411 920 1412
rect 924 1411 925 1415
rect 919 1410 925 1411
rect 983 1415 989 1416
rect 983 1411 984 1415
rect 988 1414 989 1415
rect 1047 1415 1053 1416
rect 988 1412 1042 1414
rect 988 1411 989 1412
rect 983 1410 989 1411
rect 902 1406 908 1407
rect 902 1402 903 1406
rect 907 1402 908 1406
rect 902 1401 908 1402
rect 966 1406 972 1407
rect 966 1402 967 1406
rect 971 1402 972 1406
rect 966 1401 972 1402
rect 1030 1406 1036 1407
rect 1030 1402 1031 1406
rect 1035 1402 1036 1406
rect 1030 1401 1036 1402
rect 852 1396 886 1398
rect 894 1399 900 1400
rect 852 1395 853 1396
rect 847 1394 853 1395
rect 894 1395 895 1399
rect 899 1398 900 1399
rect 919 1399 925 1400
rect 919 1398 920 1399
rect 899 1396 920 1398
rect 899 1395 900 1396
rect 894 1394 900 1395
rect 919 1395 920 1396
rect 924 1395 925 1399
rect 919 1394 925 1395
rect 983 1399 989 1400
rect 983 1395 984 1399
rect 988 1395 989 1399
rect 1040 1398 1042 1412
rect 1047 1411 1048 1415
rect 1052 1414 1053 1415
rect 1119 1415 1125 1416
rect 1052 1412 1114 1414
rect 1052 1411 1053 1412
rect 1047 1410 1053 1411
rect 1102 1406 1108 1407
rect 1102 1402 1103 1406
rect 1107 1402 1108 1406
rect 1102 1401 1108 1402
rect 1047 1399 1053 1400
rect 1047 1398 1048 1399
rect 1040 1396 1048 1398
rect 983 1394 989 1395
rect 1047 1395 1048 1396
rect 1052 1395 1053 1399
rect 1112 1398 1114 1412
rect 1119 1411 1120 1415
rect 1124 1414 1125 1415
rect 1183 1415 1189 1416
rect 1124 1412 1161 1414
rect 1124 1411 1125 1412
rect 1119 1410 1125 1411
rect 1119 1399 1125 1400
rect 1119 1398 1120 1399
rect 1112 1396 1120 1398
rect 1047 1394 1053 1395
rect 1119 1395 1120 1396
rect 1124 1395 1125 1399
rect 1159 1398 1161 1412
rect 1183 1411 1184 1415
rect 1188 1414 1189 1415
rect 1247 1415 1253 1416
rect 1188 1412 1218 1414
rect 1188 1411 1189 1412
rect 1183 1410 1189 1411
rect 1166 1406 1172 1407
rect 1166 1402 1167 1406
rect 1171 1402 1172 1406
rect 1166 1401 1172 1402
rect 1183 1399 1189 1400
rect 1183 1398 1184 1399
rect 1159 1396 1184 1398
rect 1119 1394 1125 1395
rect 1183 1395 1184 1396
rect 1188 1395 1189 1399
rect 1216 1398 1218 1412
rect 1247 1411 1248 1415
rect 1252 1414 1253 1415
rect 1304 1414 1306 1428
rect 1358 1423 1364 1424
rect 1358 1419 1359 1423
rect 1363 1419 1364 1423
rect 1358 1418 1364 1419
rect 1414 1423 1420 1424
rect 1414 1419 1415 1423
rect 1419 1419 1420 1423
rect 1414 1418 1420 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1502 1423 1508 1424
rect 1502 1419 1503 1423
rect 1507 1419 1508 1423
rect 1502 1418 1508 1419
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1590 1423 1596 1424
rect 1590 1419 1591 1423
rect 1595 1419 1596 1423
rect 1590 1418 1596 1419
rect 1622 1423 1628 1424
rect 1622 1419 1623 1423
rect 1627 1419 1628 1423
rect 1622 1418 1628 1419
rect 1662 1421 1668 1422
rect 1662 1417 1663 1421
rect 1667 1417 1668 1421
rect 1662 1416 1668 1417
rect 1311 1415 1317 1416
rect 1311 1414 1312 1415
rect 1252 1412 1282 1414
rect 1304 1412 1312 1414
rect 1252 1411 1253 1412
rect 1247 1410 1253 1411
rect 1230 1406 1236 1407
rect 1230 1402 1231 1406
rect 1235 1402 1236 1406
rect 1230 1401 1236 1402
rect 1247 1399 1253 1400
rect 1247 1398 1248 1399
rect 1216 1396 1248 1398
rect 1183 1394 1189 1395
rect 1247 1395 1248 1396
rect 1252 1395 1253 1399
rect 1280 1398 1282 1412
rect 1311 1411 1312 1412
rect 1316 1411 1317 1415
rect 1311 1410 1317 1411
rect 1375 1415 1381 1416
rect 1375 1411 1376 1415
rect 1380 1414 1381 1415
rect 1431 1415 1437 1416
rect 1380 1412 1406 1414
rect 1380 1411 1381 1412
rect 1375 1410 1381 1411
rect 1294 1406 1300 1407
rect 1294 1402 1295 1406
rect 1299 1402 1300 1406
rect 1294 1401 1300 1402
rect 1358 1406 1364 1407
rect 1358 1402 1359 1406
rect 1363 1402 1364 1406
rect 1358 1401 1364 1402
rect 1311 1399 1317 1400
rect 1311 1398 1312 1399
rect 1280 1396 1312 1398
rect 1247 1394 1253 1395
rect 1311 1395 1312 1396
rect 1316 1395 1317 1399
rect 1311 1394 1317 1395
rect 1375 1399 1381 1400
rect 1375 1395 1376 1399
rect 1380 1398 1381 1399
rect 1404 1398 1406 1412
rect 1431 1411 1432 1415
rect 1436 1414 1437 1415
rect 1479 1415 1485 1416
rect 1436 1412 1458 1414
rect 1436 1411 1437 1412
rect 1431 1410 1437 1411
rect 1414 1406 1420 1407
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1431 1399 1437 1400
rect 1431 1398 1432 1399
rect 1380 1396 1402 1398
rect 1404 1396 1432 1398
rect 1380 1395 1381 1396
rect 1375 1394 1381 1395
rect 770 1391 776 1392
rect 770 1390 771 1391
rect 560 1388 771 1390
rect 230 1387 236 1388
rect 230 1386 231 1387
rect 153 1384 231 1386
rect 153 1380 155 1384
rect 230 1383 231 1384
rect 235 1383 236 1387
rect 770 1387 771 1388
rect 775 1387 776 1391
rect 985 1390 987 1394
rect 1254 1391 1260 1392
rect 1254 1390 1255 1391
rect 985 1388 1255 1390
rect 770 1386 776 1387
rect 1254 1387 1255 1388
rect 1259 1387 1260 1391
rect 1400 1390 1402 1396
rect 1431 1395 1432 1396
rect 1436 1395 1437 1399
rect 1456 1398 1458 1412
rect 1479 1411 1480 1415
rect 1484 1414 1485 1415
rect 1487 1415 1493 1416
rect 1487 1414 1488 1415
rect 1484 1412 1488 1414
rect 1484 1411 1485 1412
rect 1479 1410 1485 1411
rect 1487 1411 1488 1412
rect 1492 1411 1493 1415
rect 1487 1410 1493 1411
rect 1495 1415 1501 1416
rect 1495 1411 1496 1415
rect 1500 1414 1501 1415
rect 1519 1415 1525 1416
rect 1519 1414 1520 1415
rect 1500 1412 1520 1414
rect 1500 1411 1501 1412
rect 1495 1410 1501 1411
rect 1519 1411 1520 1412
rect 1524 1411 1525 1415
rect 1519 1410 1525 1411
rect 1567 1415 1576 1416
rect 1567 1411 1568 1415
rect 1575 1411 1576 1415
rect 1607 1415 1613 1416
rect 1607 1414 1608 1415
rect 1567 1410 1576 1411
rect 1584 1412 1608 1414
rect 1462 1406 1468 1407
rect 1462 1402 1463 1406
rect 1467 1402 1468 1406
rect 1462 1401 1468 1402
rect 1502 1406 1508 1407
rect 1502 1402 1503 1406
rect 1507 1402 1508 1406
rect 1502 1401 1508 1402
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1479 1399 1485 1400
rect 1479 1398 1480 1399
rect 1456 1396 1480 1398
rect 1431 1394 1437 1395
rect 1479 1395 1480 1396
rect 1484 1395 1485 1399
rect 1479 1394 1485 1395
rect 1519 1399 1528 1400
rect 1519 1395 1520 1399
rect 1527 1395 1528 1399
rect 1519 1394 1528 1395
rect 1567 1399 1573 1400
rect 1567 1395 1568 1399
rect 1572 1398 1573 1399
rect 1584 1398 1586 1412
rect 1607 1411 1608 1412
rect 1612 1411 1613 1415
rect 1607 1410 1613 1411
rect 1639 1415 1645 1416
rect 1639 1411 1640 1415
rect 1644 1414 1645 1415
rect 1647 1415 1653 1416
rect 1647 1414 1648 1415
rect 1644 1412 1648 1414
rect 1644 1411 1645 1412
rect 1639 1410 1645 1411
rect 1647 1411 1648 1412
rect 1652 1411 1653 1415
rect 1647 1410 1653 1411
rect 1590 1406 1596 1407
rect 1590 1402 1591 1406
rect 1595 1402 1596 1406
rect 1590 1401 1596 1402
rect 1622 1406 1628 1407
rect 1622 1402 1623 1406
rect 1627 1402 1628 1406
rect 1622 1401 1628 1402
rect 1662 1404 1668 1405
rect 1662 1400 1663 1404
rect 1667 1400 1668 1404
rect 1572 1396 1586 1398
rect 1607 1399 1613 1400
rect 1572 1395 1573 1396
rect 1567 1394 1573 1395
rect 1607 1395 1608 1399
rect 1612 1398 1613 1399
rect 1630 1399 1636 1400
rect 1630 1398 1631 1399
rect 1612 1396 1631 1398
rect 1612 1395 1613 1396
rect 1607 1394 1613 1395
rect 1630 1395 1631 1396
rect 1635 1395 1636 1399
rect 1630 1394 1636 1395
rect 1638 1399 1645 1400
rect 1662 1399 1668 1400
rect 1638 1395 1639 1399
rect 1644 1395 1645 1399
rect 1638 1394 1645 1395
rect 1495 1391 1501 1392
rect 1495 1390 1496 1391
rect 1400 1388 1496 1390
rect 1254 1386 1260 1387
rect 1495 1387 1496 1388
rect 1500 1387 1501 1391
rect 1495 1386 1501 1387
rect 230 1382 236 1383
rect 527 1383 533 1384
rect 160 1380 187 1382
rect 241 1380 298 1382
rect 319 1380 371 1382
rect 151 1379 157 1380
rect 110 1376 116 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 151 1375 152 1379
rect 156 1375 157 1379
rect 110 1371 116 1372
rect 134 1374 140 1375
rect 151 1374 157 1375
rect 134 1370 135 1374
rect 139 1370 140 1374
rect 134 1369 140 1370
rect 151 1363 157 1364
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 151 1359 152 1363
rect 156 1362 157 1363
rect 160 1362 162 1380
rect 183 1379 189 1380
rect 183 1375 184 1379
rect 188 1375 189 1379
rect 239 1379 245 1380
rect 239 1375 240 1379
rect 244 1375 245 1379
rect 166 1374 172 1375
rect 183 1374 189 1375
rect 222 1374 228 1375
rect 239 1374 245 1375
rect 286 1374 292 1375
rect 166 1370 167 1374
rect 171 1370 172 1374
rect 166 1369 172 1370
rect 222 1370 223 1374
rect 227 1370 228 1374
rect 222 1369 228 1370
rect 286 1370 287 1374
rect 291 1370 292 1374
rect 286 1369 292 1370
rect 156 1360 162 1362
rect 183 1363 189 1364
rect 156 1359 157 1360
rect 151 1358 157 1359
rect 183 1359 184 1363
rect 188 1362 189 1363
rect 198 1363 204 1364
rect 198 1362 199 1363
rect 188 1360 199 1362
rect 188 1359 189 1360
rect 183 1358 189 1359
rect 198 1359 199 1360
rect 203 1359 204 1363
rect 198 1358 204 1359
rect 239 1363 248 1364
rect 239 1359 240 1363
rect 247 1359 248 1363
rect 296 1362 298 1380
rect 303 1379 309 1380
rect 303 1375 304 1379
rect 308 1378 309 1379
rect 319 1378 321 1380
rect 308 1376 321 1378
rect 308 1375 309 1376
rect 303 1374 309 1375
rect 358 1374 364 1375
rect 358 1370 359 1374
rect 363 1370 364 1374
rect 358 1369 364 1370
rect 303 1363 309 1364
rect 303 1362 304 1363
rect 296 1360 304 1362
rect 239 1358 248 1359
rect 303 1359 304 1360
rect 308 1359 309 1363
rect 369 1362 371 1380
rect 375 1379 381 1380
rect 375 1375 376 1379
rect 380 1378 381 1379
rect 438 1379 444 1380
rect 380 1376 418 1378
rect 380 1375 381 1376
rect 375 1374 381 1375
rect 416 1366 418 1376
rect 438 1375 439 1379
rect 443 1378 444 1379
rect 447 1379 453 1380
rect 447 1378 448 1379
rect 443 1376 448 1378
rect 443 1375 444 1376
rect 430 1374 436 1375
rect 438 1374 444 1375
rect 447 1375 448 1376
rect 452 1375 453 1379
rect 518 1379 525 1380
rect 518 1375 519 1379
rect 524 1375 525 1379
rect 527 1379 528 1383
rect 532 1382 533 1383
rect 607 1383 613 1384
rect 532 1380 594 1382
rect 532 1379 533 1380
rect 527 1378 533 1379
rect 592 1378 594 1380
rect 599 1379 605 1380
rect 599 1378 600 1379
rect 592 1376 600 1378
rect 599 1375 600 1376
rect 604 1375 605 1379
rect 607 1379 608 1383
rect 612 1382 613 1383
rect 767 1383 773 1384
rect 612 1380 683 1382
rect 612 1379 613 1380
rect 607 1378 613 1379
rect 679 1379 685 1380
rect 679 1375 680 1379
rect 684 1375 685 1379
rect 750 1379 756 1380
rect 750 1375 751 1379
rect 755 1378 756 1379
rect 759 1379 765 1380
rect 759 1378 760 1379
rect 755 1376 760 1378
rect 755 1375 756 1376
rect 447 1374 453 1375
rect 502 1374 508 1375
rect 518 1374 525 1375
rect 582 1374 588 1375
rect 599 1374 605 1375
rect 662 1374 668 1375
rect 679 1374 685 1375
rect 742 1374 748 1375
rect 750 1374 756 1375
rect 759 1375 760 1376
rect 764 1375 765 1379
rect 767 1379 768 1383
rect 772 1382 773 1383
rect 911 1383 917 1384
rect 772 1380 826 1382
rect 772 1379 773 1380
rect 767 1378 773 1379
rect 824 1378 826 1380
rect 831 1379 837 1380
rect 831 1378 832 1379
rect 824 1376 832 1378
rect 831 1375 832 1376
rect 836 1375 837 1379
rect 902 1379 909 1380
rect 902 1375 903 1379
rect 908 1375 909 1379
rect 911 1379 912 1383
rect 916 1382 917 1383
rect 983 1383 989 1384
rect 916 1380 970 1382
rect 916 1379 917 1380
rect 911 1378 917 1379
rect 968 1378 970 1380
rect 975 1379 981 1380
rect 975 1378 976 1379
rect 968 1376 976 1378
rect 975 1375 976 1376
rect 980 1375 981 1379
rect 983 1379 984 1383
rect 988 1382 989 1383
rect 1055 1383 1061 1384
rect 988 1380 1051 1382
rect 988 1379 989 1380
rect 983 1378 989 1379
rect 1047 1379 1053 1380
rect 1047 1375 1048 1379
rect 1052 1375 1053 1379
rect 1055 1379 1056 1383
rect 1060 1382 1061 1383
rect 1127 1383 1133 1384
rect 1060 1380 1114 1382
rect 1060 1379 1061 1380
rect 1055 1378 1061 1379
rect 1112 1378 1114 1380
rect 1119 1379 1125 1380
rect 1119 1378 1120 1379
rect 1112 1376 1120 1378
rect 1119 1375 1120 1376
rect 1124 1375 1125 1379
rect 1127 1379 1128 1383
rect 1132 1382 1133 1383
rect 1199 1383 1205 1384
rect 1132 1380 1186 1382
rect 1132 1379 1133 1380
rect 1127 1378 1133 1379
rect 1184 1378 1186 1380
rect 1191 1379 1197 1380
rect 1191 1378 1192 1379
rect 1184 1376 1192 1378
rect 1191 1375 1192 1376
rect 1196 1375 1197 1379
rect 1199 1379 1200 1383
rect 1204 1382 1205 1383
rect 1327 1383 1333 1384
rect 1204 1380 1250 1382
rect 1204 1379 1205 1380
rect 1199 1378 1205 1379
rect 1248 1378 1250 1380
rect 1255 1379 1261 1380
rect 1255 1378 1256 1379
rect 1248 1376 1256 1378
rect 1255 1375 1256 1376
rect 1260 1375 1261 1379
rect 1318 1379 1325 1380
rect 1318 1375 1319 1379
rect 1324 1375 1325 1379
rect 1327 1379 1328 1383
rect 1332 1382 1333 1383
rect 1391 1383 1397 1384
rect 1332 1380 1378 1382
rect 1332 1379 1333 1380
rect 1327 1378 1333 1379
rect 1376 1378 1378 1380
rect 1383 1379 1389 1380
rect 1383 1378 1384 1379
rect 1376 1376 1384 1378
rect 1383 1375 1384 1376
rect 1388 1375 1389 1379
rect 1391 1379 1392 1383
rect 1396 1382 1397 1383
rect 1487 1383 1493 1384
rect 1396 1380 1442 1382
rect 1396 1379 1397 1380
rect 1391 1378 1397 1379
rect 1440 1378 1442 1380
rect 1447 1379 1453 1380
rect 1447 1378 1448 1379
rect 1440 1376 1448 1378
rect 1447 1375 1448 1376
rect 1452 1375 1453 1379
rect 1487 1379 1488 1383
rect 1492 1382 1493 1383
rect 1519 1383 1525 1384
rect 1492 1380 1506 1382
rect 1492 1379 1493 1380
rect 1487 1378 1493 1379
rect 1504 1378 1506 1380
rect 1511 1379 1517 1380
rect 1511 1378 1512 1379
rect 1504 1376 1512 1378
rect 1511 1375 1512 1376
rect 1516 1375 1517 1379
rect 1519 1379 1520 1383
rect 1524 1382 1525 1383
rect 1524 1380 1578 1382
rect 1524 1379 1525 1380
rect 1519 1378 1525 1379
rect 1576 1378 1578 1380
rect 1583 1379 1589 1380
rect 1583 1378 1584 1379
rect 1576 1376 1584 1378
rect 1583 1375 1584 1376
rect 1588 1375 1589 1379
rect 1639 1379 1648 1380
rect 1639 1375 1640 1379
rect 1647 1375 1648 1379
rect 759 1374 765 1375
rect 814 1374 820 1375
rect 831 1374 837 1375
rect 886 1374 892 1375
rect 902 1374 909 1375
rect 958 1374 964 1375
rect 975 1374 981 1375
rect 1030 1374 1036 1375
rect 1047 1374 1053 1375
rect 1102 1374 1108 1375
rect 1119 1374 1125 1375
rect 1174 1374 1180 1375
rect 1191 1374 1197 1375
rect 1238 1374 1244 1375
rect 1255 1374 1261 1375
rect 1302 1374 1308 1375
rect 1318 1374 1325 1375
rect 1366 1374 1372 1375
rect 1383 1374 1389 1375
rect 1430 1374 1436 1375
rect 1447 1374 1453 1375
rect 1494 1374 1500 1375
rect 1511 1374 1517 1375
rect 1566 1374 1572 1375
rect 1583 1374 1589 1375
rect 1622 1374 1628 1375
rect 1639 1374 1648 1375
rect 1662 1376 1668 1377
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 502 1370 503 1374
rect 507 1370 508 1374
rect 502 1369 508 1370
rect 582 1370 583 1374
rect 587 1370 588 1374
rect 582 1369 588 1370
rect 662 1370 663 1374
rect 667 1370 668 1374
rect 662 1369 668 1370
rect 742 1370 743 1374
rect 747 1370 748 1374
rect 742 1369 748 1370
rect 814 1370 815 1374
rect 819 1370 820 1374
rect 814 1369 820 1370
rect 886 1370 887 1374
rect 891 1370 892 1374
rect 886 1369 892 1370
rect 958 1370 959 1374
rect 963 1370 964 1374
rect 958 1369 964 1370
rect 1030 1370 1031 1374
rect 1035 1370 1036 1374
rect 1030 1369 1036 1370
rect 1102 1370 1103 1374
rect 1107 1370 1108 1374
rect 1102 1369 1108 1370
rect 1174 1370 1175 1374
rect 1179 1370 1180 1374
rect 1174 1369 1180 1370
rect 1238 1370 1239 1374
rect 1243 1370 1244 1374
rect 1238 1369 1244 1370
rect 1302 1370 1303 1374
rect 1307 1370 1308 1374
rect 1302 1369 1308 1370
rect 1366 1370 1367 1374
rect 1371 1370 1372 1374
rect 1366 1369 1372 1370
rect 1430 1370 1431 1374
rect 1435 1370 1436 1374
rect 1430 1369 1436 1370
rect 1494 1370 1495 1374
rect 1499 1370 1500 1374
rect 1494 1369 1500 1370
rect 1566 1370 1567 1374
rect 1571 1370 1572 1374
rect 1566 1369 1572 1370
rect 1622 1370 1623 1374
rect 1627 1370 1628 1374
rect 1662 1372 1663 1376
rect 1667 1372 1668 1376
rect 1662 1371 1668 1372
rect 1622 1369 1628 1370
rect 416 1364 430 1366
rect 375 1363 381 1364
rect 375 1362 376 1363
rect 369 1360 376 1362
rect 303 1358 309 1359
rect 375 1359 376 1360
rect 380 1359 381 1363
rect 428 1362 442 1364
rect 447 1363 453 1364
rect 447 1362 448 1363
rect 440 1360 448 1362
rect 375 1358 381 1359
rect 447 1359 448 1360
rect 452 1359 453 1363
rect 447 1358 453 1359
rect 519 1363 525 1364
rect 519 1359 520 1363
rect 524 1362 525 1363
rect 527 1363 533 1364
rect 527 1362 528 1363
rect 524 1360 528 1362
rect 524 1359 525 1360
rect 519 1358 525 1359
rect 527 1359 528 1360
rect 532 1359 533 1363
rect 527 1358 533 1359
rect 599 1363 605 1364
rect 599 1359 600 1363
rect 604 1362 605 1363
rect 607 1363 613 1364
rect 607 1362 608 1363
rect 604 1360 608 1362
rect 604 1359 605 1360
rect 599 1358 605 1359
rect 607 1359 608 1360
rect 612 1359 613 1363
rect 607 1358 613 1359
rect 679 1363 685 1364
rect 679 1359 680 1363
rect 684 1362 685 1363
rect 710 1363 716 1364
rect 710 1362 711 1363
rect 684 1360 711 1362
rect 684 1359 685 1360
rect 679 1358 685 1359
rect 710 1359 711 1360
rect 715 1359 716 1363
rect 710 1358 716 1359
rect 759 1363 765 1364
rect 759 1359 760 1363
rect 764 1362 765 1363
rect 767 1363 773 1364
rect 767 1362 768 1363
rect 764 1360 768 1362
rect 764 1359 765 1360
rect 759 1358 765 1359
rect 767 1359 768 1360
rect 772 1359 773 1363
rect 831 1363 837 1364
rect 831 1362 832 1363
rect 767 1358 773 1359
rect 824 1360 832 1362
rect 110 1354 116 1355
rect 134 1357 140 1358
rect 134 1353 135 1357
rect 139 1353 140 1357
rect 134 1352 140 1353
rect 166 1357 172 1358
rect 166 1353 167 1357
rect 171 1353 172 1357
rect 166 1352 172 1353
rect 222 1357 228 1358
rect 222 1353 223 1357
rect 227 1353 228 1357
rect 222 1352 228 1353
rect 286 1357 292 1358
rect 286 1353 287 1357
rect 291 1353 292 1357
rect 286 1352 292 1353
rect 358 1357 364 1358
rect 358 1353 359 1357
rect 363 1353 364 1357
rect 358 1352 364 1353
rect 430 1357 436 1358
rect 430 1353 431 1357
rect 435 1353 436 1357
rect 430 1352 436 1353
rect 502 1357 508 1358
rect 502 1353 503 1357
rect 507 1353 508 1357
rect 502 1352 508 1353
rect 582 1357 588 1358
rect 582 1353 583 1357
rect 587 1353 588 1357
rect 582 1352 588 1353
rect 662 1357 668 1358
rect 662 1353 663 1357
rect 667 1353 668 1357
rect 662 1352 668 1353
rect 742 1357 748 1358
rect 742 1353 743 1357
rect 747 1353 748 1357
rect 742 1352 748 1353
rect 814 1357 820 1358
rect 814 1353 815 1357
rect 819 1353 820 1357
rect 814 1352 820 1353
rect 518 1351 524 1352
rect 518 1347 519 1351
rect 523 1350 524 1351
rect 824 1350 826 1360
rect 831 1359 832 1360
rect 836 1359 837 1363
rect 831 1358 837 1359
rect 903 1363 909 1364
rect 903 1359 904 1363
rect 908 1362 909 1363
rect 911 1363 917 1364
rect 911 1362 912 1363
rect 908 1360 912 1362
rect 908 1359 909 1360
rect 903 1358 909 1359
rect 911 1359 912 1360
rect 916 1359 917 1363
rect 911 1358 917 1359
rect 975 1363 981 1364
rect 975 1359 976 1363
rect 980 1362 981 1363
rect 983 1363 989 1364
rect 983 1362 984 1363
rect 980 1360 984 1362
rect 980 1359 981 1360
rect 975 1358 981 1359
rect 983 1359 984 1360
rect 988 1359 989 1363
rect 983 1358 989 1359
rect 1047 1363 1053 1364
rect 1047 1359 1048 1363
rect 1052 1362 1053 1363
rect 1055 1363 1061 1364
rect 1055 1362 1056 1363
rect 1052 1360 1056 1362
rect 1052 1359 1053 1360
rect 1047 1358 1053 1359
rect 1055 1359 1056 1360
rect 1060 1359 1061 1363
rect 1055 1358 1061 1359
rect 1119 1363 1125 1364
rect 1119 1359 1120 1363
rect 1124 1362 1125 1363
rect 1127 1363 1133 1364
rect 1127 1362 1128 1363
rect 1124 1360 1128 1362
rect 1124 1359 1125 1360
rect 1119 1358 1125 1359
rect 1127 1359 1128 1360
rect 1132 1359 1133 1363
rect 1127 1358 1133 1359
rect 1191 1363 1197 1364
rect 1191 1359 1192 1363
rect 1196 1362 1197 1363
rect 1199 1363 1205 1364
rect 1199 1362 1200 1363
rect 1196 1360 1200 1362
rect 1196 1359 1197 1360
rect 1191 1358 1197 1359
rect 1199 1359 1200 1360
rect 1204 1359 1205 1363
rect 1199 1358 1205 1359
rect 1254 1363 1261 1364
rect 1254 1359 1255 1363
rect 1260 1359 1261 1363
rect 1254 1358 1261 1359
rect 1319 1363 1325 1364
rect 1319 1359 1320 1363
rect 1324 1362 1325 1363
rect 1327 1363 1333 1364
rect 1327 1362 1328 1363
rect 1324 1360 1328 1362
rect 1324 1359 1325 1360
rect 1319 1358 1325 1359
rect 1327 1359 1328 1360
rect 1332 1359 1333 1363
rect 1327 1358 1333 1359
rect 1383 1363 1389 1364
rect 1383 1359 1384 1363
rect 1388 1362 1389 1363
rect 1391 1363 1397 1364
rect 1391 1362 1392 1363
rect 1388 1360 1392 1362
rect 1388 1359 1389 1360
rect 1383 1358 1389 1359
rect 1391 1359 1392 1360
rect 1396 1359 1397 1363
rect 1391 1358 1397 1359
rect 1447 1363 1453 1364
rect 1447 1359 1448 1363
rect 1452 1362 1453 1363
rect 1486 1363 1492 1364
rect 1486 1362 1487 1363
rect 1452 1360 1487 1362
rect 1452 1359 1453 1360
rect 1447 1358 1453 1359
rect 1486 1359 1487 1360
rect 1491 1359 1492 1363
rect 1486 1358 1492 1359
rect 1511 1363 1517 1364
rect 1511 1359 1512 1363
rect 1516 1362 1517 1363
rect 1519 1363 1525 1364
rect 1519 1362 1520 1363
rect 1516 1360 1520 1362
rect 1516 1359 1517 1360
rect 1511 1358 1517 1359
rect 1519 1359 1520 1360
rect 1524 1359 1525 1363
rect 1583 1363 1589 1364
rect 1583 1362 1584 1363
rect 1519 1358 1525 1359
rect 1576 1360 1584 1362
rect 886 1357 892 1358
rect 886 1353 887 1357
rect 891 1353 892 1357
rect 886 1352 892 1353
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1030 1357 1036 1358
rect 1030 1353 1031 1357
rect 1035 1353 1036 1357
rect 1030 1352 1036 1353
rect 1102 1357 1108 1358
rect 1102 1353 1103 1357
rect 1107 1353 1108 1357
rect 1102 1352 1108 1353
rect 1174 1357 1180 1358
rect 1174 1353 1175 1357
rect 1179 1353 1180 1357
rect 1174 1352 1180 1353
rect 1238 1357 1244 1358
rect 1238 1353 1239 1357
rect 1243 1353 1244 1357
rect 1238 1352 1244 1353
rect 1302 1357 1308 1358
rect 1302 1353 1303 1357
rect 1307 1353 1308 1357
rect 1302 1352 1308 1353
rect 1366 1357 1372 1358
rect 1366 1353 1367 1357
rect 1371 1353 1372 1357
rect 1366 1352 1372 1353
rect 1430 1357 1436 1358
rect 1430 1353 1431 1357
rect 1435 1353 1436 1357
rect 1430 1352 1436 1353
rect 1494 1357 1500 1358
rect 1494 1353 1495 1357
rect 1499 1353 1500 1357
rect 1494 1352 1500 1353
rect 1566 1357 1572 1358
rect 1566 1353 1567 1357
rect 1571 1353 1572 1357
rect 1566 1352 1572 1353
rect 523 1348 826 1350
rect 902 1351 908 1352
rect 523 1347 524 1348
rect 518 1346 524 1347
rect 902 1347 903 1351
rect 907 1350 908 1351
rect 1318 1351 1324 1352
rect 907 1348 1161 1350
rect 907 1347 908 1348
rect 902 1346 908 1347
rect 134 1343 140 1344
rect 110 1341 116 1342
rect 110 1337 111 1341
rect 115 1337 116 1341
rect 134 1339 135 1343
rect 139 1339 140 1343
rect 134 1338 140 1339
rect 182 1343 188 1344
rect 182 1339 183 1343
rect 187 1339 188 1343
rect 182 1338 188 1339
rect 238 1343 244 1344
rect 238 1339 239 1343
rect 243 1339 244 1343
rect 238 1338 244 1339
rect 294 1343 300 1344
rect 294 1339 295 1343
rect 299 1339 300 1343
rect 294 1338 300 1339
rect 350 1343 356 1344
rect 350 1339 351 1343
rect 355 1339 356 1343
rect 350 1338 356 1339
rect 398 1343 404 1344
rect 398 1339 399 1343
rect 403 1339 404 1343
rect 398 1338 404 1339
rect 454 1343 460 1344
rect 454 1339 455 1343
rect 459 1339 460 1343
rect 454 1338 460 1339
rect 510 1343 516 1344
rect 510 1339 511 1343
rect 515 1339 516 1343
rect 510 1338 516 1339
rect 566 1343 572 1344
rect 566 1339 567 1343
rect 571 1339 572 1343
rect 566 1338 572 1339
rect 630 1343 636 1344
rect 630 1339 631 1343
rect 635 1339 636 1343
rect 630 1338 636 1339
rect 694 1343 700 1344
rect 694 1339 695 1343
rect 699 1339 700 1343
rect 694 1338 700 1339
rect 758 1343 764 1344
rect 758 1339 759 1343
rect 763 1339 764 1343
rect 758 1338 764 1339
rect 822 1343 828 1344
rect 822 1339 823 1343
rect 827 1339 828 1343
rect 822 1338 828 1339
rect 886 1343 892 1344
rect 886 1339 887 1343
rect 891 1339 892 1343
rect 886 1338 892 1339
rect 958 1343 964 1344
rect 958 1339 959 1343
rect 963 1339 964 1343
rect 958 1338 964 1339
rect 1022 1343 1028 1344
rect 1022 1339 1023 1343
rect 1027 1339 1028 1343
rect 1022 1338 1028 1339
rect 1086 1343 1092 1344
rect 1086 1339 1087 1343
rect 1091 1339 1092 1343
rect 1086 1338 1092 1339
rect 1150 1343 1156 1344
rect 1150 1339 1151 1343
rect 1155 1339 1156 1343
rect 1150 1338 1156 1339
rect 110 1336 116 1337
rect 150 1335 157 1336
rect 150 1331 151 1335
rect 156 1331 157 1335
rect 199 1335 205 1336
rect 199 1334 200 1335
rect 150 1330 157 1331
rect 176 1332 200 1334
rect 134 1326 140 1327
rect 110 1324 116 1325
rect 110 1320 111 1324
rect 115 1320 116 1324
rect 134 1322 135 1326
rect 139 1322 140 1326
rect 134 1321 140 1322
rect 110 1319 116 1320
rect 151 1319 157 1320
rect 151 1315 152 1319
rect 156 1318 157 1319
rect 176 1318 178 1332
rect 199 1331 200 1332
rect 204 1331 205 1335
rect 199 1330 205 1331
rect 255 1335 261 1336
rect 255 1331 256 1335
rect 260 1334 261 1335
rect 311 1335 317 1336
rect 260 1332 306 1334
rect 260 1331 261 1332
rect 255 1330 261 1331
rect 182 1326 188 1327
rect 182 1322 183 1326
rect 187 1322 188 1326
rect 182 1321 188 1322
rect 238 1326 244 1327
rect 238 1322 239 1326
rect 243 1322 244 1326
rect 238 1321 244 1322
rect 294 1326 300 1327
rect 294 1322 295 1326
rect 299 1322 300 1326
rect 294 1321 300 1322
rect 156 1316 178 1318
rect 198 1319 205 1320
rect 156 1315 157 1316
rect 151 1314 157 1315
rect 198 1315 199 1319
rect 204 1315 205 1319
rect 198 1314 205 1315
rect 255 1319 261 1320
rect 255 1315 256 1319
rect 260 1318 261 1319
rect 304 1318 306 1332
rect 311 1331 312 1335
rect 316 1334 317 1335
rect 367 1335 373 1336
rect 316 1332 321 1334
rect 316 1331 317 1332
rect 311 1330 317 1331
rect 311 1319 317 1320
rect 311 1318 312 1319
rect 260 1316 290 1318
rect 304 1316 312 1318
rect 260 1315 261 1316
rect 255 1314 261 1315
rect 288 1310 290 1316
rect 311 1315 312 1316
rect 316 1315 317 1319
rect 319 1318 321 1332
rect 367 1331 368 1335
rect 372 1334 373 1335
rect 415 1335 421 1336
rect 372 1332 410 1334
rect 372 1331 373 1332
rect 367 1330 373 1331
rect 350 1326 356 1327
rect 350 1322 351 1326
rect 355 1322 356 1326
rect 350 1321 356 1322
rect 398 1326 404 1327
rect 398 1322 399 1326
rect 403 1322 404 1326
rect 398 1321 404 1322
rect 367 1319 373 1320
rect 367 1318 368 1319
rect 319 1316 368 1318
rect 311 1314 317 1315
rect 367 1315 368 1316
rect 372 1315 373 1319
rect 408 1318 410 1332
rect 415 1331 416 1335
rect 420 1334 421 1335
rect 438 1335 444 1336
rect 438 1334 439 1335
rect 420 1332 439 1334
rect 420 1331 421 1332
rect 415 1330 421 1331
rect 438 1331 439 1332
rect 443 1331 444 1335
rect 438 1330 444 1331
rect 471 1335 477 1336
rect 471 1331 472 1335
rect 476 1334 477 1335
rect 527 1335 533 1336
rect 476 1332 502 1334
rect 476 1331 477 1332
rect 471 1330 477 1331
rect 454 1326 460 1327
rect 454 1322 455 1326
rect 459 1322 460 1326
rect 454 1321 460 1322
rect 415 1319 421 1320
rect 415 1318 416 1319
rect 408 1316 416 1318
rect 367 1314 373 1315
rect 415 1315 416 1316
rect 420 1315 421 1319
rect 415 1314 421 1315
rect 471 1319 477 1320
rect 471 1315 472 1319
rect 476 1318 477 1319
rect 500 1318 502 1332
rect 527 1331 528 1335
rect 532 1334 533 1335
rect 583 1335 589 1336
rect 532 1332 558 1334
rect 532 1331 533 1332
rect 527 1330 533 1331
rect 510 1326 516 1327
rect 510 1322 511 1326
rect 515 1322 516 1326
rect 510 1321 516 1322
rect 527 1319 533 1320
rect 527 1318 528 1319
rect 476 1316 498 1318
rect 500 1316 528 1318
rect 476 1315 477 1316
rect 471 1314 477 1315
rect 390 1311 396 1312
rect 390 1310 391 1311
rect 288 1308 391 1310
rect 390 1307 391 1308
rect 395 1307 396 1311
rect 496 1310 498 1316
rect 527 1315 528 1316
rect 532 1315 533 1319
rect 556 1318 558 1332
rect 583 1331 584 1335
rect 588 1334 589 1335
rect 622 1335 628 1336
rect 622 1334 623 1335
rect 588 1332 623 1334
rect 588 1331 589 1332
rect 583 1330 589 1331
rect 622 1331 623 1332
rect 627 1331 628 1335
rect 622 1330 628 1331
rect 642 1335 653 1336
rect 642 1331 643 1335
rect 647 1331 648 1335
rect 652 1331 653 1335
rect 642 1330 653 1331
rect 711 1335 717 1336
rect 711 1331 712 1335
rect 716 1334 717 1335
rect 738 1335 744 1336
rect 738 1334 739 1335
rect 716 1332 739 1334
rect 716 1331 717 1332
rect 711 1330 717 1331
rect 738 1331 739 1332
rect 743 1331 744 1335
rect 775 1335 781 1336
rect 775 1334 776 1335
rect 738 1330 744 1331
rect 748 1332 776 1334
rect 566 1326 572 1327
rect 566 1322 567 1326
rect 571 1322 572 1326
rect 566 1321 572 1322
rect 630 1326 636 1327
rect 630 1322 631 1326
rect 635 1322 636 1326
rect 630 1321 636 1322
rect 694 1326 700 1327
rect 748 1326 750 1332
rect 775 1331 776 1332
rect 780 1331 781 1335
rect 775 1330 781 1331
rect 839 1335 845 1336
rect 839 1331 840 1335
rect 844 1334 845 1335
rect 903 1335 909 1336
rect 844 1332 874 1334
rect 844 1331 845 1332
rect 839 1330 845 1331
rect 694 1322 695 1326
rect 699 1322 700 1326
rect 694 1321 700 1322
rect 704 1324 750 1326
rect 758 1326 764 1327
rect 583 1319 589 1320
rect 583 1318 584 1319
rect 556 1316 584 1318
rect 527 1314 533 1315
rect 583 1315 584 1316
rect 588 1315 589 1319
rect 583 1314 589 1315
rect 647 1319 653 1320
rect 647 1315 648 1319
rect 652 1318 653 1319
rect 704 1318 706 1324
rect 758 1322 759 1326
rect 763 1322 764 1326
rect 758 1321 764 1322
rect 822 1326 828 1327
rect 822 1322 823 1326
rect 827 1322 828 1326
rect 822 1321 828 1322
rect 652 1316 706 1318
rect 710 1319 717 1320
rect 652 1315 653 1316
rect 647 1314 653 1315
rect 710 1315 711 1319
rect 716 1315 717 1319
rect 710 1314 717 1315
rect 738 1319 744 1320
rect 738 1315 739 1319
rect 743 1318 744 1319
rect 775 1319 781 1320
rect 775 1318 776 1319
rect 743 1316 776 1318
rect 743 1315 744 1316
rect 738 1314 744 1315
rect 775 1315 776 1316
rect 780 1315 781 1319
rect 775 1314 781 1315
rect 839 1319 845 1320
rect 839 1315 840 1319
rect 844 1318 845 1319
rect 872 1318 874 1332
rect 903 1331 904 1335
rect 908 1334 909 1335
rect 975 1335 981 1336
rect 908 1332 942 1334
rect 908 1331 909 1332
rect 903 1330 909 1331
rect 886 1326 892 1327
rect 886 1322 887 1326
rect 891 1322 892 1326
rect 886 1321 892 1322
rect 903 1319 909 1320
rect 903 1318 904 1319
rect 844 1316 870 1318
rect 872 1316 904 1318
rect 844 1315 845 1316
rect 839 1314 845 1315
rect 642 1311 648 1312
rect 642 1310 643 1311
rect 496 1308 643 1310
rect 390 1306 396 1307
rect 642 1307 643 1308
rect 647 1307 648 1311
rect 868 1310 870 1316
rect 903 1315 904 1316
rect 908 1315 909 1319
rect 940 1318 942 1332
rect 975 1331 976 1335
rect 980 1334 981 1335
rect 1039 1335 1045 1336
rect 980 1332 1010 1334
rect 980 1331 981 1332
rect 975 1330 981 1331
rect 958 1326 964 1327
rect 958 1322 959 1326
rect 963 1322 964 1326
rect 958 1321 964 1322
rect 975 1319 981 1320
rect 975 1318 976 1319
rect 940 1316 976 1318
rect 903 1314 909 1315
rect 975 1315 976 1316
rect 980 1315 981 1319
rect 1008 1318 1010 1332
rect 1039 1331 1040 1335
rect 1044 1334 1045 1335
rect 1103 1335 1109 1336
rect 1044 1332 1074 1334
rect 1044 1331 1045 1332
rect 1039 1330 1045 1331
rect 1022 1326 1028 1327
rect 1022 1322 1023 1326
rect 1027 1322 1028 1326
rect 1022 1321 1028 1322
rect 1039 1319 1045 1320
rect 1039 1318 1040 1319
rect 1008 1316 1040 1318
rect 975 1314 981 1315
rect 1039 1315 1040 1316
rect 1044 1315 1045 1319
rect 1072 1318 1074 1332
rect 1103 1331 1104 1335
rect 1108 1334 1109 1335
rect 1159 1334 1161 1348
rect 1318 1347 1319 1351
rect 1323 1350 1324 1351
rect 1576 1350 1578 1360
rect 1583 1359 1584 1360
rect 1588 1359 1589 1363
rect 1583 1358 1589 1359
rect 1634 1363 1645 1364
rect 1634 1359 1635 1363
rect 1639 1359 1640 1363
rect 1644 1359 1645 1363
rect 1634 1358 1645 1359
rect 1662 1359 1668 1360
rect 1622 1357 1628 1358
rect 1622 1353 1623 1357
rect 1627 1353 1628 1357
rect 1662 1355 1663 1359
rect 1667 1355 1668 1359
rect 1662 1354 1668 1355
rect 1622 1352 1628 1353
rect 1323 1348 1578 1350
rect 1323 1347 1324 1348
rect 1318 1346 1324 1347
rect 1214 1343 1220 1344
rect 1214 1339 1215 1343
rect 1219 1339 1220 1343
rect 1214 1338 1220 1339
rect 1278 1343 1284 1344
rect 1278 1339 1279 1343
rect 1283 1339 1284 1343
rect 1278 1338 1284 1339
rect 1342 1343 1348 1344
rect 1342 1339 1343 1343
rect 1347 1339 1348 1343
rect 1342 1338 1348 1339
rect 1406 1343 1412 1344
rect 1406 1339 1407 1343
rect 1411 1339 1412 1343
rect 1406 1338 1412 1339
rect 1478 1343 1484 1344
rect 1478 1339 1479 1343
rect 1483 1339 1484 1343
rect 1478 1338 1484 1339
rect 1558 1343 1564 1344
rect 1558 1339 1559 1343
rect 1563 1339 1564 1343
rect 1558 1338 1564 1339
rect 1622 1343 1628 1344
rect 1622 1339 1623 1343
rect 1627 1339 1628 1343
rect 1622 1338 1628 1339
rect 1662 1341 1668 1342
rect 1662 1337 1663 1341
rect 1667 1337 1668 1341
rect 1662 1336 1668 1337
rect 1167 1335 1173 1336
rect 1167 1334 1168 1335
rect 1108 1332 1134 1334
rect 1159 1332 1168 1334
rect 1108 1331 1109 1332
rect 1103 1330 1109 1331
rect 1086 1326 1092 1327
rect 1086 1322 1087 1326
rect 1091 1322 1092 1326
rect 1086 1321 1092 1322
rect 1103 1319 1109 1320
rect 1103 1318 1104 1319
rect 1072 1316 1104 1318
rect 1039 1314 1045 1315
rect 1103 1315 1104 1316
rect 1108 1315 1109 1319
rect 1132 1318 1134 1332
rect 1167 1331 1168 1332
rect 1172 1331 1173 1335
rect 1167 1330 1173 1331
rect 1231 1335 1237 1336
rect 1231 1331 1232 1335
rect 1236 1334 1237 1335
rect 1295 1335 1301 1336
rect 1236 1332 1290 1334
rect 1236 1331 1237 1332
rect 1231 1330 1237 1331
rect 1150 1326 1156 1327
rect 1150 1322 1151 1326
rect 1155 1322 1156 1326
rect 1150 1321 1156 1322
rect 1214 1326 1220 1327
rect 1214 1322 1215 1326
rect 1219 1322 1220 1326
rect 1214 1321 1220 1322
rect 1278 1326 1284 1327
rect 1278 1322 1279 1326
rect 1283 1322 1284 1326
rect 1278 1321 1284 1322
rect 1167 1319 1173 1320
rect 1167 1318 1168 1319
rect 1132 1316 1168 1318
rect 1103 1314 1109 1315
rect 1167 1315 1168 1316
rect 1172 1315 1173 1319
rect 1167 1314 1173 1315
rect 1231 1319 1237 1320
rect 1231 1315 1232 1319
rect 1236 1315 1237 1319
rect 1288 1318 1290 1332
rect 1295 1331 1296 1335
rect 1300 1334 1301 1335
rect 1359 1335 1365 1336
rect 1300 1332 1354 1334
rect 1300 1331 1301 1332
rect 1295 1330 1301 1331
rect 1342 1326 1348 1327
rect 1342 1322 1343 1326
rect 1347 1322 1348 1326
rect 1342 1321 1348 1322
rect 1295 1319 1301 1320
rect 1295 1318 1296 1319
rect 1288 1316 1296 1318
rect 1231 1314 1237 1315
rect 1295 1315 1296 1316
rect 1300 1315 1301 1319
rect 1352 1318 1354 1332
rect 1359 1331 1360 1335
rect 1364 1334 1365 1335
rect 1374 1335 1380 1336
rect 1374 1334 1375 1335
rect 1364 1332 1375 1334
rect 1364 1331 1365 1332
rect 1359 1330 1365 1331
rect 1374 1331 1375 1332
rect 1379 1331 1380 1335
rect 1374 1330 1380 1331
rect 1382 1335 1388 1336
rect 1382 1331 1383 1335
rect 1387 1334 1388 1335
rect 1423 1335 1429 1336
rect 1423 1334 1424 1335
rect 1387 1332 1424 1334
rect 1387 1331 1388 1332
rect 1382 1330 1388 1331
rect 1423 1331 1424 1332
rect 1428 1331 1429 1335
rect 1423 1330 1429 1331
rect 1495 1335 1501 1336
rect 1495 1331 1496 1335
rect 1500 1334 1501 1335
rect 1574 1335 1581 1336
rect 1500 1332 1570 1334
rect 1500 1331 1501 1332
rect 1495 1330 1501 1331
rect 1406 1326 1412 1327
rect 1406 1322 1407 1326
rect 1411 1322 1412 1326
rect 1406 1321 1412 1322
rect 1478 1326 1484 1327
rect 1478 1322 1479 1326
rect 1483 1322 1484 1326
rect 1478 1321 1484 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1359 1319 1365 1320
rect 1359 1318 1360 1319
rect 1352 1316 1360 1318
rect 1295 1314 1301 1315
rect 1359 1315 1360 1316
rect 1364 1315 1365 1319
rect 1359 1314 1365 1315
rect 1423 1319 1429 1320
rect 1423 1315 1424 1319
rect 1428 1315 1429 1319
rect 1423 1314 1429 1315
rect 1486 1319 1492 1320
rect 1486 1315 1487 1319
rect 1491 1318 1492 1319
rect 1495 1319 1501 1320
rect 1495 1318 1496 1319
rect 1491 1316 1496 1318
rect 1491 1315 1492 1316
rect 1486 1314 1492 1315
rect 1495 1315 1496 1316
rect 1500 1315 1501 1319
rect 1568 1318 1570 1332
rect 1574 1331 1575 1335
rect 1580 1331 1581 1335
rect 1574 1330 1581 1331
rect 1639 1335 1645 1336
rect 1639 1331 1640 1335
rect 1644 1334 1645 1335
rect 1650 1335 1656 1336
rect 1650 1334 1651 1335
rect 1644 1332 1651 1334
rect 1644 1331 1645 1332
rect 1639 1330 1645 1331
rect 1650 1331 1651 1332
rect 1655 1331 1656 1335
rect 1650 1330 1656 1331
rect 1622 1326 1628 1327
rect 1622 1322 1623 1326
rect 1627 1322 1628 1326
rect 1622 1321 1628 1322
rect 1662 1324 1668 1325
rect 1662 1320 1663 1324
rect 1667 1320 1668 1324
rect 1575 1319 1581 1320
rect 1575 1318 1576 1319
rect 1568 1316 1576 1318
rect 1495 1314 1501 1315
rect 1575 1315 1576 1316
rect 1580 1315 1581 1319
rect 1575 1314 1581 1315
rect 1639 1319 1645 1320
rect 1639 1315 1640 1319
rect 1644 1318 1645 1319
rect 1647 1319 1653 1320
rect 1662 1319 1668 1320
rect 1647 1318 1648 1319
rect 1644 1316 1648 1318
rect 1644 1315 1645 1316
rect 1639 1314 1645 1315
rect 1647 1315 1648 1316
rect 1652 1315 1653 1319
rect 1647 1314 1653 1315
rect 1094 1311 1100 1312
rect 1094 1310 1095 1311
rect 868 1308 1095 1310
rect 642 1306 648 1307
rect 1094 1307 1095 1308
rect 1099 1307 1100 1311
rect 1233 1310 1235 1314
rect 1382 1311 1388 1312
rect 1382 1310 1383 1311
rect 1233 1308 1383 1310
rect 1094 1306 1100 1307
rect 1382 1307 1383 1308
rect 1387 1307 1388 1311
rect 1425 1310 1427 1314
rect 1574 1311 1580 1312
rect 1574 1310 1575 1311
rect 1425 1308 1575 1310
rect 1382 1306 1388 1307
rect 1574 1307 1575 1308
rect 1579 1307 1580 1311
rect 1574 1306 1580 1307
rect 159 1299 165 1300
rect 150 1295 157 1296
rect 110 1292 116 1293
rect 110 1288 111 1292
rect 115 1288 116 1292
rect 150 1291 151 1295
rect 156 1291 157 1295
rect 159 1295 160 1299
rect 164 1298 165 1299
rect 207 1299 213 1300
rect 164 1296 203 1298
rect 164 1295 165 1296
rect 159 1294 165 1295
rect 199 1295 205 1296
rect 199 1291 200 1295
rect 204 1291 205 1295
rect 207 1295 208 1299
rect 212 1298 213 1299
rect 303 1299 309 1300
rect 212 1296 242 1298
rect 212 1295 213 1296
rect 207 1294 213 1295
rect 240 1294 242 1296
rect 247 1295 253 1296
rect 247 1294 248 1295
rect 240 1292 248 1294
rect 247 1291 248 1292
rect 252 1291 253 1295
rect 294 1295 301 1296
rect 294 1291 295 1295
rect 300 1291 301 1295
rect 303 1295 304 1299
rect 308 1298 309 1299
rect 351 1299 357 1300
rect 308 1296 338 1298
rect 308 1295 309 1296
rect 303 1294 309 1295
rect 336 1294 338 1296
rect 343 1295 349 1296
rect 343 1294 344 1295
rect 336 1292 344 1294
rect 343 1291 344 1292
rect 348 1291 349 1295
rect 351 1295 352 1299
rect 356 1298 357 1299
rect 631 1299 637 1300
rect 356 1296 386 1298
rect 536 1296 554 1298
rect 356 1295 357 1296
rect 351 1294 357 1295
rect 384 1294 386 1296
rect 391 1295 397 1296
rect 391 1294 392 1295
rect 384 1292 392 1294
rect 391 1291 392 1292
rect 396 1291 397 1295
rect 447 1295 453 1296
rect 447 1291 448 1295
rect 452 1294 453 1295
rect 503 1295 509 1296
rect 452 1292 482 1294
rect 452 1291 453 1292
rect 110 1287 116 1288
rect 134 1290 140 1291
rect 150 1290 157 1291
rect 182 1290 188 1291
rect 199 1290 205 1291
rect 230 1290 236 1291
rect 247 1290 253 1291
rect 278 1290 284 1291
rect 294 1290 301 1291
rect 326 1290 332 1291
rect 343 1290 349 1291
rect 374 1290 380 1291
rect 391 1290 397 1291
rect 430 1290 436 1291
rect 447 1290 453 1291
rect 134 1286 135 1290
rect 139 1286 140 1290
rect 134 1285 140 1286
rect 182 1286 183 1290
rect 187 1286 188 1290
rect 182 1285 188 1286
rect 230 1286 231 1290
rect 235 1286 236 1290
rect 230 1285 236 1286
rect 278 1286 279 1290
rect 283 1286 284 1290
rect 278 1285 284 1286
rect 326 1286 327 1290
rect 331 1286 332 1290
rect 326 1285 332 1286
rect 374 1286 375 1290
rect 379 1286 380 1290
rect 374 1285 380 1286
rect 430 1286 431 1290
rect 435 1286 436 1290
rect 430 1285 436 1286
rect 480 1282 482 1292
rect 503 1291 504 1295
rect 508 1294 509 1295
rect 536 1294 538 1296
rect 508 1292 538 1294
rect 508 1291 509 1292
rect 486 1290 492 1291
rect 503 1290 509 1291
rect 542 1290 548 1291
rect 486 1286 487 1290
rect 491 1286 492 1290
rect 486 1285 492 1286
rect 542 1286 543 1290
rect 547 1286 548 1290
rect 542 1285 548 1286
rect 480 1280 486 1282
rect 151 1279 157 1280
rect 110 1275 116 1276
rect 110 1271 111 1275
rect 115 1271 116 1275
rect 151 1275 152 1279
rect 156 1278 157 1279
rect 159 1279 165 1280
rect 159 1278 160 1279
rect 156 1276 160 1278
rect 156 1275 157 1276
rect 151 1274 157 1275
rect 159 1275 160 1276
rect 164 1275 165 1279
rect 159 1274 165 1275
rect 199 1279 205 1280
rect 199 1275 200 1279
rect 204 1278 205 1279
rect 207 1279 213 1280
rect 207 1278 208 1279
rect 204 1276 208 1278
rect 204 1275 205 1276
rect 199 1274 205 1275
rect 207 1275 208 1276
rect 212 1275 213 1279
rect 207 1274 213 1275
rect 242 1279 253 1280
rect 242 1275 243 1279
rect 247 1275 248 1279
rect 252 1275 253 1279
rect 242 1274 253 1275
rect 295 1279 301 1280
rect 295 1275 296 1279
rect 300 1278 301 1279
rect 303 1279 309 1280
rect 303 1278 304 1279
rect 300 1276 304 1278
rect 300 1275 301 1276
rect 295 1274 301 1275
rect 303 1275 304 1276
rect 308 1275 309 1279
rect 303 1274 309 1275
rect 343 1279 349 1280
rect 343 1275 344 1279
rect 348 1278 349 1279
rect 351 1279 357 1280
rect 351 1278 352 1279
rect 348 1276 352 1278
rect 348 1275 349 1276
rect 343 1274 349 1275
rect 351 1275 352 1276
rect 356 1275 357 1279
rect 351 1274 357 1275
rect 390 1279 397 1280
rect 390 1275 391 1279
rect 396 1275 397 1279
rect 390 1274 397 1275
rect 447 1279 456 1280
rect 447 1275 448 1279
rect 455 1275 456 1279
rect 484 1278 498 1280
rect 503 1279 509 1280
rect 503 1278 504 1279
rect 496 1276 504 1278
rect 447 1274 456 1275
rect 503 1275 504 1276
rect 508 1275 509 1279
rect 552 1278 554 1296
rect 559 1295 565 1296
rect 559 1291 560 1295
rect 564 1294 565 1295
rect 598 1295 604 1296
rect 598 1294 599 1295
rect 564 1292 599 1294
rect 564 1291 565 1292
rect 559 1290 565 1291
rect 598 1291 599 1292
rect 603 1291 604 1295
rect 622 1295 629 1296
rect 622 1291 623 1295
rect 628 1291 629 1295
rect 631 1295 632 1299
rect 636 1298 637 1299
rect 799 1299 805 1300
rect 636 1296 683 1298
rect 636 1295 637 1296
rect 631 1294 637 1295
rect 679 1295 685 1296
rect 679 1291 680 1295
rect 684 1291 685 1295
rect 734 1295 741 1296
rect 734 1291 735 1295
rect 740 1291 741 1295
rect 782 1295 788 1296
rect 782 1291 783 1295
rect 787 1294 788 1295
rect 791 1295 797 1296
rect 791 1294 792 1295
rect 787 1292 792 1294
rect 787 1291 788 1292
rect 598 1290 604 1291
rect 606 1290 612 1291
rect 622 1290 629 1291
rect 662 1290 668 1291
rect 679 1290 685 1291
rect 718 1290 724 1291
rect 734 1290 741 1291
rect 774 1290 780 1291
rect 782 1290 788 1291
rect 791 1291 792 1292
rect 796 1291 797 1295
rect 799 1295 800 1299
rect 804 1298 805 1299
rect 855 1299 861 1300
rect 804 1296 842 1298
rect 804 1295 805 1296
rect 799 1294 805 1295
rect 840 1294 842 1296
rect 847 1295 853 1296
rect 847 1294 848 1295
rect 840 1292 848 1294
rect 847 1291 848 1292
rect 852 1291 853 1295
rect 855 1295 856 1299
rect 860 1298 861 1299
rect 919 1299 925 1300
rect 860 1296 906 1298
rect 860 1295 861 1296
rect 855 1294 861 1295
rect 904 1294 906 1296
rect 911 1295 917 1296
rect 911 1294 912 1295
rect 904 1292 912 1294
rect 911 1291 912 1292
rect 916 1291 917 1295
rect 919 1295 920 1299
rect 924 1298 925 1299
rect 983 1299 989 1300
rect 924 1296 970 1298
rect 924 1295 925 1296
rect 919 1294 925 1295
rect 968 1294 970 1296
rect 975 1295 981 1296
rect 975 1294 976 1295
rect 968 1292 976 1294
rect 975 1291 976 1292
rect 980 1291 981 1295
rect 983 1295 984 1299
rect 988 1298 989 1299
rect 1047 1299 1053 1300
rect 988 1296 1034 1298
rect 988 1295 989 1296
rect 983 1294 989 1295
rect 1032 1294 1034 1296
rect 1039 1295 1045 1296
rect 1039 1294 1040 1295
rect 1032 1292 1040 1294
rect 1039 1291 1040 1292
rect 1044 1291 1045 1295
rect 1047 1295 1048 1299
rect 1052 1298 1053 1299
rect 1383 1299 1389 1300
rect 1052 1296 1090 1298
rect 1200 1296 1218 1298
rect 1272 1296 1290 1298
rect 1052 1295 1053 1296
rect 1047 1294 1053 1295
rect 1088 1294 1090 1296
rect 1095 1295 1101 1296
rect 1095 1294 1096 1295
rect 1088 1292 1096 1294
rect 1095 1291 1096 1292
rect 1100 1291 1101 1295
rect 1159 1295 1165 1296
rect 1159 1291 1160 1295
rect 1164 1294 1165 1295
rect 1200 1294 1202 1296
rect 1164 1292 1202 1294
rect 1164 1291 1165 1292
rect 791 1290 797 1291
rect 830 1290 836 1291
rect 847 1290 853 1291
rect 894 1290 900 1291
rect 911 1290 917 1291
rect 958 1290 964 1291
rect 975 1290 981 1291
rect 1022 1290 1028 1291
rect 1039 1290 1045 1291
rect 1078 1290 1084 1291
rect 1095 1290 1101 1291
rect 1142 1290 1148 1291
rect 1159 1290 1165 1291
rect 1206 1290 1212 1291
rect 606 1286 607 1290
rect 611 1286 612 1290
rect 606 1285 612 1286
rect 662 1286 663 1290
rect 667 1286 668 1290
rect 662 1285 668 1286
rect 718 1286 719 1290
rect 723 1286 724 1290
rect 718 1285 724 1286
rect 774 1286 775 1290
rect 779 1286 780 1290
rect 774 1285 780 1286
rect 830 1286 831 1290
rect 835 1286 836 1290
rect 830 1285 836 1286
rect 894 1286 895 1290
rect 899 1286 900 1290
rect 894 1285 900 1286
rect 958 1286 959 1290
rect 963 1286 964 1290
rect 958 1285 964 1286
rect 1022 1286 1023 1290
rect 1027 1286 1028 1290
rect 1022 1285 1028 1286
rect 1078 1286 1079 1290
rect 1083 1286 1084 1290
rect 1078 1285 1084 1286
rect 1142 1286 1143 1290
rect 1147 1286 1148 1290
rect 1142 1285 1148 1286
rect 1206 1286 1207 1290
rect 1211 1286 1212 1290
rect 1206 1285 1212 1286
rect 559 1279 565 1280
rect 559 1278 560 1279
rect 552 1276 560 1278
rect 503 1274 509 1275
rect 559 1275 560 1276
rect 564 1275 565 1279
rect 559 1274 565 1275
rect 623 1279 629 1280
rect 623 1275 624 1279
rect 628 1278 629 1279
rect 631 1279 637 1280
rect 631 1278 632 1279
rect 628 1276 632 1278
rect 628 1275 629 1276
rect 623 1274 629 1275
rect 631 1275 632 1276
rect 636 1275 637 1279
rect 631 1274 637 1275
rect 679 1279 685 1280
rect 679 1275 680 1279
rect 684 1275 685 1279
rect 679 1274 685 1275
rect 735 1279 741 1280
rect 735 1275 736 1279
rect 740 1278 741 1279
rect 758 1279 764 1280
rect 758 1278 759 1279
rect 740 1276 759 1278
rect 740 1275 741 1276
rect 735 1274 741 1275
rect 758 1275 759 1276
rect 763 1275 764 1279
rect 758 1274 764 1275
rect 791 1279 797 1280
rect 791 1275 792 1279
rect 796 1278 797 1279
rect 799 1279 805 1280
rect 799 1278 800 1279
rect 796 1276 800 1278
rect 796 1275 797 1276
rect 791 1274 797 1275
rect 799 1275 800 1276
rect 804 1275 805 1279
rect 799 1274 805 1275
rect 847 1279 853 1280
rect 847 1275 848 1279
rect 852 1278 853 1279
rect 855 1279 861 1280
rect 855 1278 856 1279
rect 852 1276 856 1278
rect 852 1275 853 1276
rect 847 1274 853 1275
rect 855 1275 856 1276
rect 860 1275 861 1279
rect 855 1274 861 1275
rect 911 1279 917 1280
rect 911 1275 912 1279
rect 916 1278 917 1279
rect 919 1279 925 1280
rect 919 1278 920 1279
rect 916 1276 920 1278
rect 916 1275 917 1276
rect 911 1274 917 1275
rect 919 1275 920 1276
rect 924 1275 925 1279
rect 919 1274 925 1275
rect 975 1279 981 1280
rect 975 1275 976 1279
rect 980 1278 981 1279
rect 983 1279 989 1280
rect 983 1278 984 1279
rect 980 1276 984 1278
rect 980 1275 981 1276
rect 975 1274 981 1275
rect 983 1275 984 1276
rect 988 1275 989 1279
rect 983 1274 989 1275
rect 1039 1279 1045 1280
rect 1039 1275 1040 1279
rect 1044 1278 1045 1279
rect 1047 1279 1053 1280
rect 1047 1278 1048 1279
rect 1044 1276 1048 1278
rect 1044 1275 1045 1276
rect 1039 1274 1045 1275
rect 1047 1275 1048 1276
rect 1052 1275 1053 1279
rect 1047 1274 1053 1275
rect 1094 1279 1101 1280
rect 1094 1275 1095 1279
rect 1100 1275 1101 1279
rect 1094 1274 1101 1275
rect 1154 1279 1165 1280
rect 1154 1275 1155 1279
rect 1159 1275 1160 1279
rect 1164 1275 1165 1279
rect 1216 1278 1218 1296
rect 1223 1295 1229 1296
rect 1223 1291 1224 1295
rect 1228 1294 1229 1295
rect 1272 1294 1274 1296
rect 1228 1292 1274 1294
rect 1228 1291 1229 1292
rect 1223 1290 1229 1291
rect 1278 1290 1284 1291
rect 1278 1286 1279 1290
rect 1283 1286 1284 1290
rect 1278 1285 1284 1286
rect 1223 1279 1229 1280
rect 1223 1278 1224 1279
rect 1216 1276 1224 1278
rect 1154 1274 1165 1275
rect 1223 1275 1224 1276
rect 1228 1275 1229 1279
rect 1288 1278 1290 1296
rect 1295 1295 1301 1296
rect 1295 1291 1296 1295
rect 1300 1294 1301 1295
rect 1350 1295 1356 1296
rect 1350 1294 1351 1295
rect 1300 1292 1351 1294
rect 1300 1291 1301 1292
rect 1295 1290 1301 1291
rect 1350 1291 1351 1292
rect 1355 1291 1356 1295
rect 1374 1295 1381 1296
rect 1374 1291 1375 1295
rect 1380 1291 1381 1295
rect 1383 1295 1384 1299
rect 1388 1298 1389 1299
rect 1471 1299 1477 1300
rect 1388 1296 1458 1298
rect 1388 1295 1389 1296
rect 1383 1294 1389 1295
rect 1456 1294 1458 1296
rect 1463 1295 1469 1296
rect 1463 1294 1464 1295
rect 1456 1292 1464 1294
rect 1463 1291 1464 1292
rect 1468 1291 1469 1295
rect 1471 1295 1472 1299
rect 1476 1298 1477 1299
rect 1476 1296 1554 1298
rect 1476 1295 1477 1296
rect 1471 1294 1477 1295
rect 1552 1294 1554 1296
rect 1559 1295 1565 1296
rect 1559 1294 1560 1295
rect 1552 1292 1560 1294
rect 1559 1291 1560 1292
rect 1564 1291 1565 1295
rect 1639 1295 1645 1296
rect 1639 1291 1640 1295
rect 1644 1294 1645 1295
rect 1647 1295 1653 1296
rect 1647 1294 1648 1295
rect 1644 1292 1648 1294
rect 1644 1291 1645 1292
rect 1350 1290 1356 1291
rect 1358 1290 1364 1291
rect 1374 1290 1381 1291
rect 1446 1290 1452 1291
rect 1463 1290 1469 1291
rect 1542 1290 1548 1291
rect 1559 1290 1565 1291
rect 1622 1290 1628 1291
rect 1639 1290 1645 1291
rect 1647 1291 1648 1292
rect 1652 1291 1653 1295
rect 1647 1290 1653 1291
rect 1662 1292 1668 1293
rect 1358 1286 1359 1290
rect 1363 1286 1364 1290
rect 1358 1285 1364 1286
rect 1446 1286 1447 1290
rect 1451 1286 1452 1290
rect 1446 1285 1452 1286
rect 1542 1286 1543 1290
rect 1547 1286 1548 1290
rect 1542 1285 1548 1286
rect 1622 1286 1623 1290
rect 1627 1286 1628 1290
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1622 1285 1628 1286
rect 1295 1279 1301 1280
rect 1295 1278 1296 1279
rect 1288 1276 1296 1278
rect 1223 1274 1229 1275
rect 1295 1275 1296 1276
rect 1300 1275 1301 1279
rect 1295 1274 1301 1275
rect 1375 1279 1381 1280
rect 1375 1275 1376 1279
rect 1380 1278 1381 1279
rect 1383 1279 1389 1280
rect 1383 1278 1384 1279
rect 1380 1276 1384 1278
rect 1380 1275 1381 1276
rect 1375 1274 1381 1275
rect 1383 1275 1384 1276
rect 1388 1275 1389 1279
rect 1383 1274 1389 1275
rect 1463 1279 1469 1280
rect 1463 1275 1464 1279
rect 1468 1278 1469 1279
rect 1471 1279 1477 1280
rect 1471 1278 1472 1279
rect 1468 1276 1472 1278
rect 1468 1275 1469 1276
rect 1463 1274 1469 1275
rect 1471 1275 1472 1276
rect 1476 1275 1477 1279
rect 1559 1279 1565 1280
rect 1559 1278 1560 1279
rect 1471 1274 1477 1275
rect 1552 1276 1560 1278
rect 110 1270 116 1271
rect 134 1273 140 1274
rect 134 1269 135 1273
rect 139 1269 140 1273
rect 134 1268 140 1269
rect 182 1273 188 1274
rect 182 1269 183 1273
rect 187 1269 188 1273
rect 182 1268 188 1269
rect 230 1273 236 1274
rect 230 1269 231 1273
rect 235 1269 236 1273
rect 230 1268 236 1269
rect 278 1273 284 1274
rect 278 1269 279 1273
rect 283 1269 284 1273
rect 278 1268 284 1269
rect 326 1273 332 1274
rect 326 1269 327 1273
rect 331 1269 332 1273
rect 326 1268 332 1269
rect 374 1273 380 1274
rect 374 1269 375 1273
rect 379 1269 380 1273
rect 374 1268 380 1269
rect 430 1273 436 1274
rect 430 1269 431 1273
rect 435 1269 436 1273
rect 430 1268 436 1269
rect 486 1273 492 1274
rect 486 1269 487 1273
rect 491 1269 492 1273
rect 486 1268 492 1269
rect 542 1273 548 1274
rect 542 1269 543 1273
rect 547 1269 548 1273
rect 542 1268 548 1269
rect 606 1273 612 1274
rect 606 1269 607 1273
rect 611 1269 612 1273
rect 606 1268 612 1269
rect 662 1273 668 1274
rect 662 1269 663 1273
rect 667 1269 668 1273
rect 662 1268 668 1269
rect 598 1267 604 1268
rect 598 1263 599 1267
rect 603 1266 604 1267
rect 681 1266 683 1274
rect 718 1273 724 1274
rect 718 1269 719 1273
rect 723 1269 724 1273
rect 718 1268 724 1269
rect 774 1273 780 1274
rect 774 1269 775 1273
rect 779 1269 780 1273
rect 774 1268 780 1269
rect 830 1273 836 1274
rect 830 1269 831 1273
rect 835 1269 836 1273
rect 830 1268 836 1269
rect 894 1273 900 1274
rect 894 1269 895 1273
rect 899 1269 900 1273
rect 894 1268 900 1269
rect 958 1273 964 1274
rect 958 1269 959 1273
rect 963 1269 964 1273
rect 958 1268 964 1269
rect 1022 1273 1028 1274
rect 1022 1269 1023 1273
rect 1027 1269 1028 1273
rect 1022 1268 1028 1269
rect 1078 1273 1084 1274
rect 1078 1269 1079 1273
rect 1083 1269 1084 1273
rect 1078 1268 1084 1269
rect 1142 1273 1148 1274
rect 1142 1269 1143 1273
rect 1147 1269 1148 1273
rect 1142 1268 1148 1269
rect 1206 1273 1212 1274
rect 1206 1269 1207 1273
rect 1211 1269 1212 1273
rect 1206 1268 1212 1269
rect 1278 1273 1284 1274
rect 1278 1269 1279 1273
rect 1283 1269 1284 1273
rect 1278 1268 1284 1269
rect 1358 1273 1364 1274
rect 1358 1269 1359 1273
rect 1363 1269 1364 1273
rect 1358 1268 1364 1269
rect 1446 1273 1452 1274
rect 1446 1269 1447 1273
rect 1451 1269 1452 1273
rect 1446 1268 1452 1269
rect 1542 1273 1548 1274
rect 1542 1269 1543 1273
rect 1547 1269 1548 1273
rect 1542 1268 1548 1269
rect 603 1264 683 1266
rect 1350 1267 1356 1268
rect 603 1263 604 1264
rect 598 1262 604 1263
rect 1350 1263 1351 1267
rect 1355 1266 1356 1267
rect 1552 1266 1554 1276
rect 1559 1275 1560 1276
rect 1564 1275 1565 1279
rect 1559 1274 1565 1275
rect 1639 1279 1648 1280
rect 1639 1275 1640 1279
rect 1647 1275 1648 1279
rect 1639 1274 1648 1275
rect 1662 1275 1668 1276
rect 1622 1273 1628 1274
rect 1622 1269 1623 1273
rect 1627 1269 1628 1273
rect 1662 1271 1663 1275
rect 1667 1271 1668 1275
rect 1662 1270 1668 1271
rect 1622 1268 1628 1269
rect 1355 1264 1554 1266
rect 1355 1263 1356 1264
rect 1350 1262 1356 1263
rect 134 1259 140 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 134 1255 135 1259
rect 139 1255 140 1259
rect 134 1254 140 1255
rect 166 1259 172 1260
rect 166 1255 167 1259
rect 171 1255 172 1259
rect 166 1254 172 1255
rect 222 1259 228 1260
rect 222 1255 223 1259
rect 227 1255 228 1259
rect 222 1254 228 1255
rect 278 1259 284 1260
rect 278 1255 279 1259
rect 283 1255 284 1259
rect 278 1254 284 1255
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 382 1259 388 1260
rect 382 1255 383 1259
rect 387 1255 388 1259
rect 382 1254 388 1255
rect 438 1259 444 1260
rect 438 1255 439 1259
rect 443 1255 444 1259
rect 438 1254 444 1255
rect 494 1259 500 1260
rect 494 1255 495 1259
rect 499 1255 500 1259
rect 494 1254 500 1255
rect 550 1259 556 1260
rect 550 1255 551 1259
rect 555 1255 556 1259
rect 550 1254 556 1255
rect 606 1259 612 1260
rect 606 1255 607 1259
rect 611 1255 612 1259
rect 606 1254 612 1255
rect 662 1259 668 1260
rect 662 1255 663 1259
rect 667 1255 668 1259
rect 662 1254 668 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 766 1259 772 1260
rect 766 1255 767 1259
rect 771 1255 772 1259
rect 766 1254 772 1255
rect 814 1259 820 1260
rect 814 1255 815 1259
rect 819 1255 820 1259
rect 814 1254 820 1255
rect 870 1259 876 1260
rect 870 1255 871 1259
rect 875 1255 876 1259
rect 870 1254 876 1255
rect 926 1259 932 1260
rect 926 1255 927 1259
rect 931 1255 932 1259
rect 926 1254 932 1255
rect 982 1259 988 1260
rect 982 1255 983 1259
rect 987 1255 988 1259
rect 982 1254 988 1255
rect 1038 1259 1044 1260
rect 1038 1255 1039 1259
rect 1043 1255 1044 1259
rect 1038 1254 1044 1255
rect 1094 1259 1100 1260
rect 1094 1255 1095 1259
rect 1099 1255 1100 1259
rect 1094 1254 1100 1255
rect 1158 1259 1164 1260
rect 1158 1255 1159 1259
rect 1163 1255 1164 1259
rect 1158 1254 1164 1255
rect 1230 1259 1236 1260
rect 1230 1255 1231 1259
rect 1235 1255 1236 1259
rect 1230 1254 1236 1255
rect 1318 1259 1324 1260
rect 1318 1255 1319 1259
rect 1323 1255 1324 1259
rect 1318 1254 1324 1255
rect 1422 1259 1428 1260
rect 1422 1255 1423 1259
rect 1427 1255 1428 1259
rect 1422 1254 1428 1255
rect 1534 1259 1540 1260
rect 1534 1255 1535 1259
rect 1539 1255 1540 1259
rect 1534 1254 1540 1255
rect 1622 1259 1628 1260
rect 1622 1255 1623 1259
rect 1627 1255 1628 1259
rect 1622 1254 1628 1255
rect 1662 1257 1668 1258
rect 110 1252 116 1253
rect 1662 1253 1663 1257
rect 1667 1253 1668 1257
rect 1662 1252 1668 1253
rect 150 1251 157 1252
rect 150 1247 151 1251
rect 156 1247 157 1251
rect 183 1251 189 1252
rect 183 1250 184 1251
rect 150 1246 157 1247
rect 176 1248 184 1250
rect 134 1242 140 1243
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 134 1238 135 1242
rect 139 1238 140 1242
rect 134 1237 140 1238
rect 166 1242 172 1243
rect 166 1238 167 1242
rect 171 1238 172 1242
rect 166 1237 172 1238
rect 110 1235 116 1236
rect 151 1235 157 1236
rect 151 1231 152 1235
rect 156 1234 157 1235
rect 176 1234 178 1248
rect 183 1247 184 1248
rect 188 1247 189 1251
rect 239 1251 245 1252
rect 239 1250 240 1251
rect 183 1246 189 1247
rect 212 1248 240 1250
rect 156 1232 178 1234
rect 183 1235 189 1236
rect 156 1231 157 1232
rect 151 1230 157 1231
rect 183 1231 184 1235
rect 188 1234 189 1235
rect 212 1234 214 1248
rect 239 1247 240 1248
rect 244 1247 245 1251
rect 239 1246 245 1247
rect 294 1251 301 1252
rect 294 1247 295 1251
rect 300 1247 301 1251
rect 343 1251 349 1252
rect 343 1250 344 1251
rect 294 1246 301 1247
rect 319 1248 344 1250
rect 222 1242 228 1243
rect 222 1238 223 1242
rect 227 1238 228 1242
rect 222 1237 228 1238
rect 278 1242 284 1243
rect 278 1238 279 1242
rect 283 1238 284 1242
rect 278 1237 284 1238
rect 188 1232 214 1234
rect 239 1235 248 1236
rect 188 1231 189 1232
rect 183 1230 189 1231
rect 239 1231 240 1235
rect 247 1231 248 1235
rect 239 1230 248 1231
rect 295 1235 301 1236
rect 295 1231 296 1235
rect 300 1234 301 1235
rect 319 1234 321 1248
rect 343 1247 344 1248
rect 348 1247 349 1251
rect 399 1251 405 1252
rect 399 1250 400 1251
rect 343 1246 349 1247
rect 372 1248 400 1250
rect 326 1242 332 1243
rect 326 1238 327 1242
rect 331 1238 332 1242
rect 326 1237 332 1238
rect 300 1232 321 1234
rect 343 1235 349 1236
rect 300 1231 301 1232
rect 295 1230 301 1231
rect 343 1231 344 1235
rect 348 1234 349 1235
rect 372 1234 374 1248
rect 399 1247 400 1248
rect 404 1247 405 1251
rect 399 1246 405 1247
rect 455 1251 461 1252
rect 455 1247 456 1251
rect 460 1250 461 1251
rect 511 1251 517 1252
rect 460 1248 486 1250
rect 460 1247 461 1248
rect 455 1246 461 1247
rect 382 1242 388 1243
rect 382 1238 383 1242
rect 387 1238 388 1242
rect 382 1237 388 1238
rect 438 1242 444 1243
rect 438 1238 439 1242
rect 443 1238 444 1242
rect 438 1237 444 1238
rect 348 1232 374 1234
rect 398 1235 405 1236
rect 348 1231 349 1232
rect 343 1230 349 1231
rect 398 1231 399 1235
rect 404 1231 405 1235
rect 398 1230 405 1231
rect 450 1235 461 1236
rect 450 1231 451 1235
rect 455 1231 456 1235
rect 460 1231 461 1235
rect 484 1234 486 1248
rect 511 1247 512 1251
rect 516 1250 517 1251
rect 567 1251 573 1252
rect 516 1248 542 1250
rect 516 1247 517 1248
rect 511 1246 517 1247
rect 494 1242 500 1243
rect 494 1238 495 1242
rect 499 1238 500 1242
rect 494 1237 500 1238
rect 511 1235 517 1236
rect 511 1234 512 1235
rect 484 1232 512 1234
rect 450 1230 461 1231
rect 511 1231 512 1232
rect 516 1231 517 1235
rect 540 1234 542 1248
rect 567 1247 568 1251
rect 572 1250 573 1251
rect 618 1251 629 1252
rect 572 1248 598 1250
rect 572 1247 573 1248
rect 567 1246 573 1247
rect 550 1242 556 1243
rect 550 1238 551 1242
rect 555 1238 556 1242
rect 550 1237 556 1238
rect 567 1235 573 1236
rect 567 1234 568 1235
rect 540 1232 568 1234
rect 511 1230 517 1231
rect 567 1231 568 1232
rect 572 1231 573 1235
rect 596 1234 598 1248
rect 618 1247 619 1251
rect 623 1247 624 1251
rect 628 1247 629 1251
rect 618 1246 629 1247
rect 679 1251 685 1252
rect 679 1247 680 1251
rect 684 1250 685 1251
rect 734 1251 741 1252
rect 684 1248 730 1250
rect 684 1247 685 1248
rect 679 1246 685 1247
rect 606 1242 612 1243
rect 606 1238 607 1242
rect 611 1238 612 1242
rect 606 1237 612 1238
rect 662 1242 668 1243
rect 662 1238 663 1242
rect 667 1238 668 1242
rect 662 1237 668 1238
rect 718 1242 724 1243
rect 718 1238 719 1242
rect 723 1238 724 1242
rect 718 1237 724 1238
rect 623 1235 629 1236
rect 623 1234 624 1235
rect 596 1232 624 1234
rect 567 1230 573 1231
rect 623 1231 624 1232
rect 628 1231 629 1235
rect 623 1230 629 1231
rect 679 1235 685 1236
rect 679 1231 680 1235
rect 684 1231 685 1235
rect 728 1234 730 1248
rect 734 1247 735 1251
rect 740 1247 741 1251
rect 734 1246 741 1247
rect 782 1251 789 1252
rect 782 1247 783 1251
rect 788 1247 789 1251
rect 782 1246 789 1247
rect 791 1251 797 1252
rect 791 1247 792 1251
rect 796 1250 797 1251
rect 831 1251 837 1252
rect 831 1250 832 1251
rect 796 1248 832 1250
rect 796 1247 797 1248
rect 791 1246 797 1247
rect 831 1247 832 1248
rect 836 1247 837 1251
rect 887 1251 893 1252
rect 887 1250 888 1251
rect 831 1246 837 1247
rect 860 1248 888 1250
rect 766 1242 772 1243
rect 766 1238 767 1242
rect 771 1238 772 1242
rect 766 1237 772 1238
rect 814 1242 820 1243
rect 814 1238 815 1242
rect 819 1238 820 1242
rect 814 1237 820 1238
rect 735 1235 741 1236
rect 735 1234 736 1235
rect 728 1232 736 1234
rect 679 1230 685 1231
rect 735 1231 736 1232
rect 740 1231 741 1235
rect 735 1230 741 1231
rect 758 1235 764 1236
rect 758 1231 759 1235
rect 763 1234 764 1235
rect 783 1235 789 1236
rect 783 1234 784 1235
rect 763 1232 784 1234
rect 763 1231 764 1232
rect 758 1230 764 1231
rect 783 1231 784 1232
rect 788 1231 789 1235
rect 783 1230 789 1231
rect 831 1235 837 1236
rect 831 1231 832 1235
rect 836 1234 837 1235
rect 860 1234 862 1248
rect 887 1247 888 1248
rect 892 1247 893 1251
rect 887 1246 893 1247
rect 943 1251 949 1252
rect 943 1247 944 1251
rect 948 1250 949 1251
rect 999 1251 1005 1252
rect 948 1248 974 1250
rect 948 1247 949 1248
rect 943 1246 949 1247
rect 870 1242 876 1243
rect 870 1238 871 1242
rect 875 1238 876 1242
rect 870 1237 876 1238
rect 926 1242 932 1243
rect 926 1238 927 1242
rect 931 1238 932 1242
rect 926 1237 932 1238
rect 836 1232 862 1234
rect 887 1235 893 1236
rect 836 1231 837 1232
rect 831 1230 837 1231
rect 887 1231 888 1235
rect 892 1234 893 1235
rect 906 1235 912 1236
rect 892 1232 902 1234
rect 892 1231 893 1232
rect 887 1230 893 1231
rect 681 1226 683 1230
rect 791 1227 797 1228
rect 791 1226 792 1227
rect 681 1224 792 1226
rect 618 1223 624 1224
rect 618 1222 619 1223
rect 448 1220 619 1222
rect 191 1215 197 1216
rect 160 1212 187 1214
rect 150 1211 157 1212
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 150 1207 151 1211
rect 156 1207 157 1211
rect 110 1203 116 1204
rect 134 1206 140 1207
rect 150 1206 157 1207
rect 134 1202 135 1206
rect 139 1202 140 1206
rect 134 1201 140 1202
rect 151 1195 157 1196
rect 110 1191 116 1192
rect 110 1187 111 1191
rect 115 1187 116 1191
rect 151 1191 152 1195
rect 156 1194 157 1195
rect 160 1194 162 1212
rect 183 1211 189 1212
rect 183 1207 184 1211
rect 188 1207 189 1211
rect 191 1211 192 1215
rect 196 1214 197 1215
rect 306 1215 312 1216
rect 196 1212 243 1214
rect 196 1211 197 1212
rect 191 1210 197 1211
rect 239 1211 245 1212
rect 239 1207 240 1211
rect 244 1207 245 1211
rect 295 1211 304 1212
rect 295 1207 296 1211
rect 303 1207 304 1211
rect 306 1211 307 1215
rect 311 1214 312 1215
rect 359 1215 365 1216
rect 311 1212 346 1214
rect 311 1211 312 1212
rect 306 1210 312 1211
rect 344 1210 346 1212
rect 351 1211 357 1212
rect 351 1210 352 1211
rect 344 1208 352 1210
rect 351 1207 352 1208
rect 356 1207 357 1211
rect 359 1211 360 1215
rect 364 1214 365 1215
rect 364 1212 394 1214
rect 448 1212 450 1220
rect 618 1219 619 1220
rect 623 1219 624 1223
rect 791 1223 792 1224
rect 796 1223 797 1227
rect 900 1226 902 1232
rect 906 1231 907 1235
rect 911 1234 912 1235
rect 943 1235 949 1236
rect 943 1234 944 1235
rect 911 1232 944 1234
rect 911 1231 912 1232
rect 906 1230 912 1231
rect 943 1231 944 1232
rect 948 1231 949 1235
rect 972 1234 974 1248
rect 999 1247 1000 1251
rect 1004 1250 1005 1251
rect 1050 1251 1061 1252
rect 1004 1248 1030 1250
rect 1004 1247 1005 1248
rect 999 1246 1005 1247
rect 982 1242 988 1243
rect 982 1238 983 1242
rect 987 1238 988 1242
rect 982 1237 988 1238
rect 999 1235 1005 1236
rect 999 1234 1000 1235
rect 972 1232 1000 1234
rect 943 1230 949 1231
rect 999 1231 1000 1232
rect 1004 1231 1005 1235
rect 1028 1234 1030 1248
rect 1050 1247 1051 1251
rect 1055 1247 1056 1251
rect 1060 1247 1061 1251
rect 1050 1246 1061 1247
rect 1111 1251 1117 1252
rect 1111 1247 1112 1251
rect 1116 1250 1117 1251
rect 1175 1251 1181 1252
rect 1116 1248 1170 1250
rect 1116 1247 1117 1248
rect 1111 1246 1117 1247
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1038 1237 1044 1238
rect 1094 1242 1100 1243
rect 1094 1238 1095 1242
rect 1099 1238 1100 1242
rect 1094 1237 1100 1238
rect 1158 1242 1164 1243
rect 1158 1238 1159 1242
rect 1163 1238 1164 1242
rect 1158 1237 1164 1238
rect 1055 1235 1061 1236
rect 1055 1234 1056 1235
rect 1028 1232 1056 1234
rect 999 1230 1005 1231
rect 1055 1231 1056 1232
rect 1060 1231 1061 1235
rect 1055 1230 1061 1231
rect 1111 1235 1117 1236
rect 1111 1231 1112 1235
rect 1116 1234 1117 1235
rect 1150 1235 1156 1236
rect 1150 1234 1151 1235
rect 1116 1232 1151 1234
rect 1116 1231 1117 1232
rect 1111 1230 1117 1231
rect 1150 1231 1151 1232
rect 1155 1231 1156 1235
rect 1168 1234 1170 1248
rect 1175 1247 1176 1251
rect 1180 1250 1181 1251
rect 1247 1251 1253 1252
rect 1180 1248 1242 1250
rect 1180 1247 1181 1248
rect 1175 1246 1181 1247
rect 1230 1242 1236 1243
rect 1230 1238 1231 1242
rect 1235 1238 1236 1242
rect 1230 1237 1236 1238
rect 1175 1235 1181 1236
rect 1175 1234 1176 1235
rect 1168 1232 1176 1234
rect 1150 1230 1156 1231
rect 1175 1231 1176 1232
rect 1180 1231 1181 1235
rect 1240 1234 1242 1248
rect 1247 1247 1248 1251
rect 1252 1250 1253 1251
rect 1335 1251 1341 1252
rect 1252 1248 1294 1250
rect 1252 1247 1253 1248
rect 1247 1246 1253 1247
rect 1247 1235 1253 1236
rect 1247 1234 1248 1235
rect 1240 1232 1248 1234
rect 1175 1230 1181 1231
rect 1247 1231 1248 1232
rect 1252 1231 1253 1235
rect 1292 1234 1294 1248
rect 1335 1247 1336 1251
rect 1340 1250 1341 1251
rect 1439 1251 1445 1252
rect 1340 1248 1390 1250
rect 1340 1247 1341 1248
rect 1335 1246 1341 1247
rect 1318 1242 1324 1243
rect 1318 1238 1319 1242
rect 1323 1238 1324 1242
rect 1318 1237 1324 1238
rect 1335 1235 1341 1236
rect 1335 1234 1336 1235
rect 1292 1232 1336 1234
rect 1247 1230 1253 1231
rect 1335 1231 1336 1232
rect 1340 1231 1341 1235
rect 1388 1234 1390 1248
rect 1439 1247 1440 1251
rect 1444 1250 1445 1251
rect 1502 1251 1508 1252
rect 1444 1248 1498 1250
rect 1444 1247 1445 1248
rect 1439 1246 1445 1247
rect 1422 1242 1428 1243
rect 1422 1238 1423 1242
rect 1427 1238 1428 1242
rect 1422 1237 1428 1238
rect 1439 1235 1445 1236
rect 1439 1234 1440 1235
rect 1388 1232 1440 1234
rect 1335 1230 1341 1231
rect 1439 1231 1440 1232
rect 1444 1231 1445 1235
rect 1496 1234 1498 1248
rect 1502 1247 1503 1251
rect 1507 1250 1508 1251
rect 1551 1251 1557 1252
rect 1551 1250 1552 1251
rect 1507 1248 1552 1250
rect 1507 1247 1508 1248
rect 1502 1246 1508 1247
rect 1551 1247 1552 1248
rect 1556 1247 1557 1251
rect 1551 1246 1557 1247
rect 1638 1251 1645 1252
rect 1638 1247 1639 1251
rect 1644 1247 1645 1251
rect 1638 1246 1645 1247
rect 1534 1242 1540 1243
rect 1534 1238 1535 1242
rect 1539 1238 1540 1242
rect 1534 1237 1540 1238
rect 1622 1242 1628 1243
rect 1622 1238 1623 1242
rect 1627 1238 1628 1242
rect 1622 1237 1628 1238
rect 1662 1240 1668 1241
rect 1662 1236 1663 1240
rect 1667 1236 1668 1240
rect 1551 1235 1557 1236
rect 1551 1234 1552 1235
rect 1496 1232 1552 1234
rect 1439 1230 1445 1231
rect 1551 1231 1552 1232
rect 1556 1231 1557 1235
rect 1551 1230 1557 1231
rect 1639 1235 1645 1236
rect 1639 1231 1640 1235
rect 1644 1234 1645 1235
rect 1650 1235 1656 1236
rect 1662 1235 1668 1236
rect 1650 1234 1651 1235
rect 1644 1232 1651 1234
rect 1644 1231 1645 1232
rect 1639 1230 1645 1231
rect 1650 1231 1651 1232
rect 1655 1231 1656 1235
rect 1650 1230 1656 1231
rect 1050 1227 1056 1228
rect 1050 1226 1051 1227
rect 900 1224 1051 1226
rect 791 1222 797 1223
rect 1050 1223 1051 1224
rect 1055 1223 1056 1227
rect 1050 1222 1056 1223
rect 1502 1223 1508 1224
rect 1502 1222 1503 1223
rect 618 1218 624 1219
rect 1160 1220 1503 1222
rect 455 1215 461 1216
rect 364 1211 365 1212
rect 359 1210 365 1211
rect 392 1210 394 1212
rect 399 1211 405 1212
rect 399 1210 400 1211
rect 392 1208 400 1210
rect 399 1207 400 1208
rect 404 1207 405 1211
rect 447 1211 453 1212
rect 447 1207 448 1211
rect 452 1207 453 1211
rect 455 1211 456 1215
rect 460 1214 461 1215
rect 511 1215 517 1216
rect 460 1212 498 1214
rect 460 1211 461 1212
rect 455 1210 461 1211
rect 496 1210 498 1212
rect 503 1211 509 1212
rect 503 1210 504 1211
rect 496 1208 504 1210
rect 503 1207 504 1208
rect 508 1207 509 1211
rect 511 1211 512 1215
rect 516 1214 517 1215
rect 567 1215 573 1216
rect 516 1212 554 1214
rect 516 1211 517 1212
rect 511 1210 517 1211
rect 552 1210 554 1212
rect 559 1211 565 1212
rect 559 1210 560 1211
rect 552 1208 560 1210
rect 559 1207 560 1208
rect 564 1207 565 1211
rect 567 1211 568 1215
rect 572 1214 573 1215
rect 623 1215 629 1216
rect 572 1212 619 1214
rect 572 1211 573 1212
rect 567 1210 573 1211
rect 615 1211 621 1212
rect 615 1207 616 1211
rect 620 1207 621 1211
rect 623 1211 624 1215
rect 628 1214 629 1215
rect 679 1215 685 1216
rect 628 1212 666 1214
rect 628 1211 629 1212
rect 623 1210 629 1211
rect 664 1210 666 1212
rect 671 1211 677 1212
rect 671 1210 672 1211
rect 664 1208 672 1210
rect 671 1207 672 1208
rect 676 1207 677 1211
rect 679 1211 680 1215
rect 684 1214 685 1215
rect 791 1215 797 1216
rect 684 1212 722 1214
rect 684 1211 685 1212
rect 679 1210 685 1211
rect 720 1210 722 1212
rect 727 1211 733 1212
rect 727 1210 728 1211
rect 720 1208 728 1210
rect 727 1207 728 1208
rect 732 1207 733 1211
rect 782 1211 789 1212
rect 782 1207 783 1211
rect 788 1207 789 1211
rect 791 1211 792 1215
rect 796 1214 797 1215
rect 847 1215 853 1216
rect 796 1212 834 1214
rect 796 1211 797 1212
rect 791 1210 797 1211
rect 832 1210 834 1212
rect 839 1211 845 1212
rect 839 1210 840 1211
rect 832 1208 840 1210
rect 839 1207 840 1208
rect 844 1207 845 1211
rect 847 1211 848 1215
rect 852 1214 853 1215
rect 1039 1215 1045 1216
rect 852 1212 898 1214
rect 852 1211 853 1212
rect 847 1210 853 1211
rect 896 1210 898 1212
rect 903 1211 909 1212
rect 903 1210 904 1211
rect 896 1208 904 1210
rect 903 1207 904 1208
rect 908 1207 909 1211
rect 967 1211 973 1212
rect 967 1207 968 1211
rect 972 1210 973 1211
rect 1006 1211 1012 1212
rect 1006 1210 1007 1211
rect 972 1208 1007 1210
rect 972 1207 973 1208
rect 166 1206 172 1207
rect 183 1206 189 1207
rect 222 1206 228 1207
rect 239 1206 245 1207
rect 278 1206 284 1207
rect 295 1206 304 1207
rect 334 1206 340 1207
rect 351 1206 357 1207
rect 382 1206 388 1207
rect 399 1206 405 1207
rect 430 1206 436 1207
rect 447 1206 453 1207
rect 486 1206 492 1207
rect 503 1206 509 1207
rect 542 1206 548 1207
rect 559 1206 565 1207
rect 598 1206 604 1207
rect 615 1206 621 1207
rect 654 1206 660 1207
rect 671 1206 677 1207
rect 710 1206 716 1207
rect 727 1206 733 1207
rect 766 1206 772 1207
rect 782 1206 789 1207
rect 822 1206 828 1207
rect 839 1206 845 1207
rect 886 1206 892 1207
rect 903 1206 909 1207
rect 950 1206 956 1207
rect 967 1206 973 1207
rect 1006 1207 1007 1208
rect 1011 1207 1012 1211
rect 1022 1211 1028 1212
rect 1022 1207 1023 1211
rect 1027 1210 1028 1211
rect 1031 1211 1037 1212
rect 1031 1210 1032 1211
rect 1027 1208 1032 1210
rect 1027 1207 1028 1208
rect 1006 1206 1012 1207
rect 1014 1206 1020 1207
rect 1022 1206 1028 1207
rect 1031 1207 1032 1208
rect 1036 1207 1037 1211
rect 1039 1211 1040 1215
rect 1044 1214 1045 1215
rect 1044 1212 1090 1214
rect 1160 1212 1162 1220
rect 1502 1219 1503 1220
rect 1507 1219 1508 1223
rect 1502 1218 1508 1219
rect 1167 1215 1173 1216
rect 1044 1211 1045 1212
rect 1039 1210 1045 1211
rect 1088 1210 1090 1212
rect 1095 1211 1101 1212
rect 1095 1210 1096 1211
rect 1088 1208 1096 1210
rect 1095 1207 1096 1208
rect 1100 1207 1101 1211
rect 1159 1211 1165 1212
rect 1159 1207 1160 1211
rect 1164 1207 1165 1211
rect 1167 1211 1168 1215
rect 1172 1214 1173 1215
rect 1231 1215 1237 1216
rect 1172 1212 1218 1214
rect 1172 1211 1173 1212
rect 1167 1210 1173 1211
rect 1216 1210 1218 1212
rect 1223 1211 1229 1212
rect 1223 1210 1224 1211
rect 1216 1208 1224 1210
rect 1223 1207 1224 1208
rect 1228 1207 1229 1211
rect 1231 1211 1232 1215
rect 1236 1214 1237 1215
rect 1303 1215 1309 1216
rect 1236 1212 1299 1214
rect 1236 1211 1237 1212
rect 1231 1210 1237 1211
rect 1295 1211 1301 1212
rect 1295 1207 1296 1211
rect 1300 1207 1301 1211
rect 1303 1211 1304 1215
rect 1308 1214 1309 1215
rect 1383 1215 1389 1216
rect 1308 1212 1370 1214
rect 1308 1211 1309 1212
rect 1303 1210 1309 1211
rect 1368 1210 1370 1212
rect 1375 1211 1381 1212
rect 1375 1210 1376 1211
rect 1368 1208 1376 1210
rect 1375 1207 1376 1208
rect 1380 1207 1381 1211
rect 1383 1211 1384 1215
rect 1388 1214 1389 1215
rect 1471 1215 1477 1216
rect 1388 1212 1458 1214
rect 1388 1211 1389 1212
rect 1383 1210 1389 1211
rect 1456 1210 1458 1212
rect 1463 1211 1469 1212
rect 1463 1210 1464 1211
rect 1456 1208 1464 1210
rect 1463 1207 1464 1208
rect 1468 1207 1469 1211
rect 1471 1211 1472 1215
rect 1476 1214 1477 1215
rect 1476 1212 1554 1214
rect 1476 1211 1477 1212
rect 1471 1210 1477 1211
rect 1552 1210 1554 1212
rect 1559 1211 1565 1212
rect 1559 1210 1560 1211
rect 1552 1208 1560 1210
rect 1559 1207 1560 1208
rect 1564 1207 1565 1211
rect 1638 1211 1645 1212
rect 1638 1207 1639 1211
rect 1644 1207 1645 1211
rect 1031 1206 1037 1207
rect 1078 1206 1084 1207
rect 1095 1206 1101 1207
rect 1142 1206 1148 1207
rect 1159 1206 1165 1207
rect 1206 1206 1212 1207
rect 1223 1206 1229 1207
rect 1278 1206 1284 1207
rect 1295 1206 1301 1207
rect 1358 1206 1364 1207
rect 1375 1206 1381 1207
rect 1446 1206 1452 1207
rect 1463 1206 1469 1207
rect 1542 1206 1548 1207
rect 1559 1206 1565 1207
rect 1622 1206 1628 1207
rect 1638 1206 1645 1207
rect 1662 1208 1668 1209
rect 166 1202 167 1206
rect 171 1202 172 1206
rect 166 1201 172 1202
rect 222 1202 223 1206
rect 227 1202 228 1206
rect 222 1201 228 1202
rect 278 1202 279 1206
rect 283 1202 284 1206
rect 278 1201 284 1202
rect 334 1202 335 1206
rect 339 1202 340 1206
rect 334 1201 340 1202
rect 382 1202 383 1206
rect 387 1202 388 1206
rect 382 1201 388 1202
rect 430 1202 431 1206
rect 435 1202 436 1206
rect 430 1201 436 1202
rect 486 1202 487 1206
rect 491 1202 492 1206
rect 486 1201 492 1202
rect 542 1202 543 1206
rect 547 1202 548 1206
rect 542 1201 548 1202
rect 598 1202 599 1206
rect 603 1202 604 1206
rect 598 1201 604 1202
rect 654 1202 655 1206
rect 659 1202 660 1206
rect 654 1201 660 1202
rect 710 1202 711 1206
rect 715 1202 716 1206
rect 710 1201 716 1202
rect 766 1202 767 1206
rect 771 1202 772 1206
rect 766 1201 772 1202
rect 822 1202 823 1206
rect 827 1202 828 1206
rect 822 1201 828 1202
rect 886 1202 887 1206
rect 891 1202 892 1206
rect 886 1201 892 1202
rect 950 1202 951 1206
rect 955 1202 956 1206
rect 950 1201 956 1202
rect 1014 1202 1015 1206
rect 1019 1202 1020 1206
rect 1014 1201 1020 1202
rect 1078 1202 1079 1206
rect 1083 1202 1084 1206
rect 1078 1201 1084 1202
rect 1142 1202 1143 1206
rect 1147 1202 1148 1206
rect 1142 1201 1148 1202
rect 1206 1202 1207 1206
rect 1211 1202 1212 1206
rect 1206 1201 1212 1202
rect 1278 1202 1279 1206
rect 1283 1202 1284 1206
rect 1278 1201 1284 1202
rect 1358 1202 1359 1206
rect 1363 1202 1364 1206
rect 1358 1201 1364 1202
rect 1446 1202 1447 1206
rect 1451 1202 1452 1206
rect 1446 1201 1452 1202
rect 1542 1202 1543 1206
rect 1547 1202 1548 1206
rect 1542 1201 1548 1202
rect 1622 1202 1623 1206
rect 1627 1202 1628 1206
rect 1662 1204 1663 1208
rect 1667 1204 1668 1208
rect 1662 1203 1668 1204
rect 1622 1201 1628 1202
rect 156 1192 162 1194
rect 183 1195 189 1196
rect 156 1191 157 1192
rect 151 1190 157 1191
rect 183 1191 184 1195
rect 188 1194 189 1195
rect 191 1195 197 1196
rect 191 1194 192 1195
rect 188 1192 192 1194
rect 188 1191 189 1192
rect 183 1190 189 1191
rect 191 1191 192 1192
rect 196 1191 197 1195
rect 191 1190 197 1191
rect 238 1195 245 1196
rect 238 1191 239 1195
rect 244 1191 245 1195
rect 238 1190 245 1191
rect 295 1195 301 1196
rect 295 1191 296 1195
rect 300 1194 301 1195
rect 306 1195 312 1196
rect 306 1194 307 1195
rect 300 1192 307 1194
rect 300 1191 301 1192
rect 295 1190 301 1191
rect 306 1191 307 1192
rect 311 1191 312 1195
rect 306 1190 312 1191
rect 351 1195 357 1196
rect 351 1191 352 1195
rect 356 1194 357 1195
rect 359 1195 365 1196
rect 359 1194 360 1195
rect 356 1192 360 1194
rect 356 1191 357 1192
rect 351 1190 357 1191
rect 359 1191 360 1192
rect 364 1191 365 1195
rect 359 1190 365 1191
rect 398 1195 405 1196
rect 398 1191 399 1195
rect 404 1191 405 1195
rect 398 1190 405 1191
rect 447 1195 453 1196
rect 447 1191 448 1195
rect 452 1194 453 1195
rect 455 1195 461 1196
rect 455 1194 456 1195
rect 452 1192 456 1194
rect 452 1191 453 1192
rect 447 1190 453 1191
rect 455 1191 456 1192
rect 460 1191 461 1195
rect 455 1190 461 1191
rect 503 1195 509 1196
rect 503 1191 504 1195
rect 508 1194 509 1195
rect 511 1195 517 1196
rect 511 1194 512 1195
rect 508 1192 512 1194
rect 508 1191 509 1192
rect 503 1190 509 1191
rect 511 1191 512 1192
rect 516 1191 517 1195
rect 511 1190 517 1191
rect 559 1195 565 1196
rect 559 1191 560 1195
rect 564 1194 565 1195
rect 567 1195 573 1196
rect 567 1194 568 1195
rect 564 1192 568 1194
rect 564 1191 565 1192
rect 559 1190 565 1191
rect 567 1191 568 1192
rect 572 1191 573 1195
rect 567 1190 573 1191
rect 615 1195 621 1196
rect 615 1191 616 1195
rect 620 1194 621 1195
rect 623 1195 629 1196
rect 623 1194 624 1195
rect 620 1192 624 1194
rect 620 1191 621 1192
rect 615 1190 621 1191
rect 623 1191 624 1192
rect 628 1191 629 1195
rect 623 1190 629 1191
rect 671 1195 677 1196
rect 671 1191 672 1195
rect 676 1194 677 1195
rect 679 1195 685 1196
rect 679 1194 680 1195
rect 676 1192 680 1194
rect 676 1191 677 1192
rect 671 1190 677 1191
rect 679 1191 680 1192
rect 684 1191 685 1195
rect 679 1190 685 1191
rect 727 1195 733 1196
rect 727 1191 728 1195
rect 732 1191 733 1195
rect 727 1190 733 1191
rect 783 1195 789 1196
rect 783 1191 784 1195
rect 788 1194 789 1195
rect 791 1195 797 1196
rect 791 1194 792 1195
rect 788 1192 792 1194
rect 788 1191 789 1192
rect 783 1190 789 1191
rect 791 1191 792 1192
rect 796 1191 797 1195
rect 791 1190 797 1191
rect 839 1195 845 1196
rect 839 1191 840 1195
rect 844 1194 845 1195
rect 847 1195 853 1196
rect 847 1194 848 1195
rect 844 1192 848 1194
rect 844 1191 845 1192
rect 839 1190 845 1191
rect 847 1191 848 1192
rect 852 1191 853 1195
rect 847 1190 853 1191
rect 903 1195 912 1196
rect 903 1191 904 1195
rect 911 1191 912 1195
rect 967 1195 973 1196
rect 967 1194 968 1195
rect 903 1190 912 1191
rect 960 1192 968 1194
rect 110 1186 116 1187
rect 134 1189 140 1190
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 166 1189 172 1190
rect 166 1185 167 1189
rect 171 1185 172 1189
rect 166 1184 172 1185
rect 222 1189 228 1190
rect 222 1185 223 1189
rect 227 1185 228 1189
rect 222 1184 228 1185
rect 278 1189 284 1190
rect 278 1185 279 1189
rect 283 1185 284 1189
rect 278 1184 284 1185
rect 334 1189 340 1190
rect 334 1185 335 1189
rect 339 1185 340 1189
rect 334 1184 340 1185
rect 382 1189 388 1190
rect 382 1185 383 1189
rect 387 1185 388 1189
rect 382 1184 388 1185
rect 430 1189 436 1190
rect 430 1185 431 1189
rect 435 1185 436 1189
rect 430 1184 436 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 542 1189 548 1190
rect 542 1185 543 1189
rect 547 1185 548 1189
rect 542 1184 548 1185
rect 598 1189 604 1190
rect 598 1185 599 1189
rect 603 1185 604 1189
rect 598 1184 604 1185
rect 654 1189 660 1190
rect 654 1185 655 1189
rect 659 1185 660 1189
rect 654 1184 660 1185
rect 710 1189 716 1190
rect 710 1185 711 1189
rect 715 1185 716 1189
rect 710 1184 716 1185
rect 494 1183 500 1184
rect 494 1179 495 1183
rect 499 1182 500 1183
rect 729 1182 731 1190
rect 766 1189 772 1190
rect 766 1185 767 1189
rect 771 1185 772 1189
rect 822 1189 828 1190
rect 766 1184 772 1185
rect 782 1187 788 1188
rect 782 1183 783 1187
rect 787 1183 788 1187
rect 822 1185 823 1189
rect 827 1185 828 1189
rect 822 1184 828 1185
rect 886 1189 892 1190
rect 886 1185 887 1189
rect 891 1185 892 1189
rect 886 1184 892 1185
rect 950 1189 956 1190
rect 950 1185 951 1189
rect 955 1185 956 1189
rect 950 1184 956 1185
rect 782 1182 788 1183
rect 960 1182 962 1192
rect 967 1191 968 1192
rect 972 1191 973 1195
rect 967 1190 973 1191
rect 1031 1195 1037 1196
rect 1031 1191 1032 1195
rect 1036 1194 1037 1195
rect 1039 1195 1045 1196
rect 1039 1194 1040 1195
rect 1036 1192 1040 1194
rect 1036 1191 1037 1192
rect 1031 1190 1037 1191
rect 1039 1191 1040 1192
rect 1044 1191 1045 1195
rect 1095 1195 1101 1196
rect 1095 1194 1096 1195
rect 1039 1190 1045 1191
rect 1088 1192 1096 1194
rect 1014 1189 1020 1190
rect 1014 1185 1015 1189
rect 1019 1185 1020 1189
rect 1014 1184 1020 1185
rect 1078 1189 1084 1190
rect 1078 1185 1079 1189
rect 1083 1185 1084 1189
rect 1078 1184 1084 1185
rect 499 1180 731 1182
rect 784 1180 962 1182
rect 1006 1183 1012 1184
rect 499 1179 500 1180
rect 494 1178 500 1179
rect 1006 1179 1007 1183
rect 1011 1182 1012 1183
rect 1088 1182 1090 1192
rect 1095 1191 1096 1192
rect 1100 1191 1101 1195
rect 1095 1190 1101 1191
rect 1159 1195 1165 1196
rect 1159 1191 1160 1195
rect 1164 1194 1165 1195
rect 1167 1195 1173 1196
rect 1167 1194 1168 1195
rect 1164 1192 1168 1194
rect 1164 1191 1165 1192
rect 1159 1190 1165 1191
rect 1167 1191 1168 1192
rect 1172 1191 1173 1195
rect 1167 1190 1173 1191
rect 1223 1195 1229 1196
rect 1223 1191 1224 1195
rect 1228 1194 1229 1195
rect 1231 1195 1237 1196
rect 1231 1194 1232 1195
rect 1228 1192 1232 1194
rect 1228 1191 1229 1192
rect 1223 1190 1229 1191
rect 1231 1191 1232 1192
rect 1236 1191 1237 1195
rect 1231 1190 1237 1191
rect 1295 1195 1301 1196
rect 1295 1191 1296 1195
rect 1300 1194 1301 1195
rect 1303 1195 1309 1196
rect 1303 1194 1304 1195
rect 1300 1192 1304 1194
rect 1300 1191 1301 1192
rect 1295 1190 1301 1191
rect 1303 1191 1304 1192
rect 1308 1191 1309 1195
rect 1303 1190 1309 1191
rect 1375 1195 1381 1196
rect 1375 1191 1376 1195
rect 1380 1194 1381 1195
rect 1383 1195 1389 1196
rect 1383 1194 1384 1195
rect 1380 1192 1384 1194
rect 1380 1191 1381 1192
rect 1375 1190 1381 1191
rect 1383 1191 1384 1192
rect 1388 1191 1389 1195
rect 1383 1190 1389 1191
rect 1463 1195 1469 1196
rect 1463 1191 1464 1195
rect 1468 1194 1469 1195
rect 1471 1195 1477 1196
rect 1471 1194 1472 1195
rect 1468 1192 1472 1194
rect 1468 1191 1469 1192
rect 1463 1190 1469 1191
rect 1471 1191 1472 1192
rect 1476 1191 1477 1195
rect 1559 1195 1565 1196
rect 1559 1194 1560 1195
rect 1471 1190 1477 1191
rect 1552 1192 1560 1194
rect 1142 1189 1148 1190
rect 1142 1185 1143 1189
rect 1147 1185 1148 1189
rect 1142 1184 1148 1185
rect 1206 1189 1212 1190
rect 1206 1185 1207 1189
rect 1211 1185 1212 1189
rect 1206 1184 1212 1185
rect 1278 1189 1284 1190
rect 1278 1185 1279 1189
rect 1283 1185 1284 1189
rect 1278 1184 1284 1185
rect 1358 1189 1364 1190
rect 1358 1185 1359 1189
rect 1363 1185 1364 1189
rect 1358 1184 1364 1185
rect 1446 1189 1452 1190
rect 1446 1185 1447 1189
rect 1451 1185 1452 1189
rect 1446 1184 1452 1185
rect 1542 1189 1548 1190
rect 1542 1185 1543 1189
rect 1547 1185 1548 1189
rect 1542 1184 1548 1185
rect 1011 1180 1090 1182
rect 1234 1183 1240 1184
rect 1011 1179 1012 1180
rect 1006 1178 1012 1179
rect 1234 1179 1235 1183
rect 1239 1182 1240 1183
rect 1552 1182 1554 1192
rect 1559 1191 1560 1192
rect 1564 1191 1565 1195
rect 1559 1190 1565 1191
rect 1638 1195 1645 1196
rect 1638 1191 1639 1195
rect 1644 1191 1645 1195
rect 1638 1190 1645 1191
rect 1662 1191 1668 1192
rect 1622 1189 1628 1190
rect 1622 1185 1623 1189
rect 1627 1185 1628 1189
rect 1662 1187 1663 1191
rect 1667 1187 1668 1191
rect 1662 1186 1668 1187
rect 1622 1184 1628 1185
rect 1239 1180 1554 1182
rect 1239 1179 1240 1180
rect 1234 1178 1240 1179
rect 860 1176 978 1178
rect 858 1175 864 1176
rect 134 1171 140 1172
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 134 1167 135 1171
rect 139 1167 140 1171
rect 134 1166 140 1167
rect 166 1171 172 1172
rect 166 1167 167 1171
rect 171 1167 172 1171
rect 166 1166 172 1167
rect 222 1171 228 1172
rect 222 1167 223 1171
rect 227 1167 228 1171
rect 222 1166 228 1167
rect 286 1171 292 1172
rect 286 1167 287 1171
rect 291 1167 292 1171
rect 286 1166 292 1167
rect 350 1171 356 1172
rect 350 1167 351 1171
rect 355 1167 356 1171
rect 350 1166 356 1167
rect 414 1171 420 1172
rect 414 1167 415 1171
rect 419 1167 420 1171
rect 414 1166 420 1167
rect 470 1171 476 1172
rect 470 1167 471 1171
rect 475 1167 476 1171
rect 470 1166 476 1167
rect 534 1171 540 1172
rect 534 1167 535 1171
rect 539 1167 540 1171
rect 534 1166 540 1167
rect 598 1171 604 1172
rect 598 1167 599 1171
rect 603 1167 604 1171
rect 598 1166 604 1167
rect 662 1171 668 1172
rect 662 1167 663 1171
rect 667 1167 668 1171
rect 662 1166 668 1167
rect 726 1171 732 1172
rect 726 1167 727 1171
rect 731 1167 732 1171
rect 726 1166 732 1167
rect 782 1171 788 1172
rect 782 1167 783 1171
rect 787 1167 788 1171
rect 782 1166 788 1167
rect 838 1171 844 1172
rect 838 1167 839 1171
rect 843 1167 844 1171
rect 858 1171 859 1175
rect 863 1171 864 1175
rect 976 1174 978 1176
rect 1016 1176 1179 1178
rect 1016 1174 1018 1176
rect 976 1172 1018 1174
rect 858 1170 864 1171
rect 902 1171 908 1172
rect 838 1166 844 1167
rect 902 1167 903 1171
rect 907 1167 908 1171
rect 902 1166 908 1167
rect 966 1171 972 1172
rect 966 1167 967 1171
rect 971 1167 972 1171
rect 966 1166 972 1167
rect 1030 1171 1036 1172
rect 1030 1167 1031 1171
rect 1035 1167 1036 1171
rect 1030 1166 1036 1167
rect 1094 1171 1100 1172
rect 1094 1167 1095 1171
rect 1099 1167 1100 1171
rect 1094 1166 1100 1167
rect 1158 1171 1164 1172
rect 1158 1167 1159 1171
rect 1163 1167 1164 1171
rect 1158 1166 1164 1167
rect 110 1164 116 1165
rect 1177 1164 1179 1176
rect 1214 1171 1220 1172
rect 1214 1167 1215 1171
rect 1219 1167 1220 1171
rect 1214 1166 1220 1167
rect 1278 1171 1284 1172
rect 1278 1167 1279 1171
rect 1283 1167 1284 1171
rect 1278 1166 1284 1167
rect 1342 1171 1348 1172
rect 1342 1167 1343 1171
rect 1347 1167 1348 1171
rect 1342 1166 1348 1167
rect 1406 1171 1412 1172
rect 1406 1167 1407 1171
rect 1411 1167 1412 1171
rect 1406 1166 1412 1167
rect 1478 1171 1484 1172
rect 1478 1167 1479 1171
rect 1483 1167 1484 1171
rect 1478 1166 1484 1167
rect 1558 1171 1564 1172
rect 1558 1167 1559 1171
rect 1563 1167 1564 1171
rect 1558 1166 1564 1167
rect 1622 1171 1628 1172
rect 1622 1167 1623 1171
rect 1627 1167 1628 1171
rect 1622 1166 1628 1167
rect 1662 1169 1668 1170
rect 1662 1165 1663 1169
rect 1667 1165 1668 1169
rect 1662 1164 1668 1165
rect 151 1163 160 1164
rect 151 1159 152 1163
rect 159 1159 160 1163
rect 183 1163 189 1164
rect 183 1162 184 1163
rect 151 1158 160 1159
rect 176 1160 184 1162
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 134 1150 135 1154
rect 139 1150 140 1154
rect 134 1149 140 1150
rect 166 1154 172 1155
rect 166 1150 167 1154
rect 171 1150 172 1154
rect 166 1149 172 1150
rect 110 1147 116 1148
rect 151 1147 157 1148
rect 151 1143 152 1147
rect 156 1146 157 1147
rect 176 1146 178 1160
rect 183 1159 184 1160
rect 188 1159 189 1163
rect 239 1163 245 1164
rect 239 1162 240 1163
rect 183 1158 189 1159
rect 212 1160 240 1162
rect 156 1144 178 1146
rect 183 1147 189 1148
rect 156 1143 157 1144
rect 151 1142 157 1143
rect 183 1143 184 1147
rect 188 1146 189 1147
rect 212 1146 214 1160
rect 239 1159 240 1160
rect 244 1159 245 1163
rect 239 1158 245 1159
rect 298 1163 309 1164
rect 298 1159 299 1163
rect 303 1159 304 1163
rect 308 1159 309 1163
rect 367 1163 373 1164
rect 367 1162 368 1163
rect 298 1158 309 1159
rect 340 1160 368 1162
rect 222 1154 228 1155
rect 222 1150 223 1154
rect 227 1150 228 1154
rect 222 1149 228 1150
rect 286 1154 292 1155
rect 286 1150 287 1154
rect 291 1150 292 1154
rect 286 1149 292 1150
rect 188 1144 214 1146
rect 238 1147 245 1148
rect 188 1143 189 1144
rect 183 1142 189 1143
rect 238 1143 239 1147
rect 244 1143 245 1147
rect 238 1142 245 1143
rect 303 1147 309 1148
rect 303 1143 304 1147
rect 308 1146 309 1147
rect 340 1146 342 1160
rect 367 1159 368 1160
rect 372 1159 373 1163
rect 431 1163 437 1164
rect 431 1162 432 1163
rect 367 1158 373 1159
rect 404 1160 432 1162
rect 350 1154 356 1155
rect 350 1150 351 1154
rect 355 1150 356 1154
rect 350 1149 356 1150
rect 308 1144 342 1146
rect 367 1147 373 1148
rect 308 1143 309 1144
rect 303 1142 309 1143
rect 367 1143 368 1147
rect 372 1146 373 1147
rect 404 1146 406 1160
rect 431 1159 432 1160
rect 436 1159 437 1163
rect 431 1158 437 1159
rect 487 1163 493 1164
rect 487 1159 488 1163
rect 492 1159 493 1163
rect 487 1158 493 1159
rect 551 1163 557 1164
rect 551 1159 552 1163
rect 556 1159 557 1163
rect 551 1158 557 1159
rect 615 1163 621 1164
rect 615 1159 616 1163
rect 620 1159 621 1163
rect 615 1158 621 1159
rect 679 1163 685 1164
rect 679 1159 680 1163
rect 684 1159 685 1163
rect 679 1158 685 1159
rect 743 1163 749 1164
rect 743 1159 744 1163
rect 748 1162 749 1163
rect 798 1163 805 1164
rect 748 1160 774 1162
rect 748 1159 749 1160
rect 743 1158 749 1159
rect 414 1154 420 1155
rect 414 1150 415 1154
rect 419 1150 420 1154
rect 414 1149 420 1150
rect 470 1154 476 1155
rect 470 1150 471 1154
rect 475 1150 476 1154
rect 489 1154 491 1158
rect 553 1156 586 1158
rect 617 1156 650 1158
rect 681 1156 714 1158
rect 534 1154 540 1155
rect 489 1152 522 1154
rect 470 1149 476 1150
rect 372 1144 406 1146
rect 431 1147 437 1148
rect 372 1143 373 1144
rect 367 1142 373 1143
rect 431 1143 432 1147
rect 436 1146 437 1147
rect 478 1147 484 1148
rect 478 1146 479 1147
rect 436 1144 479 1146
rect 436 1143 437 1144
rect 431 1142 437 1143
rect 478 1143 479 1144
rect 483 1143 484 1147
rect 478 1142 484 1143
rect 487 1147 493 1148
rect 487 1143 488 1147
rect 492 1143 493 1147
rect 520 1146 522 1152
rect 534 1150 535 1154
rect 539 1150 540 1154
rect 534 1149 540 1150
rect 551 1147 557 1148
rect 551 1146 552 1147
rect 520 1144 552 1146
rect 487 1142 493 1143
rect 551 1143 552 1144
rect 556 1143 557 1147
rect 584 1146 586 1156
rect 598 1154 604 1155
rect 598 1150 599 1154
rect 603 1150 604 1154
rect 598 1149 604 1150
rect 615 1147 621 1148
rect 615 1146 616 1147
rect 584 1144 616 1146
rect 551 1142 557 1143
rect 615 1143 616 1144
rect 620 1143 621 1147
rect 648 1146 650 1156
rect 662 1154 668 1155
rect 662 1150 663 1154
rect 667 1150 668 1154
rect 662 1149 668 1150
rect 679 1147 685 1148
rect 679 1146 680 1147
rect 648 1144 680 1146
rect 615 1142 621 1143
rect 679 1143 680 1144
rect 684 1143 685 1147
rect 712 1146 714 1156
rect 726 1154 732 1155
rect 726 1150 727 1154
rect 731 1150 732 1154
rect 726 1149 732 1150
rect 743 1147 749 1148
rect 743 1146 744 1147
rect 712 1144 744 1146
rect 679 1142 685 1143
rect 743 1143 744 1144
rect 748 1143 749 1147
rect 772 1146 774 1160
rect 798 1159 799 1163
rect 804 1159 805 1163
rect 798 1158 805 1159
rect 855 1163 861 1164
rect 855 1159 856 1163
rect 860 1159 861 1163
rect 855 1158 861 1159
rect 919 1163 925 1164
rect 919 1159 920 1163
rect 924 1159 925 1163
rect 919 1158 925 1159
rect 983 1163 989 1164
rect 983 1159 984 1163
rect 988 1162 989 1163
rect 1022 1163 1028 1164
rect 1022 1162 1023 1163
rect 988 1160 1023 1162
rect 988 1159 989 1160
rect 983 1158 989 1159
rect 1022 1159 1023 1160
rect 1027 1159 1028 1163
rect 1022 1158 1028 1159
rect 1047 1163 1053 1164
rect 1047 1159 1048 1163
rect 1052 1159 1053 1163
rect 1047 1158 1053 1159
rect 1111 1163 1117 1164
rect 1111 1159 1112 1163
rect 1116 1162 1117 1163
rect 1175 1163 1181 1164
rect 1116 1160 1170 1162
rect 1116 1159 1117 1160
rect 1111 1158 1117 1159
rect 782 1154 788 1155
rect 782 1150 783 1154
rect 787 1150 788 1154
rect 782 1149 788 1150
rect 838 1154 844 1155
rect 838 1150 839 1154
rect 843 1150 844 1154
rect 857 1154 859 1158
rect 921 1156 954 1158
rect 1049 1156 1082 1158
rect 902 1154 908 1155
rect 857 1152 890 1154
rect 838 1149 844 1150
rect 799 1147 805 1148
rect 799 1146 800 1147
rect 772 1144 800 1146
rect 743 1142 749 1143
rect 799 1143 800 1144
rect 804 1143 805 1147
rect 799 1142 805 1143
rect 855 1147 864 1148
rect 855 1143 856 1147
rect 863 1143 864 1147
rect 888 1146 890 1152
rect 902 1150 903 1154
rect 907 1150 908 1154
rect 902 1149 908 1150
rect 919 1147 925 1148
rect 919 1146 920 1147
rect 888 1144 920 1146
rect 855 1142 864 1143
rect 919 1143 920 1144
rect 924 1143 925 1147
rect 952 1146 954 1156
rect 966 1154 972 1155
rect 966 1150 967 1154
rect 971 1150 972 1154
rect 966 1149 972 1150
rect 1030 1154 1036 1155
rect 1030 1150 1031 1154
rect 1035 1150 1036 1154
rect 1030 1149 1036 1150
rect 983 1147 989 1148
rect 983 1146 984 1147
rect 952 1144 984 1146
rect 919 1142 925 1143
rect 983 1143 984 1144
rect 988 1143 989 1147
rect 983 1142 989 1143
rect 1042 1147 1053 1148
rect 1042 1143 1043 1147
rect 1047 1143 1048 1147
rect 1052 1143 1053 1147
rect 1080 1146 1082 1156
rect 1094 1154 1100 1155
rect 1094 1150 1095 1154
rect 1099 1150 1100 1154
rect 1094 1149 1100 1150
rect 1158 1154 1164 1155
rect 1158 1150 1159 1154
rect 1163 1150 1164 1154
rect 1158 1149 1164 1150
rect 1111 1147 1117 1148
rect 1111 1146 1112 1147
rect 1080 1144 1112 1146
rect 1042 1142 1053 1143
rect 1111 1143 1112 1144
rect 1116 1143 1117 1147
rect 1168 1146 1170 1160
rect 1175 1159 1176 1163
rect 1180 1159 1181 1163
rect 1175 1158 1181 1159
rect 1231 1163 1237 1164
rect 1231 1159 1232 1163
rect 1236 1162 1237 1163
rect 1295 1163 1301 1164
rect 1236 1160 1290 1162
rect 1236 1159 1237 1160
rect 1231 1158 1237 1159
rect 1214 1154 1220 1155
rect 1214 1150 1215 1154
rect 1219 1150 1220 1154
rect 1214 1149 1220 1150
rect 1278 1154 1284 1155
rect 1278 1150 1279 1154
rect 1283 1150 1284 1154
rect 1278 1149 1284 1150
rect 1175 1147 1181 1148
rect 1175 1146 1176 1147
rect 1168 1144 1176 1146
rect 1111 1142 1117 1143
rect 1175 1143 1176 1144
rect 1180 1143 1181 1147
rect 1175 1142 1181 1143
rect 1231 1147 1240 1148
rect 1231 1143 1232 1147
rect 1239 1143 1240 1147
rect 1288 1146 1290 1160
rect 1295 1159 1296 1163
rect 1300 1159 1301 1163
rect 1295 1158 1301 1159
rect 1359 1163 1365 1164
rect 1359 1159 1360 1163
rect 1364 1159 1365 1163
rect 1359 1158 1365 1159
rect 1423 1163 1429 1164
rect 1423 1159 1424 1163
rect 1428 1162 1429 1163
rect 1495 1163 1501 1164
rect 1428 1160 1490 1162
rect 1428 1159 1429 1160
rect 1423 1158 1429 1159
rect 1297 1156 1330 1158
rect 1295 1147 1301 1148
rect 1295 1146 1296 1147
rect 1288 1144 1296 1146
rect 1231 1142 1240 1143
rect 1295 1143 1296 1144
rect 1300 1143 1301 1147
rect 1328 1146 1330 1156
rect 1342 1154 1348 1155
rect 1342 1150 1343 1154
rect 1347 1150 1348 1154
rect 1361 1154 1363 1158
rect 1406 1154 1412 1155
rect 1361 1152 1394 1154
rect 1342 1149 1348 1150
rect 1359 1147 1365 1148
rect 1359 1146 1360 1147
rect 1328 1144 1360 1146
rect 1295 1142 1301 1143
rect 1359 1143 1360 1144
rect 1364 1143 1365 1147
rect 1392 1146 1394 1152
rect 1406 1150 1407 1154
rect 1411 1150 1412 1154
rect 1406 1149 1412 1150
rect 1478 1154 1484 1155
rect 1478 1150 1479 1154
rect 1483 1150 1484 1154
rect 1478 1149 1484 1150
rect 1423 1147 1429 1148
rect 1423 1146 1424 1147
rect 1392 1144 1424 1146
rect 1359 1142 1365 1143
rect 1423 1143 1424 1144
rect 1428 1143 1429 1147
rect 1488 1146 1490 1160
rect 1495 1159 1496 1163
rect 1500 1159 1501 1163
rect 1495 1158 1501 1159
rect 1543 1163 1549 1164
rect 1543 1159 1544 1163
rect 1548 1162 1549 1163
rect 1575 1163 1581 1164
rect 1575 1162 1576 1163
rect 1548 1160 1576 1162
rect 1548 1159 1549 1160
rect 1543 1158 1549 1159
rect 1575 1159 1576 1160
rect 1580 1159 1581 1163
rect 1575 1158 1581 1159
rect 1639 1163 1645 1164
rect 1639 1159 1640 1163
rect 1644 1162 1645 1163
rect 1647 1163 1653 1164
rect 1647 1162 1648 1163
rect 1644 1160 1648 1162
rect 1644 1159 1645 1160
rect 1639 1158 1645 1159
rect 1647 1159 1648 1160
rect 1652 1159 1653 1163
rect 1647 1158 1653 1159
rect 1497 1154 1499 1158
rect 1558 1154 1564 1155
rect 1497 1152 1538 1154
rect 1495 1147 1501 1148
rect 1495 1146 1496 1147
rect 1488 1144 1496 1146
rect 1423 1142 1429 1143
rect 1495 1143 1496 1144
rect 1500 1143 1501 1147
rect 1536 1146 1538 1152
rect 1558 1150 1559 1154
rect 1563 1150 1564 1154
rect 1558 1149 1564 1150
rect 1622 1154 1628 1155
rect 1622 1150 1623 1154
rect 1627 1150 1628 1154
rect 1622 1149 1628 1150
rect 1662 1152 1668 1153
rect 1662 1148 1663 1152
rect 1667 1148 1668 1152
rect 1575 1147 1581 1148
rect 1575 1146 1576 1147
rect 1536 1144 1576 1146
rect 1495 1142 1501 1143
rect 1575 1143 1576 1144
rect 1580 1143 1581 1147
rect 1575 1142 1581 1143
rect 1638 1147 1645 1148
rect 1662 1147 1668 1148
rect 1638 1143 1639 1147
rect 1644 1143 1645 1147
rect 1638 1142 1645 1143
rect 798 1135 804 1136
rect 798 1134 799 1135
rect 544 1132 799 1134
rect 199 1127 205 1128
rect 154 1123 165 1124
rect 110 1120 116 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 154 1119 155 1123
rect 159 1119 160 1123
rect 164 1119 165 1123
rect 191 1123 197 1124
rect 191 1122 192 1123
rect 184 1120 192 1122
rect 110 1115 116 1116
rect 142 1118 148 1119
rect 154 1118 165 1119
rect 174 1118 180 1119
rect 142 1114 143 1118
rect 147 1114 148 1118
rect 142 1113 148 1114
rect 174 1114 175 1118
rect 179 1114 180 1118
rect 174 1113 180 1114
rect 184 1108 186 1120
rect 191 1119 192 1120
rect 196 1119 197 1123
rect 199 1123 200 1127
rect 204 1126 205 1127
rect 239 1127 245 1128
rect 204 1124 226 1126
rect 204 1123 205 1124
rect 199 1122 205 1123
rect 224 1122 226 1124
rect 231 1123 237 1124
rect 231 1122 232 1123
rect 224 1120 232 1122
rect 231 1119 232 1120
rect 236 1119 237 1123
rect 239 1123 240 1127
rect 244 1126 245 1127
rect 298 1127 304 1128
rect 244 1124 282 1126
rect 244 1123 245 1124
rect 239 1122 245 1123
rect 280 1122 282 1124
rect 287 1123 293 1124
rect 287 1122 288 1123
rect 280 1120 288 1122
rect 287 1119 288 1120
rect 292 1119 293 1123
rect 298 1123 299 1127
rect 303 1126 304 1127
rect 359 1127 365 1128
rect 303 1124 346 1126
rect 303 1123 304 1124
rect 298 1122 304 1123
rect 344 1122 346 1124
rect 351 1123 357 1124
rect 351 1122 352 1123
rect 344 1120 352 1122
rect 351 1119 352 1120
rect 356 1119 357 1123
rect 359 1123 360 1127
rect 364 1126 365 1127
rect 423 1127 429 1128
rect 364 1124 410 1126
rect 364 1123 365 1124
rect 359 1122 365 1123
rect 408 1122 410 1124
rect 415 1123 421 1124
rect 415 1122 416 1123
rect 408 1120 416 1122
rect 415 1119 416 1120
rect 420 1119 421 1123
rect 423 1123 424 1127
rect 428 1126 429 1127
rect 428 1124 474 1126
rect 544 1124 546 1132
rect 798 1131 799 1132
rect 803 1131 804 1135
rect 1102 1135 1108 1136
rect 1102 1134 1103 1135
rect 798 1130 804 1131
rect 928 1132 1103 1134
rect 551 1127 557 1128
rect 428 1123 429 1124
rect 423 1122 429 1123
rect 472 1122 474 1124
rect 479 1123 485 1124
rect 479 1122 480 1123
rect 472 1120 480 1122
rect 479 1119 480 1120
rect 484 1119 485 1123
rect 543 1123 549 1124
rect 543 1119 544 1123
rect 548 1119 549 1123
rect 551 1123 552 1127
rect 556 1126 557 1127
rect 623 1127 629 1128
rect 556 1124 619 1126
rect 556 1123 557 1124
rect 551 1122 557 1123
rect 615 1123 621 1124
rect 615 1119 616 1123
rect 620 1119 621 1123
rect 623 1123 624 1127
rect 628 1126 629 1127
rect 687 1127 693 1128
rect 628 1124 683 1126
rect 628 1123 629 1124
rect 623 1122 629 1123
rect 679 1123 685 1124
rect 679 1119 680 1123
rect 684 1119 685 1123
rect 687 1123 688 1127
rect 692 1126 693 1127
rect 751 1127 757 1128
rect 692 1124 747 1126
rect 692 1123 693 1124
rect 687 1122 693 1123
rect 743 1123 749 1124
rect 743 1119 744 1123
rect 748 1119 749 1123
rect 751 1123 752 1127
rect 756 1126 757 1127
rect 815 1127 821 1128
rect 756 1124 802 1126
rect 756 1123 757 1124
rect 751 1122 757 1123
rect 800 1122 802 1124
rect 807 1123 813 1124
rect 807 1122 808 1123
rect 800 1120 808 1122
rect 807 1119 808 1120
rect 812 1119 813 1123
rect 815 1123 816 1127
rect 820 1126 821 1127
rect 820 1124 866 1126
rect 928 1124 930 1132
rect 1102 1131 1103 1132
rect 1107 1131 1108 1135
rect 1543 1135 1549 1136
rect 1543 1134 1544 1135
rect 1102 1130 1108 1131
rect 1353 1132 1544 1134
rect 935 1127 941 1128
rect 820 1123 821 1124
rect 815 1122 821 1123
rect 864 1122 866 1124
rect 871 1123 877 1124
rect 871 1122 872 1123
rect 864 1120 872 1122
rect 871 1119 872 1120
rect 876 1119 877 1123
rect 927 1123 933 1124
rect 927 1119 928 1123
rect 932 1119 933 1123
rect 935 1123 936 1127
rect 940 1126 941 1127
rect 991 1127 997 1128
rect 940 1124 987 1126
rect 940 1123 941 1124
rect 935 1122 941 1123
rect 983 1123 989 1124
rect 983 1119 984 1123
rect 988 1119 989 1123
rect 991 1123 992 1127
rect 996 1126 997 1127
rect 1175 1127 1181 1128
rect 996 1124 1034 1126
rect 996 1123 997 1124
rect 991 1122 997 1123
rect 1032 1122 1034 1124
rect 1039 1123 1045 1124
rect 1039 1122 1040 1123
rect 1032 1120 1040 1122
rect 1039 1119 1040 1120
rect 1044 1119 1045 1123
rect 1103 1123 1109 1124
rect 1103 1119 1104 1123
rect 1108 1122 1109 1123
rect 1130 1123 1136 1124
rect 1130 1122 1131 1123
rect 1108 1120 1131 1122
rect 1108 1119 1109 1120
rect 191 1118 197 1119
rect 214 1118 220 1119
rect 231 1118 237 1119
rect 270 1118 276 1119
rect 287 1118 293 1119
rect 334 1118 340 1119
rect 351 1118 357 1119
rect 398 1118 404 1119
rect 415 1118 421 1119
rect 462 1118 468 1119
rect 479 1118 485 1119
rect 526 1118 532 1119
rect 543 1118 549 1119
rect 598 1118 604 1119
rect 615 1118 621 1119
rect 662 1118 668 1119
rect 679 1118 685 1119
rect 726 1118 732 1119
rect 743 1118 749 1119
rect 790 1118 796 1119
rect 807 1118 813 1119
rect 854 1118 860 1119
rect 871 1118 877 1119
rect 910 1118 916 1119
rect 927 1118 933 1119
rect 966 1118 972 1119
rect 983 1118 989 1119
rect 1022 1118 1028 1119
rect 1039 1118 1045 1119
rect 1086 1118 1092 1119
rect 1103 1118 1109 1119
rect 1130 1119 1131 1120
rect 1135 1119 1136 1123
rect 1162 1123 1173 1124
rect 1162 1119 1163 1123
rect 1167 1119 1168 1123
rect 1172 1119 1173 1123
rect 1175 1123 1176 1127
rect 1180 1126 1181 1127
rect 1239 1127 1245 1128
rect 1180 1124 1235 1126
rect 1180 1123 1181 1124
rect 1175 1122 1181 1123
rect 1231 1123 1237 1124
rect 1231 1119 1232 1123
rect 1236 1119 1237 1123
rect 1239 1123 1240 1127
rect 1244 1126 1245 1127
rect 1244 1124 1299 1126
rect 1353 1124 1355 1132
rect 1543 1131 1544 1132
rect 1548 1131 1549 1135
rect 1543 1130 1549 1131
rect 1359 1127 1365 1128
rect 1244 1123 1245 1124
rect 1239 1122 1245 1123
rect 1295 1123 1301 1124
rect 1295 1119 1296 1123
rect 1300 1119 1301 1123
rect 1351 1123 1357 1124
rect 1351 1119 1352 1123
rect 1356 1119 1357 1123
rect 1359 1123 1360 1127
rect 1364 1126 1365 1127
rect 1415 1127 1421 1128
rect 1364 1124 1411 1126
rect 1364 1123 1365 1124
rect 1359 1122 1365 1123
rect 1407 1123 1413 1124
rect 1407 1119 1408 1123
rect 1412 1119 1413 1123
rect 1415 1123 1416 1127
rect 1420 1126 1421 1127
rect 1471 1127 1477 1128
rect 1420 1124 1467 1126
rect 1420 1123 1421 1124
rect 1415 1122 1421 1123
rect 1463 1123 1469 1124
rect 1463 1119 1464 1123
rect 1468 1119 1469 1123
rect 1471 1123 1472 1127
rect 1476 1126 1477 1127
rect 1567 1127 1573 1128
rect 1476 1124 1515 1126
rect 1476 1123 1477 1124
rect 1471 1122 1477 1123
rect 1511 1123 1517 1124
rect 1511 1119 1512 1123
rect 1516 1119 1517 1123
rect 1558 1123 1565 1124
rect 1558 1119 1559 1123
rect 1564 1119 1565 1123
rect 1567 1123 1568 1127
rect 1572 1126 1573 1127
rect 1572 1124 1611 1126
rect 1616 1124 1643 1126
rect 1572 1123 1573 1124
rect 1567 1122 1573 1123
rect 1607 1123 1613 1124
rect 1607 1119 1608 1123
rect 1612 1119 1613 1123
rect 1130 1118 1136 1119
rect 1150 1118 1156 1119
rect 1162 1118 1173 1119
rect 1214 1118 1220 1119
rect 1231 1118 1237 1119
rect 1278 1118 1284 1119
rect 1295 1118 1301 1119
rect 1334 1118 1340 1119
rect 1351 1118 1357 1119
rect 1390 1118 1396 1119
rect 1407 1118 1413 1119
rect 1446 1118 1452 1119
rect 1463 1118 1469 1119
rect 1494 1118 1500 1119
rect 1511 1118 1517 1119
rect 1542 1118 1548 1119
rect 1558 1118 1565 1119
rect 1590 1118 1596 1119
rect 1607 1118 1613 1119
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 214 1113 220 1114
rect 270 1114 271 1118
rect 275 1114 276 1118
rect 270 1113 276 1114
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 334 1113 340 1114
rect 398 1114 399 1118
rect 403 1114 404 1118
rect 398 1113 404 1114
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 462 1113 468 1114
rect 526 1114 527 1118
rect 531 1114 532 1118
rect 526 1113 532 1114
rect 598 1114 599 1118
rect 603 1114 604 1118
rect 598 1113 604 1114
rect 662 1114 663 1118
rect 667 1114 668 1118
rect 662 1113 668 1114
rect 726 1114 727 1118
rect 731 1114 732 1118
rect 726 1113 732 1114
rect 790 1114 791 1118
rect 795 1114 796 1118
rect 790 1113 796 1114
rect 854 1114 855 1118
rect 859 1114 860 1118
rect 854 1113 860 1114
rect 910 1114 911 1118
rect 915 1114 916 1118
rect 910 1113 916 1114
rect 966 1114 967 1118
rect 971 1114 972 1118
rect 966 1113 972 1114
rect 1022 1114 1023 1118
rect 1027 1114 1028 1118
rect 1022 1113 1028 1114
rect 1086 1114 1087 1118
rect 1091 1114 1092 1118
rect 1086 1113 1092 1114
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1150 1113 1156 1114
rect 1214 1114 1215 1118
rect 1219 1114 1220 1118
rect 1214 1113 1220 1114
rect 1278 1114 1279 1118
rect 1283 1114 1284 1118
rect 1278 1113 1284 1114
rect 1334 1114 1335 1118
rect 1339 1114 1340 1118
rect 1334 1113 1340 1114
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1390 1113 1396 1114
rect 1446 1114 1447 1118
rect 1451 1114 1452 1118
rect 1446 1113 1452 1114
rect 1494 1114 1495 1118
rect 1499 1114 1500 1118
rect 1494 1113 1500 1114
rect 1542 1114 1543 1118
rect 1547 1114 1548 1118
rect 1542 1113 1548 1114
rect 1590 1114 1591 1118
rect 1595 1114 1596 1118
rect 1590 1113 1596 1114
rect 159 1107 165 1108
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 159 1103 160 1107
rect 164 1106 165 1107
rect 172 1106 186 1108
rect 191 1107 197 1108
rect 164 1104 174 1106
rect 164 1103 165 1104
rect 159 1102 165 1103
rect 191 1103 192 1107
rect 196 1106 197 1107
rect 199 1107 205 1108
rect 199 1106 200 1107
rect 196 1104 200 1106
rect 196 1103 197 1104
rect 191 1102 197 1103
rect 199 1103 200 1104
rect 204 1103 205 1107
rect 199 1102 205 1103
rect 231 1107 237 1108
rect 231 1103 232 1107
rect 236 1106 237 1107
rect 239 1107 245 1108
rect 239 1106 240 1107
rect 236 1104 240 1106
rect 236 1103 237 1104
rect 231 1102 237 1103
rect 239 1103 240 1104
rect 244 1103 245 1107
rect 287 1107 293 1108
rect 287 1106 288 1107
rect 239 1102 245 1103
rect 280 1104 288 1106
rect 110 1098 116 1099
rect 142 1101 148 1102
rect 142 1097 143 1101
rect 147 1097 148 1101
rect 142 1096 148 1097
rect 174 1101 180 1102
rect 174 1097 175 1101
rect 179 1097 180 1101
rect 174 1096 180 1097
rect 214 1101 220 1102
rect 214 1097 215 1101
rect 219 1097 220 1101
rect 214 1096 220 1097
rect 270 1101 276 1102
rect 270 1097 271 1101
rect 275 1097 276 1101
rect 270 1096 276 1097
rect 234 1095 240 1096
rect 234 1091 235 1095
rect 239 1094 240 1095
rect 280 1094 282 1104
rect 287 1103 288 1104
rect 292 1103 293 1107
rect 287 1102 293 1103
rect 351 1107 357 1108
rect 351 1103 352 1107
rect 356 1106 357 1107
rect 359 1107 365 1108
rect 359 1106 360 1107
rect 356 1104 360 1106
rect 356 1103 357 1104
rect 351 1102 357 1103
rect 359 1103 360 1104
rect 364 1103 365 1107
rect 359 1102 365 1103
rect 415 1107 421 1108
rect 415 1103 416 1107
rect 420 1106 421 1107
rect 423 1107 429 1108
rect 423 1106 424 1107
rect 420 1104 424 1106
rect 420 1103 421 1104
rect 415 1102 421 1103
rect 423 1103 424 1104
rect 428 1103 429 1107
rect 423 1102 429 1103
rect 478 1107 485 1108
rect 478 1103 479 1107
rect 484 1103 485 1107
rect 478 1102 485 1103
rect 543 1107 549 1108
rect 543 1103 544 1107
rect 548 1106 549 1107
rect 551 1107 557 1108
rect 551 1106 552 1107
rect 548 1104 552 1106
rect 548 1103 549 1104
rect 543 1102 549 1103
rect 551 1103 552 1104
rect 556 1103 557 1107
rect 551 1102 557 1103
rect 615 1107 621 1108
rect 615 1103 616 1107
rect 620 1106 621 1107
rect 623 1107 629 1108
rect 623 1106 624 1107
rect 620 1104 624 1106
rect 620 1103 621 1104
rect 615 1102 621 1103
rect 623 1103 624 1104
rect 628 1103 629 1107
rect 623 1102 629 1103
rect 679 1107 685 1108
rect 679 1103 680 1107
rect 684 1106 685 1107
rect 687 1107 693 1108
rect 687 1106 688 1107
rect 684 1104 688 1106
rect 684 1103 685 1104
rect 679 1102 685 1103
rect 687 1103 688 1104
rect 692 1103 693 1107
rect 687 1102 693 1103
rect 743 1107 749 1108
rect 743 1103 744 1107
rect 748 1106 749 1107
rect 751 1107 757 1108
rect 751 1106 752 1107
rect 748 1104 752 1106
rect 748 1103 749 1104
rect 743 1102 749 1103
rect 751 1103 752 1104
rect 756 1103 757 1107
rect 751 1102 757 1103
rect 807 1107 813 1108
rect 807 1103 808 1107
rect 812 1106 813 1107
rect 815 1107 821 1108
rect 815 1106 816 1107
rect 812 1104 816 1106
rect 812 1103 813 1104
rect 807 1102 813 1103
rect 815 1103 816 1104
rect 820 1103 821 1107
rect 815 1102 821 1103
rect 871 1107 877 1108
rect 871 1103 872 1107
rect 876 1106 877 1107
rect 902 1107 908 1108
rect 902 1106 903 1107
rect 876 1104 903 1106
rect 876 1103 877 1104
rect 871 1102 877 1103
rect 902 1103 903 1104
rect 907 1103 908 1107
rect 902 1102 908 1103
rect 927 1107 933 1108
rect 927 1103 928 1107
rect 932 1106 933 1107
rect 935 1107 941 1108
rect 935 1106 936 1107
rect 932 1104 936 1106
rect 932 1103 933 1104
rect 927 1102 933 1103
rect 935 1103 936 1104
rect 940 1103 941 1107
rect 935 1102 941 1103
rect 983 1107 989 1108
rect 983 1103 984 1107
rect 988 1106 989 1107
rect 991 1107 997 1108
rect 991 1106 992 1107
rect 988 1104 992 1106
rect 988 1103 989 1104
rect 983 1102 989 1103
rect 991 1103 992 1104
rect 996 1103 997 1107
rect 991 1102 997 1103
rect 1039 1107 1048 1108
rect 1039 1103 1040 1107
rect 1047 1103 1048 1107
rect 1039 1102 1048 1103
rect 1102 1107 1109 1108
rect 1102 1103 1103 1107
rect 1108 1103 1109 1107
rect 1102 1102 1109 1103
rect 1167 1107 1173 1108
rect 1167 1103 1168 1107
rect 1172 1106 1173 1107
rect 1175 1107 1181 1108
rect 1175 1106 1176 1107
rect 1172 1104 1176 1106
rect 1172 1103 1173 1104
rect 1167 1102 1173 1103
rect 1175 1103 1176 1104
rect 1180 1103 1181 1107
rect 1175 1102 1181 1103
rect 1231 1107 1237 1108
rect 1231 1103 1232 1107
rect 1236 1106 1237 1107
rect 1239 1107 1245 1108
rect 1239 1106 1240 1107
rect 1236 1104 1240 1106
rect 1236 1103 1237 1104
rect 1231 1102 1237 1103
rect 1239 1103 1240 1104
rect 1244 1103 1245 1107
rect 1239 1102 1245 1103
rect 1295 1107 1301 1108
rect 1295 1103 1296 1107
rect 1300 1103 1301 1107
rect 1295 1102 1301 1103
rect 1351 1107 1357 1108
rect 1351 1103 1352 1107
rect 1356 1106 1357 1107
rect 1359 1107 1365 1108
rect 1359 1106 1360 1107
rect 1356 1104 1360 1106
rect 1356 1103 1357 1104
rect 1351 1102 1357 1103
rect 1359 1103 1360 1104
rect 1364 1103 1365 1107
rect 1359 1102 1365 1103
rect 1407 1107 1413 1108
rect 1407 1103 1408 1107
rect 1412 1106 1413 1107
rect 1415 1107 1421 1108
rect 1415 1106 1416 1107
rect 1412 1104 1416 1106
rect 1412 1103 1413 1104
rect 1407 1102 1413 1103
rect 1415 1103 1416 1104
rect 1420 1103 1421 1107
rect 1415 1102 1421 1103
rect 1463 1107 1469 1108
rect 1463 1103 1464 1107
rect 1468 1106 1469 1107
rect 1471 1107 1477 1108
rect 1471 1106 1472 1107
rect 1468 1104 1472 1106
rect 1468 1103 1469 1104
rect 1463 1102 1469 1103
rect 1471 1103 1472 1104
rect 1476 1103 1477 1107
rect 1471 1102 1477 1103
rect 1511 1107 1517 1108
rect 1511 1103 1512 1107
rect 1516 1103 1517 1107
rect 1511 1102 1517 1103
rect 1559 1107 1565 1108
rect 1559 1103 1560 1107
rect 1564 1106 1565 1107
rect 1567 1107 1573 1108
rect 1567 1106 1568 1107
rect 1564 1104 1568 1106
rect 1564 1103 1565 1104
rect 1559 1102 1565 1103
rect 1567 1103 1568 1104
rect 1572 1103 1573 1107
rect 1567 1102 1573 1103
rect 1607 1107 1613 1108
rect 1607 1103 1608 1107
rect 1612 1106 1613 1107
rect 1616 1106 1618 1124
rect 1639 1123 1645 1124
rect 1639 1119 1640 1123
rect 1644 1119 1645 1123
rect 1622 1118 1628 1119
rect 1639 1118 1645 1119
rect 1662 1120 1668 1121
rect 1622 1114 1623 1118
rect 1627 1114 1628 1118
rect 1662 1116 1663 1120
rect 1667 1116 1668 1120
rect 1662 1115 1668 1116
rect 1622 1113 1628 1114
rect 1612 1104 1618 1106
rect 1638 1107 1645 1108
rect 1612 1103 1613 1104
rect 1607 1102 1613 1103
rect 1638 1103 1639 1107
rect 1644 1103 1645 1107
rect 1638 1102 1645 1103
rect 1662 1103 1668 1104
rect 334 1101 340 1102
rect 334 1097 335 1101
rect 339 1097 340 1101
rect 334 1096 340 1097
rect 398 1101 404 1102
rect 398 1097 399 1101
rect 403 1097 404 1101
rect 398 1096 404 1097
rect 462 1101 468 1102
rect 462 1097 463 1101
rect 467 1097 468 1101
rect 462 1096 468 1097
rect 526 1101 532 1102
rect 526 1097 527 1101
rect 531 1097 532 1101
rect 526 1096 532 1097
rect 598 1101 604 1102
rect 598 1097 599 1101
rect 603 1097 604 1101
rect 598 1096 604 1097
rect 662 1101 668 1102
rect 662 1097 663 1101
rect 667 1097 668 1101
rect 662 1096 668 1097
rect 726 1101 732 1102
rect 726 1097 727 1101
rect 731 1097 732 1101
rect 726 1096 732 1097
rect 790 1101 796 1102
rect 790 1097 791 1101
rect 795 1097 796 1101
rect 790 1096 796 1097
rect 854 1101 860 1102
rect 854 1097 855 1101
rect 859 1097 860 1101
rect 854 1096 860 1097
rect 910 1101 916 1102
rect 910 1097 911 1101
rect 915 1097 916 1101
rect 910 1096 916 1097
rect 966 1101 972 1102
rect 966 1097 967 1101
rect 971 1097 972 1101
rect 966 1096 972 1097
rect 1022 1101 1028 1102
rect 1022 1097 1023 1101
rect 1027 1097 1028 1101
rect 1022 1096 1028 1097
rect 1086 1101 1092 1102
rect 1086 1097 1087 1101
rect 1091 1097 1092 1101
rect 1086 1096 1092 1097
rect 1150 1101 1156 1102
rect 1150 1097 1151 1101
rect 1155 1097 1156 1101
rect 1150 1096 1156 1097
rect 1214 1101 1220 1102
rect 1214 1097 1215 1101
rect 1219 1097 1220 1101
rect 1214 1096 1220 1097
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1278 1096 1284 1097
rect 239 1092 282 1094
rect 1130 1095 1136 1096
rect 239 1091 240 1092
rect 234 1090 240 1091
rect 1130 1091 1131 1095
rect 1135 1094 1136 1095
rect 1297 1094 1299 1102
rect 1334 1101 1340 1102
rect 1334 1097 1335 1101
rect 1339 1097 1340 1101
rect 1334 1096 1340 1097
rect 1390 1101 1396 1102
rect 1390 1097 1391 1101
rect 1395 1097 1396 1101
rect 1390 1096 1396 1097
rect 1446 1101 1452 1102
rect 1446 1097 1447 1101
rect 1451 1097 1452 1101
rect 1446 1096 1452 1097
rect 1494 1101 1500 1102
rect 1494 1097 1495 1101
rect 1499 1097 1500 1101
rect 1494 1096 1500 1097
rect 1135 1092 1299 1094
rect 1378 1095 1384 1096
rect 1135 1091 1136 1092
rect 1130 1090 1136 1091
rect 1378 1091 1379 1095
rect 1383 1094 1384 1095
rect 1513 1094 1515 1102
rect 1542 1101 1548 1102
rect 1542 1097 1543 1101
rect 1547 1097 1548 1101
rect 1542 1096 1548 1097
rect 1590 1101 1596 1102
rect 1590 1097 1591 1101
rect 1595 1097 1596 1101
rect 1590 1096 1596 1097
rect 1622 1101 1628 1102
rect 1622 1097 1623 1101
rect 1627 1097 1628 1101
rect 1662 1099 1663 1103
rect 1667 1099 1668 1103
rect 1662 1098 1668 1099
rect 1622 1096 1628 1097
rect 1383 1092 1515 1094
rect 1383 1091 1384 1092
rect 1378 1090 1384 1091
rect 1558 1091 1564 1092
rect 1558 1087 1559 1091
rect 1563 1090 1564 1091
rect 1563 1088 1611 1090
rect 1563 1087 1564 1088
rect 1558 1086 1564 1087
rect 214 1083 220 1084
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 214 1079 215 1083
rect 219 1079 220 1083
rect 214 1078 220 1079
rect 246 1083 252 1084
rect 246 1079 247 1083
rect 251 1079 252 1083
rect 246 1078 252 1079
rect 278 1083 284 1084
rect 278 1079 279 1083
rect 283 1079 284 1083
rect 278 1078 284 1079
rect 310 1083 316 1084
rect 310 1079 311 1083
rect 315 1079 316 1083
rect 310 1078 316 1079
rect 350 1083 356 1084
rect 350 1079 351 1083
rect 355 1079 356 1083
rect 350 1078 356 1079
rect 390 1083 396 1084
rect 390 1079 391 1083
rect 395 1079 396 1083
rect 390 1078 396 1079
rect 438 1083 444 1084
rect 438 1079 439 1083
rect 443 1079 444 1083
rect 438 1078 444 1079
rect 502 1083 508 1084
rect 502 1079 503 1083
rect 507 1079 508 1083
rect 502 1078 508 1079
rect 574 1083 580 1084
rect 574 1079 575 1083
rect 579 1079 580 1083
rect 574 1078 580 1079
rect 654 1083 660 1084
rect 654 1079 655 1083
rect 659 1079 660 1083
rect 654 1078 660 1079
rect 734 1083 740 1084
rect 734 1079 735 1083
rect 739 1079 740 1083
rect 734 1078 740 1079
rect 814 1083 820 1084
rect 814 1079 815 1083
rect 819 1079 820 1083
rect 814 1078 820 1079
rect 894 1083 900 1084
rect 894 1079 895 1083
rect 899 1079 900 1083
rect 894 1078 900 1079
rect 966 1083 972 1084
rect 966 1079 967 1083
rect 971 1079 972 1083
rect 966 1078 972 1079
rect 1038 1083 1044 1084
rect 1038 1079 1039 1083
rect 1043 1079 1044 1083
rect 1038 1078 1044 1079
rect 1110 1083 1116 1084
rect 1110 1079 1111 1083
rect 1115 1079 1116 1083
rect 1110 1078 1116 1079
rect 1174 1083 1180 1084
rect 1174 1079 1175 1083
rect 1179 1079 1180 1083
rect 1174 1078 1180 1079
rect 1238 1083 1244 1084
rect 1238 1079 1239 1083
rect 1243 1079 1244 1083
rect 1238 1078 1244 1079
rect 1302 1083 1308 1084
rect 1302 1079 1303 1083
rect 1307 1079 1308 1083
rect 1302 1078 1308 1079
rect 1358 1083 1364 1084
rect 1358 1079 1359 1083
rect 1363 1079 1364 1083
rect 1358 1078 1364 1079
rect 1414 1083 1420 1084
rect 1414 1079 1415 1083
rect 1419 1079 1420 1083
rect 1414 1078 1420 1079
rect 1462 1083 1468 1084
rect 1462 1079 1463 1083
rect 1467 1079 1468 1083
rect 1462 1078 1468 1079
rect 1502 1083 1508 1084
rect 1502 1079 1503 1083
rect 1507 1079 1508 1083
rect 1502 1078 1508 1079
rect 1550 1083 1556 1084
rect 1550 1079 1551 1083
rect 1555 1079 1556 1083
rect 1550 1078 1556 1079
rect 1590 1083 1596 1084
rect 1590 1079 1591 1083
rect 1595 1079 1596 1083
rect 1590 1078 1596 1079
rect 110 1076 116 1077
rect 1609 1076 1611 1088
rect 1622 1083 1628 1084
rect 1622 1079 1623 1083
rect 1627 1079 1628 1083
rect 1622 1078 1628 1079
rect 1662 1081 1668 1082
rect 1662 1077 1663 1081
rect 1667 1077 1668 1081
rect 1662 1076 1668 1077
rect 231 1075 237 1076
rect 231 1071 232 1075
rect 236 1074 237 1075
rect 263 1075 269 1076
rect 236 1072 258 1074
rect 236 1071 237 1072
rect 231 1070 237 1071
rect 214 1066 220 1067
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 214 1062 215 1066
rect 219 1062 220 1066
rect 214 1061 220 1062
rect 246 1066 252 1067
rect 246 1062 247 1066
rect 251 1062 252 1066
rect 246 1061 252 1062
rect 110 1059 116 1060
rect 231 1059 240 1060
rect 231 1055 232 1059
rect 239 1055 240 1059
rect 256 1058 258 1072
rect 263 1071 264 1075
rect 268 1074 269 1075
rect 295 1075 304 1076
rect 268 1072 290 1074
rect 268 1071 269 1072
rect 263 1070 269 1071
rect 278 1066 284 1067
rect 278 1062 279 1066
rect 283 1062 284 1066
rect 278 1061 284 1062
rect 263 1059 269 1060
rect 263 1058 264 1059
rect 256 1056 264 1058
rect 231 1054 240 1055
rect 263 1055 264 1056
rect 268 1055 269 1059
rect 288 1058 290 1072
rect 295 1071 296 1075
rect 303 1071 304 1075
rect 295 1070 304 1071
rect 327 1075 333 1076
rect 327 1071 328 1075
rect 332 1074 333 1075
rect 367 1075 373 1076
rect 332 1072 347 1074
rect 332 1071 333 1072
rect 327 1070 333 1071
rect 310 1066 316 1067
rect 310 1062 311 1066
rect 315 1062 316 1066
rect 310 1061 316 1062
rect 295 1059 301 1060
rect 295 1058 296 1059
rect 288 1056 296 1058
rect 263 1054 269 1055
rect 295 1055 296 1056
rect 300 1055 301 1059
rect 295 1054 301 1055
rect 327 1059 333 1060
rect 327 1055 328 1059
rect 332 1058 333 1059
rect 345 1058 347 1072
rect 367 1071 368 1075
rect 372 1074 373 1075
rect 407 1075 413 1076
rect 372 1072 387 1074
rect 372 1071 373 1072
rect 367 1070 373 1071
rect 350 1066 356 1067
rect 350 1062 351 1066
rect 355 1062 356 1066
rect 350 1061 356 1062
rect 367 1059 373 1060
rect 367 1058 368 1059
rect 332 1056 342 1058
rect 345 1056 368 1058
rect 332 1055 333 1056
rect 327 1054 333 1055
rect 340 1050 342 1056
rect 367 1055 368 1056
rect 372 1055 373 1059
rect 385 1058 387 1072
rect 407 1071 408 1075
rect 412 1074 413 1075
rect 455 1075 461 1076
rect 412 1072 435 1074
rect 412 1071 413 1072
rect 407 1070 413 1071
rect 390 1066 396 1067
rect 390 1062 391 1066
rect 395 1062 396 1066
rect 390 1061 396 1062
rect 407 1059 413 1060
rect 407 1058 408 1059
rect 385 1056 408 1058
rect 367 1054 373 1055
rect 407 1055 408 1056
rect 412 1055 413 1059
rect 433 1058 435 1072
rect 455 1071 456 1075
rect 460 1074 461 1075
rect 519 1075 525 1076
rect 460 1072 514 1074
rect 460 1071 461 1072
rect 455 1070 461 1071
rect 438 1066 444 1067
rect 438 1062 439 1066
rect 443 1062 444 1066
rect 438 1061 444 1062
rect 502 1066 508 1067
rect 502 1062 503 1066
rect 507 1062 508 1066
rect 502 1061 508 1062
rect 455 1059 461 1060
rect 455 1058 456 1059
rect 433 1056 456 1058
rect 407 1054 413 1055
rect 455 1055 456 1056
rect 460 1055 461 1059
rect 512 1058 514 1072
rect 519 1071 520 1075
rect 524 1074 525 1075
rect 591 1075 597 1076
rect 524 1072 586 1074
rect 524 1071 525 1072
rect 519 1070 525 1071
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 519 1059 525 1060
rect 519 1058 520 1059
rect 512 1056 520 1058
rect 455 1054 461 1055
rect 519 1055 520 1056
rect 524 1055 525 1059
rect 584 1058 586 1072
rect 591 1071 592 1075
rect 596 1074 597 1075
rect 666 1075 677 1076
rect 596 1072 651 1074
rect 596 1071 597 1072
rect 591 1070 597 1071
rect 591 1059 597 1060
rect 591 1058 592 1059
rect 584 1056 592 1058
rect 519 1054 525 1055
rect 591 1055 592 1056
rect 596 1055 597 1059
rect 649 1058 651 1072
rect 666 1071 667 1075
rect 671 1071 672 1075
rect 676 1071 677 1075
rect 666 1070 677 1071
rect 751 1075 757 1076
rect 751 1071 752 1075
rect 756 1074 757 1075
rect 806 1075 812 1076
rect 806 1074 807 1075
rect 756 1072 807 1074
rect 756 1071 757 1072
rect 751 1070 757 1071
rect 806 1071 807 1072
rect 811 1071 812 1075
rect 831 1075 837 1076
rect 831 1074 832 1075
rect 806 1070 812 1071
rect 824 1072 832 1074
rect 654 1066 660 1067
rect 654 1062 655 1066
rect 659 1062 660 1066
rect 654 1061 660 1062
rect 734 1066 740 1067
rect 734 1062 735 1066
rect 739 1062 740 1066
rect 734 1061 740 1062
rect 814 1066 820 1067
rect 814 1062 815 1066
rect 819 1062 820 1066
rect 814 1061 820 1062
rect 671 1059 677 1060
rect 671 1058 672 1059
rect 649 1056 672 1058
rect 591 1054 597 1055
rect 671 1055 672 1056
rect 676 1055 677 1059
rect 671 1054 677 1055
rect 751 1059 757 1060
rect 751 1055 752 1059
rect 756 1058 757 1059
rect 824 1058 826 1072
rect 831 1071 832 1072
rect 836 1071 837 1075
rect 911 1075 917 1076
rect 911 1074 912 1075
rect 831 1070 837 1071
rect 876 1072 912 1074
rect 756 1056 826 1058
rect 831 1059 837 1060
rect 756 1055 757 1056
rect 751 1054 757 1055
rect 831 1055 832 1059
rect 836 1058 837 1059
rect 876 1058 878 1072
rect 911 1071 912 1072
rect 916 1071 917 1075
rect 911 1070 917 1071
rect 983 1075 989 1076
rect 983 1071 984 1075
rect 988 1074 989 1075
rect 1055 1075 1061 1076
rect 988 1072 1050 1074
rect 988 1071 989 1072
rect 983 1070 989 1071
rect 894 1066 900 1067
rect 894 1062 895 1066
rect 899 1062 900 1066
rect 894 1061 900 1062
rect 966 1066 972 1067
rect 966 1062 967 1066
rect 971 1062 972 1066
rect 966 1061 972 1062
rect 1038 1066 1044 1067
rect 1038 1062 1039 1066
rect 1043 1062 1044 1066
rect 1038 1061 1044 1062
rect 836 1056 878 1058
rect 902 1059 908 1060
rect 836 1055 837 1056
rect 831 1054 837 1055
rect 902 1055 903 1059
rect 907 1058 908 1059
rect 911 1059 917 1060
rect 911 1058 912 1059
rect 907 1056 912 1058
rect 907 1055 908 1056
rect 902 1054 908 1055
rect 911 1055 912 1056
rect 916 1055 917 1059
rect 911 1054 917 1055
rect 983 1059 989 1060
rect 983 1055 984 1059
rect 988 1055 989 1059
rect 1048 1058 1050 1072
rect 1055 1071 1056 1075
rect 1060 1074 1061 1075
rect 1127 1075 1133 1076
rect 1060 1072 1094 1074
rect 1060 1071 1061 1072
rect 1055 1070 1061 1071
rect 1055 1059 1061 1060
rect 1055 1058 1056 1059
rect 1048 1056 1056 1058
rect 983 1054 989 1055
rect 1055 1055 1056 1056
rect 1060 1055 1061 1059
rect 1092 1058 1094 1072
rect 1127 1071 1128 1075
rect 1132 1074 1133 1075
rect 1162 1075 1168 1076
rect 1162 1074 1163 1075
rect 1132 1072 1163 1074
rect 1132 1071 1133 1072
rect 1127 1070 1133 1071
rect 1162 1071 1163 1072
rect 1167 1071 1168 1075
rect 1162 1070 1168 1071
rect 1186 1075 1197 1076
rect 1186 1071 1187 1075
rect 1191 1071 1192 1075
rect 1196 1071 1197 1075
rect 1255 1075 1261 1076
rect 1255 1074 1256 1075
rect 1186 1070 1197 1071
rect 1228 1072 1256 1074
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1174 1066 1180 1067
rect 1174 1062 1175 1066
rect 1179 1062 1180 1066
rect 1174 1061 1180 1062
rect 1127 1059 1133 1060
rect 1127 1058 1128 1059
rect 1092 1056 1128 1058
rect 1055 1054 1061 1055
rect 1127 1055 1128 1056
rect 1132 1055 1133 1059
rect 1127 1054 1133 1055
rect 1191 1059 1197 1060
rect 1191 1055 1192 1059
rect 1196 1058 1197 1059
rect 1228 1058 1230 1072
rect 1255 1071 1256 1072
rect 1260 1071 1261 1075
rect 1319 1075 1325 1076
rect 1319 1074 1320 1075
rect 1255 1070 1261 1071
rect 1289 1072 1320 1074
rect 1238 1066 1244 1067
rect 1238 1062 1239 1066
rect 1243 1062 1244 1066
rect 1238 1061 1244 1062
rect 1196 1056 1230 1058
rect 1255 1059 1261 1060
rect 1196 1055 1197 1056
rect 1191 1054 1197 1055
rect 1255 1055 1256 1059
rect 1260 1058 1261 1059
rect 1289 1058 1291 1072
rect 1319 1071 1320 1072
rect 1324 1071 1325 1075
rect 1319 1070 1325 1071
rect 1375 1075 1381 1076
rect 1375 1071 1376 1075
rect 1380 1074 1381 1075
rect 1431 1075 1437 1076
rect 1380 1072 1406 1074
rect 1380 1071 1381 1072
rect 1375 1070 1381 1071
rect 1302 1066 1308 1067
rect 1302 1062 1303 1066
rect 1307 1062 1308 1066
rect 1302 1061 1308 1062
rect 1358 1066 1364 1067
rect 1358 1062 1359 1066
rect 1363 1062 1364 1066
rect 1358 1061 1364 1062
rect 1260 1056 1291 1058
rect 1310 1059 1316 1060
rect 1260 1055 1261 1056
rect 1255 1054 1261 1055
rect 1310 1055 1311 1059
rect 1315 1058 1316 1059
rect 1319 1059 1325 1060
rect 1319 1058 1320 1059
rect 1315 1056 1320 1058
rect 1315 1055 1316 1056
rect 1310 1054 1316 1055
rect 1319 1055 1320 1056
rect 1324 1055 1325 1059
rect 1319 1054 1325 1055
rect 1375 1059 1384 1060
rect 1375 1055 1376 1059
rect 1383 1055 1384 1059
rect 1404 1058 1406 1072
rect 1431 1071 1432 1075
rect 1436 1074 1437 1075
rect 1479 1075 1485 1076
rect 1436 1072 1458 1074
rect 1436 1071 1437 1072
rect 1431 1070 1437 1071
rect 1414 1066 1420 1067
rect 1414 1062 1415 1066
rect 1419 1062 1420 1066
rect 1414 1061 1420 1062
rect 1431 1059 1437 1060
rect 1431 1058 1432 1059
rect 1404 1056 1432 1058
rect 1375 1054 1384 1055
rect 1431 1055 1432 1056
rect 1436 1055 1437 1059
rect 1456 1058 1458 1072
rect 1479 1071 1480 1075
rect 1484 1074 1485 1075
rect 1519 1075 1525 1076
rect 1484 1072 1499 1074
rect 1484 1071 1485 1072
rect 1479 1070 1485 1071
rect 1462 1066 1468 1067
rect 1462 1062 1463 1066
rect 1467 1062 1468 1066
rect 1462 1061 1468 1062
rect 1479 1059 1485 1060
rect 1479 1058 1480 1059
rect 1456 1056 1480 1058
rect 1431 1054 1437 1055
rect 1479 1055 1480 1056
rect 1484 1055 1485 1059
rect 1497 1058 1499 1072
rect 1519 1071 1520 1075
rect 1524 1074 1525 1075
rect 1567 1075 1573 1076
rect 1524 1072 1547 1074
rect 1524 1071 1525 1072
rect 1519 1070 1525 1071
rect 1502 1066 1508 1067
rect 1502 1062 1503 1066
rect 1507 1062 1508 1066
rect 1502 1061 1508 1062
rect 1519 1059 1525 1060
rect 1519 1058 1520 1059
rect 1497 1056 1520 1058
rect 1479 1054 1485 1055
rect 1519 1055 1520 1056
rect 1524 1055 1525 1059
rect 1545 1058 1547 1072
rect 1567 1071 1568 1075
rect 1572 1074 1573 1075
rect 1607 1075 1613 1076
rect 1572 1072 1586 1074
rect 1572 1071 1573 1072
rect 1567 1070 1573 1071
rect 1550 1066 1556 1067
rect 1550 1062 1551 1066
rect 1555 1062 1556 1066
rect 1550 1061 1556 1062
rect 1567 1059 1573 1060
rect 1567 1058 1568 1059
rect 1545 1056 1568 1058
rect 1519 1054 1525 1055
rect 1567 1055 1568 1056
rect 1572 1055 1573 1059
rect 1584 1058 1586 1072
rect 1607 1071 1608 1075
rect 1612 1071 1613 1075
rect 1639 1075 1645 1076
rect 1639 1074 1640 1075
rect 1607 1070 1613 1071
rect 1616 1072 1640 1074
rect 1606 1067 1612 1068
rect 1590 1066 1596 1067
rect 1590 1062 1591 1066
rect 1595 1062 1596 1066
rect 1606 1063 1607 1067
rect 1611 1066 1612 1067
rect 1616 1066 1618 1072
rect 1639 1071 1640 1072
rect 1644 1071 1645 1075
rect 1639 1070 1645 1071
rect 1611 1064 1618 1066
rect 1622 1066 1628 1067
rect 1611 1063 1612 1064
rect 1606 1062 1612 1063
rect 1622 1062 1623 1066
rect 1627 1062 1628 1066
rect 1590 1061 1596 1062
rect 1622 1061 1628 1062
rect 1662 1064 1668 1065
rect 1662 1060 1663 1064
rect 1667 1060 1668 1064
rect 1607 1059 1613 1060
rect 1607 1058 1608 1059
rect 1584 1056 1608 1058
rect 1567 1054 1573 1055
rect 1607 1055 1608 1056
rect 1612 1055 1613 1059
rect 1607 1054 1613 1055
rect 1638 1059 1645 1060
rect 1662 1059 1668 1060
rect 1638 1055 1639 1059
rect 1644 1055 1645 1059
rect 1638 1054 1645 1055
rect 470 1051 476 1052
rect 470 1050 471 1051
rect 340 1048 471 1050
rect 470 1047 471 1048
rect 475 1047 476 1051
rect 985 1050 987 1054
rect 1186 1051 1192 1052
rect 1186 1050 1187 1051
rect 985 1048 1187 1050
rect 470 1046 476 1047
rect 666 1047 672 1048
rect 666 1046 667 1047
rect 521 1044 667 1046
rect 319 1036 347 1038
rect 385 1036 411 1038
rect 448 1036 475 1038
rect 521 1036 523 1044
rect 666 1043 667 1044
rect 671 1043 672 1047
rect 1186 1047 1187 1048
rect 1191 1047 1192 1051
rect 1186 1046 1192 1047
rect 1446 1047 1452 1048
rect 1446 1046 1447 1047
rect 666 1042 672 1043
rect 1353 1044 1447 1046
rect 527 1039 533 1040
rect 302 1035 308 1036
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 302 1031 303 1035
rect 307 1034 308 1035
rect 311 1035 317 1036
rect 311 1034 312 1035
rect 307 1032 312 1034
rect 307 1031 308 1032
rect 110 1027 116 1028
rect 294 1030 300 1031
rect 302 1030 308 1031
rect 311 1031 312 1032
rect 316 1031 317 1035
rect 311 1030 317 1031
rect 294 1026 295 1030
rect 299 1026 300 1030
rect 294 1025 300 1026
rect 311 1019 317 1020
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 311 1015 312 1019
rect 316 1018 317 1019
rect 319 1018 321 1036
rect 343 1035 349 1036
rect 343 1031 344 1035
rect 348 1031 349 1035
rect 375 1035 381 1036
rect 375 1034 376 1035
rect 368 1032 376 1034
rect 326 1030 332 1031
rect 343 1030 349 1031
rect 358 1030 364 1031
rect 326 1026 327 1030
rect 331 1026 332 1030
rect 326 1025 332 1026
rect 358 1026 359 1030
rect 363 1026 364 1030
rect 358 1025 364 1026
rect 368 1020 370 1032
rect 375 1031 376 1032
rect 380 1031 381 1035
rect 375 1030 381 1031
rect 316 1016 321 1018
rect 343 1019 349 1020
rect 316 1015 317 1016
rect 311 1014 317 1015
rect 343 1015 344 1019
rect 348 1018 349 1019
rect 356 1018 370 1020
rect 375 1019 381 1020
rect 348 1016 358 1018
rect 348 1015 349 1016
rect 343 1014 349 1015
rect 375 1015 376 1019
rect 380 1018 381 1019
rect 385 1018 387 1036
rect 407 1035 413 1036
rect 407 1031 408 1035
rect 412 1031 413 1035
rect 439 1035 445 1036
rect 439 1034 440 1035
rect 432 1032 440 1034
rect 390 1030 396 1031
rect 407 1030 413 1031
rect 422 1030 428 1031
rect 390 1026 391 1030
rect 395 1026 396 1030
rect 390 1025 396 1026
rect 422 1026 423 1030
rect 427 1026 428 1030
rect 422 1025 428 1026
rect 432 1020 434 1032
rect 439 1031 440 1032
rect 444 1031 445 1035
rect 439 1030 445 1031
rect 380 1016 387 1018
rect 407 1019 413 1020
rect 380 1015 381 1016
rect 375 1014 381 1015
rect 407 1015 408 1019
rect 412 1018 413 1019
rect 420 1018 434 1020
rect 439 1019 445 1020
rect 412 1016 422 1018
rect 412 1015 413 1016
rect 407 1014 413 1015
rect 439 1015 440 1019
rect 444 1018 445 1019
rect 448 1018 450 1036
rect 471 1035 477 1036
rect 471 1031 472 1035
rect 476 1031 477 1035
rect 519 1035 525 1036
rect 519 1031 520 1035
rect 524 1031 525 1035
rect 527 1035 528 1039
rect 532 1038 533 1039
rect 583 1039 589 1040
rect 532 1036 570 1038
rect 532 1035 533 1036
rect 527 1034 533 1035
rect 568 1034 570 1036
rect 575 1035 581 1036
rect 575 1034 576 1035
rect 568 1032 576 1034
rect 575 1031 576 1032
rect 580 1031 581 1035
rect 583 1035 584 1039
rect 588 1038 589 1039
rect 655 1039 661 1040
rect 588 1036 651 1038
rect 588 1035 589 1036
rect 583 1034 589 1035
rect 647 1035 653 1036
rect 647 1031 648 1035
rect 652 1031 653 1035
rect 655 1035 656 1039
rect 660 1038 661 1039
rect 823 1039 829 1040
rect 660 1036 722 1038
rect 660 1035 661 1036
rect 655 1034 661 1035
rect 720 1034 722 1036
rect 727 1035 733 1036
rect 727 1034 728 1035
rect 720 1032 728 1034
rect 727 1031 728 1032
rect 732 1031 733 1035
rect 806 1035 812 1036
rect 806 1031 807 1035
rect 811 1034 812 1035
rect 815 1035 821 1036
rect 815 1034 816 1035
rect 811 1032 816 1034
rect 811 1031 812 1032
rect 454 1030 460 1031
rect 471 1030 477 1031
rect 502 1030 508 1031
rect 519 1030 525 1031
rect 558 1030 564 1031
rect 575 1030 581 1031
rect 630 1030 636 1031
rect 647 1030 653 1031
rect 710 1030 716 1031
rect 727 1030 733 1031
rect 798 1030 804 1031
rect 806 1030 812 1031
rect 815 1031 816 1032
rect 820 1031 821 1035
rect 823 1035 824 1039
rect 828 1038 829 1039
rect 983 1039 989 1040
rect 828 1036 899 1038
rect 828 1035 829 1036
rect 823 1034 829 1035
rect 895 1035 901 1036
rect 895 1031 896 1035
rect 900 1031 901 1035
rect 974 1035 981 1036
rect 974 1031 975 1035
rect 980 1031 981 1035
rect 983 1035 984 1039
rect 988 1038 989 1039
rect 1055 1039 1061 1040
rect 988 1036 1051 1038
rect 988 1035 989 1036
rect 983 1034 989 1035
rect 1047 1035 1053 1036
rect 1047 1031 1048 1035
rect 1052 1031 1053 1035
rect 1055 1035 1056 1039
rect 1060 1038 1061 1039
rect 1119 1039 1125 1040
rect 1060 1036 1115 1038
rect 1060 1035 1061 1036
rect 1055 1034 1061 1035
rect 1111 1035 1117 1036
rect 1111 1031 1112 1035
rect 1116 1031 1117 1035
rect 1119 1035 1120 1039
rect 1124 1038 1125 1039
rect 1183 1039 1189 1040
rect 1124 1036 1179 1038
rect 1124 1035 1125 1036
rect 1119 1034 1125 1035
rect 1175 1035 1181 1036
rect 1175 1031 1176 1035
rect 1180 1031 1181 1035
rect 1183 1035 1184 1039
rect 1188 1038 1189 1039
rect 1247 1039 1253 1040
rect 1188 1036 1234 1038
rect 1188 1035 1189 1036
rect 1183 1034 1189 1035
rect 1232 1034 1234 1036
rect 1239 1035 1245 1036
rect 1239 1034 1240 1035
rect 1232 1032 1240 1034
rect 1239 1031 1240 1032
rect 1244 1031 1245 1035
rect 1247 1035 1248 1039
rect 1252 1038 1253 1039
rect 1252 1036 1299 1038
rect 1353 1036 1355 1044
rect 1446 1043 1447 1044
rect 1451 1043 1452 1047
rect 1446 1042 1452 1043
rect 1359 1039 1365 1040
rect 1252 1035 1253 1036
rect 1247 1034 1253 1035
rect 1295 1035 1301 1036
rect 1295 1031 1296 1035
rect 1300 1031 1301 1035
rect 1351 1035 1357 1036
rect 1351 1031 1352 1035
rect 1356 1031 1357 1035
rect 1359 1035 1360 1039
rect 1364 1038 1365 1039
rect 1364 1036 1394 1038
rect 1472 1036 1490 1038
rect 1497 1036 1546 1038
rect 1616 1036 1643 1038
rect 1364 1035 1365 1036
rect 1359 1034 1365 1035
rect 1392 1034 1394 1036
rect 1399 1035 1405 1036
rect 1399 1034 1400 1035
rect 1392 1032 1400 1034
rect 1399 1031 1400 1032
rect 1404 1031 1405 1035
rect 1447 1035 1453 1036
rect 1447 1031 1448 1035
rect 1452 1034 1453 1035
rect 1472 1034 1474 1036
rect 1452 1032 1474 1034
rect 1452 1031 1453 1032
rect 815 1030 821 1031
rect 878 1030 884 1031
rect 895 1030 901 1031
rect 958 1030 964 1031
rect 974 1030 981 1031
rect 1030 1030 1036 1031
rect 1047 1030 1053 1031
rect 1094 1030 1100 1031
rect 1111 1030 1117 1031
rect 1158 1030 1164 1031
rect 1175 1030 1181 1031
rect 1222 1030 1228 1031
rect 1239 1030 1245 1031
rect 1278 1030 1284 1031
rect 1295 1030 1301 1031
rect 1334 1030 1340 1031
rect 1351 1030 1357 1031
rect 1382 1030 1388 1031
rect 1399 1030 1405 1031
rect 1430 1030 1436 1031
rect 1447 1030 1453 1031
rect 1478 1030 1484 1031
rect 454 1026 455 1030
rect 459 1026 460 1030
rect 454 1025 460 1026
rect 502 1026 503 1030
rect 507 1026 508 1030
rect 502 1025 508 1026
rect 558 1026 559 1030
rect 563 1026 564 1030
rect 558 1025 564 1026
rect 630 1026 631 1030
rect 635 1026 636 1030
rect 630 1025 636 1026
rect 710 1026 711 1030
rect 715 1026 716 1030
rect 710 1025 716 1026
rect 798 1026 799 1030
rect 803 1026 804 1030
rect 798 1025 804 1026
rect 878 1026 879 1030
rect 883 1026 884 1030
rect 878 1025 884 1026
rect 958 1026 959 1030
rect 963 1026 964 1030
rect 958 1025 964 1026
rect 1030 1026 1031 1030
rect 1035 1026 1036 1030
rect 1030 1025 1036 1026
rect 1094 1026 1095 1030
rect 1099 1026 1100 1030
rect 1094 1025 1100 1026
rect 1158 1026 1159 1030
rect 1163 1026 1164 1030
rect 1158 1025 1164 1026
rect 1222 1026 1223 1030
rect 1227 1026 1228 1030
rect 1222 1025 1228 1026
rect 1278 1026 1279 1030
rect 1283 1026 1284 1030
rect 1278 1025 1284 1026
rect 1334 1026 1335 1030
rect 1339 1026 1340 1030
rect 1334 1025 1340 1026
rect 1382 1026 1383 1030
rect 1387 1026 1388 1030
rect 1382 1025 1388 1026
rect 1430 1026 1431 1030
rect 1435 1026 1436 1030
rect 1430 1025 1436 1026
rect 1478 1026 1479 1030
rect 1483 1026 1484 1030
rect 1478 1025 1484 1026
rect 1488 1022 1490 1036
rect 1495 1035 1501 1036
rect 1495 1031 1496 1035
rect 1500 1031 1501 1035
rect 1495 1030 1501 1031
rect 1534 1030 1540 1031
rect 1534 1026 1535 1030
rect 1539 1026 1540 1030
rect 1534 1025 1540 1026
rect 1488 1020 1499 1022
rect 444 1016 450 1018
rect 470 1019 477 1020
rect 444 1015 445 1016
rect 439 1014 445 1015
rect 470 1015 471 1019
rect 476 1015 477 1019
rect 470 1014 477 1015
rect 519 1019 525 1020
rect 519 1015 520 1019
rect 524 1018 525 1019
rect 527 1019 533 1020
rect 527 1018 528 1019
rect 524 1016 528 1018
rect 524 1015 525 1016
rect 519 1014 525 1015
rect 527 1015 528 1016
rect 532 1015 533 1019
rect 527 1014 533 1015
rect 575 1019 581 1020
rect 575 1015 576 1019
rect 580 1018 581 1019
rect 583 1019 589 1020
rect 583 1018 584 1019
rect 580 1016 584 1018
rect 580 1015 581 1016
rect 575 1014 581 1015
rect 583 1015 584 1016
rect 588 1015 589 1019
rect 583 1014 589 1015
rect 647 1019 653 1020
rect 647 1015 648 1019
rect 652 1018 653 1019
rect 655 1019 661 1020
rect 655 1018 656 1019
rect 652 1016 656 1018
rect 652 1015 653 1016
rect 647 1014 653 1015
rect 655 1015 656 1016
rect 660 1015 661 1019
rect 727 1019 733 1020
rect 727 1018 728 1019
rect 655 1014 661 1015
rect 720 1016 728 1018
rect 110 1010 116 1011
rect 294 1013 300 1014
rect 294 1009 295 1013
rect 299 1009 300 1013
rect 294 1008 300 1009
rect 326 1013 332 1014
rect 326 1009 327 1013
rect 331 1009 332 1013
rect 326 1008 332 1009
rect 358 1013 364 1014
rect 358 1009 359 1013
rect 363 1009 364 1013
rect 358 1008 364 1009
rect 390 1013 396 1014
rect 390 1009 391 1013
rect 395 1009 396 1013
rect 390 1008 396 1009
rect 422 1013 428 1014
rect 422 1009 423 1013
rect 427 1009 428 1013
rect 422 1008 428 1009
rect 454 1013 460 1014
rect 454 1009 455 1013
rect 459 1009 460 1013
rect 454 1008 460 1009
rect 502 1013 508 1014
rect 502 1009 503 1013
rect 507 1009 508 1013
rect 502 1008 508 1009
rect 558 1013 564 1014
rect 558 1009 559 1013
rect 563 1009 564 1013
rect 558 1008 564 1009
rect 630 1013 636 1014
rect 630 1009 631 1013
rect 635 1009 636 1013
rect 630 1008 636 1009
rect 710 1013 716 1014
rect 710 1009 711 1013
rect 715 1009 716 1013
rect 710 1008 716 1009
rect 302 1007 308 1008
rect 302 1003 303 1007
rect 307 1006 308 1007
rect 510 1007 516 1008
rect 307 1004 434 1006
rect 307 1003 308 1004
rect 302 1002 308 1003
rect 246 999 252 1000
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 246 995 247 999
rect 251 995 252 999
rect 246 994 252 995
rect 278 999 284 1000
rect 278 995 279 999
rect 283 995 284 999
rect 278 994 284 995
rect 310 999 316 1000
rect 310 995 311 999
rect 315 995 316 999
rect 310 994 316 995
rect 342 999 348 1000
rect 342 995 343 999
rect 347 995 348 999
rect 342 994 348 995
rect 382 999 388 1000
rect 382 995 383 999
rect 387 995 388 999
rect 382 994 388 995
rect 422 999 428 1000
rect 422 995 423 999
rect 427 995 428 999
rect 422 994 428 995
rect 110 992 116 993
rect 263 991 269 992
rect 263 987 264 991
rect 268 990 269 991
rect 295 991 301 992
rect 268 988 290 990
rect 268 987 269 988
rect 263 986 269 987
rect 246 982 252 983
rect 110 980 116 981
rect 110 976 111 980
rect 115 976 116 980
rect 246 978 247 982
rect 251 978 252 982
rect 246 977 252 978
rect 278 982 284 983
rect 278 978 279 982
rect 283 978 284 982
rect 288 982 290 988
rect 295 987 296 991
rect 300 990 301 991
rect 327 991 333 992
rect 300 988 321 990
rect 300 987 301 988
rect 295 986 301 987
rect 310 982 316 983
rect 288 980 298 982
rect 296 978 298 980
rect 310 978 311 982
rect 315 978 316 982
rect 278 977 284 978
rect 295 977 301 978
rect 310 977 316 978
rect 110 975 116 976
rect 263 975 269 976
rect 263 971 264 975
rect 268 974 269 975
rect 268 972 290 974
rect 295 973 296 977
rect 300 973 301 977
rect 295 972 301 973
rect 319 974 321 988
rect 327 987 328 991
rect 332 990 333 991
rect 359 991 365 992
rect 332 988 354 990
rect 332 987 333 988
rect 327 986 333 987
rect 342 982 348 983
rect 342 978 343 982
rect 347 978 348 982
rect 342 977 348 978
rect 327 975 333 976
rect 327 974 328 975
rect 319 972 328 974
rect 268 971 269 972
rect 263 970 269 971
rect 288 966 290 972
rect 327 971 328 972
rect 332 971 333 975
rect 352 974 354 988
rect 359 987 360 991
rect 364 990 365 991
rect 399 991 405 992
rect 364 988 378 990
rect 364 987 365 988
rect 359 986 365 987
rect 359 975 365 976
rect 359 974 360 975
rect 352 972 360 974
rect 327 970 333 971
rect 359 971 360 972
rect 364 971 365 975
rect 376 974 378 988
rect 399 987 400 991
rect 404 990 405 991
rect 432 990 434 1004
rect 510 1003 511 1007
rect 515 1006 516 1007
rect 720 1006 722 1016
rect 727 1015 728 1016
rect 732 1015 733 1019
rect 727 1014 733 1015
rect 815 1019 821 1020
rect 815 1015 816 1019
rect 820 1018 821 1019
rect 823 1019 829 1020
rect 823 1018 824 1019
rect 820 1016 824 1018
rect 820 1015 821 1016
rect 815 1014 821 1015
rect 823 1015 824 1016
rect 828 1015 829 1019
rect 823 1014 829 1015
rect 890 1019 901 1020
rect 890 1015 891 1019
rect 895 1015 896 1019
rect 900 1015 901 1019
rect 890 1014 901 1015
rect 975 1019 981 1020
rect 975 1015 976 1019
rect 980 1018 981 1019
rect 983 1019 989 1020
rect 983 1018 984 1019
rect 980 1016 984 1018
rect 980 1015 981 1016
rect 975 1014 981 1015
rect 983 1015 984 1016
rect 988 1015 989 1019
rect 983 1014 989 1015
rect 1047 1019 1053 1020
rect 1047 1015 1048 1019
rect 1052 1018 1053 1019
rect 1055 1019 1061 1020
rect 1055 1018 1056 1019
rect 1052 1016 1056 1018
rect 1052 1015 1053 1016
rect 1047 1014 1053 1015
rect 1055 1015 1056 1016
rect 1060 1015 1061 1019
rect 1055 1014 1061 1015
rect 1111 1019 1117 1020
rect 1111 1015 1112 1019
rect 1116 1018 1117 1019
rect 1119 1019 1125 1020
rect 1119 1018 1120 1019
rect 1116 1016 1120 1018
rect 1116 1015 1117 1016
rect 1111 1014 1117 1015
rect 1119 1015 1120 1016
rect 1124 1015 1125 1019
rect 1119 1014 1125 1015
rect 1175 1019 1181 1020
rect 1175 1015 1176 1019
rect 1180 1018 1181 1019
rect 1183 1019 1189 1020
rect 1183 1018 1184 1019
rect 1180 1016 1184 1018
rect 1180 1015 1181 1016
rect 1175 1014 1181 1015
rect 1183 1015 1184 1016
rect 1188 1015 1189 1019
rect 1183 1014 1189 1015
rect 1239 1019 1245 1020
rect 1239 1015 1240 1019
rect 1244 1018 1245 1019
rect 1247 1019 1253 1020
rect 1247 1018 1248 1019
rect 1244 1016 1248 1018
rect 1244 1015 1245 1016
rect 1239 1014 1245 1015
rect 1247 1015 1248 1016
rect 1252 1015 1253 1019
rect 1247 1014 1253 1015
rect 1295 1019 1301 1020
rect 1295 1015 1296 1019
rect 1300 1018 1301 1019
rect 1310 1019 1316 1020
rect 1310 1018 1311 1019
rect 1300 1016 1311 1018
rect 1300 1015 1301 1016
rect 1295 1014 1301 1015
rect 1310 1015 1311 1016
rect 1315 1015 1316 1019
rect 1310 1014 1316 1015
rect 1351 1019 1357 1020
rect 1351 1015 1352 1019
rect 1356 1018 1357 1019
rect 1359 1019 1365 1020
rect 1359 1018 1360 1019
rect 1356 1016 1360 1018
rect 1356 1015 1357 1016
rect 1351 1014 1357 1015
rect 1359 1015 1360 1016
rect 1364 1015 1365 1019
rect 1359 1014 1365 1015
rect 1399 1019 1405 1020
rect 1399 1015 1400 1019
rect 1404 1018 1405 1019
rect 1414 1019 1420 1020
rect 1414 1018 1415 1019
rect 1404 1016 1415 1018
rect 1404 1015 1405 1016
rect 1399 1014 1405 1015
rect 1414 1015 1415 1016
rect 1419 1015 1420 1019
rect 1414 1014 1420 1015
rect 1446 1019 1453 1020
rect 1446 1015 1447 1019
rect 1452 1015 1453 1019
rect 1446 1014 1453 1015
rect 1495 1019 1501 1020
rect 1495 1015 1496 1019
rect 1500 1015 1501 1019
rect 1544 1018 1546 1036
rect 1551 1035 1560 1036
rect 1551 1031 1552 1035
rect 1559 1031 1560 1035
rect 1606 1035 1613 1036
rect 1606 1031 1607 1035
rect 1612 1031 1613 1035
rect 1551 1030 1560 1031
rect 1590 1030 1596 1031
rect 1606 1030 1613 1031
rect 1590 1026 1591 1030
rect 1595 1026 1596 1030
rect 1590 1025 1596 1026
rect 1551 1019 1557 1020
rect 1551 1018 1552 1019
rect 1544 1016 1552 1018
rect 1495 1014 1501 1015
rect 1551 1015 1552 1016
rect 1556 1015 1557 1019
rect 1551 1014 1557 1015
rect 1607 1019 1613 1020
rect 1607 1015 1608 1019
rect 1612 1018 1613 1019
rect 1616 1018 1618 1036
rect 1639 1035 1645 1036
rect 1639 1031 1640 1035
rect 1644 1031 1645 1035
rect 1622 1030 1628 1031
rect 1639 1030 1645 1031
rect 1662 1032 1668 1033
rect 1622 1026 1623 1030
rect 1627 1026 1628 1030
rect 1662 1028 1663 1032
rect 1667 1028 1668 1032
rect 1662 1027 1668 1028
rect 1622 1025 1628 1026
rect 1612 1016 1618 1018
rect 1638 1019 1645 1020
rect 1612 1015 1613 1016
rect 1607 1014 1613 1015
rect 1638 1015 1639 1019
rect 1644 1015 1645 1019
rect 1638 1014 1645 1015
rect 1662 1015 1668 1016
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 878 1013 884 1014
rect 878 1009 879 1013
rect 883 1009 884 1013
rect 878 1008 884 1009
rect 958 1013 964 1014
rect 958 1009 959 1013
rect 963 1009 964 1013
rect 958 1008 964 1009
rect 1030 1013 1036 1014
rect 1030 1009 1031 1013
rect 1035 1009 1036 1013
rect 1030 1008 1036 1009
rect 1094 1013 1100 1014
rect 1094 1009 1095 1013
rect 1099 1009 1100 1013
rect 1094 1008 1100 1009
rect 1158 1013 1164 1014
rect 1158 1009 1159 1013
rect 1163 1009 1164 1013
rect 1158 1008 1164 1009
rect 1222 1013 1228 1014
rect 1222 1009 1223 1013
rect 1227 1009 1228 1013
rect 1222 1008 1228 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 1334 1013 1340 1014
rect 1334 1009 1335 1013
rect 1339 1009 1340 1013
rect 1334 1008 1340 1009
rect 1382 1013 1388 1014
rect 1382 1009 1383 1013
rect 1387 1009 1388 1013
rect 1382 1008 1388 1009
rect 1430 1013 1436 1014
rect 1430 1009 1431 1013
rect 1435 1009 1436 1013
rect 1430 1008 1436 1009
rect 1478 1013 1484 1014
rect 1478 1009 1479 1013
rect 1483 1009 1484 1013
rect 1478 1008 1484 1009
rect 1534 1013 1540 1014
rect 1534 1009 1535 1013
rect 1539 1009 1540 1013
rect 1534 1008 1540 1009
rect 1590 1013 1596 1014
rect 1590 1009 1591 1013
rect 1595 1009 1596 1013
rect 1590 1008 1596 1009
rect 1622 1013 1628 1014
rect 1622 1009 1623 1013
rect 1627 1009 1628 1013
rect 1662 1011 1663 1015
rect 1667 1011 1668 1015
rect 1662 1010 1668 1011
rect 1622 1008 1628 1009
rect 515 1004 722 1006
rect 974 1007 980 1008
rect 515 1003 516 1004
rect 510 1002 516 1003
rect 974 1003 975 1007
rect 979 1006 980 1007
rect 979 1004 1234 1006
rect 979 1003 980 1004
rect 974 1002 980 1003
rect 478 999 484 1000
rect 478 995 479 999
rect 483 995 484 999
rect 478 994 484 995
rect 542 999 548 1000
rect 542 995 543 999
rect 547 995 548 999
rect 542 994 548 995
rect 614 999 620 1000
rect 614 995 615 999
rect 619 995 620 999
rect 614 994 620 995
rect 686 999 692 1000
rect 686 995 687 999
rect 691 995 692 999
rect 686 994 692 995
rect 758 999 764 1000
rect 758 995 759 999
rect 763 995 764 999
rect 758 994 764 995
rect 830 999 836 1000
rect 830 995 831 999
rect 835 995 836 999
rect 830 994 836 995
rect 902 999 908 1000
rect 902 995 903 999
rect 907 995 908 999
rect 902 994 908 995
rect 966 999 972 1000
rect 966 995 967 999
rect 971 995 972 999
rect 966 994 972 995
rect 1030 999 1036 1000
rect 1030 995 1031 999
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1094 999 1100 1000
rect 1094 995 1095 999
rect 1099 995 1100 999
rect 1094 994 1100 995
rect 1158 999 1164 1000
rect 1158 995 1159 999
rect 1163 995 1164 999
rect 1158 994 1164 995
rect 1222 999 1228 1000
rect 1222 995 1223 999
rect 1227 995 1228 999
rect 1222 994 1228 995
rect 439 991 445 992
rect 439 990 440 991
rect 404 988 418 990
rect 432 988 440 990
rect 404 987 405 988
rect 399 986 405 987
rect 382 982 388 983
rect 382 978 383 982
rect 387 978 388 982
rect 382 977 388 978
rect 399 975 405 976
rect 399 974 400 975
rect 376 972 400 974
rect 359 970 365 971
rect 399 971 400 972
rect 404 971 405 975
rect 416 974 418 988
rect 439 987 440 988
rect 444 987 445 991
rect 439 986 445 987
rect 495 991 501 992
rect 495 987 496 991
rect 500 990 501 991
rect 559 991 565 992
rect 500 988 530 990
rect 500 987 501 988
rect 495 986 501 987
rect 422 982 428 983
rect 422 978 423 982
rect 427 978 428 982
rect 422 977 428 978
rect 478 982 484 983
rect 478 978 479 982
rect 483 978 484 982
rect 478 977 484 978
rect 439 975 445 976
rect 439 974 440 975
rect 416 972 440 974
rect 399 970 405 971
rect 439 971 440 972
rect 444 971 445 975
rect 439 970 445 971
rect 495 975 501 976
rect 495 971 496 975
rect 500 974 501 975
rect 510 975 516 976
rect 510 974 511 975
rect 500 972 511 974
rect 500 971 501 972
rect 495 970 501 971
rect 510 971 511 972
rect 515 971 516 975
rect 528 974 530 988
rect 559 987 560 991
rect 564 990 565 991
rect 631 991 637 992
rect 564 988 598 990
rect 564 987 565 988
rect 559 986 565 987
rect 542 982 548 983
rect 542 978 543 982
rect 547 978 548 982
rect 542 977 548 978
rect 559 975 565 976
rect 559 974 560 975
rect 528 972 560 974
rect 510 970 516 971
rect 559 971 560 972
rect 564 971 565 975
rect 596 974 598 988
rect 631 987 632 991
rect 636 990 637 991
rect 674 991 680 992
rect 636 988 670 990
rect 636 987 637 988
rect 631 986 637 987
rect 614 982 620 983
rect 614 978 615 982
rect 619 978 620 982
rect 614 977 620 978
rect 631 975 637 976
rect 631 974 632 975
rect 596 972 632 974
rect 559 970 565 971
rect 631 971 632 972
rect 636 971 637 975
rect 668 974 670 988
rect 674 987 675 991
rect 679 990 680 991
rect 703 991 709 992
rect 703 990 704 991
rect 679 988 704 990
rect 679 987 680 988
rect 674 986 680 987
rect 703 987 704 988
rect 708 987 709 991
rect 703 986 709 987
rect 775 991 781 992
rect 775 987 776 991
rect 780 990 781 991
rect 806 991 812 992
rect 806 990 807 991
rect 780 988 807 990
rect 780 987 781 988
rect 775 986 781 987
rect 806 987 807 988
rect 811 987 812 991
rect 847 991 853 992
rect 847 990 848 991
rect 806 986 812 987
rect 816 988 848 990
rect 686 982 692 983
rect 686 978 687 982
rect 691 978 692 982
rect 686 977 692 978
rect 758 982 764 983
rect 758 978 759 982
rect 763 978 764 982
rect 758 977 764 978
rect 703 975 709 976
rect 703 974 704 975
rect 668 972 704 974
rect 631 970 637 971
rect 703 971 704 972
rect 708 971 709 975
rect 703 970 709 971
rect 775 975 781 976
rect 775 971 776 975
rect 780 974 781 975
rect 816 974 818 988
rect 847 987 848 988
rect 852 987 853 991
rect 847 986 853 987
rect 919 991 925 992
rect 919 987 920 991
rect 924 990 925 991
rect 983 991 989 992
rect 924 988 978 990
rect 924 987 925 988
rect 919 986 925 987
rect 830 982 836 983
rect 830 978 831 982
rect 835 978 836 982
rect 830 977 836 978
rect 902 982 908 983
rect 902 978 903 982
rect 907 978 908 982
rect 902 977 908 978
rect 966 982 972 983
rect 966 978 967 982
rect 971 978 972 982
rect 966 977 972 978
rect 780 972 818 974
rect 847 975 853 976
rect 780 971 781 972
rect 775 970 781 971
rect 847 971 848 975
rect 852 974 853 975
rect 890 975 896 976
rect 890 974 891 975
rect 852 972 891 974
rect 852 971 853 972
rect 847 970 853 971
rect 890 971 891 972
rect 895 971 896 975
rect 890 970 896 971
rect 919 975 925 976
rect 919 971 920 975
rect 924 971 925 975
rect 976 974 978 988
rect 983 987 984 991
rect 988 990 989 991
rect 1047 991 1053 992
rect 988 988 1042 990
rect 988 987 989 988
rect 983 986 989 987
rect 1030 982 1036 983
rect 1030 978 1031 982
rect 1035 978 1036 982
rect 1030 977 1036 978
rect 983 975 989 976
rect 983 974 984 975
rect 976 972 984 974
rect 919 970 925 971
rect 983 971 984 972
rect 988 971 989 975
rect 1040 974 1042 988
rect 1047 987 1048 991
rect 1052 990 1053 991
rect 1111 991 1117 992
rect 1052 988 1106 990
rect 1052 987 1053 988
rect 1047 986 1053 987
rect 1094 982 1100 983
rect 1094 978 1095 982
rect 1099 978 1100 982
rect 1094 977 1100 978
rect 1047 975 1053 976
rect 1047 974 1048 975
rect 1040 972 1048 974
rect 983 970 989 971
rect 1047 971 1048 972
rect 1052 971 1053 975
rect 1104 974 1106 988
rect 1111 987 1112 991
rect 1116 990 1117 991
rect 1175 991 1181 992
rect 1116 988 1170 990
rect 1116 987 1117 988
rect 1111 986 1117 987
rect 1158 982 1164 983
rect 1158 978 1159 982
rect 1163 978 1164 982
rect 1158 977 1164 978
rect 1111 975 1117 976
rect 1111 974 1112 975
rect 1104 972 1112 974
rect 1047 970 1053 971
rect 1111 971 1112 972
rect 1116 971 1117 975
rect 1168 974 1170 988
rect 1175 987 1176 991
rect 1180 990 1181 991
rect 1232 990 1234 1004
rect 1286 999 1292 1000
rect 1286 995 1287 999
rect 1291 995 1292 999
rect 1286 994 1292 995
rect 1342 999 1348 1000
rect 1342 995 1343 999
rect 1347 995 1348 999
rect 1342 994 1348 995
rect 1398 999 1404 1000
rect 1398 995 1399 999
rect 1403 995 1404 999
rect 1398 994 1404 995
rect 1446 999 1452 1000
rect 1446 995 1447 999
rect 1451 995 1452 999
rect 1446 994 1452 995
rect 1494 999 1500 1000
rect 1494 995 1495 999
rect 1499 995 1500 999
rect 1494 994 1500 995
rect 1542 999 1548 1000
rect 1542 995 1543 999
rect 1547 995 1548 999
rect 1542 994 1548 995
rect 1590 999 1596 1000
rect 1590 995 1591 999
rect 1595 995 1596 999
rect 1590 994 1596 995
rect 1622 999 1628 1000
rect 1622 995 1623 999
rect 1627 995 1628 999
rect 1622 994 1628 995
rect 1662 997 1668 998
rect 1662 993 1663 997
rect 1667 993 1668 997
rect 1662 992 1668 993
rect 1239 991 1245 992
rect 1239 990 1240 991
rect 1180 988 1219 990
rect 1232 988 1240 990
rect 1180 987 1181 988
rect 1175 986 1181 987
rect 1175 975 1181 976
rect 1175 974 1176 975
rect 1168 972 1176 974
rect 1111 970 1117 971
rect 1175 971 1176 972
rect 1180 971 1181 975
rect 1217 974 1219 988
rect 1239 987 1240 988
rect 1244 987 1245 991
rect 1239 986 1245 987
rect 1303 991 1309 992
rect 1303 987 1304 991
rect 1308 990 1309 991
rect 1322 991 1328 992
rect 1322 990 1323 991
rect 1308 988 1323 990
rect 1308 987 1309 988
rect 1303 986 1309 987
rect 1322 987 1323 988
rect 1327 987 1328 991
rect 1359 991 1365 992
rect 1359 990 1360 991
rect 1322 986 1328 987
rect 1332 988 1360 990
rect 1222 982 1228 983
rect 1222 978 1223 982
rect 1227 978 1228 982
rect 1222 977 1228 978
rect 1286 982 1292 983
rect 1286 978 1287 982
rect 1291 978 1292 982
rect 1286 977 1292 978
rect 1239 975 1245 976
rect 1239 974 1240 975
rect 1217 972 1240 974
rect 1175 970 1181 971
rect 1239 971 1240 972
rect 1244 971 1245 975
rect 1239 970 1245 971
rect 1303 975 1309 976
rect 1303 971 1304 975
rect 1308 974 1309 975
rect 1332 974 1334 988
rect 1359 987 1360 988
rect 1364 987 1365 991
rect 1415 991 1421 992
rect 1415 990 1416 991
rect 1359 986 1365 987
rect 1388 988 1416 990
rect 1342 982 1348 983
rect 1342 978 1343 982
rect 1347 978 1348 982
rect 1342 977 1348 978
rect 1308 972 1334 974
rect 1359 975 1365 976
rect 1308 971 1309 972
rect 1303 970 1309 971
rect 1359 971 1360 975
rect 1364 974 1365 975
rect 1388 974 1390 988
rect 1415 987 1416 988
rect 1420 987 1421 991
rect 1415 986 1421 987
rect 1463 991 1469 992
rect 1463 987 1464 991
rect 1468 990 1469 991
rect 1511 991 1517 992
rect 1468 988 1506 990
rect 1468 987 1469 988
rect 1463 986 1469 987
rect 1398 982 1404 983
rect 1398 978 1399 982
rect 1403 978 1404 982
rect 1398 977 1404 978
rect 1446 982 1452 983
rect 1446 978 1447 982
rect 1451 978 1452 982
rect 1446 977 1452 978
rect 1494 982 1500 983
rect 1494 978 1495 982
rect 1499 978 1500 982
rect 1494 977 1500 978
rect 1364 972 1390 974
rect 1414 975 1421 976
rect 1364 971 1365 972
rect 1359 970 1365 971
rect 1414 971 1415 975
rect 1420 971 1421 975
rect 1414 970 1421 971
rect 1458 975 1469 976
rect 1458 971 1459 975
rect 1463 971 1464 975
rect 1468 971 1469 975
rect 1504 974 1506 988
rect 1511 987 1512 991
rect 1516 990 1517 991
rect 1554 991 1565 992
rect 1516 988 1539 990
rect 1516 987 1517 988
rect 1511 986 1517 987
rect 1511 975 1517 976
rect 1511 974 1512 975
rect 1504 972 1512 974
rect 1458 970 1469 971
rect 1511 971 1512 972
rect 1516 971 1517 975
rect 1537 974 1539 988
rect 1554 987 1555 991
rect 1559 987 1560 991
rect 1564 987 1565 991
rect 1554 986 1565 987
rect 1606 991 1613 992
rect 1606 987 1607 991
rect 1612 987 1613 991
rect 1639 991 1645 992
rect 1639 990 1640 991
rect 1606 986 1613 987
rect 1632 988 1640 990
rect 1542 982 1548 983
rect 1542 978 1543 982
rect 1547 978 1548 982
rect 1542 977 1548 978
rect 1590 982 1596 983
rect 1590 978 1591 982
rect 1595 978 1596 982
rect 1590 977 1596 978
rect 1622 982 1628 983
rect 1622 978 1623 982
rect 1627 978 1628 982
rect 1622 977 1628 978
rect 1559 975 1565 976
rect 1559 974 1560 975
rect 1537 972 1560 974
rect 1511 970 1517 971
rect 1559 971 1560 972
rect 1564 971 1565 975
rect 1559 970 1565 971
rect 1607 975 1613 976
rect 1607 971 1608 975
rect 1612 974 1613 975
rect 1632 974 1634 988
rect 1639 987 1640 988
rect 1644 987 1645 991
rect 1639 986 1645 987
rect 1662 980 1668 981
rect 1662 976 1663 980
rect 1667 976 1668 980
rect 1612 972 1634 974
rect 1638 975 1645 976
rect 1662 975 1668 976
rect 1612 971 1613 972
rect 1607 970 1613 971
rect 1638 971 1639 975
rect 1644 971 1645 975
rect 1638 970 1645 971
rect 414 967 420 968
rect 414 966 415 967
rect 288 964 415 966
rect 414 963 415 964
rect 419 963 420 967
rect 674 967 680 968
rect 674 966 675 967
rect 414 962 420 963
rect 489 964 675 966
rect 223 959 229 960
rect 183 955 192 956
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 183 951 184 955
rect 191 951 192 955
rect 215 955 221 956
rect 215 954 216 955
rect 208 952 216 954
rect 110 947 116 948
rect 166 950 172 951
rect 183 950 192 951
rect 198 950 204 951
rect 166 946 167 950
rect 171 946 172 950
rect 166 945 172 946
rect 198 946 199 950
rect 203 946 204 950
rect 198 945 204 946
rect 208 940 210 952
rect 215 951 216 952
rect 220 951 221 955
rect 223 955 224 959
rect 228 958 229 959
rect 263 959 269 960
rect 228 956 250 958
rect 228 955 229 956
rect 223 954 229 955
rect 248 954 250 956
rect 255 955 261 956
rect 255 954 256 955
rect 248 952 256 954
rect 255 951 256 952
rect 260 951 261 955
rect 263 955 264 959
rect 268 958 269 959
rect 311 959 317 960
rect 268 956 307 958
rect 268 955 269 956
rect 263 954 269 955
rect 303 955 309 956
rect 303 951 304 955
rect 308 951 309 955
rect 311 955 312 959
rect 316 958 317 959
rect 367 959 373 960
rect 316 956 354 958
rect 316 955 317 956
rect 311 954 317 955
rect 352 954 354 956
rect 359 955 365 956
rect 359 954 360 955
rect 352 952 360 954
rect 359 951 360 952
rect 364 951 365 955
rect 367 955 368 959
rect 372 958 373 959
rect 372 956 418 958
rect 489 956 491 964
rect 674 963 675 964
rect 679 963 680 967
rect 921 966 923 970
rect 1182 967 1188 968
rect 1182 966 1183 967
rect 921 964 1183 966
rect 674 962 680 963
rect 1182 963 1183 964
rect 1187 963 1188 967
rect 1486 967 1492 968
rect 1486 966 1487 967
rect 1409 964 1487 966
rect 1182 962 1188 963
rect 1322 963 1328 964
rect 495 959 501 960
rect 372 955 373 956
rect 367 954 373 955
rect 416 954 418 956
rect 423 955 429 956
rect 423 954 424 955
rect 416 952 424 954
rect 423 951 424 952
rect 428 951 429 955
rect 487 955 493 956
rect 487 951 488 955
rect 492 951 493 955
rect 495 955 496 959
rect 500 958 501 959
rect 559 959 565 960
rect 500 956 555 958
rect 500 955 501 956
rect 495 954 501 955
rect 551 955 557 956
rect 551 951 552 955
rect 556 951 557 955
rect 559 955 560 959
rect 564 958 565 959
rect 623 959 629 960
rect 564 956 619 958
rect 564 955 565 956
rect 559 954 565 955
rect 615 955 621 956
rect 615 951 616 955
rect 620 951 621 955
rect 623 955 624 959
rect 628 958 629 959
rect 871 959 877 960
rect 628 956 683 958
rect 745 956 802 958
rect 628 955 629 956
rect 623 954 629 955
rect 679 955 685 956
rect 679 951 680 955
rect 684 951 685 955
rect 743 955 749 956
rect 743 951 744 955
rect 748 951 749 955
rect 215 950 221 951
rect 238 950 244 951
rect 255 950 261 951
rect 286 950 292 951
rect 303 950 309 951
rect 342 950 348 951
rect 359 950 365 951
rect 406 950 412 951
rect 423 950 429 951
rect 470 950 476 951
rect 487 950 493 951
rect 534 950 540 951
rect 551 950 557 951
rect 598 950 604 951
rect 615 950 621 951
rect 662 950 668 951
rect 679 950 685 951
rect 726 950 732 951
rect 743 950 749 951
rect 790 950 796 951
rect 238 946 239 950
rect 243 946 244 950
rect 238 945 244 946
rect 286 946 287 950
rect 291 946 292 950
rect 286 945 292 946
rect 342 946 343 950
rect 347 946 348 950
rect 342 945 348 946
rect 406 946 407 950
rect 411 946 412 950
rect 406 945 412 946
rect 470 946 471 950
rect 475 946 476 950
rect 470 945 476 946
rect 534 946 535 950
rect 539 946 540 950
rect 534 945 540 946
rect 598 946 599 950
rect 603 946 604 950
rect 598 945 604 946
rect 662 946 663 950
rect 667 946 668 950
rect 662 945 668 946
rect 726 946 727 950
rect 731 946 732 950
rect 726 945 732 946
rect 790 946 791 950
rect 795 946 796 950
rect 790 945 796 946
rect 183 939 189 940
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 183 935 184 939
rect 188 938 189 939
rect 196 938 210 940
rect 215 939 221 940
rect 188 936 198 938
rect 188 935 189 936
rect 183 934 189 935
rect 215 935 216 939
rect 220 938 221 939
rect 223 939 229 940
rect 223 938 224 939
rect 220 936 224 938
rect 220 935 221 936
rect 215 934 221 935
rect 223 935 224 936
rect 228 935 229 939
rect 223 934 229 935
rect 255 939 261 940
rect 255 935 256 939
rect 260 938 261 939
rect 263 939 269 940
rect 263 938 264 939
rect 260 936 264 938
rect 260 935 261 936
rect 255 934 261 935
rect 263 935 264 936
rect 268 935 269 939
rect 263 934 269 935
rect 303 939 309 940
rect 303 935 304 939
rect 308 938 309 939
rect 311 939 317 940
rect 311 938 312 939
rect 308 936 312 938
rect 308 935 309 936
rect 303 934 309 935
rect 311 935 312 936
rect 316 935 317 939
rect 311 934 317 935
rect 359 939 365 940
rect 359 935 360 939
rect 364 938 365 939
rect 367 939 373 940
rect 367 938 368 939
rect 364 936 368 938
rect 364 935 365 936
rect 359 934 365 935
rect 367 935 368 936
rect 372 935 373 939
rect 367 934 373 935
rect 418 939 429 940
rect 418 935 419 939
rect 423 935 424 939
rect 428 935 429 939
rect 418 934 429 935
rect 487 939 493 940
rect 487 935 488 939
rect 492 938 493 939
rect 495 939 501 940
rect 495 938 496 939
rect 492 936 496 938
rect 492 935 493 936
rect 487 934 493 935
rect 495 935 496 936
rect 500 935 501 939
rect 495 934 501 935
rect 551 939 557 940
rect 551 935 552 939
rect 556 938 557 939
rect 559 939 565 940
rect 559 938 560 939
rect 556 936 560 938
rect 556 935 557 936
rect 551 934 557 935
rect 559 935 560 936
rect 564 935 565 939
rect 559 934 565 935
rect 615 939 621 940
rect 615 935 616 939
rect 620 938 621 939
rect 623 939 629 940
rect 623 938 624 939
rect 620 936 624 938
rect 620 935 621 936
rect 615 934 621 935
rect 623 935 624 936
rect 628 935 629 939
rect 623 934 629 935
rect 674 939 685 940
rect 674 935 675 939
rect 679 935 680 939
rect 684 935 685 939
rect 674 934 685 935
rect 743 939 749 940
rect 743 935 744 939
rect 748 938 749 939
rect 758 939 764 940
rect 758 938 759 939
rect 748 936 759 938
rect 748 935 749 936
rect 743 934 749 935
rect 758 935 759 936
rect 763 935 764 939
rect 800 938 802 956
rect 806 955 813 956
rect 806 951 807 955
rect 812 951 813 955
rect 862 955 869 956
rect 862 951 863 955
rect 868 951 869 955
rect 871 955 872 959
rect 876 958 877 959
rect 935 959 941 960
rect 876 956 922 958
rect 876 955 877 956
rect 871 954 877 955
rect 920 954 922 956
rect 927 955 933 956
rect 927 954 928 955
rect 920 952 928 954
rect 927 951 928 952
rect 932 951 933 955
rect 935 955 936 959
rect 940 958 941 959
rect 999 959 1005 960
rect 940 956 986 958
rect 940 955 941 956
rect 935 954 941 955
rect 984 954 986 956
rect 991 955 997 956
rect 991 954 992 955
rect 984 952 992 954
rect 991 951 992 952
rect 996 951 997 955
rect 999 955 1000 959
rect 1004 958 1005 959
rect 1063 959 1069 960
rect 1004 956 1050 958
rect 1004 955 1005 956
rect 999 954 1005 955
rect 1048 954 1050 956
rect 1055 955 1061 956
rect 1055 954 1056 955
rect 1048 952 1056 954
rect 1055 951 1056 952
rect 1060 951 1061 955
rect 1063 955 1064 959
rect 1068 958 1069 959
rect 1127 959 1133 960
rect 1068 956 1114 958
rect 1068 955 1069 956
rect 1063 954 1069 955
rect 1112 954 1114 956
rect 1119 955 1125 956
rect 1119 954 1120 955
rect 1112 952 1120 954
rect 1119 951 1120 952
rect 1124 951 1125 955
rect 1127 955 1128 959
rect 1132 958 1133 959
rect 1322 959 1323 963
rect 1327 962 1328 963
rect 1327 960 1363 962
rect 1327 959 1328 960
rect 1322 958 1328 959
rect 1132 956 1178 958
rect 1249 956 1298 958
rect 1336 956 1354 958
rect 1361 956 1363 960
rect 1409 956 1411 964
rect 1486 963 1487 964
rect 1491 963 1492 967
rect 1486 962 1492 963
rect 1415 959 1421 960
rect 1132 955 1133 956
rect 1127 954 1133 955
rect 1176 954 1178 956
rect 1183 955 1189 956
rect 1183 954 1184 955
rect 1176 952 1184 954
rect 1183 951 1184 952
rect 1188 951 1189 955
rect 1247 955 1253 956
rect 1247 951 1248 955
rect 1252 951 1253 955
rect 806 950 813 951
rect 846 950 852 951
rect 862 950 869 951
rect 910 950 916 951
rect 927 950 933 951
rect 974 950 980 951
rect 991 950 997 951
rect 1038 950 1044 951
rect 1055 950 1061 951
rect 1102 950 1108 951
rect 1119 950 1125 951
rect 1166 950 1172 951
rect 1183 950 1189 951
rect 1230 950 1236 951
rect 1247 950 1253 951
rect 1286 950 1292 951
rect 846 946 847 950
rect 851 946 852 950
rect 846 945 852 946
rect 910 946 911 950
rect 915 946 916 950
rect 910 945 916 946
rect 974 946 975 950
rect 979 946 980 950
rect 974 945 980 946
rect 1038 946 1039 950
rect 1043 946 1044 950
rect 1038 945 1044 946
rect 1102 946 1103 950
rect 1107 946 1108 950
rect 1102 945 1108 946
rect 1166 946 1167 950
rect 1171 946 1172 950
rect 1166 945 1172 946
rect 1230 946 1231 950
rect 1235 946 1236 950
rect 1230 945 1236 946
rect 1286 946 1287 950
rect 1291 946 1292 950
rect 1286 945 1292 946
rect 807 939 813 940
rect 807 938 808 939
rect 800 936 808 938
rect 758 934 764 935
rect 807 935 808 936
rect 812 935 813 939
rect 807 934 813 935
rect 863 939 869 940
rect 863 935 864 939
rect 868 938 869 939
rect 871 939 877 940
rect 871 938 872 939
rect 868 936 872 938
rect 868 935 869 936
rect 863 934 869 935
rect 871 935 872 936
rect 876 935 877 939
rect 871 934 877 935
rect 927 939 933 940
rect 927 935 928 939
rect 932 938 933 939
rect 935 939 941 940
rect 935 938 936 939
rect 932 936 936 938
rect 932 935 933 936
rect 927 934 933 935
rect 935 935 936 936
rect 940 935 941 939
rect 935 934 941 935
rect 991 939 997 940
rect 991 935 992 939
rect 996 938 997 939
rect 999 939 1005 940
rect 999 938 1000 939
rect 996 936 1000 938
rect 996 935 997 936
rect 991 934 997 935
rect 999 935 1000 936
rect 1004 935 1005 939
rect 999 934 1005 935
rect 1055 939 1061 940
rect 1055 935 1056 939
rect 1060 938 1061 939
rect 1063 939 1069 940
rect 1063 938 1064 939
rect 1060 936 1064 938
rect 1060 935 1061 936
rect 1055 934 1061 935
rect 1063 935 1064 936
rect 1068 935 1069 939
rect 1063 934 1069 935
rect 1119 939 1125 940
rect 1119 935 1120 939
rect 1124 938 1125 939
rect 1127 939 1133 940
rect 1127 938 1128 939
rect 1124 936 1128 938
rect 1124 935 1125 936
rect 1119 934 1125 935
rect 1127 935 1128 936
rect 1132 935 1133 939
rect 1127 934 1133 935
rect 1182 939 1189 940
rect 1182 935 1183 939
rect 1188 935 1189 939
rect 1182 934 1189 935
rect 1247 939 1253 940
rect 1247 935 1248 939
rect 1252 935 1253 939
rect 1296 938 1298 956
rect 1303 955 1309 956
rect 1303 951 1304 955
rect 1308 954 1309 955
rect 1336 954 1338 956
rect 1308 952 1338 954
rect 1308 951 1309 952
rect 1303 950 1309 951
rect 1342 950 1348 951
rect 1342 946 1343 950
rect 1347 946 1348 950
rect 1342 945 1348 946
rect 1352 942 1354 956
rect 1359 955 1365 956
rect 1359 951 1360 955
rect 1364 951 1365 955
rect 1407 955 1413 956
rect 1407 951 1408 955
rect 1412 951 1413 955
rect 1415 955 1416 959
rect 1420 958 1421 959
rect 1420 956 1442 958
rect 1504 956 1522 958
rect 1545 956 1563 958
rect 1616 956 1643 958
rect 1420 955 1421 956
rect 1415 954 1421 955
rect 1440 954 1442 956
rect 1447 955 1453 956
rect 1447 954 1448 955
rect 1440 952 1448 954
rect 1447 951 1448 952
rect 1452 951 1453 955
rect 1487 955 1493 956
rect 1487 951 1488 955
rect 1492 954 1493 955
rect 1504 954 1506 956
rect 1492 952 1506 954
rect 1492 951 1493 952
rect 1359 950 1365 951
rect 1390 950 1396 951
rect 1407 950 1413 951
rect 1430 950 1436 951
rect 1447 950 1453 951
rect 1470 950 1476 951
rect 1487 950 1493 951
rect 1510 950 1516 951
rect 1390 946 1391 950
rect 1395 946 1396 950
rect 1390 945 1396 946
rect 1430 946 1431 950
rect 1435 946 1436 950
rect 1430 945 1436 946
rect 1470 946 1471 950
rect 1475 946 1476 950
rect 1470 945 1476 946
rect 1510 946 1511 950
rect 1515 946 1516 950
rect 1510 945 1516 946
rect 1458 943 1464 944
rect 1458 942 1459 943
rect 1352 940 1363 942
rect 1447 941 1459 942
rect 1303 939 1309 940
rect 1303 938 1304 939
rect 1296 936 1304 938
rect 1247 934 1253 935
rect 1303 935 1304 936
rect 1308 935 1309 939
rect 1303 934 1309 935
rect 1359 939 1365 940
rect 1359 935 1360 939
rect 1364 935 1365 939
rect 1359 934 1365 935
rect 1407 939 1413 940
rect 1407 935 1408 939
rect 1412 938 1413 939
rect 1415 939 1421 940
rect 1415 938 1416 939
rect 1412 936 1416 938
rect 1412 935 1413 936
rect 1407 934 1413 935
rect 1415 935 1416 936
rect 1420 935 1421 939
rect 1447 937 1448 941
rect 1452 940 1459 941
rect 1452 937 1453 940
rect 1458 939 1459 940
rect 1463 939 1464 943
rect 1458 938 1464 939
rect 1486 939 1493 940
rect 1447 936 1453 937
rect 1415 934 1421 935
rect 1486 935 1487 939
rect 1492 935 1493 939
rect 1520 938 1522 956
rect 1527 955 1533 956
rect 1527 951 1528 955
rect 1532 954 1533 955
rect 1545 954 1547 956
rect 1532 952 1547 954
rect 1532 951 1533 952
rect 1527 950 1533 951
rect 1550 950 1556 951
rect 1550 946 1551 950
rect 1555 946 1556 950
rect 1550 945 1556 946
rect 1527 939 1533 940
rect 1527 938 1528 939
rect 1520 936 1528 938
rect 1486 934 1493 935
rect 1527 935 1528 936
rect 1532 935 1533 939
rect 1561 938 1563 956
rect 1567 955 1573 956
rect 1567 951 1568 955
rect 1572 954 1573 955
rect 1582 955 1588 956
rect 1582 954 1583 955
rect 1572 952 1583 954
rect 1572 951 1573 952
rect 1567 950 1573 951
rect 1582 951 1583 952
rect 1587 951 1588 955
rect 1606 955 1613 956
rect 1606 951 1607 955
rect 1612 951 1613 955
rect 1582 950 1588 951
rect 1590 950 1596 951
rect 1606 950 1613 951
rect 1590 946 1591 950
rect 1595 946 1596 950
rect 1590 945 1596 946
rect 1567 939 1573 940
rect 1567 938 1568 939
rect 1561 936 1568 938
rect 1527 934 1533 935
rect 1567 935 1568 936
rect 1572 935 1573 939
rect 1567 934 1573 935
rect 1607 939 1613 940
rect 1607 935 1608 939
rect 1612 938 1613 939
rect 1616 938 1618 956
rect 1639 955 1645 956
rect 1639 951 1640 955
rect 1644 951 1645 955
rect 1622 950 1628 951
rect 1639 950 1645 951
rect 1662 952 1668 953
rect 1622 946 1623 950
rect 1627 946 1628 950
rect 1662 948 1663 952
rect 1667 948 1668 952
rect 1662 947 1668 948
rect 1622 945 1628 946
rect 1612 936 1618 938
rect 1639 939 1645 940
rect 1612 935 1613 936
rect 1607 934 1613 935
rect 1639 935 1640 939
rect 1644 935 1645 939
rect 1639 934 1645 935
rect 1662 935 1668 936
rect 110 930 116 931
rect 166 933 172 934
rect 166 929 167 933
rect 171 929 172 933
rect 166 928 172 929
rect 198 933 204 934
rect 198 929 199 933
rect 203 929 204 933
rect 198 928 204 929
rect 238 933 244 934
rect 238 929 239 933
rect 243 929 244 933
rect 238 928 244 929
rect 286 933 292 934
rect 286 929 287 933
rect 291 929 292 933
rect 286 928 292 929
rect 342 933 348 934
rect 342 929 343 933
rect 347 929 348 933
rect 342 928 348 929
rect 406 933 412 934
rect 406 929 407 933
rect 411 929 412 933
rect 406 928 412 929
rect 470 933 476 934
rect 470 929 471 933
rect 475 929 476 933
rect 470 928 476 929
rect 534 933 540 934
rect 534 929 535 933
rect 539 929 540 933
rect 534 928 540 929
rect 598 933 604 934
rect 598 929 599 933
rect 603 929 604 933
rect 598 928 604 929
rect 662 933 668 934
rect 662 929 663 933
rect 667 929 668 933
rect 662 928 668 929
rect 726 933 732 934
rect 726 929 727 933
rect 731 929 732 933
rect 726 928 732 929
rect 790 933 796 934
rect 790 929 791 933
rect 795 929 796 933
rect 790 928 796 929
rect 846 933 852 934
rect 846 929 847 933
rect 851 929 852 933
rect 846 928 852 929
rect 910 933 916 934
rect 910 929 911 933
rect 915 929 916 933
rect 910 928 916 929
rect 974 933 980 934
rect 974 929 975 933
rect 979 929 980 933
rect 974 928 980 929
rect 1038 933 1044 934
rect 1038 929 1039 933
rect 1043 929 1044 933
rect 1038 928 1044 929
rect 1102 933 1108 934
rect 1102 929 1103 933
rect 1107 929 1108 933
rect 1102 928 1108 929
rect 1166 933 1172 934
rect 1166 929 1167 933
rect 1171 929 1172 933
rect 1166 928 1172 929
rect 1230 933 1236 934
rect 1230 929 1231 933
rect 1235 929 1236 933
rect 1230 928 1236 929
rect 1174 927 1180 928
rect 186 923 192 924
rect 186 919 187 923
rect 191 922 192 923
rect 862 923 868 924
rect 191 920 418 922
rect 191 919 192 920
rect 186 918 192 919
rect 134 915 140 916
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 134 911 135 915
rect 139 911 140 915
rect 134 910 140 911
rect 166 915 172 916
rect 166 911 167 915
rect 171 911 172 915
rect 166 910 172 911
rect 206 915 212 916
rect 206 911 207 915
rect 211 911 212 915
rect 206 910 212 911
rect 270 915 276 916
rect 270 911 271 915
rect 275 911 276 915
rect 270 910 276 911
rect 334 915 340 916
rect 334 911 335 915
rect 339 911 340 915
rect 334 910 340 911
rect 406 915 412 916
rect 406 911 407 915
rect 411 911 412 915
rect 406 910 412 911
rect 110 908 116 909
rect 151 907 157 908
rect 151 903 152 907
rect 156 906 157 907
rect 183 907 189 908
rect 156 904 178 906
rect 156 903 157 904
rect 151 902 157 903
rect 134 898 140 899
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 134 894 135 898
rect 139 894 140 898
rect 134 893 140 894
rect 166 898 172 899
rect 166 894 167 898
rect 171 894 172 898
rect 166 893 172 894
rect 110 891 116 892
rect 151 891 157 892
rect 151 887 152 891
rect 156 887 157 891
rect 176 890 178 904
rect 183 903 184 907
rect 188 906 189 907
rect 223 907 229 908
rect 188 904 218 906
rect 188 903 189 904
rect 183 902 189 903
rect 206 898 212 899
rect 206 894 207 898
rect 211 894 212 898
rect 206 893 212 894
rect 183 891 189 892
rect 183 890 184 891
rect 176 888 184 890
rect 151 886 157 887
rect 183 887 184 888
rect 188 887 189 891
rect 216 890 218 904
rect 223 903 224 907
rect 228 906 229 907
rect 287 907 293 908
rect 228 904 282 906
rect 228 903 229 904
rect 223 902 229 903
rect 270 898 276 899
rect 270 894 271 898
rect 275 894 276 898
rect 270 893 276 894
rect 223 891 229 892
rect 223 890 224 891
rect 216 888 224 890
rect 183 886 189 887
rect 223 887 224 888
rect 228 887 229 891
rect 280 890 282 904
rect 287 903 288 907
rect 292 906 293 907
rect 351 907 357 908
rect 292 904 321 906
rect 292 903 293 904
rect 287 902 293 903
rect 287 891 293 892
rect 287 890 288 891
rect 280 888 288 890
rect 223 886 229 887
rect 287 887 288 888
rect 292 887 293 891
rect 319 890 321 904
rect 351 903 352 907
rect 356 906 357 907
rect 416 906 418 920
rect 862 919 863 923
rect 867 922 868 923
rect 1174 923 1175 927
rect 1179 926 1180 927
rect 1249 926 1251 934
rect 1286 933 1292 934
rect 1286 929 1287 933
rect 1291 929 1292 933
rect 1286 928 1292 929
rect 1342 933 1348 934
rect 1342 929 1343 933
rect 1347 929 1348 933
rect 1342 928 1348 929
rect 1390 933 1396 934
rect 1390 929 1391 933
rect 1395 929 1396 933
rect 1390 928 1396 929
rect 1430 933 1436 934
rect 1430 929 1431 933
rect 1435 929 1436 933
rect 1430 928 1436 929
rect 1470 933 1476 934
rect 1470 929 1471 933
rect 1475 929 1476 933
rect 1470 928 1476 929
rect 1510 933 1516 934
rect 1510 929 1511 933
rect 1515 929 1516 933
rect 1510 928 1516 929
rect 1550 933 1556 934
rect 1550 929 1551 933
rect 1555 929 1556 933
rect 1550 928 1556 929
rect 1590 933 1596 934
rect 1590 929 1591 933
rect 1595 929 1596 933
rect 1590 928 1596 929
rect 1622 933 1628 934
rect 1622 929 1623 933
rect 1627 929 1628 933
rect 1622 928 1628 929
rect 1179 924 1251 926
rect 1582 927 1588 928
rect 1179 923 1180 924
rect 1174 922 1180 923
rect 1582 923 1583 927
rect 1587 926 1588 927
rect 1641 926 1643 934
rect 1662 931 1663 935
rect 1667 931 1668 935
rect 1662 930 1668 931
rect 1587 924 1643 926
rect 1587 923 1588 924
rect 1582 922 1588 923
rect 867 920 1078 922
rect 867 919 868 920
rect 862 918 868 919
rect 470 915 476 916
rect 470 911 471 915
rect 475 911 476 915
rect 470 910 476 911
rect 534 915 540 916
rect 534 911 535 915
rect 539 911 540 915
rect 534 910 540 911
rect 590 915 596 916
rect 590 911 591 915
rect 595 911 596 915
rect 590 910 596 911
rect 646 915 652 916
rect 646 911 647 915
rect 651 911 652 915
rect 646 910 652 911
rect 702 915 708 916
rect 702 911 703 915
rect 707 911 708 915
rect 702 910 708 911
rect 750 915 756 916
rect 750 911 751 915
rect 755 911 756 915
rect 750 910 756 911
rect 798 915 804 916
rect 798 911 799 915
rect 803 911 804 915
rect 798 910 804 911
rect 846 915 852 916
rect 846 911 847 915
rect 851 911 852 915
rect 846 910 852 911
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 958 915 964 916
rect 958 911 959 915
rect 963 911 964 915
rect 958 910 964 911
rect 1022 915 1028 916
rect 1022 911 1023 915
rect 1027 911 1028 915
rect 1022 910 1028 911
rect 423 907 429 908
rect 423 906 424 907
rect 356 904 390 906
rect 416 904 424 906
rect 356 903 357 904
rect 351 902 357 903
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 351 891 357 892
rect 351 890 352 891
rect 319 888 352 890
rect 287 886 293 887
rect 351 887 352 888
rect 356 887 357 891
rect 388 890 390 904
rect 423 903 424 904
rect 428 903 429 907
rect 423 902 429 903
rect 486 907 493 908
rect 486 903 487 907
rect 492 903 493 907
rect 551 907 557 908
rect 551 906 552 907
rect 486 902 493 903
rect 521 904 552 906
rect 406 898 412 899
rect 406 894 407 898
rect 411 894 412 898
rect 406 893 412 894
rect 470 898 476 899
rect 470 894 471 898
rect 475 894 476 898
rect 470 893 476 894
rect 423 891 429 892
rect 423 890 424 891
rect 388 888 424 890
rect 351 886 357 887
rect 423 887 424 888
rect 428 887 429 891
rect 423 886 429 887
rect 487 891 493 892
rect 487 887 488 891
rect 492 890 493 891
rect 521 890 523 904
rect 551 903 552 904
rect 556 903 557 907
rect 607 907 613 908
rect 607 906 608 907
rect 551 902 557 903
rect 584 904 608 906
rect 534 898 540 899
rect 534 894 535 898
rect 539 894 540 898
rect 534 893 540 894
rect 492 888 523 890
rect 551 891 557 892
rect 492 887 493 888
rect 487 886 493 887
rect 551 887 552 891
rect 556 890 557 891
rect 584 890 586 904
rect 607 903 608 904
rect 612 903 613 907
rect 607 902 613 903
rect 663 907 672 908
rect 663 903 664 907
rect 671 903 672 907
rect 719 907 725 908
rect 719 906 720 907
rect 663 902 672 903
rect 692 904 720 906
rect 674 899 680 900
rect 590 898 596 899
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 646 898 652 899
rect 674 898 675 899
rect 646 894 647 898
rect 651 894 652 898
rect 646 893 652 894
rect 656 896 675 898
rect 556 888 586 890
rect 607 891 613 892
rect 556 887 557 888
rect 551 886 557 887
rect 607 887 608 891
rect 612 890 613 891
rect 656 890 658 896
rect 674 895 675 896
rect 679 895 680 899
rect 674 894 680 895
rect 612 888 658 890
rect 663 891 669 892
rect 612 887 613 888
rect 607 886 613 887
rect 663 887 664 891
rect 668 890 669 891
rect 692 890 694 904
rect 719 903 720 904
rect 724 903 725 907
rect 767 907 773 908
rect 767 906 768 907
rect 719 902 725 903
rect 745 904 768 906
rect 702 898 708 899
rect 702 894 703 898
rect 707 894 708 898
rect 702 893 708 894
rect 668 888 694 890
rect 719 891 725 892
rect 668 887 669 888
rect 663 886 669 887
rect 719 887 720 891
rect 724 890 725 891
rect 745 890 747 904
rect 767 903 768 904
rect 772 903 773 907
rect 767 902 773 903
rect 815 907 821 908
rect 815 903 816 907
rect 820 906 821 907
rect 863 907 869 908
rect 820 904 842 906
rect 820 903 821 904
rect 815 902 821 903
rect 750 898 756 899
rect 750 894 751 898
rect 755 894 756 898
rect 750 893 756 894
rect 798 898 804 899
rect 798 894 799 898
rect 803 894 804 898
rect 798 893 804 894
rect 724 888 747 890
rect 758 891 764 892
rect 724 887 725 888
rect 719 886 725 887
rect 758 887 759 891
rect 763 890 764 891
rect 767 891 773 892
rect 767 890 768 891
rect 763 888 768 890
rect 763 887 764 888
rect 758 886 764 887
rect 767 887 768 888
rect 772 887 773 891
rect 767 886 773 887
rect 814 891 821 892
rect 814 887 815 891
rect 820 887 821 891
rect 840 890 842 904
rect 863 903 864 907
rect 868 906 869 907
rect 919 907 925 908
rect 868 904 894 906
rect 868 903 869 904
rect 863 902 869 903
rect 846 898 852 899
rect 846 894 847 898
rect 851 894 852 898
rect 846 893 852 894
rect 863 891 869 892
rect 863 890 864 891
rect 840 888 864 890
rect 814 886 821 887
rect 863 887 864 888
rect 868 887 869 891
rect 892 890 894 904
rect 919 903 920 907
rect 924 906 925 907
rect 975 907 981 908
rect 924 904 970 906
rect 924 903 925 904
rect 919 902 925 903
rect 902 898 908 899
rect 902 894 903 898
rect 907 894 908 898
rect 902 893 908 894
rect 958 898 964 899
rect 958 894 959 898
rect 963 894 964 898
rect 958 893 964 894
rect 919 891 925 892
rect 919 890 920 891
rect 892 888 920 890
rect 863 886 869 887
rect 919 887 920 888
rect 924 887 925 891
rect 968 890 970 904
rect 975 903 976 907
rect 980 906 981 907
rect 1039 907 1045 908
rect 980 904 1034 906
rect 980 903 981 904
rect 975 902 981 903
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 975 891 981 892
rect 975 890 976 891
rect 968 888 976 890
rect 919 886 925 887
rect 975 887 976 888
rect 980 887 981 891
rect 1032 890 1034 904
rect 1039 903 1040 907
rect 1044 906 1045 907
rect 1076 906 1078 920
rect 1086 915 1092 916
rect 1086 911 1087 915
rect 1091 911 1092 915
rect 1086 910 1092 911
rect 1142 915 1148 916
rect 1142 911 1143 915
rect 1147 911 1148 915
rect 1142 910 1148 911
rect 1198 915 1204 916
rect 1198 911 1199 915
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1254 915 1260 916
rect 1254 911 1255 915
rect 1259 911 1260 915
rect 1254 910 1260 911
rect 1318 915 1324 916
rect 1318 911 1319 915
rect 1323 911 1324 915
rect 1318 910 1324 911
rect 1382 915 1388 916
rect 1382 911 1383 915
rect 1387 911 1388 915
rect 1382 910 1388 911
rect 1662 913 1668 914
rect 1662 909 1663 913
rect 1667 909 1668 913
rect 1662 908 1668 909
rect 1103 907 1109 908
rect 1103 906 1104 907
rect 1044 904 1074 906
rect 1076 904 1104 906
rect 1044 903 1045 904
rect 1039 902 1045 903
rect 1039 891 1045 892
rect 1039 890 1040 891
rect 1032 888 1040 890
rect 975 886 981 887
rect 1039 887 1040 888
rect 1044 887 1045 891
rect 1072 890 1074 904
rect 1103 903 1104 904
rect 1108 903 1109 907
rect 1103 902 1109 903
rect 1159 907 1165 908
rect 1159 903 1160 907
rect 1164 906 1165 907
rect 1215 907 1221 908
rect 1164 904 1190 906
rect 1164 903 1165 904
rect 1159 902 1165 903
rect 1086 898 1092 899
rect 1086 894 1087 898
rect 1091 894 1092 898
rect 1086 893 1092 894
rect 1142 898 1148 899
rect 1142 894 1143 898
rect 1147 894 1148 898
rect 1142 893 1148 894
rect 1103 891 1109 892
rect 1103 890 1104 891
rect 1072 888 1104 890
rect 1039 886 1045 887
rect 1103 887 1104 888
rect 1108 887 1109 891
rect 1103 886 1109 887
rect 1159 891 1165 892
rect 1159 887 1160 891
rect 1164 890 1165 891
rect 1174 891 1180 892
rect 1174 890 1175 891
rect 1164 888 1175 890
rect 1164 887 1165 888
rect 1159 886 1165 887
rect 1174 887 1175 888
rect 1179 887 1180 891
rect 1188 890 1190 904
rect 1215 903 1216 907
rect 1220 906 1221 907
rect 1271 907 1277 908
rect 1220 904 1251 906
rect 1220 903 1221 904
rect 1215 902 1221 903
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1215 891 1221 892
rect 1215 890 1216 891
rect 1188 888 1216 890
rect 1174 886 1180 887
rect 1215 887 1216 888
rect 1220 887 1221 891
rect 1249 890 1251 904
rect 1271 903 1272 907
rect 1276 906 1277 907
rect 1335 907 1341 908
rect 1276 904 1306 906
rect 1276 903 1277 904
rect 1271 902 1277 903
rect 1254 898 1260 899
rect 1254 894 1255 898
rect 1259 894 1260 898
rect 1254 893 1260 894
rect 1271 891 1277 892
rect 1271 890 1272 891
rect 1249 888 1272 890
rect 1215 886 1221 887
rect 1271 887 1272 888
rect 1276 887 1277 891
rect 1304 890 1306 904
rect 1335 903 1336 907
rect 1340 906 1341 907
rect 1374 907 1380 908
rect 1340 904 1370 906
rect 1340 903 1341 904
rect 1335 902 1341 903
rect 1318 898 1324 899
rect 1318 894 1319 898
rect 1323 894 1324 898
rect 1318 893 1324 894
rect 1335 891 1341 892
rect 1335 890 1336 891
rect 1304 888 1336 890
rect 1271 886 1277 887
rect 1335 887 1336 888
rect 1340 887 1341 891
rect 1368 890 1370 904
rect 1374 903 1375 907
rect 1379 906 1380 907
rect 1399 907 1405 908
rect 1399 906 1400 907
rect 1379 904 1400 906
rect 1379 903 1380 904
rect 1374 902 1380 903
rect 1399 903 1400 904
rect 1404 903 1405 907
rect 1399 902 1405 903
rect 1382 898 1388 899
rect 1382 894 1383 898
rect 1387 894 1388 898
rect 1382 893 1388 894
rect 1662 896 1668 897
rect 1662 892 1663 896
rect 1667 892 1668 896
rect 1399 891 1405 892
rect 1662 891 1668 892
rect 1399 890 1400 891
rect 1368 888 1400 890
rect 1335 886 1341 887
rect 1399 887 1400 888
rect 1404 887 1405 891
rect 1399 886 1405 887
rect 153 882 155 886
rect 422 883 428 884
rect 422 882 423 883
rect 153 880 423 882
rect 422 879 423 880
rect 427 879 428 883
rect 422 878 428 879
rect 1118 879 1124 880
rect 1118 878 1119 879
rect 985 876 1119 878
rect 558 875 564 876
rect 191 871 197 872
rect 160 868 187 870
rect 150 867 157 868
rect 110 864 116 865
rect 110 860 111 864
rect 115 860 116 864
rect 150 863 151 867
rect 156 863 157 867
rect 110 859 116 860
rect 134 862 140 863
rect 150 862 157 863
rect 134 858 135 862
rect 139 858 140 862
rect 134 857 140 858
rect 151 851 157 852
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 151 847 152 851
rect 156 850 157 851
rect 160 850 162 868
rect 183 867 189 868
rect 183 863 184 867
rect 188 863 189 867
rect 191 867 192 871
rect 196 870 197 871
rect 231 871 237 872
rect 196 868 227 870
rect 196 867 197 868
rect 191 866 197 867
rect 223 867 229 868
rect 223 863 224 867
rect 228 863 229 867
rect 231 867 232 871
rect 236 870 237 871
rect 295 871 301 872
rect 236 868 282 870
rect 236 867 237 868
rect 231 866 237 867
rect 280 866 282 868
rect 287 867 293 868
rect 287 866 288 867
rect 280 864 288 866
rect 287 863 288 864
rect 292 863 293 867
rect 295 867 296 871
rect 300 870 301 871
rect 359 871 365 872
rect 300 868 346 870
rect 300 867 301 868
rect 295 866 301 867
rect 344 866 346 868
rect 351 867 357 868
rect 351 866 352 867
rect 344 864 352 866
rect 351 863 352 864
rect 356 863 357 867
rect 359 867 360 871
rect 364 870 365 871
rect 495 871 501 872
rect 364 868 418 870
rect 364 867 365 868
rect 359 866 365 867
rect 416 866 418 868
rect 423 867 429 868
rect 423 866 424 867
rect 416 864 424 866
rect 423 863 424 864
rect 428 863 429 867
rect 486 867 493 868
rect 486 863 487 867
rect 492 863 493 867
rect 495 867 496 871
rect 500 870 501 871
rect 558 871 559 875
rect 563 874 564 875
rect 563 872 723 874
rect 563 871 564 872
rect 558 870 564 871
rect 500 868 555 870
rect 721 868 723 872
rect 727 871 733 872
rect 500 867 501 868
rect 495 866 501 867
rect 551 867 557 868
rect 551 863 552 867
rect 556 863 557 867
rect 615 867 621 868
rect 615 863 616 867
rect 620 866 621 867
rect 646 867 652 868
rect 646 866 647 867
rect 620 864 647 866
rect 620 863 621 864
rect 166 862 172 863
rect 183 862 189 863
rect 206 862 212 863
rect 223 862 229 863
rect 270 862 276 863
rect 287 862 293 863
rect 334 862 340 863
rect 351 862 357 863
rect 406 862 412 863
rect 423 862 429 863
rect 470 862 476 863
rect 486 862 493 863
rect 534 862 540 863
rect 551 862 557 863
rect 598 862 604 863
rect 615 862 621 863
rect 646 863 647 864
rect 651 863 652 867
rect 666 867 677 868
rect 666 863 667 867
rect 671 863 672 867
rect 676 863 677 867
rect 719 867 725 868
rect 719 863 720 867
rect 724 863 725 867
rect 727 867 728 871
rect 732 870 733 871
rect 732 868 771 870
rect 840 868 859 870
rect 897 868 914 870
rect 921 868 978 870
rect 985 868 987 876
rect 1118 875 1119 876
rect 1123 875 1124 879
rect 1374 879 1380 880
rect 1374 878 1375 879
rect 1118 874 1124 875
rect 1184 876 1375 878
rect 1063 871 1069 872
rect 732 867 733 868
rect 727 866 733 867
rect 767 867 773 868
rect 767 863 768 867
rect 772 863 773 867
rect 815 867 821 868
rect 815 863 816 867
rect 820 866 821 867
rect 840 866 842 868
rect 820 864 842 866
rect 820 863 821 864
rect 646 862 652 863
rect 654 862 660 863
rect 666 862 677 863
rect 702 862 708 863
rect 719 862 725 863
rect 750 862 756 863
rect 767 862 773 863
rect 798 862 804 863
rect 815 862 821 863
rect 846 862 852 863
rect 166 858 167 862
rect 171 858 172 862
rect 166 857 172 858
rect 206 858 207 862
rect 211 858 212 862
rect 206 857 212 858
rect 270 858 271 862
rect 275 858 276 862
rect 270 857 276 858
rect 334 858 335 862
rect 339 858 340 862
rect 334 857 340 858
rect 406 858 407 862
rect 411 858 412 862
rect 406 857 412 858
rect 470 858 471 862
rect 475 858 476 862
rect 470 857 476 858
rect 534 858 535 862
rect 539 858 540 862
rect 534 857 540 858
rect 598 858 599 862
rect 603 858 604 862
rect 598 857 604 858
rect 654 858 655 862
rect 659 858 660 862
rect 654 857 660 858
rect 702 858 703 862
rect 707 858 708 862
rect 702 857 708 858
rect 750 858 751 862
rect 755 858 756 862
rect 750 857 756 858
rect 798 858 799 862
rect 803 858 804 862
rect 798 857 804 858
rect 846 858 847 862
rect 851 858 852 862
rect 846 857 852 858
rect 156 848 162 850
rect 183 851 189 852
rect 156 847 157 848
rect 151 846 157 847
rect 183 847 184 851
rect 188 850 189 851
rect 191 851 197 852
rect 191 850 192 851
rect 188 848 192 850
rect 188 847 189 848
rect 183 846 189 847
rect 191 847 192 848
rect 196 847 197 851
rect 191 846 197 847
rect 223 851 229 852
rect 223 847 224 851
rect 228 850 229 851
rect 231 851 237 852
rect 231 850 232 851
rect 228 848 232 850
rect 228 847 229 848
rect 223 846 229 847
rect 231 847 232 848
rect 236 847 237 851
rect 231 846 237 847
rect 287 851 293 852
rect 287 847 288 851
rect 292 850 293 851
rect 295 851 301 852
rect 295 850 296 851
rect 292 848 296 850
rect 292 847 293 848
rect 287 846 293 847
rect 295 847 296 848
rect 300 847 301 851
rect 295 846 301 847
rect 351 851 357 852
rect 351 847 352 851
rect 356 850 357 851
rect 359 851 365 852
rect 359 850 360 851
rect 356 848 360 850
rect 356 847 357 848
rect 351 846 357 847
rect 359 847 360 848
rect 364 847 365 851
rect 359 846 365 847
rect 422 851 429 852
rect 422 847 423 851
rect 428 847 429 851
rect 422 846 429 847
rect 487 851 493 852
rect 487 847 488 851
rect 492 850 493 851
rect 495 851 501 852
rect 495 850 496 851
rect 492 848 496 850
rect 492 847 493 848
rect 487 846 493 847
rect 495 847 496 848
rect 500 847 501 851
rect 495 846 501 847
rect 551 851 557 852
rect 551 847 552 851
rect 556 847 557 851
rect 551 846 557 847
rect 615 851 624 852
rect 615 847 616 851
rect 623 847 624 851
rect 615 846 624 847
rect 666 851 677 852
rect 666 847 667 851
rect 671 847 672 851
rect 676 847 677 851
rect 666 846 677 847
rect 719 851 725 852
rect 719 847 720 851
rect 724 850 725 851
rect 727 851 733 852
rect 727 850 728 851
rect 724 848 728 850
rect 724 847 725 848
rect 719 846 725 847
rect 727 847 728 848
rect 732 847 733 851
rect 727 846 733 847
rect 767 851 773 852
rect 767 847 768 851
rect 772 847 773 851
rect 767 846 773 847
rect 814 851 821 852
rect 814 847 815 851
rect 820 847 821 851
rect 857 850 859 868
rect 863 867 869 868
rect 863 863 864 867
rect 868 866 869 867
rect 897 866 899 868
rect 868 864 899 866
rect 868 863 869 864
rect 863 862 869 863
rect 902 862 908 863
rect 902 858 903 862
rect 907 858 908 862
rect 902 857 908 858
rect 863 851 869 852
rect 863 850 864 851
rect 857 848 864 850
rect 814 846 821 847
rect 863 847 864 848
rect 868 847 869 851
rect 912 850 914 868
rect 919 867 925 868
rect 919 863 920 867
rect 924 863 925 867
rect 919 862 925 863
rect 966 862 972 863
rect 966 858 967 862
rect 971 858 972 862
rect 966 857 972 858
rect 919 851 925 852
rect 919 850 920 851
rect 912 848 920 850
rect 863 846 869 847
rect 919 847 920 848
rect 924 847 925 851
rect 976 850 978 868
rect 983 867 989 868
rect 983 863 984 867
rect 988 863 989 867
rect 1054 867 1061 868
rect 1054 863 1055 867
rect 1060 863 1061 867
rect 1063 867 1064 871
rect 1068 870 1069 871
rect 1068 868 1114 870
rect 1184 868 1186 876
rect 1374 875 1375 876
rect 1379 875 1380 879
rect 1374 874 1380 875
rect 1191 871 1197 872
rect 1068 867 1069 868
rect 1063 866 1069 867
rect 1112 866 1114 868
rect 1119 867 1125 868
rect 1119 866 1120 867
rect 1112 864 1120 866
rect 1119 863 1120 864
rect 1124 863 1125 867
rect 1183 867 1189 868
rect 1183 863 1184 867
rect 1188 863 1189 867
rect 1191 867 1192 871
rect 1196 870 1197 871
rect 1255 871 1261 872
rect 1196 868 1251 870
rect 1196 867 1197 868
rect 1191 866 1197 867
rect 1247 867 1253 868
rect 1247 863 1248 867
rect 1252 863 1253 867
rect 1255 867 1256 871
rect 1260 870 1261 871
rect 1311 871 1317 872
rect 1260 868 1298 870
rect 1260 867 1261 868
rect 1255 866 1261 867
rect 1296 866 1298 868
rect 1303 867 1309 868
rect 1303 866 1304 867
rect 1296 864 1304 866
rect 1303 863 1304 864
rect 1308 863 1309 867
rect 1311 867 1312 871
rect 1316 870 1317 871
rect 1367 871 1373 872
rect 1316 868 1363 870
rect 1316 867 1317 868
rect 1311 866 1317 867
rect 1359 867 1365 868
rect 1359 863 1360 867
rect 1364 863 1365 867
rect 1367 867 1368 871
rect 1372 870 1373 871
rect 1423 871 1429 872
rect 1372 868 1410 870
rect 1372 867 1373 868
rect 1367 866 1373 867
rect 1408 866 1410 868
rect 1415 867 1421 868
rect 1415 866 1416 867
rect 1408 864 1416 866
rect 1415 863 1416 864
rect 1420 863 1421 867
rect 1423 867 1424 871
rect 1428 870 1429 871
rect 1428 868 1483 870
rect 1428 867 1429 868
rect 1423 866 1429 867
rect 1479 867 1485 868
rect 1479 863 1480 867
rect 1484 863 1485 867
rect 983 862 989 863
rect 1038 862 1044 863
rect 1054 862 1061 863
rect 1102 862 1108 863
rect 1119 862 1125 863
rect 1166 862 1172 863
rect 1183 862 1189 863
rect 1230 862 1236 863
rect 1247 862 1253 863
rect 1286 862 1292 863
rect 1303 862 1309 863
rect 1342 862 1348 863
rect 1359 862 1365 863
rect 1398 862 1404 863
rect 1415 862 1421 863
rect 1462 862 1468 863
rect 1479 862 1485 863
rect 1662 864 1668 865
rect 1038 858 1039 862
rect 1043 858 1044 862
rect 1038 857 1044 858
rect 1102 858 1103 862
rect 1107 858 1108 862
rect 1102 857 1108 858
rect 1166 858 1167 862
rect 1171 858 1172 862
rect 1166 857 1172 858
rect 1230 858 1231 862
rect 1235 858 1236 862
rect 1230 857 1236 858
rect 1286 858 1287 862
rect 1291 858 1292 862
rect 1286 857 1292 858
rect 1342 858 1343 862
rect 1347 858 1348 862
rect 1342 857 1348 858
rect 1398 858 1399 862
rect 1403 858 1404 862
rect 1398 857 1404 858
rect 1462 858 1463 862
rect 1467 858 1468 862
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1462 857 1468 858
rect 983 851 989 852
rect 983 850 984 851
rect 976 848 984 850
rect 919 846 925 847
rect 983 847 984 848
rect 988 847 989 851
rect 983 846 989 847
rect 1055 851 1061 852
rect 1055 847 1056 851
rect 1060 850 1061 851
rect 1063 851 1069 852
rect 1063 850 1064 851
rect 1060 848 1064 850
rect 1060 847 1061 848
rect 1055 846 1061 847
rect 1063 847 1064 848
rect 1068 847 1069 851
rect 1063 846 1069 847
rect 1118 851 1125 852
rect 1118 847 1119 851
rect 1124 847 1125 851
rect 1118 846 1125 847
rect 1183 851 1189 852
rect 1183 847 1184 851
rect 1188 850 1189 851
rect 1191 851 1197 852
rect 1191 850 1192 851
rect 1188 848 1192 850
rect 1188 847 1189 848
rect 1183 846 1189 847
rect 1191 847 1192 848
rect 1196 847 1197 851
rect 1191 846 1197 847
rect 1247 851 1253 852
rect 1247 847 1248 851
rect 1252 850 1253 851
rect 1255 851 1261 852
rect 1255 850 1256 851
rect 1252 848 1256 850
rect 1252 847 1253 848
rect 1247 846 1253 847
rect 1255 847 1256 848
rect 1260 847 1261 851
rect 1255 846 1261 847
rect 1303 851 1309 852
rect 1303 847 1304 851
rect 1308 850 1309 851
rect 1311 851 1317 852
rect 1311 850 1312 851
rect 1308 848 1312 850
rect 1308 847 1309 848
rect 1303 846 1309 847
rect 1311 847 1312 848
rect 1316 847 1317 851
rect 1311 846 1317 847
rect 1359 851 1365 852
rect 1359 847 1360 851
rect 1364 850 1365 851
rect 1367 851 1373 852
rect 1367 850 1368 851
rect 1364 848 1368 850
rect 1364 847 1365 848
rect 1359 846 1365 847
rect 1367 847 1368 848
rect 1372 847 1373 851
rect 1367 846 1373 847
rect 1415 851 1421 852
rect 1415 847 1416 851
rect 1420 850 1421 851
rect 1423 851 1429 852
rect 1423 850 1424 851
rect 1420 848 1424 850
rect 1420 847 1421 848
rect 1415 846 1421 847
rect 1423 847 1424 848
rect 1428 847 1429 851
rect 1423 846 1429 847
rect 1479 851 1485 852
rect 1479 847 1480 851
rect 1484 847 1485 851
rect 1479 846 1485 847
rect 1662 847 1668 848
rect 110 842 116 843
rect 134 845 140 846
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 206 840 212 841
rect 270 845 276 846
rect 270 841 271 845
rect 275 841 276 845
rect 270 840 276 841
rect 334 845 340 846
rect 334 841 335 845
rect 339 841 340 845
rect 334 840 340 841
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 470 845 476 846
rect 470 841 471 845
rect 475 841 476 845
rect 470 840 476 841
rect 534 845 540 846
rect 534 841 535 845
rect 539 841 540 845
rect 534 840 540 841
rect 598 845 604 846
rect 598 841 599 845
rect 603 841 604 845
rect 598 840 604 841
rect 654 845 660 846
rect 654 841 655 845
rect 659 841 660 845
rect 654 840 660 841
rect 702 845 708 846
rect 702 841 703 845
rect 707 841 708 845
rect 702 840 708 841
rect 750 845 756 846
rect 750 841 751 845
rect 755 841 756 845
rect 750 840 756 841
rect 690 839 696 840
rect 690 835 691 839
rect 695 838 696 839
rect 769 838 771 846
rect 798 845 804 846
rect 798 841 799 845
rect 803 841 804 845
rect 798 840 804 841
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 902 845 908 846
rect 902 841 903 845
rect 907 841 908 845
rect 902 840 908 841
rect 966 845 972 846
rect 966 841 967 845
rect 971 841 972 845
rect 966 840 972 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 1102 845 1108 846
rect 1102 841 1103 845
rect 1107 841 1108 845
rect 1102 840 1108 841
rect 1166 845 1172 846
rect 1166 841 1167 845
rect 1171 841 1172 845
rect 1166 840 1172 841
rect 1230 845 1236 846
rect 1230 841 1231 845
rect 1235 841 1236 845
rect 1230 840 1236 841
rect 1286 845 1292 846
rect 1286 841 1287 845
rect 1291 841 1292 845
rect 1286 840 1292 841
rect 1342 845 1348 846
rect 1342 841 1343 845
rect 1347 841 1348 845
rect 1342 840 1348 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1462 845 1468 846
rect 1462 841 1463 845
rect 1467 841 1468 845
rect 1462 840 1468 841
rect 695 836 771 838
rect 1330 839 1336 840
rect 695 835 696 836
rect 690 834 696 835
rect 1330 835 1331 839
rect 1335 838 1336 839
rect 1481 838 1483 846
rect 1662 843 1663 847
rect 1667 843 1668 847
rect 1662 842 1668 843
rect 1335 836 1483 838
rect 1335 835 1336 836
rect 1330 834 1336 835
rect 134 831 140 832
rect 110 829 116 830
rect 110 825 111 829
rect 115 825 116 829
rect 134 827 135 831
rect 139 827 140 831
rect 134 826 140 827
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 214 831 220 832
rect 214 827 215 831
rect 219 827 220 831
rect 214 826 220 827
rect 278 831 284 832
rect 278 827 279 831
rect 283 827 284 831
rect 278 826 284 827
rect 342 831 348 832
rect 342 827 343 831
rect 347 827 348 831
rect 342 826 348 827
rect 414 831 420 832
rect 414 827 415 831
rect 419 827 420 831
rect 414 826 420 827
rect 478 831 484 832
rect 478 827 479 831
rect 483 827 484 831
rect 478 826 484 827
rect 542 831 548 832
rect 542 827 543 831
rect 547 827 548 831
rect 542 826 548 827
rect 606 831 612 832
rect 606 827 607 831
rect 611 827 612 831
rect 606 826 612 827
rect 670 831 676 832
rect 670 827 671 831
rect 675 827 676 831
rect 670 826 676 827
rect 734 831 740 832
rect 734 827 735 831
rect 739 827 740 831
rect 734 826 740 827
rect 790 831 796 832
rect 790 827 791 831
rect 795 827 796 831
rect 790 826 796 827
rect 846 831 852 832
rect 846 827 847 831
rect 851 827 852 831
rect 846 826 852 827
rect 910 831 916 832
rect 910 827 911 831
rect 915 827 916 831
rect 910 826 916 827
rect 974 831 980 832
rect 974 827 975 831
rect 979 827 980 831
rect 974 826 980 827
rect 1038 831 1044 832
rect 1038 827 1039 831
rect 1043 827 1044 831
rect 1038 826 1044 827
rect 1110 831 1116 832
rect 1110 827 1111 831
rect 1115 827 1116 831
rect 1110 826 1116 827
rect 1182 831 1188 832
rect 1182 827 1183 831
rect 1187 827 1188 831
rect 1182 826 1188 827
rect 1246 831 1252 832
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1246 826 1252 827
rect 1310 831 1316 832
rect 1310 827 1311 831
rect 1315 827 1316 831
rect 1310 826 1316 827
rect 1366 831 1372 832
rect 1366 827 1367 831
rect 1371 827 1372 831
rect 1366 826 1372 827
rect 1422 831 1428 832
rect 1422 827 1423 831
rect 1427 827 1428 831
rect 1422 826 1428 827
rect 1478 831 1484 832
rect 1478 827 1479 831
rect 1483 827 1484 831
rect 1478 826 1484 827
rect 1534 831 1540 832
rect 1534 827 1535 831
rect 1539 827 1540 831
rect 1534 826 1540 827
rect 1590 831 1596 832
rect 1590 827 1591 831
rect 1595 827 1596 831
rect 1590 826 1596 827
rect 1662 829 1668 830
rect 110 824 116 825
rect 1662 825 1663 829
rect 1667 825 1668 829
rect 1662 824 1668 825
rect 150 823 157 824
rect 150 819 151 823
rect 156 819 157 823
rect 183 823 189 824
rect 183 822 184 823
rect 150 818 157 819
rect 176 820 184 822
rect 134 814 140 815
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 134 810 135 814
rect 139 810 140 814
rect 134 809 140 810
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 110 807 116 808
rect 151 807 157 808
rect 151 803 152 807
rect 156 806 157 807
rect 176 806 178 820
rect 183 819 184 820
rect 188 819 189 823
rect 231 823 237 824
rect 231 822 232 823
rect 183 818 189 819
rect 208 820 232 822
rect 156 804 178 806
rect 183 807 189 808
rect 156 803 157 804
rect 151 802 157 803
rect 183 803 184 807
rect 188 806 189 807
rect 208 806 210 820
rect 231 819 232 820
rect 236 819 237 823
rect 231 818 237 819
rect 295 823 301 824
rect 295 819 296 823
rect 300 822 301 823
rect 359 823 365 824
rect 300 820 321 822
rect 300 819 301 820
rect 295 818 301 819
rect 214 814 220 815
rect 214 810 215 814
rect 219 810 220 814
rect 214 809 220 810
rect 278 814 284 815
rect 278 810 279 814
rect 283 810 284 814
rect 278 809 284 810
rect 188 804 210 806
rect 231 807 237 808
rect 188 803 189 804
rect 183 802 189 803
rect 231 803 232 807
rect 236 806 237 807
rect 286 807 292 808
rect 236 804 278 806
rect 236 803 237 804
rect 231 802 237 803
rect 276 798 278 804
rect 286 803 287 807
rect 291 806 292 807
rect 295 807 301 808
rect 295 806 296 807
rect 291 804 296 806
rect 291 803 292 804
rect 286 802 292 803
rect 295 803 296 804
rect 300 803 301 807
rect 319 806 321 820
rect 359 819 360 823
rect 364 822 365 823
rect 402 823 408 824
rect 364 820 398 822
rect 364 819 365 820
rect 359 818 365 819
rect 342 814 348 815
rect 342 810 343 814
rect 347 810 348 814
rect 342 809 348 810
rect 359 807 365 808
rect 359 806 360 807
rect 319 804 360 806
rect 295 802 301 803
rect 359 803 360 804
rect 364 803 365 807
rect 396 806 398 820
rect 402 819 403 823
rect 407 822 408 823
rect 431 823 437 824
rect 431 822 432 823
rect 407 820 432 822
rect 407 819 408 820
rect 402 818 408 819
rect 431 819 432 820
rect 436 819 437 823
rect 431 818 437 819
rect 495 823 501 824
rect 495 819 496 823
rect 500 822 501 823
rect 534 823 540 824
rect 534 822 535 823
rect 500 820 535 822
rect 500 819 501 820
rect 495 818 501 819
rect 534 819 535 820
rect 539 819 540 823
rect 559 823 565 824
rect 559 822 560 823
rect 534 818 540 819
rect 552 820 560 822
rect 414 814 420 815
rect 414 810 415 814
rect 419 810 420 814
rect 414 809 420 810
rect 478 814 484 815
rect 478 810 479 814
rect 483 810 484 814
rect 478 809 484 810
rect 542 814 548 815
rect 542 810 543 814
rect 547 810 548 814
rect 542 809 548 810
rect 431 807 437 808
rect 431 806 432 807
rect 396 804 432 806
rect 359 802 365 803
rect 431 803 432 804
rect 436 803 437 807
rect 431 802 437 803
rect 495 807 501 808
rect 495 803 496 807
rect 500 806 501 807
rect 552 806 554 820
rect 559 819 560 820
rect 564 819 565 823
rect 623 823 629 824
rect 623 822 624 823
rect 559 818 565 819
rect 593 820 624 822
rect 500 804 554 806
rect 559 807 565 808
rect 500 803 501 804
rect 495 802 501 803
rect 559 803 560 807
rect 564 806 565 807
rect 593 806 595 820
rect 623 819 624 820
rect 628 819 629 823
rect 623 818 629 819
rect 687 823 693 824
rect 687 819 688 823
rect 692 822 693 823
rect 751 823 757 824
rect 692 820 722 822
rect 692 819 693 820
rect 687 818 693 819
rect 606 814 612 815
rect 606 810 607 814
rect 611 810 612 814
rect 606 809 612 810
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 564 804 595 806
rect 618 807 629 808
rect 564 803 565 804
rect 559 802 565 803
rect 618 803 619 807
rect 623 803 624 807
rect 628 803 629 807
rect 618 802 629 803
rect 687 807 696 808
rect 687 803 688 807
rect 695 803 696 807
rect 720 806 722 820
rect 751 819 752 823
rect 756 822 757 823
rect 807 823 813 824
rect 756 820 782 822
rect 756 819 757 820
rect 751 818 757 819
rect 734 814 740 815
rect 734 810 735 814
rect 739 810 740 814
rect 734 809 740 810
rect 751 807 757 808
rect 751 806 752 807
rect 720 804 752 806
rect 687 802 696 803
rect 751 803 752 804
rect 756 803 757 807
rect 780 806 782 820
rect 807 819 808 823
rect 812 822 813 823
rect 858 823 869 824
rect 812 820 838 822
rect 812 819 813 820
rect 807 818 813 819
rect 790 814 796 815
rect 790 810 791 814
rect 795 810 796 814
rect 790 809 796 810
rect 807 807 813 808
rect 807 806 808 807
rect 780 804 808 806
rect 751 802 757 803
rect 807 803 808 804
rect 812 803 813 807
rect 836 806 838 820
rect 858 819 859 823
rect 863 819 864 823
rect 868 819 869 823
rect 858 818 869 819
rect 927 823 933 824
rect 927 819 928 823
rect 932 822 933 823
rect 991 823 997 824
rect 932 820 962 822
rect 932 819 933 820
rect 927 818 933 819
rect 846 814 852 815
rect 846 810 847 814
rect 851 810 852 814
rect 846 809 852 810
rect 910 814 916 815
rect 910 810 911 814
rect 915 810 916 814
rect 910 809 916 810
rect 863 807 869 808
rect 863 806 864 807
rect 836 804 864 806
rect 807 802 813 803
rect 863 803 864 804
rect 868 803 869 807
rect 863 802 869 803
rect 927 807 933 808
rect 927 803 928 807
rect 932 806 933 807
rect 960 806 962 820
rect 991 819 992 823
rect 996 822 997 823
rect 1054 823 1061 824
rect 996 820 1026 822
rect 996 819 997 820
rect 991 818 997 819
rect 974 814 980 815
rect 974 810 975 814
rect 979 810 980 814
rect 974 809 980 810
rect 991 807 997 808
rect 991 806 992 807
rect 932 804 958 806
rect 960 804 992 806
rect 932 803 933 804
rect 927 802 933 803
rect 402 799 408 800
rect 402 798 403 799
rect 276 796 403 798
rect 402 795 403 796
rect 407 795 408 799
rect 956 798 958 804
rect 991 803 992 804
rect 996 803 997 807
rect 1024 806 1026 820
rect 1054 819 1055 823
rect 1060 819 1061 823
rect 1054 818 1061 819
rect 1063 823 1069 824
rect 1063 819 1064 823
rect 1068 822 1069 823
rect 1127 823 1133 824
rect 1127 822 1128 823
rect 1068 820 1128 822
rect 1068 819 1069 820
rect 1063 818 1069 819
rect 1127 819 1128 820
rect 1132 819 1133 823
rect 1199 823 1205 824
rect 1199 822 1200 823
rect 1127 818 1133 819
rect 1159 820 1200 822
rect 1038 814 1044 815
rect 1038 810 1039 814
rect 1043 810 1044 814
rect 1038 809 1044 810
rect 1110 814 1116 815
rect 1110 810 1111 814
rect 1115 810 1116 814
rect 1110 809 1116 810
rect 1055 807 1061 808
rect 1055 806 1056 807
rect 1024 804 1056 806
rect 991 802 997 803
rect 1055 803 1056 804
rect 1060 803 1061 807
rect 1055 802 1061 803
rect 1127 807 1133 808
rect 1127 803 1128 807
rect 1132 806 1133 807
rect 1159 806 1161 820
rect 1199 819 1200 820
rect 1204 819 1205 823
rect 1263 823 1269 824
rect 1263 822 1264 823
rect 1199 818 1205 819
rect 1233 820 1264 822
rect 1182 814 1188 815
rect 1182 810 1183 814
rect 1187 810 1188 814
rect 1182 809 1188 810
rect 1132 804 1161 806
rect 1199 807 1205 808
rect 1132 803 1133 804
rect 1127 802 1133 803
rect 1199 803 1200 807
rect 1204 806 1205 807
rect 1233 806 1235 820
rect 1263 819 1264 820
rect 1268 819 1269 823
rect 1263 818 1269 819
rect 1327 823 1333 824
rect 1327 819 1328 823
rect 1332 822 1333 823
rect 1383 823 1389 824
rect 1332 820 1358 822
rect 1332 819 1333 820
rect 1327 818 1333 819
rect 1246 814 1252 815
rect 1246 810 1247 814
rect 1251 810 1252 814
rect 1246 809 1252 810
rect 1310 814 1316 815
rect 1310 810 1311 814
rect 1315 810 1316 814
rect 1310 809 1316 810
rect 1204 804 1235 806
rect 1263 807 1269 808
rect 1204 803 1205 804
rect 1199 802 1205 803
rect 1263 803 1264 807
rect 1268 806 1269 807
rect 1302 807 1308 808
rect 1302 806 1303 807
rect 1268 804 1303 806
rect 1268 803 1269 804
rect 1263 802 1269 803
rect 1302 803 1303 804
rect 1307 803 1308 807
rect 1302 802 1308 803
rect 1327 807 1336 808
rect 1327 803 1328 807
rect 1335 803 1336 807
rect 1356 806 1358 820
rect 1383 819 1384 823
rect 1388 822 1389 823
rect 1439 823 1445 824
rect 1388 820 1414 822
rect 1388 819 1389 820
rect 1383 818 1389 819
rect 1366 814 1372 815
rect 1366 810 1367 814
rect 1371 810 1372 814
rect 1366 809 1372 810
rect 1383 807 1389 808
rect 1383 806 1384 807
rect 1356 804 1384 806
rect 1327 802 1336 803
rect 1383 803 1384 804
rect 1388 803 1389 807
rect 1412 806 1414 820
rect 1439 819 1440 823
rect 1444 822 1445 823
rect 1495 823 1501 824
rect 1444 820 1470 822
rect 1444 819 1445 820
rect 1439 818 1445 819
rect 1422 814 1428 815
rect 1422 810 1423 814
rect 1427 810 1428 814
rect 1422 809 1428 810
rect 1439 807 1445 808
rect 1439 806 1440 807
rect 1412 804 1440 806
rect 1383 802 1389 803
rect 1439 803 1440 804
rect 1444 803 1445 807
rect 1468 806 1470 820
rect 1495 819 1496 823
rect 1500 822 1501 823
rect 1551 823 1557 824
rect 1500 820 1546 822
rect 1500 819 1501 820
rect 1495 818 1501 819
rect 1478 814 1484 815
rect 1478 810 1479 814
rect 1483 810 1484 814
rect 1478 809 1484 810
rect 1534 814 1540 815
rect 1534 810 1535 814
rect 1539 810 1540 814
rect 1534 809 1540 810
rect 1495 807 1501 808
rect 1495 806 1496 807
rect 1468 804 1496 806
rect 1439 802 1445 803
rect 1495 803 1496 804
rect 1500 803 1501 807
rect 1544 806 1546 820
rect 1551 819 1552 823
rect 1556 822 1557 823
rect 1606 823 1613 824
rect 1556 820 1582 822
rect 1556 819 1557 820
rect 1551 818 1557 819
rect 1551 807 1557 808
rect 1551 806 1552 807
rect 1544 804 1552 806
rect 1495 802 1501 803
rect 1551 803 1552 804
rect 1556 803 1557 807
rect 1580 806 1582 820
rect 1606 819 1607 823
rect 1612 819 1613 823
rect 1606 818 1613 819
rect 1590 814 1596 815
rect 1590 810 1591 814
rect 1595 810 1596 814
rect 1590 809 1596 810
rect 1662 812 1668 813
rect 1662 808 1663 812
rect 1667 808 1668 812
rect 1607 807 1613 808
rect 1662 807 1668 808
rect 1607 806 1608 807
rect 1580 804 1608 806
rect 1551 802 1557 803
rect 1607 803 1608 804
rect 1612 803 1613 807
rect 1607 802 1613 803
rect 1063 799 1069 800
rect 1063 798 1064 799
rect 956 796 1064 798
rect 402 794 408 795
rect 858 795 864 796
rect 858 794 859 795
rect 720 792 859 794
rect 159 787 165 788
rect 150 783 157 784
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 150 779 151 783
rect 156 779 157 783
rect 159 783 160 787
rect 164 786 165 787
rect 199 787 205 788
rect 164 784 186 786
rect 164 783 165 784
rect 159 782 165 783
rect 184 782 186 784
rect 191 783 197 784
rect 191 782 192 783
rect 184 780 192 782
rect 191 779 192 780
rect 196 779 197 783
rect 199 783 200 787
rect 204 786 205 787
rect 350 787 356 788
rect 204 784 251 786
rect 204 783 205 784
rect 199 782 205 783
rect 247 783 253 784
rect 247 779 248 783
rect 252 779 253 783
rect 306 783 317 784
rect 306 779 307 783
rect 311 779 312 783
rect 316 779 317 783
rect 350 783 351 787
rect 355 786 356 787
rect 391 787 397 788
rect 355 784 387 786
rect 355 783 356 784
rect 350 782 356 783
rect 383 783 389 784
rect 383 779 384 783
rect 388 779 389 783
rect 391 783 392 787
rect 396 786 397 787
rect 551 787 557 788
rect 396 784 458 786
rect 396 783 397 784
rect 391 782 397 783
rect 456 782 458 784
rect 463 783 469 784
rect 463 782 464 783
rect 456 780 464 782
rect 463 779 464 780
rect 468 779 469 783
rect 534 783 540 784
rect 534 779 535 783
rect 539 782 540 783
rect 543 783 549 784
rect 543 782 544 783
rect 539 780 544 782
rect 539 779 540 780
rect 110 775 116 776
rect 134 778 140 779
rect 150 778 157 779
rect 174 778 180 779
rect 191 778 197 779
rect 230 778 236 779
rect 247 778 253 779
rect 294 778 300 779
rect 306 778 317 779
rect 366 778 372 779
rect 383 778 389 779
rect 446 778 452 779
rect 463 778 469 779
rect 526 778 532 779
rect 534 778 540 779
rect 543 779 544 780
rect 548 779 549 783
rect 551 783 552 787
rect 556 786 557 787
rect 556 784 626 786
rect 720 784 722 792
rect 858 791 859 792
rect 863 791 864 795
rect 1063 795 1064 796
rect 1068 795 1069 799
rect 1063 794 1069 795
rect 858 790 864 791
rect 727 787 733 788
rect 556 783 557 784
rect 551 782 557 783
rect 624 782 626 784
rect 631 783 637 784
rect 631 782 632 783
rect 624 780 632 782
rect 631 779 632 780
rect 636 779 637 783
rect 719 783 725 784
rect 719 779 720 783
rect 724 779 725 783
rect 727 783 728 787
rect 732 786 733 787
rect 815 787 821 788
rect 732 784 802 786
rect 732 783 733 784
rect 727 782 733 783
rect 800 782 802 784
rect 807 783 813 784
rect 807 782 808 783
rect 800 780 808 782
rect 807 779 808 780
rect 812 779 813 783
rect 815 783 816 787
rect 820 786 821 787
rect 975 787 981 788
rect 820 784 882 786
rect 820 783 821 784
rect 815 782 821 783
rect 880 782 882 784
rect 887 783 893 784
rect 887 782 888 783
rect 880 780 888 782
rect 887 779 888 780
rect 892 779 893 783
rect 966 783 973 784
rect 966 779 967 783
rect 972 779 973 783
rect 975 783 976 787
rect 980 786 981 787
rect 1047 787 1053 788
rect 980 784 1034 786
rect 980 783 981 784
rect 975 782 981 783
rect 1032 782 1034 784
rect 1039 783 1045 784
rect 1039 782 1040 783
rect 1032 780 1040 782
rect 1039 779 1040 780
rect 1044 779 1045 783
rect 1047 783 1048 787
rect 1052 786 1053 787
rect 1119 787 1125 788
rect 1052 784 1115 786
rect 1052 783 1053 784
rect 1047 782 1053 783
rect 1111 783 1117 784
rect 1111 779 1112 783
rect 1116 779 1117 783
rect 1119 783 1120 787
rect 1124 786 1125 787
rect 1191 787 1197 788
rect 1124 784 1178 786
rect 1124 783 1125 784
rect 1119 782 1125 783
rect 1176 782 1178 784
rect 1183 783 1189 784
rect 1183 782 1184 783
rect 1176 780 1184 782
rect 1183 779 1184 780
rect 1188 779 1189 783
rect 1191 783 1192 787
rect 1196 786 1197 787
rect 1255 787 1261 788
rect 1196 784 1251 786
rect 1196 783 1197 784
rect 1191 782 1197 783
rect 1247 783 1253 784
rect 1247 779 1248 783
rect 1252 779 1253 783
rect 1255 783 1256 787
rect 1260 786 1261 787
rect 1383 787 1389 788
rect 1260 784 1306 786
rect 1260 783 1261 784
rect 1255 782 1261 783
rect 1304 782 1306 784
rect 1311 783 1317 784
rect 1311 782 1312 783
rect 1304 780 1312 782
rect 1311 779 1312 780
rect 1316 779 1317 783
rect 1374 783 1381 784
rect 1374 779 1375 783
rect 1380 779 1381 783
rect 1383 783 1384 787
rect 1388 786 1389 787
rect 1439 787 1445 788
rect 1388 784 1426 786
rect 1388 783 1389 784
rect 1383 782 1389 783
rect 1424 782 1426 784
rect 1431 783 1437 784
rect 1431 782 1432 783
rect 1424 780 1432 782
rect 1431 779 1432 780
rect 1436 779 1437 783
rect 1439 783 1440 787
rect 1444 786 1445 787
rect 1444 784 1482 786
rect 1545 784 1602 786
rect 1444 783 1445 784
rect 1439 782 1445 783
rect 1480 782 1482 784
rect 1487 783 1493 784
rect 1487 782 1488 783
rect 1480 780 1488 782
rect 1487 779 1488 780
rect 1492 779 1493 783
rect 1543 783 1549 784
rect 1543 779 1544 783
rect 1548 779 1549 783
rect 543 778 549 779
rect 614 778 620 779
rect 631 778 637 779
rect 702 778 708 779
rect 719 778 725 779
rect 790 778 796 779
rect 807 778 813 779
rect 870 778 876 779
rect 887 778 893 779
rect 950 778 956 779
rect 966 778 973 779
rect 1022 778 1028 779
rect 1039 778 1045 779
rect 1094 778 1100 779
rect 1111 778 1117 779
rect 1166 778 1172 779
rect 1183 778 1189 779
rect 1230 778 1236 779
rect 1247 778 1253 779
rect 1294 778 1300 779
rect 1311 778 1317 779
rect 1358 778 1364 779
rect 1374 778 1381 779
rect 1414 778 1420 779
rect 1431 778 1437 779
rect 1470 778 1476 779
rect 1487 778 1493 779
rect 1526 778 1532 779
rect 1543 778 1549 779
rect 1590 778 1596 779
rect 134 774 135 778
rect 139 774 140 778
rect 134 773 140 774
rect 174 774 175 778
rect 179 774 180 778
rect 174 773 180 774
rect 230 774 231 778
rect 235 774 236 778
rect 230 773 236 774
rect 294 774 295 778
rect 299 774 300 778
rect 294 773 300 774
rect 366 774 367 778
rect 371 774 372 778
rect 366 773 372 774
rect 446 774 447 778
rect 451 774 452 778
rect 446 773 452 774
rect 526 774 527 778
rect 531 774 532 778
rect 526 773 532 774
rect 614 774 615 778
rect 619 774 620 778
rect 614 773 620 774
rect 702 774 703 778
rect 707 774 708 778
rect 702 773 708 774
rect 790 774 791 778
rect 795 774 796 778
rect 790 773 796 774
rect 870 774 871 778
rect 875 774 876 778
rect 870 773 876 774
rect 950 774 951 778
rect 955 774 956 778
rect 950 773 956 774
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1022 773 1028 774
rect 1094 774 1095 778
rect 1099 774 1100 778
rect 1094 773 1100 774
rect 1166 774 1167 778
rect 1171 774 1172 778
rect 1166 773 1172 774
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1230 773 1236 774
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1294 773 1300 774
rect 1358 774 1359 778
rect 1363 774 1364 778
rect 1358 773 1364 774
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1414 773 1420 774
rect 1470 774 1471 778
rect 1475 774 1476 778
rect 1470 773 1476 774
rect 1526 774 1527 778
rect 1531 774 1532 778
rect 1526 773 1532 774
rect 1590 774 1591 778
rect 1595 774 1596 778
rect 1590 773 1596 774
rect 151 767 157 768
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 151 763 152 767
rect 156 766 157 767
rect 159 767 165 768
rect 159 766 160 767
rect 156 764 160 766
rect 156 763 157 764
rect 151 762 157 763
rect 159 763 160 764
rect 164 763 165 767
rect 159 762 165 763
rect 191 767 197 768
rect 191 763 192 767
rect 196 766 197 767
rect 199 767 205 768
rect 199 766 200 767
rect 196 764 200 766
rect 196 763 197 764
rect 191 762 197 763
rect 199 763 200 764
rect 204 763 205 767
rect 199 762 205 763
rect 247 767 253 768
rect 247 763 248 767
rect 252 766 253 767
rect 286 767 292 768
rect 286 766 287 767
rect 252 764 287 766
rect 252 763 253 764
rect 247 762 253 763
rect 286 763 287 764
rect 291 763 292 767
rect 286 762 292 763
rect 311 767 317 768
rect 311 763 312 767
rect 316 766 317 767
rect 350 767 356 768
rect 350 766 351 767
rect 316 764 351 766
rect 316 763 317 764
rect 311 762 317 763
rect 350 763 351 764
rect 355 763 356 767
rect 350 762 356 763
rect 383 767 389 768
rect 383 763 384 767
rect 388 766 389 767
rect 391 767 397 768
rect 391 766 392 767
rect 388 764 392 766
rect 388 763 389 764
rect 383 762 389 763
rect 391 763 392 764
rect 396 763 397 767
rect 463 767 469 768
rect 463 766 464 767
rect 391 762 397 763
rect 456 764 464 766
rect 110 758 116 759
rect 134 761 140 762
rect 134 757 135 761
rect 139 757 140 761
rect 134 756 140 757
rect 174 761 180 762
rect 174 757 175 761
rect 179 757 180 761
rect 174 756 180 757
rect 230 761 236 762
rect 230 757 231 761
rect 235 757 236 761
rect 230 756 236 757
rect 294 761 300 762
rect 294 757 295 761
rect 299 757 300 761
rect 294 756 300 757
rect 366 761 372 762
rect 366 757 367 761
rect 371 757 372 761
rect 366 756 372 757
rect 446 761 452 762
rect 446 757 447 761
rect 451 757 452 761
rect 446 756 452 757
rect 150 755 156 756
rect 150 751 151 755
rect 155 754 156 755
rect 456 754 458 764
rect 463 763 464 764
rect 468 763 469 767
rect 463 762 469 763
rect 543 767 549 768
rect 543 763 544 767
rect 548 766 549 767
rect 551 767 557 768
rect 551 766 552 767
rect 548 764 552 766
rect 548 763 549 764
rect 543 762 549 763
rect 551 763 552 764
rect 556 763 557 767
rect 551 762 557 763
rect 631 767 637 768
rect 631 763 632 767
rect 636 766 637 767
rect 686 767 692 768
rect 686 766 687 767
rect 636 764 687 766
rect 636 763 637 764
rect 631 762 637 763
rect 686 763 687 764
rect 691 763 692 767
rect 686 762 692 763
rect 719 767 725 768
rect 719 763 720 767
rect 724 766 725 767
rect 727 767 733 768
rect 727 766 728 767
rect 724 764 728 766
rect 724 763 725 764
rect 719 762 725 763
rect 727 763 728 764
rect 732 763 733 767
rect 727 762 733 763
rect 807 767 813 768
rect 807 763 808 767
rect 812 766 813 767
rect 815 767 821 768
rect 815 766 816 767
rect 812 764 816 766
rect 812 763 813 764
rect 807 762 813 763
rect 815 763 816 764
rect 820 763 821 767
rect 815 762 821 763
rect 882 767 893 768
rect 882 763 883 767
rect 887 763 888 767
rect 892 763 893 767
rect 882 762 893 763
rect 967 767 973 768
rect 967 763 968 767
rect 972 766 973 767
rect 975 767 981 768
rect 975 766 976 767
rect 972 764 976 766
rect 972 763 973 764
rect 967 762 973 763
rect 975 763 976 764
rect 980 763 981 767
rect 975 762 981 763
rect 1039 767 1045 768
rect 1039 763 1040 767
rect 1044 766 1045 767
rect 1047 767 1053 768
rect 1047 766 1048 767
rect 1044 764 1048 766
rect 1044 763 1045 764
rect 1039 762 1045 763
rect 1047 763 1048 764
rect 1052 763 1053 767
rect 1047 762 1053 763
rect 1111 767 1117 768
rect 1111 763 1112 767
rect 1116 766 1117 767
rect 1119 767 1125 768
rect 1119 766 1120 767
rect 1116 764 1120 766
rect 1116 763 1117 764
rect 1111 762 1117 763
rect 1119 763 1120 764
rect 1124 763 1125 767
rect 1119 762 1125 763
rect 1183 767 1189 768
rect 1183 763 1184 767
rect 1188 766 1189 767
rect 1191 767 1197 768
rect 1191 766 1192 767
rect 1188 764 1192 766
rect 1188 763 1189 764
rect 1183 762 1189 763
rect 1191 763 1192 764
rect 1196 763 1197 767
rect 1191 762 1197 763
rect 1247 767 1253 768
rect 1247 763 1248 767
rect 1252 766 1253 767
rect 1255 767 1261 768
rect 1255 766 1256 767
rect 1252 764 1256 766
rect 1252 763 1253 764
rect 1247 762 1253 763
rect 1255 763 1256 764
rect 1260 763 1261 767
rect 1255 762 1261 763
rect 1306 767 1317 768
rect 1306 763 1307 767
rect 1311 763 1312 767
rect 1316 763 1317 767
rect 1306 762 1317 763
rect 1375 767 1381 768
rect 1375 763 1376 767
rect 1380 766 1381 767
rect 1383 767 1389 768
rect 1383 766 1384 767
rect 1380 764 1384 766
rect 1380 763 1381 764
rect 1375 762 1381 763
rect 1383 763 1384 764
rect 1388 763 1389 767
rect 1383 762 1389 763
rect 1431 767 1437 768
rect 1431 763 1432 767
rect 1436 766 1437 767
rect 1439 767 1445 768
rect 1439 766 1440 767
rect 1436 764 1440 766
rect 1436 763 1437 764
rect 1431 762 1437 763
rect 1439 763 1440 764
rect 1444 763 1445 767
rect 1439 762 1445 763
rect 1487 767 1493 768
rect 1487 763 1488 767
rect 1492 766 1493 767
rect 1510 767 1516 768
rect 1510 766 1511 767
rect 1492 764 1511 766
rect 1492 763 1493 764
rect 1487 762 1493 763
rect 1510 763 1511 764
rect 1515 763 1516 767
rect 1510 762 1516 763
rect 1543 767 1549 768
rect 1543 763 1544 767
rect 1548 763 1549 767
rect 1600 766 1602 784
rect 1606 783 1613 784
rect 1606 779 1607 783
rect 1612 779 1613 783
rect 1606 778 1613 779
rect 1662 780 1668 781
rect 1662 776 1663 780
rect 1667 776 1668 780
rect 1662 775 1668 776
rect 1607 767 1613 768
rect 1607 766 1608 767
rect 1600 764 1608 766
rect 1543 762 1549 763
rect 1607 763 1608 764
rect 1612 763 1613 767
rect 1607 762 1613 763
rect 1662 763 1668 764
rect 526 761 532 762
rect 526 757 527 761
rect 531 757 532 761
rect 526 756 532 757
rect 614 761 620 762
rect 614 757 615 761
rect 619 757 620 761
rect 614 756 620 757
rect 702 761 708 762
rect 702 757 703 761
rect 707 757 708 761
rect 702 756 708 757
rect 790 761 796 762
rect 790 757 791 761
rect 795 757 796 761
rect 790 756 796 757
rect 870 761 876 762
rect 870 757 871 761
rect 875 757 876 761
rect 870 756 876 757
rect 950 761 956 762
rect 950 757 951 761
rect 955 757 956 761
rect 950 756 956 757
rect 1022 761 1028 762
rect 1022 757 1023 761
rect 1027 757 1028 761
rect 1022 756 1028 757
rect 1094 761 1100 762
rect 1094 757 1095 761
rect 1099 757 1100 761
rect 1094 756 1100 757
rect 1166 761 1172 762
rect 1166 757 1167 761
rect 1171 757 1172 761
rect 1166 756 1172 757
rect 1230 761 1236 762
rect 1230 757 1231 761
rect 1235 757 1236 761
rect 1230 756 1236 757
rect 1294 761 1300 762
rect 1294 757 1295 761
rect 1299 757 1300 761
rect 1294 756 1300 757
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 1526 761 1532 762
rect 1526 757 1527 761
rect 1531 757 1532 761
rect 1526 756 1532 757
rect 155 752 458 754
rect 966 755 972 756
rect 155 751 156 752
rect 150 750 156 751
rect 966 751 967 755
rect 971 754 972 755
rect 1374 755 1380 756
rect 971 752 1179 754
rect 971 751 972 752
rect 966 750 972 751
rect 214 747 220 748
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 246 747 252 748
rect 246 743 247 747
rect 251 743 252 747
rect 246 742 252 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 318 747 324 748
rect 278 742 284 743
rect 306 743 312 744
rect 306 742 307 743
rect 110 740 116 741
rect 295 741 307 742
rect 231 739 237 740
rect 231 735 232 739
rect 236 738 237 739
rect 263 739 269 740
rect 236 736 258 738
rect 236 735 237 736
rect 231 734 237 735
rect 214 730 220 731
rect 110 728 116 729
rect 110 724 111 728
rect 115 724 116 728
rect 214 726 215 730
rect 219 726 220 730
rect 214 725 220 726
rect 246 730 252 731
rect 246 726 247 730
rect 251 726 252 730
rect 246 725 252 726
rect 110 723 116 724
rect 231 723 237 724
rect 231 719 232 723
rect 236 722 237 723
rect 256 722 258 736
rect 263 735 264 739
rect 268 738 269 739
rect 268 736 290 738
rect 295 737 296 741
rect 300 740 307 741
rect 300 737 301 740
rect 306 739 307 740
rect 311 739 312 743
rect 318 743 319 747
rect 323 743 324 747
rect 318 742 324 743
rect 358 747 364 748
rect 358 743 359 747
rect 363 743 364 747
rect 358 742 364 743
rect 398 747 404 748
rect 398 743 399 747
rect 403 743 404 747
rect 398 742 404 743
rect 438 747 444 748
rect 438 743 439 747
rect 443 743 444 747
rect 438 742 444 743
rect 486 747 492 748
rect 486 743 487 747
rect 491 743 492 747
rect 486 742 492 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 606 747 612 748
rect 606 743 607 747
rect 611 743 612 747
rect 606 742 612 743
rect 670 747 676 748
rect 670 743 671 747
rect 675 743 676 747
rect 670 742 676 743
rect 734 747 740 748
rect 734 743 735 747
rect 739 743 740 747
rect 734 742 740 743
rect 798 747 804 748
rect 798 743 799 747
rect 803 743 804 747
rect 798 742 804 743
rect 862 747 868 748
rect 862 743 863 747
rect 867 743 868 747
rect 862 742 868 743
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 990 747 996 748
rect 990 743 991 747
rect 995 743 996 747
rect 990 742 996 743
rect 1054 747 1060 748
rect 1054 743 1055 747
rect 1059 743 1060 747
rect 1054 742 1060 743
rect 1118 747 1124 748
rect 1118 743 1119 747
rect 1123 743 1124 747
rect 1118 742 1124 743
rect 306 738 312 739
rect 330 739 341 740
rect 295 736 301 737
rect 268 735 269 736
rect 263 734 269 735
rect 278 730 284 731
rect 278 726 279 730
rect 283 726 284 730
rect 278 725 284 726
rect 263 723 269 724
rect 263 722 264 723
rect 236 720 254 722
rect 256 720 264 722
rect 236 719 237 720
rect 231 718 237 719
rect 252 714 254 720
rect 263 719 264 720
rect 268 719 269 723
rect 288 722 290 736
rect 330 735 331 739
rect 335 735 336 739
rect 340 735 341 739
rect 330 734 341 735
rect 375 739 381 740
rect 375 735 376 739
rect 380 738 381 739
rect 414 739 421 740
rect 380 736 394 738
rect 380 735 381 736
rect 375 734 381 735
rect 318 730 324 731
rect 318 726 319 730
rect 323 726 324 730
rect 318 725 324 726
rect 358 730 364 731
rect 358 726 359 730
rect 363 726 364 730
rect 358 725 364 726
rect 295 723 301 724
rect 295 722 296 723
rect 288 720 296 722
rect 263 718 269 719
rect 295 719 296 720
rect 300 719 301 723
rect 295 718 301 719
rect 335 723 341 724
rect 335 719 336 723
rect 340 722 341 723
rect 366 723 372 724
rect 340 720 362 722
rect 340 719 341 720
rect 335 718 341 719
rect 330 715 336 716
rect 330 714 331 715
rect 252 712 331 714
rect 330 711 331 712
rect 335 711 336 715
rect 360 714 362 720
rect 366 719 367 723
rect 371 722 372 723
rect 375 723 381 724
rect 375 722 376 723
rect 371 720 376 722
rect 371 719 372 720
rect 366 718 372 719
rect 375 719 376 720
rect 380 719 381 723
rect 392 722 394 736
rect 414 735 415 739
rect 420 735 421 739
rect 414 734 421 735
rect 455 739 461 740
rect 455 735 456 739
rect 460 738 461 739
rect 463 739 469 740
rect 463 738 464 739
rect 460 736 464 738
rect 460 735 461 736
rect 455 734 461 735
rect 463 735 464 736
rect 468 735 469 739
rect 503 739 509 740
rect 503 738 504 739
rect 463 734 469 735
rect 480 736 504 738
rect 398 730 404 731
rect 398 726 399 730
rect 403 726 404 730
rect 398 725 404 726
rect 438 730 444 731
rect 438 726 439 730
rect 443 726 444 730
rect 438 725 444 726
rect 415 723 421 724
rect 415 722 416 723
rect 392 720 416 722
rect 375 718 381 719
rect 415 719 416 720
rect 420 719 421 723
rect 415 718 421 719
rect 455 723 461 724
rect 455 719 456 723
rect 460 722 461 723
rect 480 722 482 736
rect 503 735 504 736
rect 508 735 509 739
rect 559 739 565 740
rect 559 738 560 739
rect 503 734 509 735
rect 536 736 560 738
rect 486 730 492 731
rect 486 726 487 730
rect 491 726 492 730
rect 486 725 492 726
rect 460 720 482 722
rect 503 723 509 724
rect 460 719 461 720
rect 455 718 461 719
rect 503 719 504 723
rect 508 722 509 723
rect 536 722 538 736
rect 559 735 560 736
rect 564 735 565 739
rect 623 739 629 740
rect 623 738 624 739
rect 559 734 565 735
rect 593 736 624 738
rect 542 730 548 731
rect 542 726 543 730
rect 547 726 548 730
rect 542 725 548 726
rect 508 720 538 722
rect 559 723 565 724
rect 508 719 509 720
rect 503 718 509 719
rect 559 719 560 723
rect 564 722 565 723
rect 593 722 595 736
rect 623 735 624 736
rect 628 735 629 739
rect 687 739 693 740
rect 687 738 688 739
rect 623 734 629 735
rect 657 736 688 738
rect 606 730 612 731
rect 606 726 607 730
rect 611 726 612 730
rect 606 725 612 726
rect 564 720 595 722
rect 623 723 629 724
rect 564 719 565 720
rect 559 718 565 719
rect 623 719 624 723
rect 628 722 629 723
rect 657 722 659 736
rect 687 735 688 736
rect 692 735 693 739
rect 687 734 693 735
rect 751 739 757 740
rect 751 735 752 739
rect 756 738 757 739
rect 774 739 780 740
rect 774 738 775 739
rect 756 736 775 738
rect 756 735 757 736
rect 751 734 757 735
rect 774 735 775 736
rect 779 735 780 739
rect 815 739 821 740
rect 815 738 816 739
rect 774 734 780 735
rect 785 736 816 738
rect 670 730 676 731
rect 670 726 671 730
rect 675 726 676 730
rect 670 725 676 726
rect 734 730 740 731
rect 734 726 735 730
rect 739 726 740 730
rect 734 725 740 726
rect 628 720 659 722
rect 686 723 693 724
rect 628 719 629 720
rect 623 718 629 719
rect 686 719 687 723
rect 692 719 693 723
rect 686 718 693 719
rect 751 723 757 724
rect 751 719 752 723
rect 756 722 757 723
rect 785 722 787 736
rect 815 735 816 736
rect 820 735 821 739
rect 879 739 885 740
rect 879 738 880 739
rect 815 734 821 735
rect 852 736 880 738
rect 798 730 804 731
rect 798 726 799 730
rect 803 726 804 730
rect 798 725 804 726
rect 756 720 787 722
rect 815 723 821 724
rect 756 719 757 720
rect 751 718 757 719
rect 815 719 816 723
rect 820 722 821 723
rect 852 722 854 736
rect 879 735 880 736
rect 884 735 885 739
rect 879 734 885 735
rect 943 739 949 740
rect 943 735 944 739
rect 948 738 949 739
rect 1007 739 1013 740
rect 948 736 987 738
rect 948 735 949 736
rect 943 734 949 735
rect 862 730 868 731
rect 862 726 863 730
rect 867 726 868 730
rect 862 725 868 726
rect 926 730 932 731
rect 926 726 927 730
rect 931 726 932 730
rect 926 725 932 726
rect 820 720 854 722
rect 879 723 888 724
rect 820 719 821 720
rect 815 718 821 719
rect 879 719 880 723
rect 887 719 888 723
rect 879 718 888 719
rect 943 723 949 724
rect 943 719 944 723
rect 948 722 949 723
rect 974 723 980 724
rect 974 722 975 723
rect 948 720 975 722
rect 948 719 949 720
rect 943 718 949 719
rect 974 719 975 720
rect 979 719 980 723
rect 985 722 987 736
rect 1007 735 1008 739
rect 1012 738 1013 739
rect 1071 739 1077 740
rect 1012 736 1042 738
rect 1012 735 1013 736
rect 1007 734 1013 735
rect 990 730 996 731
rect 990 726 991 730
rect 995 726 996 730
rect 990 725 996 726
rect 1007 723 1013 724
rect 1007 722 1008 723
rect 985 720 1008 722
rect 974 718 980 719
rect 1007 719 1008 720
rect 1012 719 1013 723
rect 1040 722 1042 736
rect 1071 735 1072 739
rect 1076 738 1077 739
rect 1135 739 1141 740
rect 1076 736 1106 738
rect 1076 735 1077 736
rect 1071 734 1077 735
rect 1054 730 1060 731
rect 1054 726 1055 730
rect 1059 726 1060 730
rect 1054 725 1060 726
rect 1071 723 1077 724
rect 1071 722 1072 723
rect 1040 720 1072 722
rect 1007 718 1013 719
rect 1071 719 1072 720
rect 1076 719 1077 723
rect 1104 722 1106 736
rect 1135 735 1136 739
rect 1140 738 1141 739
rect 1177 738 1179 752
rect 1374 751 1375 755
rect 1379 754 1380 755
rect 1545 754 1547 762
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1662 759 1663 763
rect 1667 759 1668 763
rect 1662 758 1668 759
rect 1590 756 1596 757
rect 1379 752 1547 754
rect 1379 751 1380 752
rect 1374 750 1380 751
rect 1182 747 1188 748
rect 1182 743 1183 747
rect 1187 743 1188 747
rect 1182 742 1188 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 743 1244 747
rect 1238 742 1244 743
rect 1294 747 1300 748
rect 1294 743 1295 747
rect 1299 743 1300 747
rect 1294 742 1300 743
rect 1350 747 1356 748
rect 1350 743 1351 747
rect 1355 743 1356 747
rect 1350 742 1356 743
rect 1406 747 1412 748
rect 1406 743 1407 747
rect 1411 743 1412 747
rect 1406 742 1412 743
rect 1462 747 1468 748
rect 1462 743 1463 747
rect 1467 743 1468 747
rect 1462 742 1468 743
rect 1518 747 1524 748
rect 1518 743 1519 747
rect 1523 743 1524 747
rect 1518 742 1524 743
rect 1582 747 1588 748
rect 1582 743 1583 747
rect 1587 743 1588 747
rect 1582 742 1588 743
rect 1622 747 1628 748
rect 1622 743 1623 747
rect 1627 743 1628 747
rect 1622 742 1628 743
rect 1662 745 1668 746
rect 1662 741 1663 745
rect 1667 741 1668 745
rect 1662 740 1668 741
rect 1199 739 1205 740
rect 1199 738 1200 739
rect 1140 736 1161 738
rect 1177 736 1200 738
rect 1140 735 1141 736
rect 1135 734 1141 735
rect 1118 730 1124 731
rect 1118 726 1119 730
rect 1123 726 1124 730
rect 1118 725 1124 726
rect 1135 723 1141 724
rect 1135 722 1136 723
rect 1104 720 1136 722
rect 1071 718 1077 719
rect 1135 719 1136 720
rect 1140 719 1141 723
rect 1159 722 1161 736
rect 1199 735 1200 736
rect 1204 735 1205 739
rect 1199 734 1205 735
rect 1207 739 1213 740
rect 1207 735 1208 739
rect 1212 738 1213 739
rect 1255 739 1261 740
rect 1255 738 1256 739
rect 1212 736 1256 738
rect 1212 735 1213 736
rect 1207 734 1213 735
rect 1255 735 1256 736
rect 1260 735 1261 739
rect 1311 739 1317 740
rect 1311 738 1312 739
rect 1255 734 1261 735
rect 1288 736 1312 738
rect 1182 730 1188 731
rect 1182 726 1183 730
rect 1187 726 1188 730
rect 1182 725 1188 726
rect 1238 730 1244 731
rect 1238 726 1239 730
rect 1243 726 1244 730
rect 1238 725 1244 726
rect 1199 723 1205 724
rect 1199 722 1200 723
rect 1159 720 1200 722
rect 1135 718 1141 719
rect 1199 719 1200 720
rect 1204 719 1205 723
rect 1199 718 1205 719
rect 1255 723 1261 724
rect 1255 719 1256 723
rect 1260 722 1261 723
rect 1288 722 1290 736
rect 1311 735 1312 736
rect 1316 735 1317 739
rect 1367 739 1373 740
rect 1367 738 1368 739
rect 1311 734 1317 735
rect 1344 736 1368 738
rect 1294 730 1300 731
rect 1294 726 1295 730
rect 1299 726 1300 730
rect 1294 725 1300 726
rect 1260 720 1290 722
rect 1311 723 1317 724
rect 1260 719 1261 720
rect 1255 718 1261 719
rect 1311 719 1312 723
rect 1316 722 1317 723
rect 1344 722 1346 736
rect 1367 735 1368 736
rect 1372 735 1373 739
rect 1423 739 1429 740
rect 1423 738 1424 739
rect 1367 734 1373 735
rect 1396 736 1424 738
rect 1350 730 1356 731
rect 1350 726 1351 730
rect 1355 726 1356 730
rect 1350 725 1356 726
rect 1316 720 1346 722
rect 1367 723 1373 724
rect 1316 719 1317 720
rect 1311 718 1317 719
rect 1367 719 1368 723
rect 1372 722 1373 723
rect 1396 722 1398 736
rect 1423 735 1424 736
rect 1428 735 1429 739
rect 1479 739 1485 740
rect 1479 738 1480 739
rect 1423 734 1429 735
rect 1452 736 1480 738
rect 1406 730 1412 731
rect 1406 726 1407 730
rect 1411 726 1412 730
rect 1406 725 1412 726
rect 1372 720 1398 722
rect 1423 723 1429 724
rect 1372 719 1373 720
rect 1367 718 1373 719
rect 1423 719 1424 723
rect 1428 722 1429 723
rect 1452 722 1454 736
rect 1479 735 1480 736
rect 1484 735 1485 739
rect 1535 739 1541 740
rect 1535 738 1536 739
rect 1479 734 1485 735
rect 1512 736 1536 738
rect 1462 730 1468 731
rect 1512 730 1514 736
rect 1535 735 1536 736
rect 1540 735 1541 739
rect 1535 734 1541 735
rect 1599 739 1605 740
rect 1599 735 1600 739
rect 1604 738 1605 739
rect 1638 739 1645 740
rect 1604 736 1634 738
rect 1604 735 1605 736
rect 1599 734 1605 735
rect 1462 726 1463 730
rect 1467 726 1468 730
rect 1462 725 1468 726
rect 1481 728 1514 730
rect 1518 730 1524 731
rect 1481 724 1483 728
rect 1518 726 1519 730
rect 1523 726 1524 730
rect 1518 725 1524 726
rect 1582 730 1588 731
rect 1582 726 1583 730
rect 1587 726 1588 730
rect 1582 725 1588 726
rect 1622 730 1628 731
rect 1622 726 1623 730
rect 1627 726 1628 730
rect 1622 725 1628 726
rect 1428 720 1454 722
rect 1479 723 1485 724
rect 1428 719 1429 720
rect 1423 718 1429 719
rect 1479 719 1480 723
rect 1484 719 1485 723
rect 1479 718 1485 719
rect 1510 723 1516 724
rect 1510 719 1511 723
rect 1515 722 1516 723
rect 1535 723 1541 724
rect 1535 722 1536 723
rect 1515 720 1536 722
rect 1515 719 1516 720
rect 1510 718 1516 719
rect 1535 719 1536 720
rect 1540 719 1541 723
rect 1535 718 1541 719
rect 1546 723 1552 724
rect 1546 719 1547 723
rect 1551 722 1552 723
rect 1599 723 1605 724
rect 1599 722 1600 723
rect 1551 720 1600 722
rect 1551 719 1552 720
rect 1546 718 1552 719
rect 1599 719 1600 720
rect 1604 719 1605 723
rect 1632 722 1634 736
rect 1638 735 1639 739
rect 1644 735 1645 739
rect 1638 734 1645 735
rect 1662 728 1668 729
rect 1662 724 1663 728
rect 1667 724 1668 728
rect 1639 723 1645 724
rect 1662 723 1668 724
rect 1639 722 1640 723
rect 1632 720 1640 722
rect 1599 718 1605 719
rect 1639 719 1640 720
rect 1644 719 1645 723
rect 1639 718 1645 719
rect 414 715 420 716
rect 414 714 415 715
rect 360 712 415 714
rect 330 710 336 711
rect 414 711 415 712
rect 419 711 420 715
rect 414 710 420 711
rect 1102 711 1108 712
rect 1102 710 1103 711
rect 977 708 1103 710
rect 390 707 396 708
rect 390 706 391 707
rect 305 704 391 706
rect 295 699 301 700
rect 110 696 116 697
rect 110 692 111 696
rect 115 692 116 696
rect 295 695 296 699
rect 300 698 301 699
rect 305 698 307 704
rect 390 703 391 704
rect 395 703 396 707
rect 390 702 396 703
rect 463 703 469 704
rect 433 700 450 702
rect 327 699 333 700
rect 327 698 328 699
rect 300 696 307 698
rect 319 696 328 698
rect 300 695 301 696
rect 110 691 116 692
rect 278 694 284 695
rect 295 694 301 695
rect 310 694 316 695
rect 278 690 279 694
rect 283 690 284 694
rect 278 689 284 690
rect 310 690 311 694
rect 315 690 316 694
rect 310 689 316 690
rect 319 684 321 696
rect 327 695 328 696
rect 332 695 333 699
rect 359 699 365 700
rect 359 698 360 699
rect 352 696 360 698
rect 327 694 333 695
rect 342 694 348 695
rect 342 690 343 694
rect 347 690 348 694
rect 342 689 348 690
rect 352 684 354 696
rect 359 695 360 696
rect 364 695 365 699
rect 391 699 397 700
rect 391 695 392 699
rect 396 698 397 699
rect 423 699 429 700
rect 396 696 402 698
rect 396 695 397 696
rect 359 694 365 695
rect 374 694 380 695
rect 391 694 397 695
rect 374 690 375 694
rect 379 690 380 694
rect 374 689 380 690
rect 400 686 402 696
rect 423 695 424 699
rect 428 698 429 699
rect 433 698 435 700
rect 428 696 435 698
rect 428 695 429 696
rect 406 694 412 695
rect 423 694 429 695
rect 438 694 444 695
rect 406 690 407 694
rect 411 690 412 694
rect 406 689 412 690
rect 438 690 439 694
rect 443 690 444 694
rect 438 689 444 690
rect 448 686 450 700
rect 455 699 461 700
rect 455 695 456 699
rect 460 695 461 699
rect 463 699 464 703
rect 468 702 469 703
rect 527 703 533 704
rect 468 700 491 702
rect 496 700 523 702
rect 468 699 469 700
rect 463 698 469 699
rect 487 699 493 700
rect 487 695 488 699
rect 492 695 493 699
rect 455 694 461 695
rect 470 694 476 695
rect 487 694 493 695
rect 457 690 459 694
rect 470 690 471 694
rect 475 690 476 694
rect 457 688 467 690
rect 470 689 476 690
rect 400 684 406 686
rect 448 684 459 686
rect 295 683 301 684
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 295 679 296 683
rect 300 682 301 683
rect 308 682 321 684
rect 327 683 333 684
rect 300 680 310 682
rect 300 679 301 680
rect 295 678 301 679
rect 327 679 328 683
rect 332 682 333 683
rect 340 682 354 684
rect 359 683 365 684
rect 332 680 342 682
rect 332 679 333 680
rect 327 678 333 679
rect 359 679 360 683
rect 364 679 365 683
rect 359 678 365 679
rect 390 683 397 684
rect 390 679 391 683
rect 396 679 397 683
rect 404 682 418 684
rect 423 683 429 684
rect 423 682 424 683
rect 416 680 424 682
rect 390 678 397 679
rect 423 679 424 680
rect 428 679 429 683
rect 423 678 429 679
rect 455 683 461 684
rect 455 679 456 683
rect 460 679 461 683
rect 455 678 461 679
rect 110 674 116 675
rect 278 677 284 678
rect 278 673 279 677
rect 283 673 284 677
rect 278 672 284 673
rect 310 677 316 678
rect 310 673 311 677
rect 315 673 316 677
rect 310 672 316 673
rect 342 677 348 678
rect 342 673 343 677
rect 347 673 348 677
rect 342 672 348 673
rect 374 677 380 678
rect 374 673 375 677
rect 379 673 380 677
rect 374 672 380 673
rect 406 677 412 678
rect 406 673 407 677
rect 411 673 412 677
rect 406 672 412 673
rect 438 677 444 678
rect 438 673 439 677
rect 443 673 444 677
rect 438 672 444 673
rect 465 670 467 688
rect 487 683 493 684
rect 487 679 488 683
rect 492 682 493 683
rect 496 682 498 700
rect 519 699 525 700
rect 519 695 520 699
rect 524 695 525 699
rect 527 699 528 703
rect 532 702 533 703
rect 567 703 573 704
rect 532 700 554 702
rect 532 699 533 700
rect 527 698 533 699
rect 552 698 554 700
rect 559 699 565 700
rect 559 698 560 699
rect 552 696 560 698
rect 559 695 560 696
rect 564 695 565 699
rect 567 699 568 703
rect 572 702 573 703
rect 615 703 621 704
rect 572 700 602 702
rect 572 699 573 700
rect 567 698 573 699
rect 600 698 602 700
rect 607 699 613 700
rect 607 698 608 699
rect 600 696 608 698
rect 607 695 608 696
rect 612 695 613 699
rect 615 699 616 703
rect 620 702 621 703
rect 671 703 677 704
rect 620 700 658 702
rect 620 699 621 700
rect 615 698 621 699
rect 656 698 658 700
rect 663 699 669 700
rect 663 698 664 699
rect 656 696 664 698
rect 663 695 664 696
rect 668 695 669 699
rect 671 699 672 703
rect 676 702 677 703
rect 783 703 789 704
rect 676 700 714 702
rect 676 699 677 700
rect 671 698 677 699
rect 712 698 714 700
rect 719 699 725 700
rect 719 698 720 699
rect 712 696 720 698
rect 719 695 720 696
rect 724 695 725 699
rect 774 699 781 700
rect 774 695 775 699
rect 780 695 781 699
rect 783 699 784 703
rect 788 702 789 703
rect 847 703 853 704
rect 788 700 834 702
rect 788 699 789 700
rect 783 698 789 699
rect 832 698 834 700
rect 839 699 845 700
rect 839 698 840 699
rect 832 696 840 698
rect 839 695 840 696
rect 844 695 845 699
rect 847 699 848 703
rect 852 702 853 703
rect 852 700 907 702
rect 977 700 979 708
rect 1102 707 1103 708
rect 1107 707 1108 711
rect 1638 711 1644 712
rect 1638 710 1639 711
rect 1102 706 1108 707
rect 1601 708 1639 710
rect 1047 703 1053 704
rect 852 699 853 700
rect 847 698 853 699
rect 903 699 909 700
rect 903 695 904 699
rect 908 695 909 699
rect 975 699 981 700
rect 975 695 976 699
rect 980 695 981 699
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 698 1036 699
rect 1039 699 1045 700
rect 1039 698 1040 699
rect 1035 696 1040 698
rect 1035 695 1036 696
rect 502 694 508 695
rect 519 694 525 695
rect 542 694 548 695
rect 559 694 565 695
rect 590 694 596 695
rect 607 694 613 695
rect 646 694 652 695
rect 663 694 669 695
rect 702 694 708 695
rect 719 694 725 695
rect 758 694 764 695
rect 774 694 781 695
rect 822 694 828 695
rect 839 694 845 695
rect 886 694 892 695
rect 903 694 909 695
rect 958 694 964 695
rect 975 694 981 695
rect 1022 694 1028 695
rect 1030 694 1036 695
rect 1039 695 1040 696
rect 1044 695 1045 699
rect 1047 699 1048 703
rect 1052 702 1053 703
rect 1183 703 1189 704
rect 1052 700 1098 702
rect 1052 699 1053 700
rect 1047 698 1053 699
rect 1096 698 1098 700
rect 1103 699 1109 700
rect 1103 698 1104 699
rect 1096 696 1104 698
rect 1103 695 1104 696
rect 1108 695 1109 699
rect 1175 699 1181 700
rect 1175 695 1176 699
rect 1180 695 1181 699
rect 1183 699 1184 703
rect 1188 702 1189 703
rect 1247 703 1253 704
rect 1188 700 1234 702
rect 1188 699 1189 700
rect 1183 698 1189 699
rect 1232 698 1234 700
rect 1239 699 1245 700
rect 1239 698 1240 699
rect 1232 696 1240 698
rect 1039 694 1045 695
rect 1086 694 1092 695
rect 1103 694 1109 695
rect 1158 694 1164 695
rect 1175 694 1181 695
rect 1207 695 1213 696
rect 1239 695 1240 696
rect 1244 695 1245 699
rect 1247 699 1248 703
rect 1252 702 1253 703
rect 1311 703 1317 704
rect 1252 700 1298 702
rect 1252 699 1253 700
rect 1247 698 1253 699
rect 1296 698 1298 700
rect 1303 699 1309 700
rect 1303 698 1304 699
rect 1296 696 1304 698
rect 1303 695 1304 696
rect 1308 695 1309 699
rect 1311 699 1312 703
rect 1316 702 1317 703
rect 1375 703 1381 704
rect 1316 700 1371 702
rect 1316 699 1317 700
rect 1311 698 1317 699
rect 1367 699 1373 700
rect 1367 695 1368 699
rect 1372 695 1373 699
rect 1375 699 1376 703
rect 1380 702 1381 703
rect 1495 703 1501 704
rect 1380 700 1426 702
rect 1380 699 1381 700
rect 1375 698 1381 699
rect 1424 698 1426 700
rect 1431 699 1437 700
rect 1431 698 1432 699
rect 1424 696 1432 698
rect 1431 695 1432 696
rect 1436 695 1437 699
rect 1486 699 1493 700
rect 1486 695 1487 699
rect 1492 695 1493 699
rect 1495 699 1496 703
rect 1500 702 1501 703
rect 1500 700 1547 702
rect 1601 700 1603 708
rect 1638 707 1639 708
rect 1643 707 1644 711
rect 1638 706 1644 707
rect 1607 703 1613 704
rect 1500 699 1501 700
rect 1495 698 1501 699
rect 1543 699 1549 700
rect 1543 695 1544 699
rect 1548 695 1549 699
rect 1599 699 1605 700
rect 1599 695 1600 699
rect 1604 695 1605 699
rect 1607 699 1608 703
rect 1612 702 1613 703
rect 1612 700 1643 702
rect 1612 699 1613 700
rect 1607 698 1613 699
rect 1639 699 1645 700
rect 1639 695 1640 699
rect 1644 695 1645 699
rect 1207 694 1208 695
rect 502 690 503 694
rect 507 690 508 694
rect 502 689 508 690
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 590 690 591 694
rect 595 690 596 694
rect 590 689 596 690
rect 646 690 647 694
rect 651 690 652 694
rect 646 689 652 690
rect 702 690 703 694
rect 707 690 708 694
rect 702 689 708 690
rect 758 690 759 694
rect 763 690 764 694
rect 758 689 764 690
rect 822 690 823 694
rect 827 690 828 694
rect 822 689 828 690
rect 886 690 887 694
rect 891 690 892 694
rect 886 689 892 690
rect 958 690 959 694
rect 963 690 964 694
rect 958 689 964 690
rect 1022 690 1023 694
rect 1027 690 1028 694
rect 1022 689 1028 690
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1086 689 1092 690
rect 1158 690 1159 694
rect 1163 690 1164 694
rect 1177 692 1208 694
rect 1207 691 1208 692
rect 1212 691 1213 695
rect 1207 690 1213 691
rect 1222 694 1228 695
rect 1239 694 1245 695
rect 1286 694 1292 695
rect 1303 694 1309 695
rect 1350 694 1356 695
rect 1367 694 1373 695
rect 1414 694 1420 695
rect 1431 694 1437 695
rect 1470 694 1476 695
rect 1486 694 1493 695
rect 1526 694 1532 695
rect 1543 694 1549 695
rect 1582 694 1588 695
rect 1599 694 1605 695
rect 1622 694 1628 695
rect 1639 694 1645 695
rect 1662 696 1668 697
rect 1222 690 1223 694
rect 1227 690 1228 694
rect 1158 689 1164 690
rect 1222 689 1228 690
rect 1286 690 1287 694
rect 1291 690 1292 694
rect 1286 689 1292 690
rect 1350 690 1351 694
rect 1355 690 1356 694
rect 1350 689 1356 690
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1414 689 1420 690
rect 1470 690 1471 694
rect 1475 690 1476 694
rect 1470 689 1476 690
rect 1526 690 1527 694
rect 1531 690 1532 694
rect 1526 689 1532 690
rect 1582 690 1583 694
rect 1587 690 1588 694
rect 1582 689 1588 690
rect 1622 690 1623 694
rect 1627 690 1628 694
rect 1662 692 1663 696
rect 1667 692 1668 696
rect 1662 691 1668 692
rect 1622 689 1628 690
rect 492 680 498 682
rect 519 683 525 684
rect 492 679 493 680
rect 487 678 493 679
rect 519 679 520 683
rect 524 682 525 683
rect 527 683 533 684
rect 527 682 528 683
rect 524 680 528 682
rect 524 679 525 680
rect 519 678 525 679
rect 527 679 528 680
rect 532 679 533 683
rect 527 678 533 679
rect 559 683 565 684
rect 559 679 560 683
rect 564 682 565 683
rect 567 683 573 684
rect 567 682 568 683
rect 564 680 568 682
rect 564 679 565 680
rect 559 678 565 679
rect 567 679 568 680
rect 572 679 573 683
rect 567 678 573 679
rect 607 683 613 684
rect 607 679 608 683
rect 612 682 613 683
rect 615 683 621 684
rect 615 682 616 683
rect 612 680 616 682
rect 612 679 613 680
rect 607 678 613 679
rect 615 679 616 680
rect 620 679 621 683
rect 615 678 621 679
rect 663 683 669 684
rect 663 679 664 683
rect 668 682 669 683
rect 671 683 677 684
rect 671 682 672 683
rect 668 680 672 682
rect 668 679 669 680
rect 663 678 669 679
rect 671 679 672 680
rect 676 679 677 683
rect 719 683 725 684
rect 719 682 720 683
rect 671 678 677 679
rect 712 680 720 682
rect 470 677 476 678
rect 470 673 471 677
rect 475 673 476 677
rect 470 672 476 673
rect 502 677 508 678
rect 502 673 503 677
rect 507 673 508 677
rect 502 672 508 673
rect 542 677 548 678
rect 542 673 543 677
rect 547 673 548 677
rect 542 672 548 673
rect 590 677 596 678
rect 590 673 591 677
rect 595 673 596 677
rect 590 672 596 673
rect 646 677 652 678
rect 646 673 647 677
rect 651 673 652 677
rect 646 672 652 673
rect 702 677 708 678
rect 702 673 703 677
rect 707 673 708 677
rect 702 672 708 673
rect 534 671 540 672
rect 465 668 507 670
rect 294 663 300 664
rect 110 661 116 662
rect 110 657 111 661
rect 115 657 116 661
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 326 663 332 664
rect 326 659 327 663
rect 331 659 332 663
rect 326 658 332 659
rect 358 663 364 664
rect 358 659 359 663
rect 363 659 364 663
rect 358 658 364 659
rect 390 663 396 664
rect 390 659 391 663
rect 395 659 396 663
rect 390 658 396 659
rect 422 663 428 664
rect 422 659 423 663
rect 427 659 428 663
rect 422 658 428 659
rect 454 663 460 664
rect 454 659 455 663
rect 459 659 460 663
rect 454 658 460 659
rect 486 663 492 664
rect 486 659 487 663
rect 491 659 492 663
rect 486 658 492 659
rect 110 656 116 657
rect 505 656 507 668
rect 534 667 535 671
rect 539 670 540 671
rect 712 670 714 680
rect 719 679 720 680
rect 724 679 725 683
rect 719 678 725 679
rect 775 683 781 684
rect 775 679 776 683
rect 780 682 781 683
rect 783 683 789 684
rect 783 682 784 683
rect 780 680 784 682
rect 780 679 781 680
rect 775 678 781 679
rect 783 679 784 680
rect 788 679 789 683
rect 783 678 789 679
rect 839 683 845 684
rect 839 679 840 683
rect 844 682 845 683
rect 847 683 853 684
rect 847 682 848 683
rect 844 680 848 682
rect 844 679 845 680
rect 839 678 845 679
rect 847 679 848 680
rect 852 679 853 683
rect 847 678 853 679
rect 903 683 909 684
rect 903 679 904 683
rect 908 682 909 683
rect 926 683 932 684
rect 926 682 927 683
rect 908 680 927 682
rect 908 679 909 680
rect 903 678 909 679
rect 926 679 927 680
rect 931 679 932 683
rect 926 678 932 679
rect 974 683 981 684
rect 974 679 975 683
rect 980 679 981 683
rect 974 678 981 679
rect 1039 683 1045 684
rect 1039 679 1040 683
rect 1044 682 1045 683
rect 1047 683 1053 684
rect 1047 682 1048 683
rect 1044 680 1048 682
rect 1044 679 1045 680
rect 1039 678 1045 679
rect 1047 679 1048 680
rect 1052 679 1053 683
rect 1047 678 1053 679
rect 1102 683 1109 684
rect 1102 679 1103 683
rect 1108 679 1109 683
rect 1102 678 1109 679
rect 1175 683 1181 684
rect 1175 679 1176 683
rect 1180 682 1181 683
rect 1183 683 1189 684
rect 1183 682 1184 683
rect 1180 680 1184 682
rect 1180 679 1181 680
rect 1175 678 1181 679
rect 1183 679 1184 680
rect 1188 679 1189 683
rect 1183 678 1189 679
rect 1239 683 1245 684
rect 1239 679 1240 683
rect 1244 682 1245 683
rect 1247 683 1253 684
rect 1247 682 1248 683
rect 1244 680 1248 682
rect 1244 679 1245 680
rect 1239 678 1245 679
rect 1247 679 1248 680
rect 1252 679 1253 683
rect 1247 678 1253 679
rect 1303 683 1309 684
rect 1303 679 1304 683
rect 1308 682 1309 683
rect 1311 683 1317 684
rect 1311 682 1312 683
rect 1308 680 1312 682
rect 1308 679 1309 680
rect 1303 678 1309 679
rect 1311 679 1312 680
rect 1316 679 1317 683
rect 1311 678 1317 679
rect 1367 683 1373 684
rect 1367 679 1368 683
rect 1372 682 1373 683
rect 1375 683 1381 684
rect 1375 682 1376 683
rect 1372 680 1376 682
rect 1372 679 1373 680
rect 1367 678 1373 679
rect 1375 679 1376 680
rect 1380 679 1381 683
rect 1375 678 1381 679
rect 1426 683 1437 684
rect 1426 679 1427 683
rect 1431 679 1432 683
rect 1436 679 1437 683
rect 1426 678 1437 679
rect 1487 683 1493 684
rect 1487 679 1488 683
rect 1492 682 1493 683
rect 1495 683 1501 684
rect 1495 682 1496 683
rect 1492 680 1496 682
rect 1492 679 1493 680
rect 1487 678 1493 679
rect 1495 679 1496 680
rect 1500 679 1501 683
rect 1495 678 1501 679
rect 1543 683 1552 684
rect 1543 679 1544 683
rect 1551 679 1552 683
rect 1543 678 1552 679
rect 1599 683 1605 684
rect 1599 679 1600 683
rect 1604 682 1605 683
rect 1607 683 1613 684
rect 1607 682 1608 683
rect 1604 680 1608 682
rect 1604 679 1605 680
rect 1599 678 1605 679
rect 1607 679 1608 680
rect 1612 679 1613 683
rect 1607 678 1613 679
rect 1638 683 1645 684
rect 1638 679 1639 683
rect 1644 679 1645 683
rect 1638 678 1645 679
rect 1662 679 1668 680
rect 758 677 764 678
rect 758 673 759 677
rect 763 673 764 677
rect 758 672 764 673
rect 822 677 828 678
rect 822 673 823 677
rect 827 673 828 677
rect 822 672 828 673
rect 886 677 892 678
rect 886 673 887 677
rect 891 673 892 677
rect 886 672 892 673
rect 958 677 964 678
rect 958 673 959 677
rect 963 673 964 677
rect 958 672 964 673
rect 1022 677 1028 678
rect 1022 673 1023 677
rect 1027 673 1028 677
rect 1022 672 1028 673
rect 1086 677 1092 678
rect 1086 673 1087 677
rect 1091 673 1092 677
rect 1086 672 1092 673
rect 1158 677 1164 678
rect 1158 673 1159 677
rect 1163 673 1164 677
rect 1158 672 1164 673
rect 1222 677 1228 678
rect 1222 673 1223 677
rect 1227 673 1228 677
rect 1222 672 1228 673
rect 1286 677 1292 678
rect 1286 673 1287 677
rect 1291 673 1292 677
rect 1286 672 1292 673
rect 1350 677 1356 678
rect 1350 673 1351 677
rect 1355 673 1356 677
rect 1350 672 1356 673
rect 1414 677 1420 678
rect 1414 673 1415 677
rect 1419 673 1420 677
rect 1414 672 1420 673
rect 1470 677 1476 678
rect 1470 673 1471 677
rect 1475 673 1476 677
rect 1470 672 1476 673
rect 1526 677 1532 678
rect 1526 673 1527 677
rect 1531 673 1532 677
rect 1526 672 1532 673
rect 1582 677 1588 678
rect 1582 673 1583 677
rect 1587 673 1588 677
rect 1582 672 1588 673
rect 1622 677 1628 678
rect 1622 673 1623 677
rect 1627 673 1628 677
rect 1662 675 1663 679
rect 1667 675 1668 679
rect 1662 674 1668 675
rect 1622 672 1628 673
rect 539 668 714 670
rect 539 667 540 668
rect 534 666 540 667
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 550 663 556 664
rect 550 659 551 663
rect 555 659 556 663
rect 550 658 556 659
rect 590 663 596 664
rect 590 659 591 663
rect 595 659 596 663
rect 590 658 596 659
rect 638 663 644 664
rect 638 659 639 663
rect 643 659 644 663
rect 638 658 644 659
rect 686 663 692 664
rect 686 659 687 663
rect 691 659 692 663
rect 686 658 692 659
rect 734 663 740 664
rect 734 659 735 663
rect 739 659 740 663
rect 734 658 740 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 659 796 663
rect 790 658 796 659
rect 846 663 852 664
rect 846 659 847 663
rect 851 659 852 663
rect 846 658 852 659
rect 910 663 916 664
rect 910 659 911 663
rect 915 659 916 663
rect 910 658 916 659
rect 974 663 980 664
rect 974 659 975 663
rect 979 659 980 663
rect 974 658 980 659
rect 1046 663 1052 664
rect 1046 659 1047 663
rect 1051 659 1052 663
rect 1046 658 1052 659
rect 1126 663 1132 664
rect 1126 659 1127 663
rect 1131 659 1132 663
rect 1126 658 1132 659
rect 1214 663 1220 664
rect 1214 659 1215 663
rect 1219 659 1220 663
rect 1214 658 1220 659
rect 1294 663 1300 664
rect 1294 659 1295 663
rect 1299 659 1300 663
rect 1294 658 1300 659
rect 1382 663 1388 664
rect 1382 659 1383 663
rect 1387 659 1388 663
rect 1382 658 1388 659
rect 1470 663 1476 664
rect 1470 659 1471 663
rect 1475 659 1476 663
rect 1470 658 1476 659
rect 1558 663 1564 664
rect 1558 659 1559 663
rect 1563 659 1564 663
rect 1558 658 1564 659
rect 1622 663 1628 664
rect 1622 659 1623 663
rect 1627 659 1628 663
rect 1622 658 1628 659
rect 1662 661 1668 662
rect 1662 657 1663 661
rect 1667 657 1668 661
rect 1662 656 1668 657
rect 311 655 317 656
rect 311 651 312 655
rect 316 654 317 655
rect 343 655 349 656
rect 316 652 338 654
rect 316 651 317 652
rect 311 650 317 651
rect 294 646 300 647
rect 110 644 116 645
rect 110 640 111 644
rect 115 640 116 644
rect 294 642 295 646
rect 299 642 300 646
rect 294 641 300 642
rect 326 646 332 647
rect 326 642 327 646
rect 331 642 332 646
rect 326 641 332 642
rect 110 639 116 640
rect 311 639 317 640
rect 311 635 312 639
rect 316 638 317 639
rect 336 638 338 652
rect 343 651 344 655
rect 348 654 349 655
rect 375 655 381 656
rect 348 652 370 654
rect 348 651 349 652
rect 343 650 349 651
rect 358 646 364 647
rect 358 642 359 646
rect 363 642 364 646
rect 358 641 364 642
rect 343 639 349 640
rect 343 638 344 639
rect 316 636 321 638
rect 336 636 344 638
rect 316 635 317 636
rect 311 634 317 635
rect 319 630 321 636
rect 343 635 344 636
rect 348 635 349 639
rect 368 638 370 652
rect 375 651 376 655
rect 380 654 381 655
rect 407 655 413 656
rect 380 652 402 654
rect 380 651 381 652
rect 375 650 381 651
rect 390 646 396 647
rect 390 642 391 646
rect 395 642 396 646
rect 390 641 396 642
rect 375 639 381 640
rect 375 638 376 639
rect 368 636 376 638
rect 343 634 349 635
rect 375 635 376 636
rect 380 635 381 639
rect 400 638 402 652
rect 407 651 408 655
rect 412 654 413 655
rect 439 655 445 656
rect 412 652 434 654
rect 412 651 413 652
rect 407 650 413 651
rect 422 646 428 647
rect 422 642 423 646
rect 427 642 428 646
rect 422 641 428 642
rect 407 639 413 640
rect 407 638 408 639
rect 400 636 408 638
rect 375 634 381 635
rect 407 635 408 636
rect 412 635 413 639
rect 432 638 434 652
rect 439 651 440 655
rect 444 654 445 655
rect 471 655 477 656
rect 444 652 466 654
rect 444 651 445 652
rect 439 650 445 651
rect 454 646 460 647
rect 454 642 455 646
rect 459 642 460 646
rect 454 641 460 642
rect 439 639 445 640
rect 439 638 440 639
rect 432 636 440 638
rect 407 634 413 635
rect 439 635 440 636
rect 444 635 445 639
rect 464 638 466 652
rect 471 651 472 655
rect 476 654 477 655
rect 503 655 509 656
rect 476 652 498 654
rect 476 651 477 652
rect 471 650 477 651
rect 486 646 492 647
rect 486 642 487 646
rect 491 642 492 646
rect 486 641 492 642
rect 471 639 477 640
rect 471 638 472 639
rect 464 636 472 638
rect 439 634 445 635
rect 471 635 472 636
rect 476 635 477 639
rect 496 638 498 652
rect 503 651 504 655
rect 508 651 509 655
rect 503 650 509 651
rect 535 655 541 656
rect 535 651 536 655
rect 540 654 541 655
rect 567 655 573 656
rect 540 652 562 654
rect 540 651 541 652
rect 535 650 541 651
rect 518 646 524 647
rect 518 642 519 646
rect 523 642 524 646
rect 518 641 524 642
rect 550 646 556 647
rect 550 642 551 646
rect 555 642 556 646
rect 550 641 556 642
rect 503 639 509 640
rect 503 638 504 639
rect 496 636 504 638
rect 471 634 477 635
rect 503 635 504 636
rect 508 635 509 639
rect 503 634 509 635
rect 534 639 541 640
rect 534 635 535 639
rect 540 635 541 639
rect 560 638 562 652
rect 567 651 568 655
rect 572 654 573 655
rect 607 655 613 656
rect 572 652 587 654
rect 572 651 573 652
rect 567 650 573 651
rect 567 639 573 640
rect 567 638 568 639
rect 560 636 568 638
rect 534 634 541 635
rect 567 635 568 636
rect 572 635 573 639
rect 585 638 587 652
rect 607 651 608 655
rect 612 654 613 655
rect 655 655 661 656
rect 612 652 634 654
rect 612 651 613 652
rect 607 650 613 651
rect 590 646 596 647
rect 590 642 591 646
rect 595 642 596 646
rect 590 641 596 642
rect 607 639 613 640
rect 607 638 608 639
rect 585 636 608 638
rect 567 634 573 635
rect 607 635 608 636
rect 612 635 613 639
rect 632 638 634 652
rect 655 651 656 655
rect 660 654 661 655
rect 703 655 709 656
rect 660 652 683 654
rect 660 651 661 652
rect 655 650 661 651
rect 638 646 644 647
rect 638 642 639 646
rect 643 642 644 646
rect 638 641 644 642
rect 655 639 661 640
rect 655 638 656 639
rect 632 636 656 638
rect 607 634 613 635
rect 655 635 656 636
rect 660 635 661 639
rect 681 638 683 652
rect 703 651 704 655
rect 708 654 709 655
rect 750 655 757 656
rect 708 652 746 654
rect 708 651 709 652
rect 703 650 709 651
rect 686 646 692 647
rect 686 642 687 646
rect 691 642 692 646
rect 686 641 692 642
rect 734 646 740 647
rect 734 642 735 646
rect 739 642 740 646
rect 734 641 740 642
rect 703 639 709 640
rect 703 638 704 639
rect 681 636 704 638
rect 655 634 661 635
rect 703 635 704 636
rect 708 635 709 639
rect 744 638 746 652
rect 750 651 751 655
rect 756 651 757 655
rect 750 650 757 651
rect 807 655 813 656
rect 807 651 808 655
rect 812 654 813 655
rect 838 655 844 656
rect 838 654 839 655
rect 812 652 839 654
rect 812 651 813 652
rect 807 650 813 651
rect 838 651 839 652
rect 843 651 844 655
rect 863 655 869 656
rect 863 654 864 655
rect 838 650 844 651
rect 856 652 864 654
rect 790 646 796 647
rect 790 642 791 646
rect 795 642 796 646
rect 790 641 796 642
rect 846 646 852 647
rect 846 642 847 646
rect 851 642 852 646
rect 846 641 852 642
rect 751 639 757 640
rect 751 638 752 639
rect 744 636 752 638
rect 703 634 709 635
rect 751 635 752 636
rect 756 635 757 639
rect 751 634 757 635
rect 807 639 813 640
rect 807 635 808 639
rect 812 638 813 639
rect 856 638 858 652
rect 863 651 864 652
rect 868 651 869 655
rect 927 655 933 656
rect 927 654 928 655
rect 863 650 869 651
rect 897 652 928 654
rect 812 636 858 638
rect 863 639 869 640
rect 812 635 813 636
rect 807 634 813 635
rect 863 635 864 639
rect 868 638 869 639
rect 897 638 899 652
rect 927 651 928 652
rect 932 651 933 655
rect 927 650 933 651
rect 991 655 997 656
rect 991 651 992 655
rect 996 654 997 655
rect 1030 655 1036 656
rect 1030 654 1031 655
rect 996 652 1031 654
rect 996 651 997 652
rect 991 650 997 651
rect 1030 651 1031 652
rect 1035 651 1036 655
rect 1063 655 1069 656
rect 1063 654 1064 655
rect 1030 650 1036 651
rect 1040 652 1064 654
rect 910 646 916 647
rect 910 642 911 646
rect 915 642 916 646
rect 910 641 916 642
rect 974 646 980 647
rect 974 642 975 646
rect 979 642 980 646
rect 974 641 980 642
rect 868 636 899 638
rect 926 639 933 640
rect 868 635 869 636
rect 863 634 869 635
rect 926 635 927 639
rect 932 635 933 639
rect 926 634 933 635
rect 991 639 997 640
rect 991 635 992 639
rect 996 638 997 639
rect 1040 638 1042 652
rect 1063 651 1064 652
rect 1068 651 1069 655
rect 1143 655 1149 656
rect 1143 654 1144 655
rect 1063 650 1069 651
rect 1108 652 1144 654
rect 1046 646 1052 647
rect 1046 642 1047 646
rect 1051 642 1052 646
rect 1046 641 1052 642
rect 996 636 1042 638
rect 1063 639 1069 640
rect 996 635 997 636
rect 991 634 997 635
rect 1063 635 1064 639
rect 1068 638 1069 639
rect 1108 638 1110 652
rect 1143 651 1144 652
rect 1148 651 1149 655
rect 1143 650 1149 651
rect 1226 655 1237 656
rect 1226 651 1227 655
rect 1231 651 1232 655
rect 1236 651 1237 655
rect 1311 655 1317 656
rect 1311 654 1312 655
rect 1226 650 1237 651
rect 1276 652 1312 654
rect 1126 646 1132 647
rect 1126 642 1127 646
rect 1131 642 1132 646
rect 1126 641 1132 642
rect 1214 646 1220 647
rect 1214 642 1215 646
rect 1219 642 1220 646
rect 1214 641 1220 642
rect 1068 636 1110 638
rect 1142 639 1149 640
rect 1068 635 1069 636
rect 1063 634 1069 635
rect 1142 635 1143 639
rect 1148 635 1149 639
rect 1142 634 1149 635
rect 1231 639 1237 640
rect 1231 635 1232 639
rect 1236 638 1237 639
rect 1276 638 1278 652
rect 1311 651 1312 652
rect 1316 651 1317 655
rect 1399 655 1405 656
rect 1399 654 1400 655
rect 1311 650 1317 651
rect 1356 652 1400 654
rect 1294 646 1300 647
rect 1294 642 1295 646
rect 1299 642 1300 646
rect 1294 641 1300 642
rect 1236 636 1278 638
rect 1311 639 1317 640
rect 1236 635 1237 636
rect 1231 634 1237 635
rect 1311 635 1312 639
rect 1316 638 1317 639
rect 1356 638 1358 652
rect 1399 651 1400 652
rect 1404 651 1405 655
rect 1399 650 1405 651
rect 1486 655 1493 656
rect 1486 651 1487 655
rect 1492 651 1493 655
rect 1575 655 1581 656
rect 1575 654 1576 655
rect 1486 650 1493 651
rect 1532 652 1576 654
rect 1382 646 1388 647
rect 1382 642 1383 646
rect 1387 642 1388 646
rect 1382 641 1388 642
rect 1470 646 1476 647
rect 1470 642 1471 646
rect 1475 642 1476 646
rect 1470 641 1476 642
rect 1316 636 1358 638
rect 1399 639 1405 640
rect 1316 635 1317 636
rect 1311 634 1317 635
rect 1399 635 1400 639
rect 1404 638 1405 639
rect 1426 639 1432 640
rect 1426 638 1427 639
rect 1404 636 1427 638
rect 1404 635 1405 636
rect 1399 634 1405 635
rect 1426 635 1427 636
rect 1431 635 1432 639
rect 1426 634 1432 635
rect 1487 639 1493 640
rect 1487 635 1488 639
rect 1492 638 1493 639
rect 1532 638 1534 652
rect 1575 651 1576 652
rect 1580 651 1581 655
rect 1575 650 1581 651
rect 1639 655 1645 656
rect 1639 651 1640 655
rect 1644 654 1645 655
rect 1647 655 1653 656
rect 1647 654 1648 655
rect 1644 652 1648 654
rect 1644 651 1645 652
rect 1639 650 1645 651
rect 1647 651 1648 652
rect 1652 651 1653 655
rect 1647 650 1653 651
rect 1558 646 1564 647
rect 1558 642 1559 646
rect 1563 642 1564 646
rect 1558 641 1564 642
rect 1622 646 1628 647
rect 1622 642 1623 646
rect 1627 642 1628 646
rect 1622 641 1628 642
rect 1662 644 1668 645
rect 1662 640 1663 644
rect 1667 640 1668 644
rect 1492 636 1534 638
rect 1575 639 1581 640
rect 1492 635 1493 636
rect 1487 634 1493 635
rect 1575 635 1576 639
rect 1580 638 1581 639
rect 1590 639 1596 640
rect 1590 638 1591 639
rect 1580 636 1591 638
rect 1580 635 1581 636
rect 1575 634 1581 635
rect 1590 635 1591 636
rect 1595 635 1596 639
rect 1590 634 1596 635
rect 1638 639 1645 640
rect 1662 639 1668 640
rect 1638 635 1639 639
rect 1644 635 1645 639
rect 1638 634 1645 635
rect 478 631 484 632
rect 478 630 479 631
rect 319 628 479 630
rect 478 627 479 628
rect 483 627 484 631
rect 750 631 756 632
rect 750 630 751 631
rect 478 626 484 627
rect 537 628 751 630
rect 303 623 309 624
rect 262 619 269 620
rect 110 616 116 617
rect 110 612 111 616
rect 115 612 116 616
rect 262 615 263 619
rect 268 615 269 619
rect 295 619 301 620
rect 295 618 296 619
rect 288 616 296 618
rect 110 611 116 612
rect 246 614 252 615
rect 262 614 269 615
rect 278 614 284 615
rect 246 610 247 614
rect 251 610 252 614
rect 246 609 252 610
rect 278 610 279 614
rect 283 610 284 614
rect 278 609 284 610
rect 288 604 290 616
rect 295 615 296 616
rect 300 615 301 619
rect 303 619 304 623
rect 308 622 309 623
rect 351 623 357 624
rect 308 620 330 622
rect 308 619 309 620
rect 303 618 309 619
rect 328 618 330 620
rect 335 619 341 620
rect 335 618 336 619
rect 328 616 336 618
rect 335 615 336 616
rect 340 615 341 619
rect 351 619 352 623
rect 356 622 357 623
rect 391 623 397 624
rect 356 620 387 622
rect 356 619 357 620
rect 351 618 357 619
rect 383 619 389 620
rect 383 615 384 619
rect 388 615 389 619
rect 391 619 392 623
rect 396 622 397 623
rect 447 623 453 624
rect 396 620 434 622
rect 396 619 397 620
rect 391 618 397 619
rect 432 618 434 620
rect 439 619 445 620
rect 439 618 440 619
rect 432 616 440 618
rect 439 615 440 616
rect 444 615 445 619
rect 447 619 448 623
rect 452 622 453 623
rect 452 620 491 622
rect 537 620 539 628
rect 750 627 751 628
rect 755 627 756 631
rect 750 626 756 627
rect 543 623 549 624
rect 452 619 453 620
rect 447 618 453 619
rect 487 619 493 620
rect 487 615 488 619
rect 492 615 493 619
rect 535 619 541 620
rect 535 615 536 619
rect 540 615 541 619
rect 543 619 544 623
rect 548 622 549 623
rect 591 623 597 624
rect 548 620 587 622
rect 548 619 549 620
rect 543 618 549 619
rect 583 619 589 620
rect 583 615 584 619
rect 588 615 589 619
rect 591 619 592 623
rect 596 622 597 623
rect 639 623 645 624
rect 596 620 626 622
rect 596 619 597 620
rect 591 618 597 619
rect 624 618 626 620
rect 631 619 637 620
rect 631 618 632 619
rect 624 616 632 618
rect 631 615 632 616
rect 636 615 637 619
rect 639 619 640 623
rect 644 622 645 623
rect 687 623 693 624
rect 644 620 683 622
rect 644 619 645 620
rect 639 618 645 619
rect 679 619 685 620
rect 679 615 680 619
rect 684 615 685 619
rect 687 619 688 623
rect 692 622 693 623
rect 743 623 749 624
rect 692 620 730 622
rect 692 619 693 620
rect 687 618 693 619
rect 728 618 730 620
rect 735 619 741 620
rect 735 618 736 619
rect 728 616 736 618
rect 735 615 736 616
rect 740 615 741 619
rect 743 619 744 623
rect 748 622 749 623
rect 855 623 861 624
rect 748 620 786 622
rect 748 619 749 620
rect 743 618 749 619
rect 784 618 786 620
rect 791 619 797 620
rect 791 618 792 619
rect 784 616 792 618
rect 791 615 792 616
rect 796 615 797 619
rect 838 619 844 620
rect 838 615 839 619
rect 843 618 844 619
rect 847 619 853 620
rect 847 618 848 619
rect 843 616 848 618
rect 843 615 844 616
rect 295 614 301 615
rect 318 614 324 615
rect 335 614 341 615
rect 366 614 372 615
rect 383 614 389 615
rect 422 614 428 615
rect 439 614 445 615
rect 470 614 476 615
rect 487 614 493 615
rect 518 614 524 615
rect 535 614 541 615
rect 566 614 572 615
rect 583 614 589 615
rect 614 614 620 615
rect 631 614 637 615
rect 662 614 668 615
rect 679 614 685 615
rect 718 614 724 615
rect 735 614 741 615
rect 774 614 780 615
rect 791 614 797 615
rect 830 614 836 615
rect 838 614 844 615
rect 847 615 848 616
rect 852 615 853 619
rect 855 619 856 623
rect 860 622 861 623
rect 919 623 925 624
rect 860 620 906 622
rect 860 619 861 620
rect 855 618 861 619
rect 904 618 906 620
rect 911 619 917 620
rect 911 618 912 619
rect 904 616 912 618
rect 911 615 912 616
rect 916 615 917 619
rect 919 619 920 623
rect 924 622 925 623
rect 1071 623 1077 624
rect 924 620 987 622
rect 924 619 925 620
rect 919 618 925 619
rect 983 619 989 620
rect 983 615 984 619
rect 988 615 989 619
rect 1063 619 1069 620
rect 1063 615 1064 619
rect 1068 615 1069 619
rect 1071 619 1072 623
rect 1076 622 1077 623
rect 1234 623 1240 624
rect 1076 620 1138 622
rect 1076 619 1077 620
rect 1071 618 1077 619
rect 1136 618 1138 620
rect 1143 619 1149 620
rect 1143 618 1144 619
rect 1136 616 1144 618
rect 847 614 853 615
rect 894 614 900 615
rect 911 614 917 615
rect 966 614 972 615
rect 983 614 989 615
rect 1046 614 1052 615
rect 1063 614 1069 615
rect 1118 615 1124 616
rect 1143 615 1144 616
rect 1148 615 1149 619
rect 1223 619 1232 620
rect 1223 615 1224 619
rect 1231 615 1232 619
rect 1234 619 1235 623
rect 1239 622 1240 623
rect 1383 623 1389 624
rect 1239 620 1298 622
rect 1239 619 1240 620
rect 1234 618 1240 619
rect 1296 618 1298 620
rect 1303 619 1309 620
rect 1303 618 1304 619
rect 1296 616 1304 618
rect 1303 615 1304 616
rect 1308 615 1309 619
rect 1374 619 1381 620
rect 1374 615 1375 619
rect 1380 615 1381 619
rect 1383 619 1384 623
rect 1388 622 1389 623
rect 1455 623 1461 624
rect 1388 620 1442 622
rect 1388 619 1389 620
rect 1383 618 1389 619
rect 1440 618 1442 620
rect 1447 619 1453 620
rect 1447 618 1448 619
rect 1440 616 1448 618
rect 1447 615 1448 616
rect 1452 615 1453 619
rect 1455 619 1456 623
rect 1460 622 1461 623
rect 1527 623 1533 624
rect 1460 620 1514 622
rect 1460 619 1461 620
rect 1455 618 1461 619
rect 1512 618 1514 620
rect 1519 619 1525 620
rect 1519 618 1520 619
rect 1512 616 1520 618
rect 1519 615 1520 616
rect 1524 615 1525 619
rect 1527 619 1528 623
rect 1532 622 1533 623
rect 1532 620 1586 622
rect 1532 619 1533 620
rect 1527 618 1533 619
rect 1584 618 1586 620
rect 1591 619 1597 620
rect 1591 618 1592 619
rect 1584 616 1592 618
rect 1591 615 1592 616
rect 1596 615 1597 619
rect 1639 619 1645 620
rect 1639 615 1640 619
rect 1644 618 1645 619
rect 1647 619 1653 620
rect 1647 618 1648 619
rect 1644 616 1648 618
rect 1644 615 1645 616
rect 1118 614 1119 615
rect 318 610 319 614
rect 323 610 324 614
rect 318 609 324 610
rect 366 610 367 614
rect 371 610 372 614
rect 366 609 372 610
rect 422 610 423 614
rect 427 610 428 614
rect 422 609 428 610
rect 470 610 471 614
rect 475 610 476 614
rect 470 609 476 610
rect 518 610 519 614
rect 523 610 524 614
rect 518 609 524 610
rect 566 610 567 614
rect 571 610 572 614
rect 566 609 572 610
rect 614 610 615 614
rect 619 610 620 614
rect 614 609 620 610
rect 662 610 663 614
rect 667 610 668 614
rect 662 609 668 610
rect 718 610 719 614
rect 723 610 724 614
rect 718 609 724 610
rect 774 610 775 614
rect 779 610 780 614
rect 774 609 780 610
rect 830 610 831 614
rect 835 610 836 614
rect 830 609 836 610
rect 894 610 895 614
rect 899 610 900 614
rect 894 609 900 610
rect 966 610 967 614
rect 971 610 972 614
rect 966 609 972 610
rect 1046 610 1047 614
rect 1051 610 1052 614
rect 1064 612 1119 614
rect 1118 611 1119 612
rect 1123 611 1124 615
rect 1118 610 1124 611
rect 1126 614 1132 615
rect 1143 614 1149 615
rect 1206 614 1212 615
rect 1223 614 1232 615
rect 1286 614 1292 615
rect 1303 614 1309 615
rect 1358 614 1364 615
rect 1374 614 1381 615
rect 1430 614 1436 615
rect 1447 614 1453 615
rect 1502 614 1508 615
rect 1519 614 1525 615
rect 1574 614 1580 615
rect 1591 614 1597 615
rect 1622 614 1628 615
rect 1639 614 1645 615
rect 1647 615 1648 616
rect 1652 615 1653 619
rect 1647 614 1653 615
rect 1662 616 1668 617
rect 1126 610 1127 614
rect 1131 610 1132 614
rect 1046 609 1052 610
rect 1126 609 1132 610
rect 1206 610 1207 614
rect 1211 610 1212 614
rect 1206 609 1212 610
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1286 609 1292 610
rect 1358 610 1359 614
rect 1363 610 1364 614
rect 1358 609 1364 610
rect 1430 610 1431 614
rect 1435 610 1436 614
rect 1430 609 1436 610
rect 1502 610 1503 614
rect 1507 610 1508 614
rect 1502 609 1508 610
rect 1574 610 1575 614
rect 1579 610 1580 614
rect 1574 609 1580 610
rect 1622 610 1623 614
rect 1627 610 1628 614
rect 1662 612 1663 616
rect 1667 612 1668 616
rect 1662 611 1668 612
rect 1622 609 1628 610
rect 263 603 269 604
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 263 599 264 603
rect 268 602 269 603
rect 276 602 290 604
rect 295 603 301 604
rect 268 600 278 602
rect 268 599 269 600
rect 263 598 269 599
rect 295 599 296 603
rect 300 602 301 603
rect 303 603 309 604
rect 303 602 304 603
rect 300 600 304 602
rect 300 599 301 600
rect 295 598 301 599
rect 303 599 304 600
rect 308 599 309 603
rect 303 598 309 599
rect 335 603 341 604
rect 335 599 336 603
rect 340 602 341 603
rect 351 603 357 604
rect 351 602 352 603
rect 340 600 352 602
rect 340 599 341 600
rect 335 598 341 599
rect 351 599 352 600
rect 356 599 357 603
rect 351 598 357 599
rect 383 603 389 604
rect 383 599 384 603
rect 388 602 389 603
rect 391 603 397 604
rect 391 602 392 603
rect 388 600 392 602
rect 388 599 389 600
rect 383 598 389 599
rect 391 599 392 600
rect 396 599 397 603
rect 391 598 397 599
rect 439 603 445 604
rect 439 599 440 603
rect 444 602 445 603
rect 447 603 453 604
rect 447 602 448 603
rect 444 600 448 602
rect 444 599 445 600
rect 439 598 445 599
rect 447 599 448 600
rect 452 599 453 603
rect 447 598 453 599
rect 482 603 493 604
rect 482 599 483 603
rect 487 599 488 603
rect 492 599 493 603
rect 482 598 493 599
rect 535 603 541 604
rect 535 599 536 603
rect 540 602 541 603
rect 543 603 549 604
rect 543 602 544 603
rect 540 600 544 602
rect 540 599 541 600
rect 535 598 541 599
rect 543 599 544 600
rect 548 599 549 603
rect 543 598 549 599
rect 583 603 589 604
rect 583 599 584 603
rect 588 602 589 603
rect 591 603 597 604
rect 591 602 592 603
rect 588 600 592 602
rect 588 599 589 600
rect 583 598 589 599
rect 591 599 592 600
rect 596 599 597 603
rect 591 598 597 599
rect 631 603 637 604
rect 631 599 632 603
rect 636 602 637 603
rect 639 603 645 604
rect 639 602 640 603
rect 636 600 640 602
rect 636 599 637 600
rect 631 598 637 599
rect 639 599 640 600
rect 644 599 645 603
rect 639 598 645 599
rect 679 603 685 604
rect 679 599 680 603
rect 684 602 685 603
rect 687 603 693 604
rect 687 602 688 603
rect 684 600 688 602
rect 684 599 685 600
rect 679 598 685 599
rect 687 599 688 600
rect 692 599 693 603
rect 687 598 693 599
rect 735 603 741 604
rect 735 599 736 603
rect 740 602 741 603
rect 743 603 749 604
rect 743 602 744 603
rect 740 600 744 602
rect 740 599 741 600
rect 735 598 741 599
rect 743 599 744 600
rect 748 599 749 603
rect 791 603 797 604
rect 791 602 792 603
rect 743 598 749 599
rect 784 600 792 602
rect 110 594 116 595
rect 246 597 252 598
rect 246 593 247 597
rect 251 593 252 597
rect 246 592 252 593
rect 278 597 284 598
rect 278 593 279 597
rect 283 593 284 597
rect 278 592 284 593
rect 318 597 324 598
rect 318 593 319 597
rect 323 593 324 597
rect 318 592 324 593
rect 366 597 372 598
rect 366 593 367 597
rect 371 593 372 597
rect 366 592 372 593
rect 422 597 428 598
rect 422 593 423 597
rect 427 593 428 597
rect 422 592 428 593
rect 470 597 476 598
rect 470 593 471 597
rect 475 593 476 597
rect 470 592 476 593
rect 518 597 524 598
rect 518 593 519 597
rect 523 593 524 597
rect 518 592 524 593
rect 566 597 572 598
rect 566 593 567 597
rect 571 593 572 597
rect 566 592 572 593
rect 614 597 620 598
rect 614 593 615 597
rect 619 593 620 597
rect 614 592 620 593
rect 662 597 668 598
rect 662 593 663 597
rect 667 593 668 597
rect 662 592 668 593
rect 718 597 724 598
rect 718 593 719 597
rect 723 593 724 597
rect 718 592 724 593
rect 774 597 780 598
rect 774 593 775 597
rect 779 593 780 597
rect 774 592 780 593
rect 262 591 268 592
rect 262 587 263 591
rect 267 590 268 591
rect 578 591 584 592
rect 267 588 475 590
rect 267 587 268 588
rect 262 586 268 587
rect 166 583 172 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 166 579 167 583
rect 171 579 172 583
rect 166 578 172 579
rect 214 583 220 584
rect 214 579 215 583
rect 219 579 220 583
rect 214 578 220 579
rect 270 583 276 584
rect 270 579 271 583
rect 275 579 276 583
rect 270 578 276 579
rect 334 583 340 584
rect 334 579 335 583
rect 339 579 340 583
rect 334 578 340 579
rect 406 583 412 584
rect 406 579 407 583
rect 411 579 412 583
rect 406 578 412 579
rect 110 576 116 577
rect 183 575 189 576
rect 183 571 184 575
rect 188 574 189 575
rect 231 575 237 576
rect 188 572 226 574
rect 188 571 189 572
rect 183 570 189 571
rect 166 566 172 567
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 166 562 167 566
rect 171 562 172 566
rect 166 561 172 562
rect 214 566 220 567
rect 214 562 215 566
rect 219 562 220 566
rect 214 561 220 562
rect 110 559 116 560
rect 183 559 189 560
rect 183 555 184 559
rect 188 555 189 559
rect 224 558 226 572
rect 231 571 232 575
rect 236 574 237 575
rect 287 575 293 576
rect 236 572 262 574
rect 236 571 237 572
rect 231 570 237 571
rect 231 559 237 560
rect 231 558 232 559
rect 224 556 232 558
rect 183 554 189 555
rect 231 555 232 556
rect 236 555 237 559
rect 260 558 262 572
rect 287 571 288 575
rect 292 574 293 575
rect 351 575 357 576
rect 292 572 321 574
rect 292 571 293 572
rect 287 570 293 571
rect 270 566 276 567
rect 270 562 271 566
rect 275 562 276 566
rect 270 561 276 562
rect 287 559 293 560
rect 287 558 288 559
rect 260 556 288 558
rect 231 554 237 555
rect 287 555 288 556
rect 292 555 293 559
rect 319 558 321 572
rect 351 571 352 575
rect 356 574 357 575
rect 423 575 429 576
rect 356 572 390 574
rect 356 571 357 572
rect 351 570 357 571
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 351 559 357 560
rect 351 558 352 559
rect 319 556 352 558
rect 287 554 293 555
rect 351 555 352 556
rect 356 555 357 559
rect 388 558 390 572
rect 423 571 424 575
rect 428 574 429 575
rect 473 574 475 588
rect 578 587 579 591
rect 583 590 584 591
rect 784 590 786 600
rect 791 599 792 600
rect 796 599 797 603
rect 791 598 797 599
rect 847 603 853 604
rect 847 599 848 603
rect 852 602 853 603
rect 855 603 861 604
rect 855 602 856 603
rect 852 600 856 602
rect 852 599 853 600
rect 847 598 853 599
rect 855 599 856 600
rect 860 599 861 603
rect 855 598 861 599
rect 911 603 917 604
rect 911 599 912 603
rect 916 602 917 603
rect 919 603 925 604
rect 919 602 920 603
rect 916 600 920 602
rect 916 599 917 600
rect 911 598 917 599
rect 919 599 920 600
rect 924 599 925 603
rect 919 598 925 599
rect 978 603 989 604
rect 978 599 979 603
rect 983 599 984 603
rect 988 599 989 603
rect 978 598 989 599
rect 1063 603 1069 604
rect 1063 599 1064 603
rect 1068 602 1069 603
rect 1071 603 1077 604
rect 1071 602 1072 603
rect 1068 600 1072 602
rect 1068 599 1069 600
rect 1063 598 1069 599
rect 1071 599 1072 600
rect 1076 599 1077 603
rect 1071 598 1077 599
rect 1142 603 1149 604
rect 1142 599 1143 603
rect 1148 599 1149 603
rect 1142 598 1149 599
rect 1223 603 1229 604
rect 1223 599 1224 603
rect 1228 602 1229 603
rect 1234 603 1240 604
rect 1234 602 1235 603
rect 1228 600 1235 602
rect 1228 599 1229 600
rect 1223 598 1229 599
rect 1234 599 1235 600
rect 1239 599 1240 603
rect 1234 598 1240 599
rect 1298 603 1309 604
rect 1298 599 1299 603
rect 1303 599 1304 603
rect 1308 599 1309 603
rect 1298 598 1309 599
rect 1375 603 1381 604
rect 1375 599 1376 603
rect 1380 602 1381 603
rect 1383 603 1389 604
rect 1383 602 1384 603
rect 1380 600 1384 602
rect 1380 599 1381 600
rect 1375 598 1381 599
rect 1383 599 1384 600
rect 1388 599 1389 603
rect 1383 598 1389 599
rect 1447 603 1453 604
rect 1447 599 1448 603
rect 1452 602 1453 603
rect 1455 603 1461 604
rect 1455 602 1456 603
rect 1452 600 1456 602
rect 1452 599 1453 600
rect 1447 598 1453 599
rect 1455 599 1456 600
rect 1460 599 1461 603
rect 1455 598 1461 599
rect 1519 603 1525 604
rect 1519 599 1520 603
rect 1524 602 1525 603
rect 1527 603 1533 604
rect 1527 602 1528 603
rect 1524 600 1528 602
rect 1524 599 1525 600
rect 1519 598 1525 599
rect 1527 599 1528 600
rect 1532 599 1533 603
rect 1527 598 1533 599
rect 1590 603 1597 604
rect 1590 599 1591 603
rect 1596 599 1597 603
rect 1590 598 1597 599
rect 1638 603 1645 604
rect 1638 599 1639 603
rect 1644 599 1645 603
rect 1638 598 1645 599
rect 1662 599 1668 600
rect 830 597 836 598
rect 830 593 831 597
rect 835 593 836 597
rect 830 592 836 593
rect 894 597 900 598
rect 894 593 895 597
rect 899 593 900 597
rect 894 592 900 593
rect 966 597 972 598
rect 966 593 967 597
rect 971 593 972 597
rect 966 592 972 593
rect 1046 597 1052 598
rect 1046 593 1047 597
rect 1051 593 1052 597
rect 1046 592 1052 593
rect 1126 597 1132 598
rect 1126 593 1127 597
rect 1131 593 1132 597
rect 1126 592 1132 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1286 597 1292 598
rect 1286 593 1287 597
rect 1291 593 1292 597
rect 1286 592 1292 593
rect 1358 597 1364 598
rect 1358 593 1359 597
rect 1363 593 1364 597
rect 1358 592 1364 593
rect 1430 597 1436 598
rect 1430 593 1431 597
rect 1435 593 1436 597
rect 1430 592 1436 593
rect 1502 597 1508 598
rect 1502 593 1503 597
rect 1507 593 1508 597
rect 1502 592 1508 593
rect 1574 597 1580 598
rect 1574 593 1575 597
rect 1579 593 1580 597
rect 1574 592 1580 593
rect 1622 597 1628 598
rect 1622 593 1623 597
rect 1627 593 1628 597
rect 1662 595 1663 599
rect 1667 595 1668 599
rect 1662 594 1668 595
rect 1622 592 1628 593
rect 583 588 786 590
rect 1374 591 1380 592
rect 583 587 584 588
rect 578 586 584 587
rect 1374 587 1375 591
rect 1379 590 1380 591
rect 1379 588 1570 590
rect 1379 587 1380 588
rect 1374 586 1380 587
rect 486 583 492 584
rect 486 579 487 583
rect 491 579 492 583
rect 486 578 492 579
rect 558 583 564 584
rect 558 579 559 583
rect 563 579 564 583
rect 558 578 564 579
rect 630 583 636 584
rect 630 579 631 583
rect 635 579 636 583
rect 630 578 636 579
rect 702 583 708 584
rect 702 579 703 583
rect 707 579 708 583
rect 702 578 708 579
rect 766 583 772 584
rect 766 579 767 583
rect 771 579 772 583
rect 766 578 772 579
rect 822 583 828 584
rect 822 579 823 583
rect 827 579 828 583
rect 822 578 828 579
rect 878 583 884 584
rect 878 579 879 583
rect 883 579 884 583
rect 878 578 884 579
rect 934 583 940 584
rect 934 579 935 583
rect 939 579 940 583
rect 934 578 940 579
rect 990 583 996 584
rect 990 579 991 583
rect 995 579 996 583
rect 990 578 996 579
rect 1046 583 1052 584
rect 1046 579 1047 583
rect 1051 579 1052 583
rect 1046 578 1052 579
rect 1102 583 1108 584
rect 1102 579 1103 583
rect 1107 579 1108 583
rect 1102 578 1108 579
rect 1158 583 1164 584
rect 1158 579 1159 583
rect 1163 579 1164 583
rect 1158 578 1164 579
rect 1214 583 1220 584
rect 1214 579 1215 583
rect 1219 579 1220 583
rect 1214 578 1220 579
rect 1270 583 1276 584
rect 1270 579 1271 583
rect 1275 579 1276 583
rect 1270 578 1276 579
rect 1326 583 1332 584
rect 1326 579 1327 583
rect 1331 579 1332 583
rect 1326 578 1332 579
rect 1382 583 1388 584
rect 1382 579 1383 583
rect 1387 579 1388 583
rect 1382 578 1388 579
rect 1446 583 1452 584
rect 1446 579 1447 583
rect 1451 579 1452 583
rect 1446 578 1452 579
rect 1510 583 1516 584
rect 1510 579 1511 583
rect 1515 579 1516 583
rect 1510 578 1516 579
rect 503 575 509 576
rect 503 574 504 575
rect 428 572 466 574
rect 473 572 504 574
rect 428 571 429 572
rect 423 570 429 571
rect 406 566 412 567
rect 406 562 407 566
rect 411 562 412 566
rect 406 561 412 562
rect 423 559 429 560
rect 423 558 424 559
rect 388 556 424 558
rect 351 554 357 555
rect 423 555 424 556
rect 428 555 429 559
rect 464 558 466 572
rect 503 571 504 572
rect 508 571 509 575
rect 503 570 509 571
rect 575 575 581 576
rect 575 571 576 575
rect 580 574 581 575
rect 647 575 653 576
rect 580 572 614 574
rect 580 571 581 572
rect 575 570 581 571
rect 486 566 492 567
rect 486 562 487 566
rect 491 562 492 566
rect 486 561 492 562
rect 558 566 564 567
rect 558 562 559 566
rect 563 562 564 566
rect 558 561 564 562
rect 503 559 509 560
rect 503 558 504 559
rect 464 556 504 558
rect 423 554 429 555
rect 503 555 504 556
rect 508 555 509 559
rect 503 554 509 555
rect 575 559 584 560
rect 575 555 576 559
rect 583 555 584 559
rect 612 558 614 572
rect 647 571 648 575
rect 652 574 653 575
rect 719 575 725 576
rect 652 572 714 574
rect 652 571 653 572
rect 647 570 653 571
rect 630 566 636 567
rect 630 562 631 566
rect 635 562 636 566
rect 630 561 636 562
rect 702 566 708 567
rect 702 562 703 566
rect 707 562 708 566
rect 702 561 708 562
rect 647 559 653 560
rect 647 558 648 559
rect 612 556 648 558
rect 575 554 584 555
rect 647 555 648 556
rect 652 555 653 559
rect 712 558 714 572
rect 719 571 720 575
rect 724 574 725 575
rect 783 575 789 576
rect 724 572 754 574
rect 724 571 725 572
rect 719 570 725 571
rect 719 559 725 560
rect 719 558 720 559
rect 712 556 720 558
rect 647 554 653 555
rect 719 555 720 556
rect 724 555 725 559
rect 752 558 754 572
rect 783 571 784 575
rect 788 574 789 575
rect 806 575 812 576
rect 806 574 807 575
rect 788 572 807 574
rect 788 571 789 572
rect 783 570 789 571
rect 806 571 807 572
rect 811 571 812 575
rect 806 570 812 571
rect 839 575 845 576
rect 839 571 840 575
rect 844 574 845 575
rect 894 575 901 576
rect 844 572 870 574
rect 844 571 845 572
rect 839 570 845 571
rect 766 566 772 567
rect 766 562 767 566
rect 771 562 772 566
rect 766 561 772 562
rect 822 566 828 567
rect 822 562 823 566
rect 827 562 828 566
rect 822 561 828 562
rect 783 559 789 560
rect 783 558 784 559
rect 752 556 784 558
rect 719 554 725 555
rect 783 555 784 556
rect 788 555 789 559
rect 783 554 789 555
rect 839 559 845 560
rect 839 555 840 559
rect 844 558 845 559
rect 868 558 870 572
rect 894 571 895 575
rect 900 571 901 575
rect 894 570 901 571
rect 903 575 909 576
rect 903 571 904 575
rect 908 574 909 575
rect 951 575 957 576
rect 951 574 952 575
rect 908 572 952 574
rect 908 571 909 572
rect 903 570 909 571
rect 951 571 952 572
rect 956 571 957 575
rect 951 570 957 571
rect 1007 575 1013 576
rect 1007 571 1008 575
rect 1012 574 1013 575
rect 1063 575 1069 576
rect 1012 572 1038 574
rect 1012 571 1013 572
rect 1007 570 1013 571
rect 878 566 884 567
rect 878 562 879 566
rect 883 562 884 566
rect 878 561 884 562
rect 934 566 940 567
rect 934 562 935 566
rect 939 562 940 566
rect 934 561 940 562
rect 990 566 996 567
rect 990 562 991 566
rect 995 562 996 566
rect 990 561 996 562
rect 895 559 901 560
rect 895 558 896 559
rect 844 556 866 558
rect 868 556 896 558
rect 844 555 845 556
rect 839 554 845 555
rect 185 550 187 554
rect 342 551 348 552
rect 342 550 343 551
rect 185 548 343 550
rect 342 547 343 548
rect 347 547 348 551
rect 864 550 866 556
rect 895 555 896 556
rect 900 555 901 559
rect 895 554 901 555
rect 951 559 957 560
rect 951 555 952 559
rect 956 558 957 559
rect 978 559 984 560
rect 978 558 979 559
rect 956 556 979 558
rect 956 555 957 556
rect 951 554 957 555
rect 978 555 979 556
rect 983 555 984 559
rect 978 554 984 555
rect 1007 559 1013 560
rect 1007 555 1008 559
rect 1012 558 1013 559
rect 1022 559 1028 560
rect 1022 558 1023 559
rect 1012 556 1023 558
rect 1012 555 1013 556
rect 1007 554 1013 555
rect 1022 555 1023 556
rect 1027 555 1028 559
rect 1036 558 1038 572
rect 1063 571 1064 575
rect 1068 574 1069 575
rect 1118 575 1125 576
rect 1068 572 1094 574
rect 1068 571 1069 572
rect 1063 570 1069 571
rect 1046 566 1052 567
rect 1046 562 1047 566
rect 1051 562 1052 566
rect 1046 561 1052 562
rect 1063 559 1069 560
rect 1063 558 1064 559
rect 1036 556 1064 558
rect 1022 554 1028 555
rect 1063 555 1064 556
rect 1068 555 1069 559
rect 1092 558 1094 572
rect 1118 571 1119 575
rect 1124 571 1125 575
rect 1118 570 1125 571
rect 1175 575 1181 576
rect 1175 571 1176 575
rect 1180 574 1181 575
rect 1198 575 1204 576
rect 1198 574 1199 575
rect 1180 572 1199 574
rect 1180 571 1181 572
rect 1175 570 1181 571
rect 1198 571 1199 572
rect 1203 571 1204 575
rect 1231 575 1237 576
rect 1231 574 1232 575
rect 1198 570 1204 571
rect 1208 572 1232 574
rect 1102 566 1108 567
rect 1102 562 1103 566
rect 1107 562 1108 566
rect 1102 561 1108 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 1119 559 1125 560
rect 1119 558 1120 559
rect 1092 556 1120 558
rect 1063 554 1069 555
rect 1119 555 1120 556
rect 1124 555 1125 559
rect 1119 554 1125 555
rect 1175 559 1181 560
rect 1175 555 1176 559
rect 1180 558 1181 559
rect 1208 558 1210 572
rect 1231 571 1232 572
rect 1236 571 1237 575
rect 1287 575 1293 576
rect 1287 574 1288 575
rect 1231 570 1237 571
rect 1260 572 1288 574
rect 1214 566 1220 567
rect 1214 562 1215 566
rect 1219 562 1220 566
rect 1214 561 1220 562
rect 1180 556 1210 558
rect 1231 559 1237 560
rect 1180 555 1181 556
rect 1175 554 1181 555
rect 1231 555 1232 559
rect 1236 558 1237 559
rect 1260 558 1262 572
rect 1287 571 1288 572
rect 1292 571 1293 575
rect 1287 570 1293 571
rect 1343 575 1349 576
rect 1343 571 1344 575
rect 1348 574 1349 575
rect 1399 575 1405 576
rect 1348 572 1394 574
rect 1348 571 1349 572
rect 1343 570 1349 571
rect 1270 566 1276 567
rect 1270 562 1271 566
rect 1275 562 1276 566
rect 1270 561 1276 562
rect 1326 566 1332 567
rect 1326 562 1327 566
rect 1331 562 1332 566
rect 1326 561 1332 562
rect 1382 566 1388 567
rect 1382 562 1383 566
rect 1387 562 1388 566
rect 1382 561 1388 562
rect 1236 556 1262 558
rect 1287 559 1293 560
rect 1236 555 1237 556
rect 1231 554 1237 555
rect 1287 555 1288 559
rect 1292 558 1293 559
rect 1298 559 1304 560
rect 1298 558 1299 559
rect 1292 556 1299 558
rect 1292 555 1293 556
rect 1287 554 1293 555
rect 1298 555 1299 556
rect 1303 555 1304 559
rect 1298 554 1304 555
rect 1343 559 1349 560
rect 1343 555 1344 559
rect 1348 555 1349 559
rect 1392 558 1394 572
rect 1399 571 1400 575
rect 1404 574 1405 575
rect 1463 575 1469 576
rect 1404 572 1434 574
rect 1404 571 1405 572
rect 1399 570 1405 571
rect 1399 559 1405 560
rect 1399 558 1400 559
rect 1392 556 1400 558
rect 1343 554 1349 555
rect 1399 555 1400 556
rect 1404 555 1405 559
rect 1432 558 1434 572
rect 1463 571 1464 575
rect 1468 574 1469 575
rect 1527 575 1533 576
rect 1468 572 1522 574
rect 1468 571 1469 572
rect 1463 570 1469 571
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1510 566 1516 567
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1463 559 1469 560
rect 1463 558 1464 559
rect 1432 556 1464 558
rect 1399 554 1405 555
rect 1463 555 1464 556
rect 1468 555 1469 559
rect 1520 558 1522 572
rect 1527 571 1528 575
rect 1532 574 1533 575
rect 1568 574 1570 588
rect 1574 583 1580 584
rect 1574 579 1575 583
rect 1579 579 1580 583
rect 1574 578 1580 579
rect 1622 583 1628 584
rect 1622 579 1623 583
rect 1627 579 1628 583
rect 1622 578 1628 579
rect 1662 581 1668 582
rect 1662 577 1663 581
rect 1667 577 1668 581
rect 1662 576 1668 577
rect 1591 575 1597 576
rect 1591 574 1592 575
rect 1532 572 1562 574
rect 1568 572 1592 574
rect 1532 571 1533 572
rect 1527 570 1533 571
rect 1527 559 1533 560
rect 1527 558 1528 559
rect 1520 556 1528 558
rect 1463 554 1469 555
rect 1527 555 1528 556
rect 1532 555 1533 559
rect 1560 558 1562 572
rect 1591 571 1592 572
rect 1596 571 1597 575
rect 1591 570 1597 571
rect 1639 575 1645 576
rect 1639 571 1640 575
rect 1644 574 1645 575
rect 1647 575 1653 576
rect 1647 574 1648 575
rect 1644 572 1648 574
rect 1644 571 1645 572
rect 1639 570 1645 571
rect 1647 571 1648 572
rect 1652 571 1653 575
rect 1647 570 1653 571
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1622 566 1628 567
rect 1622 562 1623 566
rect 1627 562 1628 566
rect 1622 561 1628 562
rect 1662 564 1668 565
rect 1662 560 1663 564
rect 1667 560 1668 564
rect 1591 559 1597 560
rect 1591 558 1592 559
rect 1560 556 1592 558
rect 1527 554 1533 555
rect 1591 555 1592 556
rect 1596 555 1597 559
rect 1591 554 1597 555
rect 1638 559 1645 560
rect 1662 559 1668 560
rect 1638 555 1639 559
rect 1644 555 1645 559
rect 1638 554 1645 555
rect 903 551 909 552
rect 903 550 904 551
rect 864 548 904 550
rect 342 546 348 547
rect 510 547 516 548
rect 510 546 511 547
rect 392 544 511 546
rect 255 539 261 540
rect 160 536 187 538
rect 225 536 251 538
rect 150 535 157 536
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 150 531 151 535
rect 156 531 157 535
rect 110 527 116 528
rect 134 530 140 531
rect 150 530 157 531
rect 134 526 135 530
rect 139 526 140 530
rect 134 525 140 526
rect 151 519 157 520
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 151 515 152 519
rect 156 518 157 519
rect 160 518 162 536
rect 183 535 189 536
rect 183 531 184 535
rect 188 531 189 535
rect 215 535 221 536
rect 215 534 216 535
rect 208 532 216 534
rect 166 530 172 531
rect 183 530 189 531
rect 198 530 204 531
rect 166 526 167 530
rect 171 526 172 530
rect 166 525 172 526
rect 198 526 199 530
rect 203 526 204 530
rect 198 525 204 526
rect 208 520 210 532
rect 215 531 216 532
rect 220 531 221 535
rect 215 530 221 531
rect 156 516 162 518
rect 183 519 189 520
rect 156 515 157 516
rect 151 514 157 515
rect 183 515 184 519
rect 188 518 189 519
rect 196 518 210 520
rect 215 519 221 520
rect 188 516 198 518
rect 188 515 189 516
rect 183 514 189 515
rect 215 515 216 519
rect 220 518 221 519
rect 225 518 227 536
rect 247 535 253 536
rect 247 531 248 535
rect 252 531 253 535
rect 255 535 256 539
rect 260 538 261 539
rect 303 539 309 540
rect 260 536 290 538
rect 260 535 261 536
rect 255 534 261 535
rect 288 534 290 536
rect 295 535 301 536
rect 295 534 296 535
rect 288 532 296 534
rect 295 531 296 532
rect 300 531 301 535
rect 303 535 304 539
rect 308 538 309 539
rect 308 536 347 538
rect 392 536 394 544
rect 510 543 511 544
rect 515 543 516 547
rect 830 547 836 548
rect 830 546 831 547
rect 705 544 831 546
rect 510 542 516 543
rect 638 543 644 544
rect 638 542 639 543
rect 617 540 639 542
rect 399 539 405 540
rect 308 535 309 536
rect 303 534 309 535
rect 343 535 349 536
rect 343 531 344 535
rect 348 531 349 535
rect 391 535 397 536
rect 391 531 392 535
rect 396 531 397 535
rect 399 535 400 539
rect 404 538 405 539
rect 404 536 442 538
rect 404 535 405 536
rect 399 534 405 535
rect 440 534 442 536
rect 447 535 453 536
rect 447 534 448 535
rect 440 532 448 534
rect 447 531 448 532
rect 452 531 453 535
rect 511 535 517 536
rect 511 531 512 535
rect 516 534 517 535
rect 575 535 581 536
rect 516 532 546 534
rect 516 531 517 532
rect 230 530 236 531
rect 247 530 253 531
rect 278 530 284 531
rect 295 530 301 531
rect 326 530 332 531
rect 343 530 349 531
rect 374 530 380 531
rect 391 530 397 531
rect 430 530 436 531
rect 447 530 453 531
rect 494 530 500 531
rect 511 530 517 531
rect 230 526 231 530
rect 235 526 236 530
rect 230 525 236 526
rect 278 526 279 530
rect 283 526 284 530
rect 278 525 284 526
rect 326 526 327 530
rect 331 526 332 530
rect 326 525 332 526
rect 374 526 375 530
rect 379 526 380 530
rect 374 525 380 526
rect 430 526 431 530
rect 435 526 436 530
rect 430 525 436 526
rect 494 526 495 530
rect 499 526 500 530
rect 494 525 500 526
rect 544 522 546 532
rect 575 531 576 535
rect 580 534 581 535
rect 617 534 619 540
rect 638 539 639 540
rect 643 539 644 543
rect 638 538 644 539
rect 705 536 707 544
rect 830 543 831 544
rect 835 543 836 547
rect 903 547 904 548
rect 908 547 909 551
rect 1345 550 1347 554
rect 1526 551 1532 552
rect 1526 550 1527 551
rect 1345 548 1527 550
rect 903 546 909 547
rect 1526 547 1527 548
rect 1531 547 1532 551
rect 1526 546 1532 547
rect 830 542 836 543
rect 711 539 717 540
rect 580 532 619 534
rect 630 535 636 536
rect 580 531 581 532
rect 630 531 631 535
rect 635 534 636 535
rect 639 535 645 536
rect 639 534 640 535
rect 635 532 640 534
rect 635 531 636 532
rect 558 530 564 531
rect 575 530 581 531
rect 622 530 628 531
rect 630 530 636 531
rect 639 531 640 532
rect 644 531 645 535
rect 703 535 709 536
rect 703 531 704 535
rect 708 531 709 535
rect 711 535 712 539
rect 716 538 717 539
rect 806 539 812 540
rect 716 536 771 538
rect 716 535 717 536
rect 711 534 717 535
rect 767 535 773 536
rect 767 531 768 535
rect 772 531 773 535
rect 806 535 807 539
rect 811 538 812 539
rect 903 539 909 540
rect 811 536 835 538
rect 811 535 812 536
rect 806 534 812 535
rect 831 535 837 536
rect 831 531 832 535
rect 836 531 837 535
rect 894 535 901 536
rect 894 531 895 535
rect 900 531 901 535
rect 903 535 904 539
rect 908 538 909 539
rect 967 539 973 540
rect 908 536 954 538
rect 908 535 909 536
rect 903 534 909 535
rect 952 534 954 536
rect 959 535 965 536
rect 959 534 960 535
rect 952 532 960 534
rect 959 531 960 532
rect 964 531 965 535
rect 967 535 968 539
rect 972 538 973 539
rect 1255 539 1261 540
rect 972 536 1018 538
rect 1120 536 1139 538
rect 1159 536 1194 538
rect 972 535 973 536
rect 967 534 973 535
rect 1016 534 1018 536
rect 1023 535 1029 536
rect 1023 534 1024 535
rect 1016 532 1024 534
rect 1023 531 1024 532
rect 1028 531 1029 535
rect 1087 535 1093 536
rect 1087 531 1088 535
rect 1092 534 1093 535
rect 1120 534 1122 536
rect 1092 532 1122 534
rect 1092 531 1093 532
rect 639 530 645 531
rect 686 530 692 531
rect 703 530 709 531
rect 750 530 756 531
rect 767 530 773 531
rect 814 530 820 531
rect 831 530 837 531
rect 878 530 884 531
rect 894 530 901 531
rect 942 530 948 531
rect 959 530 965 531
rect 1006 530 1012 531
rect 1023 530 1029 531
rect 1070 530 1076 531
rect 1087 530 1093 531
rect 1126 530 1132 531
rect 558 526 559 530
rect 563 526 564 530
rect 558 525 564 526
rect 622 526 623 530
rect 627 526 628 530
rect 622 525 628 526
rect 686 526 687 530
rect 691 526 692 530
rect 686 525 692 526
rect 750 526 751 530
rect 755 526 756 530
rect 750 525 756 526
rect 814 526 815 530
rect 819 526 820 530
rect 814 525 820 526
rect 878 526 879 530
rect 883 526 884 530
rect 878 525 884 526
rect 942 526 943 530
rect 947 526 948 530
rect 942 525 948 526
rect 1006 526 1007 530
rect 1011 526 1012 530
rect 1006 525 1012 526
rect 1070 526 1071 530
rect 1075 526 1076 530
rect 1070 525 1076 526
rect 1126 526 1127 530
rect 1131 526 1132 530
rect 1126 525 1132 526
rect 544 520 558 522
rect 220 516 227 518
rect 247 519 253 520
rect 220 515 221 516
rect 215 514 221 515
rect 247 515 248 519
rect 252 518 253 519
rect 255 519 261 520
rect 255 518 256 519
rect 252 516 256 518
rect 252 515 253 516
rect 247 514 253 515
rect 255 515 256 516
rect 260 515 261 519
rect 255 514 261 515
rect 295 519 301 520
rect 295 515 296 519
rect 300 518 301 519
rect 303 519 309 520
rect 303 518 304 519
rect 300 516 304 518
rect 300 515 301 516
rect 295 514 301 515
rect 303 515 304 516
rect 308 515 309 519
rect 303 514 309 515
rect 342 519 349 520
rect 342 515 343 519
rect 348 515 349 519
rect 342 514 349 515
rect 391 519 397 520
rect 391 515 392 519
rect 396 518 397 519
rect 399 519 405 520
rect 399 518 400 519
rect 396 516 400 518
rect 396 515 397 516
rect 391 514 397 515
rect 399 515 400 516
rect 404 515 405 519
rect 399 514 405 515
rect 447 519 453 520
rect 447 515 448 519
rect 452 518 453 519
rect 486 519 492 520
rect 486 518 487 519
rect 452 516 487 518
rect 452 515 453 516
rect 447 514 453 515
rect 486 515 487 516
rect 491 515 492 519
rect 486 514 492 515
rect 510 519 517 520
rect 510 515 511 519
rect 516 515 517 519
rect 556 518 570 520
rect 575 519 581 520
rect 575 518 576 519
rect 568 516 576 518
rect 510 514 517 515
rect 575 515 576 516
rect 580 515 581 519
rect 575 514 581 515
rect 638 519 645 520
rect 638 515 639 519
rect 644 515 645 519
rect 638 514 645 515
rect 703 519 709 520
rect 703 515 704 519
rect 708 518 709 519
rect 711 519 717 520
rect 711 518 712 519
rect 708 516 712 518
rect 708 515 709 516
rect 703 514 709 515
rect 711 515 712 516
rect 716 515 717 519
rect 711 514 717 515
rect 767 519 773 520
rect 767 515 768 519
rect 772 518 773 519
rect 790 519 796 520
rect 790 518 791 519
rect 772 516 791 518
rect 772 515 773 516
rect 767 514 773 515
rect 790 515 791 516
rect 795 515 796 519
rect 790 514 796 515
rect 830 519 837 520
rect 830 515 831 519
rect 836 515 837 519
rect 830 514 837 515
rect 895 519 901 520
rect 895 515 896 519
rect 900 518 901 519
rect 903 519 909 520
rect 903 518 904 519
rect 900 516 904 518
rect 900 515 901 516
rect 895 514 901 515
rect 903 515 904 516
rect 908 515 909 519
rect 903 514 909 515
rect 959 519 965 520
rect 959 515 960 519
rect 964 518 965 519
rect 967 519 973 520
rect 967 518 968 519
rect 964 516 968 518
rect 964 515 965 516
rect 959 514 965 515
rect 967 515 968 516
rect 972 515 973 519
rect 967 514 973 515
rect 1022 519 1029 520
rect 1022 515 1023 519
rect 1028 515 1029 519
rect 1087 519 1093 520
rect 1087 518 1088 519
rect 1022 514 1029 515
rect 1080 516 1088 518
rect 110 510 116 511
rect 134 513 140 514
rect 134 509 135 513
rect 139 509 140 513
rect 134 508 140 509
rect 166 513 172 514
rect 166 509 167 513
rect 171 509 172 513
rect 166 508 172 509
rect 198 513 204 514
rect 198 509 199 513
rect 203 509 204 513
rect 198 508 204 509
rect 230 513 236 514
rect 230 509 231 513
rect 235 509 236 513
rect 230 508 236 509
rect 278 513 284 514
rect 278 509 279 513
rect 283 509 284 513
rect 278 508 284 509
rect 326 513 332 514
rect 326 509 327 513
rect 331 509 332 513
rect 326 508 332 509
rect 374 513 380 514
rect 374 509 375 513
rect 379 509 380 513
rect 374 508 380 509
rect 430 513 436 514
rect 430 509 431 513
rect 435 509 436 513
rect 430 508 436 509
rect 494 513 500 514
rect 494 509 495 513
rect 499 509 500 513
rect 494 508 500 509
rect 558 513 564 514
rect 558 509 559 513
rect 563 509 564 513
rect 558 508 564 509
rect 622 513 628 514
rect 622 509 623 513
rect 627 509 628 513
rect 622 508 628 509
rect 686 513 692 514
rect 686 509 687 513
rect 691 509 692 513
rect 686 508 692 509
rect 750 513 756 514
rect 750 509 751 513
rect 755 509 756 513
rect 750 508 756 509
rect 814 513 820 514
rect 814 509 815 513
rect 819 509 820 513
rect 814 508 820 509
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 878 508 884 509
rect 942 513 948 514
rect 942 509 943 513
rect 947 509 948 513
rect 942 508 948 509
rect 1006 513 1012 514
rect 1006 509 1007 513
rect 1011 509 1012 513
rect 1006 508 1012 509
rect 1070 513 1076 514
rect 1070 509 1071 513
rect 1075 509 1076 513
rect 1070 508 1076 509
rect 150 507 156 508
rect 150 503 151 507
rect 155 506 156 507
rect 950 507 956 508
rect 155 504 250 506
rect 155 503 156 504
rect 150 502 156 503
rect 134 499 140 500
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 134 495 135 499
rect 139 495 140 499
rect 134 494 140 495
rect 166 499 172 500
rect 166 495 167 499
rect 171 495 172 499
rect 166 494 172 495
rect 198 499 204 500
rect 198 495 199 499
rect 203 495 204 499
rect 198 494 204 495
rect 238 499 244 500
rect 238 495 239 499
rect 243 495 244 499
rect 238 494 244 495
rect 110 492 116 493
rect 151 491 157 492
rect 151 487 152 491
rect 156 490 157 491
rect 183 491 189 492
rect 156 488 178 490
rect 156 487 157 488
rect 151 486 157 487
rect 134 482 140 483
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 134 478 135 482
rect 139 478 140 482
rect 134 477 140 478
rect 166 482 172 483
rect 166 478 167 482
rect 171 478 172 482
rect 166 477 172 478
rect 110 475 116 476
rect 151 475 157 476
rect 151 471 152 475
rect 156 471 157 475
rect 176 474 178 488
rect 183 487 184 491
rect 188 490 189 491
rect 215 491 221 492
rect 188 488 210 490
rect 188 487 189 488
rect 183 486 189 487
rect 198 482 204 483
rect 198 478 199 482
rect 203 478 204 482
rect 198 477 204 478
rect 183 475 189 476
rect 183 474 184 475
rect 176 472 184 474
rect 151 470 157 471
rect 183 471 184 472
rect 188 471 189 475
rect 208 474 210 488
rect 215 487 216 491
rect 220 490 221 491
rect 248 490 250 504
rect 950 503 951 507
rect 955 506 956 507
rect 1080 506 1082 516
rect 1087 515 1088 516
rect 1092 515 1093 519
rect 1137 518 1139 536
rect 1143 535 1149 536
rect 1143 531 1144 535
rect 1148 534 1149 535
rect 1159 534 1161 536
rect 1148 532 1161 534
rect 1148 531 1149 532
rect 1143 530 1149 531
rect 1182 530 1188 531
rect 1182 526 1183 530
rect 1187 526 1188 530
rect 1182 525 1188 526
rect 1143 519 1149 520
rect 1143 518 1144 519
rect 1137 516 1144 518
rect 1087 514 1093 515
rect 1143 515 1144 516
rect 1148 515 1149 519
rect 1192 518 1194 536
rect 1198 535 1205 536
rect 1198 531 1199 535
rect 1204 531 1205 535
rect 1246 535 1253 536
rect 1246 531 1247 535
rect 1252 531 1253 535
rect 1255 535 1256 539
rect 1260 538 1261 539
rect 1303 539 1309 540
rect 1260 536 1299 538
rect 1260 535 1261 536
rect 1255 534 1261 535
rect 1295 535 1301 536
rect 1295 531 1296 535
rect 1300 531 1301 535
rect 1303 535 1304 539
rect 1308 538 1309 539
rect 1359 539 1365 540
rect 1308 536 1355 538
rect 1308 535 1309 536
rect 1303 534 1309 535
rect 1351 535 1357 536
rect 1351 531 1352 535
rect 1356 531 1357 535
rect 1359 535 1360 539
rect 1364 538 1365 539
rect 1415 539 1421 540
rect 1364 536 1411 538
rect 1364 535 1365 536
rect 1359 534 1365 535
rect 1407 535 1413 536
rect 1407 531 1408 535
rect 1412 531 1413 535
rect 1415 535 1416 539
rect 1420 538 1421 539
rect 1471 539 1477 540
rect 1420 536 1467 538
rect 1420 535 1421 536
rect 1415 534 1421 535
rect 1463 535 1469 536
rect 1463 531 1464 535
rect 1468 531 1469 535
rect 1471 535 1472 539
rect 1476 538 1477 539
rect 1476 536 1522 538
rect 1616 536 1634 538
rect 1476 535 1477 536
rect 1471 534 1477 535
rect 1520 534 1522 536
rect 1527 535 1533 536
rect 1527 534 1528 535
rect 1520 532 1528 534
rect 1527 531 1528 532
rect 1532 531 1533 535
rect 1591 535 1597 536
rect 1591 531 1592 535
rect 1596 534 1597 535
rect 1616 534 1618 536
rect 1596 532 1618 534
rect 1596 531 1597 532
rect 1198 530 1205 531
rect 1230 530 1236 531
rect 1246 530 1253 531
rect 1278 530 1284 531
rect 1295 530 1301 531
rect 1334 530 1340 531
rect 1351 530 1357 531
rect 1390 530 1396 531
rect 1407 530 1413 531
rect 1446 530 1452 531
rect 1463 530 1469 531
rect 1510 530 1516 531
rect 1527 530 1533 531
rect 1574 530 1580 531
rect 1591 530 1597 531
rect 1622 530 1628 531
rect 1230 526 1231 530
rect 1235 526 1236 530
rect 1230 525 1236 526
rect 1278 526 1279 530
rect 1283 526 1284 530
rect 1278 525 1284 526
rect 1334 526 1335 530
rect 1339 526 1340 530
rect 1334 525 1340 526
rect 1390 526 1391 530
rect 1395 526 1396 530
rect 1390 525 1396 526
rect 1446 526 1447 530
rect 1451 526 1452 530
rect 1446 525 1452 526
rect 1510 526 1511 530
rect 1515 526 1516 530
rect 1510 525 1516 526
rect 1574 526 1575 530
rect 1579 526 1580 530
rect 1574 525 1580 526
rect 1622 526 1623 530
rect 1627 526 1628 530
rect 1622 525 1628 526
rect 1632 522 1634 536
rect 1639 535 1645 536
rect 1639 531 1640 535
rect 1644 534 1645 535
rect 1647 535 1653 536
rect 1647 534 1648 535
rect 1644 532 1648 534
rect 1644 531 1645 532
rect 1639 530 1645 531
rect 1647 531 1648 532
rect 1652 531 1653 535
rect 1647 530 1653 531
rect 1662 532 1668 533
rect 1662 528 1663 532
rect 1667 528 1668 532
rect 1662 527 1668 528
rect 1632 520 1643 522
rect 1199 519 1205 520
rect 1199 518 1200 519
rect 1192 516 1200 518
rect 1143 514 1149 515
rect 1199 515 1200 516
rect 1204 515 1205 519
rect 1199 514 1205 515
rect 1247 519 1253 520
rect 1247 515 1248 519
rect 1252 518 1253 519
rect 1255 519 1261 520
rect 1255 518 1256 519
rect 1252 516 1256 518
rect 1252 515 1253 516
rect 1247 514 1253 515
rect 1255 515 1256 516
rect 1260 515 1261 519
rect 1255 514 1261 515
rect 1295 519 1301 520
rect 1295 515 1296 519
rect 1300 518 1301 519
rect 1303 519 1309 520
rect 1303 518 1304 519
rect 1300 516 1304 518
rect 1300 515 1301 516
rect 1295 514 1301 515
rect 1303 515 1304 516
rect 1308 515 1309 519
rect 1303 514 1309 515
rect 1351 519 1357 520
rect 1351 515 1352 519
rect 1356 518 1357 519
rect 1359 519 1365 520
rect 1359 518 1360 519
rect 1356 516 1360 518
rect 1356 515 1357 516
rect 1351 514 1357 515
rect 1359 515 1360 516
rect 1364 515 1365 519
rect 1359 514 1365 515
rect 1407 519 1413 520
rect 1407 515 1408 519
rect 1412 518 1413 519
rect 1415 519 1421 520
rect 1415 518 1416 519
rect 1412 516 1416 518
rect 1412 515 1413 516
rect 1407 514 1413 515
rect 1415 515 1416 516
rect 1420 515 1421 519
rect 1415 514 1421 515
rect 1463 519 1469 520
rect 1463 515 1464 519
rect 1468 518 1469 519
rect 1471 519 1477 520
rect 1471 518 1472 519
rect 1468 516 1472 518
rect 1468 515 1469 516
rect 1463 514 1469 515
rect 1471 515 1472 516
rect 1476 515 1477 519
rect 1471 514 1477 515
rect 1526 519 1533 520
rect 1526 515 1527 519
rect 1532 515 1533 519
rect 1526 514 1533 515
rect 1591 519 1597 520
rect 1591 515 1592 519
rect 1596 518 1597 519
rect 1606 519 1612 520
rect 1606 518 1607 519
rect 1596 516 1607 518
rect 1596 515 1597 516
rect 1591 514 1597 515
rect 1606 515 1607 516
rect 1611 515 1612 519
rect 1606 514 1612 515
rect 1639 519 1645 520
rect 1639 515 1640 519
rect 1644 515 1645 519
rect 1639 514 1645 515
rect 1662 515 1668 516
rect 1126 513 1132 514
rect 1126 509 1127 513
rect 1131 509 1132 513
rect 1126 508 1132 509
rect 1182 513 1188 514
rect 1182 509 1183 513
rect 1187 509 1188 513
rect 1182 508 1188 509
rect 1230 513 1236 514
rect 1230 509 1231 513
rect 1235 509 1236 513
rect 1230 508 1236 509
rect 1278 513 1284 514
rect 1278 509 1279 513
rect 1283 509 1284 513
rect 1278 508 1284 509
rect 1334 513 1340 514
rect 1334 509 1335 513
rect 1339 509 1340 513
rect 1334 508 1340 509
rect 1390 513 1396 514
rect 1390 509 1391 513
rect 1395 509 1396 513
rect 1390 508 1396 509
rect 1446 513 1452 514
rect 1446 509 1447 513
rect 1451 509 1452 513
rect 1446 508 1452 509
rect 1510 513 1516 514
rect 1510 509 1511 513
rect 1515 509 1516 513
rect 1510 508 1516 509
rect 1574 513 1580 514
rect 1574 509 1575 513
rect 1579 509 1580 513
rect 1574 508 1580 509
rect 1622 513 1628 514
rect 1622 509 1623 513
rect 1627 509 1628 513
rect 1662 511 1663 515
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1622 508 1628 509
rect 955 504 1082 506
rect 1246 507 1252 508
rect 955 503 956 504
rect 950 502 956 503
rect 1246 503 1247 507
rect 1251 506 1252 507
rect 1251 504 1402 506
rect 1251 503 1252 504
rect 1246 502 1252 503
rect 286 499 292 500
rect 286 495 287 499
rect 291 495 292 499
rect 286 494 292 495
rect 326 499 332 500
rect 326 495 327 499
rect 331 495 332 499
rect 326 494 332 495
rect 374 499 380 500
rect 374 495 375 499
rect 379 495 380 499
rect 374 494 380 495
rect 422 499 428 500
rect 422 495 423 499
rect 427 495 428 499
rect 422 494 428 495
rect 478 499 484 500
rect 478 495 479 499
rect 483 495 484 499
rect 478 494 484 495
rect 542 499 548 500
rect 542 495 543 499
rect 547 495 548 499
rect 542 494 548 495
rect 614 499 620 500
rect 614 495 615 499
rect 619 495 620 499
rect 614 494 620 495
rect 694 499 700 500
rect 694 495 695 499
rect 699 495 700 499
rect 694 494 700 495
rect 774 499 780 500
rect 774 495 775 499
rect 779 495 780 499
rect 774 494 780 495
rect 846 499 852 500
rect 846 495 847 499
rect 851 495 852 499
rect 846 494 852 495
rect 918 499 924 500
rect 918 495 919 499
rect 923 495 924 499
rect 918 494 924 495
rect 982 499 988 500
rect 982 495 983 499
rect 987 495 988 499
rect 982 494 988 495
rect 1038 499 1044 500
rect 1038 495 1039 499
rect 1043 495 1044 499
rect 1038 494 1044 495
rect 1094 499 1100 500
rect 1094 495 1095 499
rect 1099 495 1100 499
rect 1094 494 1100 495
rect 1142 499 1148 500
rect 1142 495 1143 499
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1190 499 1196 500
rect 1190 495 1191 499
rect 1195 495 1196 499
rect 1190 494 1196 495
rect 1238 499 1244 500
rect 1238 495 1239 499
rect 1243 495 1244 499
rect 1238 494 1244 495
rect 1286 499 1292 500
rect 1286 495 1287 499
rect 1291 495 1292 499
rect 1286 494 1292 495
rect 1334 499 1340 500
rect 1334 495 1335 499
rect 1339 495 1340 499
rect 1334 494 1340 495
rect 1382 499 1388 500
rect 1382 495 1383 499
rect 1387 495 1388 499
rect 1382 494 1388 495
rect 1400 494 1402 504
rect 1430 499 1436 500
rect 1430 495 1431 499
rect 1435 495 1436 499
rect 1430 494 1436 495
rect 1478 499 1484 500
rect 1478 495 1479 499
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1534 499 1540 500
rect 1534 495 1535 499
rect 1539 495 1540 499
rect 1534 494 1540 495
rect 1590 499 1596 500
rect 1590 495 1591 499
rect 1595 495 1596 499
rect 1590 494 1596 495
rect 1622 499 1628 500
rect 1622 495 1623 499
rect 1627 495 1628 499
rect 1622 494 1628 495
rect 1662 497 1668 498
rect 1399 493 1405 494
rect 255 491 261 492
rect 255 490 256 491
rect 220 488 234 490
rect 248 488 256 490
rect 220 487 221 488
rect 215 486 221 487
rect 215 475 221 476
rect 215 474 216 475
rect 208 472 216 474
rect 183 470 189 471
rect 215 471 216 472
rect 220 471 221 475
rect 232 474 234 488
rect 255 487 256 488
rect 260 487 261 491
rect 255 486 261 487
rect 263 491 269 492
rect 263 487 264 491
rect 268 490 269 491
rect 303 491 309 492
rect 303 490 304 491
rect 268 488 304 490
rect 268 487 269 488
rect 263 486 269 487
rect 303 487 304 488
rect 308 487 309 491
rect 303 486 309 487
rect 343 491 349 492
rect 343 487 344 491
rect 348 490 349 491
rect 359 491 365 492
rect 359 490 360 491
rect 348 488 360 490
rect 348 487 349 488
rect 343 486 349 487
rect 359 487 360 488
rect 364 487 365 491
rect 391 491 397 492
rect 391 490 392 491
rect 359 486 365 487
rect 369 488 392 490
rect 238 482 244 483
rect 238 478 239 482
rect 243 478 244 482
rect 238 477 244 478
rect 286 482 292 483
rect 286 478 287 482
rect 291 478 292 482
rect 286 477 292 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 255 475 261 476
rect 255 474 256 475
rect 232 472 256 474
rect 215 470 221 471
rect 255 471 256 472
rect 260 471 261 475
rect 255 470 261 471
rect 274 475 280 476
rect 274 471 275 475
rect 279 474 280 475
rect 303 475 309 476
rect 303 474 304 475
rect 279 472 304 474
rect 279 471 280 472
rect 274 470 280 471
rect 303 471 304 472
rect 308 471 309 475
rect 303 470 309 471
rect 343 475 349 476
rect 343 471 344 475
rect 348 474 349 475
rect 369 474 371 488
rect 391 487 392 488
rect 396 487 397 491
rect 439 491 445 492
rect 439 490 440 491
rect 391 486 397 487
rect 416 488 440 490
rect 374 482 380 483
rect 374 478 375 482
rect 379 478 380 482
rect 374 477 380 478
rect 348 472 371 474
rect 391 475 397 476
rect 348 471 349 472
rect 343 470 349 471
rect 391 471 392 475
rect 396 474 397 475
rect 416 474 418 488
rect 439 487 440 488
rect 444 487 445 491
rect 495 491 501 492
rect 495 490 496 491
rect 439 486 445 487
rect 472 488 496 490
rect 422 482 428 483
rect 422 478 423 482
rect 427 478 428 482
rect 422 477 428 478
rect 396 472 418 474
rect 439 475 445 476
rect 396 471 397 472
rect 391 470 397 471
rect 439 471 440 475
rect 444 474 445 475
rect 472 474 474 488
rect 495 487 496 488
rect 500 487 501 491
rect 495 486 501 487
rect 559 491 565 492
rect 559 487 560 491
rect 564 490 565 491
rect 630 491 637 492
rect 564 488 598 490
rect 564 487 565 488
rect 559 486 565 487
rect 478 482 484 483
rect 478 478 479 482
rect 483 478 484 482
rect 478 477 484 478
rect 542 482 548 483
rect 542 478 543 482
rect 547 478 548 482
rect 542 477 548 478
rect 444 472 474 474
rect 486 475 492 476
rect 444 471 445 472
rect 439 470 445 471
rect 486 471 487 475
rect 491 474 492 475
rect 495 475 501 476
rect 495 474 496 475
rect 491 472 496 474
rect 491 471 492 472
rect 486 470 492 471
rect 495 471 496 472
rect 500 471 501 475
rect 495 470 501 471
rect 559 475 565 476
rect 559 471 560 475
rect 564 474 565 475
rect 596 474 598 488
rect 630 487 631 491
rect 636 487 637 491
rect 630 486 637 487
rect 639 491 645 492
rect 639 487 640 491
rect 644 490 645 491
rect 711 491 717 492
rect 711 490 712 491
rect 644 488 712 490
rect 644 487 645 488
rect 639 486 645 487
rect 711 487 712 488
rect 716 487 717 491
rect 711 486 717 487
rect 791 491 797 492
rect 791 487 792 491
rect 796 490 797 491
rect 834 491 840 492
rect 796 488 830 490
rect 796 487 797 488
rect 791 486 797 487
rect 614 482 620 483
rect 614 478 615 482
rect 619 478 620 482
rect 614 477 620 478
rect 694 482 700 483
rect 694 478 695 482
rect 699 478 700 482
rect 694 477 700 478
rect 774 482 780 483
rect 774 478 775 482
rect 779 478 780 482
rect 774 477 780 478
rect 631 475 637 476
rect 631 474 632 475
rect 564 472 594 474
rect 596 472 632 474
rect 564 471 565 472
rect 559 470 565 471
rect 153 466 155 470
rect 263 467 269 468
rect 263 466 264 467
rect 153 464 264 466
rect 263 463 264 464
rect 268 463 269 467
rect 592 466 594 472
rect 631 471 632 472
rect 636 471 637 475
rect 631 470 637 471
rect 702 475 708 476
rect 702 471 703 475
rect 707 474 708 475
rect 711 475 717 476
rect 711 474 712 475
rect 707 472 712 474
rect 707 471 708 472
rect 702 470 708 471
rect 711 471 712 472
rect 716 471 717 475
rect 711 470 717 471
rect 790 475 797 476
rect 790 471 791 475
rect 796 471 797 475
rect 828 474 830 488
rect 834 487 835 491
rect 839 490 840 491
rect 863 491 869 492
rect 863 490 864 491
rect 839 488 864 490
rect 839 487 840 488
rect 834 486 840 487
rect 863 487 864 488
rect 868 487 869 491
rect 863 486 869 487
rect 935 491 941 492
rect 935 487 936 491
rect 940 490 941 491
rect 999 491 1005 492
rect 940 488 970 490
rect 940 487 941 488
rect 935 486 941 487
rect 846 482 852 483
rect 846 478 847 482
rect 851 478 852 482
rect 846 477 852 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 863 475 869 476
rect 863 474 864 475
rect 828 472 864 474
rect 790 470 797 471
rect 863 471 864 472
rect 868 471 869 475
rect 863 470 869 471
rect 935 475 941 476
rect 935 471 936 475
rect 940 474 941 475
rect 950 475 956 476
rect 950 474 951 475
rect 940 472 951 474
rect 940 471 941 472
rect 935 470 941 471
rect 950 471 951 472
rect 955 471 956 475
rect 968 474 970 488
rect 999 487 1000 491
rect 1004 490 1005 491
rect 1055 491 1061 492
rect 1004 488 1030 490
rect 1004 487 1005 488
rect 999 486 1005 487
rect 982 482 988 483
rect 982 478 983 482
rect 987 478 988 482
rect 982 477 988 478
rect 999 475 1005 476
rect 999 474 1000 475
rect 968 472 1000 474
rect 950 470 956 471
rect 999 471 1000 472
rect 1004 471 1005 475
rect 1028 474 1030 488
rect 1055 487 1056 491
rect 1060 490 1061 491
rect 1111 491 1117 492
rect 1060 488 1086 490
rect 1060 487 1061 488
rect 1055 486 1061 487
rect 1038 482 1044 483
rect 1038 478 1039 482
rect 1043 478 1044 482
rect 1038 477 1044 478
rect 1055 475 1061 476
rect 1055 474 1056 475
rect 1028 472 1056 474
rect 999 470 1005 471
rect 1055 471 1056 472
rect 1060 471 1061 475
rect 1084 474 1086 488
rect 1111 487 1112 491
rect 1116 490 1117 491
rect 1159 491 1165 492
rect 1116 488 1139 490
rect 1116 487 1117 488
rect 1111 486 1117 487
rect 1094 482 1100 483
rect 1094 478 1095 482
rect 1099 478 1100 482
rect 1094 477 1100 478
rect 1111 475 1117 476
rect 1111 474 1112 475
rect 1084 472 1112 474
rect 1055 470 1061 471
rect 1111 471 1112 472
rect 1116 471 1117 475
rect 1137 474 1139 488
rect 1159 487 1160 491
rect 1164 490 1165 491
rect 1207 491 1213 492
rect 1164 488 1186 490
rect 1164 487 1165 488
rect 1159 486 1165 487
rect 1142 482 1148 483
rect 1142 478 1143 482
rect 1147 478 1148 482
rect 1142 477 1148 478
rect 1159 475 1165 476
rect 1159 474 1160 475
rect 1137 472 1160 474
rect 1111 470 1117 471
rect 1159 471 1160 472
rect 1164 471 1165 475
rect 1184 474 1186 488
rect 1207 487 1208 491
rect 1212 490 1213 491
rect 1255 491 1261 492
rect 1212 488 1235 490
rect 1212 487 1213 488
rect 1207 486 1213 487
rect 1190 482 1196 483
rect 1190 478 1191 482
rect 1195 478 1196 482
rect 1190 477 1196 478
rect 1207 475 1213 476
rect 1207 474 1208 475
rect 1184 472 1208 474
rect 1159 470 1165 471
rect 1207 471 1208 472
rect 1212 471 1213 475
rect 1233 474 1235 488
rect 1255 487 1256 491
rect 1260 490 1261 491
rect 1303 491 1309 492
rect 1260 488 1283 490
rect 1260 487 1261 488
rect 1255 486 1261 487
rect 1238 482 1244 483
rect 1238 478 1239 482
rect 1243 478 1244 482
rect 1238 477 1244 478
rect 1255 475 1261 476
rect 1255 474 1256 475
rect 1233 472 1256 474
rect 1207 470 1213 471
rect 1255 471 1256 472
rect 1260 471 1261 475
rect 1281 474 1283 488
rect 1303 487 1304 491
rect 1308 490 1309 491
rect 1351 491 1357 492
rect 1308 488 1330 490
rect 1308 487 1309 488
rect 1303 486 1309 487
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1286 477 1292 478
rect 1303 475 1309 476
rect 1303 474 1304 475
rect 1281 472 1304 474
rect 1255 470 1261 471
rect 1303 471 1304 472
rect 1308 471 1309 475
rect 1328 474 1330 488
rect 1351 487 1352 491
rect 1356 490 1357 491
rect 1356 488 1394 490
rect 1399 489 1400 493
rect 1404 489 1405 493
rect 1662 493 1663 497
rect 1667 493 1668 497
rect 1662 492 1668 493
rect 1399 488 1405 489
rect 1447 491 1453 492
rect 1356 487 1357 488
rect 1351 486 1357 487
rect 1334 482 1340 483
rect 1334 478 1335 482
rect 1339 478 1340 482
rect 1334 477 1340 478
rect 1382 482 1388 483
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1382 477 1388 478
rect 1351 475 1357 476
rect 1351 474 1352 475
rect 1328 472 1352 474
rect 1303 470 1309 471
rect 1351 471 1352 472
rect 1356 471 1357 475
rect 1392 474 1394 488
rect 1447 487 1448 491
rect 1452 490 1453 491
rect 1495 491 1501 492
rect 1452 488 1474 490
rect 1452 487 1453 488
rect 1447 486 1453 487
rect 1430 482 1436 483
rect 1430 478 1431 482
rect 1435 478 1436 482
rect 1430 477 1436 478
rect 1399 475 1405 476
rect 1399 474 1400 475
rect 1392 472 1400 474
rect 1351 470 1357 471
rect 1399 471 1400 472
rect 1404 471 1405 475
rect 1399 470 1405 471
rect 1447 475 1453 476
rect 1447 471 1448 475
rect 1452 474 1453 475
rect 1472 474 1474 488
rect 1495 487 1496 491
rect 1500 490 1501 491
rect 1510 491 1516 492
rect 1510 490 1511 491
rect 1500 488 1511 490
rect 1500 487 1501 488
rect 1495 486 1501 487
rect 1510 487 1511 488
rect 1515 487 1516 491
rect 1510 486 1516 487
rect 1518 491 1524 492
rect 1518 487 1519 491
rect 1523 490 1524 491
rect 1551 491 1557 492
rect 1551 490 1552 491
rect 1523 488 1552 490
rect 1523 487 1524 488
rect 1518 486 1524 487
rect 1551 487 1552 488
rect 1556 487 1557 491
rect 1551 486 1557 487
rect 1607 491 1613 492
rect 1607 487 1608 491
rect 1612 490 1613 491
rect 1638 491 1645 492
rect 1612 488 1634 490
rect 1612 487 1613 488
rect 1607 486 1613 487
rect 1478 482 1484 483
rect 1478 478 1479 482
rect 1483 478 1484 482
rect 1478 477 1484 478
rect 1534 482 1540 483
rect 1534 478 1535 482
rect 1539 478 1540 482
rect 1534 477 1540 478
rect 1590 482 1596 483
rect 1590 478 1591 482
rect 1595 478 1596 482
rect 1590 477 1596 478
rect 1622 482 1628 483
rect 1622 478 1623 482
rect 1627 478 1628 482
rect 1622 477 1628 478
rect 1495 475 1501 476
rect 1495 474 1496 475
rect 1452 472 1470 474
rect 1472 472 1496 474
rect 1452 471 1453 472
rect 1447 470 1453 471
rect 639 467 645 468
rect 639 466 640 467
rect 592 464 640 466
rect 263 462 269 463
rect 639 463 640 464
rect 644 463 645 467
rect 998 467 1004 468
rect 998 466 999 467
rect 639 462 645 463
rect 857 464 999 466
rect 231 459 237 460
rect 200 456 227 458
rect 167 455 173 456
rect 110 452 116 453
rect 110 448 111 452
rect 115 448 116 452
rect 167 451 168 455
rect 172 454 173 455
rect 190 455 196 456
rect 190 454 191 455
rect 172 452 191 454
rect 172 451 173 452
rect 110 447 116 448
rect 150 450 156 451
rect 167 450 173 451
rect 190 451 191 452
rect 195 451 196 455
rect 190 450 196 451
rect 150 446 151 450
rect 155 446 156 450
rect 150 445 156 446
rect 167 439 173 440
rect 110 435 116 436
rect 110 431 111 435
rect 115 431 116 435
rect 167 435 168 439
rect 172 438 173 439
rect 200 438 202 456
rect 223 455 229 456
rect 223 451 224 455
rect 228 451 229 455
rect 231 455 232 459
rect 236 458 237 459
rect 359 459 365 460
rect 236 456 266 458
rect 236 455 237 456
rect 231 454 237 455
rect 264 454 266 456
rect 271 455 277 456
rect 271 454 272 455
rect 264 452 272 454
rect 271 451 272 452
rect 276 451 277 455
rect 327 455 333 456
rect 327 451 328 455
rect 332 454 333 455
rect 351 455 357 456
rect 351 454 352 455
rect 332 452 352 454
rect 332 451 333 452
rect 206 450 212 451
rect 223 450 229 451
rect 254 450 260 451
rect 271 450 277 451
rect 310 450 316 451
rect 327 450 333 451
rect 351 451 352 452
rect 356 451 357 455
rect 359 455 360 459
rect 364 458 365 459
rect 391 459 397 460
rect 364 456 387 458
rect 364 455 365 456
rect 359 454 365 455
rect 383 455 389 456
rect 383 451 384 455
rect 388 451 389 455
rect 391 455 392 459
rect 396 458 397 459
rect 511 459 517 460
rect 396 456 459 458
rect 396 455 397 456
rect 391 454 397 455
rect 455 455 461 456
rect 455 451 456 455
rect 460 451 461 455
rect 511 455 512 459
rect 516 458 517 459
rect 543 459 549 460
rect 516 456 539 458
rect 516 455 517 456
rect 511 454 517 455
rect 535 455 541 456
rect 535 451 536 455
rect 540 451 541 455
rect 543 455 544 459
rect 548 458 549 459
rect 623 459 629 460
rect 548 456 619 458
rect 548 455 549 456
rect 543 454 549 455
rect 615 455 621 456
rect 615 451 616 455
rect 620 451 621 455
rect 623 455 624 459
rect 628 458 629 459
rect 628 456 690 458
rect 857 456 859 464
rect 998 463 999 464
rect 1003 463 1004 467
rect 1390 467 1396 468
rect 1390 466 1391 467
rect 998 462 1004 463
rect 1281 464 1391 466
rect 863 459 869 460
rect 628 455 629 456
rect 623 454 629 455
rect 688 454 690 456
rect 695 455 701 456
rect 695 454 696 455
rect 688 452 696 454
rect 695 451 696 452
rect 700 451 701 455
rect 775 455 781 456
rect 775 451 776 455
rect 780 454 781 455
rect 830 455 836 456
rect 830 454 831 455
rect 780 452 831 454
rect 780 451 781 452
rect 351 450 357 451
rect 366 450 372 451
rect 383 450 389 451
rect 438 450 444 451
rect 455 450 461 451
rect 518 450 524 451
rect 535 450 541 451
rect 598 450 604 451
rect 615 450 621 451
rect 678 450 684 451
rect 695 450 701 451
rect 758 450 764 451
rect 775 450 781 451
rect 830 451 831 452
rect 835 451 836 455
rect 855 455 861 456
rect 855 451 856 455
rect 860 451 861 455
rect 863 455 864 459
rect 868 458 869 459
rect 868 456 922 458
rect 1120 456 1139 458
rect 1159 456 1211 458
rect 1281 456 1283 464
rect 1390 463 1391 464
rect 1395 463 1396 467
rect 1468 466 1470 472
rect 1495 471 1496 472
rect 1500 471 1501 475
rect 1495 470 1501 471
rect 1551 475 1557 476
rect 1551 471 1552 475
rect 1556 474 1557 475
rect 1606 475 1613 476
rect 1556 472 1602 474
rect 1556 471 1557 472
rect 1551 470 1557 471
rect 1518 467 1524 468
rect 1518 466 1519 467
rect 1468 464 1519 466
rect 1390 462 1396 463
rect 1518 463 1519 464
rect 1523 463 1524 467
rect 1600 466 1602 472
rect 1606 471 1607 475
rect 1612 471 1613 475
rect 1632 474 1634 488
rect 1638 487 1639 491
rect 1644 487 1645 491
rect 1638 486 1645 487
rect 1662 480 1668 481
rect 1662 476 1663 480
rect 1667 476 1668 480
rect 1639 475 1645 476
rect 1662 475 1668 476
rect 1639 474 1640 475
rect 1632 472 1640 474
rect 1606 470 1613 471
rect 1639 471 1640 472
rect 1644 471 1645 475
rect 1639 470 1645 471
rect 1638 467 1644 468
rect 1638 466 1639 467
rect 1600 464 1639 466
rect 1518 462 1524 463
rect 1638 463 1639 464
rect 1643 463 1644 467
rect 1638 462 1644 463
rect 1287 459 1293 460
rect 868 455 869 456
rect 863 454 869 455
rect 920 454 922 456
rect 927 455 933 456
rect 927 454 928 455
rect 920 452 928 454
rect 927 451 928 452
rect 932 451 933 455
rect 999 455 1005 456
rect 999 451 1000 455
rect 1004 454 1005 455
rect 1071 455 1077 456
rect 1004 452 1042 454
rect 1004 451 1005 452
rect 830 450 836 451
rect 838 450 844 451
rect 855 450 861 451
rect 910 450 916 451
rect 927 450 933 451
rect 982 450 988 451
rect 999 450 1005 451
rect 206 446 207 450
rect 211 446 212 450
rect 206 445 212 446
rect 254 446 255 450
rect 259 446 260 450
rect 254 445 260 446
rect 310 446 311 450
rect 315 446 316 450
rect 310 445 316 446
rect 366 446 367 450
rect 371 446 372 450
rect 366 445 372 446
rect 438 446 439 450
rect 443 446 444 450
rect 438 445 444 446
rect 518 446 519 450
rect 523 446 524 450
rect 518 445 524 446
rect 598 446 599 450
rect 603 446 604 450
rect 598 445 604 446
rect 678 446 679 450
rect 683 446 684 450
rect 678 445 684 446
rect 758 446 759 450
rect 763 446 764 450
rect 758 445 764 446
rect 838 446 839 450
rect 843 446 844 450
rect 838 445 844 446
rect 910 446 911 450
rect 915 446 916 450
rect 910 445 916 446
rect 982 446 983 450
rect 987 446 988 450
rect 982 445 988 446
rect 1040 442 1042 452
rect 1071 451 1072 455
rect 1076 454 1077 455
rect 1120 454 1122 456
rect 1076 452 1122 454
rect 1076 451 1077 452
rect 1054 450 1060 451
rect 1071 450 1077 451
rect 1126 450 1132 451
rect 1054 446 1055 450
rect 1059 446 1060 450
rect 1054 445 1060 446
rect 1126 446 1127 450
rect 1131 446 1132 450
rect 1126 445 1132 446
rect 1040 440 1054 442
rect 172 436 202 438
rect 223 439 229 440
rect 172 435 173 436
rect 167 434 173 435
rect 223 435 224 439
rect 228 438 229 439
rect 231 439 237 440
rect 231 438 232 439
rect 228 436 232 438
rect 228 435 229 436
rect 223 434 229 435
rect 231 435 232 436
rect 236 435 237 439
rect 231 434 237 435
rect 271 439 280 440
rect 271 435 272 439
rect 279 435 280 439
rect 271 434 280 435
rect 326 439 333 440
rect 326 435 327 439
rect 332 435 333 439
rect 326 434 333 435
rect 383 439 389 440
rect 383 435 384 439
rect 388 438 389 439
rect 391 439 397 440
rect 391 438 392 439
rect 388 436 392 438
rect 388 435 389 436
rect 383 434 389 435
rect 391 435 392 436
rect 396 435 397 439
rect 391 434 397 435
rect 455 439 461 440
rect 455 435 456 439
rect 460 435 461 439
rect 455 434 461 435
rect 535 439 541 440
rect 535 435 536 439
rect 540 438 541 439
rect 543 439 549 440
rect 543 438 544 439
rect 540 436 544 438
rect 540 435 541 436
rect 535 434 541 435
rect 543 435 544 436
rect 548 435 549 439
rect 543 434 549 435
rect 615 439 621 440
rect 615 435 616 439
rect 620 438 621 439
rect 623 439 629 440
rect 623 438 624 439
rect 620 436 624 438
rect 620 435 621 436
rect 615 434 621 435
rect 623 435 624 436
rect 628 435 629 439
rect 623 434 629 435
rect 695 439 701 440
rect 695 435 696 439
rect 700 435 701 439
rect 695 434 701 435
rect 775 439 781 440
rect 775 435 776 439
rect 780 438 781 439
rect 822 439 828 440
rect 822 438 823 439
rect 780 436 823 438
rect 780 435 781 436
rect 775 434 781 435
rect 822 435 823 436
rect 827 435 828 439
rect 822 434 828 435
rect 855 439 861 440
rect 855 435 856 439
rect 860 438 861 439
rect 863 439 869 440
rect 863 438 864 439
rect 860 436 864 438
rect 860 435 861 436
rect 855 434 861 435
rect 863 435 864 436
rect 868 435 869 439
rect 863 434 869 435
rect 927 439 933 440
rect 927 435 928 439
rect 932 438 933 439
rect 950 439 956 440
rect 950 438 951 439
rect 932 436 951 438
rect 932 435 933 436
rect 927 434 933 435
rect 950 435 951 436
rect 955 435 956 439
rect 950 434 956 435
rect 998 439 1005 440
rect 998 435 999 439
rect 1004 435 1005 439
rect 1052 438 1066 440
rect 1071 439 1077 440
rect 1071 438 1072 439
rect 1064 436 1072 438
rect 998 434 1005 435
rect 1071 435 1072 436
rect 1076 435 1077 439
rect 1137 438 1139 456
rect 1143 455 1149 456
rect 1143 451 1144 455
rect 1148 454 1149 455
rect 1159 454 1161 456
rect 1148 452 1161 454
rect 1148 451 1149 452
rect 1143 450 1149 451
rect 1198 450 1204 451
rect 1198 446 1199 450
rect 1203 446 1204 450
rect 1198 445 1204 446
rect 1143 439 1149 440
rect 1143 438 1144 439
rect 1137 436 1144 438
rect 1071 434 1077 435
rect 1143 435 1144 436
rect 1148 435 1149 439
rect 1209 438 1211 456
rect 1214 455 1221 456
rect 1214 451 1215 455
rect 1220 451 1221 455
rect 1279 455 1285 456
rect 1279 451 1280 455
rect 1284 451 1285 455
rect 1287 455 1288 459
rect 1292 458 1293 459
rect 1292 456 1330 458
rect 1480 456 1506 458
rect 1292 455 1293 456
rect 1287 454 1293 455
rect 1328 454 1330 456
rect 1335 455 1341 456
rect 1335 454 1336 455
rect 1328 452 1336 454
rect 1335 451 1336 452
rect 1340 451 1341 455
rect 1391 455 1397 456
rect 1391 451 1392 455
rect 1396 454 1397 455
rect 1447 455 1453 456
rect 1396 452 1426 454
rect 1396 451 1397 452
rect 1214 450 1221 451
rect 1262 450 1268 451
rect 1279 450 1285 451
rect 1318 450 1324 451
rect 1335 450 1341 451
rect 1374 450 1380 451
rect 1391 450 1397 451
rect 1262 446 1263 450
rect 1267 446 1268 450
rect 1262 445 1268 446
rect 1318 446 1319 450
rect 1323 446 1324 450
rect 1318 445 1324 446
rect 1374 446 1375 450
rect 1379 446 1380 450
rect 1374 445 1380 446
rect 1424 442 1426 452
rect 1447 451 1448 455
rect 1452 454 1453 455
rect 1480 454 1482 456
rect 1452 452 1482 454
rect 1452 451 1453 452
rect 1430 450 1436 451
rect 1447 450 1453 451
rect 1494 450 1500 451
rect 1430 446 1431 450
rect 1435 446 1436 450
rect 1430 445 1436 446
rect 1494 446 1495 450
rect 1499 446 1500 450
rect 1494 445 1500 446
rect 1424 440 1430 442
rect 1215 439 1221 440
rect 1215 438 1216 439
rect 1209 436 1216 438
rect 1143 434 1149 435
rect 1215 435 1216 436
rect 1220 435 1221 439
rect 1215 434 1221 435
rect 1279 439 1285 440
rect 1279 435 1280 439
rect 1284 438 1285 439
rect 1287 439 1293 440
rect 1287 438 1288 439
rect 1284 436 1288 438
rect 1284 435 1285 436
rect 1279 434 1285 435
rect 1287 435 1288 436
rect 1292 435 1293 439
rect 1287 434 1293 435
rect 1335 439 1341 440
rect 1335 435 1336 439
rect 1340 438 1341 439
rect 1350 439 1356 440
rect 1350 438 1351 439
rect 1340 436 1351 438
rect 1340 435 1341 436
rect 1335 434 1341 435
rect 1350 435 1351 436
rect 1355 435 1356 439
rect 1350 434 1356 435
rect 1390 439 1397 440
rect 1390 435 1391 439
rect 1396 435 1397 439
rect 1428 438 1442 440
rect 1447 439 1453 440
rect 1447 438 1448 439
rect 1440 436 1448 438
rect 1390 434 1397 435
rect 1447 435 1448 436
rect 1452 435 1453 439
rect 1504 438 1506 456
rect 1510 455 1517 456
rect 1510 451 1511 455
rect 1516 451 1517 455
rect 1510 450 1517 451
rect 1662 452 1668 453
rect 1662 448 1663 452
rect 1667 448 1668 452
rect 1662 447 1668 448
rect 1511 439 1517 440
rect 1511 438 1512 439
rect 1504 436 1512 438
rect 1447 434 1453 435
rect 1511 435 1512 436
rect 1516 435 1517 439
rect 1511 434 1517 435
rect 1662 435 1668 436
rect 110 430 116 431
rect 150 433 156 434
rect 150 429 151 433
rect 155 429 156 433
rect 150 428 156 429
rect 206 433 212 434
rect 206 429 207 433
rect 211 429 212 433
rect 206 428 212 429
rect 254 433 260 434
rect 254 429 255 433
rect 259 429 260 433
rect 254 428 260 429
rect 310 433 316 434
rect 310 429 311 433
rect 315 429 316 433
rect 310 428 316 429
rect 366 433 372 434
rect 366 429 367 433
rect 371 429 372 433
rect 366 428 372 429
rect 438 433 444 434
rect 438 429 439 433
rect 443 429 444 433
rect 438 428 444 429
rect 351 427 357 428
rect 351 423 352 427
rect 356 426 357 427
rect 457 426 459 434
rect 518 433 524 434
rect 518 429 519 433
rect 523 429 524 433
rect 518 428 524 429
rect 598 433 604 434
rect 598 429 599 433
rect 603 429 604 433
rect 598 428 604 429
rect 678 433 684 434
rect 678 429 679 433
rect 683 429 684 433
rect 678 428 684 429
rect 758 433 764 434
rect 758 429 759 433
rect 763 429 764 433
rect 758 428 764 429
rect 838 433 844 434
rect 838 429 839 433
rect 843 429 844 433
rect 838 428 844 429
rect 910 433 916 434
rect 910 429 911 433
rect 915 429 916 433
rect 910 428 916 429
rect 982 433 988 434
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 1054 433 1060 434
rect 1054 429 1055 433
rect 1059 429 1060 433
rect 1054 428 1060 429
rect 1126 433 1132 434
rect 1126 429 1127 433
rect 1131 429 1132 433
rect 1126 428 1132 429
rect 1198 433 1204 434
rect 1198 429 1199 433
rect 1203 429 1204 433
rect 1198 428 1204 429
rect 1262 433 1268 434
rect 1262 429 1263 433
rect 1267 429 1268 433
rect 1262 428 1268 429
rect 1318 433 1324 434
rect 1318 429 1319 433
rect 1323 429 1324 433
rect 1318 428 1324 429
rect 1374 433 1380 434
rect 1374 429 1375 433
rect 1379 429 1380 433
rect 1374 428 1380 429
rect 1430 433 1436 434
rect 1430 429 1431 433
rect 1435 429 1436 433
rect 1430 428 1436 429
rect 1494 433 1500 434
rect 1494 429 1495 433
rect 1499 429 1500 433
rect 1662 431 1663 435
rect 1667 431 1668 435
rect 1662 430 1668 431
rect 1494 428 1500 429
rect 1214 427 1220 428
rect 1214 426 1215 427
rect 356 424 459 426
rect 1159 424 1215 426
rect 356 423 357 424
rect 351 422 357 423
rect 174 419 180 420
rect 110 417 116 418
rect 110 413 111 417
rect 115 413 116 417
rect 174 415 175 419
rect 179 415 180 419
rect 174 414 180 415
rect 222 419 228 420
rect 222 415 223 419
rect 227 415 228 419
rect 222 414 228 415
rect 270 419 276 420
rect 270 415 271 419
rect 275 415 276 419
rect 270 414 276 415
rect 318 419 324 420
rect 318 415 319 419
rect 323 415 324 419
rect 318 414 324 415
rect 366 419 372 420
rect 366 415 367 419
rect 371 415 372 419
rect 366 414 372 415
rect 414 419 420 420
rect 414 415 415 419
rect 419 415 420 419
rect 414 414 420 415
rect 470 419 476 420
rect 470 415 471 419
rect 475 415 476 419
rect 470 414 476 415
rect 526 419 532 420
rect 526 415 527 419
rect 531 415 532 419
rect 526 414 532 415
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 590 414 596 415
rect 662 419 668 420
rect 662 415 663 419
rect 667 415 668 419
rect 662 414 668 415
rect 734 419 740 420
rect 734 415 735 419
rect 739 415 740 419
rect 734 414 740 415
rect 806 419 812 420
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 870 419 876 420
rect 870 415 871 419
rect 875 415 876 419
rect 870 414 876 415
rect 934 419 940 420
rect 934 415 935 419
rect 939 415 940 419
rect 934 414 940 415
rect 990 419 996 420
rect 990 415 991 419
rect 995 415 996 419
rect 990 414 996 415
rect 1038 419 1044 420
rect 1038 415 1039 419
rect 1043 415 1044 419
rect 1038 414 1044 415
rect 1086 419 1092 420
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1126 419 1132 420
rect 1126 415 1127 419
rect 1131 415 1132 419
rect 1126 414 1132 415
rect 110 412 116 413
rect 190 411 197 412
rect 190 407 191 411
rect 196 407 197 411
rect 239 411 245 412
rect 239 410 240 411
rect 190 406 197 407
rect 216 408 240 410
rect 174 402 180 403
rect 110 400 116 401
rect 110 396 111 400
rect 115 396 116 400
rect 174 398 175 402
rect 179 398 180 402
rect 174 397 180 398
rect 110 395 116 396
rect 191 395 197 396
rect 191 391 192 395
rect 196 394 197 395
rect 216 394 218 408
rect 239 407 240 408
rect 244 407 245 411
rect 239 406 245 407
rect 287 411 293 412
rect 287 407 288 411
rect 292 410 293 411
rect 335 411 341 412
rect 292 408 330 410
rect 292 407 293 408
rect 287 406 293 407
rect 222 402 228 403
rect 222 398 223 402
rect 227 398 228 402
rect 222 397 228 398
rect 270 402 276 403
rect 270 398 271 402
rect 275 398 276 402
rect 270 397 276 398
rect 318 402 324 403
rect 318 398 319 402
rect 323 398 324 402
rect 328 402 330 408
rect 335 407 336 411
rect 340 410 341 411
rect 383 411 389 412
rect 340 408 362 410
rect 340 407 341 408
rect 335 406 341 407
rect 328 400 338 402
rect 318 397 324 398
rect 336 396 338 400
rect 196 392 218 394
rect 230 395 236 396
rect 196 391 197 392
rect 191 390 197 391
rect 230 391 231 395
rect 235 394 236 395
rect 239 395 245 396
rect 239 394 240 395
rect 235 392 240 394
rect 235 391 236 392
rect 230 390 236 391
rect 239 391 240 392
rect 244 391 245 395
rect 239 390 245 391
rect 287 395 293 396
rect 287 391 288 395
rect 292 394 293 395
rect 326 395 332 396
rect 326 394 327 395
rect 292 392 327 394
rect 292 391 293 392
rect 287 390 293 391
rect 326 391 327 392
rect 331 391 332 395
rect 326 390 332 391
rect 335 395 341 396
rect 335 391 336 395
rect 340 391 341 395
rect 360 394 362 408
rect 383 407 384 411
rect 388 410 389 411
rect 426 411 437 412
rect 388 408 411 410
rect 388 407 389 408
rect 383 406 389 407
rect 366 402 372 403
rect 366 398 367 402
rect 371 398 372 402
rect 366 397 372 398
rect 383 395 389 396
rect 383 394 384 395
rect 360 392 384 394
rect 335 390 341 391
rect 383 391 384 392
rect 388 391 389 395
rect 409 394 411 408
rect 426 407 427 411
rect 431 407 432 411
rect 436 407 437 411
rect 426 406 437 407
rect 487 411 493 412
rect 487 407 488 411
rect 492 410 493 411
rect 511 411 517 412
rect 511 410 512 411
rect 492 408 512 410
rect 492 407 493 408
rect 487 406 493 407
rect 511 407 512 408
rect 516 407 517 411
rect 543 411 549 412
rect 543 410 544 411
rect 511 406 517 407
rect 520 408 544 410
rect 414 402 420 403
rect 414 398 415 402
rect 419 398 420 402
rect 414 397 420 398
rect 470 402 476 403
rect 470 398 471 402
rect 475 398 476 402
rect 470 397 476 398
rect 431 395 437 396
rect 431 394 432 395
rect 409 392 432 394
rect 383 390 389 391
rect 431 391 432 392
rect 436 391 437 395
rect 431 390 437 391
rect 487 395 493 396
rect 487 391 488 395
rect 492 394 493 395
rect 520 394 522 408
rect 543 407 544 408
rect 548 407 549 411
rect 607 411 613 412
rect 607 410 608 411
rect 543 406 549 407
rect 580 408 608 410
rect 526 402 532 403
rect 526 398 527 402
rect 531 398 532 402
rect 526 397 532 398
rect 492 392 522 394
rect 543 395 549 396
rect 492 391 493 392
rect 487 390 493 391
rect 543 391 544 395
rect 548 394 549 395
rect 580 394 582 408
rect 607 407 608 408
rect 612 407 613 411
rect 679 411 685 412
rect 679 410 680 411
rect 607 406 613 407
rect 648 408 680 410
rect 590 402 596 403
rect 590 398 591 402
rect 595 398 596 402
rect 590 397 596 398
rect 548 392 582 394
rect 607 395 613 396
rect 548 391 549 392
rect 543 390 549 391
rect 607 391 608 395
rect 612 394 613 395
rect 648 394 650 408
rect 679 407 680 408
rect 684 407 685 411
rect 679 406 685 407
rect 751 411 760 412
rect 751 407 752 411
rect 759 407 760 411
rect 823 411 829 412
rect 823 410 824 411
rect 751 406 760 407
rect 788 408 824 410
rect 662 402 668 403
rect 662 398 663 402
rect 667 398 668 402
rect 662 397 668 398
rect 734 402 740 403
rect 734 398 735 402
rect 739 398 740 402
rect 734 397 740 398
rect 612 392 650 394
rect 670 395 676 396
rect 612 391 613 392
rect 607 390 613 391
rect 670 391 671 395
rect 675 394 676 395
rect 679 395 685 396
rect 679 394 680 395
rect 675 392 680 394
rect 675 391 676 392
rect 670 390 676 391
rect 679 391 680 392
rect 684 391 685 395
rect 679 390 685 391
rect 751 395 757 396
rect 751 391 752 395
rect 756 394 757 395
rect 788 394 790 408
rect 823 407 824 408
rect 828 407 829 411
rect 823 406 829 407
rect 882 411 893 412
rect 882 407 883 411
rect 887 407 888 411
rect 892 407 893 411
rect 882 406 893 407
rect 951 411 957 412
rect 951 407 952 411
rect 956 410 957 411
rect 1002 411 1013 412
rect 956 408 982 410
rect 956 407 957 408
rect 951 406 957 407
rect 806 402 812 403
rect 806 398 807 402
rect 811 398 812 402
rect 806 397 812 398
rect 870 402 876 403
rect 870 398 871 402
rect 875 398 876 402
rect 870 397 876 398
rect 934 402 940 403
rect 934 398 935 402
rect 939 398 940 402
rect 934 397 940 398
rect 756 392 790 394
rect 822 395 829 396
rect 756 391 757 392
rect 751 390 757 391
rect 822 391 823 395
rect 828 391 829 395
rect 822 390 829 391
rect 887 395 893 396
rect 887 391 888 395
rect 892 394 893 395
rect 950 395 957 396
rect 892 392 946 394
rect 892 391 893 392
rect 887 390 893 391
rect 944 386 946 392
rect 950 391 951 395
rect 956 391 957 395
rect 980 394 982 408
rect 1002 407 1003 411
rect 1007 407 1008 411
rect 1012 407 1013 411
rect 1002 406 1013 407
rect 1055 411 1061 412
rect 1055 407 1056 411
rect 1060 410 1061 411
rect 1103 411 1109 412
rect 1060 408 1082 410
rect 1060 407 1061 408
rect 1055 406 1061 407
rect 990 402 996 403
rect 990 398 991 402
rect 995 398 996 402
rect 990 397 996 398
rect 1038 402 1044 403
rect 1038 398 1039 402
rect 1043 398 1044 402
rect 1038 397 1044 398
rect 1007 395 1013 396
rect 1007 394 1008 395
rect 980 392 1008 394
rect 950 390 957 391
rect 1007 391 1008 392
rect 1012 391 1013 395
rect 1007 390 1013 391
rect 1055 395 1061 396
rect 1055 391 1056 395
rect 1060 394 1061 395
rect 1080 394 1082 408
rect 1103 407 1104 411
rect 1108 410 1109 411
rect 1143 411 1149 412
rect 1108 408 1122 410
rect 1108 407 1109 408
rect 1103 406 1109 407
rect 1086 402 1092 403
rect 1086 398 1087 402
rect 1091 398 1092 402
rect 1086 397 1092 398
rect 1103 395 1109 396
rect 1103 394 1104 395
rect 1060 392 1078 394
rect 1080 392 1104 394
rect 1060 391 1061 392
rect 1055 390 1061 391
rect 1002 387 1008 388
rect 1002 386 1003 387
rect 944 384 1003 386
rect 814 383 820 384
rect 814 382 815 383
rect 705 380 815 382
rect 487 375 493 376
rect 160 372 187 374
rect 288 372 306 374
rect 319 372 362 374
rect 369 372 418 374
rect 150 371 157 372
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 150 367 151 371
rect 156 367 157 371
rect 110 363 116 364
rect 134 366 140 367
rect 150 366 157 367
rect 134 362 135 366
rect 139 362 140 366
rect 134 361 140 362
rect 151 355 157 356
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 151 351 152 355
rect 156 354 157 355
rect 160 354 162 372
rect 183 371 189 372
rect 183 367 184 371
rect 188 367 189 371
rect 215 371 221 372
rect 215 370 216 371
rect 208 368 216 370
rect 166 366 172 367
rect 183 366 189 367
rect 198 366 204 367
rect 166 362 167 366
rect 171 362 172 366
rect 166 361 172 362
rect 198 362 199 366
rect 203 362 204 366
rect 198 361 204 362
rect 208 356 210 368
rect 215 367 216 368
rect 220 367 221 371
rect 255 371 261 372
rect 255 367 256 371
rect 260 370 261 371
rect 288 370 290 372
rect 260 368 290 370
rect 260 367 261 368
rect 215 366 221 367
rect 238 366 244 367
rect 255 366 261 367
rect 294 366 300 367
rect 238 362 239 366
rect 243 362 244 366
rect 238 361 244 362
rect 294 362 295 366
rect 299 362 300 366
rect 294 361 300 362
rect 156 352 162 354
rect 183 355 189 356
rect 156 351 157 352
rect 151 350 157 351
rect 183 351 184 355
rect 188 354 189 355
rect 196 354 210 356
rect 215 355 221 356
rect 188 352 198 354
rect 188 351 189 352
rect 183 350 189 351
rect 215 351 216 355
rect 220 354 221 355
rect 230 355 236 356
rect 230 354 231 355
rect 220 352 231 354
rect 220 351 221 352
rect 215 350 221 351
rect 230 351 231 352
rect 235 351 236 355
rect 230 350 236 351
rect 250 355 261 356
rect 250 351 251 355
rect 255 351 256 355
rect 260 351 261 355
rect 304 354 306 372
rect 311 371 317 372
rect 311 367 312 371
rect 316 370 317 371
rect 319 370 321 372
rect 316 368 321 370
rect 316 367 317 368
rect 311 366 317 367
rect 350 366 356 367
rect 350 362 351 366
rect 355 362 356 366
rect 350 361 356 362
rect 311 355 317 356
rect 311 354 312 355
rect 304 352 312 354
rect 250 350 261 351
rect 311 351 312 352
rect 316 351 317 355
rect 360 354 362 372
rect 367 371 373 372
rect 367 367 368 371
rect 372 367 373 371
rect 367 366 373 367
rect 406 366 412 367
rect 406 362 407 366
rect 411 362 412 366
rect 406 361 412 362
rect 367 355 373 356
rect 367 354 368 355
rect 360 352 368 354
rect 311 350 317 351
rect 367 351 368 352
rect 372 351 373 355
rect 416 354 418 372
rect 423 371 432 372
rect 423 367 424 371
rect 431 367 432 371
rect 474 371 485 372
rect 474 367 475 371
rect 479 367 480 371
rect 484 367 485 371
rect 487 371 488 375
rect 492 374 493 375
rect 543 375 549 376
rect 492 372 539 374
rect 492 371 493 372
rect 487 370 493 371
rect 535 371 541 372
rect 535 367 536 371
rect 540 367 541 371
rect 543 371 544 375
rect 548 374 549 375
rect 599 375 605 376
rect 548 372 595 374
rect 548 371 549 372
rect 543 370 549 371
rect 591 371 597 372
rect 591 367 592 371
rect 596 367 597 371
rect 599 371 600 375
rect 604 374 605 375
rect 604 372 651 374
rect 705 372 707 380
rect 814 379 815 380
rect 819 379 820 383
rect 1002 383 1003 384
rect 1007 383 1008 387
rect 1076 386 1078 392
rect 1103 391 1104 392
rect 1108 391 1109 395
rect 1120 394 1122 408
rect 1143 407 1144 411
rect 1148 410 1149 411
rect 1159 410 1161 424
rect 1214 423 1215 424
rect 1219 423 1220 427
rect 1214 422 1220 423
rect 1166 419 1172 420
rect 1166 415 1167 419
rect 1171 415 1172 419
rect 1166 414 1172 415
rect 1206 419 1212 420
rect 1206 415 1207 419
rect 1211 415 1212 419
rect 1206 414 1212 415
rect 1246 419 1252 420
rect 1246 415 1247 419
rect 1251 415 1252 419
rect 1246 414 1252 415
rect 1286 419 1292 420
rect 1286 415 1287 419
rect 1291 415 1292 419
rect 1286 414 1292 415
rect 1334 419 1340 420
rect 1334 415 1335 419
rect 1339 415 1340 419
rect 1334 414 1340 415
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1382 414 1388 415
rect 1662 417 1668 418
rect 1662 413 1663 417
rect 1667 413 1668 417
rect 1662 412 1668 413
rect 1148 408 1161 410
rect 1183 411 1189 412
rect 1148 407 1149 408
rect 1143 406 1149 407
rect 1183 407 1184 411
rect 1188 410 1189 411
rect 1191 411 1197 412
rect 1191 410 1192 411
rect 1188 408 1192 410
rect 1188 407 1189 408
rect 1183 406 1189 407
rect 1191 407 1192 408
rect 1196 407 1197 411
rect 1223 411 1229 412
rect 1223 410 1224 411
rect 1191 406 1197 407
rect 1200 408 1224 410
rect 1126 402 1132 403
rect 1126 398 1127 402
rect 1131 398 1132 402
rect 1126 397 1132 398
rect 1166 402 1172 403
rect 1166 398 1167 402
rect 1171 398 1172 402
rect 1166 397 1172 398
rect 1143 395 1149 396
rect 1143 394 1144 395
rect 1120 392 1144 394
rect 1103 390 1109 391
rect 1143 391 1144 392
rect 1148 391 1149 395
rect 1143 390 1149 391
rect 1183 395 1189 396
rect 1183 391 1184 395
rect 1188 394 1189 395
rect 1200 394 1202 408
rect 1223 407 1224 408
rect 1228 407 1229 411
rect 1263 411 1269 412
rect 1263 410 1264 411
rect 1223 406 1229 407
rect 1240 408 1264 410
rect 1206 402 1212 403
rect 1206 398 1207 402
rect 1211 398 1212 402
rect 1206 397 1212 398
rect 1188 392 1202 394
rect 1223 395 1229 396
rect 1188 391 1189 392
rect 1183 390 1189 391
rect 1223 391 1224 395
rect 1228 394 1229 395
rect 1240 394 1242 408
rect 1263 407 1264 408
rect 1268 407 1269 411
rect 1303 411 1309 412
rect 1303 410 1304 411
rect 1263 406 1269 407
rect 1281 408 1304 410
rect 1246 402 1252 403
rect 1246 398 1247 402
rect 1251 398 1252 402
rect 1246 397 1252 398
rect 1228 392 1242 394
rect 1263 395 1269 396
rect 1228 391 1229 392
rect 1223 390 1229 391
rect 1263 391 1264 395
rect 1268 394 1269 395
rect 1281 394 1283 408
rect 1303 407 1304 408
rect 1308 407 1309 411
rect 1303 406 1309 407
rect 1351 411 1357 412
rect 1351 407 1352 411
rect 1356 410 1357 411
rect 1399 411 1405 412
rect 1356 408 1394 410
rect 1356 407 1357 408
rect 1351 406 1357 407
rect 1286 402 1292 403
rect 1286 398 1287 402
rect 1291 398 1292 402
rect 1286 397 1292 398
rect 1334 402 1340 403
rect 1334 398 1335 402
rect 1339 398 1340 402
rect 1334 397 1340 398
rect 1382 402 1388 403
rect 1382 398 1383 402
rect 1387 398 1388 402
rect 1382 397 1388 398
rect 1268 392 1283 394
rect 1303 395 1309 396
rect 1268 391 1269 392
rect 1263 390 1269 391
rect 1303 391 1304 395
rect 1308 394 1309 395
rect 1350 395 1357 396
rect 1308 392 1347 394
rect 1308 391 1309 392
rect 1303 390 1309 391
rect 1110 387 1116 388
rect 1110 386 1111 387
rect 1076 384 1111 386
rect 1002 382 1008 383
rect 1110 383 1111 384
rect 1115 383 1116 387
rect 1345 386 1347 392
rect 1350 391 1351 395
rect 1356 391 1357 395
rect 1392 394 1394 408
rect 1399 407 1400 411
rect 1404 410 1405 411
rect 1407 411 1413 412
rect 1407 410 1408 411
rect 1404 408 1408 410
rect 1404 407 1405 408
rect 1399 406 1405 407
rect 1407 407 1408 408
rect 1412 407 1413 411
rect 1407 406 1413 407
rect 1662 400 1668 401
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1399 395 1405 396
rect 1662 395 1668 396
rect 1399 394 1400 395
rect 1392 392 1400 394
rect 1350 390 1357 391
rect 1399 391 1400 392
rect 1404 391 1405 395
rect 1399 390 1405 391
rect 1407 387 1413 388
rect 1407 386 1408 387
rect 1345 384 1408 386
rect 1110 382 1116 383
rect 1407 383 1408 384
rect 1412 383 1413 387
rect 1407 382 1413 383
rect 814 378 820 379
rect 767 375 773 376
rect 604 371 605 372
rect 599 370 605 371
rect 647 371 653 372
rect 647 367 648 371
rect 652 367 653 371
rect 703 371 709 372
rect 703 367 704 371
rect 708 367 709 371
rect 754 371 765 372
rect 754 367 755 371
rect 759 367 760 371
rect 764 367 765 371
rect 767 371 768 375
rect 772 374 773 375
rect 890 375 896 376
rect 772 372 810 374
rect 772 371 773 372
rect 767 370 773 371
rect 808 370 810 372
rect 815 371 821 372
rect 815 370 816 371
rect 808 368 816 370
rect 815 367 816 368
rect 820 367 821 371
rect 871 371 877 372
rect 871 367 872 371
rect 876 370 877 371
rect 882 371 888 372
rect 882 370 883 371
rect 876 368 883 370
rect 876 367 877 368
rect 423 366 432 367
rect 462 366 468 367
rect 474 366 485 367
rect 518 366 524 367
rect 535 366 541 367
rect 574 366 580 367
rect 591 366 597 367
rect 630 366 636 367
rect 647 366 653 367
rect 686 366 692 367
rect 703 366 709 367
rect 742 366 748 367
rect 754 366 765 367
rect 798 366 804 367
rect 815 366 821 367
rect 854 366 860 367
rect 871 366 877 367
rect 882 367 883 368
rect 887 367 888 371
rect 890 371 891 375
rect 895 374 896 375
rect 943 375 949 376
rect 895 372 930 374
rect 895 371 896 372
rect 890 370 896 371
rect 928 370 930 372
rect 935 371 941 372
rect 935 370 936 371
rect 928 368 936 370
rect 935 367 936 368
rect 940 367 941 371
rect 943 371 944 375
rect 948 374 949 375
rect 1007 375 1013 376
rect 948 372 994 374
rect 948 371 949 372
rect 943 370 949 371
rect 992 370 994 372
rect 999 371 1005 372
rect 999 370 1000 371
rect 992 368 1000 370
rect 999 367 1000 368
rect 1004 367 1005 371
rect 1007 371 1008 375
rect 1012 374 1013 375
rect 1191 375 1197 376
rect 1012 372 1050 374
rect 1012 371 1013 372
rect 1007 370 1013 371
rect 1048 370 1050 372
rect 1055 371 1061 372
rect 1055 370 1056 371
rect 1048 368 1056 370
rect 1055 367 1056 368
rect 1060 367 1061 371
rect 1111 371 1117 372
rect 1111 367 1112 371
rect 1116 367 1117 371
rect 1158 371 1164 372
rect 1158 367 1159 371
rect 1163 370 1164 371
rect 1167 371 1173 372
rect 1167 370 1168 371
rect 1163 368 1168 370
rect 1163 367 1164 368
rect 882 366 888 367
rect 918 366 924 367
rect 935 366 941 367
rect 982 366 988 367
rect 999 366 1005 367
rect 1038 366 1044 367
rect 1055 366 1061 367
rect 1094 366 1100 367
rect 1111 366 1117 367
rect 1150 366 1156 367
rect 1158 366 1164 367
rect 1167 367 1168 368
rect 1172 367 1173 371
rect 1191 371 1192 375
rect 1196 374 1197 375
rect 1238 375 1244 376
rect 1196 372 1218 374
rect 1196 371 1197 372
rect 1191 370 1197 371
rect 1216 370 1218 372
rect 1223 371 1229 372
rect 1223 370 1224 371
rect 1216 368 1224 370
rect 1223 367 1224 368
rect 1228 367 1229 371
rect 1238 371 1239 375
rect 1243 374 1244 375
rect 1279 375 1285 376
rect 1243 372 1266 374
rect 1243 371 1244 372
rect 1238 370 1244 371
rect 1264 370 1266 372
rect 1271 371 1277 372
rect 1271 370 1272 371
rect 1264 368 1272 370
rect 1271 367 1272 368
rect 1276 367 1277 371
rect 1279 371 1280 375
rect 1284 374 1285 375
rect 1327 375 1333 376
rect 1284 372 1314 374
rect 1284 371 1285 372
rect 1279 370 1285 371
rect 1312 370 1314 372
rect 1319 371 1325 372
rect 1319 370 1320 371
rect 1312 368 1320 370
rect 1319 367 1320 368
rect 1324 367 1325 371
rect 1327 371 1328 375
rect 1332 374 1333 375
rect 1375 375 1381 376
rect 1332 372 1371 374
rect 1332 371 1333 372
rect 1327 370 1333 371
rect 1367 371 1373 372
rect 1367 367 1368 371
rect 1372 367 1373 371
rect 1375 371 1376 375
rect 1380 374 1381 375
rect 1438 375 1444 376
rect 1380 372 1410 374
rect 1380 371 1381 372
rect 1375 370 1381 371
rect 1408 370 1410 372
rect 1415 371 1421 372
rect 1415 370 1416 371
rect 1408 368 1416 370
rect 1415 367 1416 368
rect 1420 367 1421 371
rect 1438 371 1439 375
rect 1443 374 1444 375
rect 1519 375 1525 376
rect 1443 372 1467 374
rect 1443 371 1444 372
rect 1438 370 1444 371
rect 1463 371 1469 372
rect 1463 367 1464 371
rect 1468 367 1469 371
rect 1511 371 1517 372
rect 1511 367 1512 371
rect 1516 367 1517 371
rect 1519 371 1520 375
rect 1524 374 1525 375
rect 1567 375 1573 376
rect 1524 372 1563 374
rect 1524 371 1525 372
rect 1519 370 1525 371
rect 1559 371 1565 372
rect 1167 366 1173 367
rect 1206 366 1212 367
rect 1223 366 1229 367
rect 1254 366 1260 367
rect 1271 366 1277 367
rect 1302 366 1308 367
rect 1319 366 1325 367
rect 1350 366 1356 367
rect 1367 366 1373 367
rect 1398 366 1404 367
rect 1415 366 1421 367
rect 1446 366 1452 367
rect 1463 366 1469 367
rect 1494 366 1500 367
rect 1511 366 1517 367
rect 1534 367 1540 368
rect 1559 367 1560 371
rect 1564 367 1565 371
rect 1567 371 1568 375
rect 1572 374 1573 375
rect 1572 372 1611 374
rect 1616 372 1643 374
rect 1572 371 1573 372
rect 1567 370 1573 371
rect 1607 371 1613 372
rect 1607 367 1608 371
rect 1612 367 1613 371
rect 1534 366 1535 367
rect 462 362 463 366
rect 467 362 468 366
rect 462 361 468 362
rect 518 362 519 366
rect 523 362 524 366
rect 518 361 524 362
rect 574 362 575 366
rect 579 362 580 366
rect 574 361 580 362
rect 630 362 631 366
rect 635 362 636 366
rect 630 361 636 362
rect 686 362 687 366
rect 691 362 692 366
rect 686 361 692 362
rect 742 362 743 366
rect 747 362 748 366
rect 742 361 748 362
rect 798 362 799 366
rect 803 362 804 366
rect 798 361 804 362
rect 854 362 855 366
rect 859 362 860 366
rect 854 361 860 362
rect 918 362 919 366
rect 923 362 924 366
rect 918 361 924 362
rect 982 362 983 366
rect 987 362 988 366
rect 982 361 988 362
rect 1038 362 1039 366
rect 1043 362 1044 366
rect 1038 361 1044 362
rect 1094 362 1095 366
rect 1099 362 1100 366
rect 1094 361 1100 362
rect 1113 362 1115 366
rect 1150 362 1151 366
rect 1155 362 1156 366
rect 1113 360 1146 362
rect 1150 361 1156 362
rect 1206 362 1207 366
rect 1211 362 1212 366
rect 1206 361 1212 362
rect 1254 362 1255 366
rect 1259 362 1260 366
rect 1254 361 1260 362
rect 1302 362 1303 366
rect 1307 362 1308 366
rect 1302 361 1308 362
rect 1350 362 1351 366
rect 1355 362 1356 366
rect 1350 361 1356 362
rect 1398 362 1399 366
rect 1403 362 1404 366
rect 1398 361 1404 362
rect 1446 362 1447 366
rect 1451 362 1452 366
rect 1446 361 1452 362
rect 1494 362 1495 366
rect 1499 362 1500 366
rect 1513 364 1535 366
rect 1534 363 1535 364
rect 1539 363 1540 367
rect 1534 362 1540 363
rect 1542 366 1548 367
rect 1559 366 1565 367
rect 1590 366 1596 367
rect 1607 366 1613 367
rect 1542 362 1543 366
rect 1547 362 1548 366
rect 1494 361 1500 362
rect 1542 361 1548 362
rect 1590 362 1591 366
rect 1595 362 1596 366
rect 1590 361 1596 362
rect 1144 358 1146 360
rect 1144 356 1150 358
rect 423 355 429 356
rect 423 354 424 355
rect 416 352 424 354
rect 367 350 373 351
rect 423 351 424 352
rect 428 351 429 355
rect 423 350 429 351
rect 479 355 485 356
rect 479 351 480 355
rect 484 354 485 355
rect 487 355 493 356
rect 487 354 488 355
rect 484 352 488 354
rect 484 351 485 352
rect 479 350 485 351
rect 487 351 488 352
rect 492 351 493 355
rect 487 350 493 351
rect 535 355 541 356
rect 535 351 536 355
rect 540 354 541 355
rect 543 355 549 356
rect 543 354 544 355
rect 540 352 544 354
rect 540 351 541 352
rect 535 350 541 351
rect 543 351 544 352
rect 548 351 549 355
rect 543 350 549 351
rect 591 355 597 356
rect 591 351 592 355
rect 596 354 597 355
rect 599 355 605 356
rect 599 354 600 355
rect 596 352 600 354
rect 596 351 597 352
rect 591 350 597 351
rect 599 351 600 352
rect 604 351 605 355
rect 599 350 605 351
rect 647 355 653 356
rect 647 351 648 355
rect 652 354 653 355
rect 670 355 676 356
rect 670 354 671 355
rect 652 352 671 354
rect 652 351 653 352
rect 647 350 653 351
rect 670 351 671 352
rect 675 351 676 355
rect 670 350 676 351
rect 698 355 709 356
rect 698 351 699 355
rect 703 351 704 355
rect 708 351 709 355
rect 698 350 709 351
rect 759 355 765 356
rect 759 351 760 355
rect 764 354 765 355
rect 767 355 773 356
rect 767 354 768 355
rect 764 352 768 354
rect 764 351 765 352
rect 759 350 765 351
rect 767 351 768 352
rect 772 351 773 355
rect 767 350 773 351
rect 814 355 821 356
rect 814 351 815 355
rect 820 351 821 355
rect 814 350 821 351
rect 871 355 877 356
rect 871 351 872 355
rect 876 354 877 355
rect 890 355 896 356
rect 890 354 891 355
rect 876 352 891 354
rect 876 351 877 352
rect 871 350 877 351
rect 890 351 891 352
rect 895 351 896 355
rect 890 350 896 351
rect 935 355 941 356
rect 935 351 936 355
rect 940 354 941 355
rect 943 355 949 356
rect 943 354 944 355
rect 940 352 944 354
rect 940 351 941 352
rect 935 350 941 351
rect 943 351 944 352
rect 948 351 949 355
rect 943 350 949 351
rect 999 355 1005 356
rect 999 351 1000 355
rect 1004 354 1005 355
rect 1007 355 1013 356
rect 1007 354 1008 355
rect 1004 352 1008 354
rect 1004 351 1005 352
rect 999 350 1005 351
rect 1007 351 1008 352
rect 1012 351 1013 355
rect 1007 350 1013 351
rect 1050 355 1061 356
rect 1050 351 1051 355
rect 1055 351 1056 355
rect 1060 351 1061 355
rect 1050 350 1061 351
rect 1110 355 1117 356
rect 1110 351 1111 355
rect 1116 351 1117 355
rect 1148 354 1161 356
rect 1167 355 1173 356
rect 1167 354 1168 355
rect 1159 352 1168 354
rect 1110 350 1117 351
rect 1167 351 1168 352
rect 1172 351 1173 355
rect 1167 350 1173 351
rect 1223 355 1229 356
rect 1223 351 1224 355
rect 1228 354 1229 355
rect 1238 355 1244 356
rect 1238 354 1239 355
rect 1228 352 1239 354
rect 1228 351 1229 352
rect 1223 350 1229 351
rect 1238 351 1239 352
rect 1243 351 1244 355
rect 1238 350 1244 351
rect 1271 355 1277 356
rect 1271 351 1272 355
rect 1276 354 1277 355
rect 1279 355 1285 356
rect 1279 354 1280 355
rect 1276 352 1280 354
rect 1276 351 1277 352
rect 1271 350 1277 351
rect 1279 351 1280 352
rect 1284 351 1285 355
rect 1279 350 1285 351
rect 1319 355 1325 356
rect 1319 351 1320 355
rect 1324 354 1325 355
rect 1327 355 1333 356
rect 1327 354 1328 355
rect 1324 352 1328 354
rect 1324 351 1325 352
rect 1319 350 1325 351
rect 1327 351 1328 352
rect 1332 351 1333 355
rect 1327 350 1333 351
rect 1367 355 1373 356
rect 1367 351 1368 355
rect 1372 354 1373 355
rect 1375 355 1381 356
rect 1375 354 1376 355
rect 1372 352 1376 354
rect 1372 351 1373 352
rect 1367 350 1373 351
rect 1375 351 1376 352
rect 1380 351 1381 355
rect 1375 350 1381 351
rect 1415 355 1421 356
rect 1415 351 1416 355
rect 1420 354 1421 355
rect 1438 355 1444 356
rect 1438 354 1439 355
rect 1420 352 1439 354
rect 1420 351 1421 352
rect 1415 350 1421 351
rect 1438 351 1439 352
rect 1443 351 1444 355
rect 1438 350 1444 351
rect 1463 355 1469 356
rect 1463 351 1464 355
rect 1468 351 1469 355
rect 1463 350 1469 351
rect 1511 355 1517 356
rect 1511 351 1512 355
rect 1516 354 1517 355
rect 1519 355 1525 356
rect 1519 354 1520 355
rect 1516 352 1520 354
rect 1516 351 1517 352
rect 1511 350 1517 351
rect 1519 351 1520 352
rect 1524 351 1525 355
rect 1519 350 1525 351
rect 1559 355 1565 356
rect 1559 351 1560 355
rect 1564 354 1565 355
rect 1567 355 1573 356
rect 1567 354 1568 355
rect 1564 352 1568 354
rect 1564 351 1565 352
rect 1559 350 1565 351
rect 1567 351 1568 352
rect 1572 351 1573 355
rect 1567 350 1573 351
rect 1607 355 1613 356
rect 1607 351 1608 355
rect 1612 354 1613 355
rect 1616 354 1618 372
rect 1639 371 1645 372
rect 1639 367 1640 371
rect 1644 367 1645 371
rect 1622 366 1628 367
rect 1639 366 1645 367
rect 1662 368 1668 369
rect 1622 362 1623 366
rect 1627 362 1628 366
rect 1662 364 1663 368
rect 1667 364 1668 368
rect 1662 363 1668 364
rect 1622 361 1628 362
rect 1612 352 1618 354
rect 1638 355 1645 356
rect 1612 351 1613 352
rect 1607 350 1613 351
rect 1638 351 1639 355
rect 1644 351 1645 355
rect 1638 350 1645 351
rect 1662 351 1668 352
rect 110 346 116 347
rect 134 349 140 350
rect 134 345 135 349
rect 139 345 140 349
rect 134 344 140 345
rect 166 349 172 350
rect 166 345 167 349
rect 171 345 172 349
rect 166 344 172 345
rect 198 349 204 350
rect 198 345 199 349
rect 203 345 204 349
rect 198 344 204 345
rect 238 349 244 350
rect 238 345 239 349
rect 243 345 244 349
rect 238 344 244 345
rect 294 349 300 350
rect 294 345 295 349
rect 299 345 300 349
rect 294 344 300 345
rect 350 349 356 350
rect 350 345 351 349
rect 355 345 356 349
rect 350 344 356 345
rect 406 349 412 350
rect 406 345 407 349
rect 411 345 412 349
rect 406 344 412 345
rect 462 349 468 350
rect 462 345 463 349
rect 467 345 468 349
rect 462 344 468 345
rect 518 349 524 350
rect 518 345 519 349
rect 523 345 524 349
rect 518 344 524 345
rect 574 349 580 350
rect 574 345 575 349
rect 579 345 580 349
rect 574 344 580 345
rect 630 349 636 350
rect 630 345 631 349
rect 635 345 636 349
rect 630 344 636 345
rect 686 349 692 350
rect 686 345 687 349
rect 691 345 692 349
rect 686 344 692 345
rect 742 349 748 350
rect 742 345 743 349
rect 747 345 748 349
rect 742 344 748 345
rect 798 349 804 350
rect 798 345 799 349
rect 803 345 804 349
rect 798 344 804 345
rect 854 349 860 350
rect 854 345 855 349
rect 859 345 860 349
rect 854 344 860 345
rect 918 349 924 350
rect 918 345 919 349
rect 923 345 924 349
rect 918 344 924 345
rect 982 349 988 350
rect 982 345 983 349
rect 987 345 988 349
rect 982 344 988 345
rect 1038 349 1044 350
rect 1038 345 1039 349
rect 1043 345 1044 349
rect 1038 344 1044 345
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1150 349 1156 350
rect 1150 345 1151 349
rect 1155 345 1156 349
rect 1150 344 1156 345
rect 1206 349 1212 350
rect 1206 345 1207 349
rect 1211 345 1212 349
rect 1206 344 1212 345
rect 1254 349 1260 350
rect 1254 345 1255 349
rect 1259 345 1260 349
rect 1254 344 1260 345
rect 1302 349 1308 350
rect 1302 345 1303 349
rect 1307 345 1308 349
rect 1302 344 1308 345
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1398 349 1404 350
rect 1398 345 1399 349
rect 1403 345 1404 349
rect 1398 344 1404 345
rect 1446 349 1452 350
rect 1446 345 1447 349
rect 1451 345 1452 349
rect 1446 344 1452 345
rect 150 343 156 344
rect 150 339 151 343
rect 155 342 156 343
rect 1367 343 1373 344
rect 155 340 187 342
rect 155 339 156 340
rect 150 338 156 339
rect 134 335 140 336
rect 110 333 116 334
rect 110 329 111 333
rect 115 329 116 333
rect 134 331 135 335
rect 139 331 140 335
rect 134 330 140 331
rect 166 335 172 336
rect 166 331 167 335
rect 171 331 172 335
rect 166 330 172 331
rect 110 328 116 329
rect 185 328 187 340
rect 1367 339 1368 343
rect 1372 342 1373 343
rect 1465 342 1467 350
rect 1494 349 1500 350
rect 1494 345 1495 349
rect 1499 345 1500 349
rect 1494 344 1500 345
rect 1542 349 1548 350
rect 1542 345 1543 349
rect 1547 345 1548 349
rect 1542 344 1548 345
rect 1590 349 1596 350
rect 1590 345 1591 349
rect 1595 345 1596 349
rect 1590 344 1596 345
rect 1622 349 1628 350
rect 1622 345 1623 349
rect 1627 345 1628 349
rect 1662 347 1663 351
rect 1667 347 1668 351
rect 1662 346 1668 347
rect 1622 344 1628 345
rect 1372 340 1467 342
rect 1372 339 1373 340
rect 1367 338 1373 339
rect 206 335 212 336
rect 206 331 207 335
rect 211 331 212 335
rect 206 330 212 331
rect 262 335 268 336
rect 262 331 263 335
rect 267 331 268 335
rect 262 330 268 331
rect 326 335 332 336
rect 326 331 327 335
rect 331 331 332 335
rect 326 330 332 331
rect 390 335 396 336
rect 390 331 391 335
rect 395 331 396 335
rect 390 330 396 331
rect 454 335 460 336
rect 454 331 455 335
rect 459 331 460 335
rect 454 330 460 331
rect 518 335 524 336
rect 518 331 519 335
rect 523 331 524 335
rect 518 330 524 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 686 335 692 336
rect 686 331 687 335
rect 691 331 692 335
rect 686 330 692 331
rect 750 335 756 336
rect 750 331 751 335
rect 755 331 756 335
rect 750 330 756 331
rect 814 335 820 336
rect 814 331 815 335
rect 819 331 820 335
rect 814 330 820 331
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 950 335 956 336
rect 950 331 951 335
rect 955 331 956 335
rect 950 330 956 331
rect 1030 335 1036 336
rect 1030 331 1031 335
rect 1035 331 1036 335
rect 1030 330 1036 331
rect 1110 335 1116 336
rect 1110 331 1111 335
rect 1115 331 1116 335
rect 1110 330 1116 331
rect 1190 335 1196 336
rect 1190 331 1191 335
rect 1195 331 1196 335
rect 1190 330 1196 331
rect 1270 335 1276 336
rect 1270 331 1271 335
rect 1275 331 1276 335
rect 1270 330 1276 331
rect 1342 335 1348 336
rect 1342 331 1343 335
rect 1347 331 1348 335
rect 1342 330 1348 331
rect 1406 335 1412 336
rect 1406 331 1407 335
rect 1411 331 1412 335
rect 1406 330 1412 331
rect 1462 335 1468 336
rect 1462 331 1463 335
rect 1467 331 1468 335
rect 1462 330 1468 331
rect 1518 335 1524 336
rect 1518 331 1519 335
rect 1523 331 1524 335
rect 1518 330 1524 331
rect 1534 335 1540 336
rect 1534 331 1535 335
rect 1539 334 1540 335
rect 1582 335 1588 336
rect 1539 332 1558 334
rect 1539 331 1540 332
rect 1534 330 1540 331
rect 151 327 157 328
rect 151 323 152 327
rect 156 326 157 327
rect 183 327 189 328
rect 156 324 178 326
rect 156 323 157 324
rect 151 322 157 323
rect 134 318 140 319
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 134 314 135 318
rect 139 314 140 318
rect 134 313 140 314
rect 166 318 172 319
rect 166 314 167 318
rect 171 314 172 318
rect 166 313 172 314
rect 110 311 116 312
rect 150 311 157 312
rect 150 307 151 311
rect 156 307 157 311
rect 176 310 178 324
rect 183 323 184 327
rect 188 323 189 327
rect 183 322 189 323
rect 223 327 229 328
rect 223 323 224 327
rect 228 326 229 327
rect 279 327 285 328
rect 228 324 274 326
rect 228 323 229 324
rect 223 322 229 323
rect 206 318 212 319
rect 206 314 207 318
rect 211 314 212 318
rect 206 313 212 314
rect 262 318 268 319
rect 262 314 263 318
rect 267 314 268 318
rect 262 313 268 314
rect 183 311 189 312
rect 183 310 184 311
rect 176 308 184 310
rect 150 306 157 307
rect 183 307 184 308
rect 188 307 189 311
rect 183 306 189 307
rect 223 311 229 312
rect 223 307 224 311
rect 228 310 229 311
rect 250 311 256 312
rect 250 310 251 311
rect 228 308 251 310
rect 228 307 229 308
rect 223 306 229 307
rect 250 307 251 308
rect 255 307 256 311
rect 272 310 274 324
rect 279 323 280 327
rect 284 323 285 327
rect 279 322 285 323
rect 343 327 349 328
rect 343 323 344 327
rect 348 323 349 327
rect 343 322 349 323
rect 407 327 413 328
rect 407 323 408 327
rect 412 326 413 327
rect 446 327 452 328
rect 446 326 447 327
rect 412 324 447 326
rect 412 323 413 324
rect 407 322 413 323
rect 446 323 447 324
rect 451 323 452 327
rect 446 322 452 323
rect 471 327 480 328
rect 471 323 472 327
rect 479 323 480 327
rect 535 327 541 328
rect 535 326 536 327
rect 471 322 480 323
rect 512 324 536 326
rect 281 318 283 322
rect 326 318 332 319
rect 281 316 314 318
rect 279 311 285 312
rect 279 310 280 311
rect 272 308 280 310
rect 250 306 256 307
rect 279 307 280 308
rect 284 307 285 311
rect 312 310 314 316
rect 326 314 327 318
rect 331 314 332 318
rect 345 318 347 322
rect 390 318 396 319
rect 345 316 378 318
rect 326 313 332 314
rect 343 311 349 312
rect 343 310 344 311
rect 312 308 344 310
rect 279 306 285 307
rect 343 307 344 308
rect 348 307 349 311
rect 376 310 378 316
rect 390 314 391 318
rect 395 314 396 318
rect 390 313 396 314
rect 454 318 460 319
rect 454 314 455 318
rect 459 314 460 318
rect 512 314 514 324
rect 535 323 536 324
rect 540 323 541 327
rect 535 322 541 323
rect 586 327 597 328
rect 586 323 587 327
rect 591 323 592 327
rect 596 323 597 327
rect 647 327 653 328
rect 647 326 648 327
rect 586 322 597 323
rect 620 324 648 326
rect 454 313 460 314
rect 508 312 514 314
rect 518 318 524 319
rect 518 314 519 318
rect 523 314 524 318
rect 518 313 524 314
rect 574 318 580 319
rect 574 314 575 318
rect 579 314 580 318
rect 574 313 580 314
rect 407 311 413 312
rect 407 310 408 311
rect 376 308 408 310
rect 343 306 349 307
rect 407 307 408 308
rect 412 307 413 311
rect 407 306 413 307
rect 471 311 477 312
rect 471 307 472 311
rect 476 310 477 311
rect 508 310 510 312
rect 476 308 510 310
rect 535 311 541 312
rect 476 307 477 308
rect 471 306 477 307
rect 535 307 536 311
rect 540 307 541 311
rect 535 306 541 307
rect 591 311 597 312
rect 591 307 592 311
rect 596 310 597 311
rect 620 310 622 324
rect 647 323 648 324
rect 652 323 653 327
rect 647 322 653 323
rect 655 327 661 328
rect 655 323 656 327
rect 660 326 661 327
rect 703 327 709 328
rect 703 326 704 327
rect 660 324 704 326
rect 660 323 661 324
rect 655 322 661 323
rect 703 323 704 324
rect 708 323 709 327
rect 767 327 773 328
rect 767 326 768 327
rect 703 322 709 323
rect 740 324 768 326
rect 630 318 636 319
rect 630 314 631 318
rect 635 314 636 318
rect 630 313 636 314
rect 686 318 692 319
rect 686 314 687 318
rect 691 314 692 318
rect 686 313 692 314
rect 596 308 622 310
rect 647 311 653 312
rect 596 307 597 308
rect 591 306 597 307
rect 647 307 648 311
rect 652 310 653 311
rect 694 311 700 312
rect 694 310 695 311
rect 652 308 695 310
rect 652 307 653 308
rect 647 306 653 307
rect 694 307 695 308
rect 699 307 700 311
rect 694 306 700 307
rect 703 311 709 312
rect 703 307 704 311
rect 708 310 709 311
rect 740 310 742 324
rect 767 323 768 324
rect 772 323 773 327
rect 767 322 773 323
rect 775 327 781 328
rect 775 323 776 327
rect 780 326 781 327
rect 831 327 837 328
rect 831 326 832 327
rect 780 324 832 326
rect 780 323 781 324
rect 775 322 781 323
rect 831 323 832 324
rect 836 323 837 327
rect 895 327 901 328
rect 895 326 896 327
rect 831 322 837 323
rect 872 324 896 326
rect 750 318 756 319
rect 750 314 751 318
rect 755 314 756 318
rect 750 313 756 314
rect 814 318 820 319
rect 814 314 815 318
rect 819 314 820 318
rect 872 314 874 324
rect 895 323 896 324
rect 900 323 901 327
rect 967 327 973 328
rect 967 326 968 327
rect 895 322 901 323
rect 932 324 968 326
rect 814 313 820 314
rect 868 312 874 314
rect 878 318 884 319
rect 878 314 879 318
rect 883 314 884 318
rect 878 313 884 314
rect 708 308 742 310
rect 767 311 773 312
rect 708 307 709 308
rect 703 306 709 307
rect 767 307 768 311
rect 772 307 773 311
rect 767 306 773 307
rect 831 311 837 312
rect 831 307 832 311
rect 836 310 837 311
rect 868 310 870 312
rect 836 308 870 310
rect 895 311 901 312
rect 836 307 837 308
rect 831 306 837 307
rect 895 307 896 311
rect 900 310 901 311
rect 932 310 934 324
rect 967 323 968 324
rect 972 323 973 327
rect 1047 327 1053 328
rect 1047 326 1048 327
rect 967 322 973 323
rect 1012 324 1048 326
rect 950 318 956 319
rect 950 314 951 318
rect 955 314 956 318
rect 950 313 956 314
rect 900 308 934 310
rect 967 311 973 312
rect 900 307 901 308
rect 895 306 901 307
rect 967 307 968 311
rect 972 310 973 311
rect 1012 310 1014 324
rect 1047 323 1048 324
rect 1052 323 1053 327
rect 1047 322 1053 323
rect 1127 327 1133 328
rect 1127 323 1128 327
rect 1132 326 1133 327
rect 1158 327 1164 328
rect 1158 326 1159 327
rect 1132 324 1159 326
rect 1132 323 1133 324
rect 1127 322 1133 323
rect 1158 323 1159 324
rect 1163 323 1164 327
rect 1207 327 1213 328
rect 1207 326 1208 327
rect 1158 322 1164 323
rect 1168 324 1208 326
rect 1030 318 1036 319
rect 1030 314 1031 318
rect 1035 314 1036 318
rect 1030 313 1036 314
rect 1110 318 1116 319
rect 1110 314 1111 318
rect 1115 314 1116 318
rect 1110 313 1116 314
rect 972 308 1014 310
rect 1047 311 1056 312
rect 972 307 973 308
rect 967 306 973 307
rect 1047 307 1048 311
rect 1055 307 1056 311
rect 1047 306 1056 307
rect 1127 311 1133 312
rect 1127 307 1128 311
rect 1132 310 1133 311
rect 1168 310 1170 324
rect 1207 323 1208 324
rect 1212 323 1213 327
rect 1287 327 1293 328
rect 1287 326 1288 327
rect 1207 322 1213 323
rect 1249 324 1288 326
rect 1190 318 1196 319
rect 1190 314 1191 318
rect 1195 314 1196 318
rect 1190 313 1196 314
rect 1132 308 1170 310
rect 1207 311 1213 312
rect 1132 307 1133 308
rect 1127 306 1133 307
rect 1207 307 1208 311
rect 1212 310 1213 311
rect 1249 310 1251 324
rect 1287 323 1288 324
rect 1292 323 1293 327
rect 1287 322 1293 323
rect 1359 327 1365 328
rect 1359 323 1360 327
rect 1364 323 1365 327
rect 1359 322 1365 323
rect 1423 327 1429 328
rect 1423 323 1424 327
rect 1428 326 1429 327
rect 1479 327 1485 328
rect 1428 324 1454 326
rect 1428 323 1429 324
rect 1423 322 1429 323
rect 1270 318 1276 319
rect 1270 314 1271 318
rect 1275 314 1276 318
rect 1270 313 1276 314
rect 1342 318 1348 319
rect 1342 314 1343 318
rect 1347 314 1348 318
rect 1361 318 1363 322
rect 1406 318 1412 319
rect 1361 316 1394 318
rect 1342 313 1348 314
rect 1212 308 1251 310
rect 1282 311 1293 312
rect 1212 307 1213 308
rect 1207 306 1213 307
rect 1282 307 1283 311
rect 1287 307 1288 311
rect 1292 307 1293 311
rect 1282 306 1293 307
rect 1359 311 1365 312
rect 1359 307 1360 311
rect 1364 310 1365 311
rect 1367 311 1373 312
rect 1367 310 1368 311
rect 1364 308 1368 310
rect 1364 307 1365 308
rect 1359 306 1365 307
rect 1367 307 1368 308
rect 1372 307 1373 311
rect 1392 310 1394 316
rect 1406 314 1407 318
rect 1411 314 1412 318
rect 1406 313 1412 314
rect 1423 311 1429 312
rect 1423 310 1424 311
rect 1392 308 1424 310
rect 1367 306 1373 307
rect 1423 307 1424 308
rect 1428 307 1429 311
rect 1452 310 1454 324
rect 1479 323 1480 327
rect 1484 323 1485 327
rect 1479 322 1485 323
rect 1535 327 1541 328
rect 1535 323 1536 327
rect 1540 323 1541 327
rect 1556 326 1558 332
rect 1582 331 1583 335
rect 1587 331 1588 335
rect 1582 330 1588 331
rect 1622 335 1628 336
rect 1622 331 1623 335
rect 1627 331 1628 335
rect 1622 330 1628 331
rect 1662 333 1668 334
rect 1662 329 1663 333
rect 1667 329 1668 333
rect 1662 328 1668 329
rect 1599 327 1605 328
rect 1599 326 1600 327
rect 1556 324 1600 326
rect 1535 322 1541 323
rect 1599 323 1600 324
rect 1604 323 1605 327
rect 1599 322 1605 323
rect 1639 327 1645 328
rect 1639 323 1640 327
rect 1644 326 1645 327
rect 1647 327 1653 328
rect 1647 326 1648 327
rect 1644 324 1648 326
rect 1644 323 1645 324
rect 1639 322 1645 323
rect 1647 323 1648 324
rect 1652 323 1653 327
rect 1647 322 1653 323
rect 1481 320 1499 322
rect 1462 318 1468 319
rect 1462 314 1463 318
rect 1467 314 1468 318
rect 1462 313 1468 314
rect 1479 311 1485 312
rect 1479 310 1480 311
rect 1452 308 1480 310
rect 1423 306 1429 307
rect 1479 307 1480 308
rect 1484 307 1485 311
rect 1497 310 1499 320
rect 1518 318 1524 319
rect 1518 314 1519 318
rect 1523 314 1524 318
rect 1537 318 1539 322
rect 1582 318 1588 319
rect 1537 316 1570 318
rect 1518 313 1524 314
rect 1535 311 1541 312
rect 1535 310 1536 311
rect 1497 308 1536 310
rect 1479 306 1485 307
rect 1535 307 1536 308
rect 1540 307 1541 311
rect 1568 310 1570 316
rect 1582 314 1583 318
rect 1587 314 1588 318
rect 1582 313 1588 314
rect 1622 318 1628 319
rect 1622 314 1623 318
rect 1627 314 1628 318
rect 1622 313 1628 314
rect 1662 316 1668 317
rect 1662 312 1663 316
rect 1667 312 1668 316
rect 1599 311 1605 312
rect 1599 310 1600 311
rect 1568 308 1600 310
rect 1535 306 1541 307
rect 1599 307 1600 308
rect 1604 307 1605 311
rect 1599 306 1605 307
rect 1638 311 1645 312
rect 1662 311 1668 312
rect 1638 307 1639 311
rect 1644 307 1645 311
rect 1638 306 1645 307
rect 537 302 539 306
rect 655 303 661 304
rect 655 302 656 303
rect 537 300 656 302
rect 246 299 252 300
rect 246 298 247 299
rect 185 296 247 298
rect 153 292 178 294
rect 185 292 187 296
rect 246 295 247 296
rect 251 295 252 299
rect 655 299 656 300
rect 660 299 661 303
rect 655 298 661 299
rect 706 303 712 304
rect 706 299 707 303
rect 711 302 712 303
rect 769 302 771 306
rect 711 300 771 302
rect 711 299 712 300
rect 706 298 712 299
rect 246 294 252 295
rect 783 295 789 296
rect 319 292 378 294
rect 151 291 157 292
rect 110 288 116 289
rect 110 284 111 288
rect 115 284 116 288
rect 151 287 152 291
rect 156 287 157 291
rect 110 283 116 284
rect 134 286 140 287
rect 151 286 157 287
rect 166 286 172 287
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 150 275 157 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 150 271 151 275
rect 156 271 157 275
rect 176 274 178 292
rect 183 291 189 292
rect 183 287 184 291
rect 188 287 189 291
rect 238 291 244 292
rect 238 287 239 291
rect 243 290 244 291
rect 247 291 253 292
rect 247 290 248 291
rect 243 288 248 290
rect 243 287 244 288
rect 183 286 189 287
rect 230 286 236 287
rect 238 286 244 287
rect 247 287 248 288
rect 252 287 253 291
rect 311 291 317 292
rect 311 287 312 291
rect 316 290 317 291
rect 319 290 321 292
rect 316 288 321 290
rect 316 287 317 288
rect 247 286 253 287
rect 294 286 300 287
rect 311 286 317 287
rect 366 286 372 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 366 282 367 286
rect 371 282 372 286
rect 366 281 372 282
rect 183 275 189 276
rect 183 274 184 275
rect 176 272 184 274
rect 150 270 157 271
rect 183 271 184 272
rect 188 271 189 275
rect 183 270 189 271
rect 246 275 253 276
rect 246 271 247 275
rect 252 271 253 275
rect 246 270 253 271
rect 306 275 317 276
rect 306 271 307 275
rect 311 271 312 275
rect 316 271 317 275
rect 376 274 378 292
rect 383 291 389 292
rect 383 287 384 291
rect 388 290 389 291
rect 446 291 452 292
rect 388 288 426 290
rect 388 287 389 288
rect 383 286 389 287
rect 424 278 426 288
rect 446 287 447 291
rect 451 290 452 291
rect 455 291 461 292
rect 455 290 456 291
rect 451 288 456 290
rect 451 287 452 288
rect 438 286 444 287
rect 446 286 452 287
rect 455 287 456 288
rect 460 287 461 291
rect 519 291 525 292
rect 519 287 520 291
rect 524 290 525 291
rect 583 291 592 292
rect 524 288 562 290
rect 524 287 525 288
rect 455 286 461 287
rect 502 286 508 287
rect 519 286 525 287
rect 438 282 439 286
rect 443 282 444 286
rect 438 281 444 282
rect 502 282 503 286
rect 507 282 508 286
rect 502 281 508 282
rect 560 278 562 288
rect 583 287 584 291
rect 591 287 592 291
rect 647 291 653 292
rect 647 287 648 291
rect 652 290 653 291
rect 678 291 684 292
rect 678 290 679 291
rect 652 288 679 290
rect 652 287 653 288
rect 566 286 572 287
rect 583 286 592 287
rect 630 286 636 287
rect 647 286 653 287
rect 678 287 679 288
rect 683 287 684 291
rect 703 291 709 292
rect 703 290 704 291
rect 696 288 704 290
rect 678 286 684 287
rect 686 286 692 287
rect 566 282 567 286
rect 571 282 572 286
rect 566 281 572 282
rect 630 282 631 286
rect 635 282 636 286
rect 630 281 636 282
rect 686 282 687 286
rect 691 282 692 286
rect 686 281 692 282
rect 424 276 438 278
rect 560 276 566 278
rect 696 276 698 288
rect 703 287 704 288
rect 708 287 709 291
rect 759 291 765 292
rect 759 287 760 291
rect 764 290 765 291
rect 775 291 781 292
rect 775 290 776 291
rect 764 288 776 290
rect 764 287 765 288
rect 703 286 709 287
rect 742 286 748 287
rect 759 286 765 287
rect 775 287 776 288
rect 780 287 781 291
rect 783 291 784 295
rect 788 294 789 295
rect 831 295 837 296
rect 788 292 818 294
rect 788 291 789 292
rect 783 290 789 291
rect 816 290 818 292
rect 823 291 829 292
rect 823 290 824 291
rect 816 288 824 290
rect 823 287 824 288
rect 828 287 829 291
rect 831 291 832 295
rect 836 294 837 295
rect 903 295 909 296
rect 836 292 899 294
rect 836 291 837 292
rect 831 290 837 291
rect 895 291 901 292
rect 895 287 896 291
rect 900 287 901 291
rect 903 291 904 295
rect 908 294 909 295
rect 975 295 981 296
rect 908 292 971 294
rect 908 291 909 292
rect 903 290 909 291
rect 967 291 973 292
rect 967 287 968 291
rect 972 287 973 291
rect 975 291 976 295
rect 980 294 981 295
rect 1135 295 1141 296
rect 980 292 1051 294
rect 980 291 981 292
rect 975 290 981 291
rect 1047 291 1053 292
rect 1047 287 1048 291
rect 1052 287 1053 291
rect 1126 291 1133 292
rect 1126 287 1127 291
rect 1132 287 1133 291
rect 1135 291 1136 295
rect 1140 294 1141 295
rect 1215 295 1221 296
rect 1140 292 1211 294
rect 1140 291 1141 292
rect 1135 290 1141 291
rect 1207 291 1213 292
rect 1207 287 1208 291
rect 1212 287 1213 291
rect 1215 291 1216 295
rect 1220 294 1221 295
rect 1351 295 1357 296
rect 1220 292 1274 294
rect 1220 291 1221 292
rect 1215 290 1221 291
rect 1272 290 1274 292
rect 1279 291 1285 292
rect 1279 290 1280 291
rect 1272 288 1280 290
rect 1279 287 1280 288
rect 1284 287 1285 291
rect 1342 291 1349 292
rect 1342 287 1343 291
rect 1348 287 1349 291
rect 1351 291 1352 295
rect 1356 294 1357 295
rect 1356 292 1402 294
rect 1488 292 1506 294
rect 1537 292 1554 294
rect 1584 292 1602 294
rect 1616 292 1634 294
rect 1356 291 1357 292
rect 1351 290 1357 291
rect 1400 290 1402 292
rect 1407 291 1413 292
rect 1407 290 1408 291
rect 1400 288 1408 290
rect 1407 287 1408 288
rect 1412 287 1413 291
rect 1463 291 1469 292
rect 1463 287 1464 291
rect 1468 290 1469 291
rect 1488 290 1490 292
rect 1468 288 1490 290
rect 1468 287 1469 288
rect 775 286 781 287
rect 806 286 812 287
rect 823 286 829 287
rect 878 286 884 287
rect 895 286 901 287
rect 950 286 956 287
rect 967 286 973 287
rect 1030 286 1036 287
rect 1047 286 1053 287
rect 1110 286 1116 287
rect 1126 286 1133 287
rect 1190 286 1196 287
rect 1207 286 1213 287
rect 1262 286 1268 287
rect 1279 286 1285 287
rect 1326 286 1332 287
rect 1342 286 1349 287
rect 1390 286 1396 287
rect 1407 286 1413 287
rect 1446 286 1452 287
rect 1463 286 1469 287
rect 1494 286 1500 287
rect 742 282 743 286
rect 747 282 748 286
rect 742 281 748 282
rect 806 282 807 286
rect 811 282 812 286
rect 806 281 812 282
rect 878 282 879 286
rect 883 282 884 286
rect 878 281 884 282
rect 950 282 951 286
rect 955 282 956 286
rect 950 281 956 282
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1110 282 1111 286
rect 1115 282 1116 286
rect 1110 281 1116 282
rect 1190 282 1191 286
rect 1195 282 1196 286
rect 1190 281 1196 282
rect 1262 282 1263 286
rect 1267 282 1268 286
rect 1262 281 1268 282
rect 1326 282 1327 286
rect 1331 282 1332 286
rect 1326 281 1332 282
rect 1390 282 1391 286
rect 1395 282 1396 286
rect 1390 281 1396 282
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1494 282 1495 286
rect 1499 282 1500 286
rect 1494 281 1500 282
rect 383 275 389 276
rect 383 274 384 275
rect 376 272 384 274
rect 306 270 317 271
rect 383 271 384 272
rect 388 271 389 275
rect 436 274 450 276
rect 455 275 461 276
rect 455 274 456 275
rect 448 272 456 274
rect 383 270 389 271
rect 455 271 456 272
rect 460 271 461 275
rect 455 270 461 271
rect 519 275 525 276
rect 519 271 520 275
rect 524 274 525 275
rect 534 275 540 276
rect 534 274 535 275
rect 524 272 535 274
rect 524 271 525 272
rect 519 270 525 271
rect 534 271 535 272
rect 539 271 540 275
rect 564 274 578 276
rect 583 275 589 276
rect 583 274 584 275
rect 576 272 584 274
rect 534 270 540 271
rect 583 271 584 272
rect 588 271 589 275
rect 583 270 589 271
rect 647 275 653 276
rect 647 271 648 275
rect 652 274 653 275
rect 684 274 698 276
rect 703 275 712 276
rect 652 272 686 274
rect 652 271 653 272
rect 647 270 653 271
rect 703 271 704 275
rect 711 271 712 275
rect 703 270 712 271
rect 759 275 765 276
rect 759 271 760 275
rect 764 274 765 275
rect 783 275 789 276
rect 783 274 784 275
rect 764 272 784 274
rect 764 271 765 272
rect 759 270 765 271
rect 783 271 784 272
rect 788 271 789 275
rect 783 270 789 271
rect 823 275 829 276
rect 823 271 824 275
rect 828 274 829 275
rect 831 275 837 276
rect 831 274 832 275
rect 828 272 832 274
rect 828 271 829 272
rect 823 270 829 271
rect 831 271 832 272
rect 836 271 837 275
rect 831 270 837 271
rect 895 275 901 276
rect 895 271 896 275
rect 900 274 901 275
rect 903 275 909 276
rect 903 274 904 275
rect 900 272 904 274
rect 900 271 901 272
rect 895 270 901 271
rect 903 271 904 272
rect 908 271 909 275
rect 903 270 909 271
rect 967 275 973 276
rect 967 271 968 275
rect 972 274 973 275
rect 975 275 981 276
rect 975 274 976 275
rect 972 272 976 274
rect 972 271 973 272
rect 967 270 973 271
rect 975 271 976 272
rect 980 271 981 275
rect 975 270 981 271
rect 1047 275 1053 276
rect 1047 271 1048 275
rect 1052 271 1053 275
rect 1047 270 1053 271
rect 1127 275 1133 276
rect 1127 271 1128 275
rect 1132 274 1133 275
rect 1135 275 1141 276
rect 1135 274 1136 275
rect 1132 272 1136 274
rect 1132 271 1133 272
rect 1127 270 1133 271
rect 1135 271 1136 272
rect 1140 271 1141 275
rect 1135 270 1141 271
rect 1207 275 1213 276
rect 1207 271 1208 275
rect 1212 274 1213 275
rect 1215 275 1221 276
rect 1215 274 1216 275
rect 1212 272 1216 274
rect 1212 271 1213 272
rect 1207 270 1213 271
rect 1215 271 1216 272
rect 1220 271 1221 275
rect 1215 270 1221 271
rect 1279 275 1288 276
rect 1279 271 1280 275
rect 1287 271 1288 275
rect 1279 270 1288 271
rect 1343 275 1349 276
rect 1343 271 1344 275
rect 1348 274 1349 275
rect 1351 275 1357 276
rect 1351 274 1352 275
rect 1348 272 1352 274
rect 1348 271 1349 272
rect 1343 270 1349 271
rect 1351 271 1352 272
rect 1356 271 1357 275
rect 1351 270 1357 271
rect 1407 275 1413 276
rect 1407 271 1408 275
rect 1412 274 1413 275
rect 1430 275 1436 276
rect 1430 274 1431 275
rect 1412 272 1431 274
rect 1412 271 1413 272
rect 1407 270 1413 271
rect 1430 271 1431 272
rect 1435 271 1436 275
rect 1463 275 1469 276
rect 1463 274 1464 275
rect 1430 270 1436 271
rect 1456 272 1464 274
rect 110 266 116 267
rect 134 269 140 270
rect 134 265 135 269
rect 139 265 140 269
rect 134 264 140 265
rect 166 269 172 270
rect 166 265 167 269
rect 171 265 172 269
rect 166 264 172 265
rect 230 269 236 270
rect 230 265 231 269
rect 235 265 236 269
rect 230 264 236 265
rect 294 269 300 270
rect 294 265 295 269
rect 299 265 300 269
rect 294 264 300 265
rect 366 269 372 270
rect 366 265 367 269
rect 371 265 372 269
rect 366 264 372 265
rect 438 269 444 270
rect 438 265 439 269
rect 443 265 444 269
rect 438 264 444 265
rect 502 269 508 270
rect 502 265 503 269
rect 507 265 508 269
rect 502 264 508 265
rect 566 269 572 270
rect 566 265 567 269
rect 571 265 572 269
rect 566 264 572 265
rect 630 269 636 270
rect 630 265 631 269
rect 635 265 636 269
rect 630 264 636 265
rect 686 269 692 270
rect 686 265 687 269
rect 691 265 692 269
rect 686 264 692 265
rect 742 269 748 270
rect 742 265 743 269
rect 747 265 748 269
rect 742 264 748 265
rect 806 269 812 270
rect 806 265 807 269
rect 811 265 812 269
rect 806 264 812 265
rect 878 269 884 270
rect 878 265 879 269
rect 883 265 884 269
rect 878 264 884 265
rect 950 269 956 270
rect 950 265 951 269
rect 955 265 956 269
rect 950 264 956 265
rect 1030 269 1036 270
rect 1030 265 1031 269
rect 1035 265 1036 269
rect 1030 264 1036 265
rect 914 263 920 264
rect 914 259 915 263
rect 919 262 920 263
rect 1049 262 1051 270
rect 1110 269 1116 270
rect 1110 265 1111 269
rect 1115 265 1116 269
rect 1110 264 1116 265
rect 1190 269 1196 270
rect 1190 265 1191 269
rect 1195 265 1196 269
rect 1190 264 1196 265
rect 1262 269 1268 270
rect 1262 265 1263 269
rect 1267 265 1268 269
rect 1262 264 1268 265
rect 1326 269 1332 270
rect 1326 265 1327 269
rect 1331 265 1332 269
rect 1326 264 1332 265
rect 1390 269 1396 270
rect 1390 265 1391 269
rect 1395 265 1396 269
rect 1390 264 1396 265
rect 1446 269 1452 270
rect 1446 265 1447 269
rect 1451 265 1452 269
rect 1446 264 1452 265
rect 919 260 1051 262
rect 1342 263 1348 264
rect 919 259 920 260
rect 914 258 920 259
rect 1126 259 1132 260
rect 1126 255 1127 259
rect 1131 258 1132 259
rect 1342 259 1343 263
rect 1347 262 1348 263
rect 1456 262 1458 272
rect 1463 271 1464 272
rect 1468 271 1469 275
rect 1504 274 1506 292
rect 1511 291 1517 292
rect 1511 287 1512 291
rect 1516 290 1517 291
rect 1537 290 1539 292
rect 1516 288 1539 290
rect 1516 287 1517 288
rect 1511 286 1517 287
rect 1542 286 1548 287
rect 1542 282 1543 286
rect 1547 282 1548 286
rect 1542 281 1548 282
rect 1511 275 1517 276
rect 1511 274 1512 275
rect 1504 272 1512 274
rect 1463 270 1469 271
rect 1511 271 1512 272
rect 1516 271 1517 275
rect 1552 274 1554 292
rect 1559 291 1565 292
rect 1559 287 1560 291
rect 1564 290 1565 291
rect 1584 290 1586 292
rect 1564 288 1586 290
rect 1564 287 1565 288
rect 1559 286 1565 287
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1559 275 1565 276
rect 1559 274 1560 275
rect 1552 272 1560 274
rect 1511 270 1517 271
rect 1559 271 1560 272
rect 1564 271 1565 275
rect 1600 274 1602 292
rect 1607 291 1613 292
rect 1607 287 1608 291
rect 1612 290 1613 291
rect 1616 290 1618 292
rect 1612 288 1618 290
rect 1612 287 1613 288
rect 1607 286 1613 287
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1622 281 1628 282
rect 1632 278 1634 292
rect 1639 291 1645 292
rect 1639 287 1640 291
rect 1644 290 1645 291
rect 1647 291 1653 292
rect 1647 290 1648 291
rect 1644 288 1648 290
rect 1644 287 1645 288
rect 1639 286 1645 287
rect 1647 287 1648 288
rect 1652 287 1653 291
rect 1647 286 1653 287
rect 1662 288 1668 289
rect 1662 284 1663 288
rect 1667 284 1668 288
rect 1662 283 1668 284
rect 1632 276 1643 278
rect 1607 275 1613 276
rect 1607 274 1608 275
rect 1600 272 1608 274
rect 1559 270 1565 271
rect 1607 271 1608 272
rect 1612 271 1613 275
rect 1607 270 1613 271
rect 1639 275 1645 276
rect 1639 271 1640 275
rect 1644 271 1645 275
rect 1639 270 1645 271
rect 1662 271 1668 272
rect 1494 269 1500 270
rect 1494 265 1495 269
rect 1499 265 1500 269
rect 1494 264 1500 265
rect 1542 269 1548 270
rect 1542 265 1543 269
rect 1547 265 1548 269
rect 1542 264 1548 265
rect 1590 269 1596 270
rect 1590 265 1591 269
rect 1595 265 1596 269
rect 1590 264 1596 265
rect 1622 269 1628 270
rect 1622 265 1623 269
rect 1627 265 1628 269
rect 1662 267 1663 271
rect 1667 267 1668 271
rect 1662 266 1668 267
rect 1622 264 1628 265
rect 1347 260 1458 262
rect 1347 259 1348 260
rect 1342 258 1348 259
rect 1131 256 1251 258
rect 1131 255 1132 256
rect 1126 254 1132 255
rect 134 251 140 252
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 247 135 251
rect 139 247 140 251
rect 134 246 140 247
rect 174 251 180 252
rect 174 247 175 251
rect 179 247 180 251
rect 174 246 180 247
rect 246 251 252 252
rect 246 247 247 251
rect 251 247 252 251
rect 246 246 252 247
rect 318 251 324 252
rect 318 247 319 251
rect 323 247 324 251
rect 318 246 324 247
rect 382 251 388 252
rect 382 247 383 251
rect 387 247 388 251
rect 382 246 388 247
rect 446 251 452 252
rect 446 247 447 251
rect 451 247 452 251
rect 446 246 452 247
rect 518 251 524 252
rect 518 247 519 251
rect 523 247 524 251
rect 518 246 524 247
rect 590 251 596 252
rect 590 247 591 251
rect 595 247 596 251
rect 590 246 596 247
rect 662 251 668 252
rect 662 247 663 251
rect 667 247 668 251
rect 662 246 668 247
rect 742 251 748 252
rect 742 247 743 251
rect 747 247 748 251
rect 742 246 748 247
rect 822 251 828 252
rect 822 247 823 251
rect 827 247 828 251
rect 822 246 828 247
rect 894 251 900 252
rect 894 247 895 251
rect 899 247 900 251
rect 894 246 900 247
rect 966 251 972 252
rect 966 247 967 251
rect 971 247 972 251
rect 966 246 972 247
rect 1030 251 1036 252
rect 1030 247 1031 251
rect 1035 247 1036 251
rect 1030 246 1036 247
rect 1086 251 1092 252
rect 1086 247 1087 251
rect 1091 247 1092 251
rect 1086 246 1092 247
rect 1142 251 1148 252
rect 1142 247 1143 251
rect 1147 247 1148 251
rect 1142 246 1148 247
rect 1198 251 1204 252
rect 1198 247 1199 251
rect 1203 247 1204 251
rect 1198 246 1204 247
rect 110 244 116 245
rect 151 243 157 244
rect 151 239 152 243
rect 156 242 157 243
rect 191 243 197 244
rect 156 240 186 242
rect 156 239 157 240
rect 151 238 157 239
rect 134 234 140 235
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 134 230 135 234
rect 139 230 140 234
rect 134 229 140 230
rect 174 234 180 235
rect 174 230 175 234
rect 179 230 180 234
rect 174 229 180 230
rect 110 227 116 228
rect 150 227 157 228
rect 150 223 151 227
rect 156 223 157 227
rect 184 226 186 240
rect 191 239 192 243
rect 196 242 197 243
rect 238 243 244 244
rect 238 242 239 243
rect 196 240 239 242
rect 196 239 197 240
rect 191 238 197 239
rect 238 239 239 240
rect 243 239 244 243
rect 238 238 244 239
rect 263 243 269 244
rect 263 239 264 243
rect 268 242 269 243
rect 335 243 341 244
rect 268 240 330 242
rect 268 239 269 240
rect 263 238 269 239
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 318 234 324 235
rect 318 230 319 234
rect 323 230 324 234
rect 318 229 324 230
rect 191 227 197 228
rect 191 226 192 227
rect 184 224 192 226
rect 150 222 157 223
rect 191 223 192 224
rect 196 223 197 227
rect 191 222 197 223
rect 263 227 269 228
rect 263 223 264 227
rect 268 226 269 227
rect 306 227 312 228
rect 306 226 307 227
rect 268 224 307 226
rect 268 223 269 224
rect 263 222 269 223
rect 306 223 307 224
rect 311 223 312 227
rect 328 226 330 240
rect 335 239 336 243
rect 340 242 341 243
rect 399 243 405 244
rect 340 240 370 242
rect 340 239 341 240
rect 335 238 341 239
rect 335 227 341 228
rect 335 226 336 227
rect 328 224 336 226
rect 306 222 312 223
rect 335 223 336 224
rect 340 223 341 227
rect 368 226 370 240
rect 399 239 400 243
rect 404 242 405 243
rect 438 243 444 244
rect 404 240 434 242
rect 404 239 405 240
rect 399 238 405 239
rect 382 234 388 235
rect 382 230 383 234
rect 387 230 388 234
rect 382 229 388 230
rect 399 227 405 228
rect 399 226 400 227
rect 368 224 400 226
rect 335 222 341 223
rect 399 223 400 224
rect 404 223 405 227
rect 432 226 434 240
rect 438 239 439 243
rect 443 242 444 243
rect 463 243 469 244
rect 463 242 464 243
rect 443 240 464 242
rect 443 239 444 240
rect 438 238 444 239
rect 463 239 464 240
rect 468 239 469 243
rect 463 238 469 239
rect 535 243 541 244
rect 535 239 536 243
rect 540 239 541 243
rect 535 238 541 239
rect 574 243 580 244
rect 574 239 575 243
rect 579 242 580 243
rect 607 243 613 244
rect 607 242 608 243
rect 579 240 608 242
rect 579 239 580 240
rect 574 238 580 239
rect 607 239 608 240
rect 612 239 613 243
rect 607 238 613 239
rect 678 243 685 244
rect 678 239 679 243
rect 684 239 685 243
rect 759 243 765 244
rect 759 242 760 243
rect 678 238 685 239
rect 724 240 760 242
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 518 234 524 235
rect 518 230 519 234
rect 523 230 524 234
rect 537 234 539 238
rect 590 234 596 235
rect 537 232 574 234
rect 518 229 524 230
rect 463 227 469 228
rect 463 226 464 227
rect 432 224 464 226
rect 399 222 405 223
rect 463 223 464 224
rect 468 223 469 227
rect 463 222 469 223
rect 534 227 541 228
rect 534 223 535 227
rect 540 223 541 227
rect 572 226 574 232
rect 590 230 591 234
rect 595 230 596 234
rect 590 229 596 230
rect 662 234 668 235
rect 662 230 663 234
rect 667 230 668 234
rect 662 229 668 230
rect 607 227 613 228
rect 607 226 608 227
rect 572 224 608 226
rect 534 222 541 223
rect 607 223 608 224
rect 612 223 613 227
rect 607 222 613 223
rect 679 227 685 228
rect 679 223 680 227
rect 684 226 685 227
rect 724 226 726 240
rect 759 239 760 240
rect 764 239 765 243
rect 839 243 845 244
rect 839 242 840 243
rect 759 238 765 239
rect 804 240 840 242
rect 742 234 748 235
rect 742 230 743 234
rect 747 230 748 234
rect 742 229 748 230
rect 684 224 726 226
rect 759 227 765 228
rect 684 223 685 224
rect 679 222 685 223
rect 759 223 760 227
rect 764 226 765 227
rect 804 226 806 240
rect 839 239 840 240
rect 844 239 845 243
rect 911 243 917 244
rect 911 242 912 243
rect 839 238 845 239
rect 876 240 912 242
rect 822 234 828 235
rect 822 230 823 234
rect 827 230 828 234
rect 822 229 828 230
rect 764 224 806 226
rect 839 227 845 228
rect 764 223 765 224
rect 759 222 765 223
rect 839 223 840 227
rect 844 226 845 227
rect 876 226 878 240
rect 911 239 912 240
rect 916 239 917 243
rect 911 238 917 239
rect 983 243 989 244
rect 983 239 984 243
rect 988 242 989 243
rect 1047 243 1053 244
rect 988 240 1018 242
rect 988 239 989 240
rect 983 238 989 239
rect 894 234 900 235
rect 894 230 895 234
rect 899 230 900 234
rect 894 229 900 230
rect 966 234 972 235
rect 966 230 967 234
rect 971 230 972 234
rect 966 229 972 230
rect 844 224 878 226
rect 911 227 920 228
rect 844 223 845 224
rect 839 222 845 223
rect 911 223 912 227
rect 919 223 920 227
rect 911 222 920 223
rect 983 227 989 228
rect 983 223 984 227
rect 988 226 989 227
rect 1016 226 1018 240
rect 1047 239 1048 243
rect 1052 242 1053 243
rect 1103 243 1109 244
rect 1052 240 1098 242
rect 1052 239 1053 240
rect 1047 238 1053 239
rect 1030 234 1036 235
rect 1030 230 1031 234
rect 1035 230 1036 234
rect 1030 229 1036 230
rect 1086 234 1092 235
rect 1086 230 1087 234
rect 1091 230 1092 234
rect 1086 229 1092 230
rect 1047 227 1053 228
rect 1047 226 1048 227
rect 988 224 1014 226
rect 1016 224 1048 226
rect 988 223 989 224
rect 983 222 989 223
rect 438 219 444 220
rect 438 218 439 219
rect 368 216 439 218
rect 153 208 178 210
rect 185 208 218 210
rect 296 208 314 210
rect 151 207 157 208
rect 110 204 116 205
rect 110 200 111 204
rect 115 200 116 204
rect 151 203 152 207
rect 156 203 157 207
rect 110 199 116 200
rect 134 202 140 203
rect 151 202 157 203
rect 166 202 172 203
rect 134 198 135 202
rect 139 198 140 202
rect 134 197 140 198
rect 166 198 167 202
rect 171 198 172 202
rect 166 197 172 198
rect 150 191 157 192
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 150 187 151 191
rect 156 187 157 191
rect 176 190 178 208
rect 183 207 189 208
rect 183 203 184 207
rect 188 203 189 207
rect 183 202 189 203
rect 206 202 212 203
rect 206 198 207 202
rect 211 198 212 202
rect 206 197 212 198
rect 183 191 189 192
rect 183 190 184 191
rect 176 188 184 190
rect 150 186 157 187
rect 183 187 184 188
rect 188 187 189 191
rect 216 190 218 208
rect 223 207 229 208
rect 223 203 224 207
rect 228 206 229 207
rect 246 207 252 208
rect 246 206 247 207
rect 228 204 247 206
rect 228 203 229 204
rect 223 202 229 203
rect 246 203 247 204
rect 251 203 252 207
rect 271 207 277 208
rect 271 203 272 207
rect 276 206 277 207
rect 296 206 298 208
rect 276 204 298 206
rect 276 203 277 204
rect 246 202 252 203
rect 254 202 260 203
rect 271 202 277 203
rect 302 202 308 203
rect 254 198 255 202
rect 259 198 260 202
rect 254 197 260 198
rect 302 198 303 202
rect 307 198 308 202
rect 302 197 308 198
rect 223 191 229 192
rect 223 190 224 191
rect 216 188 224 190
rect 183 186 189 187
rect 223 187 224 188
rect 228 187 229 191
rect 223 186 229 187
rect 271 191 277 192
rect 271 187 272 191
rect 276 190 277 191
rect 294 191 300 192
rect 294 190 295 191
rect 276 188 295 190
rect 276 187 277 188
rect 271 186 277 187
rect 294 187 295 188
rect 299 187 300 191
rect 312 190 314 208
rect 319 207 325 208
rect 319 203 320 207
rect 324 206 325 207
rect 359 207 365 208
rect 324 204 338 206
rect 324 203 325 204
rect 319 202 325 203
rect 336 194 338 204
rect 359 203 360 207
rect 364 206 365 207
rect 368 206 370 216
rect 438 215 439 216
rect 443 215 444 219
rect 1012 218 1014 224
rect 1047 223 1048 224
rect 1052 223 1053 227
rect 1096 226 1098 240
rect 1103 239 1104 243
rect 1108 242 1109 243
rect 1159 243 1165 244
rect 1108 240 1131 242
rect 1108 239 1109 240
rect 1103 238 1109 239
rect 1103 227 1109 228
rect 1103 226 1104 227
rect 1096 224 1104 226
rect 1047 222 1053 223
rect 1103 223 1104 224
rect 1108 223 1109 227
rect 1129 226 1131 240
rect 1159 239 1160 243
rect 1164 242 1165 243
rect 1215 243 1221 244
rect 1164 240 1190 242
rect 1164 239 1165 240
rect 1159 238 1165 239
rect 1142 234 1148 235
rect 1142 230 1143 234
rect 1147 230 1148 234
rect 1142 229 1148 230
rect 1159 227 1165 228
rect 1159 226 1160 227
rect 1129 224 1160 226
rect 1103 222 1109 223
rect 1159 223 1160 224
rect 1164 223 1165 227
rect 1188 226 1190 240
rect 1215 239 1216 243
rect 1220 242 1221 243
rect 1249 242 1251 256
rect 1254 251 1260 252
rect 1254 247 1255 251
rect 1259 247 1260 251
rect 1254 246 1260 247
rect 1310 251 1316 252
rect 1310 247 1311 251
rect 1315 247 1316 251
rect 1310 246 1316 247
rect 1366 251 1372 252
rect 1366 247 1367 251
rect 1371 247 1372 251
rect 1366 246 1372 247
rect 1414 251 1420 252
rect 1414 247 1415 251
rect 1419 247 1420 251
rect 1414 246 1420 247
rect 1462 251 1468 252
rect 1462 247 1463 251
rect 1467 247 1468 251
rect 1462 246 1468 247
rect 1518 251 1524 252
rect 1518 247 1519 251
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1574 251 1580 252
rect 1574 247 1575 251
rect 1579 247 1580 251
rect 1574 246 1580 247
rect 1622 251 1628 252
rect 1622 247 1623 251
rect 1627 247 1628 251
rect 1622 246 1628 247
rect 1662 249 1668 250
rect 1662 245 1663 249
rect 1667 245 1668 249
rect 1662 244 1668 245
rect 1271 243 1277 244
rect 1271 242 1272 243
rect 1220 240 1246 242
rect 1249 240 1272 242
rect 1220 239 1221 240
rect 1215 238 1221 239
rect 1198 234 1204 235
rect 1198 230 1199 234
rect 1203 230 1204 234
rect 1198 229 1204 230
rect 1215 227 1221 228
rect 1215 226 1216 227
rect 1188 224 1216 226
rect 1159 222 1165 223
rect 1215 223 1216 224
rect 1220 223 1221 227
rect 1244 226 1246 240
rect 1271 239 1272 240
rect 1276 239 1277 243
rect 1271 238 1277 239
rect 1322 243 1333 244
rect 1322 239 1323 243
rect 1327 239 1328 243
rect 1332 239 1333 243
rect 1383 243 1389 244
rect 1383 242 1384 243
rect 1322 238 1333 239
rect 1356 240 1384 242
rect 1254 234 1260 235
rect 1254 230 1255 234
rect 1259 230 1260 234
rect 1254 229 1260 230
rect 1310 234 1316 235
rect 1310 230 1311 234
rect 1315 230 1316 234
rect 1310 229 1316 230
rect 1271 227 1277 228
rect 1271 226 1272 227
rect 1244 224 1272 226
rect 1215 222 1221 223
rect 1271 223 1272 224
rect 1276 223 1277 227
rect 1271 222 1277 223
rect 1327 227 1333 228
rect 1327 223 1328 227
rect 1332 226 1333 227
rect 1356 226 1358 240
rect 1383 239 1384 240
rect 1388 239 1389 243
rect 1431 243 1437 244
rect 1431 242 1432 243
rect 1383 238 1389 239
rect 1408 240 1432 242
rect 1366 234 1372 235
rect 1366 230 1367 234
rect 1371 230 1372 234
rect 1366 229 1372 230
rect 1332 224 1358 226
rect 1383 227 1389 228
rect 1332 223 1333 224
rect 1327 222 1333 223
rect 1383 223 1384 227
rect 1388 226 1389 227
rect 1408 226 1410 240
rect 1431 239 1432 240
rect 1436 239 1437 243
rect 1431 238 1437 239
rect 1479 243 1485 244
rect 1479 239 1480 243
rect 1484 242 1485 243
rect 1535 243 1541 244
rect 1484 240 1530 242
rect 1484 239 1485 240
rect 1479 238 1485 239
rect 1414 234 1420 235
rect 1414 230 1415 234
rect 1419 230 1420 234
rect 1414 229 1420 230
rect 1462 234 1468 235
rect 1462 230 1463 234
rect 1467 230 1468 234
rect 1462 229 1468 230
rect 1518 234 1524 235
rect 1518 230 1519 234
rect 1523 230 1524 234
rect 1518 229 1524 230
rect 1388 224 1410 226
rect 1430 227 1437 228
rect 1388 223 1389 224
rect 1383 222 1389 223
rect 1430 223 1431 227
rect 1436 223 1437 227
rect 1430 222 1437 223
rect 1479 227 1488 228
rect 1479 223 1480 227
rect 1487 223 1488 227
rect 1528 226 1530 240
rect 1535 239 1536 243
rect 1540 242 1541 243
rect 1591 243 1597 244
rect 1540 240 1586 242
rect 1540 239 1541 240
rect 1535 238 1541 239
rect 1574 234 1580 235
rect 1574 230 1575 234
rect 1579 230 1580 234
rect 1574 229 1580 230
rect 1535 227 1541 228
rect 1535 226 1536 227
rect 1528 224 1536 226
rect 1479 222 1488 223
rect 1535 223 1536 224
rect 1540 223 1541 227
rect 1584 226 1586 240
rect 1591 239 1592 243
rect 1596 242 1597 243
rect 1634 243 1645 244
rect 1596 240 1618 242
rect 1596 239 1597 240
rect 1591 238 1597 239
rect 1591 227 1597 228
rect 1591 226 1592 227
rect 1584 224 1592 226
rect 1535 222 1541 223
rect 1591 223 1592 224
rect 1596 223 1597 227
rect 1616 226 1618 240
rect 1634 239 1635 243
rect 1639 239 1640 243
rect 1644 239 1645 243
rect 1634 238 1645 239
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1662 232 1668 233
rect 1662 228 1663 232
rect 1667 228 1668 232
rect 1639 227 1645 228
rect 1662 227 1668 228
rect 1639 226 1640 227
rect 1616 224 1640 226
rect 1591 222 1597 223
rect 1639 223 1640 224
rect 1644 223 1645 227
rect 1639 222 1645 223
rect 1230 219 1236 220
rect 1230 218 1231 219
rect 1012 216 1231 218
rect 438 214 444 215
rect 490 215 496 216
rect 399 211 405 212
rect 364 204 370 206
rect 390 207 397 208
rect 364 203 365 204
rect 390 203 391 207
rect 396 203 397 207
rect 399 207 400 211
rect 404 210 405 211
rect 439 211 445 212
rect 404 208 426 210
rect 404 207 405 208
rect 399 206 405 207
rect 424 206 426 208
rect 431 207 437 208
rect 431 206 432 207
rect 424 204 432 206
rect 431 203 432 204
rect 436 203 437 207
rect 439 207 440 211
rect 444 210 445 211
rect 490 211 491 215
rect 495 214 496 215
rect 1230 215 1231 216
rect 1235 215 1236 219
rect 1634 219 1640 220
rect 1634 218 1635 219
rect 1230 214 1236 215
rect 1544 216 1635 218
rect 495 212 626 214
rect 495 211 496 212
rect 490 210 496 211
rect 444 208 482 210
rect 444 207 445 208
rect 439 206 445 207
rect 480 206 482 208
rect 487 207 493 208
rect 487 206 488 207
rect 480 204 488 206
rect 487 203 488 204
rect 492 203 493 207
rect 551 207 557 208
rect 551 203 552 207
rect 556 206 557 207
rect 574 207 580 208
rect 574 206 575 207
rect 556 204 575 206
rect 556 203 557 204
rect 342 202 348 203
rect 359 202 365 203
rect 374 202 380 203
rect 390 202 397 203
rect 414 202 420 203
rect 431 202 437 203
rect 470 202 476 203
rect 487 202 493 203
rect 534 202 540 203
rect 551 202 557 203
rect 574 203 575 204
rect 579 203 580 207
rect 624 206 626 212
rect 639 211 645 212
rect 631 207 637 208
rect 631 206 632 207
rect 624 204 632 206
rect 631 203 632 204
rect 636 203 637 207
rect 639 207 640 211
rect 644 210 645 211
rect 719 211 725 212
rect 644 208 706 210
rect 644 207 645 208
rect 639 206 645 207
rect 704 206 706 208
rect 711 207 717 208
rect 711 206 712 207
rect 704 204 712 206
rect 711 203 712 204
rect 716 203 717 207
rect 719 207 720 211
rect 724 210 725 211
rect 879 211 885 212
rect 724 208 786 210
rect 724 207 725 208
rect 719 206 725 207
rect 784 206 786 208
rect 791 207 797 208
rect 791 206 792 207
rect 784 204 792 206
rect 791 203 792 204
rect 796 203 797 207
rect 870 207 877 208
rect 870 203 871 207
rect 876 203 877 207
rect 879 207 880 211
rect 884 210 885 211
rect 951 211 957 212
rect 884 208 938 210
rect 884 207 885 208
rect 879 206 885 207
rect 936 206 938 208
rect 943 207 949 208
rect 943 206 944 207
rect 936 204 944 206
rect 943 203 944 204
rect 948 203 949 207
rect 951 207 952 211
rect 956 210 957 211
rect 1023 211 1029 212
rect 956 208 1010 210
rect 956 207 957 208
rect 951 206 957 207
rect 1008 206 1010 208
rect 1015 207 1021 208
rect 1015 206 1016 207
rect 1008 204 1016 206
rect 1015 203 1016 204
rect 1020 203 1021 207
rect 1023 207 1024 211
rect 1028 210 1029 211
rect 1095 211 1101 212
rect 1028 208 1082 210
rect 1028 207 1029 208
rect 1023 206 1029 207
rect 1080 206 1082 208
rect 1087 207 1093 208
rect 1087 206 1088 207
rect 1080 204 1088 206
rect 1087 203 1088 204
rect 1092 203 1093 207
rect 1095 207 1096 211
rect 1100 210 1101 211
rect 1167 211 1173 212
rect 1100 208 1161 210
rect 1100 207 1101 208
rect 1095 206 1101 207
rect 1159 207 1165 208
rect 1159 203 1160 207
rect 1164 203 1165 207
rect 1167 207 1168 211
rect 1172 210 1173 211
rect 1330 211 1336 212
rect 1172 208 1226 210
rect 1172 207 1173 208
rect 1167 206 1173 207
rect 1224 206 1226 208
rect 1231 207 1237 208
rect 1231 206 1232 207
rect 1224 204 1232 206
rect 1231 203 1232 204
rect 1236 203 1237 207
rect 1303 207 1309 208
rect 1303 203 1304 207
rect 1308 206 1309 207
rect 1322 207 1328 208
rect 1322 206 1323 207
rect 1308 204 1323 206
rect 1308 203 1309 204
rect 574 202 580 203
rect 614 202 620 203
rect 631 202 637 203
rect 694 202 700 203
rect 711 202 717 203
rect 774 202 780 203
rect 791 202 797 203
rect 854 202 860 203
rect 870 202 877 203
rect 926 202 932 203
rect 943 202 949 203
rect 998 202 1004 203
rect 1015 202 1021 203
rect 1070 202 1076 203
rect 1087 202 1093 203
rect 1142 202 1148 203
rect 1159 202 1165 203
rect 1214 202 1220 203
rect 1231 202 1237 203
rect 1286 202 1292 203
rect 1303 202 1309 203
rect 1322 203 1323 204
rect 1327 203 1328 207
rect 1330 207 1331 211
rect 1335 210 1336 211
rect 1454 211 1460 212
rect 1335 208 1362 210
rect 1335 207 1336 208
rect 1330 206 1336 207
rect 1360 206 1362 208
rect 1367 207 1373 208
rect 1367 206 1368 207
rect 1360 204 1368 206
rect 1367 203 1368 204
rect 1372 203 1373 207
rect 1431 207 1440 208
rect 1431 203 1432 207
rect 1439 203 1440 207
rect 1454 207 1455 211
rect 1459 210 1460 211
rect 1459 208 1482 210
rect 1544 208 1546 216
rect 1634 215 1635 216
rect 1639 215 1640 219
rect 1634 214 1640 215
rect 1551 211 1557 212
rect 1459 207 1460 208
rect 1454 206 1460 207
rect 1480 206 1482 208
rect 1487 207 1493 208
rect 1487 206 1488 207
rect 1480 204 1488 206
rect 1487 203 1488 204
rect 1492 203 1493 207
rect 1543 207 1549 208
rect 1543 203 1544 207
rect 1548 203 1549 207
rect 1551 207 1552 211
rect 1556 210 1557 211
rect 1607 211 1613 212
rect 1556 208 1603 210
rect 1556 207 1557 208
rect 1551 206 1557 207
rect 1599 207 1605 208
rect 1599 203 1600 207
rect 1604 203 1605 207
rect 1607 207 1608 211
rect 1612 210 1613 211
rect 1612 208 1643 210
rect 1612 207 1613 208
rect 1607 206 1613 207
rect 1639 207 1645 208
rect 1639 203 1640 207
rect 1644 203 1645 207
rect 1322 202 1328 203
rect 1350 202 1356 203
rect 1367 202 1373 203
rect 1414 202 1420 203
rect 1431 202 1440 203
rect 1470 202 1476 203
rect 1487 202 1493 203
rect 1526 202 1532 203
rect 1543 202 1549 203
rect 1582 202 1588 203
rect 1599 202 1605 203
rect 1622 202 1628 203
rect 1639 202 1645 203
rect 1662 204 1668 205
rect 342 198 343 202
rect 347 198 348 202
rect 342 197 348 198
rect 374 198 375 202
rect 379 198 380 202
rect 374 197 380 198
rect 414 198 415 202
rect 419 198 420 202
rect 414 197 420 198
rect 470 198 471 202
rect 475 198 476 202
rect 470 197 476 198
rect 534 198 535 202
rect 539 198 540 202
rect 534 197 540 198
rect 614 198 615 202
rect 619 198 620 202
rect 614 197 620 198
rect 694 198 695 202
rect 699 198 700 202
rect 694 197 700 198
rect 774 198 775 202
rect 779 198 780 202
rect 774 197 780 198
rect 854 198 855 202
rect 859 198 860 202
rect 854 197 860 198
rect 926 198 927 202
rect 931 198 932 202
rect 926 197 932 198
rect 998 198 999 202
rect 1003 198 1004 202
rect 998 197 1004 198
rect 1070 198 1071 202
rect 1075 198 1076 202
rect 1070 197 1076 198
rect 1142 198 1143 202
rect 1147 198 1148 202
rect 1142 197 1148 198
rect 1214 198 1215 202
rect 1219 198 1220 202
rect 1214 197 1220 198
rect 1286 198 1287 202
rect 1291 198 1292 202
rect 1286 197 1292 198
rect 1350 198 1351 202
rect 1355 198 1356 202
rect 1350 197 1356 198
rect 1414 198 1415 202
rect 1419 198 1420 202
rect 1414 197 1420 198
rect 1470 198 1471 202
rect 1475 198 1476 202
rect 1470 197 1476 198
rect 1526 198 1527 202
rect 1531 198 1532 202
rect 1526 197 1532 198
rect 1582 198 1583 202
rect 1587 198 1588 202
rect 1582 197 1588 198
rect 1622 198 1623 202
rect 1627 198 1628 202
rect 1662 200 1663 204
rect 1667 200 1668 204
rect 1662 199 1668 200
rect 1622 197 1628 198
rect 336 192 342 194
rect 319 191 325 192
rect 319 190 320 191
rect 312 188 320 190
rect 294 186 300 187
rect 319 187 320 188
rect 324 187 325 191
rect 340 190 354 192
rect 359 191 365 192
rect 359 190 360 191
rect 352 188 360 190
rect 319 186 325 187
rect 359 187 360 188
rect 364 187 365 191
rect 359 186 365 187
rect 391 191 397 192
rect 391 187 392 191
rect 396 190 397 191
rect 399 191 405 192
rect 399 190 400 191
rect 396 188 400 190
rect 396 187 397 188
rect 391 186 397 187
rect 399 187 400 188
rect 404 187 405 191
rect 399 186 405 187
rect 431 191 437 192
rect 431 187 432 191
rect 436 190 437 191
rect 439 191 445 192
rect 439 190 440 191
rect 436 188 440 190
rect 436 187 437 188
rect 431 186 437 187
rect 439 187 440 188
rect 444 187 445 191
rect 439 186 445 187
rect 487 191 496 192
rect 487 187 488 191
rect 495 187 496 191
rect 551 191 557 192
rect 551 190 552 191
rect 487 186 496 187
rect 544 188 552 190
rect 110 182 116 183
rect 134 185 140 186
rect 134 181 135 185
rect 139 181 140 185
rect 134 180 140 181
rect 166 185 172 186
rect 166 181 167 185
rect 171 181 172 185
rect 166 180 172 181
rect 206 185 212 186
rect 206 181 207 185
rect 211 181 212 185
rect 206 180 212 181
rect 254 185 260 186
rect 254 181 255 185
rect 259 181 260 185
rect 254 180 260 181
rect 302 185 308 186
rect 302 181 303 185
rect 307 181 308 185
rect 302 180 308 181
rect 342 185 348 186
rect 342 181 343 185
rect 347 181 348 185
rect 342 180 348 181
rect 374 185 380 186
rect 374 181 375 185
rect 379 181 380 185
rect 374 180 380 181
rect 414 185 420 186
rect 414 181 415 185
rect 419 181 420 185
rect 414 180 420 181
rect 470 185 476 186
rect 470 181 471 185
rect 475 181 476 185
rect 470 180 476 181
rect 534 185 540 186
rect 534 181 535 185
rect 539 181 540 185
rect 534 180 540 181
rect 390 179 396 180
rect 390 175 391 179
rect 395 178 396 179
rect 544 178 546 188
rect 551 187 552 188
rect 556 187 557 191
rect 551 186 557 187
rect 631 191 637 192
rect 631 187 632 191
rect 636 190 637 191
rect 639 191 645 192
rect 639 190 640 191
rect 636 188 640 190
rect 636 187 637 188
rect 631 186 637 187
rect 639 187 640 188
rect 644 187 645 191
rect 639 186 645 187
rect 711 191 717 192
rect 711 187 712 191
rect 716 190 717 191
rect 719 191 725 192
rect 719 190 720 191
rect 716 188 720 190
rect 716 187 717 188
rect 711 186 717 187
rect 719 187 720 188
rect 724 187 725 191
rect 719 186 725 187
rect 786 191 797 192
rect 786 187 787 191
rect 791 187 792 191
rect 796 187 797 191
rect 786 186 797 187
rect 871 191 877 192
rect 871 187 872 191
rect 876 190 877 191
rect 879 191 885 192
rect 879 190 880 191
rect 876 188 880 190
rect 876 187 877 188
rect 871 186 877 187
rect 879 187 880 188
rect 884 187 885 191
rect 879 186 885 187
rect 943 191 949 192
rect 943 187 944 191
rect 948 190 949 191
rect 951 191 957 192
rect 951 190 952 191
rect 948 188 952 190
rect 948 187 949 188
rect 943 186 949 187
rect 951 187 952 188
rect 956 187 957 191
rect 951 186 957 187
rect 1015 191 1021 192
rect 1015 187 1016 191
rect 1020 190 1021 191
rect 1023 191 1029 192
rect 1023 190 1024 191
rect 1020 188 1024 190
rect 1020 187 1021 188
rect 1015 186 1021 187
rect 1023 187 1024 188
rect 1028 187 1029 191
rect 1023 186 1029 187
rect 1087 191 1093 192
rect 1087 187 1088 191
rect 1092 190 1093 191
rect 1095 191 1101 192
rect 1095 190 1096 191
rect 1092 188 1096 190
rect 1092 187 1093 188
rect 1087 186 1093 187
rect 1095 187 1096 188
rect 1100 187 1101 191
rect 1095 186 1101 187
rect 1159 191 1165 192
rect 1159 187 1160 191
rect 1164 190 1165 191
rect 1167 191 1173 192
rect 1167 190 1168 191
rect 1164 188 1168 190
rect 1164 187 1165 188
rect 1159 186 1165 187
rect 1167 187 1168 188
rect 1172 187 1173 191
rect 1167 186 1173 187
rect 1230 191 1237 192
rect 1230 187 1231 191
rect 1236 187 1237 191
rect 1230 186 1237 187
rect 1303 191 1309 192
rect 1303 187 1304 191
rect 1308 190 1309 191
rect 1330 191 1336 192
rect 1330 190 1331 191
rect 1308 188 1331 190
rect 1308 187 1309 188
rect 1303 186 1309 187
rect 1330 187 1331 188
rect 1335 187 1336 191
rect 1330 186 1336 187
rect 1366 191 1373 192
rect 1366 187 1367 191
rect 1372 187 1373 191
rect 1366 186 1373 187
rect 1431 191 1437 192
rect 1431 187 1432 191
rect 1436 190 1437 191
rect 1454 191 1460 192
rect 1454 190 1455 191
rect 1436 188 1455 190
rect 1436 187 1437 188
rect 1431 186 1437 187
rect 1454 187 1455 188
rect 1459 187 1460 191
rect 1454 186 1460 187
rect 1482 191 1493 192
rect 1482 187 1483 191
rect 1487 187 1488 191
rect 1492 187 1493 191
rect 1482 186 1493 187
rect 1543 191 1549 192
rect 1543 187 1544 191
rect 1548 190 1549 191
rect 1551 191 1557 192
rect 1551 190 1552 191
rect 1548 188 1552 190
rect 1548 187 1549 188
rect 1543 186 1549 187
rect 1551 187 1552 188
rect 1556 187 1557 191
rect 1551 186 1557 187
rect 1599 191 1605 192
rect 1599 187 1600 191
rect 1604 190 1605 191
rect 1607 191 1613 192
rect 1607 190 1608 191
rect 1604 188 1608 190
rect 1604 187 1605 188
rect 1599 186 1605 187
rect 1607 187 1608 188
rect 1612 187 1613 191
rect 1607 186 1613 187
rect 1638 191 1645 192
rect 1638 187 1639 191
rect 1644 187 1645 191
rect 1638 186 1645 187
rect 1662 187 1668 188
rect 614 185 620 186
rect 614 181 615 185
rect 619 181 620 185
rect 614 180 620 181
rect 694 185 700 186
rect 694 181 695 185
rect 699 181 700 185
rect 694 180 700 181
rect 774 185 780 186
rect 774 181 775 185
rect 779 181 780 185
rect 774 180 780 181
rect 854 185 860 186
rect 854 181 855 185
rect 859 181 860 185
rect 854 180 860 181
rect 926 185 932 186
rect 926 181 927 185
rect 931 181 932 185
rect 926 180 932 181
rect 998 185 1004 186
rect 998 181 999 185
rect 1003 181 1004 185
rect 998 180 1004 181
rect 1070 185 1076 186
rect 1070 181 1071 185
rect 1075 181 1076 185
rect 1070 180 1076 181
rect 1142 185 1148 186
rect 1142 181 1143 185
rect 1147 181 1148 185
rect 1142 180 1148 181
rect 1214 185 1220 186
rect 1214 181 1215 185
rect 1219 181 1220 185
rect 1214 180 1220 181
rect 1286 185 1292 186
rect 1286 181 1287 185
rect 1291 181 1292 185
rect 1286 180 1292 181
rect 1350 185 1356 186
rect 1350 181 1351 185
rect 1355 181 1356 185
rect 1350 180 1356 181
rect 1414 185 1420 186
rect 1414 181 1415 185
rect 1419 181 1420 185
rect 1414 180 1420 181
rect 1470 185 1476 186
rect 1470 181 1471 185
rect 1475 181 1476 185
rect 1470 180 1476 181
rect 1526 185 1532 186
rect 1526 181 1527 185
rect 1531 181 1532 185
rect 1526 180 1532 181
rect 1582 185 1588 186
rect 1582 181 1583 185
rect 1587 181 1588 185
rect 1582 180 1588 181
rect 1622 185 1628 186
rect 1622 181 1623 185
rect 1627 181 1628 185
rect 1662 183 1663 187
rect 1667 183 1668 187
rect 1662 182 1668 183
rect 1622 180 1628 181
rect 395 176 546 178
rect 870 179 876 180
rect 395 175 396 176
rect 390 174 396 175
rect 870 175 871 179
rect 875 178 876 179
rect 875 176 1161 178
rect 875 175 876 176
rect 870 174 876 175
rect 134 171 140 172
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 134 167 135 171
rect 139 167 140 171
rect 134 166 140 167
rect 174 171 180 172
rect 174 167 175 171
rect 179 167 180 171
rect 174 166 180 167
rect 230 171 236 172
rect 230 167 231 171
rect 235 167 236 171
rect 230 166 236 167
rect 286 171 292 172
rect 286 167 287 171
rect 291 167 292 171
rect 286 166 292 167
rect 342 171 348 172
rect 342 167 343 171
rect 347 167 348 171
rect 342 166 348 167
rect 398 171 404 172
rect 398 167 399 171
rect 403 167 404 171
rect 398 166 404 167
rect 454 171 460 172
rect 454 167 455 171
rect 459 167 460 171
rect 454 166 460 167
rect 510 171 516 172
rect 510 167 511 171
rect 515 167 516 171
rect 510 166 516 167
rect 574 171 580 172
rect 574 167 575 171
rect 579 167 580 171
rect 574 166 580 167
rect 638 171 644 172
rect 638 167 639 171
rect 643 167 644 171
rect 638 166 644 167
rect 702 171 708 172
rect 702 167 703 171
rect 707 167 708 171
rect 702 166 708 167
rect 766 171 772 172
rect 766 167 767 171
rect 771 167 772 171
rect 766 166 772 167
rect 830 171 836 172
rect 830 167 831 171
rect 835 167 836 171
rect 830 166 836 167
rect 894 171 900 172
rect 894 167 895 171
rect 899 167 900 171
rect 894 166 900 167
rect 950 171 956 172
rect 950 167 951 171
rect 955 167 956 171
rect 950 166 956 167
rect 1014 171 1020 172
rect 1014 167 1015 171
rect 1019 167 1020 171
rect 1014 166 1020 167
rect 1078 171 1084 172
rect 1078 167 1079 171
rect 1083 167 1084 171
rect 1078 166 1084 167
rect 1142 171 1148 172
rect 1142 167 1143 171
rect 1147 167 1148 171
rect 1142 166 1148 167
rect 110 164 116 165
rect 1159 164 1161 176
rect 1206 171 1212 172
rect 1206 167 1207 171
rect 1211 167 1212 171
rect 1206 166 1212 167
rect 1278 171 1284 172
rect 1278 167 1279 171
rect 1283 167 1284 171
rect 1278 166 1284 167
rect 1350 171 1356 172
rect 1350 167 1351 171
rect 1355 167 1356 171
rect 1350 166 1356 167
rect 1422 171 1428 172
rect 1422 167 1423 171
rect 1427 167 1428 171
rect 1422 166 1428 167
rect 1494 171 1500 172
rect 1494 167 1495 171
rect 1499 167 1500 171
rect 1494 166 1500 167
rect 1566 171 1572 172
rect 1566 167 1567 171
rect 1571 167 1572 171
rect 1566 166 1572 167
rect 1622 171 1628 172
rect 1622 167 1623 171
rect 1627 167 1628 171
rect 1622 166 1628 167
rect 1662 169 1668 170
rect 1662 165 1663 169
rect 1667 165 1668 169
rect 1662 164 1668 165
rect 151 163 157 164
rect 151 159 152 163
rect 156 162 157 163
rect 191 163 197 164
rect 156 160 186 162
rect 156 159 157 160
rect 151 158 157 159
rect 134 154 140 155
rect 110 152 116 153
rect 110 148 111 152
rect 115 148 116 152
rect 134 150 135 154
rect 139 150 140 154
rect 134 149 140 150
rect 174 154 180 155
rect 174 150 175 154
rect 179 150 180 154
rect 174 149 180 150
rect 110 147 116 148
rect 150 147 157 148
rect 150 143 151 147
rect 156 143 157 147
rect 184 146 186 160
rect 191 159 192 163
rect 196 162 197 163
rect 246 163 253 164
rect 196 160 222 162
rect 196 159 197 160
rect 191 158 197 159
rect 191 147 197 148
rect 191 146 192 147
rect 184 144 192 146
rect 150 142 157 143
rect 191 143 192 144
rect 196 143 197 147
rect 220 146 222 160
rect 246 159 247 163
rect 252 159 253 163
rect 246 158 253 159
rect 303 163 309 164
rect 303 159 304 163
rect 308 162 309 163
rect 359 163 365 164
rect 308 160 321 162
rect 308 159 309 160
rect 303 158 309 159
rect 230 154 236 155
rect 230 150 231 154
rect 235 150 236 154
rect 230 149 236 150
rect 286 154 292 155
rect 286 150 287 154
rect 291 150 292 154
rect 286 149 292 150
rect 247 147 253 148
rect 247 146 248 147
rect 220 144 248 146
rect 191 142 197 143
rect 247 143 248 144
rect 252 143 253 147
rect 247 142 253 143
rect 294 147 300 148
rect 294 143 295 147
rect 299 146 300 147
rect 303 147 309 148
rect 303 146 304 147
rect 299 144 304 146
rect 299 143 300 144
rect 294 142 300 143
rect 303 143 304 144
rect 308 143 309 147
rect 319 146 321 160
rect 359 159 360 163
rect 364 162 365 163
rect 415 163 421 164
rect 364 160 390 162
rect 364 159 365 160
rect 359 158 365 159
rect 342 154 348 155
rect 342 150 343 154
rect 347 150 348 154
rect 342 149 348 150
rect 359 147 365 148
rect 359 146 360 147
rect 319 144 360 146
rect 303 142 309 143
rect 359 143 360 144
rect 364 143 365 147
rect 388 146 390 160
rect 415 159 416 163
rect 420 162 421 163
rect 438 163 444 164
rect 438 162 439 163
rect 420 160 439 162
rect 420 159 421 160
rect 415 158 421 159
rect 438 159 439 160
rect 443 159 444 163
rect 438 158 444 159
rect 471 163 477 164
rect 471 159 472 163
rect 476 162 477 163
rect 527 163 533 164
rect 476 160 522 162
rect 476 159 477 160
rect 471 158 477 159
rect 398 154 404 155
rect 398 150 399 154
rect 403 150 404 154
rect 398 149 404 150
rect 454 154 460 155
rect 454 150 455 154
rect 459 150 460 154
rect 454 149 460 150
rect 510 154 516 155
rect 510 150 511 154
rect 515 150 516 154
rect 510 149 516 150
rect 415 147 421 148
rect 415 146 416 147
rect 388 144 416 146
rect 359 142 365 143
rect 415 143 416 144
rect 420 143 421 147
rect 415 142 421 143
rect 471 147 477 148
rect 471 143 472 147
rect 476 143 477 147
rect 520 146 522 160
rect 527 159 528 163
rect 532 162 533 163
rect 591 163 597 164
rect 532 160 562 162
rect 532 159 533 160
rect 527 158 533 159
rect 527 147 533 148
rect 527 146 528 147
rect 520 144 528 146
rect 471 142 477 143
rect 527 143 528 144
rect 532 143 533 147
rect 560 146 562 160
rect 591 159 592 163
rect 596 162 597 163
rect 655 163 661 164
rect 596 160 650 162
rect 596 159 597 160
rect 591 158 597 159
rect 574 154 580 155
rect 574 150 575 154
rect 579 150 580 154
rect 574 149 580 150
rect 638 154 644 155
rect 638 150 639 154
rect 643 150 644 154
rect 638 149 644 150
rect 591 147 597 148
rect 591 146 592 147
rect 560 144 592 146
rect 527 142 533 143
rect 591 143 592 144
rect 596 143 597 147
rect 648 146 650 160
rect 655 159 656 163
rect 660 162 661 163
rect 719 163 725 164
rect 660 160 714 162
rect 660 159 661 160
rect 655 158 661 159
rect 702 154 708 155
rect 702 150 703 154
rect 707 150 708 154
rect 702 149 708 150
rect 655 147 661 148
rect 655 146 656 147
rect 648 144 656 146
rect 591 142 597 143
rect 655 143 656 144
rect 660 143 661 147
rect 712 146 714 160
rect 719 159 720 163
rect 724 162 725 163
rect 758 163 764 164
rect 724 160 754 162
rect 724 159 725 160
rect 719 158 725 159
rect 719 147 725 148
rect 719 146 720 147
rect 712 144 720 146
rect 655 142 661 143
rect 719 143 720 144
rect 724 143 725 147
rect 752 146 754 160
rect 758 159 759 163
rect 763 162 764 163
rect 783 163 789 164
rect 783 162 784 163
rect 763 160 784 162
rect 763 159 764 160
rect 758 158 764 159
rect 783 159 784 160
rect 788 159 789 163
rect 783 158 789 159
rect 847 163 853 164
rect 847 159 848 163
rect 852 162 853 163
rect 911 163 917 164
rect 852 160 882 162
rect 852 159 853 160
rect 847 158 853 159
rect 766 154 772 155
rect 766 150 767 154
rect 771 150 772 154
rect 766 149 772 150
rect 830 154 836 155
rect 830 150 831 154
rect 835 150 836 154
rect 830 149 836 150
rect 783 147 789 148
rect 783 146 784 147
rect 752 144 784 146
rect 719 142 725 143
rect 783 143 784 144
rect 788 143 789 147
rect 783 142 789 143
rect 847 147 853 148
rect 847 143 848 147
rect 852 146 853 147
rect 880 146 882 160
rect 911 159 912 163
rect 916 162 917 163
rect 967 163 973 164
rect 916 160 942 162
rect 916 159 917 160
rect 911 158 917 159
rect 894 154 900 155
rect 894 150 895 154
rect 899 150 900 154
rect 894 149 900 150
rect 911 147 917 148
rect 911 146 912 147
rect 852 144 878 146
rect 880 144 912 146
rect 852 143 853 144
rect 847 142 853 143
rect 473 138 475 142
rect 786 139 792 140
rect 786 138 787 139
rect 473 136 787 138
rect 786 135 787 136
rect 791 135 792 139
rect 876 138 878 144
rect 911 143 912 144
rect 916 143 917 147
rect 940 146 942 160
rect 967 159 968 163
rect 972 162 973 163
rect 1031 163 1037 164
rect 972 160 1026 162
rect 972 159 973 160
rect 967 158 973 159
rect 950 154 956 155
rect 950 150 951 154
rect 955 150 956 154
rect 950 149 956 150
rect 1014 154 1020 155
rect 1014 150 1015 154
rect 1019 150 1020 154
rect 1014 149 1020 150
rect 967 147 973 148
rect 967 146 968 147
rect 940 144 968 146
rect 911 142 917 143
rect 967 143 968 144
rect 972 143 973 147
rect 1024 146 1026 160
rect 1031 159 1032 163
rect 1036 162 1037 163
rect 1095 163 1101 164
rect 1036 160 1066 162
rect 1036 159 1037 160
rect 1031 158 1037 159
rect 1031 147 1037 148
rect 1031 146 1032 147
rect 1024 144 1032 146
rect 967 142 973 143
rect 1031 143 1032 144
rect 1036 143 1037 147
rect 1064 146 1066 160
rect 1095 159 1096 163
rect 1100 162 1101 163
rect 1159 163 1165 164
rect 1100 160 1130 162
rect 1100 159 1101 160
rect 1095 158 1101 159
rect 1078 154 1084 155
rect 1078 150 1079 154
rect 1083 150 1084 154
rect 1078 149 1084 150
rect 1095 147 1101 148
rect 1095 146 1096 147
rect 1064 144 1096 146
rect 1031 142 1037 143
rect 1095 143 1096 144
rect 1100 143 1101 147
rect 1128 146 1130 160
rect 1159 159 1160 163
rect 1164 159 1165 163
rect 1159 158 1165 159
rect 1198 163 1204 164
rect 1198 159 1199 163
rect 1203 162 1204 163
rect 1223 163 1229 164
rect 1223 162 1224 163
rect 1203 160 1224 162
rect 1203 159 1204 160
rect 1198 158 1204 159
rect 1223 159 1224 160
rect 1228 159 1229 163
rect 1295 163 1301 164
rect 1295 162 1296 163
rect 1223 158 1229 159
rect 1260 160 1296 162
rect 1142 154 1148 155
rect 1142 150 1143 154
rect 1147 150 1148 154
rect 1142 149 1148 150
rect 1206 154 1212 155
rect 1206 150 1207 154
rect 1211 150 1212 154
rect 1206 149 1212 150
rect 1159 147 1165 148
rect 1159 146 1160 147
rect 1128 144 1160 146
rect 1095 142 1101 143
rect 1159 143 1160 144
rect 1164 143 1165 147
rect 1159 142 1165 143
rect 1223 147 1229 148
rect 1223 143 1224 147
rect 1228 146 1229 147
rect 1260 146 1262 160
rect 1295 159 1296 160
rect 1300 159 1301 163
rect 1367 163 1373 164
rect 1367 162 1368 163
rect 1295 158 1301 159
rect 1332 160 1368 162
rect 1278 154 1284 155
rect 1278 150 1279 154
rect 1283 150 1284 154
rect 1278 149 1284 150
rect 1228 144 1262 146
rect 1295 147 1301 148
rect 1228 143 1229 144
rect 1223 142 1229 143
rect 1295 143 1296 147
rect 1300 146 1301 147
rect 1332 146 1334 160
rect 1367 159 1368 160
rect 1372 159 1373 163
rect 1367 158 1373 159
rect 1434 163 1445 164
rect 1434 159 1435 163
rect 1439 159 1440 163
rect 1444 159 1445 163
rect 1511 163 1517 164
rect 1511 162 1512 163
rect 1434 158 1445 159
rect 1480 160 1512 162
rect 1350 154 1356 155
rect 1350 150 1351 154
rect 1355 150 1356 154
rect 1350 149 1356 150
rect 1422 154 1428 155
rect 1422 150 1423 154
rect 1427 150 1428 154
rect 1422 149 1428 150
rect 1300 144 1334 146
rect 1366 147 1373 148
rect 1300 143 1301 144
rect 1295 142 1301 143
rect 1366 143 1367 147
rect 1372 143 1373 147
rect 1366 142 1373 143
rect 1439 147 1445 148
rect 1439 143 1440 147
rect 1444 146 1445 147
rect 1480 146 1482 160
rect 1511 159 1512 160
rect 1516 159 1517 163
rect 1583 163 1589 164
rect 1583 162 1584 163
rect 1511 158 1517 159
rect 1548 160 1584 162
rect 1494 154 1500 155
rect 1494 150 1495 154
rect 1499 150 1500 154
rect 1494 149 1500 150
rect 1444 144 1482 146
rect 1511 147 1517 148
rect 1444 143 1445 144
rect 1439 142 1445 143
rect 1511 143 1512 147
rect 1516 146 1517 147
rect 1548 146 1550 160
rect 1583 159 1584 160
rect 1588 159 1589 163
rect 1583 158 1589 159
rect 1639 163 1645 164
rect 1639 159 1640 163
rect 1644 162 1645 163
rect 1647 163 1653 164
rect 1647 162 1648 163
rect 1644 160 1648 162
rect 1644 159 1645 160
rect 1639 158 1645 159
rect 1647 159 1648 160
rect 1652 159 1653 163
rect 1647 158 1653 159
rect 1566 154 1572 155
rect 1566 150 1567 154
rect 1571 150 1572 154
rect 1566 149 1572 150
rect 1622 154 1628 155
rect 1622 150 1623 154
rect 1627 150 1628 154
rect 1622 149 1628 150
rect 1662 152 1668 153
rect 1662 148 1663 152
rect 1667 148 1668 152
rect 1516 144 1550 146
rect 1574 147 1580 148
rect 1516 143 1517 144
rect 1511 142 1517 143
rect 1574 143 1575 147
rect 1579 146 1580 147
rect 1583 147 1589 148
rect 1583 146 1584 147
rect 1579 144 1584 146
rect 1579 143 1580 144
rect 1574 142 1580 143
rect 1583 143 1584 144
rect 1588 143 1589 147
rect 1583 142 1589 143
rect 1638 147 1645 148
rect 1662 147 1668 148
rect 1638 143 1639 147
rect 1644 143 1645 147
rect 1638 142 1645 143
rect 1158 139 1164 140
rect 1158 138 1159 139
rect 876 136 1159 138
rect 786 134 792 135
rect 1158 135 1159 136
rect 1163 135 1164 139
rect 1158 134 1164 135
rect 480 132 762 134
rect 478 131 484 132
rect 478 127 479 131
rect 483 127 484 131
rect 478 126 484 127
rect 758 131 764 132
rect 758 127 759 131
rect 763 127 764 131
rect 758 126 764 127
rect 487 115 493 116
rect 153 112 178 114
rect 185 112 210 114
rect 225 112 242 114
rect 256 112 274 114
rect 281 112 306 114
rect 319 112 338 114
rect 345 112 370 114
rect 384 112 402 114
rect 409 112 434 114
rect 151 111 157 112
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 151 107 152 111
rect 156 107 157 111
rect 110 103 116 104
rect 134 106 140 107
rect 151 106 157 107
rect 166 106 172 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 150 95 157 96
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 150 91 151 95
rect 156 91 157 95
rect 176 94 178 112
rect 183 111 189 112
rect 183 107 184 111
rect 188 107 189 111
rect 183 106 189 107
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 183 95 189 96
rect 183 94 184 95
rect 176 92 184 94
rect 150 90 157 91
rect 183 91 184 92
rect 188 91 189 95
rect 208 94 210 112
rect 215 111 221 112
rect 215 107 216 111
rect 220 110 221 111
rect 225 110 227 112
rect 220 108 227 110
rect 220 107 221 108
rect 215 106 221 107
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 215 95 221 96
rect 215 94 216 95
rect 208 92 216 94
rect 183 90 189 91
rect 215 91 216 92
rect 220 91 221 95
rect 240 94 242 112
rect 247 111 253 112
rect 247 107 248 111
rect 252 110 253 111
rect 256 110 258 112
rect 252 108 258 110
rect 252 107 253 108
rect 247 106 253 107
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 247 95 253 96
rect 247 94 248 95
rect 240 92 248 94
rect 215 90 221 91
rect 247 91 248 92
rect 252 91 253 95
rect 272 94 274 112
rect 279 111 285 112
rect 279 107 280 111
rect 284 107 285 111
rect 279 106 285 107
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 279 95 285 96
rect 279 94 280 95
rect 272 92 280 94
rect 247 90 253 91
rect 279 91 280 92
rect 284 91 285 95
rect 304 94 306 112
rect 311 111 317 112
rect 311 107 312 111
rect 316 110 317 111
rect 319 110 321 112
rect 316 108 321 110
rect 316 107 317 108
rect 311 106 317 107
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 336 102 338 112
rect 343 111 349 112
rect 343 107 344 111
rect 348 107 349 111
rect 343 106 349 107
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 336 100 347 102
rect 358 101 364 102
rect 345 96 347 100
rect 311 95 317 96
rect 311 94 312 95
rect 304 92 312 94
rect 279 90 285 91
rect 311 91 312 92
rect 316 91 317 95
rect 311 90 317 91
rect 343 95 349 96
rect 343 91 344 95
rect 348 91 349 95
rect 368 94 370 112
rect 375 111 381 112
rect 375 107 376 111
rect 380 110 381 111
rect 384 110 386 112
rect 380 108 386 110
rect 380 107 381 108
rect 375 106 381 107
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 400 98 402 112
rect 407 111 413 112
rect 407 107 408 111
rect 412 107 413 111
rect 407 106 413 107
rect 422 106 428 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 400 96 411 98
rect 375 95 381 96
rect 375 94 376 95
rect 368 92 376 94
rect 343 90 349 91
rect 375 91 376 92
rect 380 91 381 95
rect 375 90 381 91
rect 407 95 413 96
rect 407 91 408 95
rect 412 91 413 95
rect 432 94 434 112
rect 438 111 445 112
rect 438 107 439 111
rect 444 107 445 111
rect 478 111 485 112
rect 478 107 479 111
rect 484 107 485 111
rect 487 111 488 115
rect 492 114 493 115
rect 527 115 533 116
rect 492 112 514 114
rect 492 111 493 112
rect 487 110 493 111
rect 512 110 514 112
rect 519 111 525 112
rect 519 110 520 111
rect 512 108 520 110
rect 519 107 520 108
rect 524 107 525 111
rect 527 111 528 115
rect 532 114 533 115
rect 919 115 925 116
rect 532 112 554 114
rect 568 112 595 114
rect 632 112 659 114
rect 532 111 533 112
rect 527 110 533 111
rect 552 110 554 112
rect 559 111 565 112
rect 559 110 560 111
rect 552 108 560 110
rect 559 107 560 108
rect 564 107 565 111
rect 438 106 445 107
rect 462 106 468 107
rect 478 106 485 107
rect 502 106 508 107
rect 519 106 525 107
rect 542 106 548 107
rect 559 106 565 107
rect 462 102 463 106
rect 467 102 468 106
rect 462 101 468 102
rect 502 102 503 106
rect 507 102 508 106
rect 502 101 508 102
rect 542 102 543 106
rect 547 102 548 106
rect 542 101 548 102
rect 439 95 445 96
rect 439 94 440 95
rect 432 92 440 94
rect 407 90 413 91
rect 439 91 440 92
rect 444 91 445 95
rect 439 90 445 91
rect 479 95 485 96
rect 479 91 480 95
rect 484 94 485 95
rect 487 95 493 96
rect 487 94 488 95
rect 484 92 488 94
rect 484 91 485 92
rect 479 90 485 91
rect 487 91 488 92
rect 492 91 493 95
rect 487 90 493 91
rect 519 95 525 96
rect 519 91 520 95
rect 524 94 525 95
rect 527 95 533 96
rect 527 94 528 95
rect 524 92 528 94
rect 524 91 525 92
rect 519 90 525 91
rect 527 91 528 92
rect 532 91 533 95
rect 527 90 533 91
rect 559 95 565 96
rect 559 91 560 95
rect 564 94 565 95
rect 568 94 570 112
rect 591 111 597 112
rect 591 107 592 111
rect 596 107 597 111
rect 623 111 629 112
rect 623 110 624 111
rect 616 108 624 110
rect 574 106 580 107
rect 591 106 597 107
rect 606 106 612 107
rect 574 102 575 106
rect 579 102 580 106
rect 574 101 580 102
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 616 96 618 108
rect 623 107 624 108
rect 628 107 629 111
rect 623 106 629 107
rect 564 92 570 94
rect 591 95 597 96
rect 564 91 565 92
rect 559 90 565 91
rect 591 91 592 95
rect 596 94 597 95
rect 604 94 618 96
rect 623 95 629 96
rect 596 92 606 94
rect 596 91 597 92
rect 591 90 597 91
rect 623 91 624 95
rect 628 94 629 95
rect 632 94 634 112
rect 655 111 661 112
rect 655 107 656 111
rect 660 107 661 111
rect 687 111 693 112
rect 687 110 688 111
rect 680 108 688 110
rect 638 106 644 107
rect 655 106 661 107
rect 670 106 676 107
rect 638 102 639 106
rect 643 102 644 106
rect 638 101 644 102
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 680 96 682 108
rect 687 107 688 108
rect 692 107 693 111
rect 719 111 725 112
rect 719 110 720 111
rect 712 108 720 110
rect 687 106 693 107
rect 702 106 708 107
rect 702 102 703 106
rect 707 102 708 106
rect 702 101 708 102
rect 712 96 714 108
rect 719 107 720 108
rect 724 107 725 111
rect 751 111 757 112
rect 751 110 752 111
rect 744 108 752 110
rect 719 106 725 107
rect 734 106 740 107
rect 734 102 735 106
rect 739 102 740 106
rect 734 101 740 102
rect 744 96 746 108
rect 751 107 752 108
rect 756 107 757 111
rect 783 111 789 112
rect 783 110 784 111
rect 776 108 784 110
rect 751 106 757 107
rect 766 106 772 107
rect 766 102 767 106
rect 771 102 772 106
rect 766 101 772 102
rect 776 96 778 108
rect 783 107 784 108
rect 788 107 789 111
rect 815 111 821 112
rect 815 110 816 111
rect 808 108 816 110
rect 783 106 789 107
rect 798 106 804 107
rect 798 102 799 106
rect 803 102 804 106
rect 798 101 804 102
rect 808 96 810 108
rect 815 107 816 108
rect 820 107 821 111
rect 847 111 853 112
rect 847 110 848 111
rect 840 108 848 110
rect 815 106 821 107
rect 830 106 836 107
rect 830 102 831 106
rect 835 102 836 106
rect 830 101 836 102
rect 840 96 842 108
rect 847 107 848 108
rect 852 107 853 111
rect 879 111 885 112
rect 879 110 880 111
rect 872 108 880 110
rect 847 106 853 107
rect 862 106 868 107
rect 862 102 863 106
rect 867 102 868 106
rect 862 101 868 102
rect 872 96 874 108
rect 879 107 880 108
rect 884 107 885 111
rect 911 111 917 112
rect 911 110 912 111
rect 904 108 912 110
rect 879 106 885 107
rect 894 106 900 107
rect 894 102 895 106
rect 899 102 900 106
rect 894 101 900 102
rect 904 96 906 108
rect 911 107 912 108
rect 916 107 917 111
rect 919 111 920 115
rect 924 114 925 115
rect 959 115 965 116
rect 924 112 946 114
rect 924 111 925 112
rect 919 110 925 111
rect 944 110 946 112
rect 951 111 957 112
rect 951 110 952 111
rect 944 108 952 110
rect 951 107 952 108
rect 956 107 957 111
rect 959 111 960 115
rect 964 114 965 115
rect 999 115 1005 116
rect 964 112 986 114
rect 964 111 965 112
rect 959 110 965 111
rect 984 110 986 112
rect 991 111 997 112
rect 991 110 992 111
rect 984 108 992 110
rect 991 107 992 108
rect 996 107 997 111
rect 999 111 1000 115
rect 1004 114 1005 115
rect 1039 115 1045 116
rect 1004 112 1026 114
rect 1004 111 1005 112
rect 999 110 1005 111
rect 1024 110 1026 112
rect 1031 111 1037 112
rect 1031 110 1032 111
rect 1024 108 1032 110
rect 1031 107 1032 108
rect 1036 107 1037 111
rect 1039 111 1040 115
rect 1044 114 1045 115
rect 1087 115 1093 116
rect 1044 112 1074 114
rect 1044 111 1045 112
rect 1039 110 1045 111
rect 1072 110 1074 112
rect 1079 111 1085 112
rect 1079 110 1080 111
rect 1072 108 1080 110
rect 1079 107 1080 108
rect 1084 107 1085 111
rect 1087 111 1088 115
rect 1092 114 1093 115
rect 1127 115 1133 116
rect 1092 112 1114 114
rect 1092 111 1093 112
rect 1087 110 1093 111
rect 1112 110 1114 112
rect 1119 111 1125 112
rect 1119 110 1120 111
rect 1112 108 1120 110
rect 1119 107 1120 108
rect 1124 107 1125 111
rect 1127 111 1128 115
rect 1132 114 1133 115
rect 1207 115 1213 116
rect 1132 112 1161 114
rect 1132 111 1133 112
rect 1127 110 1133 111
rect 1159 111 1165 112
rect 1159 107 1160 111
rect 1164 107 1165 111
rect 1198 111 1205 112
rect 1198 107 1199 111
rect 1204 107 1205 111
rect 1207 111 1208 115
rect 1212 114 1213 115
rect 1247 115 1253 116
rect 1212 112 1234 114
rect 1212 111 1213 112
rect 1207 110 1213 111
rect 1232 110 1234 112
rect 1239 111 1245 112
rect 1239 110 1240 111
rect 1232 108 1240 110
rect 1239 107 1240 108
rect 1244 107 1245 111
rect 1247 111 1248 115
rect 1252 114 1253 115
rect 1319 115 1325 116
rect 1252 112 1274 114
rect 1252 111 1253 112
rect 1247 110 1253 111
rect 1272 110 1274 112
rect 1279 111 1285 112
rect 1279 110 1280 111
rect 1272 108 1280 110
rect 1279 107 1280 108
rect 1284 107 1285 111
rect 1311 111 1317 112
rect 1311 110 1312 111
rect 1304 108 1312 110
rect 911 106 917 107
rect 934 106 940 107
rect 951 106 957 107
rect 974 106 980 107
rect 991 106 997 107
rect 1014 106 1020 107
rect 1031 106 1037 107
rect 1062 106 1068 107
rect 1079 106 1085 107
rect 1102 106 1108 107
rect 1119 106 1125 107
rect 1142 106 1148 107
rect 1159 106 1165 107
rect 1182 106 1188 107
rect 1198 106 1205 107
rect 1222 106 1228 107
rect 1239 106 1245 107
rect 1262 106 1268 107
rect 1279 106 1285 107
rect 1294 106 1300 107
rect 934 102 935 106
rect 939 102 940 106
rect 934 101 940 102
rect 974 102 975 106
rect 979 102 980 106
rect 974 101 980 102
rect 1014 102 1015 106
rect 1019 102 1020 106
rect 1014 101 1020 102
rect 1062 102 1063 106
rect 1067 102 1068 106
rect 1062 101 1068 102
rect 1102 102 1103 106
rect 1107 102 1108 106
rect 1102 101 1108 102
rect 1142 102 1143 106
rect 1147 102 1148 106
rect 1142 101 1148 102
rect 1182 102 1183 106
rect 1187 102 1188 106
rect 1182 101 1188 102
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1262 102 1263 106
rect 1267 102 1268 106
rect 1262 101 1268 102
rect 1294 102 1295 106
rect 1299 102 1300 106
rect 1294 101 1300 102
rect 1304 96 1306 108
rect 1311 107 1312 108
rect 1316 107 1317 111
rect 1319 111 1320 115
rect 1324 114 1325 115
rect 1359 115 1365 116
rect 1324 112 1346 114
rect 1324 111 1325 112
rect 1319 110 1325 111
rect 1344 110 1346 112
rect 1351 111 1357 112
rect 1351 110 1352 111
rect 1344 108 1352 110
rect 1351 107 1352 108
rect 1356 107 1357 111
rect 1359 111 1360 115
rect 1364 114 1365 115
rect 1399 115 1405 116
rect 1364 112 1386 114
rect 1364 111 1365 112
rect 1359 110 1365 111
rect 1384 110 1386 112
rect 1391 111 1397 112
rect 1391 110 1392 111
rect 1384 108 1392 110
rect 1391 107 1392 108
rect 1396 107 1397 111
rect 1399 111 1400 115
rect 1404 114 1405 115
rect 1439 115 1445 116
rect 1404 112 1426 114
rect 1404 111 1405 112
rect 1399 110 1405 111
rect 1424 110 1426 112
rect 1431 111 1437 112
rect 1431 110 1432 111
rect 1424 108 1432 110
rect 1431 107 1432 108
rect 1436 107 1437 111
rect 1439 111 1440 115
rect 1444 114 1445 115
rect 1479 115 1485 116
rect 1444 112 1466 114
rect 1444 111 1445 112
rect 1439 110 1445 111
rect 1464 110 1466 112
rect 1471 111 1477 112
rect 1471 110 1472 111
rect 1464 108 1472 110
rect 1471 107 1472 108
rect 1476 107 1477 111
rect 1479 111 1480 115
rect 1484 114 1485 115
rect 1527 115 1533 116
rect 1484 112 1514 114
rect 1484 111 1485 112
rect 1479 110 1485 111
rect 1512 110 1514 112
rect 1519 111 1525 112
rect 1519 110 1520 111
rect 1512 108 1520 110
rect 1519 107 1520 108
rect 1524 107 1525 111
rect 1527 111 1528 115
rect 1532 114 1533 115
rect 1532 112 1562 114
rect 1616 112 1634 114
rect 1532 111 1533 112
rect 1527 110 1533 111
rect 1560 110 1562 112
rect 1567 111 1573 112
rect 1567 110 1568 111
rect 1560 108 1568 110
rect 1567 107 1568 108
rect 1572 107 1573 111
rect 1607 111 1613 112
rect 1607 107 1608 111
rect 1612 110 1613 111
rect 1616 110 1618 112
rect 1612 108 1618 110
rect 1612 107 1613 108
rect 1311 106 1317 107
rect 1334 106 1340 107
rect 1351 106 1357 107
rect 1374 106 1380 107
rect 1391 106 1397 107
rect 1414 106 1420 107
rect 1431 106 1437 107
rect 1454 106 1460 107
rect 1471 106 1477 107
rect 1502 106 1508 107
rect 1519 106 1525 107
rect 1550 106 1556 107
rect 1567 106 1573 107
rect 1590 106 1596 107
rect 1607 106 1613 107
rect 1622 106 1628 107
rect 1334 102 1335 106
rect 1339 102 1340 106
rect 1334 101 1340 102
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1454 102 1455 106
rect 1459 102 1460 106
rect 1454 101 1460 102
rect 1502 102 1503 106
rect 1507 102 1508 106
rect 1502 101 1508 102
rect 1550 102 1551 106
rect 1555 102 1556 106
rect 1550 101 1556 102
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1622 101 1628 102
rect 628 92 634 94
rect 655 95 661 96
rect 628 91 629 92
rect 623 90 629 91
rect 655 91 656 95
rect 660 94 661 95
rect 668 94 682 96
rect 687 95 693 96
rect 660 92 670 94
rect 660 91 661 92
rect 655 90 661 91
rect 687 91 688 95
rect 692 94 693 95
rect 700 94 714 96
rect 719 95 725 96
rect 692 92 702 94
rect 692 91 693 92
rect 687 90 693 91
rect 719 91 720 95
rect 724 94 725 95
rect 732 94 746 96
rect 751 95 757 96
rect 724 92 734 94
rect 724 91 725 92
rect 719 90 725 91
rect 751 91 752 95
rect 756 94 757 95
rect 764 94 778 96
rect 783 95 789 96
rect 756 92 766 94
rect 756 91 757 92
rect 751 90 757 91
rect 783 91 784 95
rect 788 94 789 95
rect 796 94 810 96
rect 815 95 821 96
rect 788 92 798 94
rect 788 91 789 92
rect 783 90 789 91
rect 815 91 816 95
rect 820 94 821 95
rect 828 94 842 96
rect 847 95 853 96
rect 820 92 830 94
rect 820 91 821 92
rect 815 90 821 91
rect 847 91 848 95
rect 852 94 853 95
rect 860 94 874 96
rect 879 95 885 96
rect 852 92 862 94
rect 852 91 853 92
rect 847 90 853 91
rect 879 91 880 95
rect 884 94 885 95
rect 892 94 906 96
rect 911 95 917 96
rect 884 92 894 94
rect 884 91 885 92
rect 879 90 885 91
rect 911 91 912 95
rect 916 94 917 95
rect 919 95 925 96
rect 919 94 920 95
rect 916 92 920 94
rect 916 91 917 92
rect 911 90 917 91
rect 919 91 920 92
rect 924 91 925 95
rect 919 90 925 91
rect 951 95 957 96
rect 951 91 952 95
rect 956 94 957 95
rect 959 95 965 96
rect 959 94 960 95
rect 956 92 960 94
rect 956 91 957 92
rect 951 90 957 91
rect 959 91 960 92
rect 964 91 965 95
rect 959 90 965 91
rect 991 95 997 96
rect 991 91 992 95
rect 996 94 997 95
rect 999 95 1005 96
rect 999 94 1000 95
rect 996 92 1000 94
rect 996 91 997 92
rect 991 90 997 91
rect 999 91 1000 92
rect 1004 91 1005 95
rect 999 90 1005 91
rect 1031 95 1037 96
rect 1031 91 1032 95
rect 1036 94 1037 95
rect 1039 95 1045 96
rect 1039 94 1040 95
rect 1036 92 1040 94
rect 1036 91 1037 92
rect 1031 90 1037 91
rect 1039 91 1040 92
rect 1044 91 1045 95
rect 1039 90 1045 91
rect 1079 95 1085 96
rect 1079 91 1080 95
rect 1084 94 1085 95
rect 1087 95 1093 96
rect 1087 94 1088 95
rect 1084 92 1088 94
rect 1084 91 1085 92
rect 1079 90 1085 91
rect 1087 91 1088 92
rect 1092 91 1093 95
rect 1087 90 1093 91
rect 1119 95 1125 96
rect 1119 91 1120 95
rect 1124 94 1125 95
rect 1127 95 1133 96
rect 1127 94 1128 95
rect 1124 92 1128 94
rect 1124 91 1125 92
rect 1119 90 1125 91
rect 1127 91 1128 92
rect 1132 91 1133 95
rect 1127 90 1133 91
rect 1158 95 1165 96
rect 1158 91 1159 95
rect 1164 91 1165 95
rect 1158 90 1165 91
rect 1199 95 1205 96
rect 1199 91 1200 95
rect 1204 94 1205 95
rect 1207 95 1213 96
rect 1207 94 1208 95
rect 1204 92 1208 94
rect 1204 91 1205 92
rect 1199 90 1205 91
rect 1207 91 1208 92
rect 1212 91 1213 95
rect 1207 90 1213 91
rect 1239 95 1245 96
rect 1239 91 1240 95
rect 1244 94 1245 95
rect 1247 95 1253 96
rect 1247 94 1248 95
rect 1244 92 1248 94
rect 1244 91 1245 92
rect 1239 90 1245 91
rect 1247 91 1248 92
rect 1252 91 1253 95
rect 1247 90 1253 91
rect 1279 95 1285 96
rect 1279 91 1280 95
rect 1284 94 1285 95
rect 1292 94 1306 96
rect 1311 95 1317 96
rect 1284 92 1294 94
rect 1284 91 1285 92
rect 1279 90 1285 91
rect 1311 91 1312 95
rect 1316 94 1317 95
rect 1319 95 1325 96
rect 1319 94 1320 95
rect 1316 92 1320 94
rect 1316 91 1317 92
rect 1311 90 1317 91
rect 1319 91 1320 92
rect 1324 91 1325 95
rect 1319 90 1325 91
rect 1351 95 1357 96
rect 1351 91 1352 95
rect 1356 94 1357 95
rect 1359 95 1365 96
rect 1359 94 1360 95
rect 1356 92 1360 94
rect 1356 91 1357 92
rect 1351 90 1357 91
rect 1359 91 1360 92
rect 1364 91 1365 95
rect 1359 90 1365 91
rect 1391 95 1397 96
rect 1391 91 1392 95
rect 1396 94 1397 95
rect 1399 95 1405 96
rect 1399 94 1400 95
rect 1396 92 1400 94
rect 1396 91 1397 92
rect 1391 90 1397 91
rect 1399 91 1400 92
rect 1404 91 1405 95
rect 1399 90 1405 91
rect 1431 95 1437 96
rect 1431 91 1432 95
rect 1436 94 1437 95
rect 1439 95 1445 96
rect 1439 94 1440 95
rect 1436 92 1440 94
rect 1436 91 1437 92
rect 1431 90 1437 91
rect 1439 91 1440 92
rect 1444 91 1445 95
rect 1439 90 1445 91
rect 1471 95 1477 96
rect 1471 91 1472 95
rect 1476 94 1477 95
rect 1479 95 1485 96
rect 1479 94 1480 95
rect 1476 92 1480 94
rect 1476 91 1477 92
rect 1471 90 1477 91
rect 1479 91 1480 92
rect 1484 91 1485 95
rect 1479 90 1485 91
rect 1519 95 1525 96
rect 1519 91 1520 95
rect 1524 94 1525 95
rect 1527 95 1533 96
rect 1527 94 1528 95
rect 1524 92 1528 94
rect 1524 91 1525 92
rect 1519 90 1525 91
rect 1527 91 1528 92
rect 1532 91 1533 95
rect 1527 90 1533 91
rect 1567 95 1573 96
rect 1567 91 1568 95
rect 1572 91 1573 95
rect 1632 94 1634 112
rect 1639 111 1645 112
rect 1639 107 1640 111
rect 1644 110 1645 111
rect 1647 111 1653 112
rect 1647 110 1648 111
rect 1644 108 1648 110
rect 1644 107 1645 108
rect 1639 106 1645 107
rect 1647 107 1648 108
rect 1652 107 1653 111
rect 1647 106 1653 107
rect 1662 108 1668 109
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1639 95 1645 96
rect 1639 94 1640 95
rect 1632 92 1640 94
rect 1567 90 1573 91
rect 1639 91 1640 92
rect 1644 91 1645 95
rect 1639 90 1645 91
rect 1662 91 1668 92
rect 110 86 116 87
rect 134 89 140 90
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 462 89 468 90
rect 462 85 463 89
rect 467 85 468 89
rect 462 84 468 85
rect 502 89 508 90
rect 502 85 503 89
rect 507 85 508 89
rect 502 84 508 85
rect 542 89 548 90
rect 542 85 543 89
rect 547 85 548 89
rect 542 84 548 85
rect 574 89 580 90
rect 574 85 575 89
rect 579 85 580 89
rect 574 84 580 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 638 89 644 90
rect 638 85 639 89
rect 643 85 644 89
rect 638 84 644 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 702 89 708 90
rect 702 85 703 89
rect 707 85 708 89
rect 702 84 708 85
rect 734 89 740 90
rect 734 85 735 89
rect 739 85 740 89
rect 734 84 740 85
rect 766 89 772 90
rect 766 85 767 89
rect 771 85 772 89
rect 766 84 772 85
rect 798 89 804 90
rect 798 85 799 89
rect 803 85 804 89
rect 798 84 804 85
rect 830 89 836 90
rect 830 85 831 89
rect 835 85 836 89
rect 830 84 836 85
rect 862 89 868 90
rect 862 85 863 89
rect 867 85 868 89
rect 862 84 868 85
rect 894 89 900 90
rect 894 85 895 89
rect 899 85 900 89
rect 894 84 900 85
rect 934 89 940 90
rect 934 85 935 89
rect 939 85 940 89
rect 934 84 940 85
rect 974 89 980 90
rect 974 85 975 89
rect 979 85 980 89
rect 974 84 980 85
rect 1014 89 1020 90
rect 1014 85 1015 89
rect 1019 85 1020 89
rect 1014 84 1020 85
rect 1062 89 1068 90
rect 1062 85 1063 89
rect 1067 85 1068 89
rect 1062 84 1068 85
rect 1102 89 1108 90
rect 1102 85 1103 89
rect 1107 85 1108 89
rect 1102 84 1108 85
rect 1142 89 1148 90
rect 1142 85 1143 89
rect 1147 85 1148 89
rect 1142 84 1148 85
rect 1182 89 1188 90
rect 1182 85 1183 89
rect 1187 85 1188 89
rect 1182 84 1188 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1262 89 1268 90
rect 1262 85 1263 89
rect 1267 85 1268 89
rect 1262 84 1268 85
rect 1294 89 1300 90
rect 1294 85 1295 89
rect 1299 85 1300 89
rect 1294 84 1300 85
rect 1334 89 1340 90
rect 1334 85 1335 89
rect 1339 85 1340 89
rect 1334 84 1340 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1414 89 1420 90
rect 1414 85 1415 89
rect 1419 85 1420 89
rect 1414 84 1420 85
rect 1454 89 1460 90
rect 1454 85 1455 89
rect 1459 85 1460 89
rect 1454 84 1460 85
rect 1502 89 1508 90
rect 1502 85 1503 89
rect 1507 85 1508 89
rect 1502 84 1508 85
rect 1550 89 1556 90
rect 1550 85 1551 89
rect 1555 85 1556 89
rect 1550 84 1556 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1662 87 1663 91
rect 1667 87 1668 91
rect 1662 86 1668 87
rect 1622 84 1628 85
<< m3c >>
rect 375 1711 379 1715
rect 111 1700 115 1704
rect 255 1698 259 1702
rect 111 1683 115 1687
rect 287 1698 291 1702
rect 319 1698 323 1702
rect 359 1698 363 1702
rect 407 1698 411 1702
rect 471 1707 475 1711
rect 515 1703 519 1707
rect 539 1707 543 1711
rect 455 1698 459 1702
rect 887 1703 891 1707
rect 503 1698 507 1702
rect 551 1698 555 1702
rect 607 1698 611 1702
rect 663 1698 667 1702
rect 727 1698 731 1702
rect 783 1698 787 1702
rect 839 1698 843 1702
rect 895 1698 899 1702
rect 1107 1707 1111 1711
rect 1139 1711 1143 1715
rect 951 1698 955 1702
rect 1007 1698 1011 1702
rect 1063 1698 1067 1702
rect 1119 1698 1123 1702
rect 1175 1698 1179 1702
rect 1263 1703 1267 1707
rect 1271 1707 1275 1711
rect 1459 1707 1463 1711
rect 1231 1698 1235 1702
rect 1287 1698 1291 1702
rect 1335 1698 1339 1702
rect 1375 1698 1379 1702
rect 1423 1698 1427 1702
rect 1471 1698 1475 1702
rect 1519 1698 1523 1702
rect 1663 1700 1667 1704
rect 351 1687 355 1691
rect 375 1687 376 1691
rect 376 1687 379 1691
rect 471 1687 472 1691
rect 472 1687 475 1691
rect 539 1687 543 1691
rect 803 1687 804 1691
rect 804 1687 807 1691
rect 1107 1687 1111 1691
rect 1139 1687 1140 1691
rect 1140 1687 1143 1691
rect 1191 1687 1192 1691
rect 1192 1687 1195 1691
rect 1271 1687 1275 1691
rect 1459 1687 1463 1691
rect 255 1681 259 1685
rect 287 1681 291 1685
rect 319 1681 323 1685
rect 359 1681 363 1685
rect 407 1681 411 1685
rect 455 1681 459 1685
rect 503 1681 507 1685
rect 551 1681 555 1685
rect 607 1681 611 1685
rect 663 1681 667 1685
rect 727 1681 731 1685
rect 783 1681 787 1685
rect 839 1681 843 1685
rect 895 1681 899 1685
rect 951 1681 955 1685
rect 1007 1681 1011 1685
rect 1063 1681 1067 1685
rect 1119 1681 1123 1685
rect 1175 1681 1179 1685
rect 1231 1681 1235 1685
rect 1287 1681 1291 1685
rect 1335 1681 1339 1685
rect 1375 1681 1379 1685
rect 1423 1681 1427 1685
rect 1471 1681 1475 1685
rect 1519 1681 1523 1685
rect 1411 1675 1415 1679
rect 1663 1683 1667 1687
rect 111 1665 115 1669
rect 135 1667 139 1671
rect 167 1667 171 1671
rect 215 1667 219 1671
rect 279 1667 283 1671
rect 343 1667 347 1671
rect 415 1667 419 1671
rect 487 1667 491 1671
rect 151 1659 152 1663
rect 152 1659 155 1663
rect 111 1648 115 1652
rect 135 1650 139 1654
rect 167 1650 171 1654
rect 215 1650 219 1654
rect 279 1650 283 1654
rect 515 1663 519 1667
rect 559 1667 563 1671
rect 631 1667 635 1671
rect 711 1667 715 1671
rect 791 1667 795 1671
rect 871 1667 875 1671
rect 951 1667 955 1671
rect 1031 1667 1035 1671
rect 1103 1667 1107 1671
rect 1175 1667 1179 1671
rect 1247 1667 1251 1671
rect 1319 1667 1323 1671
rect 1391 1667 1395 1671
rect 1455 1667 1459 1671
rect 1519 1667 1523 1671
rect 1583 1667 1587 1671
rect 1623 1667 1627 1671
rect 1663 1665 1667 1669
rect 343 1650 347 1654
rect 415 1650 419 1654
rect 351 1643 355 1647
rect 523 1659 527 1663
rect 679 1659 683 1663
rect 487 1650 491 1654
rect 559 1650 563 1654
rect 631 1650 635 1654
rect 615 1643 619 1647
rect 711 1650 715 1654
rect 887 1659 888 1663
rect 888 1659 891 1663
rect 791 1650 795 1654
rect 871 1650 875 1654
rect 803 1643 807 1647
rect 951 1650 955 1654
rect 1031 1650 1035 1654
rect 1103 1650 1107 1654
rect 963 1643 967 1647
rect 1147 1659 1151 1663
rect 1263 1659 1264 1663
rect 1264 1659 1267 1663
rect 1167 1651 1171 1655
rect 1175 1650 1179 1654
rect 1247 1650 1251 1654
rect 1191 1643 1192 1647
rect 1192 1643 1195 1647
rect 1319 1650 1323 1654
rect 1391 1650 1395 1654
rect 1335 1643 1336 1647
rect 1336 1643 1339 1647
rect 1411 1643 1412 1647
rect 1412 1643 1415 1647
rect 1455 1650 1459 1654
rect 1519 1650 1523 1654
rect 1575 1659 1579 1663
rect 1583 1650 1587 1654
rect 1547 1643 1551 1647
rect 1639 1659 1640 1663
rect 1640 1659 1643 1663
rect 1623 1650 1627 1654
rect 1663 1648 1667 1652
rect 523 1635 527 1639
rect 1147 1635 1151 1639
rect 111 1620 115 1624
rect 151 1623 152 1627
rect 152 1623 155 1627
rect 199 1623 200 1627
rect 200 1623 203 1627
rect 491 1623 492 1627
rect 492 1623 495 1627
rect 499 1627 503 1631
rect 679 1623 680 1627
rect 680 1623 683 1627
rect 815 1623 816 1627
rect 816 1623 819 1627
rect 135 1618 139 1622
rect 183 1618 187 1622
rect 247 1618 251 1622
rect 303 1618 307 1622
rect 359 1618 363 1622
rect 415 1618 419 1622
rect 471 1618 475 1622
rect 535 1618 539 1622
rect 599 1618 603 1622
rect 663 1618 667 1622
rect 727 1618 731 1622
rect 799 1618 803 1622
rect 871 1618 875 1622
rect 943 1618 947 1622
rect 1023 1618 1027 1622
rect 1103 1618 1107 1622
rect 111 1603 115 1607
rect 151 1607 152 1611
rect 152 1607 155 1611
rect 447 1607 451 1611
rect 499 1607 503 1611
rect 615 1607 616 1611
rect 616 1607 619 1611
rect 743 1607 744 1611
rect 744 1607 747 1611
rect 963 1607 964 1611
rect 964 1607 967 1611
rect 1035 1607 1039 1611
rect 1167 1627 1171 1631
rect 1295 1623 1299 1627
rect 1303 1627 1307 1631
rect 1175 1618 1179 1622
rect 1247 1618 1251 1622
rect 1319 1618 1323 1622
rect 1399 1618 1403 1622
rect 1479 1618 1483 1622
rect 1303 1607 1307 1611
rect 1335 1607 1336 1611
rect 1336 1607 1339 1611
rect 1431 1607 1435 1611
rect 1559 1618 1563 1622
rect 1575 1623 1576 1627
rect 1576 1623 1579 1627
rect 1639 1623 1640 1627
rect 1640 1623 1643 1627
rect 1623 1618 1627 1622
rect 1663 1620 1667 1624
rect 1639 1607 1640 1611
rect 1640 1607 1643 1611
rect 135 1601 139 1605
rect 183 1601 187 1605
rect 247 1601 251 1605
rect 303 1601 307 1605
rect 359 1601 363 1605
rect 415 1601 419 1605
rect 471 1601 475 1605
rect 535 1601 539 1605
rect 599 1601 603 1605
rect 663 1601 667 1605
rect 727 1601 731 1605
rect 799 1601 803 1605
rect 871 1601 875 1605
rect 943 1601 947 1605
rect 1023 1601 1027 1605
rect 1103 1601 1107 1605
rect 1175 1601 1179 1605
rect 1247 1601 1251 1605
rect 1319 1601 1323 1605
rect 1399 1601 1403 1605
rect 1479 1601 1483 1605
rect 1559 1601 1563 1605
rect 1623 1601 1627 1605
rect 1663 1603 1667 1607
rect 199 1595 203 1599
rect 111 1585 115 1589
rect 135 1587 139 1591
rect 167 1587 171 1591
rect 223 1587 227 1591
rect 279 1587 283 1591
rect 335 1587 339 1591
rect 383 1587 387 1591
rect 431 1587 435 1591
rect 479 1587 483 1591
rect 535 1587 539 1591
rect 599 1587 603 1591
rect 663 1587 667 1591
rect 727 1587 731 1591
rect 799 1587 803 1591
rect 871 1587 875 1591
rect 951 1587 955 1591
rect 1039 1587 1043 1591
rect 1119 1587 1123 1591
rect 1199 1587 1203 1591
rect 1279 1587 1283 1591
rect 1351 1587 1355 1591
rect 1415 1587 1419 1591
rect 1471 1587 1475 1591
rect 1527 1587 1531 1591
rect 1583 1587 1587 1591
rect 1623 1587 1627 1591
rect 111 1568 115 1572
rect 135 1570 139 1574
rect 167 1570 171 1574
rect 151 1563 152 1567
rect 152 1563 155 1567
rect 183 1579 184 1583
rect 184 1579 187 1583
rect 1663 1585 1667 1589
rect 223 1570 227 1574
rect 279 1570 283 1574
rect 235 1563 239 1567
rect 375 1579 379 1583
rect 335 1570 339 1574
rect 383 1570 387 1574
rect 491 1579 495 1583
rect 431 1570 435 1574
rect 479 1570 483 1574
rect 447 1563 448 1567
rect 448 1563 451 1567
rect 535 1570 539 1574
rect 599 1570 603 1574
rect 663 1570 667 1574
rect 587 1563 591 1567
rect 815 1579 816 1583
rect 816 1579 819 1583
rect 727 1570 731 1574
rect 799 1570 803 1574
rect 871 1570 875 1574
rect 951 1570 955 1574
rect 1039 1570 1043 1574
rect 743 1563 744 1567
rect 744 1563 747 1567
rect 851 1563 855 1567
rect 1031 1563 1035 1567
rect 1119 1570 1123 1574
rect 1211 1579 1215 1583
rect 1295 1579 1296 1583
rect 1296 1579 1299 1583
rect 1363 1579 1367 1583
rect 1199 1570 1203 1574
rect 1279 1570 1283 1574
rect 1351 1570 1355 1574
rect 1415 1570 1419 1574
rect 1287 1563 1291 1567
rect 1431 1563 1432 1567
rect 1432 1563 1435 1567
rect 1483 1579 1487 1583
rect 1547 1579 1548 1583
rect 1548 1579 1551 1583
rect 1471 1570 1475 1574
rect 1527 1570 1531 1574
rect 1583 1570 1587 1574
rect 1623 1570 1627 1574
rect 1663 1568 1667 1572
rect 1599 1563 1600 1567
rect 1600 1563 1603 1567
rect 1639 1563 1640 1567
rect 1640 1563 1643 1567
rect 1483 1555 1487 1559
rect 111 1540 115 1544
rect 135 1538 139 1542
rect 167 1538 171 1542
rect 111 1523 115 1527
rect 151 1527 152 1531
rect 152 1527 155 1531
rect 183 1543 184 1547
rect 184 1543 187 1547
rect 215 1538 219 1542
rect 263 1538 267 1542
rect 235 1527 236 1531
rect 236 1527 239 1531
rect 311 1538 315 1542
rect 351 1543 355 1547
rect 375 1543 376 1547
rect 376 1543 379 1547
rect 895 1543 899 1547
rect 359 1538 363 1542
rect 407 1538 411 1542
rect 455 1538 459 1542
rect 511 1538 515 1542
rect 567 1538 571 1542
rect 631 1538 635 1542
rect 695 1538 699 1542
rect 759 1538 763 1542
rect 831 1538 835 1542
rect 919 1538 923 1542
rect 1007 1538 1011 1542
rect 587 1527 588 1531
rect 588 1527 591 1531
rect 771 1527 775 1531
rect 851 1527 852 1531
rect 852 1527 855 1531
rect 959 1527 963 1531
rect 1095 1538 1099 1542
rect 1183 1538 1187 1542
rect 1211 1543 1215 1547
rect 1327 1543 1331 1547
rect 1363 1543 1367 1547
rect 1371 1547 1375 1551
rect 1263 1538 1267 1542
rect 1335 1538 1339 1542
rect 1407 1538 1411 1542
rect 1471 1538 1475 1542
rect 1527 1538 1531 1542
rect 1583 1538 1587 1542
rect 1623 1538 1627 1542
rect 1663 1540 1667 1544
rect 1280 1527 1284 1531
rect 1371 1527 1375 1531
rect 1599 1527 1600 1531
rect 1600 1527 1603 1531
rect 1639 1527 1640 1531
rect 1640 1527 1643 1531
rect 135 1521 139 1525
rect 167 1521 171 1525
rect 215 1521 219 1525
rect 263 1521 267 1525
rect 311 1521 315 1525
rect 359 1521 363 1525
rect 407 1521 411 1525
rect 455 1521 459 1525
rect 511 1521 515 1525
rect 567 1521 571 1525
rect 631 1521 635 1525
rect 695 1521 699 1525
rect 759 1521 763 1525
rect 831 1521 835 1525
rect 919 1521 923 1525
rect 1007 1521 1011 1525
rect 1095 1521 1099 1525
rect 1183 1521 1187 1525
rect 1263 1521 1267 1525
rect 1335 1521 1339 1525
rect 1407 1521 1411 1525
rect 1471 1521 1475 1525
rect 1527 1521 1531 1525
rect 1583 1521 1587 1525
rect 1623 1521 1627 1525
rect 1663 1523 1667 1527
rect 351 1511 355 1515
rect 111 1501 115 1505
rect 135 1503 139 1507
rect 167 1503 171 1507
rect 223 1503 227 1507
rect 295 1503 299 1507
rect 375 1503 379 1507
rect 111 1484 115 1488
rect 135 1486 139 1490
rect 167 1486 171 1490
rect 183 1487 187 1491
rect 223 1486 227 1490
rect 151 1479 152 1483
rect 152 1479 155 1483
rect 295 1486 299 1490
rect 1327 1511 1331 1515
rect 455 1503 459 1507
rect 527 1503 531 1507
rect 599 1503 603 1507
rect 671 1503 675 1507
rect 743 1503 747 1507
rect 815 1503 819 1507
rect 879 1503 883 1507
rect 943 1503 947 1507
rect 1007 1503 1011 1507
rect 1063 1503 1067 1507
rect 1111 1503 1115 1507
rect 1151 1503 1155 1507
rect 1183 1503 1187 1507
rect 1215 1503 1219 1507
rect 1255 1503 1259 1507
rect 1295 1503 1299 1507
rect 1351 1503 1355 1507
rect 1415 1503 1419 1507
rect 1487 1503 1491 1507
rect 375 1486 379 1490
rect 543 1495 544 1499
rect 544 1495 547 1499
rect 455 1486 459 1490
rect 527 1486 531 1490
rect 599 1486 603 1490
rect 671 1486 675 1490
rect 743 1486 747 1490
rect 771 1487 775 1491
rect 799 1479 803 1483
rect 815 1486 819 1490
rect 895 1495 896 1499
rect 896 1495 899 1499
rect 975 1495 979 1499
rect 879 1486 883 1490
rect 943 1486 947 1490
rect 1007 1486 1011 1490
rect 959 1479 960 1483
rect 960 1479 963 1483
rect 1027 1479 1028 1483
rect 1028 1479 1031 1483
rect 1063 1486 1067 1490
rect 1111 1486 1115 1490
rect 1151 1486 1155 1490
rect 1183 1486 1187 1490
rect 1215 1486 1219 1490
rect 1231 1495 1232 1499
rect 1232 1495 1235 1499
rect 1255 1486 1259 1490
rect 1295 1486 1299 1490
rect 239 1471 243 1475
rect 111 1456 115 1460
rect 135 1454 139 1458
rect 167 1454 171 1458
rect 111 1439 115 1443
rect 151 1443 152 1447
rect 152 1443 155 1447
rect 183 1459 184 1463
rect 184 1459 187 1463
rect 223 1454 227 1458
rect 295 1454 299 1458
rect 239 1443 240 1447
rect 240 1443 243 1447
rect 375 1454 379 1458
rect 463 1459 467 1463
rect 543 1459 544 1463
rect 544 1459 547 1463
rect 1231 1471 1235 1475
rect 1351 1486 1355 1490
rect 1415 1486 1419 1490
rect 1567 1503 1571 1507
rect 1623 1503 1627 1507
rect 1663 1501 1667 1505
rect 1487 1486 1491 1490
rect 1567 1486 1571 1490
rect 1623 1486 1627 1490
rect 1663 1484 1667 1488
rect 1639 1479 1640 1483
rect 1640 1479 1643 1483
rect 1495 1471 1499 1475
rect 455 1454 459 1458
rect 527 1454 531 1458
rect 599 1454 603 1458
rect 663 1454 667 1458
rect 719 1454 723 1458
rect 783 1454 787 1458
rect 847 1454 851 1458
rect 903 1454 907 1458
rect 959 1454 963 1458
rect 799 1443 800 1447
rect 800 1443 803 1447
rect 895 1443 899 1447
rect 975 1459 976 1463
rect 976 1459 979 1463
rect 1015 1454 1019 1458
rect 1071 1454 1075 1458
rect 1027 1443 1031 1447
rect 1119 1454 1123 1458
rect 1147 1459 1151 1463
rect 1571 1459 1575 1463
rect 1159 1454 1163 1458
rect 1207 1454 1211 1458
rect 1263 1454 1267 1458
rect 1327 1454 1331 1458
rect 1399 1454 1403 1458
rect 1479 1454 1483 1458
rect 1559 1454 1563 1458
rect 1623 1454 1627 1458
rect 1663 1456 1667 1460
rect 1495 1443 1496 1447
rect 1496 1443 1499 1447
rect 1639 1443 1640 1447
rect 1640 1443 1643 1447
rect 135 1437 139 1441
rect 167 1437 171 1441
rect 223 1437 227 1441
rect 295 1437 299 1441
rect 375 1437 379 1441
rect 455 1437 459 1441
rect 527 1437 531 1441
rect 599 1437 603 1441
rect 663 1437 667 1441
rect 719 1437 723 1441
rect 783 1437 787 1441
rect 847 1437 851 1441
rect 903 1437 907 1441
rect 959 1437 963 1441
rect 1015 1437 1019 1441
rect 1071 1437 1075 1441
rect 1119 1437 1123 1441
rect 1159 1437 1163 1441
rect 1207 1437 1211 1441
rect 1263 1437 1267 1441
rect 1327 1437 1331 1441
rect 1399 1437 1403 1441
rect 1479 1437 1483 1441
rect 1559 1437 1563 1441
rect 1147 1427 1151 1431
rect 1523 1431 1527 1435
rect 1623 1437 1627 1441
rect 1663 1439 1667 1443
rect 111 1417 115 1421
rect 135 1419 139 1423
rect 167 1419 171 1423
rect 215 1419 219 1423
rect 287 1419 291 1423
rect 359 1419 363 1423
rect 439 1419 443 1423
rect 519 1419 523 1423
rect 599 1419 603 1423
rect 679 1419 683 1423
rect 759 1419 763 1423
rect 831 1419 835 1423
rect 903 1419 907 1423
rect 967 1419 971 1423
rect 1031 1419 1035 1423
rect 1103 1419 1107 1423
rect 1167 1419 1171 1423
rect 1231 1419 1235 1423
rect 1295 1419 1299 1423
rect 111 1400 115 1404
rect 135 1402 139 1406
rect 167 1402 171 1406
rect 151 1395 152 1399
rect 152 1395 155 1399
rect 215 1402 219 1406
rect 231 1411 232 1415
rect 232 1411 235 1415
rect 287 1402 291 1406
rect 243 1395 247 1399
rect 359 1402 363 1406
rect 456 1411 460 1415
rect 439 1402 443 1406
rect 519 1402 523 1406
rect 599 1402 603 1406
rect 679 1402 683 1406
rect 751 1411 755 1415
rect 771 1411 775 1415
rect 759 1402 763 1406
rect 831 1402 835 1406
rect 903 1402 907 1406
rect 967 1402 971 1406
rect 1031 1402 1035 1406
rect 895 1395 899 1399
rect 1103 1402 1107 1406
rect 1167 1402 1171 1406
rect 1359 1419 1363 1423
rect 1415 1419 1419 1423
rect 1463 1419 1467 1423
rect 1503 1419 1507 1423
rect 1551 1419 1555 1423
rect 1591 1419 1595 1423
rect 1623 1419 1627 1423
rect 1663 1417 1667 1421
rect 1231 1402 1235 1406
rect 1295 1402 1299 1406
rect 1359 1402 1363 1406
rect 1415 1402 1419 1406
rect 231 1383 235 1387
rect 771 1387 775 1391
rect 1255 1387 1259 1391
rect 1571 1411 1572 1415
rect 1572 1411 1575 1415
rect 1463 1402 1467 1406
rect 1503 1402 1507 1406
rect 1551 1402 1555 1406
rect 1523 1395 1524 1399
rect 1524 1395 1527 1399
rect 1591 1402 1595 1406
rect 1623 1402 1627 1406
rect 1663 1400 1667 1404
rect 1631 1395 1635 1399
rect 1639 1395 1640 1399
rect 1640 1395 1643 1399
rect 111 1372 115 1376
rect 135 1370 139 1374
rect 111 1355 115 1359
rect 167 1370 171 1374
rect 223 1370 227 1374
rect 287 1370 291 1374
rect 199 1359 203 1363
rect 243 1359 244 1363
rect 244 1359 247 1363
rect 359 1370 363 1374
rect 439 1375 443 1379
rect 519 1375 520 1379
rect 520 1375 523 1379
rect 751 1375 755 1379
rect 903 1375 904 1379
rect 904 1375 907 1379
rect 1319 1375 1320 1379
rect 1320 1375 1323 1379
rect 1643 1375 1644 1379
rect 1644 1375 1647 1379
rect 431 1370 435 1374
rect 503 1370 507 1374
rect 583 1370 587 1374
rect 663 1370 667 1374
rect 743 1370 747 1374
rect 815 1370 819 1374
rect 887 1370 891 1374
rect 959 1370 963 1374
rect 1031 1370 1035 1374
rect 1103 1370 1107 1374
rect 1175 1370 1179 1374
rect 1239 1370 1243 1374
rect 1303 1370 1307 1374
rect 1367 1370 1371 1374
rect 1431 1370 1435 1374
rect 1495 1370 1499 1374
rect 1567 1370 1571 1374
rect 1623 1370 1627 1374
rect 1663 1372 1667 1376
rect 711 1359 715 1363
rect 135 1353 139 1357
rect 167 1353 171 1357
rect 223 1353 227 1357
rect 287 1353 291 1357
rect 359 1353 363 1357
rect 431 1353 435 1357
rect 503 1353 507 1357
rect 583 1353 587 1357
rect 663 1353 667 1357
rect 743 1353 747 1357
rect 815 1353 819 1357
rect 519 1347 523 1351
rect 1255 1359 1256 1363
rect 1256 1359 1259 1363
rect 1487 1359 1491 1363
rect 887 1353 891 1357
rect 959 1353 963 1357
rect 1031 1353 1035 1357
rect 1103 1353 1107 1357
rect 1175 1353 1179 1357
rect 1239 1353 1243 1357
rect 1303 1353 1307 1357
rect 1367 1353 1371 1357
rect 1431 1353 1435 1357
rect 1495 1353 1499 1357
rect 1567 1353 1571 1357
rect 903 1347 907 1351
rect 111 1337 115 1341
rect 135 1339 139 1343
rect 183 1339 187 1343
rect 239 1339 243 1343
rect 295 1339 299 1343
rect 351 1339 355 1343
rect 399 1339 403 1343
rect 455 1339 459 1343
rect 511 1339 515 1343
rect 567 1339 571 1343
rect 631 1339 635 1343
rect 695 1339 699 1343
rect 759 1339 763 1343
rect 823 1339 827 1343
rect 887 1339 891 1343
rect 959 1339 963 1343
rect 1023 1339 1027 1343
rect 1087 1339 1091 1343
rect 1151 1339 1155 1343
rect 151 1331 152 1335
rect 152 1331 155 1335
rect 111 1320 115 1324
rect 135 1322 139 1326
rect 183 1322 187 1326
rect 239 1322 243 1326
rect 295 1322 299 1326
rect 199 1315 200 1319
rect 200 1315 203 1319
rect 351 1322 355 1326
rect 399 1322 403 1326
rect 439 1331 443 1335
rect 455 1322 459 1326
rect 511 1322 515 1326
rect 391 1307 395 1311
rect 623 1331 627 1335
rect 643 1331 647 1335
rect 739 1331 743 1335
rect 567 1322 571 1326
rect 631 1322 635 1326
rect 695 1322 699 1326
rect 759 1322 763 1326
rect 823 1322 827 1326
rect 711 1315 712 1319
rect 712 1315 715 1319
rect 739 1315 743 1319
rect 887 1322 891 1326
rect 643 1307 647 1311
rect 959 1322 963 1326
rect 1023 1322 1027 1326
rect 1319 1347 1323 1351
rect 1635 1359 1639 1363
rect 1623 1353 1627 1357
rect 1663 1355 1667 1359
rect 1215 1339 1219 1343
rect 1279 1339 1283 1343
rect 1343 1339 1347 1343
rect 1407 1339 1411 1343
rect 1479 1339 1483 1343
rect 1559 1339 1563 1343
rect 1623 1339 1627 1343
rect 1663 1337 1667 1341
rect 1087 1322 1091 1326
rect 1151 1322 1155 1326
rect 1215 1322 1219 1326
rect 1279 1322 1283 1326
rect 1343 1322 1347 1326
rect 1375 1331 1379 1335
rect 1383 1331 1387 1335
rect 1407 1322 1411 1326
rect 1479 1322 1483 1326
rect 1559 1322 1563 1326
rect 1487 1315 1491 1319
rect 1575 1331 1576 1335
rect 1576 1331 1579 1335
rect 1651 1331 1655 1335
rect 1623 1322 1627 1326
rect 1663 1320 1667 1324
rect 1095 1307 1099 1311
rect 1383 1307 1387 1311
rect 1575 1307 1579 1311
rect 111 1288 115 1292
rect 151 1291 152 1295
rect 152 1291 155 1295
rect 295 1291 296 1295
rect 296 1291 299 1295
rect 135 1286 139 1290
rect 183 1286 187 1290
rect 231 1286 235 1290
rect 279 1286 283 1290
rect 327 1286 331 1290
rect 375 1286 379 1290
rect 431 1286 435 1290
rect 487 1286 491 1290
rect 543 1286 547 1290
rect 111 1271 115 1275
rect 243 1275 247 1279
rect 391 1275 392 1279
rect 392 1275 395 1279
rect 451 1275 452 1279
rect 452 1275 455 1279
rect 599 1291 603 1295
rect 623 1291 624 1295
rect 624 1291 627 1295
rect 735 1291 736 1295
rect 736 1291 739 1295
rect 783 1291 787 1295
rect 607 1286 611 1290
rect 663 1286 667 1290
rect 719 1286 723 1290
rect 775 1286 779 1290
rect 831 1286 835 1290
rect 895 1286 899 1290
rect 959 1286 963 1290
rect 1023 1286 1027 1290
rect 1079 1286 1083 1290
rect 1143 1286 1147 1290
rect 1207 1286 1211 1290
rect 759 1275 763 1279
rect 1095 1275 1096 1279
rect 1096 1275 1099 1279
rect 1155 1275 1159 1279
rect 1279 1286 1283 1290
rect 1351 1291 1355 1295
rect 1375 1291 1376 1295
rect 1376 1291 1379 1295
rect 1359 1286 1363 1290
rect 1447 1286 1451 1290
rect 1543 1286 1547 1290
rect 1623 1286 1627 1290
rect 1663 1288 1667 1292
rect 135 1269 139 1273
rect 183 1269 187 1273
rect 231 1269 235 1273
rect 279 1269 283 1273
rect 327 1269 331 1273
rect 375 1269 379 1273
rect 431 1269 435 1273
rect 487 1269 491 1273
rect 543 1269 547 1273
rect 607 1269 611 1273
rect 663 1269 667 1273
rect 599 1263 603 1267
rect 719 1269 723 1273
rect 775 1269 779 1273
rect 831 1269 835 1273
rect 895 1269 899 1273
rect 959 1269 963 1273
rect 1023 1269 1027 1273
rect 1079 1269 1083 1273
rect 1143 1269 1147 1273
rect 1207 1269 1211 1273
rect 1279 1269 1283 1273
rect 1359 1269 1363 1273
rect 1447 1269 1451 1273
rect 1543 1269 1547 1273
rect 1351 1263 1355 1267
rect 1643 1275 1644 1279
rect 1644 1275 1647 1279
rect 1623 1269 1627 1273
rect 1663 1271 1667 1275
rect 111 1253 115 1257
rect 135 1255 139 1259
rect 167 1255 171 1259
rect 223 1255 227 1259
rect 279 1255 283 1259
rect 327 1255 331 1259
rect 383 1255 387 1259
rect 439 1255 443 1259
rect 495 1255 499 1259
rect 551 1255 555 1259
rect 607 1255 611 1259
rect 663 1255 667 1259
rect 719 1255 723 1259
rect 767 1255 771 1259
rect 815 1255 819 1259
rect 871 1255 875 1259
rect 927 1255 931 1259
rect 983 1255 987 1259
rect 1039 1255 1043 1259
rect 1095 1255 1099 1259
rect 1159 1255 1163 1259
rect 1231 1255 1235 1259
rect 1319 1255 1323 1259
rect 1423 1255 1427 1259
rect 1535 1255 1539 1259
rect 1623 1255 1627 1259
rect 1663 1253 1667 1257
rect 151 1247 152 1251
rect 152 1247 155 1251
rect 111 1236 115 1240
rect 135 1238 139 1242
rect 167 1238 171 1242
rect 295 1247 296 1251
rect 296 1247 299 1251
rect 223 1238 227 1242
rect 279 1238 283 1242
rect 243 1231 244 1235
rect 244 1231 247 1235
rect 327 1238 331 1242
rect 383 1238 387 1242
rect 439 1238 443 1242
rect 399 1231 400 1235
rect 400 1231 403 1235
rect 451 1231 455 1235
rect 495 1238 499 1242
rect 551 1238 555 1242
rect 619 1247 623 1251
rect 607 1238 611 1242
rect 663 1238 667 1242
rect 719 1238 723 1242
rect 735 1247 736 1251
rect 736 1247 739 1251
rect 783 1247 784 1251
rect 784 1247 787 1251
rect 767 1238 771 1242
rect 815 1238 819 1242
rect 759 1231 763 1235
rect 871 1238 875 1242
rect 927 1238 931 1242
rect 111 1204 115 1208
rect 151 1207 152 1211
rect 152 1207 155 1211
rect 135 1202 139 1206
rect 111 1187 115 1191
rect 299 1207 300 1211
rect 300 1207 303 1211
rect 307 1211 311 1215
rect 619 1219 623 1223
rect 907 1231 911 1235
rect 983 1238 987 1242
rect 1051 1247 1055 1251
rect 1039 1238 1043 1242
rect 1095 1238 1099 1242
rect 1159 1238 1163 1242
rect 1151 1231 1155 1235
rect 1231 1238 1235 1242
rect 1319 1238 1323 1242
rect 1423 1238 1427 1242
rect 1503 1247 1507 1251
rect 1639 1247 1640 1251
rect 1640 1247 1643 1251
rect 1535 1238 1539 1242
rect 1623 1238 1627 1242
rect 1663 1236 1667 1240
rect 1651 1231 1655 1235
rect 1051 1223 1055 1227
rect 783 1207 784 1211
rect 784 1207 787 1211
rect 1007 1207 1011 1211
rect 1023 1207 1027 1211
rect 1503 1219 1507 1223
rect 1639 1207 1640 1211
rect 1640 1207 1643 1211
rect 167 1202 171 1206
rect 223 1202 227 1206
rect 279 1202 283 1206
rect 335 1202 339 1206
rect 383 1202 387 1206
rect 431 1202 435 1206
rect 487 1202 491 1206
rect 543 1202 547 1206
rect 599 1202 603 1206
rect 655 1202 659 1206
rect 711 1202 715 1206
rect 767 1202 771 1206
rect 823 1202 827 1206
rect 887 1202 891 1206
rect 951 1202 955 1206
rect 1015 1202 1019 1206
rect 1079 1202 1083 1206
rect 1143 1202 1147 1206
rect 1207 1202 1211 1206
rect 1279 1202 1283 1206
rect 1359 1202 1363 1206
rect 1447 1202 1451 1206
rect 1543 1202 1547 1206
rect 1623 1202 1627 1206
rect 1663 1204 1667 1208
rect 239 1191 240 1195
rect 240 1191 243 1195
rect 307 1191 311 1195
rect 399 1191 400 1195
rect 400 1191 403 1195
rect 907 1191 908 1195
rect 908 1191 911 1195
rect 135 1185 139 1189
rect 167 1185 171 1189
rect 223 1185 227 1189
rect 279 1185 283 1189
rect 335 1185 339 1189
rect 383 1185 387 1189
rect 431 1185 435 1189
rect 487 1185 491 1189
rect 543 1185 547 1189
rect 599 1185 603 1189
rect 655 1185 659 1189
rect 711 1185 715 1189
rect 495 1179 499 1183
rect 767 1185 771 1189
rect 783 1183 787 1187
rect 823 1185 827 1189
rect 887 1185 891 1189
rect 951 1185 955 1189
rect 1015 1185 1019 1189
rect 1079 1185 1083 1189
rect 1007 1179 1011 1183
rect 1143 1185 1147 1189
rect 1207 1185 1211 1189
rect 1279 1185 1283 1189
rect 1359 1185 1363 1189
rect 1447 1185 1451 1189
rect 1543 1185 1547 1189
rect 1235 1179 1239 1183
rect 1639 1191 1640 1195
rect 1640 1191 1643 1195
rect 1623 1185 1627 1189
rect 1663 1187 1667 1191
rect 111 1165 115 1169
rect 135 1167 139 1171
rect 167 1167 171 1171
rect 223 1167 227 1171
rect 287 1167 291 1171
rect 351 1167 355 1171
rect 415 1167 419 1171
rect 471 1167 475 1171
rect 535 1167 539 1171
rect 599 1167 603 1171
rect 663 1167 667 1171
rect 727 1167 731 1171
rect 783 1167 787 1171
rect 839 1167 843 1171
rect 859 1171 863 1175
rect 903 1167 907 1171
rect 967 1167 971 1171
rect 1031 1167 1035 1171
rect 1095 1167 1099 1171
rect 1159 1167 1163 1171
rect 1215 1167 1219 1171
rect 1279 1167 1283 1171
rect 1343 1167 1347 1171
rect 1407 1167 1411 1171
rect 1479 1167 1483 1171
rect 1559 1167 1563 1171
rect 1623 1167 1627 1171
rect 1663 1165 1667 1169
rect 155 1159 156 1163
rect 156 1159 159 1163
rect 111 1148 115 1152
rect 135 1150 139 1154
rect 167 1150 171 1154
rect 299 1159 303 1163
rect 223 1150 227 1154
rect 287 1150 291 1154
rect 239 1143 240 1147
rect 240 1143 243 1147
rect 351 1150 355 1154
rect 415 1150 419 1154
rect 471 1150 475 1154
rect 479 1143 483 1147
rect 488 1143 492 1147
rect 535 1150 539 1154
rect 599 1150 603 1154
rect 663 1150 667 1154
rect 727 1150 731 1154
rect 799 1159 800 1163
rect 800 1159 803 1163
rect 1023 1159 1027 1163
rect 783 1150 787 1154
rect 839 1150 843 1154
rect 859 1143 860 1147
rect 860 1143 863 1147
rect 903 1150 907 1154
rect 967 1150 971 1154
rect 1031 1150 1035 1154
rect 1043 1143 1047 1147
rect 1095 1150 1099 1154
rect 1159 1150 1163 1154
rect 1215 1150 1219 1154
rect 1279 1150 1283 1154
rect 1235 1143 1236 1147
rect 1236 1143 1239 1147
rect 1343 1150 1347 1154
rect 1407 1150 1411 1154
rect 1479 1150 1483 1154
rect 1559 1150 1563 1154
rect 1623 1150 1627 1154
rect 1663 1148 1667 1152
rect 1639 1143 1640 1147
rect 1640 1143 1643 1147
rect 111 1116 115 1120
rect 155 1119 159 1123
rect 143 1114 147 1118
rect 175 1114 179 1118
rect 299 1123 303 1127
rect 799 1131 803 1135
rect 1103 1131 1107 1135
rect 1131 1119 1135 1123
rect 1163 1119 1167 1123
rect 1559 1119 1560 1123
rect 1560 1119 1563 1123
rect 215 1114 219 1118
rect 271 1114 275 1118
rect 335 1114 339 1118
rect 399 1114 403 1118
rect 463 1114 467 1118
rect 527 1114 531 1118
rect 599 1114 603 1118
rect 663 1114 667 1118
rect 727 1114 731 1118
rect 791 1114 795 1118
rect 855 1114 859 1118
rect 911 1114 915 1118
rect 967 1114 971 1118
rect 1023 1114 1027 1118
rect 1087 1114 1091 1118
rect 1151 1114 1155 1118
rect 1215 1114 1219 1118
rect 1279 1114 1283 1118
rect 1335 1114 1339 1118
rect 1391 1114 1395 1118
rect 1447 1114 1451 1118
rect 1495 1114 1499 1118
rect 1543 1114 1547 1118
rect 1591 1114 1595 1118
rect 111 1099 115 1103
rect 143 1097 147 1101
rect 175 1097 179 1101
rect 215 1097 219 1101
rect 271 1097 275 1101
rect 235 1091 239 1095
rect 479 1103 480 1107
rect 480 1103 483 1107
rect 903 1103 907 1107
rect 1043 1103 1044 1107
rect 1044 1103 1047 1107
rect 1103 1103 1104 1107
rect 1104 1103 1107 1107
rect 1623 1114 1627 1118
rect 1663 1116 1667 1120
rect 1639 1103 1640 1107
rect 1640 1103 1643 1107
rect 335 1097 339 1101
rect 399 1097 403 1101
rect 463 1097 467 1101
rect 527 1097 531 1101
rect 599 1097 603 1101
rect 663 1097 667 1101
rect 727 1097 731 1101
rect 791 1097 795 1101
rect 855 1097 859 1101
rect 911 1097 915 1101
rect 967 1097 971 1101
rect 1023 1097 1027 1101
rect 1087 1097 1091 1101
rect 1151 1097 1155 1101
rect 1215 1097 1219 1101
rect 1279 1097 1283 1101
rect 1131 1091 1135 1095
rect 1335 1097 1339 1101
rect 1391 1097 1395 1101
rect 1447 1097 1451 1101
rect 1495 1097 1499 1101
rect 1379 1091 1383 1095
rect 1543 1097 1547 1101
rect 1591 1097 1595 1101
rect 1623 1097 1627 1101
rect 1663 1099 1667 1103
rect 1559 1087 1563 1091
rect 111 1077 115 1081
rect 215 1079 219 1083
rect 247 1079 251 1083
rect 279 1079 283 1083
rect 311 1079 315 1083
rect 351 1079 355 1083
rect 391 1079 395 1083
rect 439 1079 443 1083
rect 503 1079 507 1083
rect 575 1079 579 1083
rect 655 1079 659 1083
rect 735 1079 739 1083
rect 815 1079 819 1083
rect 895 1079 899 1083
rect 967 1079 971 1083
rect 1039 1079 1043 1083
rect 1111 1079 1115 1083
rect 1175 1079 1179 1083
rect 1239 1079 1243 1083
rect 1303 1079 1307 1083
rect 1359 1079 1363 1083
rect 1415 1079 1419 1083
rect 1463 1079 1467 1083
rect 1503 1079 1507 1083
rect 1551 1079 1555 1083
rect 1591 1079 1595 1083
rect 1623 1079 1627 1083
rect 1663 1077 1667 1081
rect 111 1060 115 1064
rect 215 1062 219 1066
rect 247 1062 251 1066
rect 235 1055 236 1059
rect 236 1055 239 1059
rect 279 1062 283 1066
rect 299 1071 300 1075
rect 300 1071 303 1075
rect 311 1062 315 1066
rect 351 1062 355 1066
rect 391 1062 395 1066
rect 439 1062 443 1066
rect 503 1062 507 1066
rect 575 1062 579 1066
rect 667 1071 671 1075
rect 807 1071 811 1075
rect 655 1062 659 1066
rect 735 1062 739 1066
rect 815 1062 819 1066
rect 895 1062 899 1066
rect 967 1062 971 1066
rect 1039 1062 1043 1066
rect 903 1055 907 1059
rect 1163 1071 1167 1075
rect 1187 1071 1191 1075
rect 1111 1062 1115 1066
rect 1175 1062 1179 1066
rect 1239 1062 1243 1066
rect 1303 1062 1307 1066
rect 1359 1062 1363 1066
rect 1311 1055 1315 1059
rect 1379 1055 1380 1059
rect 1380 1055 1383 1059
rect 1415 1062 1419 1066
rect 1463 1062 1467 1066
rect 1503 1062 1507 1066
rect 1551 1062 1555 1066
rect 1591 1062 1595 1066
rect 1607 1063 1611 1067
rect 1623 1062 1627 1066
rect 1663 1060 1667 1064
rect 1639 1055 1640 1059
rect 1640 1055 1643 1059
rect 471 1047 475 1051
rect 667 1043 671 1047
rect 1187 1047 1191 1051
rect 111 1028 115 1032
rect 303 1031 307 1035
rect 295 1026 299 1030
rect 111 1011 115 1015
rect 327 1026 331 1030
rect 359 1026 363 1030
rect 391 1026 395 1030
rect 423 1026 427 1030
rect 807 1031 811 1035
rect 975 1031 976 1035
rect 976 1031 979 1035
rect 1447 1043 1451 1047
rect 455 1026 459 1030
rect 503 1026 507 1030
rect 559 1026 563 1030
rect 631 1026 635 1030
rect 711 1026 715 1030
rect 799 1026 803 1030
rect 879 1026 883 1030
rect 959 1026 963 1030
rect 1031 1026 1035 1030
rect 1095 1026 1099 1030
rect 1159 1026 1163 1030
rect 1223 1026 1227 1030
rect 1279 1026 1283 1030
rect 1335 1026 1339 1030
rect 1383 1026 1387 1030
rect 1431 1026 1435 1030
rect 1479 1026 1483 1030
rect 1535 1026 1539 1030
rect 471 1015 472 1019
rect 472 1015 475 1019
rect 295 1009 299 1013
rect 327 1009 331 1013
rect 359 1009 363 1013
rect 391 1009 395 1013
rect 423 1009 427 1013
rect 455 1009 459 1013
rect 503 1009 507 1013
rect 559 1009 563 1013
rect 631 1009 635 1013
rect 711 1009 715 1013
rect 303 1003 307 1007
rect 111 993 115 997
rect 247 995 251 999
rect 279 995 283 999
rect 311 995 315 999
rect 343 995 347 999
rect 383 995 387 999
rect 423 995 427 999
rect 111 976 115 980
rect 247 978 251 982
rect 279 978 283 982
rect 311 978 315 982
rect 343 978 347 982
rect 511 1003 515 1007
rect 891 1015 895 1019
rect 1311 1015 1315 1019
rect 1415 1015 1419 1019
rect 1447 1015 1448 1019
rect 1448 1015 1451 1019
rect 1555 1031 1556 1035
rect 1556 1031 1559 1035
rect 1607 1031 1608 1035
rect 1608 1031 1611 1035
rect 1591 1026 1595 1030
rect 1623 1026 1627 1030
rect 1663 1028 1667 1032
rect 1639 1015 1640 1019
rect 1640 1015 1643 1019
rect 799 1009 803 1013
rect 879 1009 883 1013
rect 959 1009 963 1013
rect 1031 1009 1035 1013
rect 1095 1009 1099 1013
rect 1159 1009 1163 1013
rect 1223 1009 1227 1013
rect 1279 1009 1283 1013
rect 1335 1009 1339 1013
rect 1383 1009 1387 1013
rect 1431 1009 1435 1013
rect 1479 1009 1483 1013
rect 1535 1009 1539 1013
rect 1591 1009 1595 1013
rect 1623 1009 1627 1013
rect 1663 1011 1667 1015
rect 975 1003 979 1007
rect 479 995 483 999
rect 543 995 547 999
rect 615 995 619 999
rect 687 995 691 999
rect 759 995 763 999
rect 831 995 835 999
rect 903 995 907 999
rect 967 995 971 999
rect 1031 995 1035 999
rect 1095 995 1099 999
rect 1159 995 1163 999
rect 1223 995 1227 999
rect 383 978 387 982
rect 423 978 427 982
rect 479 978 483 982
rect 511 971 515 975
rect 543 978 547 982
rect 615 978 619 982
rect 675 987 679 991
rect 807 987 811 991
rect 687 978 691 982
rect 759 978 763 982
rect 831 978 835 982
rect 903 978 907 982
rect 967 978 971 982
rect 891 971 895 975
rect 1031 978 1035 982
rect 1095 978 1099 982
rect 1159 978 1163 982
rect 1287 995 1291 999
rect 1343 995 1347 999
rect 1399 995 1403 999
rect 1447 995 1451 999
rect 1495 995 1499 999
rect 1543 995 1547 999
rect 1591 995 1595 999
rect 1623 995 1627 999
rect 1663 993 1667 997
rect 1323 987 1327 991
rect 1223 978 1227 982
rect 1287 978 1291 982
rect 1343 978 1347 982
rect 1399 978 1403 982
rect 1447 978 1451 982
rect 1495 978 1499 982
rect 1415 971 1416 975
rect 1416 971 1419 975
rect 1459 971 1463 975
rect 1555 987 1559 991
rect 1607 987 1608 991
rect 1608 987 1611 991
rect 1543 978 1547 982
rect 1591 978 1595 982
rect 1623 978 1627 982
rect 1663 976 1667 980
rect 1639 971 1640 975
rect 1640 971 1643 975
rect 415 963 419 967
rect 111 948 115 952
rect 187 951 188 955
rect 188 951 191 955
rect 167 946 171 950
rect 199 946 203 950
rect 675 963 679 967
rect 1183 963 1187 967
rect 239 946 243 950
rect 287 946 291 950
rect 343 946 347 950
rect 407 946 411 950
rect 471 946 475 950
rect 535 946 539 950
rect 599 946 603 950
rect 663 946 667 950
rect 727 946 731 950
rect 791 946 795 950
rect 111 931 115 935
rect 419 935 423 939
rect 675 935 679 939
rect 759 935 763 939
rect 807 951 808 955
rect 808 951 811 955
rect 863 951 864 955
rect 864 951 867 955
rect 1323 959 1327 963
rect 1487 963 1491 967
rect 847 946 851 950
rect 911 946 915 950
rect 975 946 979 950
rect 1039 946 1043 950
rect 1103 946 1107 950
rect 1167 946 1171 950
rect 1231 946 1235 950
rect 1287 946 1291 950
rect 1183 935 1184 939
rect 1184 935 1187 939
rect 1343 946 1347 950
rect 1391 946 1395 950
rect 1431 946 1435 950
rect 1471 946 1475 950
rect 1511 946 1515 950
rect 1459 939 1463 943
rect 1487 935 1488 939
rect 1488 935 1491 939
rect 1551 946 1555 950
rect 1583 951 1587 955
rect 1607 951 1608 955
rect 1608 951 1611 955
rect 1591 946 1595 950
rect 1623 946 1627 950
rect 1663 948 1667 952
rect 167 929 171 933
rect 199 929 203 933
rect 239 929 243 933
rect 287 929 291 933
rect 343 929 347 933
rect 407 929 411 933
rect 471 929 475 933
rect 535 929 539 933
rect 599 929 603 933
rect 663 929 667 933
rect 727 929 731 933
rect 791 929 795 933
rect 847 929 851 933
rect 911 929 915 933
rect 975 929 979 933
rect 1039 929 1043 933
rect 1103 929 1107 933
rect 1167 929 1171 933
rect 1231 929 1235 933
rect 187 919 191 923
rect 111 909 115 913
rect 135 911 139 915
rect 167 911 171 915
rect 207 911 211 915
rect 271 911 275 915
rect 335 911 339 915
rect 407 911 411 915
rect 111 892 115 896
rect 135 894 139 898
rect 167 894 171 898
rect 207 894 211 898
rect 271 894 275 898
rect 863 919 867 923
rect 1175 923 1179 927
rect 1287 929 1291 933
rect 1343 929 1347 933
rect 1391 929 1395 933
rect 1431 929 1435 933
rect 1471 929 1475 933
rect 1511 929 1515 933
rect 1551 929 1555 933
rect 1591 929 1595 933
rect 1623 929 1627 933
rect 1583 923 1587 927
rect 1663 931 1667 935
rect 471 911 475 915
rect 535 911 539 915
rect 591 911 595 915
rect 647 911 651 915
rect 703 911 707 915
rect 751 911 755 915
rect 799 911 803 915
rect 847 911 851 915
rect 903 911 907 915
rect 959 911 963 915
rect 1023 911 1027 915
rect 335 894 339 898
rect 487 903 488 907
rect 488 903 491 907
rect 407 894 411 898
rect 471 894 475 898
rect 535 894 539 898
rect 667 903 668 907
rect 668 903 671 907
rect 591 894 595 898
rect 647 894 651 898
rect 675 895 679 899
rect 703 894 707 898
rect 751 894 755 898
rect 799 894 803 898
rect 759 887 763 891
rect 815 887 816 891
rect 816 887 819 891
rect 847 894 851 898
rect 903 894 907 898
rect 959 894 963 898
rect 1023 894 1027 898
rect 1087 911 1091 915
rect 1143 911 1147 915
rect 1199 911 1203 915
rect 1255 911 1259 915
rect 1319 911 1323 915
rect 1383 911 1387 915
rect 1663 909 1667 913
rect 1087 894 1091 898
rect 1143 894 1147 898
rect 1175 887 1179 891
rect 1199 894 1203 898
rect 1255 894 1259 898
rect 1319 894 1323 898
rect 1375 903 1379 907
rect 1383 894 1387 898
rect 1663 892 1667 896
rect 423 879 427 883
rect 111 860 115 864
rect 151 863 152 867
rect 152 863 155 867
rect 135 858 139 862
rect 111 843 115 847
rect 487 863 488 867
rect 488 863 491 867
rect 559 871 563 875
rect 647 863 651 867
rect 667 863 671 867
rect 1119 875 1123 879
rect 167 858 171 862
rect 207 858 211 862
rect 271 858 275 862
rect 335 858 339 862
rect 407 858 411 862
rect 471 858 475 862
rect 535 858 539 862
rect 599 858 603 862
rect 655 858 659 862
rect 703 858 707 862
rect 751 858 755 862
rect 799 858 803 862
rect 847 858 851 862
rect 423 847 424 851
rect 424 847 427 851
rect 552 847 556 851
rect 619 847 620 851
rect 620 847 623 851
rect 667 847 671 851
rect 815 847 816 851
rect 816 847 819 851
rect 903 858 907 862
rect 967 858 971 862
rect 1055 863 1056 867
rect 1056 863 1059 867
rect 1375 875 1379 879
rect 1039 858 1043 862
rect 1103 858 1107 862
rect 1167 858 1171 862
rect 1231 858 1235 862
rect 1287 858 1291 862
rect 1343 858 1347 862
rect 1399 858 1403 862
rect 1463 858 1467 862
rect 1663 860 1667 864
rect 1119 847 1120 851
rect 1120 847 1123 851
rect 135 841 139 845
rect 167 841 171 845
rect 207 841 211 845
rect 271 841 275 845
rect 335 841 339 845
rect 407 841 411 845
rect 471 841 475 845
rect 535 841 539 845
rect 599 841 603 845
rect 655 841 659 845
rect 703 841 707 845
rect 751 841 755 845
rect 691 835 695 839
rect 799 841 803 845
rect 847 841 851 845
rect 903 841 907 845
rect 967 841 971 845
rect 1039 841 1043 845
rect 1103 841 1107 845
rect 1167 841 1171 845
rect 1231 841 1235 845
rect 1287 841 1291 845
rect 1343 841 1347 845
rect 1399 841 1403 845
rect 1463 841 1467 845
rect 1331 835 1335 839
rect 1663 843 1667 847
rect 111 825 115 829
rect 135 827 139 831
rect 167 827 171 831
rect 215 827 219 831
rect 279 827 283 831
rect 343 827 347 831
rect 415 827 419 831
rect 479 827 483 831
rect 543 827 547 831
rect 607 827 611 831
rect 671 827 675 831
rect 735 827 739 831
rect 791 827 795 831
rect 847 827 851 831
rect 911 827 915 831
rect 975 827 979 831
rect 1039 827 1043 831
rect 1111 827 1115 831
rect 1183 827 1187 831
rect 1247 827 1251 831
rect 1311 827 1315 831
rect 1367 827 1371 831
rect 1423 827 1427 831
rect 1479 827 1483 831
rect 1535 827 1539 831
rect 1591 827 1595 831
rect 1663 825 1667 829
rect 151 819 152 823
rect 152 819 155 823
rect 111 808 115 812
rect 135 810 139 814
rect 167 810 171 814
rect 215 810 219 814
rect 279 810 283 814
rect 287 803 291 807
rect 343 810 347 814
rect 403 819 407 823
rect 535 819 539 823
rect 415 810 419 814
rect 479 810 483 814
rect 543 810 547 814
rect 607 810 611 814
rect 671 810 675 814
rect 619 803 623 807
rect 691 803 692 807
rect 692 803 695 807
rect 735 810 739 814
rect 791 810 795 814
rect 859 819 863 823
rect 847 810 851 814
rect 911 810 915 814
rect 975 810 979 814
rect 403 795 407 799
rect 1055 819 1056 823
rect 1056 819 1059 823
rect 1039 810 1043 814
rect 1111 810 1115 814
rect 1183 810 1187 814
rect 1247 810 1251 814
rect 1311 810 1315 814
rect 1303 803 1307 807
rect 1331 803 1332 807
rect 1332 803 1335 807
rect 1367 810 1371 814
rect 1423 810 1427 814
rect 1479 810 1483 814
rect 1535 810 1539 814
rect 1607 819 1608 823
rect 1608 819 1611 823
rect 1591 810 1595 814
rect 1663 808 1667 812
rect 111 776 115 780
rect 151 779 152 783
rect 152 779 155 783
rect 307 779 311 783
rect 351 783 355 787
rect 535 779 539 783
rect 859 791 863 795
rect 967 779 968 783
rect 968 779 971 783
rect 1375 779 1376 783
rect 1376 779 1379 783
rect 135 774 139 778
rect 175 774 179 778
rect 231 774 235 778
rect 295 774 299 778
rect 367 774 371 778
rect 447 774 451 778
rect 527 774 531 778
rect 615 774 619 778
rect 703 774 707 778
rect 791 774 795 778
rect 871 774 875 778
rect 951 774 955 778
rect 1023 774 1027 778
rect 1095 774 1099 778
rect 1167 774 1171 778
rect 1231 774 1235 778
rect 1295 774 1299 778
rect 1359 774 1363 778
rect 1415 774 1419 778
rect 1471 774 1475 778
rect 1527 774 1531 778
rect 1591 774 1595 778
rect 111 759 115 763
rect 287 763 291 767
rect 351 763 355 767
rect 135 757 139 761
rect 175 757 179 761
rect 231 757 235 761
rect 295 757 299 761
rect 367 757 371 761
rect 447 757 451 761
rect 151 751 155 755
rect 687 763 691 767
rect 883 763 887 767
rect 1307 763 1311 767
rect 1511 763 1515 767
rect 1607 779 1608 783
rect 1608 779 1611 783
rect 1663 776 1667 780
rect 527 757 531 761
rect 615 757 619 761
rect 703 757 707 761
rect 791 757 795 761
rect 871 757 875 761
rect 951 757 955 761
rect 1023 757 1027 761
rect 1095 757 1099 761
rect 1167 757 1171 761
rect 1231 757 1235 761
rect 1295 757 1299 761
rect 1359 757 1363 761
rect 1415 757 1419 761
rect 1471 757 1475 761
rect 1527 757 1531 761
rect 967 751 971 755
rect 111 741 115 745
rect 215 743 219 747
rect 247 743 251 747
rect 279 743 283 747
rect 111 724 115 728
rect 215 726 219 730
rect 247 726 251 730
rect 307 739 311 743
rect 319 743 323 747
rect 359 743 363 747
rect 399 743 403 747
rect 439 743 443 747
rect 487 743 491 747
rect 543 743 547 747
rect 607 743 611 747
rect 671 743 675 747
rect 735 743 739 747
rect 799 743 803 747
rect 863 743 867 747
rect 927 743 931 747
rect 991 743 995 747
rect 1055 743 1059 747
rect 1119 743 1123 747
rect 279 726 283 730
rect 331 735 335 739
rect 319 726 323 730
rect 359 726 363 730
rect 331 711 335 715
rect 367 719 371 723
rect 415 735 416 739
rect 416 735 419 739
rect 399 726 403 730
rect 439 726 443 730
rect 487 726 491 730
rect 543 726 547 730
rect 607 726 611 730
rect 775 735 779 739
rect 671 726 675 730
rect 735 726 739 730
rect 687 719 688 723
rect 688 719 691 723
rect 799 726 803 730
rect 863 726 867 730
rect 927 726 931 730
rect 883 719 884 723
rect 884 719 887 723
rect 975 719 979 723
rect 991 726 995 730
rect 1055 726 1059 730
rect 1375 751 1379 755
rect 1591 757 1595 761
rect 1663 759 1667 763
rect 1183 743 1187 747
rect 1239 743 1243 747
rect 1295 743 1299 747
rect 1351 743 1355 747
rect 1407 743 1411 747
rect 1463 743 1467 747
rect 1519 743 1523 747
rect 1583 743 1587 747
rect 1623 743 1627 747
rect 1663 741 1667 745
rect 1119 726 1123 730
rect 1183 726 1187 730
rect 1239 726 1243 730
rect 1295 726 1299 730
rect 1351 726 1355 730
rect 1407 726 1411 730
rect 1463 726 1467 730
rect 1519 726 1523 730
rect 1583 726 1587 730
rect 1623 726 1627 730
rect 1511 719 1515 723
rect 1547 719 1551 723
rect 1639 735 1640 739
rect 1640 735 1643 739
rect 1663 724 1667 728
rect 415 711 419 715
rect 111 692 115 696
rect 391 703 395 707
rect 279 690 283 694
rect 311 690 315 694
rect 343 690 347 694
rect 375 690 379 694
rect 407 690 411 694
rect 439 690 443 694
rect 471 690 475 694
rect 111 675 115 679
rect 360 679 364 683
rect 391 679 392 683
rect 392 679 395 683
rect 279 673 283 677
rect 311 673 315 677
rect 343 673 347 677
rect 375 673 379 677
rect 407 673 411 677
rect 439 673 443 677
rect 775 695 776 699
rect 776 695 779 699
rect 1103 707 1107 711
rect 1031 695 1035 699
rect 1487 695 1488 699
rect 1488 695 1491 699
rect 1639 707 1643 711
rect 503 690 507 694
rect 543 690 547 694
rect 591 690 595 694
rect 647 690 651 694
rect 703 690 707 694
rect 759 690 763 694
rect 823 690 827 694
rect 887 690 891 694
rect 959 690 963 694
rect 1023 690 1027 694
rect 1087 690 1091 694
rect 1159 690 1163 694
rect 1223 690 1227 694
rect 1287 690 1291 694
rect 1351 690 1355 694
rect 1415 690 1419 694
rect 1471 690 1475 694
rect 1527 690 1531 694
rect 1583 690 1587 694
rect 1623 690 1627 694
rect 1663 692 1667 696
rect 471 673 475 677
rect 503 673 507 677
rect 543 673 547 677
rect 591 673 595 677
rect 647 673 651 677
rect 703 673 707 677
rect 111 657 115 661
rect 295 659 299 663
rect 327 659 331 663
rect 359 659 363 663
rect 391 659 395 663
rect 423 659 427 663
rect 455 659 459 663
rect 487 659 491 663
rect 535 667 539 671
rect 927 679 931 683
rect 975 679 976 683
rect 976 679 979 683
rect 1103 679 1104 683
rect 1104 679 1107 683
rect 1427 679 1431 683
rect 1547 679 1548 683
rect 1548 679 1551 683
rect 1639 679 1640 683
rect 1640 679 1643 683
rect 759 673 763 677
rect 823 673 827 677
rect 887 673 891 677
rect 959 673 963 677
rect 1023 673 1027 677
rect 1087 673 1091 677
rect 1159 673 1163 677
rect 1223 673 1227 677
rect 1287 673 1291 677
rect 1351 673 1355 677
rect 1415 673 1419 677
rect 1471 673 1475 677
rect 1527 673 1531 677
rect 1583 673 1587 677
rect 1623 673 1627 677
rect 1663 675 1667 679
rect 519 659 523 663
rect 551 659 555 663
rect 591 659 595 663
rect 639 659 643 663
rect 687 659 691 663
rect 735 659 739 663
rect 791 659 795 663
rect 847 659 851 663
rect 911 659 915 663
rect 975 659 979 663
rect 1047 659 1051 663
rect 1127 659 1131 663
rect 1215 659 1219 663
rect 1295 659 1299 663
rect 1383 659 1387 663
rect 1471 659 1475 663
rect 1559 659 1563 663
rect 1623 659 1627 663
rect 1663 657 1667 661
rect 111 640 115 644
rect 295 642 299 646
rect 327 642 331 646
rect 359 642 363 646
rect 391 642 395 646
rect 423 642 427 646
rect 455 642 459 646
rect 487 642 491 646
rect 519 642 523 646
rect 551 642 555 646
rect 535 635 536 639
rect 536 635 539 639
rect 591 642 595 646
rect 639 642 643 646
rect 687 642 691 646
rect 735 642 739 646
rect 751 651 752 655
rect 752 651 755 655
rect 839 651 843 655
rect 791 642 795 646
rect 847 642 851 646
rect 1031 651 1035 655
rect 911 642 915 646
rect 975 642 979 646
rect 927 635 928 639
rect 928 635 931 639
rect 1047 642 1051 646
rect 1227 651 1231 655
rect 1127 642 1131 646
rect 1215 642 1219 646
rect 1143 635 1144 639
rect 1144 635 1147 639
rect 1295 642 1299 646
rect 1487 651 1488 655
rect 1488 651 1491 655
rect 1383 642 1387 646
rect 1471 642 1475 646
rect 1427 635 1431 639
rect 1559 642 1563 646
rect 1623 642 1627 646
rect 1663 640 1667 644
rect 1591 635 1595 639
rect 1639 635 1640 639
rect 1640 635 1643 639
rect 479 627 483 631
rect 111 612 115 616
rect 263 615 264 619
rect 264 615 267 619
rect 247 610 251 614
rect 279 610 283 614
rect 751 627 755 631
rect 839 615 843 619
rect 1227 615 1228 619
rect 1228 615 1231 619
rect 1235 619 1239 623
rect 1375 615 1376 619
rect 1376 615 1379 619
rect 319 610 323 614
rect 367 610 371 614
rect 423 610 427 614
rect 471 610 475 614
rect 519 610 523 614
rect 567 610 571 614
rect 615 610 619 614
rect 663 610 667 614
rect 719 610 723 614
rect 775 610 779 614
rect 831 610 835 614
rect 895 610 899 614
rect 967 610 971 614
rect 1047 610 1051 614
rect 1119 611 1123 615
rect 1127 610 1131 614
rect 1207 610 1211 614
rect 1287 610 1291 614
rect 1359 610 1363 614
rect 1431 610 1435 614
rect 1503 610 1507 614
rect 1575 610 1579 614
rect 1623 610 1627 614
rect 1663 612 1667 616
rect 111 595 115 599
rect 483 599 487 603
rect 247 593 251 597
rect 279 593 283 597
rect 319 593 323 597
rect 367 593 371 597
rect 423 593 427 597
rect 471 593 475 597
rect 519 593 523 597
rect 567 593 571 597
rect 615 593 619 597
rect 663 593 667 597
rect 719 593 723 597
rect 775 593 779 597
rect 263 587 267 591
rect 111 577 115 581
rect 167 579 171 583
rect 215 579 219 583
rect 271 579 275 583
rect 335 579 339 583
rect 407 579 411 583
rect 111 560 115 564
rect 167 562 171 566
rect 215 562 219 566
rect 271 562 275 566
rect 335 562 339 566
rect 579 587 583 591
rect 979 599 983 603
rect 1143 599 1144 603
rect 1144 599 1147 603
rect 1235 599 1239 603
rect 1299 599 1303 603
rect 1591 599 1592 603
rect 1592 599 1595 603
rect 1639 599 1640 603
rect 1640 599 1643 603
rect 831 593 835 597
rect 895 593 899 597
rect 967 593 971 597
rect 1047 593 1051 597
rect 1127 593 1131 597
rect 1207 593 1211 597
rect 1287 593 1291 597
rect 1359 593 1363 597
rect 1431 593 1435 597
rect 1503 593 1507 597
rect 1575 593 1579 597
rect 1623 593 1627 597
rect 1663 595 1667 599
rect 1375 587 1379 591
rect 487 579 491 583
rect 559 579 563 583
rect 631 579 635 583
rect 703 579 707 583
rect 767 579 771 583
rect 823 579 827 583
rect 879 579 883 583
rect 935 579 939 583
rect 991 579 995 583
rect 1047 579 1051 583
rect 1103 579 1107 583
rect 1159 579 1163 583
rect 1215 579 1219 583
rect 1271 579 1275 583
rect 1327 579 1331 583
rect 1383 579 1387 583
rect 1447 579 1451 583
rect 1511 579 1515 583
rect 407 562 411 566
rect 487 562 491 566
rect 559 562 563 566
rect 579 555 580 559
rect 580 555 583 559
rect 631 562 635 566
rect 703 562 707 566
rect 807 571 811 575
rect 767 562 771 566
rect 823 562 827 566
rect 895 571 896 575
rect 896 571 899 575
rect 879 562 883 566
rect 935 562 939 566
rect 991 562 995 566
rect 343 547 347 551
rect 979 555 983 559
rect 1023 555 1027 559
rect 1047 562 1051 566
rect 1119 571 1120 575
rect 1120 571 1123 575
rect 1199 571 1203 575
rect 1103 562 1107 566
rect 1159 562 1163 566
rect 1215 562 1219 566
rect 1271 562 1275 566
rect 1327 562 1331 566
rect 1383 562 1387 566
rect 1299 555 1303 559
rect 1447 562 1451 566
rect 1511 562 1515 566
rect 1575 579 1579 583
rect 1623 579 1627 583
rect 1663 577 1667 581
rect 1575 562 1579 566
rect 1623 562 1627 566
rect 1663 560 1667 564
rect 1639 555 1640 559
rect 1640 555 1643 559
rect 111 528 115 532
rect 151 531 152 535
rect 152 531 155 535
rect 135 526 139 530
rect 111 511 115 515
rect 167 526 171 530
rect 199 526 203 530
rect 511 543 515 547
rect 231 526 235 530
rect 279 526 283 530
rect 327 526 331 530
rect 375 526 379 530
rect 431 526 435 530
rect 495 526 499 530
rect 639 539 643 543
rect 831 543 835 547
rect 1527 547 1531 551
rect 631 531 635 535
rect 807 535 811 539
rect 895 531 896 535
rect 896 531 899 535
rect 559 526 563 530
rect 623 526 627 530
rect 687 526 691 530
rect 751 526 755 530
rect 815 526 819 530
rect 879 526 883 530
rect 943 526 947 530
rect 1007 526 1011 530
rect 1071 526 1075 530
rect 1127 526 1131 530
rect 343 515 344 519
rect 344 515 347 519
rect 487 515 491 519
rect 511 515 512 519
rect 512 515 515 519
rect 639 515 640 519
rect 640 515 643 519
rect 791 515 795 519
rect 831 515 832 519
rect 832 515 835 519
rect 1023 515 1024 519
rect 1024 515 1027 519
rect 135 509 139 513
rect 167 509 171 513
rect 199 509 203 513
rect 231 509 235 513
rect 279 509 283 513
rect 327 509 331 513
rect 375 509 379 513
rect 431 509 435 513
rect 495 509 499 513
rect 559 509 563 513
rect 623 509 627 513
rect 687 509 691 513
rect 751 509 755 513
rect 815 509 819 513
rect 879 509 883 513
rect 943 509 947 513
rect 1007 509 1011 513
rect 1071 509 1075 513
rect 151 503 155 507
rect 111 493 115 497
rect 135 495 139 499
rect 167 495 171 499
rect 199 495 203 499
rect 239 495 243 499
rect 111 476 115 480
rect 135 478 139 482
rect 167 478 171 482
rect 199 478 203 482
rect 951 503 955 507
rect 1183 526 1187 530
rect 1199 531 1200 535
rect 1200 531 1203 535
rect 1247 531 1248 535
rect 1248 531 1251 535
rect 1231 526 1235 530
rect 1279 526 1283 530
rect 1335 526 1339 530
rect 1391 526 1395 530
rect 1447 526 1451 530
rect 1511 526 1515 530
rect 1575 526 1579 530
rect 1623 526 1627 530
rect 1663 528 1667 532
rect 1527 515 1528 519
rect 1528 515 1531 519
rect 1607 515 1611 519
rect 1127 509 1131 513
rect 1183 509 1187 513
rect 1231 509 1235 513
rect 1279 509 1283 513
rect 1335 509 1339 513
rect 1391 509 1395 513
rect 1447 509 1451 513
rect 1511 509 1515 513
rect 1575 509 1579 513
rect 1623 509 1627 513
rect 1663 511 1667 515
rect 1247 503 1251 507
rect 287 495 291 499
rect 327 495 331 499
rect 375 495 379 499
rect 423 495 427 499
rect 479 495 483 499
rect 543 495 547 499
rect 615 495 619 499
rect 695 495 699 499
rect 775 495 779 499
rect 847 495 851 499
rect 919 495 923 499
rect 983 495 987 499
rect 1039 495 1043 499
rect 1095 495 1099 499
rect 1143 495 1147 499
rect 1191 495 1195 499
rect 1239 495 1243 499
rect 1287 495 1291 499
rect 1335 495 1339 499
rect 1383 495 1387 499
rect 1431 495 1435 499
rect 1479 495 1483 499
rect 1535 495 1539 499
rect 1591 495 1595 499
rect 1623 495 1627 499
rect 239 478 243 482
rect 287 478 291 482
rect 327 478 331 482
rect 275 471 279 475
rect 375 478 379 482
rect 423 478 427 482
rect 479 478 483 482
rect 543 478 547 482
rect 487 471 491 475
rect 631 487 632 491
rect 632 487 635 491
rect 615 478 619 482
rect 695 478 699 482
rect 775 478 779 482
rect 703 471 707 475
rect 791 471 792 475
rect 792 471 795 475
rect 835 487 839 491
rect 847 478 851 482
rect 919 478 923 482
rect 951 471 955 475
rect 983 478 987 482
rect 1039 478 1043 482
rect 1095 478 1099 482
rect 1143 478 1147 482
rect 1191 478 1195 482
rect 1239 478 1243 482
rect 1287 478 1291 482
rect 1663 493 1667 497
rect 1335 478 1339 482
rect 1383 478 1387 482
rect 1431 478 1435 482
rect 1511 487 1515 491
rect 1519 487 1523 491
rect 1479 478 1483 482
rect 1535 478 1539 482
rect 1591 478 1595 482
rect 1623 478 1627 482
rect 111 448 115 452
rect 191 451 195 455
rect 151 446 155 450
rect 111 431 115 435
rect 999 463 1003 467
rect 831 451 835 455
rect 1391 463 1395 467
rect 1519 463 1523 467
rect 1607 471 1608 475
rect 1608 471 1611 475
rect 1639 487 1640 491
rect 1640 487 1643 491
rect 1663 476 1667 480
rect 1639 463 1643 467
rect 207 446 211 450
rect 255 446 259 450
rect 311 446 315 450
rect 367 446 371 450
rect 439 446 443 450
rect 519 446 523 450
rect 599 446 603 450
rect 679 446 683 450
rect 759 446 763 450
rect 839 446 843 450
rect 911 446 915 450
rect 983 446 987 450
rect 1055 446 1059 450
rect 1127 446 1131 450
rect 275 435 276 439
rect 276 435 279 439
rect 327 435 328 439
rect 328 435 331 439
rect 696 435 700 439
rect 823 435 827 439
rect 951 435 955 439
rect 999 435 1000 439
rect 1000 435 1003 439
rect 1199 446 1203 450
rect 1215 451 1216 455
rect 1216 451 1219 455
rect 1263 446 1267 450
rect 1319 446 1323 450
rect 1375 446 1379 450
rect 1431 446 1435 450
rect 1495 446 1499 450
rect 1351 435 1355 439
rect 1391 435 1392 439
rect 1392 435 1395 439
rect 1511 451 1512 455
rect 1512 451 1515 455
rect 1663 448 1667 452
rect 151 429 155 433
rect 207 429 211 433
rect 255 429 259 433
rect 311 429 315 433
rect 367 429 371 433
rect 439 429 443 433
rect 519 429 523 433
rect 599 429 603 433
rect 679 429 683 433
rect 759 429 763 433
rect 839 429 843 433
rect 911 429 915 433
rect 983 429 987 433
rect 1055 429 1059 433
rect 1127 429 1131 433
rect 1199 429 1203 433
rect 1263 429 1267 433
rect 1319 429 1323 433
rect 1375 429 1379 433
rect 1431 429 1435 433
rect 1495 429 1499 433
rect 1663 431 1667 435
rect 111 413 115 417
rect 175 415 179 419
rect 223 415 227 419
rect 271 415 275 419
rect 319 415 323 419
rect 367 415 371 419
rect 415 415 419 419
rect 471 415 475 419
rect 527 415 531 419
rect 591 415 595 419
rect 663 415 667 419
rect 735 415 739 419
rect 807 415 811 419
rect 871 415 875 419
rect 935 415 939 419
rect 991 415 995 419
rect 1039 415 1043 419
rect 1087 415 1091 419
rect 1127 415 1131 419
rect 191 407 192 411
rect 192 407 195 411
rect 111 396 115 400
rect 175 398 179 402
rect 223 398 227 402
rect 271 398 275 402
rect 319 398 323 402
rect 231 391 235 395
rect 327 391 331 395
rect 367 398 371 402
rect 427 407 431 411
rect 415 398 419 402
rect 471 398 475 402
rect 527 398 531 402
rect 591 398 595 402
rect 755 407 756 411
rect 756 407 759 411
rect 663 398 667 402
rect 735 398 739 402
rect 671 391 675 395
rect 883 407 887 411
rect 807 398 811 402
rect 871 398 875 402
rect 935 398 939 402
rect 823 391 824 395
rect 824 391 827 395
rect 951 391 952 395
rect 952 391 955 395
rect 1003 407 1007 411
rect 991 398 995 402
rect 1039 398 1043 402
rect 1087 398 1091 402
rect 111 364 115 368
rect 151 367 152 371
rect 152 367 155 371
rect 135 362 139 366
rect 111 347 115 351
rect 167 362 171 366
rect 199 362 203 366
rect 239 362 243 366
rect 295 362 299 366
rect 231 351 235 355
rect 251 351 255 355
rect 351 362 355 366
rect 407 362 411 366
rect 427 367 428 371
rect 428 367 431 371
rect 475 367 479 371
rect 815 379 819 383
rect 1003 383 1007 387
rect 1215 423 1219 427
rect 1167 415 1171 419
rect 1207 415 1211 419
rect 1247 415 1251 419
rect 1287 415 1291 419
rect 1335 415 1339 419
rect 1383 415 1387 419
rect 1663 413 1667 417
rect 1127 398 1131 402
rect 1167 398 1171 402
rect 1207 398 1211 402
rect 1247 398 1251 402
rect 1287 398 1291 402
rect 1335 398 1339 402
rect 1383 398 1387 402
rect 1111 383 1115 387
rect 1351 391 1352 395
rect 1352 391 1355 395
rect 1663 396 1667 400
rect 755 367 759 371
rect 883 367 887 371
rect 891 371 895 375
rect 1159 367 1163 371
rect 1239 371 1243 375
rect 1439 371 1443 375
rect 463 362 467 366
rect 519 362 523 366
rect 575 362 579 366
rect 631 362 635 366
rect 687 362 691 366
rect 743 362 747 366
rect 799 362 803 366
rect 855 362 859 366
rect 919 362 923 366
rect 983 362 987 366
rect 1039 362 1043 366
rect 1095 362 1099 366
rect 1151 362 1155 366
rect 1207 362 1211 366
rect 1255 362 1259 366
rect 1303 362 1307 366
rect 1351 362 1355 366
rect 1399 362 1403 366
rect 1447 362 1451 366
rect 1495 362 1499 366
rect 1535 363 1539 367
rect 1543 362 1547 366
rect 1591 362 1595 366
rect 671 351 675 355
rect 699 351 703 355
rect 815 351 816 355
rect 816 351 819 355
rect 891 351 895 355
rect 1051 351 1055 355
rect 1111 351 1112 355
rect 1112 351 1115 355
rect 1239 351 1243 355
rect 1439 351 1443 355
rect 1623 362 1627 366
rect 1663 364 1667 368
rect 1639 351 1640 355
rect 1640 351 1643 355
rect 135 345 139 349
rect 167 345 171 349
rect 199 345 203 349
rect 239 345 243 349
rect 295 345 299 349
rect 351 345 355 349
rect 407 345 411 349
rect 463 345 467 349
rect 519 345 523 349
rect 575 345 579 349
rect 631 345 635 349
rect 687 345 691 349
rect 743 345 747 349
rect 799 345 803 349
rect 855 345 859 349
rect 919 345 923 349
rect 983 345 987 349
rect 1039 345 1043 349
rect 1095 345 1099 349
rect 1151 345 1155 349
rect 1207 345 1211 349
rect 1255 345 1259 349
rect 1303 345 1307 349
rect 1351 345 1355 349
rect 1399 345 1403 349
rect 1447 345 1451 349
rect 151 339 155 343
rect 111 329 115 333
rect 135 331 139 335
rect 167 331 171 335
rect 1495 345 1499 349
rect 1543 345 1547 349
rect 1591 345 1595 349
rect 1623 345 1627 349
rect 1663 347 1667 351
rect 207 331 211 335
rect 263 331 267 335
rect 327 331 331 335
rect 391 331 395 335
rect 455 331 459 335
rect 519 331 523 335
rect 575 331 579 335
rect 631 331 635 335
rect 687 331 691 335
rect 751 331 755 335
rect 815 331 819 335
rect 879 331 883 335
rect 951 331 955 335
rect 1031 331 1035 335
rect 1111 331 1115 335
rect 1191 331 1195 335
rect 1271 331 1275 335
rect 1343 331 1347 335
rect 1407 331 1411 335
rect 1463 331 1467 335
rect 1519 331 1523 335
rect 1535 331 1539 335
rect 111 312 115 316
rect 135 314 139 318
rect 167 314 171 318
rect 151 307 152 311
rect 152 307 155 311
rect 207 314 211 318
rect 263 314 267 318
rect 251 307 255 311
rect 447 323 451 327
rect 475 323 476 327
rect 476 323 479 327
rect 327 314 331 318
rect 391 314 395 318
rect 455 314 459 318
rect 587 323 591 327
rect 519 314 523 318
rect 575 314 579 318
rect 631 314 635 318
rect 687 314 691 318
rect 695 307 699 311
rect 751 314 755 318
rect 815 314 819 318
rect 879 314 883 318
rect 951 314 955 318
rect 1159 323 1163 327
rect 1031 314 1035 318
rect 1111 314 1115 318
rect 1051 307 1052 311
rect 1052 307 1055 311
rect 1191 314 1195 318
rect 1271 314 1275 318
rect 1343 314 1347 318
rect 1283 307 1287 311
rect 1407 314 1411 318
rect 1583 331 1587 335
rect 1623 331 1627 335
rect 1663 329 1667 333
rect 1463 314 1467 318
rect 1519 314 1523 318
rect 1583 314 1587 318
rect 1623 314 1627 318
rect 1663 312 1667 316
rect 1639 307 1640 311
rect 1640 307 1643 311
rect 247 295 251 299
rect 707 299 711 303
rect 111 284 115 288
rect 135 282 139 286
rect 167 282 171 286
rect 111 267 115 271
rect 151 271 152 275
rect 152 271 155 275
rect 239 287 243 291
rect 231 282 235 286
rect 295 282 299 286
rect 367 282 371 286
rect 247 271 248 275
rect 248 271 251 275
rect 307 271 311 275
rect 447 287 451 291
rect 439 282 443 286
rect 503 282 507 286
rect 587 287 588 291
rect 588 287 591 291
rect 679 287 683 291
rect 567 282 571 286
rect 631 282 635 286
rect 687 282 691 286
rect 1127 287 1128 291
rect 1128 287 1131 291
rect 1343 287 1344 291
rect 1344 287 1347 291
rect 743 282 747 286
rect 807 282 811 286
rect 879 282 883 286
rect 951 282 955 286
rect 1031 282 1035 286
rect 1111 282 1115 286
rect 1191 282 1195 286
rect 1263 282 1267 286
rect 1327 282 1331 286
rect 1391 282 1395 286
rect 1447 282 1451 286
rect 1495 282 1499 286
rect 535 271 539 275
rect 707 271 708 275
rect 708 271 711 275
rect 1283 271 1284 275
rect 1284 271 1287 275
rect 1431 271 1435 275
rect 135 265 139 269
rect 167 265 171 269
rect 231 265 235 269
rect 295 265 299 269
rect 367 265 371 269
rect 439 265 443 269
rect 503 265 507 269
rect 567 265 571 269
rect 631 265 635 269
rect 687 265 691 269
rect 743 265 747 269
rect 807 265 811 269
rect 879 265 883 269
rect 951 265 955 269
rect 1031 265 1035 269
rect 915 259 919 263
rect 1111 265 1115 269
rect 1191 265 1195 269
rect 1263 265 1267 269
rect 1327 265 1331 269
rect 1391 265 1395 269
rect 1447 265 1451 269
rect 1127 255 1131 259
rect 1343 259 1347 263
rect 1543 282 1547 286
rect 1591 282 1595 286
rect 1623 282 1627 286
rect 1663 284 1667 288
rect 1495 265 1499 269
rect 1543 265 1547 269
rect 1591 265 1595 269
rect 1623 265 1627 269
rect 1663 267 1667 271
rect 111 245 115 249
rect 135 247 139 251
rect 175 247 179 251
rect 247 247 251 251
rect 319 247 323 251
rect 383 247 387 251
rect 447 247 451 251
rect 519 247 523 251
rect 591 247 595 251
rect 663 247 667 251
rect 743 247 747 251
rect 823 247 827 251
rect 895 247 899 251
rect 967 247 971 251
rect 1031 247 1035 251
rect 1087 247 1091 251
rect 1143 247 1147 251
rect 1199 247 1203 251
rect 111 228 115 232
rect 135 230 139 234
rect 175 230 179 234
rect 151 223 152 227
rect 152 223 155 227
rect 239 239 243 243
rect 247 230 251 234
rect 319 230 323 234
rect 307 223 311 227
rect 383 230 387 234
rect 439 239 443 243
rect 575 239 579 243
rect 679 239 680 243
rect 680 239 683 243
rect 447 230 451 234
rect 519 230 523 234
rect 535 223 536 227
rect 536 223 539 227
rect 591 230 595 234
rect 663 230 667 234
rect 743 230 747 234
rect 823 230 827 234
rect 895 230 899 234
rect 967 230 971 234
rect 915 223 916 227
rect 916 223 919 227
rect 1031 230 1035 234
rect 1087 230 1091 234
rect 111 200 115 204
rect 135 198 139 202
rect 167 198 171 202
rect 111 183 115 187
rect 151 187 152 191
rect 152 187 155 191
rect 207 198 211 202
rect 247 203 251 207
rect 255 198 259 202
rect 303 198 307 202
rect 295 187 299 191
rect 439 215 443 219
rect 1143 230 1147 234
rect 1255 247 1259 251
rect 1311 247 1315 251
rect 1367 247 1371 251
rect 1415 247 1419 251
rect 1463 247 1467 251
rect 1519 247 1523 251
rect 1575 247 1579 251
rect 1623 247 1627 251
rect 1663 245 1667 249
rect 1199 230 1203 234
rect 1323 239 1327 243
rect 1255 230 1259 234
rect 1311 230 1315 234
rect 1367 230 1371 234
rect 1415 230 1419 234
rect 1463 230 1467 234
rect 1519 230 1523 234
rect 1431 223 1432 227
rect 1432 223 1435 227
rect 1483 223 1484 227
rect 1484 223 1487 227
rect 1575 230 1579 234
rect 1635 239 1639 243
rect 1623 230 1627 234
rect 1663 228 1667 232
rect 391 203 392 207
rect 392 203 395 207
rect 491 211 495 215
rect 1231 215 1235 219
rect 575 203 579 207
rect 871 203 872 207
rect 872 203 875 207
rect 1323 203 1327 207
rect 1331 207 1335 211
rect 1435 203 1436 207
rect 1436 203 1439 207
rect 1455 207 1459 211
rect 1635 215 1639 219
rect 343 198 347 202
rect 375 198 379 202
rect 415 198 419 202
rect 471 198 475 202
rect 535 198 539 202
rect 615 198 619 202
rect 695 198 699 202
rect 775 198 779 202
rect 855 198 859 202
rect 927 198 931 202
rect 999 198 1003 202
rect 1071 198 1075 202
rect 1143 198 1147 202
rect 1215 198 1219 202
rect 1287 198 1291 202
rect 1351 198 1355 202
rect 1415 198 1419 202
rect 1471 198 1475 202
rect 1527 198 1531 202
rect 1583 198 1587 202
rect 1623 198 1627 202
rect 1663 200 1667 204
rect 491 187 492 191
rect 492 187 495 191
rect 135 181 139 185
rect 167 181 171 185
rect 207 181 211 185
rect 255 181 259 185
rect 303 181 307 185
rect 343 181 347 185
rect 375 181 379 185
rect 415 181 419 185
rect 471 181 475 185
rect 535 181 539 185
rect 391 175 395 179
rect 787 187 791 191
rect 1231 187 1232 191
rect 1232 187 1235 191
rect 1331 187 1335 191
rect 1367 187 1368 191
rect 1368 187 1371 191
rect 1455 187 1459 191
rect 1483 187 1487 191
rect 1639 187 1640 191
rect 1640 187 1643 191
rect 615 181 619 185
rect 695 181 699 185
rect 775 181 779 185
rect 855 181 859 185
rect 927 181 931 185
rect 999 181 1003 185
rect 1071 181 1075 185
rect 1143 181 1147 185
rect 1215 181 1219 185
rect 1287 181 1291 185
rect 1351 181 1355 185
rect 1415 181 1419 185
rect 1471 181 1475 185
rect 1527 181 1531 185
rect 1583 181 1587 185
rect 1623 181 1627 185
rect 1663 183 1667 187
rect 871 175 875 179
rect 111 165 115 169
rect 135 167 139 171
rect 175 167 179 171
rect 231 167 235 171
rect 287 167 291 171
rect 343 167 347 171
rect 399 167 403 171
rect 455 167 459 171
rect 511 167 515 171
rect 575 167 579 171
rect 639 167 643 171
rect 703 167 707 171
rect 767 167 771 171
rect 831 167 835 171
rect 895 167 899 171
rect 951 167 955 171
rect 1015 167 1019 171
rect 1079 167 1083 171
rect 1143 167 1147 171
rect 1207 167 1211 171
rect 1279 167 1283 171
rect 1351 167 1355 171
rect 1423 167 1427 171
rect 1495 167 1499 171
rect 1567 167 1571 171
rect 1623 167 1627 171
rect 1663 165 1667 169
rect 111 148 115 152
rect 135 150 139 154
rect 175 150 179 154
rect 151 143 152 147
rect 152 143 155 147
rect 247 159 248 163
rect 248 159 251 163
rect 231 150 235 154
rect 287 150 291 154
rect 295 143 299 147
rect 343 150 347 154
rect 439 159 443 163
rect 399 150 403 154
rect 455 150 459 154
rect 511 150 515 154
rect 575 150 579 154
rect 639 150 643 154
rect 703 150 707 154
rect 759 159 763 163
rect 767 150 771 154
rect 831 150 835 154
rect 895 150 899 154
rect 787 135 791 139
rect 951 150 955 154
rect 1015 150 1019 154
rect 1079 150 1083 154
rect 1199 159 1203 163
rect 1143 150 1147 154
rect 1207 150 1211 154
rect 1279 150 1283 154
rect 1435 159 1439 163
rect 1351 150 1355 154
rect 1423 150 1427 154
rect 1367 143 1368 147
rect 1368 143 1371 147
rect 1495 150 1499 154
rect 1567 150 1571 154
rect 1623 150 1627 154
rect 1663 148 1667 152
rect 1575 143 1579 147
rect 1639 143 1640 147
rect 1640 143 1643 147
rect 1159 135 1163 139
rect 479 127 483 131
rect 759 127 763 131
rect 111 104 115 108
rect 135 102 139 106
rect 167 102 171 106
rect 111 87 115 91
rect 151 91 152 95
rect 152 91 155 95
rect 199 102 203 106
rect 231 102 235 106
rect 263 102 267 106
rect 295 102 299 106
rect 327 102 331 106
rect 359 102 363 106
rect 391 102 395 106
rect 423 102 427 106
rect 439 107 440 111
rect 440 107 443 111
rect 479 107 480 111
rect 480 107 483 111
rect 463 102 467 106
rect 503 102 507 106
rect 543 102 547 106
rect 575 102 579 106
rect 607 102 611 106
rect 639 102 643 106
rect 671 102 675 106
rect 703 102 707 106
rect 735 102 739 106
rect 767 102 771 106
rect 799 102 803 106
rect 831 102 835 106
rect 863 102 867 106
rect 895 102 899 106
rect 1199 107 1200 111
rect 1200 107 1203 111
rect 935 102 939 106
rect 975 102 979 106
rect 1015 102 1019 106
rect 1063 102 1067 106
rect 1103 102 1107 106
rect 1143 102 1147 106
rect 1183 102 1187 106
rect 1223 102 1227 106
rect 1263 102 1267 106
rect 1295 102 1299 106
rect 1335 102 1339 106
rect 1375 102 1379 106
rect 1415 102 1419 106
rect 1455 102 1459 106
rect 1503 102 1507 106
rect 1551 102 1555 106
rect 1591 102 1595 106
rect 1623 102 1627 106
rect 1159 91 1160 95
rect 1160 91 1163 95
rect 1568 91 1572 95
rect 1663 104 1667 108
rect 135 85 139 89
rect 167 85 171 89
rect 199 85 203 89
rect 231 85 235 89
rect 263 85 267 89
rect 295 85 299 89
rect 327 85 331 89
rect 359 85 363 89
rect 391 85 395 89
rect 423 85 427 89
rect 463 85 467 89
rect 503 85 507 89
rect 543 85 547 89
rect 575 85 579 89
rect 607 85 611 89
rect 639 85 643 89
rect 671 85 675 89
rect 703 85 707 89
rect 735 85 739 89
rect 767 85 771 89
rect 799 85 803 89
rect 831 85 835 89
rect 863 85 867 89
rect 895 85 899 89
rect 935 85 939 89
rect 975 85 979 89
rect 1015 85 1019 89
rect 1063 85 1067 89
rect 1103 85 1107 89
rect 1143 85 1147 89
rect 1183 85 1187 89
rect 1223 85 1227 89
rect 1263 85 1267 89
rect 1295 85 1299 89
rect 1335 85 1339 89
rect 1375 85 1379 89
rect 1415 85 1419 89
rect 1455 85 1459 89
rect 1503 85 1507 89
rect 1551 85 1555 89
rect 1591 85 1595 89
rect 1623 85 1627 89
rect 1663 87 1667 91
<< m3 >>
rect 111 1718 115 1719
rect 111 1713 115 1714
rect 255 1718 259 1719
rect 255 1713 259 1714
rect 287 1718 291 1719
rect 287 1713 291 1714
rect 319 1718 323 1719
rect 319 1713 323 1714
rect 359 1718 363 1719
rect 407 1718 411 1719
rect 359 1713 363 1714
rect 374 1715 380 1716
rect 112 1705 114 1713
rect 110 1704 116 1705
rect 110 1700 111 1704
rect 115 1700 116 1704
rect 256 1703 258 1713
rect 288 1703 290 1713
rect 320 1703 322 1713
rect 360 1703 362 1713
rect 374 1711 375 1715
rect 379 1711 380 1715
rect 407 1713 411 1714
rect 455 1718 459 1719
rect 455 1713 459 1714
rect 503 1718 507 1719
rect 503 1713 507 1714
rect 551 1718 555 1719
rect 551 1713 555 1714
rect 607 1718 611 1719
rect 607 1713 611 1714
rect 663 1718 667 1719
rect 663 1713 667 1714
rect 727 1718 731 1719
rect 727 1713 731 1714
rect 783 1718 787 1719
rect 783 1713 787 1714
rect 839 1718 843 1719
rect 839 1713 843 1714
rect 895 1718 899 1719
rect 895 1713 899 1714
rect 951 1718 955 1719
rect 951 1713 955 1714
rect 1007 1718 1011 1719
rect 1007 1713 1011 1714
rect 1063 1718 1067 1719
rect 1063 1713 1067 1714
rect 1119 1718 1123 1719
rect 1175 1718 1179 1719
rect 1119 1713 1123 1714
rect 1138 1715 1144 1716
rect 374 1710 380 1711
rect 110 1699 116 1700
rect 254 1702 260 1703
rect 254 1698 255 1702
rect 259 1698 260 1702
rect 254 1697 260 1698
rect 286 1702 292 1703
rect 286 1698 287 1702
rect 291 1698 292 1702
rect 286 1697 292 1698
rect 318 1702 324 1703
rect 318 1698 319 1702
rect 323 1698 324 1702
rect 318 1697 324 1698
rect 358 1702 364 1703
rect 358 1698 359 1702
rect 363 1698 364 1702
rect 358 1697 364 1698
rect 376 1692 378 1710
rect 408 1703 410 1713
rect 456 1703 458 1713
rect 470 1711 476 1712
rect 470 1707 471 1711
rect 475 1707 476 1711
rect 470 1706 476 1707
rect 406 1702 412 1703
rect 406 1698 407 1702
rect 411 1698 412 1702
rect 406 1697 412 1698
rect 454 1702 460 1703
rect 454 1698 455 1702
rect 459 1698 460 1702
rect 454 1697 460 1698
rect 472 1692 474 1706
rect 504 1703 506 1713
rect 538 1711 544 1712
rect 514 1707 520 1708
rect 514 1703 515 1707
rect 519 1703 520 1707
rect 538 1707 539 1711
rect 543 1707 544 1711
rect 538 1706 544 1707
rect 502 1702 508 1703
rect 514 1702 520 1703
rect 502 1698 503 1702
rect 507 1698 508 1702
rect 502 1697 508 1698
rect 350 1691 356 1692
rect 110 1687 116 1688
rect 110 1683 111 1687
rect 115 1683 116 1687
rect 350 1687 351 1691
rect 355 1687 356 1691
rect 350 1686 356 1687
rect 374 1691 380 1692
rect 374 1687 375 1691
rect 379 1687 380 1691
rect 374 1686 380 1687
rect 470 1691 476 1692
rect 470 1687 471 1691
rect 475 1687 476 1691
rect 470 1686 476 1687
rect 110 1682 116 1683
rect 254 1685 260 1686
rect 112 1679 114 1682
rect 254 1681 255 1685
rect 259 1681 260 1685
rect 254 1680 260 1681
rect 286 1685 292 1686
rect 286 1681 287 1685
rect 291 1681 292 1685
rect 286 1680 292 1681
rect 318 1685 324 1686
rect 318 1681 319 1685
rect 323 1681 324 1685
rect 318 1680 324 1681
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 135 1678 139 1679
rect 112 1670 114 1673
rect 135 1672 139 1674
rect 167 1678 171 1679
rect 167 1672 171 1674
rect 215 1678 219 1679
rect 215 1672 219 1674
rect 255 1678 259 1680
rect 255 1673 259 1674
rect 279 1678 283 1679
rect 279 1672 283 1674
rect 287 1678 291 1680
rect 287 1673 291 1674
rect 319 1678 323 1680
rect 319 1673 323 1674
rect 343 1678 347 1679
rect 343 1672 347 1674
rect 134 1671 140 1672
rect 110 1669 116 1670
rect 110 1665 111 1669
rect 115 1665 116 1669
rect 134 1667 135 1671
rect 139 1667 140 1671
rect 134 1666 140 1667
rect 166 1671 172 1672
rect 166 1667 167 1671
rect 171 1667 172 1671
rect 166 1666 172 1667
rect 214 1671 220 1672
rect 214 1667 215 1671
rect 219 1667 220 1671
rect 214 1666 220 1667
rect 278 1671 284 1672
rect 278 1667 279 1671
rect 283 1667 284 1671
rect 278 1666 284 1667
rect 342 1671 348 1672
rect 342 1667 343 1671
rect 347 1667 348 1671
rect 342 1666 348 1667
rect 110 1664 116 1665
rect 150 1663 156 1664
rect 150 1659 151 1663
rect 155 1659 156 1663
rect 150 1658 156 1659
rect 134 1654 140 1655
rect 110 1652 116 1653
rect 110 1648 111 1652
rect 115 1648 116 1652
rect 134 1650 135 1654
rect 139 1650 140 1654
rect 134 1649 140 1650
rect 110 1647 116 1648
rect 112 1639 114 1647
rect 136 1639 138 1649
rect 111 1638 115 1639
rect 111 1633 115 1634
rect 135 1638 139 1639
rect 135 1633 139 1634
rect 112 1625 114 1633
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 136 1623 138 1633
rect 152 1628 154 1658
rect 166 1654 172 1655
rect 166 1650 167 1654
rect 171 1650 172 1654
rect 166 1649 172 1650
rect 214 1654 220 1655
rect 214 1650 215 1654
rect 219 1650 220 1654
rect 214 1649 220 1650
rect 278 1654 284 1655
rect 278 1650 279 1654
rect 283 1650 284 1654
rect 278 1649 284 1650
rect 342 1654 348 1655
rect 342 1650 343 1654
rect 347 1650 348 1654
rect 342 1649 348 1650
rect 168 1639 170 1649
rect 216 1639 218 1649
rect 280 1639 282 1649
rect 344 1639 346 1649
rect 352 1648 354 1686
rect 358 1685 364 1686
rect 358 1681 359 1685
rect 363 1681 364 1685
rect 358 1680 364 1681
rect 406 1685 412 1686
rect 406 1681 407 1685
rect 411 1681 412 1685
rect 406 1680 412 1681
rect 454 1685 460 1686
rect 454 1681 455 1685
rect 459 1681 460 1685
rect 454 1680 460 1681
rect 502 1685 508 1686
rect 502 1681 503 1685
rect 507 1681 508 1685
rect 502 1680 508 1681
rect 359 1678 363 1680
rect 359 1673 363 1674
rect 407 1678 411 1680
rect 407 1673 411 1674
rect 415 1678 419 1679
rect 415 1672 419 1674
rect 455 1678 459 1680
rect 455 1673 459 1674
rect 487 1678 491 1679
rect 487 1672 491 1674
rect 503 1678 507 1680
rect 503 1673 507 1674
rect 414 1671 420 1672
rect 414 1667 415 1671
rect 419 1667 420 1671
rect 414 1666 420 1667
rect 486 1671 492 1672
rect 486 1667 487 1671
rect 491 1667 492 1671
rect 516 1668 518 1702
rect 540 1692 542 1706
rect 552 1703 554 1713
rect 608 1703 610 1713
rect 664 1703 666 1713
rect 728 1703 730 1713
rect 784 1703 786 1713
rect 840 1703 842 1713
rect 886 1707 892 1708
rect 886 1703 887 1707
rect 891 1703 892 1707
rect 896 1703 898 1713
rect 952 1703 954 1713
rect 1008 1703 1010 1713
rect 1064 1703 1066 1713
rect 1106 1711 1112 1712
rect 1106 1707 1107 1711
rect 1111 1707 1112 1711
rect 1106 1706 1112 1707
rect 550 1702 556 1703
rect 550 1698 551 1702
rect 555 1698 556 1702
rect 550 1697 556 1698
rect 606 1702 612 1703
rect 606 1698 607 1702
rect 611 1698 612 1702
rect 606 1697 612 1698
rect 662 1702 668 1703
rect 662 1698 663 1702
rect 667 1698 668 1702
rect 662 1697 668 1698
rect 726 1702 732 1703
rect 726 1698 727 1702
rect 731 1698 732 1702
rect 726 1697 732 1698
rect 782 1702 788 1703
rect 782 1698 783 1702
rect 787 1698 788 1702
rect 782 1697 788 1698
rect 838 1702 844 1703
rect 886 1702 892 1703
rect 894 1702 900 1703
rect 838 1698 839 1702
rect 843 1698 844 1702
rect 838 1697 844 1698
rect 538 1691 544 1692
rect 538 1687 539 1691
rect 543 1687 544 1691
rect 538 1686 544 1687
rect 802 1691 808 1692
rect 802 1687 803 1691
rect 807 1687 808 1691
rect 802 1686 808 1687
rect 550 1685 556 1686
rect 550 1681 551 1685
rect 555 1681 556 1685
rect 550 1680 556 1681
rect 606 1685 612 1686
rect 606 1681 607 1685
rect 611 1681 612 1685
rect 606 1680 612 1681
rect 662 1685 668 1686
rect 662 1681 663 1685
rect 667 1681 668 1685
rect 662 1680 668 1681
rect 726 1685 732 1686
rect 726 1681 727 1685
rect 731 1681 732 1685
rect 726 1680 732 1681
rect 782 1685 788 1686
rect 782 1681 783 1685
rect 787 1681 788 1685
rect 782 1680 788 1681
rect 551 1678 555 1680
rect 551 1673 555 1674
rect 559 1678 563 1679
rect 559 1672 563 1674
rect 607 1678 611 1680
rect 607 1673 611 1674
rect 631 1678 635 1679
rect 631 1672 635 1674
rect 663 1678 667 1680
rect 663 1673 667 1674
rect 711 1678 715 1679
rect 711 1672 715 1674
rect 727 1678 731 1680
rect 727 1673 731 1674
rect 783 1678 787 1680
rect 783 1673 787 1674
rect 791 1678 795 1679
rect 791 1672 795 1674
rect 558 1671 564 1672
rect 486 1666 492 1667
rect 514 1667 520 1668
rect 514 1663 515 1667
rect 519 1663 520 1667
rect 558 1667 559 1671
rect 563 1667 564 1671
rect 558 1666 564 1667
rect 630 1671 636 1672
rect 630 1667 631 1671
rect 635 1667 636 1671
rect 630 1666 636 1667
rect 710 1671 716 1672
rect 710 1667 711 1671
rect 715 1667 716 1671
rect 710 1666 716 1667
rect 790 1671 796 1672
rect 790 1667 791 1671
rect 795 1667 796 1671
rect 790 1666 796 1667
rect 514 1662 520 1663
rect 522 1663 528 1664
rect 522 1659 523 1663
rect 527 1659 528 1663
rect 522 1658 528 1659
rect 678 1663 684 1664
rect 678 1659 679 1663
rect 683 1659 684 1663
rect 678 1658 684 1659
rect 414 1654 420 1655
rect 414 1650 415 1654
rect 419 1650 420 1654
rect 414 1649 420 1650
rect 486 1654 492 1655
rect 486 1650 487 1654
rect 491 1650 492 1654
rect 486 1649 492 1650
rect 350 1647 356 1648
rect 350 1643 351 1647
rect 355 1643 356 1647
rect 350 1642 356 1643
rect 416 1639 418 1649
rect 488 1639 490 1649
rect 524 1640 526 1658
rect 558 1654 564 1655
rect 558 1650 559 1654
rect 563 1650 564 1654
rect 558 1649 564 1650
rect 630 1654 636 1655
rect 630 1650 631 1654
rect 635 1650 636 1654
rect 630 1649 636 1650
rect 522 1639 528 1640
rect 560 1639 562 1649
rect 614 1647 620 1648
rect 614 1643 615 1647
rect 619 1643 620 1647
rect 614 1642 620 1643
rect 167 1638 171 1639
rect 167 1633 171 1634
rect 183 1638 187 1639
rect 183 1633 187 1634
rect 215 1638 219 1639
rect 215 1633 219 1634
rect 247 1638 251 1639
rect 247 1633 251 1634
rect 279 1638 283 1639
rect 279 1633 283 1634
rect 303 1638 307 1639
rect 303 1633 307 1634
rect 343 1638 347 1639
rect 343 1633 347 1634
rect 359 1638 363 1639
rect 359 1633 363 1634
rect 415 1638 419 1639
rect 415 1633 419 1634
rect 471 1638 475 1639
rect 471 1633 475 1634
rect 487 1638 491 1639
rect 522 1635 523 1639
rect 527 1635 528 1639
rect 522 1634 528 1635
rect 535 1638 539 1639
rect 487 1633 491 1634
rect 535 1633 539 1634
rect 559 1638 563 1639
rect 559 1633 563 1634
rect 599 1638 603 1639
rect 599 1633 603 1634
rect 150 1627 156 1628
rect 150 1623 151 1627
rect 155 1623 156 1627
rect 184 1623 186 1633
rect 198 1627 204 1628
rect 198 1623 199 1627
rect 203 1623 204 1627
rect 248 1623 250 1633
rect 304 1623 306 1633
rect 360 1623 362 1633
rect 416 1623 418 1633
rect 472 1623 474 1633
rect 498 1631 504 1632
rect 490 1627 496 1628
rect 490 1623 491 1627
rect 495 1623 496 1627
rect 498 1627 499 1631
rect 503 1627 504 1631
rect 498 1626 504 1627
rect 110 1619 116 1620
rect 134 1622 140 1623
rect 150 1622 156 1623
rect 182 1622 188 1623
rect 198 1622 204 1623
rect 246 1622 252 1623
rect 134 1618 135 1622
rect 139 1618 140 1622
rect 134 1617 140 1618
rect 182 1618 183 1622
rect 187 1618 188 1622
rect 182 1617 188 1618
rect 150 1611 156 1612
rect 110 1607 116 1608
rect 110 1603 111 1607
rect 115 1603 116 1607
rect 150 1607 151 1611
rect 155 1607 156 1611
rect 150 1606 156 1607
rect 110 1602 116 1603
rect 134 1605 140 1606
rect 112 1599 114 1602
rect 134 1601 135 1605
rect 139 1601 140 1605
rect 134 1600 140 1601
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 135 1598 139 1600
rect 112 1590 114 1593
rect 135 1592 139 1594
rect 134 1591 140 1592
rect 110 1589 116 1590
rect 110 1585 111 1589
rect 115 1585 116 1589
rect 134 1587 135 1591
rect 139 1587 140 1591
rect 134 1586 140 1587
rect 110 1584 116 1585
rect 134 1574 140 1575
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 134 1570 135 1574
rect 139 1570 140 1574
rect 134 1569 140 1570
rect 110 1567 116 1568
rect 112 1559 114 1567
rect 136 1559 138 1569
rect 152 1568 154 1606
rect 182 1605 188 1606
rect 182 1601 183 1605
rect 187 1601 188 1605
rect 182 1600 188 1601
rect 200 1600 202 1622
rect 246 1618 247 1622
rect 251 1618 252 1622
rect 246 1617 252 1618
rect 302 1622 308 1623
rect 302 1618 303 1622
rect 307 1618 308 1622
rect 302 1617 308 1618
rect 358 1622 364 1623
rect 358 1618 359 1622
rect 363 1618 364 1622
rect 358 1617 364 1618
rect 414 1622 420 1623
rect 414 1618 415 1622
rect 419 1618 420 1622
rect 414 1617 420 1618
rect 470 1622 476 1623
rect 490 1622 496 1623
rect 470 1618 471 1622
rect 475 1618 476 1622
rect 470 1617 476 1618
rect 446 1611 452 1612
rect 446 1607 447 1611
rect 451 1607 452 1611
rect 446 1606 452 1607
rect 246 1605 252 1606
rect 246 1601 247 1605
rect 251 1601 252 1605
rect 246 1600 252 1601
rect 302 1605 308 1606
rect 302 1601 303 1605
rect 307 1601 308 1605
rect 302 1600 308 1601
rect 358 1605 364 1606
rect 358 1601 359 1605
rect 363 1601 364 1605
rect 358 1600 364 1601
rect 414 1605 420 1606
rect 414 1601 415 1605
rect 419 1601 420 1605
rect 414 1600 420 1601
rect 167 1598 171 1599
rect 167 1592 171 1594
rect 183 1598 187 1600
rect 198 1599 204 1600
rect 198 1595 199 1599
rect 203 1595 204 1599
rect 198 1594 204 1595
rect 223 1598 227 1599
rect 183 1593 187 1594
rect 223 1592 227 1594
rect 247 1598 251 1600
rect 247 1593 251 1594
rect 279 1598 283 1599
rect 279 1592 283 1594
rect 303 1598 307 1600
rect 303 1593 307 1594
rect 335 1598 339 1599
rect 335 1592 339 1594
rect 359 1598 363 1600
rect 359 1593 363 1594
rect 383 1598 387 1599
rect 383 1592 387 1594
rect 415 1598 419 1600
rect 415 1593 419 1594
rect 431 1598 435 1599
rect 431 1592 435 1594
rect 166 1591 172 1592
rect 166 1587 167 1591
rect 171 1587 172 1591
rect 166 1586 172 1587
rect 222 1591 228 1592
rect 222 1587 223 1591
rect 227 1587 228 1591
rect 222 1586 228 1587
rect 278 1591 284 1592
rect 278 1587 279 1591
rect 283 1587 284 1591
rect 278 1586 284 1587
rect 334 1591 340 1592
rect 334 1587 335 1591
rect 339 1587 340 1591
rect 334 1586 340 1587
rect 382 1591 388 1592
rect 382 1587 383 1591
rect 387 1587 388 1591
rect 382 1586 388 1587
rect 430 1591 436 1592
rect 430 1587 431 1591
rect 435 1587 436 1591
rect 430 1586 436 1587
rect 182 1583 188 1584
rect 182 1579 183 1583
rect 187 1579 188 1583
rect 182 1578 188 1579
rect 374 1583 380 1584
rect 374 1579 375 1583
rect 379 1579 380 1583
rect 374 1578 380 1579
rect 166 1574 172 1575
rect 166 1570 167 1574
rect 171 1570 172 1574
rect 166 1569 172 1570
rect 150 1567 156 1568
rect 150 1563 151 1567
rect 155 1563 156 1567
rect 150 1562 156 1563
rect 168 1559 170 1569
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 135 1558 139 1559
rect 135 1553 139 1554
rect 167 1558 171 1559
rect 167 1553 171 1554
rect 112 1545 114 1553
rect 110 1544 116 1545
rect 110 1540 111 1544
rect 115 1540 116 1544
rect 136 1543 138 1553
rect 168 1543 170 1553
rect 184 1548 186 1578
rect 222 1574 228 1575
rect 222 1570 223 1574
rect 227 1570 228 1574
rect 222 1569 228 1570
rect 278 1574 284 1575
rect 278 1570 279 1574
rect 283 1570 284 1574
rect 278 1569 284 1570
rect 334 1574 340 1575
rect 334 1570 335 1574
rect 339 1570 340 1574
rect 334 1569 340 1570
rect 224 1559 226 1569
rect 234 1567 240 1568
rect 234 1563 235 1567
rect 239 1563 240 1567
rect 234 1562 240 1563
rect 215 1558 219 1559
rect 215 1553 219 1554
rect 223 1558 227 1559
rect 223 1553 227 1554
rect 182 1547 188 1548
rect 182 1543 183 1547
rect 187 1543 188 1547
rect 216 1543 218 1553
rect 110 1539 116 1540
rect 134 1542 140 1543
rect 134 1538 135 1542
rect 139 1538 140 1542
rect 134 1537 140 1538
rect 166 1542 172 1543
rect 182 1542 188 1543
rect 214 1542 220 1543
rect 166 1538 167 1542
rect 171 1538 172 1542
rect 166 1537 172 1538
rect 214 1538 215 1542
rect 219 1538 220 1542
rect 214 1537 220 1538
rect 236 1532 238 1562
rect 280 1559 282 1569
rect 336 1559 338 1569
rect 263 1558 267 1559
rect 263 1553 267 1554
rect 279 1558 283 1559
rect 279 1553 283 1554
rect 311 1558 315 1559
rect 311 1553 315 1554
rect 335 1558 339 1559
rect 335 1553 339 1554
rect 359 1558 363 1559
rect 359 1553 363 1554
rect 264 1543 266 1553
rect 312 1543 314 1553
rect 350 1547 356 1548
rect 350 1543 351 1547
rect 355 1543 356 1547
rect 360 1543 362 1553
rect 376 1548 378 1578
rect 382 1574 388 1575
rect 382 1570 383 1574
rect 387 1570 388 1574
rect 382 1569 388 1570
rect 430 1574 436 1575
rect 430 1570 431 1574
rect 435 1570 436 1574
rect 430 1569 436 1570
rect 384 1559 386 1569
rect 432 1559 434 1569
rect 448 1568 450 1606
rect 470 1605 476 1606
rect 470 1601 471 1605
rect 475 1601 476 1605
rect 470 1600 476 1601
rect 471 1598 475 1600
rect 471 1593 475 1594
rect 479 1598 483 1599
rect 479 1592 483 1594
rect 478 1591 484 1592
rect 478 1587 479 1591
rect 483 1587 484 1591
rect 478 1586 484 1587
rect 492 1584 494 1622
rect 500 1612 502 1626
rect 536 1623 538 1633
rect 600 1623 602 1633
rect 534 1622 540 1623
rect 534 1618 535 1622
rect 539 1618 540 1622
rect 534 1617 540 1618
rect 598 1622 604 1623
rect 598 1618 599 1622
rect 603 1618 604 1622
rect 598 1617 604 1618
rect 616 1612 618 1642
rect 632 1639 634 1649
rect 631 1638 635 1639
rect 631 1633 635 1634
rect 663 1638 667 1639
rect 663 1633 667 1634
rect 664 1623 666 1633
rect 680 1628 682 1658
rect 710 1654 716 1655
rect 710 1650 711 1654
rect 715 1650 716 1654
rect 710 1649 716 1650
rect 790 1654 796 1655
rect 790 1650 791 1654
rect 795 1650 796 1654
rect 790 1649 796 1650
rect 712 1639 714 1649
rect 792 1639 794 1649
rect 804 1648 806 1686
rect 838 1685 844 1686
rect 838 1681 839 1685
rect 843 1681 844 1685
rect 838 1680 844 1681
rect 839 1678 843 1680
rect 839 1673 843 1674
rect 871 1678 875 1679
rect 871 1672 875 1674
rect 870 1671 876 1672
rect 870 1667 871 1671
rect 875 1667 876 1671
rect 870 1666 876 1667
rect 888 1664 890 1702
rect 894 1698 895 1702
rect 899 1698 900 1702
rect 894 1697 900 1698
rect 950 1702 956 1703
rect 950 1698 951 1702
rect 955 1698 956 1702
rect 950 1697 956 1698
rect 1006 1702 1012 1703
rect 1006 1698 1007 1702
rect 1011 1698 1012 1702
rect 1006 1697 1012 1698
rect 1062 1702 1068 1703
rect 1062 1698 1063 1702
rect 1067 1698 1068 1702
rect 1062 1697 1068 1698
rect 1108 1692 1110 1706
rect 1120 1703 1122 1713
rect 1138 1711 1139 1715
rect 1143 1711 1144 1715
rect 1175 1713 1179 1714
rect 1231 1718 1235 1719
rect 1231 1713 1235 1714
rect 1287 1718 1291 1719
rect 1287 1713 1291 1714
rect 1335 1718 1339 1719
rect 1335 1713 1339 1714
rect 1375 1718 1379 1719
rect 1375 1713 1379 1714
rect 1423 1718 1427 1719
rect 1423 1713 1427 1714
rect 1471 1718 1475 1719
rect 1471 1713 1475 1714
rect 1519 1718 1523 1719
rect 1519 1713 1523 1714
rect 1663 1718 1667 1719
rect 1663 1713 1667 1714
rect 1138 1710 1144 1711
rect 1118 1702 1124 1703
rect 1118 1698 1119 1702
rect 1123 1698 1124 1702
rect 1118 1697 1124 1698
rect 1140 1692 1142 1710
rect 1176 1703 1178 1713
rect 1232 1703 1234 1713
rect 1270 1711 1276 1712
rect 1262 1707 1268 1708
rect 1262 1703 1263 1707
rect 1267 1703 1268 1707
rect 1270 1707 1271 1711
rect 1275 1707 1276 1711
rect 1270 1706 1276 1707
rect 1174 1702 1180 1703
rect 1174 1698 1175 1702
rect 1179 1698 1180 1702
rect 1174 1697 1180 1698
rect 1230 1702 1236 1703
rect 1262 1702 1268 1703
rect 1230 1698 1231 1702
rect 1235 1698 1236 1702
rect 1230 1697 1236 1698
rect 1106 1691 1112 1692
rect 1106 1687 1107 1691
rect 1111 1687 1112 1691
rect 1106 1686 1112 1687
rect 1138 1691 1144 1692
rect 1138 1687 1139 1691
rect 1143 1687 1144 1691
rect 1138 1686 1144 1687
rect 1190 1691 1196 1692
rect 1190 1687 1191 1691
rect 1195 1687 1196 1691
rect 1190 1686 1196 1687
rect 894 1685 900 1686
rect 894 1681 895 1685
rect 899 1681 900 1685
rect 894 1680 900 1681
rect 950 1685 956 1686
rect 950 1681 951 1685
rect 955 1681 956 1685
rect 950 1680 956 1681
rect 1006 1685 1012 1686
rect 1006 1681 1007 1685
rect 1011 1681 1012 1685
rect 1006 1680 1012 1681
rect 1062 1685 1068 1686
rect 1062 1681 1063 1685
rect 1067 1681 1068 1685
rect 1062 1680 1068 1681
rect 1118 1685 1124 1686
rect 1118 1681 1119 1685
rect 1123 1681 1124 1685
rect 1118 1680 1124 1681
rect 1174 1685 1180 1686
rect 1174 1681 1175 1685
rect 1179 1681 1180 1685
rect 1174 1680 1180 1681
rect 895 1678 899 1680
rect 895 1673 899 1674
rect 951 1678 955 1680
rect 951 1672 955 1674
rect 1007 1678 1011 1680
rect 1007 1673 1011 1674
rect 1031 1678 1035 1679
rect 1031 1672 1035 1674
rect 1063 1678 1067 1680
rect 1063 1673 1067 1674
rect 1103 1678 1107 1679
rect 1103 1672 1107 1674
rect 1119 1678 1123 1680
rect 1119 1673 1123 1674
rect 1175 1678 1179 1680
rect 1175 1672 1179 1674
rect 950 1671 956 1672
rect 950 1667 951 1671
rect 955 1667 956 1671
rect 950 1666 956 1667
rect 1030 1671 1036 1672
rect 1030 1667 1031 1671
rect 1035 1667 1036 1671
rect 1030 1666 1036 1667
rect 1102 1671 1108 1672
rect 1102 1667 1103 1671
rect 1107 1667 1108 1671
rect 1102 1666 1108 1667
rect 1174 1671 1180 1672
rect 1174 1667 1175 1671
rect 1179 1667 1180 1671
rect 1174 1666 1180 1667
rect 886 1663 892 1664
rect 886 1659 887 1663
rect 891 1659 892 1663
rect 886 1658 892 1659
rect 1146 1663 1152 1664
rect 1146 1659 1147 1663
rect 1151 1659 1152 1663
rect 1146 1658 1152 1659
rect 870 1654 876 1655
rect 870 1650 871 1654
rect 875 1650 876 1654
rect 870 1649 876 1650
rect 950 1654 956 1655
rect 950 1650 951 1654
rect 955 1650 956 1654
rect 950 1649 956 1650
rect 1030 1654 1036 1655
rect 1030 1650 1031 1654
rect 1035 1650 1036 1654
rect 1030 1649 1036 1650
rect 1102 1654 1108 1655
rect 1102 1650 1103 1654
rect 1107 1650 1108 1654
rect 1102 1649 1108 1650
rect 802 1647 808 1648
rect 802 1643 803 1647
rect 807 1643 808 1647
rect 802 1642 808 1643
rect 872 1639 874 1649
rect 952 1639 954 1649
rect 962 1647 968 1648
rect 962 1643 963 1647
rect 967 1643 968 1647
rect 962 1642 968 1643
rect 711 1638 715 1639
rect 711 1633 715 1634
rect 727 1638 731 1639
rect 727 1633 731 1634
rect 791 1638 795 1639
rect 791 1633 795 1634
rect 799 1638 803 1639
rect 799 1633 803 1634
rect 871 1638 875 1639
rect 871 1633 875 1634
rect 943 1638 947 1639
rect 943 1633 947 1634
rect 951 1638 955 1639
rect 951 1633 955 1634
rect 678 1627 684 1628
rect 678 1623 679 1627
rect 683 1623 684 1627
rect 728 1623 730 1633
rect 800 1623 802 1633
rect 814 1627 820 1628
rect 814 1623 815 1627
rect 819 1623 820 1627
rect 872 1623 874 1633
rect 944 1623 946 1633
rect 662 1622 668 1623
rect 678 1622 684 1623
rect 726 1622 732 1623
rect 662 1618 663 1622
rect 667 1618 668 1622
rect 662 1617 668 1618
rect 726 1618 727 1622
rect 731 1618 732 1622
rect 726 1617 732 1618
rect 798 1622 804 1623
rect 814 1622 820 1623
rect 870 1622 876 1623
rect 798 1618 799 1622
rect 803 1618 804 1622
rect 798 1617 804 1618
rect 498 1611 504 1612
rect 498 1607 499 1611
rect 503 1607 504 1611
rect 498 1606 504 1607
rect 614 1611 620 1612
rect 614 1607 615 1611
rect 619 1607 620 1611
rect 614 1606 620 1607
rect 742 1611 748 1612
rect 742 1607 743 1611
rect 747 1607 748 1611
rect 742 1606 748 1607
rect 534 1605 540 1606
rect 534 1601 535 1605
rect 539 1601 540 1605
rect 534 1600 540 1601
rect 598 1605 604 1606
rect 598 1601 599 1605
rect 603 1601 604 1605
rect 598 1600 604 1601
rect 662 1605 668 1606
rect 662 1601 663 1605
rect 667 1601 668 1605
rect 662 1600 668 1601
rect 726 1605 732 1606
rect 726 1601 727 1605
rect 731 1601 732 1605
rect 726 1600 732 1601
rect 535 1598 539 1600
rect 535 1592 539 1594
rect 599 1598 603 1600
rect 599 1592 603 1594
rect 663 1598 667 1600
rect 663 1592 667 1594
rect 727 1598 731 1600
rect 727 1592 731 1594
rect 534 1591 540 1592
rect 534 1587 535 1591
rect 539 1587 540 1591
rect 534 1586 540 1587
rect 598 1591 604 1592
rect 598 1587 599 1591
rect 603 1587 604 1591
rect 598 1586 604 1587
rect 662 1591 668 1592
rect 662 1587 663 1591
rect 667 1587 668 1591
rect 662 1586 668 1587
rect 726 1591 732 1592
rect 726 1587 727 1591
rect 731 1587 732 1591
rect 726 1586 732 1587
rect 490 1583 496 1584
rect 490 1579 491 1583
rect 495 1579 496 1583
rect 490 1578 496 1579
rect 478 1574 484 1575
rect 478 1570 479 1574
rect 483 1570 484 1574
rect 478 1569 484 1570
rect 534 1574 540 1575
rect 534 1570 535 1574
rect 539 1570 540 1574
rect 534 1569 540 1570
rect 598 1574 604 1575
rect 598 1570 599 1574
rect 603 1570 604 1574
rect 598 1569 604 1570
rect 662 1574 668 1575
rect 662 1570 663 1574
rect 667 1570 668 1574
rect 662 1569 668 1570
rect 726 1574 732 1575
rect 726 1570 727 1574
rect 731 1570 732 1574
rect 726 1569 732 1570
rect 446 1567 452 1568
rect 446 1563 447 1567
rect 451 1563 452 1567
rect 446 1562 452 1563
rect 480 1559 482 1569
rect 536 1559 538 1569
rect 586 1567 592 1568
rect 586 1563 587 1567
rect 591 1563 592 1567
rect 586 1562 592 1563
rect 383 1558 387 1559
rect 383 1553 387 1554
rect 407 1558 411 1559
rect 407 1553 411 1554
rect 431 1558 435 1559
rect 431 1553 435 1554
rect 455 1558 459 1559
rect 455 1553 459 1554
rect 479 1558 483 1559
rect 479 1553 483 1554
rect 511 1558 515 1559
rect 511 1553 515 1554
rect 535 1558 539 1559
rect 535 1553 539 1554
rect 567 1558 571 1559
rect 567 1553 571 1554
rect 374 1547 380 1548
rect 374 1543 375 1547
rect 379 1543 380 1547
rect 408 1543 410 1553
rect 456 1543 458 1553
rect 512 1543 514 1553
rect 568 1543 570 1553
rect 262 1542 268 1543
rect 262 1538 263 1542
rect 267 1538 268 1542
rect 262 1537 268 1538
rect 310 1542 316 1543
rect 350 1542 356 1543
rect 358 1542 364 1543
rect 374 1542 380 1543
rect 406 1542 412 1543
rect 310 1538 311 1542
rect 315 1538 316 1542
rect 310 1537 316 1538
rect 150 1531 156 1532
rect 110 1527 116 1528
rect 110 1523 111 1527
rect 115 1523 116 1527
rect 150 1527 151 1531
rect 155 1527 156 1531
rect 150 1526 156 1527
rect 234 1531 240 1532
rect 234 1527 235 1531
rect 239 1527 240 1531
rect 234 1526 240 1527
rect 110 1522 116 1523
rect 134 1525 140 1526
rect 112 1515 114 1522
rect 134 1521 135 1525
rect 139 1521 140 1525
rect 134 1520 140 1521
rect 136 1515 138 1520
rect 111 1514 115 1515
rect 111 1509 115 1510
rect 135 1514 139 1515
rect 112 1506 114 1509
rect 135 1508 139 1510
rect 134 1507 140 1508
rect 110 1505 116 1506
rect 110 1501 111 1505
rect 115 1501 116 1505
rect 134 1503 135 1507
rect 139 1503 140 1507
rect 134 1502 140 1503
rect 110 1500 116 1501
rect 134 1490 140 1491
rect 110 1488 116 1489
rect 110 1484 111 1488
rect 115 1484 116 1488
rect 134 1486 135 1490
rect 139 1486 140 1490
rect 134 1485 140 1486
rect 110 1483 116 1484
rect 112 1475 114 1483
rect 136 1475 138 1485
rect 152 1484 154 1526
rect 166 1525 172 1526
rect 166 1521 167 1525
rect 171 1521 172 1525
rect 166 1520 172 1521
rect 214 1525 220 1526
rect 214 1521 215 1525
rect 219 1521 220 1525
rect 214 1520 220 1521
rect 262 1525 268 1526
rect 262 1521 263 1525
rect 267 1521 268 1525
rect 262 1520 268 1521
rect 310 1525 316 1526
rect 310 1521 311 1525
rect 315 1521 316 1525
rect 310 1520 316 1521
rect 168 1515 170 1520
rect 216 1515 218 1520
rect 264 1515 266 1520
rect 312 1515 314 1520
rect 352 1516 354 1542
rect 358 1538 359 1542
rect 363 1538 364 1542
rect 358 1537 364 1538
rect 406 1538 407 1542
rect 411 1538 412 1542
rect 406 1537 412 1538
rect 454 1542 460 1543
rect 454 1538 455 1542
rect 459 1538 460 1542
rect 454 1537 460 1538
rect 510 1542 516 1543
rect 510 1538 511 1542
rect 515 1538 516 1542
rect 510 1537 516 1538
rect 566 1542 572 1543
rect 566 1538 567 1542
rect 571 1538 572 1542
rect 566 1537 572 1538
rect 588 1532 590 1562
rect 600 1559 602 1569
rect 664 1559 666 1569
rect 728 1559 730 1569
rect 744 1568 746 1606
rect 798 1605 804 1606
rect 798 1601 799 1605
rect 803 1601 804 1605
rect 798 1600 804 1601
rect 799 1598 803 1600
rect 799 1592 803 1594
rect 798 1591 804 1592
rect 798 1587 799 1591
rect 803 1587 804 1591
rect 798 1586 804 1587
rect 816 1584 818 1622
rect 870 1618 871 1622
rect 875 1618 876 1622
rect 870 1617 876 1618
rect 942 1622 948 1623
rect 942 1618 943 1622
rect 947 1618 948 1622
rect 942 1617 948 1618
rect 964 1612 966 1642
rect 1032 1639 1034 1649
rect 1104 1639 1106 1649
rect 1148 1640 1150 1658
rect 1166 1655 1172 1656
rect 1166 1651 1167 1655
rect 1171 1651 1172 1655
rect 1166 1650 1172 1651
rect 1174 1654 1180 1655
rect 1174 1650 1175 1654
rect 1179 1650 1180 1654
rect 1146 1639 1152 1640
rect 1023 1638 1027 1639
rect 1023 1633 1027 1634
rect 1031 1638 1035 1639
rect 1031 1633 1035 1634
rect 1103 1638 1107 1639
rect 1146 1635 1147 1639
rect 1151 1635 1152 1639
rect 1146 1634 1152 1635
rect 1103 1633 1107 1634
rect 1024 1623 1026 1633
rect 1104 1623 1106 1633
rect 1168 1632 1170 1650
rect 1174 1649 1180 1650
rect 1176 1639 1178 1649
rect 1192 1648 1194 1686
rect 1230 1685 1236 1686
rect 1230 1681 1231 1685
rect 1235 1681 1236 1685
rect 1230 1680 1236 1681
rect 1231 1678 1235 1680
rect 1231 1673 1235 1674
rect 1247 1678 1251 1679
rect 1247 1672 1251 1674
rect 1246 1671 1252 1672
rect 1246 1667 1247 1671
rect 1251 1667 1252 1671
rect 1246 1666 1252 1667
rect 1264 1664 1266 1702
rect 1272 1692 1274 1706
rect 1288 1703 1290 1713
rect 1336 1703 1338 1713
rect 1376 1703 1378 1713
rect 1424 1703 1426 1713
rect 1458 1711 1464 1712
rect 1458 1707 1459 1711
rect 1463 1707 1464 1711
rect 1458 1706 1464 1707
rect 1286 1702 1292 1703
rect 1286 1698 1287 1702
rect 1291 1698 1292 1702
rect 1286 1697 1292 1698
rect 1334 1702 1340 1703
rect 1334 1698 1335 1702
rect 1339 1698 1340 1702
rect 1334 1697 1340 1698
rect 1374 1702 1380 1703
rect 1374 1698 1375 1702
rect 1379 1698 1380 1702
rect 1374 1697 1380 1698
rect 1422 1702 1428 1703
rect 1422 1698 1423 1702
rect 1427 1698 1428 1702
rect 1422 1697 1428 1698
rect 1460 1692 1462 1706
rect 1472 1703 1474 1713
rect 1520 1703 1522 1713
rect 1664 1705 1666 1713
rect 1662 1704 1668 1705
rect 1470 1702 1476 1703
rect 1470 1698 1471 1702
rect 1475 1698 1476 1702
rect 1470 1697 1476 1698
rect 1518 1702 1524 1703
rect 1518 1698 1519 1702
rect 1523 1698 1524 1702
rect 1662 1700 1663 1704
rect 1667 1700 1668 1704
rect 1662 1699 1668 1700
rect 1518 1697 1524 1698
rect 1270 1691 1276 1692
rect 1270 1687 1271 1691
rect 1275 1687 1276 1691
rect 1270 1686 1276 1687
rect 1458 1691 1464 1692
rect 1458 1687 1459 1691
rect 1463 1687 1464 1691
rect 1458 1686 1464 1687
rect 1662 1687 1668 1688
rect 1286 1685 1292 1686
rect 1286 1681 1287 1685
rect 1291 1681 1292 1685
rect 1286 1680 1292 1681
rect 1334 1685 1340 1686
rect 1334 1681 1335 1685
rect 1339 1681 1340 1685
rect 1334 1680 1340 1681
rect 1374 1685 1380 1686
rect 1374 1681 1375 1685
rect 1379 1681 1380 1685
rect 1374 1680 1380 1681
rect 1422 1685 1428 1686
rect 1422 1681 1423 1685
rect 1427 1681 1428 1685
rect 1422 1680 1428 1681
rect 1470 1685 1476 1686
rect 1470 1681 1471 1685
rect 1475 1681 1476 1685
rect 1470 1680 1476 1681
rect 1518 1685 1524 1686
rect 1518 1681 1519 1685
rect 1523 1681 1524 1685
rect 1662 1683 1663 1687
rect 1667 1683 1668 1687
rect 1662 1682 1668 1683
rect 1518 1680 1524 1681
rect 1287 1678 1291 1680
rect 1287 1673 1291 1674
rect 1319 1678 1323 1679
rect 1319 1672 1323 1674
rect 1335 1678 1339 1680
rect 1335 1673 1339 1674
rect 1375 1678 1379 1680
rect 1410 1679 1416 1680
rect 1375 1673 1379 1674
rect 1391 1678 1395 1679
rect 1410 1675 1411 1679
rect 1415 1675 1416 1679
rect 1410 1674 1416 1675
rect 1423 1678 1427 1680
rect 1391 1672 1395 1674
rect 1318 1671 1324 1672
rect 1318 1667 1319 1671
rect 1323 1667 1324 1671
rect 1318 1666 1324 1667
rect 1390 1671 1396 1672
rect 1390 1667 1391 1671
rect 1395 1667 1396 1671
rect 1390 1666 1396 1667
rect 1262 1663 1268 1664
rect 1262 1659 1263 1663
rect 1267 1659 1268 1663
rect 1262 1658 1268 1659
rect 1246 1654 1252 1655
rect 1246 1650 1247 1654
rect 1251 1650 1252 1654
rect 1246 1649 1252 1650
rect 1318 1654 1324 1655
rect 1318 1650 1319 1654
rect 1323 1650 1324 1654
rect 1318 1649 1324 1650
rect 1390 1654 1396 1655
rect 1390 1650 1391 1654
rect 1395 1650 1396 1654
rect 1390 1649 1396 1650
rect 1190 1647 1196 1648
rect 1190 1643 1191 1647
rect 1195 1643 1196 1647
rect 1190 1642 1196 1643
rect 1248 1639 1250 1649
rect 1320 1639 1322 1649
rect 1334 1647 1340 1648
rect 1334 1643 1335 1647
rect 1339 1643 1340 1647
rect 1334 1642 1340 1643
rect 1175 1638 1179 1639
rect 1175 1633 1179 1634
rect 1247 1638 1251 1639
rect 1247 1633 1251 1634
rect 1319 1638 1323 1639
rect 1319 1633 1323 1634
rect 1166 1631 1172 1632
rect 1166 1627 1167 1631
rect 1171 1627 1172 1631
rect 1166 1626 1172 1627
rect 1176 1623 1178 1633
rect 1248 1623 1250 1633
rect 1302 1631 1308 1632
rect 1294 1627 1300 1628
rect 1294 1623 1295 1627
rect 1299 1623 1300 1627
rect 1302 1627 1303 1631
rect 1307 1627 1308 1631
rect 1302 1626 1308 1627
rect 1022 1622 1028 1623
rect 1022 1618 1023 1622
rect 1027 1618 1028 1622
rect 1022 1617 1028 1618
rect 1102 1622 1108 1623
rect 1102 1618 1103 1622
rect 1107 1618 1108 1622
rect 1102 1617 1108 1618
rect 1174 1622 1180 1623
rect 1174 1618 1175 1622
rect 1179 1618 1180 1622
rect 1174 1617 1180 1618
rect 1246 1622 1252 1623
rect 1294 1622 1300 1623
rect 1246 1618 1247 1622
rect 1251 1618 1252 1622
rect 1246 1617 1252 1618
rect 962 1611 968 1612
rect 962 1607 963 1611
rect 967 1607 968 1611
rect 962 1606 968 1607
rect 1034 1611 1040 1612
rect 1034 1607 1035 1611
rect 1039 1607 1040 1611
rect 1034 1606 1040 1607
rect 870 1605 876 1606
rect 870 1601 871 1605
rect 875 1601 876 1605
rect 870 1600 876 1601
rect 942 1605 948 1606
rect 942 1601 943 1605
rect 947 1601 948 1605
rect 942 1600 948 1601
rect 1022 1605 1028 1606
rect 1022 1601 1023 1605
rect 1027 1601 1028 1605
rect 1036 1603 1038 1606
rect 1022 1600 1028 1601
rect 1032 1601 1038 1603
rect 1102 1605 1108 1606
rect 1102 1601 1103 1605
rect 1107 1601 1108 1605
rect 871 1598 875 1600
rect 871 1592 875 1594
rect 943 1598 947 1600
rect 943 1593 947 1594
rect 951 1598 955 1599
rect 951 1592 955 1594
rect 1023 1598 1027 1600
rect 1023 1593 1027 1594
rect 870 1591 876 1592
rect 870 1587 871 1591
rect 875 1587 876 1591
rect 870 1586 876 1587
rect 950 1591 956 1592
rect 950 1587 951 1591
rect 955 1587 956 1591
rect 950 1586 956 1587
rect 814 1583 820 1584
rect 814 1579 815 1583
rect 819 1579 820 1583
rect 814 1578 820 1579
rect 798 1574 804 1575
rect 798 1570 799 1574
rect 803 1570 804 1574
rect 798 1569 804 1570
rect 870 1574 876 1575
rect 870 1570 871 1574
rect 875 1570 876 1574
rect 870 1569 876 1570
rect 950 1574 956 1575
rect 950 1570 951 1574
rect 955 1570 956 1574
rect 950 1569 956 1570
rect 742 1567 748 1568
rect 742 1563 743 1567
rect 747 1563 748 1567
rect 742 1562 748 1563
rect 800 1559 802 1569
rect 850 1567 856 1568
rect 850 1563 851 1567
rect 855 1563 856 1567
rect 850 1562 856 1563
rect 599 1558 603 1559
rect 599 1553 603 1554
rect 631 1558 635 1559
rect 631 1553 635 1554
rect 663 1558 667 1559
rect 663 1553 667 1554
rect 695 1558 699 1559
rect 695 1553 699 1554
rect 727 1558 731 1559
rect 727 1553 731 1554
rect 759 1558 763 1559
rect 759 1553 763 1554
rect 799 1558 803 1559
rect 799 1553 803 1554
rect 831 1558 835 1559
rect 831 1553 835 1554
rect 632 1543 634 1553
rect 696 1543 698 1553
rect 760 1543 762 1553
rect 832 1543 834 1553
rect 630 1542 636 1543
rect 630 1538 631 1542
rect 635 1538 636 1542
rect 630 1537 636 1538
rect 694 1542 700 1543
rect 694 1538 695 1542
rect 699 1538 700 1542
rect 694 1537 700 1538
rect 758 1542 764 1543
rect 758 1538 759 1542
rect 763 1538 764 1542
rect 758 1537 764 1538
rect 830 1542 836 1543
rect 830 1538 831 1542
rect 835 1538 836 1542
rect 830 1537 836 1538
rect 852 1532 854 1562
rect 872 1559 874 1569
rect 952 1559 954 1569
rect 1032 1568 1034 1601
rect 1102 1600 1108 1601
rect 1174 1605 1180 1606
rect 1174 1601 1175 1605
rect 1179 1601 1180 1605
rect 1174 1600 1180 1601
rect 1246 1605 1252 1606
rect 1246 1601 1247 1605
rect 1251 1601 1252 1605
rect 1246 1600 1252 1601
rect 1039 1598 1043 1599
rect 1039 1592 1043 1594
rect 1103 1598 1107 1600
rect 1103 1593 1107 1594
rect 1119 1598 1123 1599
rect 1119 1592 1123 1594
rect 1175 1598 1179 1600
rect 1175 1593 1179 1594
rect 1199 1598 1203 1599
rect 1199 1592 1203 1594
rect 1247 1598 1251 1600
rect 1247 1593 1251 1594
rect 1279 1598 1283 1599
rect 1279 1592 1283 1594
rect 1038 1591 1044 1592
rect 1038 1587 1039 1591
rect 1043 1587 1044 1591
rect 1038 1586 1044 1587
rect 1118 1591 1124 1592
rect 1118 1587 1119 1591
rect 1123 1587 1124 1591
rect 1118 1586 1124 1587
rect 1198 1591 1204 1592
rect 1198 1587 1199 1591
rect 1203 1587 1204 1591
rect 1198 1586 1204 1587
rect 1278 1591 1284 1592
rect 1278 1587 1279 1591
rect 1283 1587 1284 1591
rect 1278 1586 1284 1587
rect 1296 1584 1298 1622
rect 1304 1612 1306 1626
rect 1320 1623 1322 1633
rect 1318 1622 1324 1623
rect 1318 1618 1319 1622
rect 1323 1618 1324 1622
rect 1318 1617 1324 1618
rect 1336 1612 1338 1642
rect 1392 1639 1394 1649
rect 1412 1648 1414 1674
rect 1423 1673 1427 1674
rect 1455 1678 1459 1679
rect 1455 1672 1459 1674
rect 1471 1678 1475 1680
rect 1471 1673 1475 1674
rect 1519 1678 1523 1680
rect 1664 1679 1666 1682
rect 1519 1672 1523 1674
rect 1583 1678 1587 1679
rect 1583 1672 1587 1674
rect 1623 1678 1627 1679
rect 1623 1672 1627 1674
rect 1663 1678 1667 1679
rect 1663 1673 1667 1674
rect 1454 1671 1460 1672
rect 1454 1667 1455 1671
rect 1459 1667 1460 1671
rect 1454 1666 1460 1667
rect 1518 1671 1524 1672
rect 1518 1667 1519 1671
rect 1523 1667 1524 1671
rect 1518 1666 1524 1667
rect 1582 1671 1588 1672
rect 1582 1667 1583 1671
rect 1587 1667 1588 1671
rect 1582 1666 1588 1667
rect 1622 1671 1628 1672
rect 1622 1667 1623 1671
rect 1627 1667 1628 1671
rect 1664 1670 1666 1673
rect 1622 1666 1628 1667
rect 1662 1669 1668 1670
rect 1662 1665 1663 1669
rect 1667 1665 1668 1669
rect 1662 1664 1668 1665
rect 1574 1663 1580 1664
rect 1574 1659 1575 1663
rect 1579 1659 1580 1663
rect 1574 1658 1580 1659
rect 1638 1663 1644 1664
rect 1638 1659 1639 1663
rect 1643 1659 1644 1663
rect 1638 1658 1644 1659
rect 1454 1654 1460 1655
rect 1454 1650 1455 1654
rect 1459 1650 1460 1654
rect 1454 1649 1460 1650
rect 1518 1654 1524 1655
rect 1518 1650 1519 1654
rect 1523 1650 1524 1654
rect 1518 1649 1524 1650
rect 1410 1647 1416 1648
rect 1410 1643 1411 1647
rect 1415 1643 1416 1647
rect 1410 1642 1416 1643
rect 1456 1639 1458 1649
rect 1520 1639 1522 1649
rect 1546 1647 1552 1648
rect 1546 1643 1547 1647
rect 1551 1643 1552 1647
rect 1546 1642 1552 1643
rect 1391 1638 1395 1639
rect 1391 1633 1395 1634
rect 1399 1638 1403 1639
rect 1399 1633 1403 1634
rect 1455 1638 1459 1639
rect 1455 1633 1459 1634
rect 1479 1638 1483 1639
rect 1479 1633 1483 1634
rect 1519 1638 1523 1639
rect 1519 1633 1523 1634
rect 1400 1623 1402 1633
rect 1480 1623 1482 1633
rect 1398 1622 1404 1623
rect 1398 1618 1399 1622
rect 1403 1618 1404 1622
rect 1398 1617 1404 1618
rect 1478 1622 1484 1623
rect 1478 1618 1479 1622
rect 1483 1618 1484 1622
rect 1478 1617 1484 1618
rect 1302 1611 1308 1612
rect 1302 1607 1303 1611
rect 1307 1607 1308 1611
rect 1302 1606 1308 1607
rect 1334 1611 1340 1612
rect 1334 1607 1335 1611
rect 1339 1607 1340 1611
rect 1334 1606 1340 1607
rect 1430 1611 1436 1612
rect 1430 1607 1431 1611
rect 1435 1607 1436 1611
rect 1430 1606 1436 1607
rect 1318 1605 1324 1606
rect 1318 1601 1319 1605
rect 1323 1601 1324 1605
rect 1318 1600 1324 1601
rect 1398 1605 1404 1606
rect 1398 1601 1399 1605
rect 1403 1601 1404 1605
rect 1398 1600 1404 1601
rect 1319 1598 1323 1600
rect 1319 1593 1323 1594
rect 1351 1598 1355 1599
rect 1351 1592 1355 1594
rect 1399 1598 1403 1600
rect 1399 1593 1403 1594
rect 1415 1598 1419 1599
rect 1415 1592 1419 1594
rect 1350 1591 1356 1592
rect 1350 1587 1351 1591
rect 1355 1587 1356 1591
rect 1350 1586 1356 1587
rect 1414 1591 1420 1592
rect 1414 1587 1415 1591
rect 1419 1587 1420 1591
rect 1414 1586 1420 1587
rect 1210 1583 1216 1584
rect 1210 1579 1211 1583
rect 1215 1579 1216 1583
rect 1210 1578 1216 1579
rect 1294 1583 1300 1584
rect 1294 1579 1295 1583
rect 1299 1579 1300 1583
rect 1294 1578 1300 1579
rect 1362 1583 1368 1584
rect 1362 1579 1363 1583
rect 1367 1579 1368 1583
rect 1362 1578 1368 1579
rect 1038 1574 1044 1575
rect 1038 1570 1039 1574
rect 1043 1570 1044 1574
rect 1038 1569 1044 1570
rect 1118 1574 1124 1575
rect 1118 1570 1119 1574
rect 1123 1570 1124 1574
rect 1118 1569 1124 1570
rect 1198 1574 1204 1575
rect 1198 1570 1199 1574
rect 1203 1570 1204 1574
rect 1198 1569 1204 1570
rect 1030 1567 1036 1568
rect 1030 1563 1031 1567
rect 1035 1563 1036 1567
rect 1030 1562 1036 1563
rect 1040 1559 1042 1569
rect 1120 1559 1122 1569
rect 1200 1559 1202 1569
rect 871 1558 875 1559
rect 871 1553 875 1554
rect 919 1558 923 1559
rect 919 1553 923 1554
rect 951 1558 955 1559
rect 951 1553 955 1554
rect 1007 1558 1011 1559
rect 1007 1553 1011 1554
rect 1039 1558 1043 1559
rect 1039 1553 1043 1554
rect 1095 1558 1099 1559
rect 1095 1553 1099 1554
rect 1119 1558 1123 1559
rect 1119 1553 1123 1554
rect 1183 1558 1187 1559
rect 1183 1553 1187 1554
rect 1199 1558 1203 1559
rect 1199 1553 1203 1554
rect 894 1547 900 1548
rect 894 1543 895 1547
rect 899 1543 900 1547
rect 920 1543 922 1553
rect 1008 1543 1010 1553
rect 1096 1543 1098 1553
rect 1184 1543 1186 1553
rect 1212 1548 1214 1578
rect 1278 1574 1284 1575
rect 1278 1570 1279 1574
rect 1283 1570 1284 1574
rect 1278 1569 1284 1570
rect 1350 1574 1356 1575
rect 1350 1570 1351 1574
rect 1355 1570 1356 1574
rect 1350 1569 1356 1570
rect 1280 1559 1282 1569
rect 1286 1567 1292 1568
rect 1286 1563 1287 1567
rect 1291 1563 1292 1567
rect 1286 1562 1292 1563
rect 1263 1558 1267 1559
rect 1263 1553 1267 1554
rect 1279 1558 1283 1559
rect 1279 1553 1283 1554
rect 1210 1547 1216 1548
rect 1210 1543 1211 1547
rect 1215 1543 1216 1547
rect 1264 1543 1266 1553
rect 894 1542 900 1543
rect 918 1542 924 1543
rect 586 1531 592 1532
rect 586 1527 587 1531
rect 591 1527 592 1531
rect 586 1526 592 1527
rect 770 1531 776 1532
rect 770 1527 771 1531
rect 775 1527 776 1531
rect 770 1526 776 1527
rect 850 1531 856 1532
rect 850 1527 851 1531
rect 855 1527 856 1531
rect 850 1526 856 1527
rect 358 1525 364 1526
rect 358 1521 359 1525
rect 363 1521 364 1525
rect 358 1520 364 1521
rect 406 1525 412 1526
rect 406 1521 407 1525
rect 411 1521 412 1525
rect 406 1520 412 1521
rect 454 1525 460 1526
rect 454 1521 455 1525
rect 459 1521 460 1525
rect 454 1520 460 1521
rect 510 1525 516 1526
rect 510 1521 511 1525
rect 515 1521 516 1525
rect 510 1520 516 1521
rect 566 1525 572 1526
rect 566 1521 567 1525
rect 571 1521 572 1525
rect 566 1520 572 1521
rect 630 1525 636 1526
rect 630 1521 631 1525
rect 635 1521 636 1525
rect 630 1520 636 1521
rect 694 1525 700 1526
rect 694 1521 695 1525
rect 699 1521 700 1525
rect 694 1520 700 1521
rect 758 1525 764 1526
rect 758 1521 759 1525
rect 763 1521 764 1525
rect 758 1520 764 1521
rect 350 1515 356 1516
rect 360 1515 362 1520
rect 408 1515 410 1520
rect 456 1515 458 1520
rect 512 1515 514 1520
rect 568 1515 570 1520
rect 632 1515 634 1520
rect 696 1515 698 1520
rect 760 1515 762 1520
rect 167 1514 171 1515
rect 167 1508 171 1510
rect 215 1514 219 1515
rect 215 1509 219 1510
rect 223 1514 227 1515
rect 223 1508 227 1510
rect 263 1514 267 1515
rect 263 1509 267 1510
rect 295 1514 299 1515
rect 295 1508 299 1510
rect 311 1514 315 1515
rect 350 1511 351 1515
rect 355 1511 356 1515
rect 350 1510 356 1511
rect 359 1514 363 1515
rect 311 1509 315 1510
rect 359 1509 363 1510
rect 375 1514 379 1515
rect 375 1508 379 1510
rect 407 1514 411 1515
rect 407 1509 411 1510
rect 455 1514 459 1515
rect 455 1508 459 1510
rect 511 1514 515 1515
rect 511 1509 515 1510
rect 527 1514 531 1515
rect 527 1508 531 1510
rect 567 1514 571 1515
rect 567 1509 571 1510
rect 599 1514 603 1515
rect 599 1508 603 1510
rect 631 1514 635 1515
rect 631 1509 635 1510
rect 671 1514 675 1515
rect 671 1508 675 1510
rect 695 1514 699 1515
rect 695 1509 699 1510
rect 743 1514 747 1515
rect 743 1508 747 1510
rect 759 1514 763 1515
rect 759 1509 763 1510
rect 166 1507 172 1508
rect 166 1503 167 1507
rect 171 1503 172 1507
rect 166 1502 172 1503
rect 222 1507 228 1508
rect 222 1503 223 1507
rect 227 1503 228 1507
rect 222 1502 228 1503
rect 294 1507 300 1508
rect 294 1503 295 1507
rect 299 1503 300 1507
rect 294 1502 300 1503
rect 374 1507 380 1508
rect 374 1503 375 1507
rect 379 1503 380 1507
rect 374 1502 380 1503
rect 454 1507 460 1508
rect 454 1503 455 1507
rect 459 1503 460 1507
rect 454 1502 460 1503
rect 526 1507 532 1508
rect 526 1503 527 1507
rect 531 1503 532 1507
rect 526 1502 532 1503
rect 598 1507 604 1508
rect 598 1503 599 1507
rect 603 1503 604 1507
rect 598 1502 604 1503
rect 670 1507 676 1508
rect 670 1503 671 1507
rect 675 1503 676 1507
rect 670 1502 676 1503
rect 742 1507 748 1508
rect 742 1503 743 1507
rect 747 1503 748 1507
rect 742 1502 748 1503
rect 542 1499 548 1500
rect 542 1495 543 1499
rect 547 1495 548 1499
rect 542 1494 548 1495
rect 182 1491 188 1492
rect 166 1490 172 1491
rect 166 1486 167 1490
rect 171 1486 172 1490
rect 182 1487 183 1491
rect 187 1487 188 1491
rect 182 1486 188 1487
rect 222 1490 228 1491
rect 222 1486 223 1490
rect 227 1486 228 1490
rect 166 1485 172 1486
rect 150 1483 156 1484
rect 150 1479 151 1483
rect 155 1479 156 1483
rect 150 1478 156 1479
rect 168 1475 170 1485
rect 111 1474 115 1475
rect 111 1469 115 1470
rect 135 1474 139 1475
rect 135 1469 139 1470
rect 167 1474 171 1475
rect 167 1469 171 1470
rect 112 1461 114 1469
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 136 1459 138 1469
rect 168 1459 170 1469
rect 184 1464 186 1486
rect 222 1485 228 1486
rect 294 1490 300 1491
rect 294 1486 295 1490
rect 299 1486 300 1490
rect 294 1485 300 1486
rect 374 1490 380 1491
rect 374 1486 375 1490
rect 379 1486 380 1490
rect 374 1485 380 1486
rect 454 1490 460 1491
rect 454 1486 455 1490
rect 459 1486 460 1490
rect 454 1485 460 1486
rect 526 1490 532 1491
rect 526 1486 527 1490
rect 531 1486 532 1490
rect 526 1485 532 1486
rect 224 1475 226 1485
rect 238 1475 244 1476
rect 296 1475 298 1485
rect 376 1475 378 1485
rect 456 1475 458 1485
rect 528 1475 530 1485
rect 223 1474 227 1475
rect 238 1471 239 1475
rect 243 1471 244 1475
rect 238 1470 244 1471
rect 295 1474 299 1475
rect 223 1469 227 1470
rect 182 1463 188 1464
rect 182 1459 183 1463
rect 187 1459 188 1463
rect 224 1459 226 1469
rect 110 1455 116 1456
rect 134 1458 140 1459
rect 134 1454 135 1458
rect 139 1454 140 1458
rect 134 1453 140 1454
rect 166 1458 172 1459
rect 182 1458 188 1459
rect 222 1458 228 1459
rect 166 1454 167 1458
rect 171 1454 172 1458
rect 166 1453 172 1454
rect 222 1454 223 1458
rect 227 1454 228 1458
rect 222 1453 228 1454
rect 240 1448 242 1470
rect 295 1469 299 1470
rect 375 1474 379 1475
rect 375 1469 379 1470
rect 455 1474 459 1475
rect 455 1469 459 1470
rect 527 1474 531 1475
rect 527 1469 531 1470
rect 296 1459 298 1469
rect 376 1459 378 1469
rect 456 1459 458 1469
rect 462 1463 468 1464
rect 462 1459 463 1463
rect 467 1459 468 1463
rect 528 1459 530 1469
rect 544 1464 546 1494
rect 772 1492 774 1526
rect 830 1525 836 1526
rect 830 1521 831 1525
rect 835 1521 836 1525
rect 830 1520 836 1521
rect 832 1515 834 1520
rect 815 1514 819 1515
rect 815 1508 819 1510
rect 831 1514 835 1515
rect 831 1509 835 1510
rect 879 1514 883 1515
rect 879 1508 883 1510
rect 814 1507 820 1508
rect 814 1503 815 1507
rect 819 1503 820 1507
rect 814 1502 820 1503
rect 878 1507 884 1508
rect 878 1503 879 1507
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 896 1500 898 1542
rect 918 1538 919 1542
rect 923 1538 924 1542
rect 918 1537 924 1538
rect 1006 1542 1012 1543
rect 1006 1538 1007 1542
rect 1011 1538 1012 1542
rect 1006 1537 1012 1538
rect 1094 1542 1100 1543
rect 1094 1538 1095 1542
rect 1099 1538 1100 1542
rect 1094 1537 1100 1538
rect 1182 1542 1188 1543
rect 1210 1542 1216 1543
rect 1262 1542 1268 1543
rect 1182 1538 1183 1542
rect 1187 1538 1188 1542
rect 1182 1537 1188 1538
rect 1262 1538 1263 1542
rect 1267 1538 1268 1542
rect 1262 1537 1268 1538
rect 958 1531 964 1532
rect 958 1527 959 1531
rect 963 1527 964 1531
rect 958 1526 964 1527
rect 1279 1531 1285 1532
rect 1279 1527 1280 1531
rect 1284 1530 1285 1531
rect 1288 1530 1290 1562
rect 1352 1559 1354 1569
rect 1335 1558 1339 1559
rect 1335 1553 1339 1554
rect 1351 1558 1355 1559
rect 1351 1553 1355 1554
rect 1326 1547 1332 1548
rect 1326 1543 1327 1547
rect 1331 1543 1332 1547
rect 1336 1543 1338 1553
rect 1364 1548 1366 1578
rect 1414 1574 1420 1575
rect 1414 1570 1415 1574
rect 1419 1570 1420 1574
rect 1414 1569 1420 1570
rect 1416 1559 1418 1569
rect 1432 1568 1434 1606
rect 1478 1605 1484 1606
rect 1478 1601 1479 1605
rect 1483 1601 1484 1605
rect 1478 1600 1484 1601
rect 1471 1598 1475 1599
rect 1471 1592 1475 1594
rect 1479 1598 1483 1600
rect 1479 1593 1483 1594
rect 1527 1598 1531 1599
rect 1527 1592 1531 1594
rect 1470 1591 1476 1592
rect 1470 1587 1471 1591
rect 1475 1587 1476 1591
rect 1470 1586 1476 1587
rect 1526 1591 1532 1592
rect 1526 1587 1527 1591
rect 1531 1587 1532 1591
rect 1526 1586 1532 1587
rect 1548 1584 1550 1642
rect 1559 1638 1563 1639
rect 1559 1633 1563 1634
rect 1560 1623 1562 1633
rect 1576 1628 1578 1658
rect 1582 1654 1588 1655
rect 1582 1650 1583 1654
rect 1587 1650 1588 1654
rect 1582 1649 1588 1650
rect 1622 1654 1628 1655
rect 1622 1650 1623 1654
rect 1627 1650 1628 1654
rect 1622 1649 1628 1650
rect 1584 1639 1586 1649
rect 1624 1639 1626 1649
rect 1583 1638 1587 1639
rect 1583 1633 1587 1634
rect 1623 1638 1627 1639
rect 1623 1633 1627 1634
rect 1574 1627 1580 1628
rect 1574 1623 1575 1627
rect 1579 1623 1580 1627
rect 1624 1623 1626 1633
rect 1640 1628 1642 1658
rect 1662 1652 1668 1653
rect 1662 1648 1663 1652
rect 1667 1648 1668 1652
rect 1662 1647 1668 1648
rect 1664 1639 1666 1647
rect 1663 1638 1667 1639
rect 1663 1633 1667 1634
rect 1638 1627 1644 1628
rect 1638 1623 1639 1627
rect 1643 1623 1644 1627
rect 1664 1625 1666 1633
rect 1558 1622 1564 1623
rect 1574 1622 1580 1623
rect 1622 1622 1628 1623
rect 1638 1622 1644 1623
rect 1662 1624 1668 1625
rect 1558 1618 1559 1622
rect 1563 1618 1564 1622
rect 1558 1617 1564 1618
rect 1622 1618 1623 1622
rect 1627 1618 1628 1622
rect 1662 1620 1663 1624
rect 1667 1620 1668 1624
rect 1662 1619 1668 1620
rect 1622 1617 1628 1618
rect 1638 1611 1644 1612
rect 1638 1607 1639 1611
rect 1643 1607 1644 1611
rect 1638 1606 1644 1607
rect 1662 1607 1668 1608
rect 1558 1605 1564 1606
rect 1558 1601 1559 1605
rect 1563 1601 1564 1605
rect 1558 1600 1564 1601
rect 1622 1605 1628 1606
rect 1622 1601 1623 1605
rect 1627 1601 1628 1605
rect 1622 1600 1628 1601
rect 1559 1598 1563 1600
rect 1559 1593 1563 1594
rect 1583 1598 1587 1599
rect 1583 1592 1587 1594
rect 1623 1598 1627 1600
rect 1623 1592 1627 1594
rect 1582 1591 1588 1592
rect 1582 1587 1583 1591
rect 1587 1587 1588 1591
rect 1582 1586 1588 1587
rect 1622 1591 1628 1592
rect 1622 1587 1623 1591
rect 1627 1587 1628 1591
rect 1622 1586 1628 1587
rect 1482 1583 1488 1584
rect 1482 1579 1483 1583
rect 1487 1579 1488 1583
rect 1482 1578 1488 1579
rect 1546 1583 1552 1584
rect 1546 1579 1547 1583
rect 1551 1579 1552 1583
rect 1546 1578 1552 1579
rect 1470 1574 1476 1575
rect 1470 1570 1471 1574
rect 1475 1570 1476 1574
rect 1470 1569 1476 1570
rect 1430 1567 1436 1568
rect 1430 1563 1431 1567
rect 1435 1563 1436 1567
rect 1430 1562 1436 1563
rect 1472 1559 1474 1569
rect 1484 1560 1486 1578
rect 1526 1574 1532 1575
rect 1526 1570 1527 1574
rect 1531 1570 1532 1574
rect 1526 1569 1532 1570
rect 1582 1574 1588 1575
rect 1582 1570 1583 1574
rect 1587 1570 1588 1574
rect 1582 1569 1588 1570
rect 1622 1574 1628 1575
rect 1622 1570 1623 1574
rect 1627 1570 1628 1574
rect 1622 1569 1628 1570
rect 1482 1559 1488 1560
rect 1528 1559 1530 1569
rect 1584 1559 1586 1569
rect 1598 1567 1604 1568
rect 1598 1563 1599 1567
rect 1603 1563 1604 1567
rect 1598 1562 1604 1563
rect 1407 1558 1411 1559
rect 1407 1553 1411 1554
rect 1415 1558 1419 1559
rect 1415 1553 1419 1554
rect 1471 1558 1475 1559
rect 1482 1555 1483 1559
rect 1487 1555 1488 1559
rect 1482 1554 1488 1555
rect 1527 1558 1531 1559
rect 1471 1553 1475 1554
rect 1527 1553 1531 1554
rect 1583 1558 1587 1559
rect 1583 1553 1587 1554
rect 1370 1551 1376 1552
rect 1362 1547 1368 1548
rect 1362 1543 1363 1547
rect 1367 1543 1368 1547
rect 1370 1547 1371 1551
rect 1375 1547 1376 1551
rect 1370 1546 1376 1547
rect 1326 1542 1332 1543
rect 1334 1542 1340 1543
rect 1362 1542 1368 1543
rect 1284 1528 1290 1530
rect 1284 1527 1285 1528
rect 1279 1526 1285 1527
rect 918 1525 924 1526
rect 918 1521 919 1525
rect 923 1521 924 1525
rect 918 1520 924 1521
rect 920 1515 922 1520
rect 919 1514 923 1515
rect 919 1509 923 1510
rect 943 1514 947 1515
rect 943 1508 947 1510
rect 942 1507 948 1508
rect 942 1503 943 1507
rect 947 1503 948 1507
rect 942 1502 948 1503
rect 894 1499 900 1500
rect 894 1495 895 1499
rect 899 1495 900 1499
rect 894 1494 900 1495
rect 770 1491 776 1492
rect 598 1490 604 1491
rect 598 1486 599 1490
rect 603 1486 604 1490
rect 598 1485 604 1486
rect 670 1490 676 1491
rect 670 1486 671 1490
rect 675 1486 676 1490
rect 670 1485 676 1486
rect 742 1490 748 1491
rect 742 1486 743 1490
rect 747 1486 748 1490
rect 770 1487 771 1491
rect 775 1487 776 1491
rect 770 1486 776 1487
rect 814 1490 820 1491
rect 814 1486 815 1490
rect 819 1486 820 1490
rect 742 1485 748 1486
rect 814 1485 820 1486
rect 878 1490 884 1491
rect 878 1486 879 1490
rect 883 1486 884 1490
rect 878 1485 884 1486
rect 942 1490 948 1491
rect 942 1486 943 1490
rect 947 1486 948 1490
rect 942 1485 948 1486
rect 600 1475 602 1485
rect 672 1475 674 1485
rect 744 1475 746 1485
rect 798 1483 804 1484
rect 798 1479 799 1483
rect 803 1479 804 1483
rect 798 1478 804 1479
rect 599 1474 603 1475
rect 599 1469 603 1470
rect 663 1474 667 1475
rect 663 1469 667 1470
rect 671 1474 675 1475
rect 671 1469 675 1470
rect 719 1474 723 1475
rect 719 1469 723 1470
rect 743 1474 747 1475
rect 743 1469 747 1470
rect 783 1474 787 1475
rect 783 1469 787 1470
rect 542 1463 548 1464
rect 542 1459 543 1463
rect 547 1459 548 1463
rect 600 1459 602 1469
rect 664 1459 666 1469
rect 720 1459 722 1469
rect 784 1459 786 1469
rect 294 1458 300 1459
rect 294 1454 295 1458
rect 299 1454 300 1458
rect 294 1453 300 1454
rect 374 1458 380 1459
rect 374 1454 375 1458
rect 379 1454 380 1458
rect 374 1453 380 1454
rect 454 1458 460 1459
rect 462 1458 468 1459
rect 526 1458 532 1459
rect 542 1458 548 1459
rect 598 1458 604 1459
rect 454 1454 455 1458
rect 459 1454 460 1458
rect 454 1453 460 1454
rect 150 1447 156 1448
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 150 1443 151 1447
rect 155 1443 156 1447
rect 150 1442 156 1443
rect 238 1447 244 1448
rect 238 1443 239 1447
rect 243 1443 244 1447
rect 238 1442 244 1443
rect 110 1438 116 1439
rect 134 1441 140 1442
rect 112 1431 114 1438
rect 134 1437 135 1441
rect 139 1437 140 1441
rect 134 1436 140 1437
rect 136 1431 138 1436
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 135 1430 139 1431
rect 112 1422 114 1425
rect 135 1424 139 1426
rect 134 1423 140 1424
rect 110 1421 116 1422
rect 110 1417 111 1421
rect 115 1417 116 1421
rect 134 1419 135 1423
rect 139 1419 140 1423
rect 134 1418 140 1419
rect 110 1416 116 1417
rect 134 1406 140 1407
rect 110 1404 116 1405
rect 110 1400 111 1404
rect 115 1400 116 1404
rect 134 1402 135 1406
rect 139 1402 140 1406
rect 134 1401 140 1402
rect 110 1399 116 1400
rect 112 1391 114 1399
rect 136 1391 138 1401
rect 152 1400 154 1442
rect 166 1441 172 1442
rect 166 1437 167 1441
rect 171 1437 172 1441
rect 166 1436 172 1437
rect 222 1441 228 1442
rect 222 1437 223 1441
rect 227 1437 228 1441
rect 222 1436 228 1437
rect 294 1441 300 1442
rect 294 1437 295 1441
rect 299 1437 300 1441
rect 294 1436 300 1437
rect 374 1441 380 1442
rect 374 1437 375 1441
rect 379 1437 380 1441
rect 374 1436 380 1437
rect 454 1441 460 1442
rect 454 1437 455 1441
rect 459 1437 460 1441
rect 454 1436 460 1437
rect 168 1431 170 1436
rect 224 1431 226 1436
rect 296 1431 298 1436
rect 376 1431 378 1436
rect 456 1431 458 1436
rect 167 1430 171 1431
rect 167 1424 171 1426
rect 215 1430 219 1431
rect 215 1424 219 1426
rect 223 1430 227 1431
rect 223 1425 227 1426
rect 287 1430 291 1431
rect 287 1424 291 1426
rect 295 1430 299 1431
rect 295 1425 299 1426
rect 359 1430 363 1431
rect 359 1424 363 1426
rect 375 1430 379 1431
rect 375 1425 379 1426
rect 439 1430 443 1431
rect 439 1424 443 1426
rect 455 1430 459 1431
rect 455 1425 459 1426
rect 166 1423 172 1424
rect 166 1419 167 1423
rect 171 1419 172 1423
rect 166 1418 172 1419
rect 214 1423 220 1424
rect 214 1419 215 1423
rect 219 1419 220 1423
rect 214 1418 220 1419
rect 286 1423 292 1424
rect 286 1419 287 1423
rect 291 1419 292 1423
rect 286 1418 292 1419
rect 358 1423 364 1424
rect 358 1419 359 1423
rect 363 1419 364 1423
rect 358 1418 364 1419
rect 438 1423 444 1424
rect 438 1419 439 1423
rect 443 1419 444 1423
rect 438 1418 444 1419
rect 230 1415 236 1416
rect 230 1411 231 1415
rect 235 1411 236 1415
rect 230 1410 236 1411
rect 455 1415 461 1416
rect 455 1411 456 1415
rect 460 1414 461 1415
rect 464 1414 466 1458
rect 526 1454 527 1458
rect 531 1454 532 1458
rect 526 1453 532 1454
rect 598 1454 599 1458
rect 603 1454 604 1458
rect 598 1453 604 1454
rect 662 1458 668 1459
rect 662 1454 663 1458
rect 667 1454 668 1458
rect 662 1453 668 1454
rect 718 1458 724 1459
rect 718 1454 719 1458
rect 723 1454 724 1458
rect 718 1453 724 1454
rect 782 1458 788 1459
rect 782 1454 783 1458
rect 787 1454 788 1458
rect 782 1453 788 1454
rect 800 1448 802 1478
rect 816 1475 818 1485
rect 880 1475 882 1485
rect 944 1475 946 1485
rect 960 1484 962 1526
rect 1006 1525 1012 1526
rect 1006 1521 1007 1525
rect 1011 1521 1012 1525
rect 1006 1520 1012 1521
rect 1094 1525 1100 1526
rect 1094 1521 1095 1525
rect 1099 1521 1100 1525
rect 1094 1520 1100 1521
rect 1182 1525 1188 1526
rect 1182 1521 1183 1525
rect 1187 1521 1188 1525
rect 1182 1520 1188 1521
rect 1262 1525 1268 1526
rect 1262 1521 1263 1525
rect 1267 1521 1268 1525
rect 1262 1520 1268 1521
rect 1008 1515 1010 1520
rect 1096 1515 1098 1520
rect 1184 1515 1186 1520
rect 1264 1515 1266 1520
rect 1328 1516 1330 1542
rect 1334 1538 1335 1542
rect 1339 1538 1340 1542
rect 1334 1537 1340 1538
rect 1372 1532 1374 1546
rect 1408 1543 1410 1553
rect 1472 1543 1474 1553
rect 1528 1543 1530 1553
rect 1584 1543 1586 1553
rect 1406 1542 1412 1543
rect 1406 1538 1407 1542
rect 1411 1538 1412 1542
rect 1406 1537 1412 1538
rect 1470 1542 1476 1543
rect 1470 1538 1471 1542
rect 1475 1538 1476 1542
rect 1470 1537 1476 1538
rect 1526 1542 1532 1543
rect 1526 1538 1527 1542
rect 1531 1538 1532 1542
rect 1526 1537 1532 1538
rect 1582 1542 1588 1543
rect 1582 1538 1583 1542
rect 1587 1538 1588 1542
rect 1582 1537 1588 1538
rect 1600 1532 1602 1562
rect 1624 1559 1626 1569
rect 1640 1568 1642 1606
rect 1662 1603 1663 1607
rect 1667 1603 1668 1607
rect 1662 1602 1668 1603
rect 1664 1599 1666 1602
rect 1663 1598 1667 1599
rect 1663 1593 1667 1594
rect 1664 1590 1666 1593
rect 1662 1589 1668 1590
rect 1662 1585 1663 1589
rect 1667 1585 1668 1589
rect 1662 1584 1668 1585
rect 1662 1572 1668 1573
rect 1662 1568 1663 1572
rect 1667 1568 1668 1572
rect 1638 1567 1644 1568
rect 1662 1567 1668 1568
rect 1638 1563 1639 1567
rect 1643 1563 1644 1567
rect 1638 1562 1644 1563
rect 1664 1559 1666 1567
rect 1623 1558 1627 1559
rect 1623 1553 1627 1554
rect 1663 1558 1667 1559
rect 1663 1553 1667 1554
rect 1624 1543 1626 1553
rect 1664 1545 1666 1553
rect 1662 1544 1668 1545
rect 1622 1542 1628 1543
rect 1622 1538 1623 1542
rect 1627 1538 1628 1542
rect 1662 1540 1663 1544
rect 1667 1540 1668 1544
rect 1662 1539 1668 1540
rect 1622 1537 1628 1538
rect 1370 1531 1376 1532
rect 1370 1527 1371 1531
rect 1375 1527 1376 1531
rect 1370 1526 1376 1527
rect 1598 1531 1604 1532
rect 1598 1527 1599 1531
rect 1603 1527 1604 1531
rect 1598 1526 1604 1527
rect 1638 1531 1644 1532
rect 1638 1527 1639 1531
rect 1643 1527 1644 1531
rect 1638 1526 1644 1527
rect 1662 1527 1668 1528
rect 1334 1525 1340 1526
rect 1334 1521 1335 1525
rect 1339 1521 1340 1525
rect 1334 1520 1340 1521
rect 1406 1525 1412 1526
rect 1406 1521 1407 1525
rect 1411 1521 1412 1525
rect 1406 1520 1412 1521
rect 1470 1525 1476 1526
rect 1470 1521 1471 1525
rect 1475 1521 1476 1525
rect 1470 1520 1476 1521
rect 1526 1525 1532 1526
rect 1526 1521 1527 1525
rect 1531 1521 1532 1525
rect 1526 1520 1532 1521
rect 1582 1525 1588 1526
rect 1582 1521 1583 1525
rect 1587 1521 1588 1525
rect 1582 1520 1588 1521
rect 1622 1525 1628 1526
rect 1622 1521 1623 1525
rect 1627 1521 1628 1525
rect 1622 1520 1628 1521
rect 1326 1515 1332 1516
rect 1336 1515 1338 1520
rect 1408 1515 1410 1520
rect 1472 1515 1474 1520
rect 1528 1515 1530 1520
rect 1584 1515 1586 1520
rect 1624 1515 1626 1520
rect 1007 1514 1011 1515
rect 1007 1508 1011 1510
rect 1063 1514 1067 1515
rect 1063 1508 1067 1510
rect 1095 1514 1099 1515
rect 1095 1509 1099 1510
rect 1111 1514 1115 1515
rect 1111 1508 1115 1510
rect 1151 1514 1155 1515
rect 1151 1508 1155 1510
rect 1183 1514 1187 1515
rect 1183 1508 1187 1510
rect 1215 1514 1219 1515
rect 1215 1508 1219 1510
rect 1255 1514 1259 1515
rect 1255 1508 1259 1510
rect 1263 1514 1267 1515
rect 1263 1509 1267 1510
rect 1295 1514 1299 1515
rect 1326 1511 1327 1515
rect 1331 1511 1332 1515
rect 1326 1510 1332 1511
rect 1335 1514 1339 1515
rect 1295 1508 1299 1510
rect 1335 1509 1339 1510
rect 1351 1514 1355 1515
rect 1351 1508 1355 1510
rect 1407 1514 1411 1515
rect 1407 1509 1411 1510
rect 1415 1514 1419 1515
rect 1415 1508 1419 1510
rect 1471 1514 1475 1515
rect 1471 1509 1475 1510
rect 1487 1514 1491 1515
rect 1487 1508 1491 1510
rect 1527 1514 1531 1515
rect 1527 1509 1531 1510
rect 1567 1514 1571 1515
rect 1567 1508 1571 1510
rect 1583 1514 1587 1515
rect 1583 1509 1587 1510
rect 1623 1514 1627 1515
rect 1623 1508 1627 1510
rect 1006 1507 1012 1508
rect 1006 1503 1007 1507
rect 1011 1503 1012 1507
rect 1006 1502 1012 1503
rect 1062 1507 1068 1508
rect 1062 1503 1063 1507
rect 1067 1503 1068 1507
rect 1062 1502 1068 1503
rect 1110 1507 1116 1508
rect 1110 1503 1111 1507
rect 1115 1503 1116 1507
rect 1110 1502 1116 1503
rect 1150 1507 1156 1508
rect 1150 1503 1151 1507
rect 1155 1503 1156 1507
rect 1150 1502 1156 1503
rect 1182 1507 1188 1508
rect 1182 1503 1183 1507
rect 1187 1503 1188 1507
rect 1182 1502 1188 1503
rect 1214 1507 1220 1508
rect 1214 1503 1215 1507
rect 1219 1503 1220 1507
rect 1214 1502 1220 1503
rect 1254 1507 1260 1508
rect 1254 1503 1255 1507
rect 1259 1503 1260 1507
rect 1254 1502 1260 1503
rect 1294 1507 1300 1508
rect 1294 1503 1295 1507
rect 1299 1503 1300 1507
rect 1294 1502 1300 1503
rect 1350 1507 1356 1508
rect 1350 1503 1351 1507
rect 1355 1503 1356 1507
rect 1350 1502 1356 1503
rect 1414 1507 1420 1508
rect 1414 1503 1415 1507
rect 1419 1503 1420 1507
rect 1414 1502 1420 1503
rect 1486 1507 1492 1508
rect 1486 1503 1487 1507
rect 1491 1503 1492 1507
rect 1486 1502 1492 1503
rect 1566 1507 1572 1508
rect 1566 1503 1567 1507
rect 1571 1503 1572 1507
rect 1566 1502 1572 1503
rect 1622 1507 1628 1508
rect 1622 1503 1623 1507
rect 1627 1503 1628 1507
rect 1622 1502 1628 1503
rect 974 1499 980 1500
rect 974 1495 975 1499
rect 979 1495 980 1499
rect 974 1494 980 1495
rect 1230 1499 1236 1500
rect 1230 1495 1231 1499
rect 1235 1495 1236 1499
rect 1230 1494 1236 1495
rect 958 1483 964 1484
rect 958 1479 959 1483
rect 963 1479 964 1483
rect 958 1478 964 1479
rect 815 1474 819 1475
rect 815 1469 819 1470
rect 847 1474 851 1475
rect 847 1469 851 1470
rect 879 1474 883 1475
rect 879 1469 883 1470
rect 903 1474 907 1475
rect 903 1469 907 1470
rect 943 1474 947 1475
rect 943 1469 947 1470
rect 959 1474 963 1475
rect 959 1469 963 1470
rect 848 1459 850 1469
rect 904 1459 906 1469
rect 960 1459 962 1469
rect 976 1464 978 1494
rect 1006 1490 1012 1491
rect 1006 1486 1007 1490
rect 1011 1486 1012 1490
rect 1006 1485 1012 1486
rect 1062 1490 1068 1491
rect 1062 1486 1063 1490
rect 1067 1486 1068 1490
rect 1062 1485 1068 1486
rect 1110 1490 1116 1491
rect 1110 1486 1111 1490
rect 1115 1486 1116 1490
rect 1110 1485 1116 1486
rect 1150 1490 1156 1491
rect 1150 1486 1151 1490
rect 1155 1486 1156 1490
rect 1150 1485 1156 1486
rect 1182 1490 1188 1491
rect 1182 1486 1183 1490
rect 1187 1486 1188 1490
rect 1182 1485 1188 1486
rect 1214 1490 1220 1491
rect 1214 1486 1215 1490
rect 1219 1486 1220 1490
rect 1214 1485 1220 1486
rect 1008 1475 1010 1485
rect 1026 1483 1032 1484
rect 1026 1479 1027 1483
rect 1031 1479 1032 1483
rect 1026 1478 1032 1479
rect 1007 1474 1011 1475
rect 1007 1469 1011 1470
rect 1015 1474 1019 1475
rect 1015 1469 1019 1470
rect 974 1463 980 1464
rect 974 1459 975 1463
rect 979 1459 980 1463
rect 1016 1459 1018 1469
rect 846 1458 852 1459
rect 846 1454 847 1458
rect 851 1454 852 1458
rect 846 1453 852 1454
rect 902 1458 908 1459
rect 902 1454 903 1458
rect 907 1454 908 1458
rect 902 1453 908 1454
rect 958 1458 964 1459
rect 974 1458 980 1459
rect 1014 1458 1020 1459
rect 958 1454 959 1458
rect 963 1454 964 1458
rect 958 1453 964 1454
rect 1014 1454 1015 1458
rect 1019 1454 1020 1458
rect 1014 1453 1020 1454
rect 1028 1448 1030 1478
rect 1064 1475 1066 1485
rect 1112 1475 1114 1485
rect 1152 1475 1154 1485
rect 1184 1475 1186 1485
rect 1216 1475 1218 1485
rect 1232 1476 1234 1494
rect 1254 1490 1260 1491
rect 1254 1486 1255 1490
rect 1259 1486 1260 1490
rect 1254 1485 1260 1486
rect 1294 1490 1300 1491
rect 1294 1486 1295 1490
rect 1299 1486 1300 1490
rect 1294 1485 1300 1486
rect 1350 1490 1356 1491
rect 1350 1486 1351 1490
rect 1355 1486 1356 1490
rect 1350 1485 1356 1486
rect 1414 1490 1420 1491
rect 1414 1486 1415 1490
rect 1419 1486 1420 1490
rect 1414 1485 1420 1486
rect 1486 1490 1492 1491
rect 1486 1486 1487 1490
rect 1491 1486 1492 1490
rect 1486 1485 1492 1486
rect 1566 1490 1572 1491
rect 1566 1486 1567 1490
rect 1571 1486 1572 1490
rect 1566 1485 1572 1486
rect 1622 1490 1628 1491
rect 1622 1486 1623 1490
rect 1627 1486 1628 1490
rect 1622 1485 1628 1486
rect 1230 1475 1236 1476
rect 1256 1475 1258 1485
rect 1296 1475 1298 1485
rect 1352 1475 1354 1485
rect 1416 1475 1418 1485
rect 1488 1475 1490 1485
rect 1494 1475 1500 1476
rect 1568 1475 1570 1485
rect 1624 1475 1626 1485
rect 1640 1484 1642 1526
rect 1662 1523 1663 1527
rect 1667 1523 1668 1527
rect 1662 1522 1668 1523
rect 1664 1515 1666 1522
rect 1663 1514 1667 1515
rect 1663 1509 1667 1510
rect 1664 1506 1666 1509
rect 1662 1505 1668 1506
rect 1662 1501 1663 1505
rect 1667 1501 1668 1505
rect 1662 1500 1668 1501
rect 1662 1488 1668 1489
rect 1662 1484 1663 1488
rect 1667 1484 1668 1488
rect 1638 1483 1644 1484
rect 1662 1483 1668 1484
rect 1638 1479 1639 1483
rect 1643 1479 1644 1483
rect 1638 1478 1644 1479
rect 1664 1475 1666 1483
rect 1063 1474 1067 1475
rect 1063 1469 1067 1470
rect 1071 1474 1075 1475
rect 1071 1469 1075 1470
rect 1111 1474 1115 1475
rect 1111 1469 1115 1470
rect 1119 1474 1123 1475
rect 1119 1469 1123 1470
rect 1151 1474 1155 1475
rect 1151 1469 1155 1470
rect 1159 1474 1163 1475
rect 1159 1469 1163 1470
rect 1183 1474 1187 1475
rect 1183 1469 1187 1470
rect 1207 1474 1211 1475
rect 1207 1469 1211 1470
rect 1215 1474 1219 1475
rect 1230 1471 1231 1475
rect 1235 1471 1236 1475
rect 1230 1470 1236 1471
rect 1255 1474 1259 1475
rect 1215 1469 1219 1470
rect 1255 1469 1259 1470
rect 1263 1474 1267 1475
rect 1263 1469 1267 1470
rect 1295 1474 1299 1475
rect 1295 1469 1299 1470
rect 1327 1474 1331 1475
rect 1327 1469 1331 1470
rect 1351 1474 1355 1475
rect 1351 1469 1355 1470
rect 1399 1474 1403 1475
rect 1399 1469 1403 1470
rect 1415 1474 1419 1475
rect 1415 1469 1419 1470
rect 1479 1474 1483 1475
rect 1479 1469 1483 1470
rect 1487 1474 1491 1475
rect 1494 1471 1495 1475
rect 1499 1471 1500 1475
rect 1494 1470 1500 1471
rect 1559 1474 1563 1475
rect 1487 1469 1491 1470
rect 1072 1459 1074 1469
rect 1120 1459 1122 1469
rect 1146 1463 1152 1464
rect 1146 1459 1147 1463
rect 1151 1459 1152 1463
rect 1160 1459 1162 1469
rect 1208 1459 1210 1469
rect 1264 1459 1266 1469
rect 1328 1459 1330 1469
rect 1400 1459 1402 1469
rect 1480 1459 1482 1469
rect 1070 1458 1076 1459
rect 1070 1454 1071 1458
rect 1075 1454 1076 1458
rect 1070 1453 1076 1454
rect 1118 1458 1124 1459
rect 1146 1458 1152 1459
rect 1158 1458 1164 1459
rect 1118 1454 1119 1458
rect 1123 1454 1124 1458
rect 1118 1453 1124 1454
rect 798 1447 804 1448
rect 798 1443 799 1447
rect 803 1443 804 1447
rect 798 1442 804 1443
rect 894 1447 900 1448
rect 894 1443 895 1447
rect 899 1443 900 1447
rect 894 1442 900 1443
rect 1026 1447 1032 1448
rect 1026 1443 1027 1447
rect 1031 1443 1032 1447
rect 1026 1442 1032 1443
rect 526 1441 532 1442
rect 526 1437 527 1441
rect 531 1437 532 1441
rect 526 1436 532 1437
rect 598 1441 604 1442
rect 598 1437 599 1441
rect 603 1437 604 1441
rect 598 1436 604 1437
rect 662 1441 668 1442
rect 662 1437 663 1441
rect 667 1437 668 1441
rect 662 1436 668 1437
rect 718 1441 724 1442
rect 718 1437 719 1441
rect 723 1437 724 1441
rect 718 1436 724 1437
rect 782 1441 788 1442
rect 782 1437 783 1441
rect 787 1437 788 1441
rect 782 1436 788 1437
rect 846 1441 852 1442
rect 846 1437 847 1441
rect 851 1437 852 1441
rect 846 1436 852 1437
rect 528 1431 530 1436
rect 600 1431 602 1436
rect 664 1431 666 1436
rect 720 1431 722 1436
rect 784 1431 786 1436
rect 848 1431 850 1436
rect 519 1430 523 1431
rect 519 1424 523 1426
rect 527 1430 531 1431
rect 527 1425 531 1426
rect 599 1430 603 1431
rect 599 1424 603 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 679 1430 683 1431
rect 679 1424 683 1426
rect 719 1430 723 1431
rect 719 1425 723 1426
rect 759 1430 763 1431
rect 759 1424 763 1426
rect 783 1430 787 1431
rect 783 1425 787 1426
rect 831 1430 835 1431
rect 831 1424 835 1426
rect 847 1430 851 1431
rect 847 1425 851 1426
rect 518 1423 524 1424
rect 518 1419 519 1423
rect 523 1419 524 1423
rect 518 1418 524 1419
rect 598 1423 604 1424
rect 598 1419 599 1423
rect 603 1419 604 1423
rect 598 1418 604 1419
rect 678 1423 684 1424
rect 678 1419 679 1423
rect 683 1419 684 1423
rect 678 1418 684 1419
rect 758 1423 764 1424
rect 758 1419 759 1423
rect 763 1419 764 1423
rect 758 1418 764 1419
rect 830 1423 836 1424
rect 830 1419 831 1423
rect 835 1419 836 1423
rect 830 1418 836 1419
rect 460 1412 466 1414
rect 750 1415 756 1416
rect 460 1411 461 1412
rect 455 1410 461 1411
rect 750 1411 751 1415
rect 755 1411 756 1415
rect 750 1410 756 1411
rect 770 1415 776 1416
rect 770 1411 771 1415
rect 775 1411 776 1415
rect 770 1410 776 1411
rect 166 1406 172 1407
rect 166 1402 167 1406
rect 171 1402 172 1406
rect 166 1401 172 1402
rect 214 1406 220 1407
rect 214 1402 215 1406
rect 219 1402 220 1406
rect 214 1401 220 1402
rect 150 1399 156 1400
rect 150 1395 151 1399
rect 155 1395 156 1399
rect 150 1394 156 1395
rect 168 1391 170 1401
rect 216 1391 218 1401
rect 111 1390 115 1391
rect 111 1385 115 1386
rect 135 1390 139 1391
rect 135 1385 139 1386
rect 167 1390 171 1391
rect 167 1385 171 1386
rect 215 1390 219 1391
rect 215 1385 219 1386
rect 223 1390 227 1391
rect 232 1388 234 1410
rect 286 1406 292 1407
rect 286 1402 287 1406
rect 291 1402 292 1406
rect 286 1401 292 1402
rect 358 1406 364 1407
rect 358 1402 359 1406
rect 363 1402 364 1406
rect 358 1401 364 1402
rect 438 1406 444 1407
rect 438 1402 439 1406
rect 443 1402 444 1406
rect 438 1401 444 1402
rect 518 1406 524 1407
rect 518 1402 519 1406
rect 523 1402 524 1406
rect 518 1401 524 1402
rect 598 1406 604 1407
rect 598 1402 599 1406
rect 603 1402 604 1406
rect 598 1401 604 1402
rect 678 1406 684 1407
rect 678 1402 679 1406
rect 683 1402 684 1406
rect 678 1401 684 1402
rect 242 1399 248 1400
rect 242 1395 243 1399
rect 247 1395 248 1399
rect 242 1394 248 1395
rect 223 1385 227 1386
rect 230 1387 236 1388
rect 112 1377 114 1385
rect 110 1376 116 1377
rect 110 1372 111 1376
rect 115 1372 116 1376
rect 136 1375 138 1385
rect 168 1375 170 1385
rect 224 1375 226 1385
rect 230 1383 231 1387
rect 235 1383 236 1387
rect 230 1382 236 1383
rect 110 1371 116 1372
rect 134 1374 140 1375
rect 134 1370 135 1374
rect 139 1370 140 1374
rect 134 1369 140 1370
rect 166 1374 172 1375
rect 166 1370 167 1374
rect 171 1370 172 1374
rect 166 1369 172 1370
rect 222 1374 228 1375
rect 222 1370 223 1374
rect 227 1370 228 1374
rect 222 1369 228 1370
rect 244 1364 246 1394
rect 288 1391 290 1401
rect 360 1391 362 1401
rect 440 1391 442 1401
rect 520 1391 522 1401
rect 600 1391 602 1401
rect 680 1391 682 1401
rect 287 1390 291 1391
rect 287 1385 291 1386
rect 359 1390 363 1391
rect 359 1385 363 1386
rect 431 1390 435 1391
rect 431 1385 435 1386
rect 439 1390 443 1391
rect 439 1385 443 1386
rect 503 1390 507 1391
rect 503 1385 507 1386
rect 519 1390 523 1391
rect 519 1385 523 1386
rect 583 1390 587 1391
rect 583 1385 587 1386
rect 599 1390 603 1391
rect 599 1385 603 1386
rect 663 1390 667 1391
rect 663 1385 667 1386
rect 679 1390 683 1391
rect 679 1385 683 1386
rect 743 1390 747 1391
rect 743 1385 747 1386
rect 288 1375 290 1385
rect 360 1375 362 1385
rect 432 1375 434 1385
rect 438 1379 444 1380
rect 438 1375 439 1379
rect 443 1375 444 1379
rect 504 1375 506 1385
rect 518 1379 524 1380
rect 518 1375 519 1379
rect 523 1375 524 1379
rect 584 1375 586 1385
rect 664 1375 666 1385
rect 744 1375 746 1385
rect 752 1380 754 1410
rect 758 1406 764 1407
rect 758 1402 759 1406
rect 763 1402 764 1406
rect 758 1401 764 1402
rect 760 1391 762 1401
rect 772 1392 774 1410
rect 830 1406 836 1407
rect 830 1402 831 1406
rect 835 1402 836 1406
rect 830 1401 836 1402
rect 770 1391 776 1392
rect 832 1391 834 1401
rect 896 1400 898 1442
rect 902 1441 908 1442
rect 902 1437 903 1441
rect 907 1437 908 1441
rect 902 1436 908 1437
rect 958 1441 964 1442
rect 958 1437 959 1441
rect 963 1437 964 1441
rect 958 1436 964 1437
rect 1014 1441 1020 1442
rect 1014 1437 1015 1441
rect 1019 1437 1020 1441
rect 1014 1436 1020 1437
rect 1070 1441 1076 1442
rect 1070 1437 1071 1441
rect 1075 1437 1076 1441
rect 1070 1436 1076 1437
rect 1118 1441 1124 1442
rect 1118 1437 1119 1441
rect 1123 1437 1124 1441
rect 1118 1436 1124 1437
rect 904 1431 906 1436
rect 960 1431 962 1436
rect 1016 1431 1018 1436
rect 1072 1431 1074 1436
rect 1120 1431 1122 1436
rect 1148 1432 1150 1458
rect 1158 1454 1159 1458
rect 1163 1454 1164 1458
rect 1158 1453 1164 1454
rect 1206 1458 1212 1459
rect 1206 1454 1207 1458
rect 1211 1454 1212 1458
rect 1206 1453 1212 1454
rect 1262 1458 1268 1459
rect 1262 1454 1263 1458
rect 1267 1454 1268 1458
rect 1262 1453 1268 1454
rect 1326 1458 1332 1459
rect 1326 1454 1327 1458
rect 1331 1454 1332 1458
rect 1326 1453 1332 1454
rect 1398 1458 1404 1459
rect 1398 1454 1399 1458
rect 1403 1454 1404 1458
rect 1398 1453 1404 1454
rect 1478 1458 1484 1459
rect 1478 1454 1479 1458
rect 1483 1454 1484 1458
rect 1478 1453 1484 1454
rect 1496 1448 1498 1470
rect 1559 1469 1563 1470
rect 1567 1474 1571 1475
rect 1567 1469 1571 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1663 1474 1667 1475
rect 1663 1469 1667 1470
rect 1560 1459 1562 1469
rect 1570 1463 1576 1464
rect 1570 1459 1571 1463
rect 1575 1459 1576 1463
rect 1624 1459 1626 1469
rect 1664 1461 1666 1469
rect 1662 1460 1668 1461
rect 1558 1458 1564 1459
rect 1570 1458 1576 1459
rect 1622 1458 1628 1459
rect 1558 1454 1559 1458
rect 1563 1454 1564 1458
rect 1558 1453 1564 1454
rect 1494 1447 1500 1448
rect 1494 1443 1495 1447
rect 1499 1443 1500 1447
rect 1494 1442 1500 1443
rect 1158 1441 1164 1442
rect 1158 1437 1159 1441
rect 1163 1437 1164 1441
rect 1158 1436 1164 1437
rect 1206 1441 1212 1442
rect 1206 1437 1207 1441
rect 1211 1437 1212 1441
rect 1206 1436 1212 1437
rect 1262 1441 1268 1442
rect 1262 1437 1263 1441
rect 1267 1437 1268 1441
rect 1262 1436 1268 1437
rect 1326 1441 1332 1442
rect 1326 1437 1327 1441
rect 1331 1437 1332 1441
rect 1326 1436 1332 1437
rect 1398 1441 1404 1442
rect 1398 1437 1399 1441
rect 1403 1437 1404 1441
rect 1398 1436 1404 1437
rect 1478 1441 1484 1442
rect 1478 1437 1479 1441
rect 1483 1437 1484 1441
rect 1478 1436 1484 1437
rect 1558 1441 1564 1442
rect 1558 1437 1559 1441
rect 1563 1437 1564 1441
rect 1558 1436 1564 1437
rect 1146 1431 1152 1432
rect 1160 1431 1162 1436
rect 1208 1431 1210 1436
rect 1264 1431 1266 1436
rect 1328 1431 1330 1436
rect 1400 1431 1402 1436
rect 1480 1431 1482 1436
rect 1522 1435 1528 1436
rect 1522 1431 1523 1435
rect 1527 1431 1528 1435
rect 1560 1431 1562 1436
rect 903 1430 907 1431
rect 903 1424 907 1426
rect 959 1430 963 1431
rect 959 1425 963 1426
rect 967 1430 971 1431
rect 967 1424 971 1426
rect 1015 1430 1019 1431
rect 1015 1425 1019 1426
rect 1031 1430 1035 1431
rect 1031 1424 1035 1426
rect 1071 1430 1075 1431
rect 1071 1425 1075 1426
rect 1103 1430 1107 1431
rect 1103 1424 1107 1426
rect 1119 1430 1123 1431
rect 1146 1427 1147 1431
rect 1151 1427 1152 1431
rect 1146 1426 1152 1427
rect 1159 1430 1163 1431
rect 1119 1425 1123 1426
rect 1159 1425 1163 1426
rect 1167 1430 1171 1431
rect 1167 1424 1171 1426
rect 1207 1430 1211 1431
rect 1207 1425 1211 1426
rect 1231 1430 1235 1431
rect 1231 1424 1235 1426
rect 1263 1430 1267 1431
rect 1263 1425 1267 1426
rect 1295 1430 1299 1431
rect 1295 1424 1299 1426
rect 1327 1430 1331 1431
rect 1327 1425 1331 1426
rect 1359 1430 1363 1431
rect 1359 1424 1363 1426
rect 1399 1430 1403 1431
rect 1399 1425 1403 1426
rect 1415 1430 1419 1431
rect 1415 1424 1419 1426
rect 1463 1430 1467 1431
rect 1463 1424 1467 1426
rect 1479 1430 1483 1431
rect 1479 1425 1483 1426
rect 1503 1430 1507 1431
rect 1522 1430 1528 1431
rect 1551 1430 1555 1431
rect 1503 1424 1507 1426
rect 902 1423 908 1424
rect 902 1419 903 1423
rect 907 1419 908 1423
rect 902 1418 908 1419
rect 966 1423 972 1424
rect 966 1419 967 1423
rect 971 1419 972 1423
rect 966 1418 972 1419
rect 1030 1423 1036 1424
rect 1030 1419 1031 1423
rect 1035 1419 1036 1423
rect 1030 1418 1036 1419
rect 1102 1423 1108 1424
rect 1102 1419 1103 1423
rect 1107 1419 1108 1423
rect 1102 1418 1108 1419
rect 1166 1423 1172 1424
rect 1166 1419 1167 1423
rect 1171 1419 1172 1423
rect 1166 1418 1172 1419
rect 1230 1423 1236 1424
rect 1230 1419 1231 1423
rect 1235 1419 1236 1423
rect 1230 1418 1236 1419
rect 1294 1423 1300 1424
rect 1294 1419 1295 1423
rect 1299 1419 1300 1423
rect 1294 1418 1300 1419
rect 1358 1423 1364 1424
rect 1358 1419 1359 1423
rect 1363 1419 1364 1423
rect 1358 1418 1364 1419
rect 1414 1423 1420 1424
rect 1414 1419 1415 1423
rect 1419 1419 1420 1423
rect 1414 1418 1420 1419
rect 1462 1423 1468 1424
rect 1462 1419 1463 1423
rect 1467 1419 1468 1423
rect 1462 1418 1468 1419
rect 1502 1423 1508 1424
rect 1502 1419 1503 1423
rect 1507 1419 1508 1423
rect 1502 1418 1508 1419
rect 902 1406 908 1407
rect 902 1402 903 1406
rect 907 1402 908 1406
rect 902 1401 908 1402
rect 966 1406 972 1407
rect 966 1402 967 1406
rect 971 1402 972 1406
rect 966 1401 972 1402
rect 1030 1406 1036 1407
rect 1030 1402 1031 1406
rect 1035 1402 1036 1406
rect 1030 1401 1036 1402
rect 1102 1406 1108 1407
rect 1102 1402 1103 1406
rect 1107 1402 1108 1406
rect 1102 1401 1108 1402
rect 1166 1406 1172 1407
rect 1166 1402 1167 1406
rect 1171 1402 1172 1406
rect 1166 1401 1172 1402
rect 1230 1406 1236 1407
rect 1230 1402 1231 1406
rect 1235 1402 1236 1406
rect 1230 1401 1236 1402
rect 1294 1406 1300 1407
rect 1294 1402 1295 1406
rect 1299 1402 1300 1406
rect 1294 1401 1300 1402
rect 1358 1406 1364 1407
rect 1358 1402 1359 1406
rect 1363 1402 1364 1406
rect 1358 1401 1364 1402
rect 1414 1406 1420 1407
rect 1414 1402 1415 1406
rect 1419 1402 1420 1406
rect 1414 1401 1420 1402
rect 1462 1406 1468 1407
rect 1462 1402 1463 1406
rect 1467 1402 1468 1406
rect 1462 1401 1468 1402
rect 1502 1406 1508 1407
rect 1502 1402 1503 1406
rect 1507 1402 1508 1406
rect 1502 1401 1508 1402
rect 894 1399 900 1400
rect 894 1395 895 1399
rect 899 1395 900 1399
rect 894 1394 900 1395
rect 904 1391 906 1401
rect 968 1391 970 1401
rect 1032 1391 1034 1401
rect 1104 1391 1106 1401
rect 1168 1391 1170 1401
rect 1232 1391 1234 1401
rect 1254 1391 1260 1392
rect 1296 1391 1298 1401
rect 1360 1391 1362 1401
rect 1416 1391 1418 1401
rect 1464 1391 1466 1401
rect 1504 1391 1506 1401
rect 1524 1400 1526 1430
rect 1551 1424 1555 1426
rect 1559 1430 1563 1431
rect 1559 1425 1563 1426
rect 1550 1423 1556 1424
rect 1550 1419 1551 1423
rect 1555 1419 1556 1423
rect 1550 1418 1556 1419
rect 1572 1416 1574 1458
rect 1622 1454 1623 1458
rect 1627 1454 1628 1458
rect 1662 1456 1663 1460
rect 1667 1456 1668 1460
rect 1662 1455 1668 1456
rect 1622 1453 1628 1454
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1662 1443 1668 1444
rect 1622 1441 1628 1442
rect 1622 1437 1623 1441
rect 1627 1437 1628 1441
rect 1622 1436 1628 1437
rect 1624 1431 1626 1436
rect 1591 1430 1595 1431
rect 1591 1424 1595 1426
rect 1623 1430 1627 1431
rect 1623 1424 1627 1426
rect 1590 1423 1596 1424
rect 1590 1419 1591 1423
rect 1595 1419 1596 1423
rect 1590 1418 1596 1419
rect 1622 1423 1628 1424
rect 1622 1419 1623 1423
rect 1627 1419 1628 1423
rect 1622 1418 1628 1419
rect 1570 1415 1576 1416
rect 1570 1411 1571 1415
rect 1575 1411 1576 1415
rect 1570 1410 1576 1411
rect 1550 1406 1556 1407
rect 1550 1402 1551 1406
rect 1555 1402 1556 1406
rect 1550 1401 1556 1402
rect 1590 1406 1596 1407
rect 1590 1402 1591 1406
rect 1595 1402 1596 1406
rect 1590 1401 1596 1402
rect 1622 1406 1628 1407
rect 1622 1402 1623 1406
rect 1627 1402 1628 1406
rect 1622 1401 1628 1402
rect 1522 1399 1528 1400
rect 1522 1395 1523 1399
rect 1527 1395 1528 1399
rect 1522 1394 1528 1395
rect 1552 1391 1554 1401
rect 1592 1391 1594 1401
rect 1624 1391 1626 1401
rect 1640 1400 1642 1442
rect 1662 1439 1663 1443
rect 1667 1439 1668 1443
rect 1662 1438 1668 1439
rect 1664 1431 1666 1438
rect 1663 1430 1667 1431
rect 1663 1425 1667 1426
rect 1664 1422 1666 1425
rect 1662 1421 1668 1422
rect 1662 1417 1663 1421
rect 1667 1417 1668 1421
rect 1662 1416 1668 1417
rect 1662 1404 1668 1405
rect 1662 1400 1663 1404
rect 1667 1400 1668 1404
rect 1630 1399 1636 1400
rect 1630 1395 1631 1399
rect 1635 1395 1636 1399
rect 1630 1394 1636 1395
rect 1638 1399 1644 1400
rect 1662 1399 1668 1400
rect 1638 1395 1639 1399
rect 1643 1395 1644 1399
rect 1638 1394 1644 1395
rect 759 1390 763 1391
rect 770 1387 771 1391
rect 775 1387 776 1391
rect 770 1386 776 1387
rect 815 1390 819 1391
rect 759 1385 763 1386
rect 815 1385 819 1386
rect 831 1390 835 1391
rect 831 1385 835 1386
rect 887 1390 891 1391
rect 887 1385 891 1386
rect 903 1390 907 1391
rect 903 1385 907 1386
rect 959 1390 963 1391
rect 959 1385 963 1386
rect 967 1390 971 1391
rect 967 1385 971 1386
rect 1031 1390 1035 1391
rect 1031 1385 1035 1386
rect 1103 1390 1107 1391
rect 1103 1385 1107 1386
rect 1167 1390 1171 1391
rect 1167 1385 1171 1386
rect 1175 1390 1179 1391
rect 1175 1385 1179 1386
rect 1231 1390 1235 1391
rect 1231 1385 1235 1386
rect 1239 1390 1243 1391
rect 1254 1387 1255 1391
rect 1259 1387 1260 1391
rect 1254 1386 1260 1387
rect 1295 1390 1299 1391
rect 1239 1385 1243 1386
rect 750 1379 756 1380
rect 750 1375 751 1379
rect 755 1375 756 1379
rect 816 1375 818 1385
rect 888 1375 890 1385
rect 902 1379 908 1380
rect 902 1375 903 1379
rect 907 1375 908 1379
rect 960 1375 962 1385
rect 1032 1375 1034 1385
rect 1104 1375 1106 1385
rect 1176 1375 1178 1385
rect 1240 1375 1242 1385
rect 286 1374 292 1375
rect 286 1370 287 1374
rect 291 1370 292 1374
rect 286 1369 292 1370
rect 358 1374 364 1375
rect 358 1370 359 1374
rect 363 1370 364 1374
rect 358 1369 364 1370
rect 430 1374 436 1375
rect 438 1374 444 1375
rect 502 1374 508 1375
rect 518 1374 524 1375
rect 582 1374 588 1375
rect 430 1370 431 1374
rect 435 1370 436 1374
rect 430 1369 436 1370
rect 198 1363 204 1364
rect 110 1359 116 1360
rect 110 1355 111 1359
rect 115 1355 116 1359
rect 198 1359 199 1363
rect 203 1359 204 1363
rect 198 1358 204 1359
rect 242 1363 248 1364
rect 242 1359 243 1363
rect 247 1359 248 1363
rect 242 1358 248 1359
rect 110 1354 116 1355
rect 134 1357 140 1358
rect 112 1351 114 1354
rect 134 1353 135 1357
rect 139 1353 140 1357
rect 134 1352 140 1353
rect 166 1357 172 1358
rect 166 1353 167 1357
rect 171 1353 172 1357
rect 166 1352 172 1353
rect 111 1350 115 1351
rect 111 1345 115 1346
rect 135 1350 139 1352
rect 112 1342 114 1345
rect 135 1344 139 1346
rect 167 1350 171 1352
rect 167 1345 171 1346
rect 183 1350 187 1351
rect 183 1344 187 1346
rect 134 1343 140 1344
rect 110 1341 116 1342
rect 110 1337 111 1341
rect 115 1337 116 1341
rect 134 1339 135 1343
rect 139 1339 140 1343
rect 134 1338 140 1339
rect 182 1343 188 1344
rect 182 1339 183 1343
rect 187 1339 188 1343
rect 182 1338 188 1339
rect 110 1336 116 1337
rect 150 1335 156 1336
rect 150 1331 151 1335
rect 155 1331 156 1335
rect 150 1330 156 1331
rect 134 1326 140 1327
rect 110 1324 116 1325
rect 110 1320 111 1324
rect 115 1320 116 1324
rect 134 1322 135 1326
rect 139 1322 140 1326
rect 134 1321 140 1322
rect 110 1319 116 1320
rect 112 1307 114 1319
rect 136 1307 138 1321
rect 111 1306 115 1307
rect 111 1301 115 1302
rect 135 1306 139 1307
rect 135 1301 139 1302
rect 112 1293 114 1301
rect 110 1292 116 1293
rect 110 1288 111 1292
rect 115 1288 116 1292
rect 136 1291 138 1301
rect 152 1296 154 1330
rect 182 1326 188 1327
rect 182 1322 183 1326
rect 187 1322 188 1326
rect 182 1321 188 1322
rect 184 1307 186 1321
rect 200 1320 202 1358
rect 222 1357 228 1358
rect 222 1353 223 1357
rect 227 1353 228 1357
rect 222 1352 228 1353
rect 286 1357 292 1358
rect 286 1353 287 1357
rect 291 1353 292 1357
rect 286 1352 292 1353
rect 358 1357 364 1358
rect 358 1353 359 1357
rect 363 1353 364 1357
rect 358 1352 364 1353
rect 430 1357 436 1358
rect 430 1353 431 1357
rect 435 1353 436 1357
rect 430 1352 436 1353
rect 223 1350 227 1352
rect 223 1345 227 1346
rect 239 1350 243 1351
rect 239 1344 243 1346
rect 287 1350 291 1352
rect 287 1345 291 1346
rect 295 1350 299 1351
rect 295 1344 299 1346
rect 351 1350 355 1351
rect 351 1344 355 1346
rect 359 1350 363 1352
rect 359 1345 363 1346
rect 399 1350 403 1351
rect 399 1344 403 1346
rect 431 1350 435 1352
rect 431 1345 435 1346
rect 238 1343 244 1344
rect 238 1339 239 1343
rect 243 1339 244 1343
rect 238 1338 244 1339
rect 294 1343 300 1344
rect 294 1339 295 1343
rect 299 1339 300 1343
rect 294 1338 300 1339
rect 350 1343 356 1344
rect 350 1339 351 1343
rect 355 1339 356 1343
rect 350 1338 356 1339
rect 398 1343 404 1344
rect 398 1339 399 1343
rect 403 1339 404 1343
rect 398 1338 404 1339
rect 440 1336 442 1374
rect 502 1370 503 1374
rect 507 1370 508 1374
rect 502 1369 508 1370
rect 502 1357 508 1358
rect 502 1353 503 1357
rect 507 1353 508 1357
rect 502 1352 508 1353
rect 520 1352 522 1374
rect 582 1370 583 1374
rect 587 1370 588 1374
rect 582 1369 588 1370
rect 662 1374 668 1375
rect 662 1370 663 1374
rect 667 1370 668 1374
rect 662 1369 668 1370
rect 742 1374 748 1375
rect 750 1374 756 1375
rect 814 1374 820 1375
rect 742 1370 743 1374
rect 747 1370 748 1374
rect 742 1369 748 1370
rect 814 1370 815 1374
rect 819 1370 820 1374
rect 814 1369 820 1370
rect 886 1374 892 1375
rect 902 1374 908 1375
rect 958 1374 964 1375
rect 886 1370 887 1374
rect 891 1370 892 1374
rect 886 1369 892 1370
rect 710 1363 716 1364
rect 710 1359 711 1363
rect 715 1359 716 1363
rect 710 1358 716 1359
rect 582 1357 588 1358
rect 582 1353 583 1357
rect 587 1353 588 1357
rect 582 1352 588 1353
rect 662 1357 668 1358
rect 662 1353 663 1357
rect 667 1353 668 1357
rect 662 1352 668 1353
rect 455 1350 459 1351
rect 455 1344 459 1346
rect 503 1350 507 1352
rect 518 1351 524 1352
rect 503 1345 507 1346
rect 511 1350 515 1351
rect 518 1347 519 1351
rect 523 1347 524 1351
rect 518 1346 524 1347
rect 567 1350 571 1351
rect 511 1344 515 1346
rect 567 1344 571 1346
rect 583 1350 587 1352
rect 583 1345 587 1346
rect 631 1350 635 1351
rect 631 1344 635 1346
rect 663 1350 667 1352
rect 663 1345 667 1346
rect 695 1350 699 1351
rect 695 1344 699 1346
rect 454 1343 460 1344
rect 454 1339 455 1343
rect 459 1339 460 1343
rect 454 1338 460 1339
rect 510 1343 516 1344
rect 510 1339 511 1343
rect 515 1339 516 1343
rect 510 1338 516 1339
rect 566 1343 572 1344
rect 566 1339 567 1343
rect 571 1339 572 1343
rect 566 1338 572 1339
rect 630 1343 636 1344
rect 630 1339 631 1343
rect 635 1339 636 1343
rect 630 1338 636 1339
rect 694 1343 700 1344
rect 694 1339 695 1343
rect 699 1339 700 1343
rect 694 1338 700 1339
rect 438 1335 444 1336
rect 438 1331 439 1335
rect 443 1331 444 1335
rect 438 1330 444 1331
rect 622 1335 628 1336
rect 622 1331 623 1335
rect 627 1331 628 1335
rect 622 1330 628 1331
rect 642 1335 648 1336
rect 642 1331 643 1335
rect 647 1331 648 1335
rect 642 1330 648 1331
rect 238 1326 244 1327
rect 238 1322 239 1326
rect 243 1322 244 1326
rect 238 1321 244 1322
rect 294 1326 300 1327
rect 294 1322 295 1326
rect 299 1322 300 1326
rect 294 1321 300 1322
rect 350 1326 356 1327
rect 350 1322 351 1326
rect 355 1322 356 1326
rect 350 1321 356 1322
rect 398 1326 404 1327
rect 398 1322 399 1326
rect 403 1322 404 1326
rect 398 1321 404 1322
rect 454 1326 460 1327
rect 454 1322 455 1326
rect 459 1322 460 1326
rect 454 1321 460 1322
rect 510 1326 516 1327
rect 510 1322 511 1326
rect 515 1322 516 1326
rect 510 1321 516 1322
rect 566 1326 572 1327
rect 566 1322 567 1326
rect 571 1322 572 1326
rect 566 1321 572 1322
rect 198 1319 204 1320
rect 198 1315 199 1319
rect 203 1315 204 1319
rect 198 1314 204 1315
rect 240 1307 242 1321
rect 296 1307 298 1321
rect 352 1307 354 1321
rect 390 1311 396 1312
rect 390 1307 391 1311
rect 395 1307 396 1311
rect 400 1307 402 1321
rect 456 1307 458 1321
rect 512 1307 514 1321
rect 568 1307 570 1321
rect 183 1306 187 1307
rect 183 1301 187 1302
rect 231 1306 235 1307
rect 231 1301 235 1302
rect 239 1306 243 1307
rect 239 1301 243 1302
rect 279 1306 283 1307
rect 279 1301 283 1302
rect 295 1306 299 1307
rect 295 1301 299 1302
rect 327 1306 331 1307
rect 327 1301 331 1302
rect 351 1306 355 1307
rect 351 1301 355 1302
rect 375 1306 379 1307
rect 390 1306 396 1307
rect 399 1306 403 1307
rect 375 1301 379 1302
rect 150 1295 156 1296
rect 150 1291 151 1295
rect 155 1291 156 1295
rect 184 1291 186 1301
rect 232 1291 234 1301
rect 280 1291 282 1301
rect 294 1295 300 1296
rect 294 1291 295 1295
rect 299 1291 300 1295
rect 328 1291 330 1301
rect 376 1291 378 1301
rect 110 1287 116 1288
rect 134 1290 140 1291
rect 150 1290 156 1291
rect 182 1290 188 1291
rect 134 1286 135 1290
rect 139 1286 140 1290
rect 134 1285 140 1286
rect 182 1286 183 1290
rect 187 1286 188 1290
rect 182 1285 188 1286
rect 230 1290 236 1291
rect 230 1286 231 1290
rect 235 1286 236 1290
rect 230 1285 236 1286
rect 278 1290 284 1291
rect 294 1290 300 1291
rect 326 1290 332 1291
rect 278 1286 279 1290
rect 283 1286 284 1290
rect 278 1285 284 1286
rect 242 1279 248 1280
rect 110 1275 116 1276
rect 110 1271 111 1275
rect 115 1271 116 1275
rect 242 1275 243 1279
rect 247 1275 248 1279
rect 242 1274 248 1275
rect 110 1270 116 1271
rect 134 1273 140 1274
rect 112 1267 114 1270
rect 134 1269 135 1273
rect 139 1269 140 1273
rect 134 1268 140 1269
rect 182 1273 188 1274
rect 182 1269 183 1273
rect 187 1269 188 1273
rect 182 1268 188 1269
rect 230 1273 236 1274
rect 230 1269 231 1273
rect 235 1269 236 1273
rect 230 1268 236 1269
rect 111 1266 115 1267
rect 111 1261 115 1262
rect 135 1266 139 1268
rect 112 1258 114 1261
rect 135 1260 139 1262
rect 167 1266 171 1267
rect 167 1260 171 1262
rect 183 1266 187 1268
rect 183 1261 187 1262
rect 223 1266 227 1267
rect 223 1260 227 1262
rect 231 1266 235 1268
rect 231 1261 235 1262
rect 134 1259 140 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 134 1255 135 1259
rect 139 1255 140 1259
rect 134 1254 140 1255
rect 166 1259 172 1260
rect 166 1255 167 1259
rect 171 1255 172 1259
rect 166 1254 172 1255
rect 222 1259 228 1260
rect 222 1255 223 1259
rect 227 1255 228 1259
rect 222 1254 228 1255
rect 110 1252 116 1253
rect 150 1251 156 1252
rect 150 1247 151 1251
rect 155 1247 156 1251
rect 150 1246 156 1247
rect 134 1242 140 1243
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 134 1238 135 1242
rect 139 1238 140 1242
rect 134 1237 140 1238
rect 110 1235 116 1236
rect 112 1223 114 1235
rect 136 1223 138 1237
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 135 1222 139 1223
rect 135 1217 139 1218
rect 112 1209 114 1217
rect 110 1208 116 1209
rect 110 1204 111 1208
rect 115 1204 116 1208
rect 136 1207 138 1217
rect 152 1212 154 1246
rect 166 1242 172 1243
rect 166 1238 167 1242
rect 171 1238 172 1242
rect 166 1237 172 1238
rect 222 1242 228 1243
rect 222 1238 223 1242
rect 227 1238 228 1242
rect 222 1237 228 1238
rect 168 1223 170 1237
rect 224 1223 226 1237
rect 244 1236 246 1274
rect 278 1273 284 1274
rect 278 1269 279 1273
rect 283 1269 284 1273
rect 278 1268 284 1269
rect 279 1266 283 1268
rect 279 1260 283 1262
rect 278 1259 284 1260
rect 278 1255 279 1259
rect 283 1255 284 1259
rect 278 1254 284 1255
rect 296 1252 298 1290
rect 326 1286 327 1290
rect 331 1286 332 1290
rect 326 1285 332 1286
rect 374 1290 380 1291
rect 374 1286 375 1290
rect 379 1286 380 1290
rect 374 1285 380 1286
rect 392 1280 394 1306
rect 399 1301 403 1302
rect 431 1306 435 1307
rect 431 1301 435 1302
rect 455 1306 459 1307
rect 455 1301 459 1302
rect 487 1306 491 1307
rect 487 1301 491 1302
rect 511 1306 515 1307
rect 511 1301 515 1302
rect 543 1306 547 1307
rect 543 1301 547 1302
rect 567 1306 571 1307
rect 567 1301 571 1302
rect 607 1306 611 1307
rect 607 1301 611 1302
rect 432 1291 434 1301
rect 488 1291 490 1301
rect 544 1291 546 1301
rect 598 1295 604 1296
rect 598 1291 599 1295
rect 603 1291 604 1295
rect 608 1291 610 1301
rect 624 1296 626 1330
rect 630 1326 636 1327
rect 630 1322 631 1326
rect 635 1322 636 1326
rect 630 1321 636 1322
rect 632 1307 634 1321
rect 644 1312 646 1330
rect 694 1326 700 1327
rect 694 1322 695 1326
rect 699 1322 700 1326
rect 694 1321 700 1322
rect 642 1311 648 1312
rect 642 1307 643 1311
rect 647 1307 648 1311
rect 696 1307 698 1321
rect 712 1320 714 1358
rect 742 1357 748 1358
rect 742 1353 743 1357
rect 747 1353 748 1357
rect 742 1352 748 1353
rect 814 1357 820 1358
rect 814 1353 815 1357
rect 819 1353 820 1357
rect 814 1352 820 1353
rect 886 1357 892 1358
rect 886 1353 887 1357
rect 891 1353 892 1357
rect 886 1352 892 1353
rect 904 1352 906 1374
rect 958 1370 959 1374
rect 963 1370 964 1374
rect 958 1369 964 1370
rect 1030 1374 1036 1375
rect 1030 1370 1031 1374
rect 1035 1370 1036 1374
rect 1030 1369 1036 1370
rect 1102 1374 1108 1375
rect 1102 1370 1103 1374
rect 1107 1370 1108 1374
rect 1102 1369 1108 1370
rect 1174 1374 1180 1375
rect 1174 1370 1175 1374
rect 1179 1370 1180 1374
rect 1174 1369 1180 1370
rect 1238 1374 1244 1375
rect 1238 1370 1239 1374
rect 1243 1370 1244 1374
rect 1238 1369 1244 1370
rect 1256 1364 1258 1386
rect 1295 1385 1299 1386
rect 1303 1390 1307 1391
rect 1303 1385 1307 1386
rect 1359 1390 1363 1391
rect 1359 1385 1363 1386
rect 1367 1390 1371 1391
rect 1367 1385 1371 1386
rect 1415 1390 1419 1391
rect 1415 1385 1419 1386
rect 1431 1390 1435 1391
rect 1431 1385 1435 1386
rect 1463 1390 1467 1391
rect 1463 1385 1467 1386
rect 1495 1390 1499 1391
rect 1495 1385 1499 1386
rect 1503 1390 1507 1391
rect 1503 1385 1507 1386
rect 1551 1390 1555 1391
rect 1551 1385 1555 1386
rect 1567 1390 1571 1391
rect 1567 1385 1571 1386
rect 1591 1390 1595 1391
rect 1591 1385 1595 1386
rect 1623 1390 1627 1391
rect 1623 1385 1627 1386
rect 1304 1375 1306 1385
rect 1318 1379 1324 1380
rect 1318 1375 1319 1379
rect 1323 1375 1324 1379
rect 1368 1375 1370 1385
rect 1432 1375 1434 1385
rect 1496 1375 1498 1385
rect 1568 1375 1570 1385
rect 1624 1375 1626 1385
rect 1302 1374 1308 1375
rect 1318 1374 1324 1375
rect 1366 1374 1372 1375
rect 1302 1370 1303 1374
rect 1307 1370 1308 1374
rect 1302 1369 1308 1370
rect 1254 1363 1260 1364
rect 1254 1359 1255 1363
rect 1259 1359 1260 1363
rect 1254 1358 1260 1359
rect 958 1357 964 1358
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 1030 1357 1036 1358
rect 1030 1353 1031 1357
rect 1035 1353 1036 1357
rect 1030 1352 1036 1353
rect 1102 1357 1108 1358
rect 1102 1353 1103 1357
rect 1107 1353 1108 1357
rect 1102 1352 1108 1353
rect 1174 1357 1180 1358
rect 1174 1353 1175 1357
rect 1179 1353 1180 1357
rect 1174 1352 1180 1353
rect 1238 1357 1244 1358
rect 1238 1353 1239 1357
rect 1243 1353 1244 1357
rect 1238 1352 1244 1353
rect 1302 1357 1308 1358
rect 1302 1353 1303 1357
rect 1307 1353 1308 1357
rect 1302 1352 1308 1353
rect 1320 1352 1322 1374
rect 1366 1370 1367 1374
rect 1371 1370 1372 1374
rect 1366 1369 1372 1370
rect 1430 1374 1436 1375
rect 1430 1370 1431 1374
rect 1435 1370 1436 1374
rect 1430 1369 1436 1370
rect 1494 1374 1500 1375
rect 1494 1370 1495 1374
rect 1499 1370 1500 1374
rect 1494 1369 1500 1370
rect 1566 1374 1572 1375
rect 1566 1370 1567 1374
rect 1571 1370 1572 1374
rect 1566 1369 1572 1370
rect 1622 1374 1628 1375
rect 1622 1370 1623 1374
rect 1627 1370 1628 1374
rect 1622 1369 1628 1370
rect 1632 1364 1634 1394
rect 1664 1391 1666 1399
rect 1663 1390 1667 1391
rect 1663 1385 1667 1386
rect 1642 1379 1648 1380
rect 1642 1375 1643 1379
rect 1647 1375 1648 1379
rect 1664 1377 1666 1385
rect 1642 1374 1648 1375
rect 1662 1376 1668 1377
rect 1486 1363 1492 1364
rect 1486 1359 1487 1363
rect 1491 1359 1492 1363
rect 1632 1363 1640 1364
rect 1632 1361 1635 1363
rect 1486 1358 1492 1359
rect 1634 1359 1635 1361
rect 1639 1359 1640 1363
rect 1634 1358 1640 1359
rect 1366 1357 1372 1358
rect 1366 1353 1367 1357
rect 1371 1353 1372 1357
rect 1366 1352 1372 1353
rect 1430 1357 1436 1358
rect 1430 1353 1431 1357
rect 1435 1353 1436 1357
rect 1430 1352 1436 1353
rect 743 1350 747 1352
rect 743 1345 747 1346
rect 759 1350 763 1351
rect 759 1344 763 1346
rect 815 1350 819 1352
rect 815 1345 819 1346
rect 823 1350 827 1351
rect 823 1344 827 1346
rect 887 1350 891 1352
rect 902 1351 908 1352
rect 902 1347 903 1351
rect 907 1347 908 1351
rect 902 1346 908 1347
rect 959 1350 963 1352
rect 887 1344 891 1346
rect 959 1344 963 1346
rect 1023 1350 1027 1351
rect 1023 1344 1027 1346
rect 1031 1350 1035 1352
rect 1031 1345 1035 1346
rect 1087 1350 1091 1351
rect 1087 1344 1091 1346
rect 1103 1350 1107 1352
rect 1103 1345 1107 1346
rect 1151 1350 1155 1351
rect 1151 1344 1155 1346
rect 1175 1350 1179 1352
rect 1175 1345 1179 1346
rect 1215 1350 1219 1351
rect 1215 1344 1219 1346
rect 1239 1350 1243 1352
rect 1239 1345 1243 1346
rect 1279 1350 1283 1351
rect 1279 1344 1283 1346
rect 1303 1350 1307 1352
rect 1318 1351 1324 1352
rect 1318 1347 1319 1351
rect 1323 1347 1324 1351
rect 1318 1346 1324 1347
rect 1343 1350 1347 1351
rect 1303 1345 1307 1346
rect 1343 1344 1347 1346
rect 1367 1350 1371 1352
rect 1367 1345 1371 1346
rect 1407 1350 1411 1351
rect 1407 1344 1411 1346
rect 1431 1350 1435 1352
rect 1431 1345 1435 1346
rect 1479 1350 1483 1351
rect 1479 1344 1483 1346
rect 758 1343 764 1344
rect 758 1339 759 1343
rect 763 1339 764 1343
rect 758 1338 764 1339
rect 822 1343 828 1344
rect 822 1339 823 1343
rect 827 1339 828 1343
rect 822 1338 828 1339
rect 886 1343 892 1344
rect 886 1339 887 1343
rect 891 1339 892 1343
rect 886 1338 892 1339
rect 958 1343 964 1344
rect 958 1339 959 1343
rect 963 1339 964 1343
rect 958 1338 964 1339
rect 1022 1343 1028 1344
rect 1022 1339 1023 1343
rect 1027 1339 1028 1343
rect 1022 1338 1028 1339
rect 1086 1343 1092 1344
rect 1086 1339 1087 1343
rect 1091 1339 1092 1343
rect 1086 1338 1092 1339
rect 1150 1343 1156 1344
rect 1150 1339 1151 1343
rect 1155 1339 1156 1343
rect 1150 1338 1156 1339
rect 1214 1343 1220 1344
rect 1214 1339 1215 1343
rect 1219 1339 1220 1343
rect 1214 1338 1220 1339
rect 1278 1343 1284 1344
rect 1278 1339 1279 1343
rect 1283 1339 1284 1343
rect 1278 1338 1284 1339
rect 1342 1343 1348 1344
rect 1342 1339 1343 1343
rect 1347 1339 1348 1343
rect 1342 1338 1348 1339
rect 1406 1343 1412 1344
rect 1406 1339 1407 1343
rect 1411 1339 1412 1343
rect 1406 1338 1412 1339
rect 1478 1343 1484 1344
rect 1478 1339 1479 1343
rect 1483 1339 1484 1343
rect 1478 1338 1484 1339
rect 738 1335 744 1336
rect 738 1331 739 1335
rect 743 1331 744 1335
rect 738 1330 744 1331
rect 1374 1335 1380 1336
rect 1374 1331 1375 1335
rect 1379 1331 1380 1335
rect 1374 1330 1380 1331
rect 1382 1335 1388 1336
rect 1382 1331 1383 1335
rect 1387 1331 1388 1335
rect 1382 1330 1388 1331
rect 740 1320 742 1330
rect 758 1326 764 1327
rect 758 1322 759 1326
rect 763 1322 764 1326
rect 758 1321 764 1322
rect 822 1326 828 1327
rect 822 1322 823 1326
rect 827 1322 828 1326
rect 822 1321 828 1322
rect 886 1326 892 1327
rect 886 1322 887 1326
rect 891 1322 892 1326
rect 886 1321 892 1322
rect 958 1326 964 1327
rect 958 1322 959 1326
rect 963 1322 964 1326
rect 958 1321 964 1322
rect 1022 1326 1028 1327
rect 1022 1322 1023 1326
rect 1027 1322 1028 1326
rect 1022 1321 1028 1322
rect 1086 1326 1092 1327
rect 1086 1322 1087 1326
rect 1091 1322 1092 1326
rect 1086 1321 1092 1322
rect 1150 1326 1156 1327
rect 1150 1322 1151 1326
rect 1155 1322 1156 1326
rect 1150 1321 1156 1322
rect 1214 1326 1220 1327
rect 1214 1322 1215 1326
rect 1219 1322 1220 1326
rect 1214 1321 1220 1322
rect 1278 1326 1284 1327
rect 1278 1322 1279 1326
rect 1283 1322 1284 1326
rect 1278 1321 1284 1322
rect 1342 1326 1348 1327
rect 1342 1322 1343 1326
rect 1347 1322 1348 1326
rect 1342 1321 1348 1322
rect 710 1319 716 1320
rect 710 1315 711 1319
rect 715 1315 716 1319
rect 710 1314 716 1315
rect 738 1319 744 1320
rect 738 1315 739 1319
rect 743 1315 744 1319
rect 738 1314 744 1315
rect 760 1307 762 1321
rect 824 1307 826 1321
rect 888 1307 890 1321
rect 960 1307 962 1321
rect 1024 1307 1026 1321
rect 1088 1307 1090 1321
rect 1094 1311 1100 1312
rect 1094 1307 1095 1311
rect 1099 1307 1100 1311
rect 1152 1307 1154 1321
rect 1216 1307 1218 1321
rect 1280 1307 1282 1321
rect 1344 1307 1346 1321
rect 631 1306 635 1307
rect 642 1306 648 1307
rect 663 1306 667 1307
rect 631 1301 635 1302
rect 663 1301 667 1302
rect 695 1306 699 1307
rect 695 1301 699 1302
rect 719 1306 723 1307
rect 719 1301 723 1302
rect 759 1306 763 1307
rect 759 1301 763 1302
rect 775 1306 779 1307
rect 775 1301 779 1302
rect 823 1306 827 1307
rect 823 1301 827 1302
rect 831 1306 835 1307
rect 831 1301 835 1302
rect 887 1306 891 1307
rect 887 1301 891 1302
rect 895 1306 899 1307
rect 895 1301 899 1302
rect 959 1306 963 1307
rect 959 1301 963 1302
rect 1023 1306 1027 1307
rect 1023 1301 1027 1302
rect 1079 1306 1083 1307
rect 1079 1301 1083 1302
rect 1087 1306 1091 1307
rect 1094 1306 1100 1307
rect 1143 1306 1147 1307
rect 1087 1301 1091 1302
rect 622 1295 628 1296
rect 622 1291 623 1295
rect 627 1291 628 1295
rect 664 1291 666 1301
rect 720 1291 722 1301
rect 734 1295 740 1296
rect 734 1291 735 1295
rect 739 1291 740 1295
rect 776 1291 778 1301
rect 782 1295 788 1296
rect 782 1291 783 1295
rect 787 1291 788 1295
rect 832 1291 834 1301
rect 896 1291 898 1301
rect 960 1291 962 1301
rect 1024 1291 1026 1301
rect 1080 1291 1082 1301
rect 430 1290 436 1291
rect 430 1286 431 1290
rect 435 1286 436 1290
rect 430 1285 436 1286
rect 486 1290 492 1291
rect 486 1286 487 1290
rect 491 1286 492 1290
rect 486 1285 492 1286
rect 542 1290 548 1291
rect 598 1290 604 1291
rect 606 1290 612 1291
rect 622 1290 628 1291
rect 662 1290 668 1291
rect 542 1286 543 1290
rect 547 1286 548 1290
rect 542 1285 548 1286
rect 390 1279 396 1280
rect 390 1275 391 1279
rect 395 1275 396 1279
rect 390 1274 396 1275
rect 450 1279 456 1280
rect 450 1275 451 1279
rect 455 1275 456 1279
rect 450 1274 456 1275
rect 326 1273 332 1274
rect 326 1269 327 1273
rect 331 1269 332 1273
rect 326 1268 332 1269
rect 374 1273 380 1274
rect 374 1269 375 1273
rect 379 1269 380 1273
rect 374 1268 380 1269
rect 430 1273 436 1274
rect 430 1269 431 1273
rect 435 1269 436 1273
rect 430 1268 436 1269
rect 327 1266 331 1268
rect 327 1260 331 1262
rect 375 1266 379 1268
rect 375 1261 379 1262
rect 383 1266 387 1267
rect 383 1260 387 1262
rect 431 1266 435 1268
rect 431 1261 435 1262
rect 439 1266 443 1267
rect 439 1260 443 1262
rect 326 1259 332 1260
rect 326 1255 327 1259
rect 331 1255 332 1259
rect 326 1254 332 1255
rect 382 1259 388 1260
rect 382 1255 383 1259
rect 387 1255 388 1259
rect 382 1254 388 1255
rect 438 1259 444 1260
rect 438 1255 439 1259
rect 443 1255 444 1259
rect 438 1254 444 1255
rect 294 1251 300 1252
rect 294 1247 295 1251
rect 299 1247 300 1251
rect 294 1246 300 1247
rect 278 1242 284 1243
rect 278 1238 279 1242
rect 283 1238 284 1242
rect 278 1237 284 1238
rect 326 1242 332 1243
rect 326 1238 327 1242
rect 331 1238 332 1242
rect 326 1237 332 1238
rect 382 1242 388 1243
rect 382 1238 383 1242
rect 387 1238 388 1242
rect 382 1237 388 1238
rect 438 1242 444 1243
rect 438 1238 439 1242
rect 443 1238 444 1242
rect 438 1237 444 1238
rect 242 1235 248 1236
rect 242 1231 243 1235
rect 247 1231 248 1235
rect 242 1230 248 1231
rect 280 1223 282 1237
rect 328 1223 330 1237
rect 384 1223 386 1237
rect 398 1235 404 1236
rect 398 1231 399 1235
rect 403 1231 404 1235
rect 398 1230 404 1231
rect 167 1222 171 1223
rect 167 1217 171 1218
rect 223 1222 227 1223
rect 223 1217 227 1218
rect 279 1222 283 1223
rect 279 1217 283 1218
rect 327 1222 331 1223
rect 327 1217 331 1218
rect 335 1222 339 1223
rect 335 1217 339 1218
rect 383 1222 387 1223
rect 383 1217 387 1218
rect 150 1211 156 1212
rect 150 1207 151 1211
rect 155 1207 156 1211
rect 168 1207 170 1217
rect 224 1207 226 1217
rect 280 1207 282 1217
rect 306 1215 312 1216
rect 298 1211 304 1212
rect 298 1207 299 1211
rect 303 1207 304 1211
rect 306 1211 307 1215
rect 311 1211 312 1215
rect 306 1210 312 1211
rect 110 1203 116 1204
rect 134 1206 140 1207
rect 150 1206 156 1207
rect 166 1206 172 1207
rect 134 1202 135 1206
rect 139 1202 140 1206
rect 134 1201 140 1202
rect 166 1202 167 1206
rect 171 1202 172 1206
rect 166 1201 172 1202
rect 222 1206 228 1207
rect 222 1202 223 1206
rect 227 1202 228 1206
rect 222 1201 228 1202
rect 278 1206 284 1207
rect 298 1206 304 1207
rect 278 1202 279 1206
rect 283 1202 284 1206
rect 278 1201 284 1202
rect 238 1195 244 1196
rect 110 1191 116 1192
rect 110 1187 111 1191
rect 115 1187 116 1191
rect 238 1191 239 1195
rect 243 1191 244 1195
rect 238 1190 244 1191
rect 110 1186 116 1187
rect 134 1189 140 1190
rect 112 1179 114 1186
rect 134 1185 135 1189
rect 139 1185 140 1189
rect 134 1184 140 1185
rect 166 1189 172 1190
rect 166 1185 167 1189
rect 171 1185 172 1189
rect 166 1184 172 1185
rect 222 1189 228 1190
rect 222 1185 223 1189
rect 227 1185 228 1189
rect 222 1184 228 1185
rect 136 1179 138 1184
rect 168 1179 170 1184
rect 224 1179 226 1184
rect 111 1178 115 1179
rect 111 1173 115 1174
rect 135 1178 139 1179
rect 112 1170 114 1173
rect 135 1172 139 1174
rect 167 1178 171 1179
rect 167 1172 171 1174
rect 223 1178 227 1179
rect 223 1172 227 1174
rect 134 1171 140 1172
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 134 1167 135 1171
rect 139 1167 140 1171
rect 134 1166 140 1167
rect 166 1171 172 1172
rect 166 1167 167 1171
rect 171 1167 172 1171
rect 166 1166 172 1167
rect 222 1171 228 1172
rect 222 1167 223 1171
rect 227 1167 228 1171
rect 222 1166 228 1167
rect 110 1164 116 1165
rect 154 1163 160 1164
rect 154 1159 155 1163
rect 159 1159 160 1163
rect 154 1158 160 1159
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 134 1150 135 1154
rect 139 1150 140 1154
rect 134 1149 140 1150
rect 110 1147 116 1148
rect 112 1135 114 1147
rect 136 1135 138 1149
rect 111 1134 115 1135
rect 111 1129 115 1130
rect 135 1134 139 1135
rect 135 1129 139 1130
rect 143 1134 147 1135
rect 143 1129 147 1130
rect 112 1121 114 1129
rect 110 1120 116 1121
rect 110 1116 111 1120
rect 115 1116 116 1120
rect 144 1119 146 1129
rect 156 1124 158 1158
rect 166 1154 172 1155
rect 166 1150 167 1154
rect 171 1150 172 1154
rect 166 1149 172 1150
rect 222 1154 228 1155
rect 222 1150 223 1154
rect 227 1150 228 1154
rect 222 1149 228 1150
rect 168 1135 170 1149
rect 224 1135 226 1149
rect 240 1148 242 1190
rect 278 1189 284 1190
rect 278 1185 279 1189
rect 283 1185 284 1189
rect 278 1184 284 1185
rect 280 1179 282 1184
rect 279 1178 283 1179
rect 279 1173 283 1174
rect 287 1178 291 1179
rect 287 1172 291 1174
rect 286 1171 292 1172
rect 286 1167 287 1171
rect 291 1167 292 1171
rect 286 1166 292 1167
rect 300 1164 302 1206
rect 308 1196 310 1210
rect 336 1207 338 1217
rect 384 1207 386 1217
rect 334 1206 340 1207
rect 334 1202 335 1206
rect 339 1202 340 1206
rect 334 1201 340 1202
rect 382 1206 388 1207
rect 382 1202 383 1206
rect 387 1202 388 1206
rect 382 1201 388 1202
rect 400 1196 402 1230
rect 440 1223 442 1237
rect 452 1236 454 1274
rect 486 1273 492 1274
rect 486 1269 487 1273
rect 491 1269 492 1273
rect 486 1268 492 1269
rect 542 1273 548 1274
rect 542 1269 543 1273
rect 547 1269 548 1273
rect 542 1268 548 1269
rect 600 1268 602 1290
rect 606 1286 607 1290
rect 611 1286 612 1290
rect 606 1285 612 1286
rect 662 1286 663 1290
rect 667 1286 668 1290
rect 662 1285 668 1286
rect 718 1290 724 1291
rect 734 1290 740 1291
rect 774 1290 780 1291
rect 782 1290 788 1291
rect 830 1290 836 1291
rect 718 1286 719 1290
rect 723 1286 724 1290
rect 718 1285 724 1286
rect 606 1273 612 1274
rect 606 1269 607 1273
rect 611 1269 612 1273
rect 606 1268 612 1269
rect 662 1273 668 1274
rect 662 1269 663 1273
rect 667 1269 668 1273
rect 662 1268 668 1269
rect 718 1273 724 1274
rect 718 1269 719 1273
rect 723 1269 724 1273
rect 718 1268 724 1269
rect 487 1266 491 1268
rect 487 1261 491 1262
rect 495 1266 499 1267
rect 495 1260 499 1262
rect 543 1266 547 1268
rect 598 1267 604 1268
rect 543 1261 547 1262
rect 551 1266 555 1267
rect 598 1263 599 1267
rect 603 1263 604 1267
rect 598 1262 604 1263
rect 607 1266 611 1268
rect 551 1260 555 1262
rect 607 1260 611 1262
rect 663 1266 667 1268
rect 663 1260 667 1262
rect 719 1266 723 1268
rect 719 1260 723 1262
rect 494 1259 500 1260
rect 494 1255 495 1259
rect 499 1255 500 1259
rect 494 1254 500 1255
rect 550 1259 556 1260
rect 550 1255 551 1259
rect 555 1255 556 1259
rect 550 1254 556 1255
rect 606 1259 612 1260
rect 606 1255 607 1259
rect 611 1255 612 1259
rect 606 1254 612 1255
rect 662 1259 668 1260
rect 662 1255 663 1259
rect 667 1255 668 1259
rect 662 1254 668 1255
rect 718 1259 724 1260
rect 718 1255 719 1259
rect 723 1255 724 1259
rect 718 1254 724 1255
rect 736 1252 738 1290
rect 774 1286 775 1290
rect 779 1286 780 1290
rect 774 1285 780 1286
rect 758 1279 764 1280
rect 758 1275 759 1279
rect 763 1275 764 1279
rect 758 1274 764 1275
rect 618 1251 624 1252
rect 618 1247 619 1251
rect 623 1247 624 1251
rect 618 1246 624 1247
rect 734 1251 740 1252
rect 734 1247 735 1251
rect 739 1247 740 1251
rect 734 1246 740 1247
rect 494 1242 500 1243
rect 494 1238 495 1242
rect 499 1238 500 1242
rect 494 1237 500 1238
rect 550 1242 556 1243
rect 550 1238 551 1242
rect 555 1238 556 1242
rect 550 1237 556 1238
rect 606 1242 612 1243
rect 606 1238 607 1242
rect 611 1238 612 1242
rect 606 1237 612 1238
rect 450 1235 456 1236
rect 450 1231 451 1235
rect 455 1231 456 1235
rect 450 1230 456 1231
rect 496 1223 498 1237
rect 552 1223 554 1237
rect 608 1223 610 1237
rect 620 1224 622 1246
rect 662 1242 668 1243
rect 662 1238 663 1242
rect 667 1238 668 1242
rect 662 1237 668 1238
rect 718 1242 724 1243
rect 718 1238 719 1242
rect 723 1238 724 1242
rect 718 1237 724 1238
rect 618 1223 624 1224
rect 664 1223 666 1237
rect 720 1223 722 1237
rect 760 1236 762 1274
rect 774 1273 780 1274
rect 774 1269 775 1273
rect 779 1269 780 1273
rect 774 1268 780 1269
rect 767 1266 771 1267
rect 767 1260 771 1262
rect 775 1266 779 1268
rect 775 1261 779 1262
rect 766 1259 772 1260
rect 766 1255 767 1259
rect 771 1255 772 1259
rect 766 1254 772 1255
rect 784 1252 786 1290
rect 830 1286 831 1290
rect 835 1286 836 1290
rect 830 1285 836 1286
rect 894 1290 900 1291
rect 894 1286 895 1290
rect 899 1286 900 1290
rect 894 1285 900 1286
rect 958 1290 964 1291
rect 958 1286 959 1290
rect 963 1286 964 1290
rect 958 1285 964 1286
rect 1022 1290 1028 1291
rect 1022 1286 1023 1290
rect 1027 1286 1028 1290
rect 1022 1285 1028 1286
rect 1078 1290 1084 1291
rect 1078 1286 1079 1290
rect 1083 1286 1084 1290
rect 1078 1285 1084 1286
rect 1096 1280 1098 1306
rect 1143 1301 1147 1302
rect 1151 1306 1155 1307
rect 1151 1301 1155 1302
rect 1207 1306 1211 1307
rect 1207 1301 1211 1302
rect 1215 1306 1219 1307
rect 1215 1301 1219 1302
rect 1279 1306 1283 1307
rect 1279 1301 1283 1302
rect 1343 1306 1347 1307
rect 1343 1301 1347 1302
rect 1359 1306 1363 1307
rect 1359 1301 1363 1302
rect 1144 1291 1146 1301
rect 1208 1291 1210 1301
rect 1280 1291 1282 1301
rect 1350 1295 1356 1296
rect 1350 1291 1351 1295
rect 1355 1291 1356 1295
rect 1360 1291 1362 1301
rect 1376 1296 1378 1330
rect 1384 1312 1386 1330
rect 1406 1326 1412 1327
rect 1406 1322 1407 1326
rect 1411 1322 1412 1326
rect 1406 1321 1412 1322
rect 1478 1326 1484 1327
rect 1478 1322 1479 1326
rect 1483 1322 1484 1326
rect 1478 1321 1484 1322
rect 1382 1311 1388 1312
rect 1382 1307 1383 1311
rect 1387 1307 1388 1311
rect 1408 1307 1410 1321
rect 1480 1307 1482 1321
rect 1488 1320 1490 1358
rect 1494 1357 1500 1358
rect 1494 1353 1495 1357
rect 1499 1353 1500 1357
rect 1494 1352 1500 1353
rect 1566 1357 1572 1358
rect 1566 1353 1567 1357
rect 1571 1353 1572 1357
rect 1566 1352 1572 1353
rect 1622 1357 1628 1358
rect 1622 1353 1623 1357
rect 1627 1353 1628 1357
rect 1622 1352 1628 1353
rect 1495 1350 1499 1352
rect 1495 1345 1499 1346
rect 1559 1350 1563 1351
rect 1559 1344 1563 1346
rect 1567 1350 1571 1352
rect 1567 1345 1571 1346
rect 1623 1350 1627 1352
rect 1623 1344 1627 1346
rect 1558 1343 1564 1344
rect 1558 1339 1559 1343
rect 1563 1339 1564 1343
rect 1558 1338 1564 1339
rect 1622 1343 1628 1344
rect 1622 1339 1623 1343
rect 1627 1339 1628 1343
rect 1622 1338 1628 1339
rect 1574 1335 1580 1336
rect 1574 1331 1575 1335
rect 1579 1331 1580 1335
rect 1574 1330 1580 1331
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1486 1319 1492 1320
rect 1486 1315 1487 1319
rect 1491 1315 1492 1319
rect 1486 1314 1492 1315
rect 1560 1307 1562 1321
rect 1576 1312 1578 1330
rect 1622 1326 1628 1327
rect 1622 1322 1623 1326
rect 1627 1322 1628 1326
rect 1622 1321 1628 1322
rect 1574 1311 1580 1312
rect 1574 1307 1575 1311
rect 1579 1307 1580 1311
rect 1624 1307 1626 1321
rect 1382 1306 1388 1307
rect 1407 1306 1411 1307
rect 1407 1301 1411 1302
rect 1447 1306 1451 1307
rect 1447 1301 1451 1302
rect 1479 1306 1483 1307
rect 1479 1301 1483 1302
rect 1543 1306 1547 1307
rect 1543 1301 1547 1302
rect 1559 1306 1563 1307
rect 1574 1306 1580 1307
rect 1623 1306 1627 1307
rect 1559 1301 1563 1302
rect 1623 1301 1627 1302
rect 1374 1295 1380 1296
rect 1374 1291 1375 1295
rect 1379 1291 1380 1295
rect 1448 1291 1450 1301
rect 1544 1291 1546 1301
rect 1624 1291 1626 1301
rect 1142 1290 1148 1291
rect 1142 1286 1143 1290
rect 1147 1286 1148 1290
rect 1142 1285 1148 1286
rect 1206 1290 1212 1291
rect 1206 1286 1207 1290
rect 1211 1286 1212 1290
rect 1206 1285 1212 1286
rect 1278 1290 1284 1291
rect 1350 1290 1356 1291
rect 1358 1290 1364 1291
rect 1374 1290 1380 1291
rect 1446 1290 1452 1291
rect 1278 1286 1279 1290
rect 1283 1286 1284 1290
rect 1278 1285 1284 1286
rect 1094 1279 1100 1280
rect 1094 1275 1095 1279
rect 1099 1275 1100 1279
rect 1154 1279 1160 1280
rect 1154 1275 1155 1279
rect 1159 1275 1160 1279
rect 1094 1274 1100 1275
rect 1152 1274 1160 1275
rect 830 1273 836 1274
rect 830 1269 831 1273
rect 835 1269 836 1273
rect 830 1268 836 1269
rect 894 1273 900 1274
rect 894 1269 895 1273
rect 899 1269 900 1273
rect 894 1268 900 1269
rect 958 1273 964 1274
rect 958 1269 959 1273
rect 963 1269 964 1273
rect 958 1268 964 1269
rect 1022 1273 1028 1274
rect 1022 1269 1023 1273
rect 1027 1269 1028 1273
rect 1022 1268 1028 1269
rect 1078 1273 1084 1274
rect 1078 1269 1079 1273
rect 1083 1269 1084 1273
rect 1078 1268 1084 1269
rect 1142 1273 1148 1274
rect 1142 1269 1143 1273
rect 1147 1269 1148 1273
rect 1142 1268 1148 1269
rect 1152 1273 1158 1274
rect 1206 1273 1212 1274
rect 815 1266 819 1267
rect 815 1260 819 1262
rect 831 1266 835 1268
rect 831 1261 835 1262
rect 871 1266 875 1267
rect 871 1260 875 1262
rect 895 1266 899 1268
rect 895 1261 899 1262
rect 927 1266 931 1267
rect 927 1260 931 1262
rect 959 1266 963 1268
rect 959 1261 963 1262
rect 983 1266 987 1267
rect 983 1260 987 1262
rect 1023 1266 1027 1268
rect 1023 1261 1027 1262
rect 1039 1266 1043 1267
rect 1039 1260 1043 1262
rect 1079 1266 1083 1268
rect 1079 1261 1083 1262
rect 1095 1266 1099 1267
rect 1095 1260 1099 1262
rect 1143 1266 1147 1268
rect 1143 1261 1147 1262
rect 814 1259 820 1260
rect 814 1255 815 1259
rect 819 1255 820 1259
rect 814 1254 820 1255
rect 870 1259 876 1260
rect 870 1255 871 1259
rect 875 1255 876 1259
rect 870 1254 876 1255
rect 926 1259 932 1260
rect 926 1255 927 1259
rect 931 1255 932 1259
rect 926 1254 932 1255
rect 982 1259 988 1260
rect 982 1255 983 1259
rect 987 1255 988 1259
rect 982 1254 988 1255
rect 1038 1259 1044 1260
rect 1038 1255 1039 1259
rect 1043 1255 1044 1259
rect 1038 1254 1044 1255
rect 1094 1259 1100 1260
rect 1094 1255 1095 1259
rect 1099 1255 1100 1259
rect 1094 1254 1100 1255
rect 782 1251 788 1252
rect 782 1247 783 1251
rect 787 1247 788 1251
rect 782 1246 788 1247
rect 1050 1251 1056 1252
rect 1050 1247 1051 1251
rect 1055 1247 1056 1251
rect 1050 1246 1056 1247
rect 766 1242 772 1243
rect 766 1238 767 1242
rect 771 1238 772 1242
rect 766 1237 772 1238
rect 814 1242 820 1243
rect 814 1238 815 1242
rect 819 1238 820 1242
rect 814 1237 820 1238
rect 870 1242 876 1243
rect 870 1238 871 1242
rect 875 1238 876 1242
rect 870 1237 876 1238
rect 926 1242 932 1243
rect 926 1238 927 1242
rect 931 1238 932 1242
rect 926 1237 932 1238
rect 982 1242 988 1243
rect 982 1238 983 1242
rect 987 1238 988 1242
rect 982 1237 988 1238
rect 1038 1242 1044 1243
rect 1038 1238 1039 1242
rect 1043 1238 1044 1242
rect 1038 1237 1044 1238
rect 758 1235 764 1236
rect 758 1231 759 1235
rect 763 1231 764 1235
rect 758 1230 764 1231
rect 768 1223 770 1237
rect 816 1223 818 1237
rect 872 1223 874 1237
rect 906 1235 912 1236
rect 906 1231 907 1235
rect 911 1231 912 1235
rect 906 1230 912 1231
rect 431 1222 435 1223
rect 431 1217 435 1218
rect 439 1222 443 1223
rect 439 1217 443 1218
rect 487 1222 491 1223
rect 487 1217 491 1218
rect 495 1222 499 1223
rect 495 1217 499 1218
rect 543 1222 547 1223
rect 543 1217 547 1218
rect 551 1222 555 1223
rect 551 1217 555 1218
rect 599 1222 603 1223
rect 599 1217 603 1218
rect 607 1222 611 1223
rect 618 1219 619 1223
rect 623 1219 624 1223
rect 618 1218 624 1219
rect 655 1222 659 1223
rect 607 1217 611 1218
rect 655 1217 659 1218
rect 663 1222 667 1223
rect 663 1217 667 1218
rect 711 1222 715 1223
rect 711 1217 715 1218
rect 719 1222 723 1223
rect 719 1217 723 1218
rect 767 1222 771 1223
rect 767 1217 771 1218
rect 815 1222 819 1223
rect 815 1217 819 1218
rect 823 1222 827 1223
rect 823 1217 827 1218
rect 871 1222 875 1223
rect 871 1217 875 1218
rect 887 1222 891 1223
rect 887 1217 891 1218
rect 432 1207 434 1217
rect 488 1207 490 1217
rect 544 1207 546 1217
rect 600 1207 602 1217
rect 656 1207 658 1217
rect 712 1207 714 1217
rect 768 1207 770 1217
rect 782 1211 788 1212
rect 782 1207 783 1211
rect 787 1207 788 1211
rect 824 1207 826 1217
rect 888 1207 890 1217
rect 430 1206 436 1207
rect 430 1202 431 1206
rect 435 1202 436 1206
rect 430 1201 436 1202
rect 486 1206 492 1207
rect 486 1202 487 1206
rect 491 1202 492 1206
rect 486 1201 492 1202
rect 542 1206 548 1207
rect 542 1202 543 1206
rect 547 1202 548 1206
rect 542 1201 548 1202
rect 598 1206 604 1207
rect 598 1202 599 1206
rect 603 1202 604 1206
rect 598 1201 604 1202
rect 654 1206 660 1207
rect 654 1202 655 1206
rect 659 1202 660 1206
rect 654 1201 660 1202
rect 710 1206 716 1207
rect 710 1202 711 1206
rect 715 1202 716 1206
rect 710 1201 716 1202
rect 766 1206 772 1207
rect 782 1206 788 1207
rect 822 1206 828 1207
rect 766 1202 767 1206
rect 771 1202 772 1206
rect 766 1201 772 1202
rect 306 1195 312 1196
rect 306 1191 307 1195
rect 311 1191 312 1195
rect 306 1190 312 1191
rect 398 1195 404 1196
rect 398 1191 399 1195
rect 403 1191 404 1195
rect 398 1190 404 1191
rect 334 1189 340 1190
rect 334 1185 335 1189
rect 339 1185 340 1189
rect 334 1184 340 1185
rect 382 1189 388 1190
rect 382 1185 383 1189
rect 387 1185 388 1189
rect 382 1184 388 1185
rect 430 1189 436 1190
rect 430 1185 431 1189
rect 435 1185 436 1189
rect 430 1184 436 1185
rect 486 1189 492 1190
rect 486 1185 487 1189
rect 491 1185 492 1189
rect 486 1184 492 1185
rect 542 1189 548 1190
rect 542 1185 543 1189
rect 547 1185 548 1189
rect 542 1184 548 1185
rect 598 1189 604 1190
rect 598 1185 599 1189
rect 603 1185 604 1189
rect 598 1184 604 1185
rect 654 1189 660 1190
rect 654 1185 655 1189
rect 659 1185 660 1189
rect 654 1184 660 1185
rect 710 1189 716 1190
rect 710 1185 711 1189
rect 715 1185 716 1189
rect 710 1184 716 1185
rect 766 1189 772 1190
rect 766 1185 767 1189
rect 771 1185 772 1189
rect 784 1188 786 1206
rect 822 1202 823 1206
rect 827 1202 828 1206
rect 822 1201 828 1202
rect 886 1206 892 1207
rect 886 1202 887 1206
rect 891 1202 892 1206
rect 886 1201 892 1202
rect 908 1196 910 1230
rect 928 1223 930 1237
rect 984 1223 986 1237
rect 1040 1223 1042 1237
rect 1052 1228 1054 1246
rect 1094 1242 1100 1243
rect 1094 1238 1095 1242
rect 1099 1238 1100 1242
rect 1094 1237 1100 1238
rect 1050 1227 1056 1228
rect 1050 1223 1051 1227
rect 1055 1223 1056 1227
rect 1096 1223 1098 1237
rect 1152 1236 1154 1273
rect 1206 1269 1207 1273
rect 1211 1269 1212 1273
rect 1206 1268 1212 1269
rect 1278 1273 1284 1274
rect 1278 1269 1279 1273
rect 1283 1269 1284 1273
rect 1278 1268 1284 1269
rect 1352 1268 1354 1290
rect 1358 1286 1359 1290
rect 1363 1286 1364 1290
rect 1358 1285 1364 1286
rect 1446 1286 1447 1290
rect 1451 1286 1452 1290
rect 1446 1285 1452 1286
rect 1542 1290 1548 1291
rect 1542 1286 1543 1290
rect 1547 1286 1548 1290
rect 1542 1285 1548 1286
rect 1622 1290 1628 1291
rect 1622 1286 1623 1290
rect 1627 1286 1628 1290
rect 1622 1285 1628 1286
rect 1644 1280 1646 1374
rect 1662 1372 1663 1376
rect 1667 1372 1668 1376
rect 1662 1371 1668 1372
rect 1662 1359 1668 1360
rect 1662 1355 1663 1359
rect 1667 1355 1668 1359
rect 1662 1354 1668 1355
rect 1664 1351 1666 1354
rect 1663 1350 1667 1351
rect 1663 1345 1667 1346
rect 1664 1342 1666 1345
rect 1662 1341 1668 1342
rect 1662 1337 1663 1341
rect 1667 1337 1668 1341
rect 1662 1336 1668 1337
rect 1650 1335 1656 1336
rect 1650 1331 1651 1335
rect 1655 1331 1656 1335
rect 1650 1330 1656 1331
rect 1642 1279 1648 1280
rect 1642 1275 1643 1279
rect 1647 1275 1648 1279
rect 1642 1274 1648 1275
rect 1358 1273 1364 1274
rect 1358 1269 1359 1273
rect 1363 1269 1364 1273
rect 1358 1268 1364 1269
rect 1446 1273 1452 1274
rect 1446 1269 1447 1273
rect 1451 1269 1452 1273
rect 1446 1268 1452 1269
rect 1542 1273 1548 1274
rect 1542 1269 1543 1273
rect 1547 1269 1548 1273
rect 1542 1268 1548 1269
rect 1622 1273 1628 1274
rect 1622 1269 1623 1273
rect 1627 1269 1628 1273
rect 1622 1268 1628 1269
rect 1159 1266 1163 1267
rect 1159 1260 1163 1262
rect 1207 1266 1211 1268
rect 1207 1261 1211 1262
rect 1231 1266 1235 1267
rect 1231 1260 1235 1262
rect 1279 1266 1283 1268
rect 1350 1267 1356 1268
rect 1279 1261 1283 1262
rect 1319 1266 1323 1267
rect 1350 1263 1351 1267
rect 1355 1263 1356 1267
rect 1350 1262 1356 1263
rect 1359 1266 1363 1268
rect 1319 1260 1323 1262
rect 1359 1261 1363 1262
rect 1423 1266 1427 1267
rect 1423 1260 1427 1262
rect 1447 1266 1451 1268
rect 1447 1261 1451 1262
rect 1535 1266 1539 1267
rect 1535 1260 1539 1262
rect 1543 1266 1547 1268
rect 1543 1261 1547 1262
rect 1623 1266 1627 1268
rect 1623 1260 1627 1262
rect 1158 1259 1164 1260
rect 1158 1255 1159 1259
rect 1163 1255 1164 1259
rect 1158 1254 1164 1255
rect 1230 1259 1236 1260
rect 1230 1255 1231 1259
rect 1235 1255 1236 1259
rect 1230 1254 1236 1255
rect 1318 1259 1324 1260
rect 1318 1255 1319 1259
rect 1323 1255 1324 1259
rect 1318 1254 1324 1255
rect 1422 1259 1428 1260
rect 1422 1255 1423 1259
rect 1427 1255 1428 1259
rect 1422 1254 1428 1255
rect 1534 1259 1540 1260
rect 1534 1255 1535 1259
rect 1539 1255 1540 1259
rect 1534 1254 1540 1255
rect 1622 1259 1628 1260
rect 1622 1255 1623 1259
rect 1627 1255 1628 1259
rect 1622 1254 1628 1255
rect 1502 1251 1508 1252
rect 1502 1247 1503 1251
rect 1507 1247 1508 1251
rect 1502 1246 1508 1247
rect 1638 1251 1644 1252
rect 1638 1247 1639 1251
rect 1643 1247 1644 1251
rect 1638 1246 1644 1247
rect 1158 1242 1164 1243
rect 1158 1238 1159 1242
rect 1163 1238 1164 1242
rect 1158 1237 1164 1238
rect 1230 1242 1236 1243
rect 1230 1238 1231 1242
rect 1235 1238 1236 1242
rect 1230 1237 1236 1238
rect 1318 1242 1324 1243
rect 1318 1238 1319 1242
rect 1323 1238 1324 1242
rect 1318 1237 1324 1238
rect 1422 1242 1428 1243
rect 1422 1238 1423 1242
rect 1427 1238 1428 1242
rect 1422 1237 1428 1238
rect 1150 1235 1156 1236
rect 1150 1231 1151 1235
rect 1155 1231 1156 1235
rect 1150 1230 1156 1231
rect 1160 1223 1162 1237
rect 1232 1223 1234 1237
rect 1320 1223 1322 1237
rect 1424 1223 1426 1237
rect 1504 1224 1506 1246
rect 1534 1242 1540 1243
rect 1534 1238 1535 1242
rect 1539 1238 1540 1242
rect 1534 1237 1540 1238
rect 1622 1242 1628 1243
rect 1622 1238 1623 1242
rect 1627 1238 1628 1242
rect 1622 1237 1628 1238
rect 1502 1223 1508 1224
rect 1536 1223 1538 1237
rect 1624 1223 1626 1237
rect 927 1222 931 1223
rect 927 1217 931 1218
rect 951 1222 955 1223
rect 951 1217 955 1218
rect 983 1222 987 1223
rect 983 1217 987 1218
rect 1015 1222 1019 1223
rect 1015 1217 1019 1218
rect 1039 1222 1043 1223
rect 1050 1222 1056 1223
rect 1079 1222 1083 1223
rect 1039 1217 1043 1218
rect 1079 1217 1083 1218
rect 1095 1222 1099 1223
rect 1095 1217 1099 1218
rect 1143 1222 1147 1223
rect 1143 1217 1147 1218
rect 1159 1222 1163 1223
rect 1159 1217 1163 1218
rect 1207 1222 1211 1223
rect 1207 1217 1211 1218
rect 1231 1222 1235 1223
rect 1231 1217 1235 1218
rect 1279 1222 1283 1223
rect 1279 1217 1283 1218
rect 1319 1222 1323 1223
rect 1319 1217 1323 1218
rect 1359 1222 1363 1223
rect 1359 1217 1363 1218
rect 1423 1222 1427 1223
rect 1423 1217 1427 1218
rect 1447 1222 1451 1223
rect 1502 1219 1503 1223
rect 1507 1219 1508 1223
rect 1502 1218 1508 1219
rect 1535 1222 1539 1223
rect 1447 1217 1451 1218
rect 1535 1217 1539 1218
rect 1543 1222 1547 1223
rect 1543 1217 1547 1218
rect 1623 1222 1627 1223
rect 1623 1217 1627 1218
rect 952 1207 954 1217
rect 1006 1211 1012 1212
rect 1006 1207 1007 1211
rect 1011 1207 1012 1211
rect 1016 1207 1018 1217
rect 1022 1211 1028 1212
rect 1022 1207 1023 1211
rect 1027 1207 1028 1211
rect 1080 1207 1082 1217
rect 1144 1207 1146 1217
rect 1208 1207 1210 1217
rect 1280 1207 1282 1217
rect 1360 1207 1362 1217
rect 1448 1207 1450 1217
rect 1544 1207 1546 1217
rect 1624 1207 1626 1217
rect 1640 1212 1642 1246
rect 1652 1236 1654 1330
rect 1662 1324 1668 1325
rect 1662 1320 1663 1324
rect 1667 1320 1668 1324
rect 1662 1319 1668 1320
rect 1664 1307 1666 1319
rect 1663 1306 1667 1307
rect 1663 1301 1667 1302
rect 1664 1293 1666 1301
rect 1662 1292 1668 1293
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1662 1275 1668 1276
rect 1662 1271 1663 1275
rect 1667 1271 1668 1275
rect 1662 1270 1668 1271
rect 1664 1267 1666 1270
rect 1663 1266 1667 1267
rect 1663 1261 1667 1262
rect 1664 1258 1666 1261
rect 1662 1257 1668 1258
rect 1662 1253 1663 1257
rect 1667 1253 1668 1257
rect 1662 1252 1668 1253
rect 1662 1240 1668 1241
rect 1662 1236 1663 1240
rect 1667 1236 1668 1240
rect 1650 1235 1656 1236
rect 1662 1235 1668 1236
rect 1650 1231 1651 1235
rect 1655 1231 1656 1235
rect 1650 1230 1656 1231
rect 1664 1223 1666 1235
rect 1663 1222 1667 1223
rect 1663 1217 1667 1218
rect 1638 1211 1644 1212
rect 1638 1207 1639 1211
rect 1643 1207 1644 1211
rect 1664 1209 1666 1217
rect 950 1206 956 1207
rect 1006 1206 1012 1207
rect 1014 1206 1020 1207
rect 1022 1206 1028 1207
rect 1078 1206 1084 1207
rect 950 1202 951 1206
rect 955 1202 956 1206
rect 950 1201 956 1202
rect 906 1195 912 1196
rect 906 1191 907 1195
rect 911 1191 912 1195
rect 906 1190 912 1191
rect 822 1189 828 1190
rect 766 1184 772 1185
rect 782 1187 788 1188
rect 336 1179 338 1184
rect 384 1179 386 1184
rect 432 1179 434 1184
rect 488 1179 490 1184
rect 494 1183 500 1184
rect 494 1179 495 1183
rect 499 1179 500 1183
rect 544 1179 546 1184
rect 600 1179 602 1184
rect 656 1179 658 1184
rect 712 1179 714 1184
rect 768 1179 770 1184
rect 782 1183 783 1187
rect 787 1183 788 1187
rect 822 1185 823 1189
rect 827 1185 828 1189
rect 822 1184 828 1185
rect 886 1189 892 1190
rect 886 1185 887 1189
rect 891 1185 892 1189
rect 886 1184 892 1185
rect 950 1189 956 1190
rect 950 1185 951 1189
rect 955 1185 956 1189
rect 950 1184 956 1185
rect 1008 1184 1010 1206
rect 1014 1202 1015 1206
rect 1019 1202 1020 1206
rect 1014 1201 1020 1202
rect 1014 1189 1020 1190
rect 1014 1185 1015 1189
rect 1019 1185 1020 1189
rect 1014 1184 1020 1185
rect 782 1182 788 1183
rect 824 1179 826 1184
rect 888 1179 890 1184
rect 952 1179 954 1184
rect 1006 1183 1012 1184
rect 1006 1179 1007 1183
rect 1011 1179 1012 1183
rect 1016 1179 1018 1184
rect 335 1178 339 1179
rect 335 1173 339 1174
rect 351 1178 355 1179
rect 351 1172 355 1174
rect 383 1178 387 1179
rect 383 1173 387 1174
rect 415 1178 419 1179
rect 415 1172 419 1174
rect 431 1178 435 1179
rect 431 1173 435 1174
rect 471 1178 475 1179
rect 471 1172 475 1174
rect 487 1178 491 1179
rect 494 1178 500 1179
rect 535 1178 539 1179
rect 487 1173 491 1174
rect 350 1171 356 1172
rect 350 1167 351 1171
rect 355 1167 356 1171
rect 350 1166 356 1167
rect 414 1171 420 1172
rect 414 1167 415 1171
rect 419 1167 420 1171
rect 414 1166 420 1167
rect 470 1171 476 1172
rect 470 1167 471 1171
rect 475 1167 476 1171
rect 470 1166 476 1167
rect 298 1163 304 1164
rect 298 1159 299 1163
rect 303 1159 304 1163
rect 298 1158 304 1159
rect 286 1154 292 1155
rect 286 1150 287 1154
rect 291 1150 292 1154
rect 286 1149 292 1150
rect 350 1154 356 1155
rect 350 1150 351 1154
rect 355 1150 356 1154
rect 350 1149 356 1150
rect 414 1154 420 1155
rect 414 1150 415 1154
rect 419 1150 420 1154
rect 414 1149 420 1150
rect 470 1154 476 1155
rect 470 1150 471 1154
rect 475 1150 476 1154
rect 470 1149 476 1150
rect 238 1147 244 1148
rect 238 1143 239 1147
rect 243 1143 244 1147
rect 238 1142 244 1143
rect 288 1135 290 1149
rect 352 1135 354 1149
rect 416 1135 418 1149
rect 472 1135 474 1149
rect 478 1147 484 1148
rect 478 1143 479 1147
rect 483 1143 484 1147
rect 478 1142 484 1143
rect 487 1147 493 1148
rect 487 1143 488 1147
rect 492 1146 493 1147
rect 496 1146 498 1178
rect 535 1172 539 1174
rect 543 1178 547 1179
rect 543 1173 547 1174
rect 599 1178 603 1179
rect 599 1172 603 1174
rect 655 1178 659 1179
rect 655 1173 659 1174
rect 663 1178 667 1179
rect 663 1172 667 1174
rect 711 1178 715 1179
rect 711 1173 715 1174
rect 727 1178 731 1179
rect 727 1172 731 1174
rect 767 1178 771 1179
rect 767 1173 771 1174
rect 783 1178 787 1179
rect 783 1172 787 1174
rect 823 1178 827 1179
rect 823 1173 827 1174
rect 839 1178 843 1179
rect 887 1178 891 1179
rect 839 1172 843 1174
rect 858 1175 864 1176
rect 534 1171 540 1172
rect 534 1167 535 1171
rect 539 1167 540 1171
rect 534 1166 540 1167
rect 598 1171 604 1172
rect 598 1167 599 1171
rect 603 1167 604 1171
rect 598 1166 604 1167
rect 662 1171 668 1172
rect 662 1167 663 1171
rect 667 1167 668 1171
rect 662 1166 668 1167
rect 726 1171 732 1172
rect 726 1167 727 1171
rect 731 1167 732 1171
rect 726 1166 732 1167
rect 782 1171 788 1172
rect 782 1167 783 1171
rect 787 1167 788 1171
rect 782 1166 788 1167
rect 838 1171 844 1172
rect 838 1167 839 1171
rect 843 1167 844 1171
rect 858 1171 859 1175
rect 863 1171 864 1175
rect 887 1173 891 1174
rect 903 1178 907 1179
rect 903 1172 907 1174
rect 951 1178 955 1179
rect 951 1173 955 1174
rect 967 1178 971 1179
rect 1006 1178 1012 1179
rect 1015 1178 1019 1179
rect 967 1172 971 1174
rect 1015 1173 1019 1174
rect 858 1170 864 1171
rect 902 1171 908 1172
rect 838 1166 844 1167
rect 798 1163 804 1164
rect 798 1159 799 1163
rect 803 1159 804 1163
rect 798 1158 804 1159
rect 534 1154 540 1155
rect 534 1150 535 1154
rect 539 1150 540 1154
rect 534 1149 540 1150
rect 598 1154 604 1155
rect 598 1150 599 1154
rect 603 1150 604 1154
rect 598 1149 604 1150
rect 662 1154 668 1155
rect 662 1150 663 1154
rect 667 1150 668 1154
rect 662 1149 668 1150
rect 726 1154 732 1155
rect 726 1150 727 1154
rect 731 1150 732 1154
rect 726 1149 732 1150
rect 782 1154 788 1155
rect 782 1150 783 1154
rect 787 1150 788 1154
rect 782 1149 788 1150
rect 492 1144 498 1146
rect 492 1143 493 1144
rect 487 1142 493 1143
rect 167 1134 171 1135
rect 167 1129 171 1130
rect 175 1134 179 1135
rect 175 1129 179 1130
rect 215 1134 219 1135
rect 215 1129 219 1130
rect 223 1134 227 1135
rect 223 1129 227 1130
rect 271 1134 275 1135
rect 271 1129 275 1130
rect 287 1134 291 1135
rect 287 1129 291 1130
rect 335 1134 339 1135
rect 335 1129 339 1130
rect 351 1134 355 1135
rect 351 1129 355 1130
rect 399 1134 403 1135
rect 399 1129 403 1130
rect 415 1134 419 1135
rect 415 1129 419 1130
rect 463 1134 467 1135
rect 463 1129 467 1130
rect 471 1134 475 1135
rect 471 1129 475 1130
rect 154 1123 160 1124
rect 154 1119 155 1123
rect 159 1119 160 1123
rect 176 1119 178 1129
rect 216 1119 218 1129
rect 272 1119 274 1129
rect 298 1127 304 1128
rect 298 1123 299 1127
rect 303 1123 304 1127
rect 298 1122 304 1123
rect 110 1115 116 1116
rect 142 1118 148 1119
rect 154 1118 160 1119
rect 174 1118 180 1119
rect 142 1114 143 1118
rect 147 1114 148 1118
rect 142 1113 148 1114
rect 174 1114 175 1118
rect 179 1114 180 1118
rect 174 1113 180 1114
rect 214 1118 220 1119
rect 214 1114 215 1118
rect 219 1114 220 1118
rect 214 1113 220 1114
rect 270 1118 276 1119
rect 270 1114 271 1118
rect 275 1114 276 1118
rect 270 1113 276 1114
rect 110 1103 116 1104
rect 110 1099 111 1103
rect 115 1099 116 1103
rect 110 1098 116 1099
rect 142 1101 148 1102
rect 112 1091 114 1098
rect 142 1097 143 1101
rect 147 1097 148 1101
rect 142 1096 148 1097
rect 174 1101 180 1102
rect 174 1097 175 1101
rect 179 1097 180 1101
rect 174 1096 180 1097
rect 214 1101 220 1102
rect 214 1097 215 1101
rect 219 1097 220 1101
rect 214 1096 220 1097
rect 270 1101 276 1102
rect 270 1097 271 1101
rect 275 1097 276 1101
rect 270 1096 276 1097
rect 144 1091 146 1096
rect 176 1091 178 1096
rect 216 1091 218 1096
rect 234 1095 240 1096
rect 234 1091 235 1095
rect 239 1091 240 1095
rect 272 1091 274 1096
rect 111 1090 115 1091
rect 111 1085 115 1086
rect 143 1090 147 1091
rect 143 1085 147 1086
rect 175 1090 179 1091
rect 175 1085 179 1086
rect 215 1090 219 1091
rect 234 1090 240 1091
rect 247 1090 251 1091
rect 112 1082 114 1085
rect 215 1084 219 1086
rect 214 1083 220 1084
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 214 1079 215 1083
rect 219 1079 220 1083
rect 214 1078 220 1079
rect 110 1076 116 1077
rect 214 1066 220 1067
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 214 1062 215 1066
rect 219 1062 220 1066
rect 214 1061 220 1062
rect 110 1059 116 1060
rect 112 1047 114 1059
rect 216 1047 218 1061
rect 236 1060 238 1090
rect 247 1084 251 1086
rect 271 1090 275 1091
rect 271 1085 275 1086
rect 279 1090 283 1091
rect 279 1084 283 1086
rect 246 1083 252 1084
rect 246 1079 247 1083
rect 251 1079 252 1083
rect 246 1078 252 1079
rect 278 1083 284 1084
rect 278 1079 279 1083
rect 283 1079 284 1083
rect 278 1078 284 1079
rect 300 1076 302 1122
rect 336 1119 338 1129
rect 400 1119 402 1129
rect 464 1119 466 1129
rect 334 1118 340 1119
rect 334 1114 335 1118
rect 339 1114 340 1118
rect 334 1113 340 1114
rect 398 1118 404 1119
rect 398 1114 399 1118
rect 403 1114 404 1118
rect 398 1113 404 1114
rect 462 1118 468 1119
rect 462 1114 463 1118
rect 467 1114 468 1118
rect 462 1113 468 1114
rect 480 1108 482 1142
rect 536 1135 538 1149
rect 600 1135 602 1149
rect 664 1135 666 1149
rect 728 1135 730 1149
rect 784 1135 786 1149
rect 800 1136 802 1158
rect 838 1154 844 1155
rect 838 1150 839 1154
rect 843 1150 844 1154
rect 838 1149 844 1150
rect 798 1135 804 1136
rect 840 1135 842 1149
rect 860 1148 862 1170
rect 902 1167 903 1171
rect 907 1167 908 1171
rect 902 1166 908 1167
rect 966 1171 972 1172
rect 966 1167 967 1171
rect 971 1167 972 1171
rect 966 1166 972 1167
rect 1024 1164 1026 1206
rect 1078 1202 1079 1206
rect 1083 1202 1084 1206
rect 1078 1201 1084 1202
rect 1142 1206 1148 1207
rect 1142 1202 1143 1206
rect 1147 1202 1148 1206
rect 1142 1201 1148 1202
rect 1206 1206 1212 1207
rect 1206 1202 1207 1206
rect 1211 1202 1212 1206
rect 1206 1201 1212 1202
rect 1278 1206 1284 1207
rect 1278 1202 1279 1206
rect 1283 1202 1284 1206
rect 1278 1201 1284 1202
rect 1358 1206 1364 1207
rect 1358 1202 1359 1206
rect 1363 1202 1364 1206
rect 1358 1201 1364 1202
rect 1446 1206 1452 1207
rect 1446 1202 1447 1206
rect 1451 1202 1452 1206
rect 1446 1201 1452 1202
rect 1542 1206 1548 1207
rect 1542 1202 1543 1206
rect 1547 1202 1548 1206
rect 1542 1201 1548 1202
rect 1622 1206 1628 1207
rect 1638 1206 1644 1207
rect 1662 1208 1668 1209
rect 1622 1202 1623 1206
rect 1627 1202 1628 1206
rect 1662 1204 1663 1208
rect 1667 1204 1668 1208
rect 1662 1203 1668 1204
rect 1622 1201 1628 1202
rect 1638 1195 1644 1196
rect 1638 1191 1639 1195
rect 1643 1191 1644 1195
rect 1638 1190 1644 1191
rect 1662 1191 1668 1192
rect 1078 1189 1084 1190
rect 1078 1185 1079 1189
rect 1083 1185 1084 1189
rect 1078 1184 1084 1185
rect 1142 1189 1148 1190
rect 1142 1185 1143 1189
rect 1147 1185 1148 1189
rect 1142 1184 1148 1185
rect 1206 1189 1212 1190
rect 1206 1185 1207 1189
rect 1211 1185 1212 1189
rect 1206 1184 1212 1185
rect 1278 1189 1284 1190
rect 1278 1185 1279 1189
rect 1283 1185 1284 1189
rect 1278 1184 1284 1185
rect 1358 1189 1364 1190
rect 1358 1185 1359 1189
rect 1363 1185 1364 1189
rect 1358 1184 1364 1185
rect 1446 1189 1452 1190
rect 1446 1185 1447 1189
rect 1451 1185 1452 1189
rect 1446 1184 1452 1185
rect 1542 1189 1548 1190
rect 1542 1185 1543 1189
rect 1547 1185 1548 1189
rect 1542 1184 1548 1185
rect 1622 1189 1628 1190
rect 1622 1185 1623 1189
rect 1627 1185 1628 1189
rect 1622 1184 1628 1185
rect 1080 1179 1082 1184
rect 1144 1179 1146 1184
rect 1208 1179 1210 1184
rect 1234 1183 1240 1184
rect 1234 1179 1235 1183
rect 1239 1179 1240 1183
rect 1280 1179 1282 1184
rect 1360 1179 1362 1184
rect 1448 1179 1450 1184
rect 1544 1179 1546 1184
rect 1624 1179 1626 1184
rect 1031 1178 1035 1179
rect 1031 1172 1035 1174
rect 1079 1178 1083 1179
rect 1079 1173 1083 1174
rect 1095 1178 1099 1179
rect 1095 1172 1099 1174
rect 1143 1178 1147 1179
rect 1143 1173 1147 1174
rect 1159 1178 1163 1179
rect 1159 1172 1163 1174
rect 1207 1178 1211 1179
rect 1207 1173 1211 1174
rect 1215 1178 1219 1179
rect 1234 1178 1240 1179
rect 1279 1178 1283 1179
rect 1215 1172 1219 1174
rect 1030 1171 1036 1172
rect 1030 1167 1031 1171
rect 1035 1167 1036 1171
rect 1030 1166 1036 1167
rect 1094 1171 1100 1172
rect 1094 1167 1095 1171
rect 1099 1167 1100 1171
rect 1094 1166 1100 1167
rect 1158 1171 1164 1172
rect 1158 1167 1159 1171
rect 1163 1167 1164 1171
rect 1158 1166 1164 1167
rect 1214 1171 1220 1172
rect 1214 1167 1215 1171
rect 1219 1167 1220 1171
rect 1214 1166 1220 1167
rect 1022 1163 1028 1164
rect 1022 1159 1023 1163
rect 1027 1159 1028 1163
rect 1022 1158 1028 1159
rect 902 1154 908 1155
rect 902 1150 903 1154
rect 907 1150 908 1154
rect 902 1149 908 1150
rect 966 1154 972 1155
rect 966 1150 967 1154
rect 971 1150 972 1154
rect 966 1149 972 1150
rect 1030 1154 1036 1155
rect 1030 1150 1031 1154
rect 1035 1150 1036 1154
rect 1030 1149 1036 1150
rect 1094 1154 1100 1155
rect 1094 1150 1095 1154
rect 1099 1150 1100 1154
rect 1094 1149 1100 1150
rect 1158 1154 1164 1155
rect 1158 1150 1159 1154
rect 1163 1150 1164 1154
rect 1158 1149 1164 1150
rect 1214 1154 1220 1155
rect 1214 1150 1215 1154
rect 1219 1150 1220 1154
rect 1214 1149 1220 1150
rect 858 1147 864 1148
rect 858 1143 859 1147
rect 863 1143 864 1147
rect 858 1142 864 1143
rect 904 1135 906 1149
rect 968 1135 970 1149
rect 1032 1135 1034 1149
rect 1042 1147 1048 1148
rect 1042 1143 1043 1147
rect 1047 1143 1048 1147
rect 1042 1142 1048 1143
rect 527 1134 531 1135
rect 527 1129 531 1130
rect 535 1134 539 1135
rect 535 1129 539 1130
rect 599 1134 603 1135
rect 599 1129 603 1130
rect 663 1134 667 1135
rect 663 1129 667 1130
rect 727 1134 731 1135
rect 727 1129 731 1130
rect 783 1134 787 1135
rect 783 1129 787 1130
rect 791 1134 795 1135
rect 798 1131 799 1135
rect 803 1131 804 1135
rect 798 1130 804 1131
rect 839 1134 843 1135
rect 791 1129 795 1130
rect 839 1129 843 1130
rect 855 1134 859 1135
rect 855 1129 859 1130
rect 903 1134 907 1135
rect 903 1129 907 1130
rect 911 1134 915 1135
rect 911 1129 915 1130
rect 967 1134 971 1135
rect 967 1129 971 1130
rect 1023 1134 1027 1135
rect 1023 1129 1027 1130
rect 1031 1134 1035 1135
rect 1031 1129 1035 1130
rect 528 1119 530 1129
rect 600 1119 602 1129
rect 664 1119 666 1129
rect 728 1119 730 1129
rect 792 1119 794 1129
rect 856 1119 858 1129
rect 912 1119 914 1129
rect 968 1119 970 1129
rect 1024 1119 1026 1129
rect 526 1118 532 1119
rect 526 1114 527 1118
rect 531 1114 532 1118
rect 526 1113 532 1114
rect 598 1118 604 1119
rect 598 1114 599 1118
rect 603 1114 604 1118
rect 598 1113 604 1114
rect 662 1118 668 1119
rect 662 1114 663 1118
rect 667 1114 668 1118
rect 662 1113 668 1114
rect 726 1118 732 1119
rect 726 1114 727 1118
rect 731 1114 732 1118
rect 726 1113 732 1114
rect 790 1118 796 1119
rect 790 1114 791 1118
rect 795 1114 796 1118
rect 790 1113 796 1114
rect 854 1118 860 1119
rect 854 1114 855 1118
rect 859 1114 860 1118
rect 854 1113 860 1114
rect 910 1118 916 1119
rect 910 1114 911 1118
rect 915 1114 916 1118
rect 910 1113 916 1114
rect 966 1118 972 1119
rect 966 1114 967 1118
rect 971 1114 972 1118
rect 966 1113 972 1114
rect 1022 1118 1028 1119
rect 1022 1114 1023 1118
rect 1027 1114 1028 1118
rect 1022 1113 1028 1114
rect 1044 1108 1046 1142
rect 1096 1135 1098 1149
rect 1102 1135 1108 1136
rect 1160 1135 1162 1149
rect 1216 1135 1218 1149
rect 1236 1148 1238 1178
rect 1279 1172 1283 1174
rect 1343 1178 1347 1179
rect 1343 1172 1347 1174
rect 1359 1178 1363 1179
rect 1359 1173 1363 1174
rect 1407 1178 1411 1179
rect 1407 1172 1411 1174
rect 1447 1178 1451 1179
rect 1447 1173 1451 1174
rect 1479 1178 1483 1179
rect 1479 1172 1483 1174
rect 1543 1178 1547 1179
rect 1543 1173 1547 1174
rect 1559 1178 1563 1179
rect 1559 1172 1563 1174
rect 1623 1178 1627 1179
rect 1623 1172 1627 1174
rect 1278 1171 1284 1172
rect 1278 1167 1279 1171
rect 1283 1167 1284 1171
rect 1278 1166 1284 1167
rect 1342 1171 1348 1172
rect 1342 1167 1343 1171
rect 1347 1167 1348 1171
rect 1342 1166 1348 1167
rect 1406 1171 1412 1172
rect 1406 1167 1407 1171
rect 1411 1167 1412 1171
rect 1406 1166 1412 1167
rect 1478 1171 1484 1172
rect 1478 1167 1479 1171
rect 1483 1167 1484 1171
rect 1478 1166 1484 1167
rect 1558 1171 1564 1172
rect 1558 1167 1559 1171
rect 1563 1167 1564 1171
rect 1558 1166 1564 1167
rect 1622 1171 1628 1172
rect 1622 1167 1623 1171
rect 1627 1167 1628 1171
rect 1622 1166 1628 1167
rect 1278 1154 1284 1155
rect 1278 1150 1279 1154
rect 1283 1150 1284 1154
rect 1278 1149 1284 1150
rect 1342 1154 1348 1155
rect 1342 1150 1343 1154
rect 1347 1150 1348 1154
rect 1342 1149 1348 1150
rect 1406 1154 1412 1155
rect 1406 1150 1407 1154
rect 1411 1150 1412 1154
rect 1406 1149 1412 1150
rect 1478 1154 1484 1155
rect 1478 1150 1479 1154
rect 1483 1150 1484 1154
rect 1478 1149 1484 1150
rect 1558 1154 1564 1155
rect 1558 1150 1559 1154
rect 1563 1150 1564 1154
rect 1558 1149 1564 1150
rect 1622 1154 1628 1155
rect 1622 1150 1623 1154
rect 1627 1150 1628 1154
rect 1622 1149 1628 1150
rect 1234 1147 1240 1148
rect 1234 1143 1235 1147
rect 1239 1143 1240 1147
rect 1234 1142 1240 1143
rect 1280 1135 1282 1149
rect 1344 1135 1346 1149
rect 1408 1135 1410 1149
rect 1480 1135 1482 1149
rect 1560 1135 1562 1149
rect 1624 1135 1626 1149
rect 1640 1148 1642 1190
rect 1662 1187 1663 1191
rect 1667 1187 1668 1191
rect 1662 1186 1668 1187
rect 1664 1179 1666 1186
rect 1663 1178 1667 1179
rect 1663 1173 1667 1174
rect 1664 1170 1666 1173
rect 1662 1169 1668 1170
rect 1662 1165 1663 1169
rect 1667 1165 1668 1169
rect 1662 1164 1668 1165
rect 1662 1152 1668 1153
rect 1662 1148 1663 1152
rect 1667 1148 1668 1152
rect 1638 1147 1644 1148
rect 1662 1147 1668 1148
rect 1638 1143 1639 1147
rect 1643 1143 1644 1147
rect 1638 1142 1644 1143
rect 1664 1135 1666 1147
rect 1087 1134 1091 1135
rect 1087 1129 1091 1130
rect 1095 1134 1099 1135
rect 1102 1131 1103 1135
rect 1107 1131 1108 1135
rect 1102 1130 1108 1131
rect 1151 1134 1155 1135
rect 1095 1129 1099 1130
rect 1088 1119 1090 1129
rect 1086 1118 1092 1119
rect 1086 1114 1087 1118
rect 1091 1114 1092 1118
rect 1086 1113 1092 1114
rect 1104 1108 1106 1130
rect 1151 1129 1155 1130
rect 1159 1134 1163 1135
rect 1159 1129 1163 1130
rect 1215 1134 1219 1135
rect 1215 1129 1219 1130
rect 1279 1134 1283 1135
rect 1279 1129 1283 1130
rect 1335 1134 1339 1135
rect 1335 1129 1339 1130
rect 1343 1134 1347 1135
rect 1343 1129 1347 1130
rect 1391 1134 1395 1135
rect 1391 1129 1395 1130
rect 1407 1134 1411 1135
rect 1407 1129 1411 1130
rect 1447 1134 1451 1135
rect 1447 1129 1451 1130
rect 1479 1134 1483 1135
rect 1479 1129 1483 1130
rect 1495 1134 1499 1135
rect 1495 1129 1499 1130
rect 1543 1134 1547 1135
rect 1543 1129 1547 1130
rect 1559 1134 1563 1135
rect 1559 1129 1563 1130
rect 1591 1134 1595 1135
rect 1591 1129 1595 1130
rect 1623 1134 1627 1135
rect 1623 1129 1627 1130
rect 1663 1134 1667 1135
rect 1663 1129 1667 1130
rect 1130 1123 1136 1124
rect 1130 1119 1131 1123
rect 1135 1119 1136 1123
rect 1152 1119 1154 1129
rect 1162 1123 1168 1124
rect 1162 1119 1163 1123
rect 1167 1119 1168 1123
rect 1216 1119 1218 1129
rect 1280 1119 1282 1129
rect 1336 1119 1338 1129
rect 1392 1119 1394 1129
rect 1448 1119 1450 1129
rect 1496 1119 1498 1129
rect 1544 1119 1546 1129
rect 1558 1123 1564 1124
rect 1558 1119 1559 1123
rect 1563 1119 1564 1123
rect 1592 1119 1594 1129
rect 1624 1119 1626 1129
rect 1664 1121 1666 1129
rect 1662 1120 1668 1121
rect 1130 1118 1136 1119
rect 1150 1118 1156 1119
rect 1162 1118 1168 1119
rect 1214 1118 1220 1119
rect 478 1107 484 1108
rect 478 1103 479 1107
rect 483 1103 484 1107
rect 478 1102 484 1103
rect 902 1107 908 1108
rect 902 1103 903 1107
rect 907 1103 908 1107
rect 902 1102 908 1103
rect 1042 1107 1048 1108
rect 1042 1103 1043 1107
rect 1047 1103 1048 1107
rect 1042 1102 1048 1103
rect 1102 1107 1108 1108
rect 1102 1103 1103 1107
rect 1107 1103 1108 1107
rect 1102 1102 1108 1103
rect 334 1101 340 1102
rect 334 1097 335 1101
rect 339 1097 340 1101
rect 334 1096 340 1097
rect 398 1101 404 1102
rect 398 1097 399 1101
rect 403 1097 404 1101
rect 398 1096 404 1097
rect 462 1101 468 1102
rect 462 1097 463 1101
rect 467 1097 468 1101
rect 462 1096 468 1097
rect 526 1101 532 1102
rect 526 1097 527 1101
rect 531 1097 532 1101
rect 526 1096 532 1097
rect 598 1101 604 1102
rect 598 1097 599 1101
rect 603 1097 604 1101
rect 598 1096 604 1097
rect 662 1101 668 1102
rect 662 1097 663 1101
rect 667 1097 668 1101
rect 662 1096 668 1097
rect 726 1101 732 1102
rect 726 1097 727 1101
rect 731 1097 732 1101
rect 726 1096 732 1097
rect 790 1101 796 1102
rect 790 1097 791 1101
rect 795 1097 796 1101
rect 790 1096 796 1097
rect 854 1101 860 1102
rect 854 1097 855 1101
rect 859 1097 860 1101
rect 854 1096 860 1097
rect 336 1091 338 1096
rect 400 1091 402 1096
rect 464 1091 466 1096
rect 528 1091 530 1096
rect 600 1091 602 1096
rect 664 1091 666 1096
rect 728 1091 730 1096
rect 792 1091 794 1096
rect 856 1091 858 1096
rect 311 1090 315 1091
rect 311 1084 315 1086
rect 335 1090 339 1091
rect 335 1085 339 1086
rect 351 1090 355 1091
rect 351 1084 355 1086
rect 391 1090 395 1091
rect 391 1084 395 1086
rect 399 1090 403 1091
rect 399 1085 403 1086
rect 439 1090 443 1091
rect 439 1084 443 1086
rect 463 1090 467 1091
rect 463 1085 467 1086
rect 503 1090 507 1091
rect 503 1084 507 1086
rect 527 1090 531 1091
rect 527 1085 531 1086
rect 575 1090 579 1091
rect 575 1084 579 1086
rect 599 1090 603 1091
rect 599 1085 603 1086
rect 655 1090 659 1091
rect 655 1084 659 1086
rect 663 1090 667 1091
rect 663 1085 667 1086
rect 727 1090 731 1091
rect 727 1085 731 1086
rect 735 1090 739 1091
rect 735 1084 739 1086
rect 791 1090 795 1091
rect 791 1085 795 1086
rect 815 1090 819 1091
rect 815 1084 819 1086
rect 855 1090 859 1091
rect 855 1085 859 1086
rect 895 1090 899 1091
rect 895 1084 899 1086
rect 310 1083 316 1084
rect 310 1079 311 1083
rect 315 1079 316 1083
rect 310 1078 316 1079
rect 350 1083 356 1084
rect 350 1079 351 1083
rect 355 1079 356 1083
rect 350 1078 356 1079
rect 390 1083 396 1084
rect 390 1079 391 1083
rect 395 1079 396 1083
rect 390 1078 396 1079
rect 438 1083 444 1084
rect 438 1079 439 1083
rect 443 1079 444 1083
rect 438 1078 444 1079
rect 502 1083 508 1084
rect 502 1079 503 1083
rect 507 1079 508 1083
rect 502 1078 508 1079
rect 574 1083 580 1084
rect 574 1079 575 1083
rect 579 1079 580 1083
rect 574 1078 580 1079
rect 654 1083 660 1084
rect 654 1079 655 1083
rect 659 1079 660 1083
rect 654 1078 660 1079
rect 734 1083 740 1084
rect 734 1079 735 1083
rect 739 1079 740 1083
rect 734 1078 740 1079
rect 814 1083 820 1084
rect 814 1079 815 1083
rect 819 1079 820 1083
rect 814 1078 820 1079
rect 894 1083 900 1084
rect 894 1079 895 1083
rect 899 1079 900 1083
rect 894 1078 900 1079
rect 298 1075 304 1076
rect 298 1071 299 1075
rect 303 1071 304 1075
rect 298 1070 304 1071
rect 666 1075 672 1076
rect 666 1071 667 1075
rect 671 1071 672 1075
rect 666 1070 672 1071
rect 806 1075 812 1076
rect 806 1071 807 1075
rect 811 1071 812 1075
rect 806 1070 812 1071
rect 246 1066 252 1067
rect 246 1062 247 1066
rect 251 1062 252 1066
rect 246 1061 252 1062
rect 278 1066 284 1067
rect 278 1062 279 1066
rect 283 1062 284 1066
rect 278 1061 284 1062
rect 310 1066 316 1067
rect 310 1062 311 1066
rect 315 1062 316 1066
rect 310 1061 316 1062
rect 350 1066 356 1067
rect 350 1062 351 1066
rect 355 1062 356 1066
rect 350 1061 356 1062
rect 390 1066 396 1067
rect 390 1062 391 1066
rect 395 1062 396 1066
rect 390 1061 396 1062
rect 438 1066 444 1067
rect 438 1062 439 1066
rect 443 1062 444 1066
rect 438 1061 444 1062
rect 502 1066 508 1067
rect 502 1062 503 1066
rect 507 1062 508 1066
rect 502 1061 508 1062
rect 574 1066 580 1067
rect 574 1062 575 1066
rect 579 1062 580 1066
rect 574 1061 580 1062
rect 654 1066 660 1067
rect 654 1062 655 1066
rect 659 1062 660 1066
rect 654 1061 660 1062
rect 234 1059 240 1060
rect 234 1055 235 1059
rect 239 1055 240 1059
rect 234 1054 240 1055
rect 248 1047 250 1061
rect 280 1047 282 1061
rect 312 1047 314 1061
rect 352 1047 354 1061
rect 392 1047 394 1061
rect 440 1047 442 1061
rect 470 1051 476 1052
rect 470 1047 471 1051
rect 475 1047 476 1051
rect 504 1047 506 1061
rect 576 1047 578 1061
rect 656 1047 658 1061
rect 668 1048 670 1070
rect 734 1066 740 1067
rect 734 1062 735 1066
rect 739 1062 740 1066
rect 734 1061 740 1062
rect 666 1047 672 1048
rect 736 1047 738 1061
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 215 1046 219 1047
rect 215 1041 219 1042
rect 247 1046 251 1047
rect 247 1041 251 1042
rect 279 1046 283 1047
rect 279 1041 283 1042
rect 295 1046 299 1047
rect 295 1041 299 1042
rect 311 1046 315 1047
rect 311 1041 315 1042
rect 327 1046 331 1047
rect 327 1041 331 1042
rect 351 1046 355 1047
rect 351 1041 355 1042
rect 359 1046 363 1047
rect 359 1041 363 1042
rect 391 1046 395 1047
rect 391 1041 395 1042
rect 423 1046 427 1047
rect 423 1041 427 1042
rect 439 1046 443 1047
rect 439 1041 443 1042
rect 455 1046 459 1047
rect 470 1046 476 1047
rect 503 1046 507 1047
rect 455 1041 459 1042
rect 112 1033 114 1041
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 296 1031 298 1041
rect 302 1035 308 1036
rect 302 1031 303 1035
rect 307 1031 308 1035
rect 328 1031 330 1041
rect 360 1031 362 1041
rect 392 1031 394 1041
rect 424 1031 426 1041
rect 456 1031 458 1041
rect 110 1027 116 1028
rect 294 1030 300 1031
rect 302 1030 308 1031
rect 326 1030 332 1031
rect 294 1026 295 1030
rect 299 1026 300 1030
rect 294 1025 300 1026
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 110 1010 116 1011
rect 294 1013 300 1014
rect 112 1007 114 1010
rect 294 1009 295 1013
rect 299 1009 300 1013
rect 294 1008 300 1009
rect 304 1008 306 1030
rect 326 1026 327 1030
rect 331 1026 332 1030
rect 326 1025 332 1026
rect 358 1030 364 1031
rect 358 1026 359 1030
rect 363 1026 364 1030
rect 358 1025 364 1026
rect 390 1030 396 1031
rect 390 1026 391 1030
rect 395 1026 396 1030
rect 390 1025 396 1026
rect 422 1030 428 1031
rect 422 1026 423 1030
rect 427 1026 428 1030
rect 422 1025 428 1026
rect 454 1030 460 1031
rect 454 1026 455 1030
rect 459 1026 460 1030
rect 454 1025 460 1026
rect 472 1020 474 1046
rect 503 1041 507 1042
rect 559 1046 563 1047
rect 559 1041 563 1042
rect 575 1046 579 1047
rect 575 1041 579 1042
rect 631 1046 635 1047
rect 631 1041 635 1042
rect 655 1046 659 1047
rect 666 1043 667 1047
rect 671 1043 672 1047
rect 666 1042 672 1043
rect 711 1046 715 1047
rect 655 1041 659 1042
rect 711 1041 715 1042
rect 735 1046 739 1047
rect 735 1041 739 1042
rect 799 1046 803 1047
rect 799 1041 803 1042
rect 504 1031 506 1041
rect 560 1031 562 1041
rect 632 1031 634 1041
rect 712 1031 714 1041
rect 800 1031 802 1041
rect 808 1036 810 1070
rect 814 1066 820 1067
rect 814 1062 815 1066
rect 819 1062 820 1066
rect 814 1061 820 1062
rect 894 1066 900 1067
rect 894 1062 895 1066
rect 899 1062 900 1066
rect 894 1061 900 1062
rect 816 1047 818 1061
rect 896 1047 898 1061
rect 904 1060 906 1102
rect 910 1101 916 1102
rect 910 1097 911 1101
rect 915 1097 916 1101
rect 910 1096 916 1097
rect 966 1101 972 1102
rect 966 1097 967 1101
rect 971 1097 972 1101
rect 966 1096 972 1097
rect 1022 1101 1028 1102
rect 1022 1097 1023 1101
rect 1027 1097 1028 1101
rect 1022 1096 1028 1097
rect 1086 1101 1092 1102
rect 1086 1097 1087 1101
rect 1091 1097 1092 1101
rect 1086 1096 1092 1097
rect 1132 1096 1134 1118
rect 1150 1114 1151 1118
rect 1155 1114 1156 1118
rect 1150 1113 1156 1114
rect 1150 1101 1156 1102
rect 1150 1097 1151 1101
rect 1155 1097 1156 1101
rect 1150 1096 1156 1097
rect 912 1091 914 1096
rect 968 1091 970 1096
rect 1024 1091 1026 1096
rect 1088 1091 1090 1096
rect 1130 1095 1136 1096
rect 1130 1091 1131 1095
rect 1135 1091 1136 1095
rect 1152 1091 1154 1096
rect 911 1090 915 1091
rect 911 1085 915 1086
rect 967 1090 971 1091
rect 967 1084 971 1086
rect 1023 1090 1027 1091
rect 1023 1085 1027 1086
rect 1039 1090 1043 1091
rect 1039 1084 1043 1086
rect 1087 1090 1091 1091
rect 1087 1085 1091 1086
rect 1111 1090 1115 1091
rect 1130 1090 1136 1091
rect 1151 1090 1155 1091
rect 1111 1084 1115 1086
rect 1151 1085 1155 1086
rect 966 1083 972 1084
rect 966 1079 967 1083
rect 971 1079 972 1083
rect 966 1078 972 1079
rect 1038 1083 1044 1084
rect 1038 1079 1039 1083
rect 1043 1079 1044 1083
rect 1038 1078 1044 1079
rect 1110 1083 1116 1084
rect 1110 1079 1111 1083
rect 1115 1079 1116 1083
rect 1110 1078 1116 1079
rect 1164 1076 1166 1118
rect 1214 1114 1215 1118
rect 1219 1114 1220 1118
rect 1214 1113 1220 1114
rect 1278 1118 1284 1119
rect 1278 1114 1279 1118
rect 1283 1114 1284 1118
rect 1278 1113 1284 1114
rect 1334 1118 1340 1119
rect 1334 1114 1335 1118
rect 1339 1114 1340 1118
rect 1334 1113 1340 1114
rect 1390 1118 1396 1119
rect 1390 1114 1391 1118
rect 1395 1114 1396 1118
rect 1390 1113 1396 1114
rect 1446 1118 1452 1119
rect 1446 1114 1447 1118
rect 1451 1114 1452 1118
rect 1446 1113 1452 1114
rect 1494 1118 1500 1119
rect 1494 1114 1495 1118
rect 1499 1114 1500 1118
rect 1494 1113 1500 1114
rect 1542 1118 1548 1119
rect 1558 1118 1564 1119
rect 1590 1118 1596 1119
rect 1542 1114 1543 1118
rect 1547 1114 1548 1118
rect 1542 1113 1548 1114
rect 1214 1101 1220 1102
rect 1214 1097 1215 1101
rect 1219 1097 1220 1101
rect 1214 1096 1220 1097
rect 1278 1101 1284 1102
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1278 1096 1284 1097
rect 1334 1101 1340 1102
rect 1334 1097 1335 1101
rect 1339 1097 1340 1101
rect 1334 1096 1340 1097
rect 1390 1101 1396 1102
rect 1390 1097 1391 1101
rect 1395 1097 1396 1101
rect 1390 1096 1396 1097
rect 1446 1101 1452 1102
rect 1446 1097 1447 1101
rect 1451 1097 1452 1101
rect 1446 1096 1452 1097
rect 1494 1101 1500 1102
rect 1494 1097 1495 1101
rect 1499 1097 1500 1101
rect 1494 1096 1500 1097
rect 1542 1101 1548 1102
rect 1542 1097 1543 1101
rect 1547 1097 1548 1101
rect 1542 1096 1548 1097
rect 1216 1091 1218 1096
rect 1280 1091 1282 1096
rect 1336 1091 1338 1096
rect 1378 1095 1384 1096
rect 1378 1091 1379 1095
rect 1383 1091 1384 1095
rect 1392 1091 1394 1096
rect 1448 1091 1450 1096
rect 1496 1091 1498 1096
rect 1544 1091 1546 1096
rect 1560 1092 1562 1118
rect 1590 1114 1591 1118
rect 1595 1114 1596 1118
rect 1590 1113 1596 1114
rect 1622 1118 1628 1119
rect 1622 1114 1623 1118
rect 1627 1114 1628 1118
rect 1662 1116 1663 1120
rect 1667 1116 1668 1120
rect 1662 1115 1668 1116
rect 1622 1113 1628 1114
rect 1638 1107 1644 1108
rect 1638 1103 1639 1107
rect 1643 1103 1644 1107
rect 1638 1102 1644 1103
rect 1662 1103 1668 1104
rect 1590 1101 1596 1102
rect 1590 1097 1591 1101
rect 1595 1097 1596 1101
rect 1590 1096 1596 1097
rect 1622 1101 1628 1102
rect 1622 1097 1623 1101
rect 1627 1097 1628 1101
rect 1622 1096 1628 1097
rect 1558 1091 1564 1092
rect 1592 1091 1594 1096
rect 1624 1091 1626 1096
rect 1175 1090 1179 1091
rect 1175 1084 1179 1086
rect 1215 1090 1219 1091
rect 1215 1085 1219 1086
rect 1239 1090 1243 1091
rect 1239 1084 1243 1086
rect 1279 1090 1283 1091
rect 1279 1085 1283 1086
rect 1303 1090 1307 1091
rect 1303 1084 1307 1086
rect 1335 1090 1339 1091
rect 1335 1085 1339 1086
rect 1359 1090 1363 1091
rect 1378 1090 1384 1091
rect 1391 1090 1395 1091
rect 1359 1084 1363 1086
rect 1174 1083 1180 1084
rect 1174 1079 1175 1083
rect 1179 1079 1180 1083
rect 1174 1078 1180 1079
rect 1238 1083 1244 1084
rect 1238 1079 1239 1083
rect 1243 1079 1244 1083
rect 1238 1078 1244 1079
rect 1302 1083 1308 1084
rect 1302 1079 1303 1083
rect 1307 1079 1308 1083
rect 1302 1078 1308 1079
rect 1358 1083 1364 1084
rect 1358 1079 1359 1083
rect 1363 1079 1364 1083
rect 1358 1078 1364 1079
rect 1162 1075 1168 1076
rect 1162 1071 1163 1075
rect 1167 1071 1168 1075
rect 1162 1070 1168 1071
rect 1186 1075 1192 1076
rect 1186 1071 1187 1075
rect 1191 1071 1192 1075
rect 1186 1070 1192 1071
rect 966 1066 972 1067
rect 966 1062 967 1066
rect 971 1062 972 1066
rect 966 1061 972 1062
rect 1038 1066 1044 1067
rect 1038 1062 1039 1066
rect 1043 1062 1044 1066
rect 1038 1061 1044 1062
rect 1110 1066 1116 1067
rect 1110 1062 1111 1066
rect 1115 1062 1116 1066
rect 1110 1061 1116 1062
rect 1174 1066 1180 1067
rect 1174 1062 1175 1066
rect 1179 1062 1180 1066
rect 1174 1061 1180 1062
rect 902 1059 908 1060
rect 902 1055 903 1059
rect 907 1055 908 1059
rect 902 1054 908 1055
rect 968 1047 970 1061
rect 1040 1047 1042 1061
rect 1112 1047 1114 1061
rect 1176 1047 1178 1061
rect 1188 1052 1190 1070
rect 1238 1066 1244 1067
rect 1238 1062 1239 1066
rect 1243 1062 1244 1066
rect 1238 1061 1244 1062
rect 1302 1066 1308 1067
rect 1302 1062 1303 1066
rect 1307 1062 1308 1066
rect 1302 1061 1308 1062
rect 1358 1066 1364 1067
rect 1358 1062 1359 1066
rect 1363 1062 1364 1066
rect 1358 1061 1364 1062
rect 1186 1051 1192 1052
rect 1186 1047 1187 1051
rect 1191 1047 1192 1051
rect 1240 1047 1242 1061
rect 1304 1047 1306 1061
rect 1310 1059 1316 1060
rect 1310 1055 1311 1059
rect 1315 1055 1316 1059
rect 1310 1054 1316 1055
rect 815 1046 819 1047
rect 815 1041 819 1042
rect 879 1046 883 1047
rect 879 1041 883 1042
rect 895 1046 899 1047
rect 895 1041 899 1042
rect 959 1046 963 1047
rect 959 1041 963 1042
rect 967 1046 971 1047
rect 967 1041 971 1042
rect 1031 1046 1035 1047
rect 1031 1041 1035 1042
rect 1039 1046 1043 1047
rect 1039 1041 1043 1042
rect 1095 1046 1099 1047
rect 1095 1041 1099 1042
rect 1111 1046 1115 1047
rect 1111 1041 1115 1042
rect 1159 1046 1163 1047
rect 1159 1041 1163 1042
rect 1175 1046 1179 1047
rect 1186 1046 1192 1047
rect 1223 1046 1227 1047
rect 1175 1041 1179 1042
rect 1223 1041 1227 1042
rect 1239 1046 1243 1047
rect 1239 1041 1243 1042
rect 1279 1046 1283 1047
rect 1279 1041 1283 1042
rect 1303 1046 1307 1047
rect 1303 1041 1307 1042
rect 806 1035 812 1036
rect 806 1031 807 1035
rect 811 1031 812 1035
rect 880 1031 882 1041
rect 960 1031 962 1041
rect 974 1035 980 1036
rect 974 1031 975 1035
rect 979 1031 980 1035
rect 1032 1031 1034 1041
rect 1096 1031 1098 1041
rect 1160 1031 1162 1041
rect 1224 1031 1226 1041
rect 1280 1031 1282 1041
rect 502 1030 508 1031
rect 502 1026 503 1030
rect 507 1026 508 1030
rect 502 1025 508 1026
rect 558 1030 564 1031
rect 558 1026 559 1030
rect 563 1026 564 1030
rect 558 1025 564 1026
rect 630 1030 636 1031
rect 630 1026 631 1030
rect 635 1026 636 1030
rect 630 1025 636 1026
rect 710 1030 716 1031
rect 710 1026 711 1030
rect 715 1026 716 1030
rect 710 1025 716 1026
rect 798 1030 804 1031
rect 806 1030 812 1031
rect 878 1030 884 1031
rect 798 1026 799 1030
rect 803 1026 804 1030
rect 798 1025 804 1026
rect 878 1026 879 1030
rect 883 1026 884 1030
rect 878 1025 884 1026
rect 958 1030 964 1031
rect 974 1030 980 1031
rect 1030 1030 1036 1031
rect 958 1026 959 1030
rect 963 1026 964 1030
rect 958 1025 964 1026
rect 470 1019 476 1020
rect 470 1015 471 1019
rect 475 1015 476 1019
rect 470 1014 476 1015
rect 890 1019 896 1020
rect 890 1015 891 1019
rect 895 1015 896 1019
rect 890 1014 896 1015
rect 326 1013 332 1014
rect 326 1009 327 1013
rect 331 1009 332 1013
rect 326 1008 332 1009
rect 358 1013 364 1014
rect 358 1009 359 1013
rect 363 1009 364 1013
rect 358 1008 364 1009
rect 390 1013 396 1014
rect 390 1009 391 1013
rect 395 1009 396 1013
rect 390 1008 396 1009
rect 422 1013 428 1014
rect 422 1009 423 1013
rect 427 1009 428 1013
rect 422 1008 428 1009
rect 454 1013 460 1014
rect 454 1009 455 1013
rect 459 1009 460 1013
rect 454 1008 460 1009
rect 502 1013 508 1014
rect 502 1009 503 1013
rect 507 1009 508 1013
rect 502 1008 508 1009
rect 558 1013 564 1014
rect 558 1009 559 1013
rect 563 1009 564 1013
rect 558 1008 564 1009
rect 630 1013 636 1014
rect 630 1009 631 1013
rect 635 1009 636 1013
rect 630 1008 636 1009
rect 710 1013 716 1014
rect 710 1009 711 1013
rect 715 1009 716 1013
rect 710 1008 716 1009
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 878 1013 884 1014
rect 878 1009 879 1013
rect 883 1009 884 1013
rect 878 1008 884 1009
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 247 1006 251 1007
rect 112 998 114 1001
rect 247 1000 251 1002
rect 279 1006 283 1007
rect 279 1000 283 1002
rect 295 1006 299 1008
rect 302 1007 308 1008
rect 302 1003 303 1007
rect 307 1003 308 1007
rect 302 1002 308 1003
rect 311 1006 315 1007
rect 295 1001 299 1002
rect 311 1000 315 1002
rect 327 1006 331 1008
rect 327 1001 331 1002
rect 343 1006 347 1007
rect 343 1000 347 1002
rect 359 1006 363 1008
rect 359 1001 363 1002
rect 383 1006 387 1007
rect 383 1000 387 1002
rect 391 1006 395 1008
rect 391 1001 395 1002
rect 423 1006 427 1008
rect 423 1000 427 1002
rect 455 1006 459 1008
rect 455 1001 459 1002
rect 479 1006 483 1007
rect 479 1000 483 1002
rect 503 1006 507 1008
rect 510 1007 516 1008
rect 510 1003 511 1007
rect 515 1003 516 1007
rect 510 1002 516 1003
rect 543 1006 547 1007
rect 503 1001 507 1002
rect 246 999 252 1000
rect 110 997 116 998
rect 110 993 111 997
rect 115 993 116 997
rect 246 995 247 999
rect 251 995 252 999
rect 246 994 252 995
rect 278 999 284 1000
rect 278 995 279 999
rect 283 995 284 999
rect 278 994 284 995
rect 310 999 316 1000
rect 310 995 311 999
rect 315 995 316 999
rect 310 994 316 995
rect 342 999 348 1000
rect 342 995 343 999
rect 347 995 348 999
rect 342 994 348 995
rect 382 999 388 1000
rect 382 995 383 999
rect 387 995 388 999
rect 382 994 388 995
rect 422 999 428 1000
rect 422 995 423 999
rect 427 995 428 999
rect 422 994 428 995
rect 478 999 484 1000
rect 478 995 479 999
rect 483 995 484 999
rect 478 994 484 995
rect 110 992 116 993
rect 246 982 252 983
rect 110 980 116 981
rect 110 976 111 980
rect 115 976 116 980
rect 246 978 247 982
rect 251 978 252 982
rect 246 977 252 978
rect 278 982 284 983
rect 278 978 279 982
rect 283 978 284 982
rect 278 977 284 978
rect 310 982 316 983
rect 310 978 311 982
rect 315 978 316 982
rect 310 977 316 978
rect 342 982 348 983
rect 342 978 343 982
rect 347 978 348 982
rect 342 977 348 978
rect 382 982 388 983
rect 382 978 383 982
rect 387 978 388 982
rect 382 977 388 978
rect 422 982 428 983
rect 422 978 423 982
rect 427 978 428 982
rect 422 977 428 978
rect 478 982 484 983
rect 478 978 479 982
rect 483 978 484 982
rect 478 977 484 978
rect 110 975 116 976
rect 112 967 114 975
rect 248 967 250 977
rect 280 967 282 977
rect 312 967 314 977
rect 344 967 346 977
rect 384 967 386 977
rect 414 967 420 968
rect 424 967 426 977
rect 480 967 482 977
rect 512 976 514 1002
rect 543 1000 547 1002
rect 559 1006 563 1008
rect 559 1001 563 1002
rect 615 1006 619 1007
rect 615 1000 619 1002
rect 631 1006 635 1008
rect 631 1001 635 1002
rect 687 1006 691 1007
rect 687 1000 691 1002
rect 711 1006 715 1008
rect 711 1001 715 1002
rect 759 1006 763 1007
rect 759 1000 763 1002
rect 799 1006 803 1008
rect 799 1001 803 1002
rect 831 1006 835 1007
rect 831 1000 835 1002
rect 879 1006 883 1008
rect 879 1001 883 1002
rect 542 999 548 1000
rect 542 995 543 999
rect 547 995 548 999
rect 542 994 548 995
rect 614 999 620 1000
rect 614 995 615 999
rect 619 995 620 999
rect 614 994 620 995
rect 686 999 692 1000
rect 686 995 687 999
rect 691 995 692 999
rect 686 994 692 995
rect 758 999 764 1000
rect 758 995 759 999
rect 763 995 764 999
rect 758 994 764 995
rect 830 999 836 1000
rect 830 995 831 999
rect 835 995 836 999
rect 830 994 836 995
rect 674 991 680 992
rect 674 987 675 991
rect 679 987 680 991
rect 674 986 680 987
rect 806 991 812 992
rect 806 987 807 991
rect 811 987 812 991
rect 806 986 812 987
rect 542 982 548 983
rect 542 978 543 982
rect 547 978 548 982
rect 542 977 548 978
rect 614 982 620 983
rect 614 978 615 982
rect 619 978 620 982
rect 614 977 620 978
rect 510 975 516 976
rect 510 971 511 975
rect 515 971 516 975
rect 510 970 516 971
rect 544 967 546 977
rect 616 967 618 977
rect 676 968 678 986
rect 686 982 692 983
rect 686 978 687 982
rect 691 978 692 982
rect 686 977 692 978
rect 758 982 764 983
rect 758 978 759 982
rect 763 978 764 982
rect 758 977 764 978
rect 674 967 680 968
rect 688 967 690 977
rect 760 967 762 977
rect 111 966 115 967
rect 111 961 115 962
rect 167 966 171 967
rect 167 961 171 962
rect 199 966 203 967
rect 199 961 203 962
rect 239 966 243 967
rect 239 961 243 962
rect 247 966 251 967
rect 247 961 251 962
rect 279 966 283 967
rect 279 961 283 962
rect 287 966 291 967
rect 287 961 291 962
rect 311 966 315 967
rect 311 961 315 962
rect 343 966 347 967
rect 343 961 347 962
rect 383 966 387 967
rect 383 961 387 962
rect 407 966 411 967
rect 414 963 415 967
rect 419 963 420 967
rect 414 962 420 963
rect 423 966 427 967
rect 407 961 411 962
rect 112 953 114 961
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 168 951 170 961
rect 186 955 192 956
rect 186 951 187 955
rect 191 951 192 955
rect 200 951 202 961
rect 240 951 242 961
rect 288 951 290 961
rect 344 951 346 961
rect 408 951 410 961
rect 110 947 116 948
rect 166 950 172 951
rect 186 950 192 951
rect 198 950 204 951
rect 166 946 167 950
rect 171 946 172 950
rect 166 945 172 946
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 110 930 116 931
rect 166 933 172 934
rect 112 923 114 930
rect 166 929 167 933
rect 171 929 172 933
rect 166 928 172 929
rect 168 923 170 928
rect 188 924 190 950
rect 198 946 199 950
rect 203 946 204 950
rect 198 945 204 946
rect 238 950 244 951
rect 238 946 239 950
rect 243 946 244 950
rect 238 945 244 946
rect 286 950 292 951
rect 286 946 287 950
rect 291 946 292 950
rect 286 945 292 946
rect 342 950 348 951
rect 342 946 343 950
rect 347 946 348 950
rect 342 945 348 946
rect 406 950 412 951
rect 406 946 407 950
rect 411 946 412 950
rect 406 945 412 946
rect 416 940 418 962
rect 423 961 427 962
rect 471 966 475 967
rect 471 961 475 962
rect 479 966 483 967
rect 479 961 483 962
rect 535 966 539 967
rect 535 961 539 962
rect 543 966 547 967
rect 543 961 547 962
rect 599 966 603 967
rect 599 961 603 962
rect 615 966 619 967
rect 615 961 619 962
rect 663 966 667 967
rect 674 963 675 967
rect 679 963 680 967
rect 674 962 680 963
rect 687 966 691 967
rect 663 961 667 962
rect 687 961 691 962
rect 727 966 731 967
rect 727 961 731 962
rect 759 966 763 967
rect 759 961 763 962
rect 791 966 795 967
rect 791 961 795 962
rect 472 951 474 961
rect 536 951 538 961
rect 600 951 602 961
rect 664 951 666 961
rect 728 951 730 961
rect 792 951 794 961
rect 808 956 810 986
rect 830 982 836 983
rect 830 978 831 982
rect 835 978 836 982
rect 830 977 836 978
rect 832 967 834 977
rect 892 976 894 1014
rect 958 1013 964 1014
rect 958 1009 959 1013
rect 963 1009 964 1013
rect 958 1008 964 1009
rect 976 1008 978 1030
rect 1030 1026 1031 1030
rect 1035 1026 1036 1030
rect 1030 1025 1036 1026
rect 1094 1030 1100 1031
rect 1094 1026 1095 1030
rect 1099 1026 1100 1030
rect 1094 1025 1100 1026
rect 1158 1030 1164 1031
rect 1158 1026 1159 1030
rect 1163 1026 1164 1030
rect 1158 1025 1164 1026
rect 1222 1030 1228 1031
rect 1222 1026 1223 1030
rect 1227 1026 1228 1030
rect 1222 1025 1228 1026
rect 1278 1030 1284 1031
rect 1278 1026 1279 1030
rect 1283 1026 1284 1030
rect 1278 1025 1284 1026
rect 1312 1020 1314 1054
rect 1360 1047 1362 1061
rect 1380 1060 1382 1090
rect 1391 1085 1395 1086
rect 1415 1090 1419 1091
rect 1415 1084 1419 1086
rect 1447 1090 1451 1091
rect 1447 1085 1451 1086
rect 1463 1090 1467 1091
rect 1463 1084 1467 1086
rect 1495 1090 1499 1091
rect 1495 1085 1499 1086
rect 1503 1090 1507 1091
rect 1503 1084 1507 1086
rect 1543 1090 1547 1091
rect 1543 1085 1547 1086
rect 1551 1090 1555 1091
rect 1558 1087 1559 1091
rect 1563 1087 1564 1091
rect 1558 1086 1564 1087
rect 1591 1090 1595 1091
rect 1551 1084 1555 1086
rect 1591 1084 1595 1086
rect 1623 1090 1627 1091
rect 1623 1084 1627 1086
rect 1414 1083 1420 1084
rect 1414 1079 1415 1083
rect 1419 1079 1420 1083
rect 1414 1078 1420 1079
rect 1462 1083 1468 1084
rect 1462 1079 1463 1083
rect 1467 1079 1468 1083
rect 1462 1078 1468 1079
rect 1502 1083 1508 1084
rect 1502 1079 1503 1083
rect 1507 1079 1508 1083
rect 1502 1078 1508 1079
rect 1550 1083 1556 1084
rect 1550 1079 1551 1083
rect 1555 1079 1556 1083
rect 1550 1078 1556 1079
rect 1590 1083 1596 1084
rect 1590 1079 1591 1083
rect 1595 1079 1596 1083
rect 1590 1078 1596 1079
rect 1622 1083 1628 1084
rect 1622 1079 1623 1083
rect 1627 1079 1628 1083
rect 1622 1078 1628 1079
rect 1606 1067 1612 1068
rect 1414 1066 1420 1067
rect 1414 1062 1415 1066
rect 1419 1062 1420 1066
rect 1414 1061 1420 1062
rect 1462 1066 1468 1067
rect 1462 1062 1463 1066
rect 1467 1062 1468 1066
rect 1462 1061 1468 1062
rect 1502 1066 1508 1067
rect 1502 1062 1503 1066
rect 1507 1062 1508 1066
rect 1502 1061 1508 1062
rect 1550 1066 1556 1067
rect 1550 1062 1551 1066
rect 1555 1062 1556 1066
rect 1550 1061 1556 1062
rect 1590 1066 1596 1067
rect 1590 1062 1591 1066
rect 1595 1062 1596 1066
rect 1606 1063 1607 1067
rect 1611 1063 1612 1067
rect 1606 1062 1612 1063
rect 1622 1066 1628 1067
rect 1622 1062 1623 1066
rect 1627 1062 1628 1066
rect 1590 1061 1596 1062
rect 1378 1059 1384 1060
rect 1378 1055 1379 1059
rect 1383 1055 1384 1059
rect 1378 1054 1384 1055
rect 1416 1047 1418 1061
rect 1446 1047 1452 1048
rect 1464 1047 1466 1061
rect 1504 1047 1506 1061
rect 1552 1047 1554 1061
rect 1592 1047 1594 1061
rect 1335 1046 1339 1047
rect 1335 1041 1339 1042
rect 1359 1046 1363 1047
rect 1359 1041 1363 1042
rect 1383 1046 1387 1047
rect 1383 1041 1387 1042
rect 1415 1046 1419 1047
rect 1415 1041 1419 1042
rect 1431 1046 1435 1047
rect 1446 1043 1447 1047
rect 1451 1043 1452 1047
rect 1446 1042 1452 1043
rect 1463 1046 1467 1047
rect 1431 1041 1435 1042
rect 1336 1031 1338 1041
rect 1384 1031 1386 1041
rect 1432 1031 1434 1041
rect 1334 1030 1340 1031
rect 1334 1026 1335 1030
rect 1339 1026 1340 1030
rect 1334 1025 1340 1026
rect 1382 1030 1388 1031
rect 1382 1026 1383 1030
rect 1387 1026 1388 1030
rect 1382 1025 1388 1026
rect 1430 1030 1436 1031
rect 1430 1026 1431 1030
rect 1435 1026 1436 1030
rect 1430 1025 1436 1026
rect 1448 1020 1450 1042
rect 1463 1041 1467 1042
rect 1479 1046 1483 1047
rect 1479 1041 1483 1042
rect 1503 1046 1507 1047
rect 1503 1041 1507 1042
rect 1535 1046 1539 1047
rect 1535 1041 1539 1042
rect 1551 1046 1555 1047
rect 1551 1041 1555 1042
rect 1591 1046 1595 1047
rect 1591 1041 1595 1042
rect 1480 1031 1482 1041
rect 1536 1031 1538 1041
rect 1554 1035 1560 1036
rect 1554 1031 1555 1035
rect 1559 1031 1560 1035
rect 1592 1031 1594 1041
rect 1608 1036 1610 1062
rect 1622 1061 1628 1062
rect 1624 1047 1626 1061
rect 1640 1060 1642 1102
rect 1662 1099 1663 1103
rect 1667 1099 1668 1103
rect 1662 1098 1668 1099
rect 1664 1091 1666 1098
rect 1663 1090 1667 1091
rect 1663 1085 1667 1086
rect 1664 1082 1666 1085
rect 1662 1081 1668 1082
rect 1662 1077 1663 1081
rect 1667 1077 1668 1081
rect 1662 1076 1668 1077
rect 1662 1064 1668 1065
rect 1662 1060 1663 1064
rect 1667 1060 1668 1064
rect 1638 1059 1644 1060
rect 1662 1059 1668 1060
rect 1638 1055 1639 1059
rect 1643 1055 1644 1059
rect 1638 1054 1644 1055
rect 1664 1047 1666 1059
rect 1623 1046 1627 1047
rect 1623 1041 1627 1042
rect 1663 1046 1667 1047
rect 1663 1041 1667 1042
rect 1606 1035 1612 1036
rect 1606 1031 1607 1035
rect 1611 1031 1612 1035
rect 1624 1031 1626 1041
rect 1664 1033 1666 1041
rect 1662 1032 1668 1033
rect 1478 1030 1484 1031
rect 1478 1026 1479 1030
rect 1483 1026 1484 1030
rect 1478 1025 1484 1026
rect 1534 1030 1540 1031
rect 1554 1030 1560 1031
rect 1590 1030 1596 1031
rect 1606 1030 1612 1031
rect 1622 1030 1628 1031
rect 1534 1026 1535 1030
rect 1539 1026 1540 1030
rect 1534 1025 1540 1026
rect 1310 1019 1316 1020
rect 1310 1015 1311 1019
rect 1315 1015 1316 1019
rect 1310 1014 1316 1015
rect 1414 1019 1420 1020
rect 1414 1015 1415 1019
rect 1419 1015 1420 1019
rect 1414 1014 1420 1015
rect 1446 1019 1452 1020
rect 1446 1015 1447 1019
rect 1451 1015 1452 1019
rect 1446 1014 1452 1015
rect 1030 1013 1036 1014
rect 1030 1009 1031 1013
rect 1035 1009 1036 1013
rect 1030 1008 1036 1009
rect 1094 1013 1100 1014
rect 1094 1009 1095 1013
rect 1099 1009 1100 1013
rect 1094 1008 1100 1009
rect 1158 1013 1164 1014
rect 1158 1009 1159 1013
rect 1163 1009 1164 1013
rect 1158 1008 1164 1009
rect 1222 1013 1228 1014
rect 1222 1009 1223 1013
rect 1227 1009 1228 1013
rect 1222 1008 1228 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 1334 1013 1340 1014
rect 1334 1009 1335 1013
rect 1339 1009 1340 1013
rect 1334 1008 1340 1009
rect 1382 1013 1388 1014
rect 1382 1009 1383 1013
rect 1387 1009 1388 1013
rect 1382 1008 1388 1009
rect 903 1006 907 1007
rect 903 1000 907 1002
rect 959 1006 963 1008
rect 974 1007 980 1008
rect 959 1001 963 1002
rect 967 1006 971 1007
rect 974 1003 975 1007
rect 979 1003 980 1007
rect 974 1002 980 1003
rect 1031 1006 1035 1008
rect 967 1000 971 1002
rect 1031 1000 1035 1002
rect 1095 1006 1099 1008
rect 1095 1000 1099 1002
rect 1159 1006 1163 1008
rect 1159 1000 1163 1002
rect 1223 1006 1227 1008
rect 1223 1000 1227 1002
rect 1279 1006 1283 1008
rect 1279 1001 1283 1002
rect 1287 1006 1291 1007
rect 1287 1000 1291 1002
rect 1335 1006 1339 1008
rect 1335 1001 1339 1002
rect 1343 1006 1347 1007
rect 1343 1000 1347 1002
rect 1383 1006 1387 1008
rect 1383 1001 1387 1002
rect 1399 1006 1403 1007
rect 1399 1000 1403 1002
rect 902 999 908 1000
rect 902 995 903 999
rect 907 995 908 999
rect 902 994 908 995
rect 966 999 972 1000
rect 966 995 967 999
rect 971 995 972 999
rect 966 994 972 995
rect 1030 999 1036 1000
rect 1030 995 1031 999
rect 1035 995 1036 999
rect 1030 994 1036 995
rect 1094 999 1100 1000
rect 1094 995 1095 999
rect 1099 995 1100 999
rect 1094 994 1100 995
rect 1158 999 1164 1000
rect 1158 995 1159 999
rect 1163 995 1164 999
rect 1158 994 1164 995
rect 1222 999 1228 1000
rect 1222 995 1223 999
rect 1227 995 1228 999
rect 1222 994 1228 995
rect 1286 999 1292 1000
rect 1286 995 1287 999
rect 1291 995 1292 999
rect 1286 994 1292 995
rect 1342 999 1348 1000
rect 1342 995 1343 999
rect 1347 995 1348 999
rect 1342 994 1348 995
rect 1398 999 1404 1000
rect 1398 995 1399 999
rect 1403 995 1404 999
rect 1398 994 1404 995
rect 1322 991 1328 992
rect 1322 987 1323 991
rect 1327 987 1328 991
rect 1322 986 1328 987
rect 902 982 908 983
rect 902 978 903 982
rect 907 978 908 982
rect 902 977 908 978
rect 966 982 972 983
rect 966 978 967 982
rect 971 978 972 982
rect 966 977 972 978
rect 1030 982 1036 983
rect 1030 978 1031 982
rect 1035 978 1036 982
rect 1030 977 1036 978
rect 1094 982 1100 983
rect 1094 978 1095 982
rect 1099 978 1100 982
rect 1094 977 1100 978
rect 1158 982 1164 983
rect 1158 978 1159 982
rect 1163 978 1164 982
rect 1158 977 1164 978
rect 1222 982 1228 983
rect 1222 978 1223 982
rect 1227 978 1228 982
rect 1222 977 1228 978
rect 1286 982 1292 983
rect 1286 978 1287 982
rect 1291 978 1292 982
rect 1286 977 1292 978
rect 890 975 896 976
rect 890 971 891 975
rect 895 971 896 975
rect 890 970 896 971
rect 904 967 906 977
rect 968 967 970 977
rect 1032 967 1034 977
rect 1096 967 1098 977
rect 1160 967 1162 977
rect 1182 967 1188 968
rect 1224 967 1226 977
rect 1288 967 1290 977
rect 831 966 835 967
rect 831 961 835 962
rect 847 966 851 967
rect 847 961 851 962
rect 903 966 907 967
rect 903 961 907 962
rect 911 966 915 967
rect 911 961 915 962
rect 967 966 971 967
rect 967 961 971 962
rect 975 966 979 967
rect 975 961 979 962
rect 1031 966 1035 967
rect 1031 961 1035 962
rect 1039 966 1043 967
rect 1039 961 1043 962
rect 1095 966 1099 967
rect 1095 961 1099 962
rect 1103 966 1107 967
rect 1103 961 1107 962
rect 1159 966 1163 967
rect 1159 961 1163 962
rect 1167 966 1171 967
rect 1182 963 1183 967
rect 1187 963 1188 967
rect 1182 962 1188 963
rect 1223 966 1227 967
rect 1167 961 1171 962
rect 806 955 812 956
rect 806 951 807 955
rect 811 951 812 955
rect 848 951 850 961
rect 862 955 868 956
rect 862 951 863 955
rect 867 951 868 955
rect 912 951 914 961
rect 976 951 978 961
rect 1040 951 1042 961
rect 1104 951 1106 961
rect 1168 951 1170 961
rect 470 950 476 951
rect 470 946 471 950
rect 475 946 476 950
rect 470 945 476 946
rect 534 950 540 951
rect 534 946 535 950
rect 539 946 540 950
rect 534 945 540 946
rect 598 950 604 951
rect 598 946 599 950
rect 603 946 604 950
rect 598 945 604 946
rect 662 950 668 951
rect 662 946 663 950
rect 667 946 668 950
rect 662 945 668 946
rect 726 950 732 951
rect 726 946 727 950
rect 731 946 732 950
rect 726 945 732 946
rect 790 950 796 951
rect 806 950 812 951
rect 846 950 852 951
rect 862 950 868 951
rect 910 950 916 951
rect 790 946 791 950
rect 795 946 796 950
rect 790 945 796 946
rect 846 946 847 950
rect 851 946 852 950
rect 846 945 852 946
rect 416 939 424 940
rect 416 936 419 939
rect 418 935 419 936
rect 423 935 424 939
rect 418 934 424 935
rect 674 939 680 940
rect 674 935 675 939
rect 679 935 680 939
rect 674 934 680 935
rect 758 939 764 940
rect 758 935 759 939
rect 763 935 764 939
rect 758 934 764 935
rect 198 933 204 934
rect 198 929 199 933
rect 203 929 204 933
rect 198 928 204 929
rect 238 933 244 934
rect 238 929 239 933
rect 243 929 244 933
rect 238 928 244 929
rect 286 933 292 934
rect 286 929 287 933
rect 291 929 292 933
rect 286 928 292 929
rect 342 933 348 934
rect 342 929 343 933
rect 347 929 348 933
rect 342 928 348 929
rect 406 933 412 934
rect 406 929 407 933
rect 411 929 412 933
rect 406 928 412 929
rect 470 933 476 934
rect 470 929 471 933
rect 475 929 476 933
rect 470 928 476 929
rect 534 933 540 934
rect 534 929 535 933
rect 539 929 540 933
rect 534 928 540 929
rect 598 933 604 934
rect 598 929 599 933
rect 603 929 604 933
rect 598 928 604 929
rect 662 933 668 934
rect 662 929 663 933
rect 667 929 668 933
rect 662 928 668 929
rect 186 923 192 924
rect 200 923 202 928
rect 240 923 242 928
rect 288 923 290 928
rect 344 923 346 928
rect 408 923 410 928
rect 472 923 474 928
rect 536 923 538 928
rect 600 923 602 928
rect 664 923 666 928
rect 111 922 115 923
rect 111 917 115 918
rect 135 922 139 923
rect 112 914 114 917
rect 135 916 139 918
rect 167 922 171 923
rect 186 919 187 923
rect 191 919 192 923
rect 186 918 192 919
rect 199 922 203 923
rect 167 916 171 918
rect 199 917 203 918
rect 207 922 211 923
rect 207 916 211 918
rect 239 922 243 923
rect 239 917 243 918
rect 271 922 275 923
rect 271 916 275 918
rect 287 922 291 923
rect 287 917 291 918
rect 335 922 339 923
rect 335 916 339 918
rect 343 922 347 923
rect 343 917 347 918
rect 407 922 411 923
rect 407 916 411 918
rect 471 922 475 923
rect 471 916 475 918
rect 535 922 539 923
rect 535 916 539 918
rect 591 922 595 923
rect 591 916 595 918
rect 599 922 603 923
rect 599 917 603 918
rect 647 922 651 923
rect 647 916 651 918
rect 663 922 667 923
rect 663 917 667 918
rect 134 915 140 916
rect 110 913 116 914
rect 110 909 111 913
rect 115 909 116 913
rect 134 911 135 915
rect 139 911 140 915
rect 134 910 140 911
rect 166 915 172 916
rect 166 911 167 915
rect 171 911 172 915
rect 166 910 172 911
rect 206 915 212 916
rect 206 911 207 915
rect 211 911 212 915
rect 206 910 212 911
rect 270 915 276 916
rect 270 911 271 915
rect 275 911 276 915
rect 270 910 276 911
rect 334 915 340 916
rect 334 911 335 915
rect 339 911 340 915
rect 334 910 340 911
rect 406 915 412 916
rect 406 911 407 915
rect 411 911 412 915
rect 406 910 412 911
rect 470 915 476 916
rect 470 911 471 915
rect 475 911 476 915
rect 470 910 476 911
rect 534 915 540 916
rect 534 911 535 915
rect 539 911 540 915
rect 534 910 540 911
rect 590 915 596 916
rect 590 911 591 915
rect 595 911 596 915
rect 590 910 596 911
rect 646 915 652 916
rect 646 911 647 915
rect 651 911 652 915
rect 646 910 652 911
rect 110 908 116 909
rect 486 907 492 908
rect 486 903 487 907
rect 491 903 492 907
rect 486 902 492 903
rect 666 907 672 908
rect 666 903 667 907
rect 671 903 672 907
rect 666 902 672 903
rect 134 898 140 899
rect 110 896 116 897
rect 110 892 111 896
rect 115 892 116 896
rect 134 894 135 898
rect 139 894 140 898
rect 134 893 140 894
rect 166 898 172 899
rect 166 894 167 898
rect 171 894 172 898
rect 166 893 172 894
rect 206 898 212 899
rect 206 894 207 898
rect 211 894 212 898
rect 206 893 212 894
rect 270 898 276 899
rect 270 894 271 898
rect 275 894 276 898
rect 270 893 276 894
rect 334 898 340 899
rect 334 894 335 898
rect 339 894 340 898
rect 334 893 340 894
rect 406 898 412 899
rect 406 894 407 898
rect 411 894 412 898
rect 406 893 412 894
rect 470 898 476 899
rect 470 894 471 898
rect 475 894 476 898
rect 470 893 476 894
rect 110 891 116 892
rect 112 879 114 891
rect 136 879 138 893
rect 168 879 170 893
rect 208 879 210 893
rect 272 879 274 893
rect 336 879 338 893
rect 408 879 410 893
rect 422 883 428 884
rect 422 879 423 883
rect 427 879 428 883
rect 472 879 474 893
rect 111 878 115 879
rect 111 873 115 874
rect 135 878 139 879
rect 135 873 139 874
rect 167 878 171 879
rect 167 873 171 874
rect 207 878 211 879
rect 207 873 211 874
rect 271 878 275 879
rect 271 873 275 874
rect 335 878 339 879
rect 335 873 339 874
rect 407 878 411 879
rect 422 878 428 879
rect 471 878 475 879
rect 407 873 411 874
rect 112 865 114 873
rect 110 864 116 865
rect 110 860 111 864
rect 115 860 116 864
rect 136 863 138 873
rect 150 867 156 868
rect 150 863 151 867
rect 155 863 156 867
rect 168 863 170 873
rect 208 863 210 873
rect 272 863 274 873
rect 336 863 338 873
rect 408 863 410 873
rect 110 859 116 860
rect 134 862 140 863
rect 150 862 156 863
rect 166 862 172 863
rect 134 858 135 862
rect 139 858 140 862
rect 134 857 140 858
rect 110 847 116 848
rect 110 843 111 847
rect 115 843 116 847
rect 110 842 116 843
rect 134 845 140 846
rect 112 839 114 842
rect 134 841 135 845
rect 139 841 140 845
rect 134 840 140 841
rect 111 838 115 839
rect 111 833 115 834
rect 135 838 139 840
rect 112 830 114 833
rect 135 832 139 834
rect 134 831 140 832
rect 110 829 116 830
rect 110 825 111 829
rect 115 825 116 829
rect 134 827 135 831
rect 139 827 140 831
rect 134 826 140 827
rect 110 824 116 825
rect 152 824 154 862
rect 166 858 167 862
rect 171 858 172 862
rect 166 857 172 858
rect 206 862 212 863
rect 206 858 207 862
rect 211 858 212 862
rect 206 857 212 858
rect 270 862 276 863
rect 270 858 271 862
rect 275 858 276 862
rect 270 857 276 858
rect 334 862 340 863
rect 334 858 335 862
rect 339 858 340 862
rect 334 857 340 858
rect 406 862 412 863
rect 406 858 407 862
rect 411 858 412 862
rect 406 857 412 858
rect 424 852 426 878
rect 471 873 475 874
rect 472 863 474 873
rect 488 868 490 902
rect 534 898 540 899
rect 534 894 535 898
rect 539 894 540 898
rect 534 893 540 894
rect 590 898 596 899
rect 590 894 591 898
rect 595 894 596 898
rect 590 893 596 894
rect 646 898 652 899
rect 646 894 647 898
rect 651 894 652 898
rect 646 893 652 894
rect 536 879 538 893
rect 592 879 594 893
rect 648 879 650 893
rect 535 878 539 879
rect 591 878 595 879
rect 535 873 539 874
rect 558 875 564 876
rect 486 867 492 868
rect 486 863 487 867
rect 491 863 492 867
rect 536 863 538 873
rect 558 871 559 875
rect 563 871 564 875
rect 591 873 595 874
rect 599 878 603 879
rect 599 873 603 874
rect 647 878 651 879
rect 647 873 651 874
rect 655 878 659 879
rect 655 873 659 874
rect 558 870 564 871
rect 470 862 476 863
rect 486 862 492 863
rect 534 862 540 863
rect 470 858 471 862
rect 475 858 476 862
rect 470 857 476 858
rect 534 858 535 862
rect 539 858 540 862
rect 534 857 540 858
rect 422 851 428 852
rect 422 847 423 851
rect 427 847 428 851
rect 422 846 428 847
rect 551 851 557 852
rect 551 847 552 851
rect 556 850 557 851
rect 560 850 562 870
rect 600 863 602 873
rect 646 867 652 868
rect 646 863 647 867
rect 651 863 652 867
rect 656 863 658 873
rect 668 868 670 902
rect 676 900 678 934
rect 726 933 732 934
rect 726 929 727 933
rect 731 929 732 933
rect 726 928 732 929
rect 728 923 730 928
rect 703 922 707 923
rect 703 916 707 918
rect 727 922 731 923
rect 727 917 731 918
rect 751 922 755 923
rect 751 916 755 918
rect 702 915 708 916
rect 702 911 703 915
rect 707 911 708 915
rect 702 910 708 911
rect 750 915 756 916
rect 750 911 751 915
rect 755 911 756 915
rect 750 910 756 911
rect 674 899 680 900
rect 674 895 675 899
rect 679 895 680 899
rect 674 894 680 895
rect 702 898 708 899
rect 702 894 703 898
rect 707 894 708 898
rect 702 893 708 894
rect 750 898 756 899
rect 750 894 751 898
rect 755 894 756 898
rect 750 893 756 894
rect 704 879 706 893
rect 752 879 754 893
rect 760 892 762 934
rect 790 933 796 934
rect 790 929 791 933
rect 795 929 796 933
rect 790 928 796 929
rect 846 933 852 934
rect 846 929 847 933
rect 851 929 852 933
rect 846 928 852 929
rect 792 923 794 928
rect 848 923 850 928
rect 864 924 866 950
rect 910 946 911 950
rect 915 946 916 950
rect 910 945 916 946
rect 974 950 980 951
rect 974 946 975 950
rect 979 946 980 950
rect 974 945 980 946
rect 1038 950 1044 951
rect 1038 946 1039 950
rect 1043 946 1044 950
rect 1038 945 1044 946
rect 1102 950 1108 951
rect 1102 946 1103 950
rect 1107 946 1108 950
rect 1102 945 1108 946
rect 1166 950 1172 951
rect 1166 946 1167 950
rect 1171 946 1172 950
rect 1166 945 1172 946
rect 1184 940 1186 962
rect 1223 961 1227 962
rect 1231 966 1235 967
rect 1231 961 1235 962
rect 1287 966 1291 967
rect 1324 964 1326 986
rect 1342 982 1348 983
rect 1342 978 1343 982
rect 1347 978 1348 982
rect 1342 977 1348 978
rect 1398 982 1404 983
rect 1398 978 1399 982
rect 1403 978 1404 982
rect 1398 977 1404 978
rect 1344 967 1346 977
rect 1400 967 1402 977
rect 1416 976 1418 1014
rect 1430 1013 1436 1014
rect 1430 1009 1431 1013
rect 1435 1009 1436 1013
rect 1430 1008 1436 1009
rect 1478 1013 1484 1014
rect 1478 1009 1479 1013
rect 1483 1009 1484 1013
rect 1478 1008 1484 1009
rect 1534 1013 1540 1014
rect 1534 1009 1535 1013
rect 1539 1009 1540 1013
rect 1534 1008 1540 1009
rect 1431 1006 1435 1008
rect 1431 1001 1435 1002
rect 1447 1006 1451 1007
rect 1447 1000 1451 1002
rect 1479 1006 1483 1008
rect 1479 1001 1483 1002
rect 1495 1006 1499 1007
rect 1495 1000 1499 1002
rect 1535 1006 1539 1008
rect 1535 1001 1539 1002
rect 1543 1006 1547 1007
rect 1543 1000 1547 1002
rect 1446 999 1452 1000
rect 1446 995 1447 999
rect 1451 995 1452 999
rect 1446 994 1452 995
rect 1494 999 1500 1000
rect 1494 995 1495 999
rect 1499 995 1500 999
rect 1494 994 1500 995
rect 1542 999 1548 1000
rect 1542 995 1543 999
rect 1547 995 1548 999
rect 1542 994 1548 995
rect 1556 992 1558 1030
rect 1590 1026 1591 1030
rect 1595 1026 1596 1030
rect 1590 1025 1596 1026
rect 1622 1026 1623 1030
rect 1627 1026 1628 1030
rect 1662 1028 1663 1032
rect 1667 1028 1668 1032
rect 1662 1027 1668 1028
rect 1622 1025 1628 1026
rect 1638 1019 1644 1020
rect 1638 1015 1639 1019
rect 1643 1015 1644 1019
rect 1638 1014 1644 1015
rect 1662 1015 1668 1016
rect 1590 1013 1596 1014
rect 1590 1009 1591 1013
rect 1595 1009 1596 1013
rect 1590 1008 1596 1009
rect 1622 1013 1628 1014
rect 1622 1009 1623 1013
rect 1627 1009 1628 1013
rect 1622 1008 1628 1009
rect 1591 1006 1595 1008
rect 1591 1000 1595 1002
rect 1623 1006 1627 1008
rect 1623 1000 1627 1002
rect 1590 999 1596 1000
rect 1590 995 1591 999
rect 1595 995 1596 999
rect 1590 994 1596 995
rect 1622 999 1628 1000
rect 1622 995 1623 999
rect 1627 995 1628 999
rect 1622 994 1628 995
rect 1554 991 1560 992
rect 1554 987 1555 991
rect 1559 987 1560 991
rect 1554 986 1560 987
rect 1606 991 1612 992
rect 1606 987 1607 991
rect 1611 987 1612 991
rect 1606 986 1612 987
rect 1446 982 1452 983
rect 1446 978 1447 982
rect 1451 978 1452 982
rect 1446 977 1452 978
rect 1494 982 1500 983
rect 1494 978 1495 982
rect 1499 978 1500 982
rect 1494 977 1500 978
rect 1542 982 1548 983
rect 1542 978 1543 982
rect 1547 978 1548 982
rect 1542 977 1548 978
rect 1590 982 1596 983
rect 1590 978 1591 982
rect 1595 978 1596 982
rect 1590 977 1596 978
rect 1414 975 1420 976
rect 1414 971 1415 975
rect 1419 971 1420 975
rect 1414 970 1420 971
rect 1448 967 1450 977
rect 1458 975 1464 976
rect 1458 971 1459 975
rect 1463 971 1464 975
rect 1458 970 1464 971
rect 1343 966 1347 967
rect 1287 961 1291 962
rect 1322 963 1328 964
rect 1232 951 1234 961
rect 1288 951 1290 961
rect 1322 959 1323 963
rect 1327 959 1328 963
rect 1343 961 1347 962
rect 1391 966 1395 967
rect 1391 961 1395 962
rect 1399 966 1403 967
rect 1399 961 1403 962
rect 1431 966 1435 967
rect 1431 961 1435 962
rect 1447 966 1451 967
rect 1447 961 1451 962
rect 1322 958 1328 959
rect 1344 951 1346 961
rect 1392 951 1394 961
rect 1432 951 1434 961
rect 1230 950 1236 951
rect 1230 946 1231 950
rect 1235 946 1236 950
rect 1230 945 1236 946
rect 1286 950 1292 951
rect 1286 946 1287 950
rect 1291 946 1292 950
rect 1286 945 1292 946
rect 1342 950 1348 951
rect 1342 946 1343 950
rect 1347 946 1348 950
rect 1342 945 1348 946
rect 1390 950 1396 951
rect 1390 946 1391 950
rect 1395 946 1396 950
rect 1390 945 1396 946
rect 1430 950 1436 951
rect 1430 946 1431 950
rect 1435 946 1436 950
rect 1430 945 1436 946
rect 1460 944 1462 970
rect 1486 967 1492 968
rect 1496 967 1498 977
rect 1544 967 1546 977
rect 1592 967 1594 977
rect 1471 966 1475 967
rect 1486 963 1487 967
rect 1491 963 1492 967
rect 1486 962 1492 963
rect 1495 966 1499 967
rect 1471 961 1475 962
rect 1472 951 1474 961
rect 1470 950 1476 951
rect 1470 946 1471 950
rect 1475 946 1476 950
rect 1470 945 1476 946
rect 1458 943 1464 944
rect 1182 939 1188 940
rect 1182 935 1183 939
rect 1187 935 1188 939
rect 1458 939 1459 943
rect 1463 939 1464 943
rect 1488 940 1490 962
rect 1495 961 1499 962
rect 1511 966 1515 967
rect 1511 961 1515 962
rect 1543 966 1547 967
rect 1543 961 1547 962
rect 1551 966 1555 967
rect 1551 961 1555 962
rect 1591 966 1595 967
rect 1591 961 1595 962
rect 1512 951 1514 961
rect 1552 951 1554 961
rect 1582 955 1588 956
rect 1582 951 1583 955
rect 1587 951 1588 955
rect 1592 951 1594 961
rect 1608 956 1610 986
rect 1622 982 1628 983
rect 1622 978 1623 982
rect 1627 978 1628 982
rect 1622 977 1628 978
rect 1624 967 1626 977
rect 1640 976 1642 1014
rect 1662 1011 1663 1015
rect 1667 1011 1668 1015
rect 1662 1010 1668 1011
rect 1664 1007 1666 1010
rect 1663 1006 1667 1007
rect 1663 1001 1667 1002
rect 1664 998 1666 1001
rect 1662 997 1668 998
rect 1662 993 1663 997
rect 1667 993 1668 997
rect 1662 992 1668 993
rect 1662 980 1668 981
rect 1662 976 1663 980
rect 1667 976 1668 980
rect 1638 975 1644 976
rect 1662 975 1668 976
rect 1638 971 1639 975
rect 1643 971 1644 975
rect 1638 970 1644 971
rect 1664 967 1666 975
rect 1623 966 1627 967
rect 1623 961 1627 962
rect 1663 966 1667 967
rect 1663 961 1667 962
rect 1606 955 1612 956
rect 1606 951 1607 955
rect 1611 951 1612 955
rect 1624 951 1626 961
rect 1664 953 1666 961
rect 1662 952 1668 953
rect 1510 950 1516 951
rect 1510 946 1511 950
rect 1515 946 1516 950
rect 1510 945 1516 946
rect 1550 950 1556 951
rect 1582 950 1588 951
rect 1590 950 1596 951
rect 1606 950 1612 951
rect 1622 950 1628 951
rect 1550 946 1551 950
rect 1555 946 1556 950
rect 1550 945 1556 946
rect 1458 938 1464 939
rect 1486 939 1492 940
rect 1182 934 1188 935
rect 1486 935 1487 939
rect 1491 935 1492 939
rect 1486 934 1492 935
rect 910 933 916 934
rect 910 929 911 933
rect 915 929 916 933
rect 910 928 916 929
rect 974 933 980 934
rect 974 929 975 933
rect 979 929 980 933
rect 974 928 980 929
rect 1038 933 1044 934
rect 1038 929 1039 933
rect 1043 929 1044 933
rect 1038 928 1044 929
rect 1102 933 1108 934
rect 1102 929 1103 933
rect 1107 929 1108 933
rect 1102 928 1108 929
rect 1166 933 1172 934
rect 1166 929 1167 933
rect 1171 929 1172 933
rect 1166 928 1172 929
rect 1230 933 1236 934
rect 1230 929 1231 933
rect 1235 929 1236 933
rect 1230 928 1236 929
rect 1286 933 1292 934
rect 1286 929 1287 933
rect 1291 929 1292 933
rect 1286 928 1292 929
rect 1342 933 1348 934
rect 1342 929 1343 933
rect 1347 929 1348 933
rect 1342 928 1348 929
rect 1390 933 1396 934
rect 1390 929 1391 933
rect 1395 929 1396 933
rect 1390 928 1396 929
rect 1430 933 1436 934
rect 1430 929 1431 933
rect 1435 929 1436 933
rect 1430 928 1436 929
rect 1470 933 1476 934
rect 1470 929 1471 933
rect 1475 929 1476 933
rect 1470 928 1476 929
rect 1510 933 1516 934
rect 1510 929 1511 933
rect 1515 929 1516 933
rect 1510 928 1516 929
rect 1550 933 1556 934
rect 1550 929 1551 933
rect 1555 929 1556 933
rect 1550 928 1556 929
rect 1584 928 1586 950
rect 1590 946 1591 950
rect 1595 946 1596 950
rect 1590 945 1596 946
rect 1622 946 1623 950
rect 1627 946 1628 950
rect 1662 948 1663 952
rect 1667 948 1668 952
rect 1662 947 1668 948
rect 1622 945 1628 946
rect 1662 935 1668 936
rect 1590 933 1596 934
rect 1590 929 1591 933
rect 1595 929 1596 933
rect 1590 928 1596 929
rect 1622 933 1628 934
rect 1622 929 1623 933
rect 1627 929 1628 933
rect 1662 931 1663 935
rect 1667 931 1668 935
rect 1662 930 1668 931
rect 1622 928 1628 929
rect 862 923 868 924
rect 912 923 914 928
rect 976 923 978 928
rect 1040 923 1042 928
rect 1104 923 1106 928
rect 1168 923 1170 928
rect 1174 927 1180 928
rect 1174 923 1175 927
rect 1179 923 1180 927
rect 1232 923 1234 928
rect 1288 923 1290 928
rect 1344 923 1346 928
rect 1392 923 1394 928
rect 1432 923 1434 928
rect 1472 923 1474 928
rect 1512 923 1514 928
rect 1552 923 1554 928
rect 1582 927 1588 928
rect 1582 923 1583 927
rect 1587 923 1588 927
rect 1592 923 1594 928
rect 1624 923 1626 928
rect 1664 923 1666 930
rect 791 922 795 923
rect 791 917 795 918
rect 799 922 803 923
rect 799 916 803 918
rect 847 922 851 923
rect 862 919 863 923
rect 867 919 868 923
rect 862 918 868 919
rect 903 922 907 923
rect 847 916 851 918
rect 903 916 907 918
rect 911 922 915 923
rect 911 917 915 918
rect 959 922 963 923
rect 959 916 963 918
rect 975 922 979 923
rect 975 917 979 918
rect 1023 922 1027 923
rect 1023 916 1027 918
rect 1039 922 1043 923
rect 1039 917 1043 918
rect 1087 922 1091 923
rect 1087 916 1091 918
rect 1103 922 1107 923
rect 1103 917 1107 918
rect 1143 922 1147 923
rect 1143 916 1147 918
rect 1167 922 1171 923
rect 1174 922 1180 923
rect 1199 922 1203 923
rect 1167 917 1171 918
rect 798 915 804 916
rect 798 911 799 915
rect 803 911 804 915
rect 798 910 804 911
rect 846 915 852 916
rect 846 911 847 915
rect 851 911 852 915
rect 846 910 852 911
rect 902 915 908 916
rect 902 911 903 915
rect 907 911 908 915
rect 902 910 908 911
rect 958 915 964 916
rect 958 911 959 915
rect 963 911 964 915
rect 958 910 964 911
rect 1022 915 1028 916
rect 1022 911 1023 915
rect 1027 911 1028 915
rect 1022 910 1028 911
rect 1086 915 1092 916
rect 1086 911 1087 915
rect 1091 911 1092 915
rect 1086 910 1092 911
rect 1142 915 1148 916
rect 1142 911 1143 915
rect 1147 911 1148 915
rect 1142 910 1148 911
rect 798 898 804 899
rect 798 894 799 898
rect 803 894 804 898
rect 798 893 804 894
rect 846 898 852 899
rect 846 894 847 898
rect 851 894 852 898
rect 846 893 852 894
rect 902 898 908 899
rect 902 894 903 898
rect 907 894 908 898
rect 902 893 908 894
rect 958 898 964 899
rect 958 894 959 898
rect 963 894 964 898
rect 958 893 964 894
rect 1022 898 1028 899
rect 1022 894 1023 898
rect 1027 894 1028 898
rect 1022 893 1028 894
rect 1086 898 1092 899
rect 1086 894 1087 898
rect 1091 894 1092 898
rect 1086 893 1092 894
rect 1142 898 1148 899
rect 1142 894 1143 898
rect 1147 894 1148 898
rect 1142 893 1148 894
rect 758 891 764 892
rect 758 887 759 891
rect 763 887 764 891
rect 758 886 764 887
rect 800 879 802 893
rect 814 891 820 892
rect 814 887 815 891
rect 819 887 820 891
rect 814 886 820 887
rect 703 878 707 879
rect 703 873 707 874
rect 751 878 755 879
rect 751 873 755 874
rect 799 878 803 879
rect 799 873 803 874
rect 666 867 672 868
rect 666 863 667 867
rect 671 863 672 867
rect 704 863 706 873
rect 752 863 754 873
rect 800 863 802 873
rect 598 862 604 863
rect 646 862 652 863
rect 654 862 660 863
rect 666 862 672 863
rect 702 862 708 863
rect 598 858 599 862
rect 603 858 604 862
rect 598 857 604 858
rect 556 848 562 850
rect 618 851 624 852
rect 556 847 557 848
rect 551 846 557 847
rect 618 847 619 851
rect 623 847 624 851
rect 648 851 650 862
rect 654 858 655 862
rect 659 858 660 862
rect 654 857 660 858
rect 702 858 703 862
rect 707 858 708 862
rect 702 857 708 858
rect 750 862 756 863
rect 750 858 751 862
rect 755 858 756 862
rect 750 857 756 858
rect 798 862 804 863
rect 798 858 799 862
rect 803 858 804 862
rect 798 857 804 858
rect 816 852 818 886
rect 848 879 850 893
rect 904 879 906 893
rect 960 879 962 893
rect 1024 879 1026 893
rect 1088 879 1090 893
rect 1118 879 1124 880
rect 1144 879 1146 893
rect 1176 892 1178 922
rect 1199 916 1203 918
rect 1231 922 1235 923
rect 1231 917 1235 918
rect 1255 922 1259 923
rect 1255 916 1259 918
rect 1287 922 1291 923
rect 1287 917 1291 918
rect 1319 922 1323 923
rect 1319 916 1323 918
rect 1343 922 1347 923
rect 1343 917 1347 918
rect 1383 922 1387 923
rect 1383 916 1387 918
rect 1391 922 1395 923
rect 1391 917 1395 918
rect 1431 922 1435 923
rect 1431 917 1435 918
rect 1471 922 1475 923
rect 1471 917 1475 918
rect 1511 922 1515 923
rect 1511 917 1515 918
rect 1551 922 1555 923
rect 1582 922 1588 923
rect 1591 922 1595 923
rect 1551 917 1555 918
rect 1591 917 1595 918
rect 1623 922 1627 923
rect 1623 917 1627 918
rect 1663 922 1667 923
rect 1663 917 1667 918
rect 1198 915 1204 916
rect 1198 911 1199 915
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1254 915 1260 916
rect 1254 911 1255 915
rect 1259 911 1260 915
rect 1254 910 1260 911
rect 1318 915 1324 916
rect 1318 911 1319 915
rect 1323 911 1324 915
rect 1318 910 1324 911
rect 1382 915 1388 916
rect 1382 911 1383 915
rect 1387 911 1388 915
rect 1664 914 1666 917
rect 1382 910 1388 911
rect 1662 913 1668 914
rect 1662 909 1663 913
rect 1667 909 1668 913
rect 1662 908 1668 909
rect 1374 907 1380 908
rect 1374 903 1375 907
rect 1379 903 1380 907
rect 1374 902 1380 903
rect 1198 898 1204 899
rect 1198 894 1199 898
rect 1203 894 1204 898
rect 1198 893 1204 894
rect 1254 898 1260 899
rect 1254 894 1255 898
rect 1259 894 1260 898
rect 1254 893 1260 894
rect 1318 898 1324 899
rect 1318 894 1319 898
rect 1323 894 1324 898
rect 1318 893 1324 894
rect 1174 891 1180 892
rect 1174 887 1175 891
rect 1179 887 1180 891
rect 1174 886 1180 887
rect 1200 879 1202 893
rect 1256 879 1258 893
rect 1320 879 1322 893
rect 1376 880 1378 902
rect 1382 898 1388 899
rect 1382 894 1383 898
rect 1387 894 1388 898
rect 1382 893 1388 894
rect 1662 896 1668 897
rect 1374 879 1380 880
rect 1384 879 1386 893
rect 1662 892 1663 896
rect 1667 892 1668 896
rect 1662 891 1668 892
rect 1664 879 1666 891
rect 847 878 851 879
rect 847 873 851 874
rect 903 878 907 879
rect 903 873 907 874
rect 959 878 963 879
rect 959 873 963 874
rect 967 878 971 879
rect 967 873 971 874
rect 1023 878 1027 879
rect 1023 873 1027 874
rect 1039 878 1043 879
rect 1039 873 1043 874
rect 1087 878 1091 879
rect 1087 873 1091 874
rect 1103 878 1107 879
rect 1118 875 1119 879
rect 1123 875 1124 879
rect 1118 874 1124 875
rect 1143 878 1147 879
rect 1103 873 1107 874
rect 848 863 850 873
rect 904 863 906 873
rect 968 863 970 873
rect 1040 863 1042 873
rect 1054 867 1060 868
rect 1054 863 1055 867
rect 1059 863 1060 867
rect 1104 863 1106 873
rect 846 862 852 863
rect 846 858 847 862
rect 851 858 852 862
rect 846 857 852 858
rect 902 862 908 863
rect 902 858 903 862
rect 907 858 908 862
rect 902 857 908 858
rect 966 862 972 863
rect 966 858 967 862
rect 971 858 972 862
rect 966 857 972 858
rect 1038 862 1044 863
rect 1054 862 1060 863
rect 1102 862 1108 863
rect 1038 858 1039 862
rect 1043 858 1044 862
rect 1038 857 1044 858
rect 666 851 672 852
rect 648 849 667 851
rect 618 846 624 847
rect 666 847 667 849
rect 671 847 672 851
rect 666 846 672 847
rect 814 851 820 852
rect 814 847 815 851
rect 819 847 820 851
rect 814 846 820 847
rect 166 845 172 846
rect 166 841 167 845
rect 171 841 172 845
rect 166 840 172 841
rect 206 845 212 846
rect 206 841 207 845
rect 211 841 212 845
rect 206 840 212 841
rect 270 845 276 846
rect 270 841 271 845
rect 275 841 276 845
rect 270 840 276 841
rect 334 845 340 846
rect 334 841 335 845
rect 339 841 340 845
rect 334 840 340 841
rect 406 845 412 846
rect 406 841 407 845
rect 411 841 412 845
rect 406 840 412 841
rect 470 845 476 846
rect 470 841 471 845
rect 475 841 476 845
rect 470 840 476 841
rect 534 845 540 846
rect 534 841 535 845
rect 539 841 540 845
rect 534 840 540 841
rect 598 845 604 846
rect 598 841 599 845
rect 603 841 604 845
rect 598 840 604 841
rect 167 838 171 840
rect 167 832 171 834
rect 207 838 211 840
rect 207 833 211 834
rect 215 838 219 839
rect 215 832 219 834
rect 271 838 275 840
rect 271 833 275 834
rect 279 838 283 839
rect 279 832 283 834
rect 335 838 339 840
rect 335 833 339 834
rect 343 838 347 839
rect 343 832 347 834
rect 407 838 411 840
rect 407 833 411 834
rect 415 838 419 839
rect 415 832 419 834
rect 471 838 475 840
rect 471 833 475 834
rect 479 838 483 839
rect 479 832 483 834
rect 535 838 539 840
rect 535 833 539 834
rect 543 838 547 839
rect 543 832 547 834
rect 599 838 603 840
rect 599 833 603 834
rect 607 838 611 839
rect 607 832 611 834
rect 166 831 172 832
rect 166 827 167 831
rect 171 827 172 831
rect 166 826 172 827
rect 214 831 220 832
rect 214 827 215 831
rect 219 827 220 831
rect 214 826 220 827
rect 278 831 284 832
rect 278 827 279 831
rect 283 827 284 831
rect 278 826 284 827
rect 342 831 348 832
rect 342 827 343 831
rect 347 827 348 831
rect 342 826 348 827
rect 414 831 420 832
rect 414 827 415 831
rect 419 827 420 831
rect 414 826 420 827
rect 478 831 484 832
rect 478 827 479 831
rect 483 827 484 831
rect 478 826 484 827
rect 542 831 548 832
rect 542 827 543 831
rect 547 827 548 831
rect 542 826 548 827
rect 606 831 612 832
rect 606 827 607 831
rect 611 827 612 831
rect 606 826 612 827
rect 150 823 156 824
rect 150 819 151 823
rect 155 819 156 823
rect 150 818 156 819
rect 402 823 408 824
rect 402 819 403 823
rect 407 819 408 823
rect 402 818 408 819
rect 534 823 540 824
rect 534 819 535 823
rect 539 819 540 823
rect 534 818 540 819
rect 134 814 140 815
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 134 810 135 814
rect 139 810 140 814
rect 134 809 140 810
rect 166 814 172 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 214 814 220 815
rect 214 810 215 814
rect 219 810 220 814
rect 214 809 220 810
rect 278 814 284 815
rect 278 810 279 814
rect 283 810 284 814
rect 278 809 284 810
rect 342 814 348 815
rect 342 810 343 814
rect 347 810 348 814
rect 342 809 348 810
rect 110 807 116 808
rect 112 795 114 807
rect 136 795 138 809
rect 168 795 170 809
rect 216 795 218 809
rect 280 795 282 809
rect 286 807 292 808
rect 286 803 287 807
rect 291 803 292 807
rect 286 802 292 803
rect 111 794 115 795
rect 111 789 115 790
rect 135 794 139 795
rect 135 789 139 790
rect 167 794 171 795
rect 167 789 171 790
rect 175 794 179 795
rect 175 789 179 790
rect 215 794 219 795
rect 215 789 219 790
rect 231 794 235 795
rect 231 789 235 790
rect 279 794 283 795
rect 279 789 283 790
rect 112 781 114 789
rect 110 780 116 781
rect 110 776 111 780
rect 115 776 116 780
rect 136 779 138 789
rect 150 783 156 784
rect 150 779 151 783
rect 155 779 156 783
rect 176 779 178 789
rect 232 779 234 789
rect 110 775 116 776
rect 134 778 140 779
rect 150 778 156 779
rect 174 778 180 779
rect 134 774 135 778
rect 139 774 140 778
rect 134 773 140 774
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 110 758 116 759
rect 134 761 140 762
rect 112 755 114 758
rect 134 757 135 761
rect 139 757 140 761
rect 134 756 140 757
rect 152 756 154 778
rect 174 774 175 778
rect 179 774 180 778
rect 174 773 180 774
rect 230 778 236 779
rect 230 774 231 778
rect 235 774 236 778
rect 230 773 236 774
rect 288 768 290 802
rect 344 795 346 809
rect 404 800 406 818
rect 414 814 420 815
rect 414 810 415 814
rect 419 810 420 814
rect 414 809 420 810
rect 478 814 484 815
rect 478 810 479 814
rect 483 810 484 814
rect 478 809 484 810
rect 402 799 408 800
rect 402 795 403 799
rect 407 795 408 799
rect 416 795 418 809
rect 480 795 482 809
rect 295 794 299 795
rect 295 789 299 790
rect 343 794 347 795
rect 343 789 347 790
rect 367 794 371 795
rect 402 794 408 795
rect 415 794 419 795
rect 367 789 371 790
rect 415 789 419 790
rect 447 794 451 795
rect 447 789 451 790
rect 479 794 483 795
rect 479 789 483 790
rect 527 794 531 795
rect 527 789 531 790
rect 296 779 298 789
rect 350 787 356 788
rect 306 783 312 784
rect 306 779 307 783
rect 311 779 312 783
rect 350 783 351 787
rect 355 783 356 787
rect 350 782 356 783
rect 294 778 300 779
rect 306 778 312 779
rect 294 774 295 778
rect 299 774 300 778
rect 294 773 300 774
rect 286 767 292 768
rect 286 763 287 767
rect 291 763 292 767
rect 286 762 292 763
rect 174 761 180 762
rect 174 757 175 761
rect 179 757 180 761
rect 174 756 180 757
rect 230 761 236 762
rect 230 757 231 761
rect 235 757 236 761
rect 230 756 236 757
rect 294 761 300 762
rect 294 757 295 761
rect 299 757 300 761
rect 294 756 300 757
rect 111 754 115 755
rect 111 749 115 750
rect 135 754 139 756
rect 150 755 156 756
rect 150 751 151 755
rect 155 751 156 755
rect 150 750 156 751
rect 175 754 179 756
rect 135 749 139 750
rect 175 749 179 750
rect 215 754 219 755
rect 112 746 114 749
rect 215 748 219 750
rect 231 754 235 756
rect 231 749 235 750
rect 247 754 251 755
rect 247 748 251 750
rect 279 754 283 755
rect 279 748 283 750
rect 295 754 299 756
rect 295 749 299 750
rect 214 747 220 748
rect 110 745 116 746
rect 110 741 111 745
rect 115 741 116 745
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 246 747 252 748
rect 246 743 247 747
rect 251 743 252 747
rect 246 742 252 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 308 744 310 778
rect 352 768 354 782
rect 368 779 370 789
rect 448 779 450 789
rect 528 779 530 789
rect 536 784 538 818
rect 542 814 548 815
rect 542 810 543 814
rect 547 810 548 814
rect 542 809 548 810
rect 606 814 612 815
rect 606 810 607 814
rect 611 810 612 814
rect 606 809 612 810
rect 544 795 546 809
rect 608 795 610 809
rect 620 808 622 846
rect 654 845 660 846
rect 654 841 655 845
rect 659 841 660 845
rect 654 840 660 841
rect 702 845 708 846
rect 702 841 703 845
rect 707 841 708 845
rect 702 840 708 841
rect 750 845 756 846
rect 750 841 751 845
rect 755 841 756 845
rect 750 840 756 841
rect 798 845 804 846
rect 798 841 799 845
rect 803 841 804 845
rect 798 840 804 841
rect 846 845 852 846
rect 846 841 847 845
rect 851 841 852 845
rect 846 840 852 841
rect 902 845 908 846
rect 902 841 903 845
rect 907 841 908 845
rect 902 840 908 841
rect 966 845 972 846
rect 966 841 967 845
rect 971 841 972 845
rect 966 840 972 841
rect 1038 845 1044 846
rect 1038 841 1039 845
rect 1043 841 1044 845
rect 1038 840 1044 841
rect 655 838 659 840
rect 690 839 696 840
rect 655 833 659 834
rect 671 838 675 839
rect 690 835 691 839
rect 695 835 696 839
rect 690 834 696 835
rect 703 838 707 840
rect 671 832 675 834
rect 670 831 676 832
rect 670 827 671 831
rect 675 827 676 831
rect 670 826 676 827
rect 670 814 676 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 618 807 624 808
rect 618 803 619 807
rect 623 803 624 807
rect 618 802 624 803
rect 672 795 674 809
rect 692 808 694 834
rect 703 833 707 834
rect 735 838 739 839
rect 735 832 739 834
rect 751 838 755 840
rect 751 833 755 834
rect 791 838 795 839
rect 791 832 795 834
rect 799 838 803 840
rect 799 833 803 834
rect 847 838 851 840
rect 847 832 851 834
rect 903 838 907 840
rect 903 833 907 834
rect 911 838 915 839
rect 911 832 915 834
rect 967 838 971 840
rect 967 833 971 834
rect 975 838 979 839
rect 975 832 979 834
rect 1039 838 1043 840
rect 1039 832 1043 834
rect 734 831 740 832
rect 734 827 735 831
rect 739 827 740 831
rect 734 826 740 827
rect 790 831 796 832
rect 790 827 791 831
rect 795 827 796 831
rect 790 826 796 827
rect 846 831 852 832
rect 846 827 847 831
rect 851 827 852 831
rect 846 826 852 827
rect 910 831 916 832
rect 910 827 911 831
rect 915 827 916 831
rect 910 826 916 827
rect 974 831 980 832
rect 974 827 975 831
rect 979 827 980 831
rect 974 826 980 827
rect 1038 831 1044 832
rect 1038 827 1039 831
rect 1043 827 1044 831
rect 1038 826 1044 827
rect 1056 824 1058 862
rect 1102 858 1103 862
rect 1107 858 1108 862
rect 1102 857 1108 858
rect 1120 852 1122 874
rect 1143 873 1147 874
rect 1167 878 1171 879
rect 1167 873 1171 874
rect 1199 878 1203 879
rect 1199 873 1203 874
rect 1231 878 1235 879
rect 1231 873 1235 874
rect 1255 878 1259 879
rect 1255 873 1259 874
rect 1287 878 1291 879
rect 1287 873 1291 874
rect 1319 878 1323 879
rect 1319 873 1323 874
rect 1343 878 1347 879
rect 1374 875 1375 879
rect 1379 875 1380 879
rect 1374 874 1380 875
rect 1383 878 1387 879
rect 1343 873 1347 874
rect 1383 873 1387 874
rect 1399 878 1403 879
rect 1399 873 1403 874
rect 1463 878 1467 879
rect 1463 873 1467 874
rect 1663 878 1667 879
rect 1663 873 1667 874
rect 1168 863 1170 873
rect 1232 863 1234 873
rect 1288 863 1290 873
rect 1344 863 1346 873
rect 1400 863 1402 873
rect 1464 863 1466 873
rect 1664 865 1666 873
rect 1662 864 1668 865
rect 1166 862 1172 863
rect 1166 858 1167 862
rect 1171 858 1172 862
rect 1166 857 1172 858
rect 1230 862 1236 863
rect 1230 858 1231 862
rect 1235 858 1236 862
rect 1230 857 1236 858
rect 1286 862 1292 863
rect 1286 858 1287 862
rect 1291 858 1292 862
rect 1286 857 1292 858
rect 1342 862 1348 863
rect 1342 858 1343 862
rect 1347 858 1348 862
rect 1342 857 1348 858
rect 1398 862 1404 863
rect 1398 858 1399 862
rect 1403 858 1404 862
rect 1398 857 1404 858
rect 1462 862 1468 863
rect 1462 858 1463 862
rect 1467 858 1468 862
rect 1662 860 1663 864
rect 1667 860 1668 864
rect 1662 859 1668 860
rect 1462 857 1468 858
rect 1118 851 1124 852
rect 1118 847 1119 851
rect 1123 847 1124 851
rect 1118 846 1124 847
rect 1662 847 1668 848
rect 1102 845 1108 846
rect 1102 841 1103 845
rect 1107 841 1108 845
rect 1102 840 1108 841
rect 1166 845 1172 846
rect 1166 841 1167 845
rect 1171 841 1172 845
rect 1166 840 1172 841
rect 1230 845 1236 846
rect 1230 841 1231 845
rect 1235 841 1236 845
rect 1230 840 1236 841
rect 1286 845 1292 846
rect 1286 841 1287 845
rect 1291 841 1292 845
rect 1286 840 1292 841
rect 1342 845 1348 846
rect 1342 841 1343 845
rect 1347 841 1348 845
rect 1342 840 1348 841
rect 1398 845 1404 846
rect 1398 841 1399 845
rect 1403 841 1404 845
rect 1398 840 1404 841
rect 1462 845 1468 846
rect 1462 841 1463 845
rect 1467 841 1468 845
rect 1662 843 1663 847
rect 1667 843 1668 847
rect 1662 842 1668 843
rect 1462 840 1468 841
rect 1103 838 1107 840
rect 1103 833 1107 834
rect 1111 838 1115 839
rect 1111 832 1115 834
rect 1167 838 1171 840
rect 1167 833 1171 834
rect 1183 838 1187 839
rect 1183 832 1187 834
rect 1231 838 1235 840
rect 1231 833 1235 834
rect 1247 838 1251 839
rect 1247 832 1251 834
rect 1287 838 1291 840
rect 1330 839 1336 840
rect 1287 833 1291 834
rect 1311 838 1315 839
rect 1330 835 1331 839
rect 1335 835 1336 839
rect 1330 834 1336 835
rect 1343 838 1347 840
rect 1311 832 1315 834
rect 1110 831 1116 832
rect 1110 827 1111 831
rect 1115 827 1116 831
rect 1110 826 1116 827
rect 1182 831 1188 832
rect 1182 827 1183 831
rect 1187 827 1188 831
rect 1182 826 1188 827
rect 1246 831 1252 832
rect 1246 827 1247 831
rect 1251 827 1252 831
rect 1246 826 1252 827
rect 1310 831 1316 832
rect 1310 827 1311 831
rect 1315 827 1316 831
rect 1310 826 1316 827
rect 858 823 864 824
rect 858 819 859 823
rect 863 819 864 823
rect 858 818 864 819
rect 1054 823 1060 824
rect 1054 819 1055 823
rect 1059 819 1060 823
rect 1054 818 1060 819
rect 734 814 740 815
rect 734 810 735 814
rect 739 810 740 814
rect 734 809 740 810
rect 790 814 796 815
rect 790 810 791 814
rect 795 810 796 814
rect 790 809 796 810
rect 846 814 852 815
rect 846 810 847 814
rect 851 810 852 814
rect 846 809 852 810
rect 690 807 696 808
rect 690 803 691 807
rect 695 803 696 807
rect 690 802 696 803
rect 736 795 738 809
rect 792 795 794 809
rect 848 795 850 809
rect 860 796 862 818
rect 910 814 916 815
rect 910 810 911 814
rect 915 810 916 814
rect 910 809 916 810
rect 974 814 980 815
rect 974 810 975 814
rect 979 810 980 814
rect 974 809 980 810
rect 1038 814 1044 815
rect 1038 810 1039 814
rect 1043 810 1044 814
rect 1038 809 1044 810
rect 1110 814 1116 815
rect 1110 810 1111 814
rect 1115 810 1116 814
rect 1110 809 1116 810
rect 1182 814 1188 815
rect 1182 810 1183 814
rect 1187 810 1188 814
rect 1182 809 1188 810
rect 1246 814 1252 815
rect 1246 810 1247 814
rect 1251 810 1252 814
rect 1246 809 1252 810
rect 1310 814 1316 815
rect 1310 810 1311 814
rect 1315 810 1316 814
rect 1310 809 1316 810
rect 858 795 864 796
rect 912 795 914 809
rect 976 795 978 809
rect 1040 795 1042 809
rect 1112 795 1114 809
rect 1184 795 1186 809
rect 1248 795 1250 809
rect 1302 807 1308 808
rect 1302 803 1303 807
rect 1307 803 1308 807
rect 1302 802 1308 803
rect 543 794 547 795
rect 543 789 547 790
rect 607 794 611 795
rect 607 789 611 790
rect 615 794 619 795
rect 615 789 619 790
rect 671 794 675 795
rect 671 789 675 790
rect 703 794 707 795
rect 703 789 707 790
rect 735 794 739 795
rect 735 789 739 790
rect 791 794 795 795
rect 791 789 795 790
rect 847 794 851 795
rect 858 791 859 795
rect 863 791 864 795
rect 858 790 864 791
rect 871 794 875 795
rect 847 789 851 790
rect 871 789 875 790
rect 911 794 915 795
rect 911 789 915 790
rect 951 794 955 795
rect 951 789 955 790
rect 975 794 979 795
rect 975 789 979 790
rect 1023 794 1027 795
rect 1023 789 1027 790
rect 1039 794 1043 795
rect 1039 789 1043 790
rect 1095 794 1099 795
rect 1095 789 1099 790
rect 1111 794 1115 795
rect 1111 789 1115 790
rect 1167 794 1171 795
rect 1167 789 1171 790
rect 1183 794 1187 795
rect 1183 789 1187 790
rect 1231 794 1235 795
rect 1231 789 1235 790
rect 1247 794 1251 795
rect 1247 789 1251 790
rect 1295 794 1299 795
rect 1295 789 1299 790
rect 534 783 540 784
rect 534 779 535 783
rect 539 779 540 783
rect 616 779 618 789
rect 704 779 706 789
rect 792 779 794 789
rect 872 779 874 789
rect 952 779 954 789
rect 966 783 972 784
rect 966 779 967 783
rect 971 779 972 783
rect 1024 779 1026 789
rect 1096 779 1098 789
rect 1168 779 1170 789
rect 1232 779 1234 789
rect 1296 779 1298 789
rect 366 778 372 779
rect 366 774 367 778
rect 371 774 372 778
rect 366 773 372 774
rect 446 778 452 779
rect 446 774 447 778
rect 451 774 452 778
rect 446 773 452 774
rect 526 778 532 779
rect 534 778 540 779
rect 614 778 620 779
rect 526 774 527 778
rect 531 774 532 778
rect 526 773 532 774
rect 614 774 615 778
rect 619 774 620 778
rect 614 773 620 774
rect 702 778 708 779
rect 702 774 703 778
rect 707 774 708 778
rect 702 773 708 774
rect 790 778 796 779
rect 790 774 791 778
rect 795 774 796 778
rect 790 773 796 774
rect 870 778 876 779
rect 870 774 871 778
rect 875 774 876 778
rect 870 773 876 774
rect 950 778 956 779
rect 966 778 972 779
rect 1022 778 1028 779
rect 950 774 951 778
rect 955 774 956 778
rect 950 773 956 774
rect 350 767 356 768
rect 350 763 351 767
rect 355 763 356 767
rect 350 762 356 763
rect 686 767 692 768
rect 686 763 687 767
rect 691 763 692 767
rect 686 762 692 763
rect 882 767 888 768
rect 882 763 883 767
rect 887 763 888 767
rect 882 762 888 763
rect 366 761 372 762
rect 366 757 367 761
rect 371 757 372 761
rect 366 756 372 757
rect 446 761 452 762
rect 446 757 447 761
rect 451 757 452 761
rect 446 756 452 757
rect 526 761 532 762
rect 526 757 527 761
rect 531 757 532 761
rect 526 756 532 757
rect 614 761 620 762
rect 614 757 615 761
rect 619 757 620 761
rect 614 756 620 757
rect 319 754 323 755
rect 319 748 323 750
rect 359 754 363 755
rect 359 748 363 750
rect 367 754 371 756
rect 367 749 371 750
rect 399 754 403 755
rect 399 748 403 750
rect 439 754 443 755
rect 439 748 443 750
rect 447 754 451 756
rect 447 749 451 750
rect 487 754 491 755
rect 487 748 491 750
rect 527 754 531 756
rect 527 749 531 750
rect 543 754 547 755
rect 543 748 547 750
rect 607 754 611 755
rect 607 748 611 750
rect 615 754 619 756
rect 615 749 619 750
rect 671 754 675 755
rect 671 748 675 750
rect 318 747 324 748
rect 278 742 284 743
rect 306 743 312 744
rect 110 740 116 741
rect 306 739 307 743
rect 311 739 312 743
rect 318 743 319 747
rect 323 743 324 747
rect 318 742 324 743
rect 358 747 364 748
rect 358 743 359 747
rect 363 743 364 747
rect 358 742 364 743
rect 398 747 404 748
rect 398 743 399 747
rect 403 743 404 747
rect 398 742 404 743
rect 438 747 444 748
rect 438 743 439 747
rect 443 743 444 747
rect 438 742 444 743
rect 486 747 492 748
rect 486 743 487 747
rect 491 743 492 747
rect 486 742 492 743
rect 542 747 548 748
rect 542 743 543 747
rect 547 743 548 747
rect 542 742 548 743
rect 606 747 612 748
rect 606 743 607 747
rect 611 743 612 747
rect 606 742 612 743
rect 670 747 676 748
rect 670 743 671 747
rect 675 743 676 747
rect 670 742 676 743
rect 306 738 312 739
rect 330 739 336 740
rect 330 735 331 739
rect 335 735 336 739
rect 330 734 336 735
rect 414 739 420 740
rect 414 735 415 739
rect 419 735 420 739
rect 414 734 420 735
rect 214 730 220 731
rect 110 728 116 729
rect 110 724 111 728
rect 115 724 116 728
rect 214 726 215 730
rect 219 726 220 730
rect 214 725 220 726
rect 246 730 252 731
rect 246 726 247 730
rect 251 726 252 730
rect 246 725 252 726
rect 278 730 284 731
rect 278 726 279 730
rect 283 726 284 730
rect 278 725 284 726
rect 318 730 324 731
rect 318 726 319 730
rect 323 726 324 730
rect 318 725 324 726
rect 110 723 116 724
rect 112 711 114 723
rect 216 711 218 725
rect 248 711 250 725
rect 280 711 282 725
rect 320 711 322 725
rect 332 716 334 734
rect 358 730 364 731
rect 358 726 359 730
rect 363 726 364 730
rect 358 725 364 726
rect 398 730 404 731
rect 398 726 399 730
rect 403 726 404 730
rect 398 725 404 726
rect 330 715 336 716
rect 330 711 331 715
rect 335 711 336 715
rect 360 711 362 725
rect 366 723 372 724
rect 366 719 367 723
rect 371 719 372 723
rect 366 718 372 719
rect 111 710 115 711
rect 111 705 115 706
rect 215 710 219 711
rect 215 705 219 706
rect 247 710 251 711
rect 247 705 251 706
rect 279 710 283 711
rect 279 705 283 706
rect 311 710 315 711
rect 311 705 315 706
rect 319 710 323 711
rect 330 710 336 711
rect 343 710 347 711
rect 319 705 323 706
rect 343 705 347 706
rect 359 710 363 711
rect 359 705 363 706
rect 112 697 114 705
rect 110 696 116 697
rect 110 692 111 696
rect 115 692 116 696
rect 280 695 282 705
rect 312 695 314 705
rect 344 695 346 705
rect 110 691 116 692
rect 278 694 284 695
rect 278 690 279 694
rect 283 690 284 694
rect 278 689 284 690
rect 310 694 316 695
rect 310 690 311 694
rect 315 690 316 694
rect 310 689 316 690
rect 342 694 348 695
rect 342 690 343 694
rect 347 690 348 694
rect 342 689 348 690
rect 359 683 365 684
rect 110 679 116 680
rect 110 675 111 679
rect 115 675 116 679
rect 359 679 360 683
rect 364 682 365 683
rect 368 682 370 718
rect 400 711 402 725
rect 416 716 418 734
rect 438 730 444 731
rect 438 726 439 730
rect 443 726 444 730
rect 438 725 444 726
rect 486 730 492 731
rect 486 726 487 730
rect 491 726 492 730
rect 486 725 492 726
rect 542 730 548 731
rect 542 726 543 730
rect 547 726 548 730
rect 542 725 548 726
rect 606 730 612 731
rect 606 726 607 730
rect 611 726 612 730
rect 606 725 612 726
rect 670 730 676 731
rect 670 726 671 730
rect 675 726 676 730
rect 670 725 676 726
rect 414 715 420 716
rect 414 711 415 715
rect 419 711 420 715
rect 440 711 442 725
rect 488 711 490 725
rect 544 711 546 725
rect 608 711 610 725
rect 672 711 674 725
rect 688 724 690 762
rect 702 761 708 762
rect 702 757 703 761
rect 707 757 708 761
rect 702 756 708 757
rect 790 761 796 762
rect 790 757 791 761
rect 795 757 796 761
rect 790 756 796 757
rect 870 761 876 762
rect 870 757 871 761
rect 875 757 876 761
rect 870 756 876 757
rect 703 754 707 756
rect 703 749 707 750
rect 735 754 739 755
rect 735 748 739 750
rect 791 754 795 756
rect 791 749 795 750
rect 799 754 803 755
rect 799 748 803 750
rect 863 754 867 755
rect 863 748 867 750
rect 871 754 875 756
rect 871 749 875 750
rect 734 747 740 748
rect 734 743 735 747
rect 739 743 740 747
rect 734 742 740 743
rect 798 747 804 748
rect 798 743 799 747
rect 803 743 804 747
rect 798 742 804 743
rect 862 747 868 748
rect 862 743 863 747
rect 867 743 868 747
rect 862 742 868 743
rect 774 739 780 740
rect 774 735 775 739
rect 779 735 780 739
rect 774 734 780 735
rect 734 730 740 731
rect 734 726 735 730
rect 739 726 740 730
rect 734 725 740 726
rect 686 723 692 724
rect 686 719 687 723
rect 691 719 692 723
rect 686 718 692 719
rect 736 711 738 725
rect 375 710 379 711
rect 399 710 403 711
rect 375 705 379 706
rect 390 707 396 708
rect 376 695 378 705
rect 390 703 391 707
rect 395 703 396 707
rect 399 705 403 706
rect 407 710 411 711
rect 414 710 420 711
rect 439 710 443 711
rect 407 705 411 706
rect 439 705 443 706
rect 471 710 475 711
rect 471 705 475 706
rect 487 710 491 711
rect 487 705 491 706
rect 503 710 507 711
rect 503 705 507 706
rect 543 710 547 711
rect 543 705 547 706
rect 591 710 595 711
rect 591 705 595 706
rect 607 710 611 711
rect 607 705 611 706
rect 647 710 651 711
rect 647 705 651 706
rect 671 710 675 711
rect 671 705 675 706
rect 703 710 707 711
rect 703 705 707 706
rect 735 710 739 711
rect 735 705 739 706
rect 759 710 763 711
rect 759 705 763 706
rect 390 702 396 703
rect 374 694 380 695
rect 374 690 375 694
rect 379 690 380 694
rect 374 689 380 690
rect 392 684 394 702
rect 408 695 410 705
rect 440 695 442 705
rect 472 695 474 705
rect 504 695 506 705
rect 544 695 546 705
rect 592 695 594 705
rect 648 695 650 705
rect 704 695 706 705
rect 760 695 762 705
rect 776 700 778 734
rect 798 730 804 731
rect 798 726 799 730
rect 803 726 804 730
rect 798 725 804 726
rect 862 730 868 731
rect 862 726 863 730
rect 867 726 868 730
rect 862 725 868 726
rect 800 711 802 725
rect 864 711 866 725
rect 884 724 886 762
rect 950 761 956 762
rect 950 757 951 761
rect 955 757 956 761
rect 950 756 956 757
rect 968 756 970 778
rect 1022 774 1023 778
rect 1027 774 1028 778
rect 1022 773 1028 774
rect 1094 778 1100 779
rect 1094 774 1095 778
rect 1099 774 1100 778
rect 1094 773 1100 774
rect 1166 778 1172 779
rect 1166 774 1167 778
rect 1171 774 1172 778
rect 1166 773 1172 774
rect 1230 778 1236 779
rect 1230 774 1231 778
rect 1235 774 1236 778
rect 1230 773 1236 774
rect 1294 778 1300 779
rect 1294 774 1295 778
rect 1299 774 1300 778
rect 1294 773 1300 774
rect 1304 768 1306 802
rect 1312 795 1314 809
rect 1332 808 1334 834
rect 1343 833 1347 834
rect 1367 838 1371 839
rect 1367 832 1371 834
rect 1399 838 1403 840
rect 1399 833 1403 834
rect 1423 838 1427 839
rect 1423 832 1427 834
rect 1463 838 1467 840
rect 1664 839 1666 842
rect 1463 833 1467 834
rect 1479 838 1483 839
rect 1479 832 1483 834
rect 1535 838 1539 839
rect 1535 832 1539 834
rect 1591 838 1595 839
rect 1591 832 1595 834
rect 1663 838 1667 839
rect 1663 833 1667 834
rect 1366 831 1372 832
rect 1366 827 1367 831
rect 1371 827 1372 831
rect 1366 826 1372 827
rect 1422 831 1428 832
rect 1422 827 1423 831
rect 1427 827 1428 831
rect 1422 826 1428 827
rect 1478 831 1484 832
rect 1478 827 1479 831
rect 1483 827 1484 831
rect 1478 826 1484 827
rect 1534 831 1540 832
rect 1534 827 1535 831
rect 1539 827 1540 831
rect 1534 826 1540 827
rect 1590 831 1596 832
rect 1590 827 1591 831
rect 1595 827 1596 831
rect 1664 830 1666 833
rect 1590 826 1596 827
rect 1662 829 1668 830
rect 1662 825 1663 829
rect 1667 825 1668 829
rect 1662 824 1668 825
rect 1606 823 1612 824
rect 1606 819 1607 823
rect 1611 819 1612 823
rect 1606 818 1612 819
rect 1366 814 1372 815
rect 1366 810 1367 814
rect 1371 810 1372 814
rect 1366 809 1372 810
rect 1422 814 1428 815
rect 1422 810 1423 814
rect 1427 810 1428 814
rect 1422 809 1428 810
rect 1478 814 1484 815
rect 1478 810 1479 814
rect 1483 810 1484 814
rect 1478 809 1484 810
rect 1534 814 1540 815
rect 1534 810 1535 814
rect 1539 810 1540 814
rect 1534 809 1540 810
rect 1590 814 1596 815
rect 1590 810 1591 814
rect 1595 810 1596 814
rect 1590 809 1596 810
rect 1330 807 1336 808
rect 1330 803 1331 807
rect 1335 803 1336 807
rect 1330 802 1336 803
rect 1368 795 1370 809
rect 1424 795 1426 809
rect 1480 795 1482 809
rect 1536 795 1538 809
rect 1592 795 1594 809
rect 1311 794 1315 795
rect 1311 789 1315 790
rect 1359 794 1363 795
rect 1359 789 1363 790
rect 1367 794 1371 795
rect 1367 789 1371 790
rect 1415 794 1419 795
rect 1415 789 1419 790
rect 1423 794 1427 795
rect 1423 789 1427 790
rect 1471 794 1475 795
rect 1471 789 1475 790
rect 1479 794 1483 795
rect 1479 789 1483 790
rect 1527 794 1531 795
rect 1527 789 1531 790
rect 1535 794 1539 795
rect 1535 789 1539 790
rect 1591 794 1595 795
rect 1591 789 1595 790
rect 1360 779 1362 789
rect 1374 783 1380 784
rect 1374 779 1375 783
rect 1379 779 1380 783
rect 1416 779 1418 789
rect 1472 779 1474 789
rect 1528 779 1530 789
rect 1592 779 1594 789
rect 1608 784 1610 818
rect 1662 812 1668 813
rect 1662 808 1663 812
rect 1667 808 1668 812
rect 1662 807 1668 808
rect 1664 795 1666 807
rect 1663 794 1667 795
rect 1663 789 1667 790
rect 1606 783 1612 784
rect 1606 779 1607 783
rect 1611 779 1612 783
rect 1664 781 1666 789
rect 1358 778 1364 779
rect 1374 778 1380 779
rect 1414 778 1420 779
rect 1358 774 1359 778
rect 1363 774 1364 778
rect 1358 773 1364 774
rect 1304 767 1312 768
rect 1304 764 1307 767
rect 1306 763 1307 764
rect 1311 763 1312 767
rect 1306 762 1312 763
rect 1022 761 1028 762
rect 1022 757 1023 761
rect 1027 757 1028 761
rect 1022 756 1028 757
rect 1094 761 1100 762
rect 1094 757 1095 761
rect 1099 757 1100 761
rect 1094 756 1100 757
rect 1166 761 1172 762
rect 1166 757 1167 761
rect 1171 757 1172 761
rect 1166 756 1172 757
rect 1230 761 1236 762
rect 1230 757 1231 761
rect 1235 757 1236 761
rect 1230 756 1236 757
rect 1294 761 1300 762
rect 1294 757 1295 761
rect 1299 757 1300 761
rect 1294 756 1300 757
rect 1358 761 1364 762
rect 1358 757 1359 761
rect 1363 757 1364 761
rect 1358 756 1364 757
rect 1376 756 1378 778
rect 1414 774 1415 778
rect 1419 774 1420 778
rect 1414 773 1420 774
rect 1470 778 1476 779
rect 1470 774 1471 778
rect 1475 774 1476 778
rect 1470 773 1476 774
rect 1526 778 1532 779
rect 1526 774 1527 778
rect 1531 774 1532 778
rect 1526 773 1532 774
rect 1590 778 1596 779
rect 1606 778 1612 779
rect 1662 780 1668 781
rect 1590 774 1591 778
rect 1595 774 1596 778
rect 1662 776 1663 780
rect 1667 776 1668 780
rect 1662 775 1668 776
rect 1590 773 1596 774
rect 1510 767 1516 768
rect 1510 763 1511 767
rect 1515 763 1516 767
rect 1510 762 1516 763
rect 1662 763 1668 764
rect 1414 761 1420 762
rect 1414 757 1415 761
rect 1419 757 1420 761
rect 1414 756 1420 757
rect 1470 761 1476 762
rect 1470 757 1471 761
rect 1475 757 1476 761
rect 1470 756 1476 757
rect 927 754 931 755
rect 927 748 931 750
rect 951 754 955 756
rect 966 755 972 756
rect 966 751 967 755
rect 971 751 972 755
rect 966 750 972 751
rect 991 754 995 755
rect 951 749 955 750
rect 991 748 995 750
rect 1023 754 1027 756
rect 1023 749 1027 750
rect 1055 754 1059 755
rect 1055 748 1059 750
rect 1095 754 1099 756
rect 1095 749 1099 750
rect 1119 754 1123 755
rect 1119 748 1123 750
rect 1167 754 1171 756
rect 1167 749 1171 750
rect 1183 754 1187 755
rect 1183 748 1187 750
rect 1231 754 1235 756
rect 1231 749 1235 750
rect 1239 754 1243 755
rect 1239 748 1243 750
rect 1295 754 1299 756
rect 1295 748 1299 750
rect 1351 754 1355 755
rect 1351 748 1355 750
rect 1359 754 1363 756
rect 1374 755 1380 756
rect 1374 751 1375 755
rect 1379 751 1380 755
rect 1374 750 1380 751
rect 1407 754 1411 755
rect 1359 749 1363 750
rect 1407 748 1411 750
rect 1415 754 1419 756
rect 1415 749 1419 750
rect 1463 754 1467 755
rect 1463 748 1467 750
rect 1471 754 1475 756
rect 1471 749 1475 750
rect 926 747 932 748
rect 926 743 927 747
rect 931 743 932 747
rect 926 742 932 743
rect 990 747 996 748
rect 990 743 991 747
rect 995 743 996 747
rect 990 742 996 743
rect 1054 747 1060 748
rect 1054 743 1055 747
rect 1059 743 1060 747
rect 1054 742 1060 743
rect 1118 747 1124 748
rect 1118 743 1119 747
rect 1123 743 1124 747
rect 1118 742 1124 743
rect 1182 747 1188 748
rect 1182 743 1183 747
rect 1187 743 1188 747
rect 1182 742 1188 743
rect 1238 747 1244 748
rect 1238 743 1239 747
rect 1243 743 1244 747
rect 1238 742 1244 743
rect 1294 747 1300 748
rect 1294 743 1295 747
rect 1299 743 1300 747
rect 1294 742 1300 743
rect 1350 747 1356 748
rect 1350 743 1351 747
rect 1355 743 1356 747
rect 1350 742 1356 743
rect 1406 747 1412 748
rect 1406 743 1407 747
rect 1411 743 1412 747
rect 1406 742 1412 743
rect 1462 747 1468 748
rect 1462 743 1463 747
rect 1467 743 1468 747
rect 1462 742 1468 743
rect 926 730 932 731
rect 926 726 927 730
rect 931 726 932 730
rect 926 725 932 726
rect 990 730 996 731
rect 990 726 991 730
rect 995 726 996 730
rect 990 725 996 726
rect 1054 730 1060 731
rect 1054 726 1055 730
rect 1059 726 1060 730
rect 1054 725 1060 726
rect 1118 730 1124 731
rect 1118 726 1119 730
rect 1123 726 1124 730
rect 1118 725 1124 726
rect 1182 730 1188 731
rect 1182 726 1183 730
rect 1187 726 1188 730
rect 1182 725 1188 726
rect 1238 730 1244 731
rect 1238 726 1239 730
rect 1243 726 1244 730
rect 1238 725 1244 726
rect 1294 730 1300 731
rect 1294 726 1295 730
rect 1299 726 1300 730
rect 1294 725 1300 726
rect 1350 730 1356 731
rect 1350 726 1351 730
rect 1355 726 1356 730
rect 1350 725 1356 726
rect 1406 730 1412 731
rect 1406 726 1407 730
rect 1411 726 1412 730
rect 1406 725 1412 726
rect 1462 730 1468 731
rect 1462 726 1463 730
rect 1467 726 1468 730
rect 1462 725 1468 726
rect 882 723 888 724
rect 882 719 883 723
rect 887 719 888 723
rect 882 718 888 719
rect 928 711 930 725
rect 974 723 980 724
rect 974 719 975 723
rect 979 719 980 723
rect 974 718 980 719
rect 799 710 803 711
rect 799 705 803 706
rect 823 710 827 711
rect 823 705 827 706
rect 863 710 867 711
rect 863 705 867 706
rect 887 710 891 711
rect 887 705 891 706
rect 927 710 931 711
rect 927 705 931 706
rect 959 710 963 711
rect 959 705 963 706
rect 774 699 780 700
rect 774 695 775 699
rect 779 695 780 699
rect 824 695 826 705
rect 888 695 890 705
rect 960 695 962 705
rect 406 694 412 695
rect 406 690 407 694
rect 411 690 412 694
rect 406 689 412 690
rect 438 694 444 695
rect 438 690 439 694
rect 443 690 444 694
rect 438 689 444 690
rect 470 694 476 695
rect 470 690 471 694
rect 475 690 476 694
rect 470 689 476 690
rect 502 694 508 695
rect 502 690 503 694
rect 507 690 508 694
rect 502 689 508 690
rect 542 694 548 695
rect 542 690 543 694
rect 547 690 548 694
rect 542 689 548 690
rect 590 694 596 695
rect 590 690 591 694
rect 595 690 596 694
rect 590 689 596 690
rect 646 694 652 695
rect 646 690 647 694
rect 651 690 652 694
rect 646 689 652 690
rect 702 694 708 695
rect 702 690 703 694
rect 707 690 708 694
rect 702 689 708 690
rect 758 694 764 695
rect 774 694 780 695
rect 822 694 828 695
rect 758 690 759 694
rect 763 690 764 694
rect 758 689 764 690
rect 822 690 823 694
rect 827 690 828 694
rect 822 689 828 690
rect 886 694 892 695
rect 886 690 887 694
rect 891 690 892 694
rect 886 689 892 690
rect 958 694 964 695
rect 958 690 959 694
rect 963 690 964 694
rect 958 689 964 690
rect 976 684 978 718
rect 992 711 994 725
rect 1056 711 1058 725
rect 1102 711 1108 712
rect 1120 711 1122 725
rect 1184 711 1186 725
rect 1240 711 1242 725
rect 1296 711 1298 725
rect 1352 711 1354 725
rect 1408 711 1410 725
rect 1464 711 1466 725
rect 1512 724 1514 762
rect 1526 761 1532 762
rect 1526 757 1527 761
rect 1531 757 1532 761
rect 1526 756 1532 757
rect 1590 761 1596 762
rect 1590 757 1591 761
rect 1595 757 1596 761
rect 1662 759 1663 763
rect 1667 759 1668 763
rect 1662 758 1668 759
rect 1590 756 1596 757
rect 1519 754 1523 755
rect 1519 748 1523 750
rect 1527 754 1531 756
rect 1527 749 1531 750
rect 1583 754 1587 755
rect 1583 748 1587 750
rect 1591 754 1595 756
rect 1664 755 1666 758
rect 1591 749 1595 750
rect 1623 754 1627 755
rect 1623 748 1627 750
rect 1663 754 1667 755
rect 1663 749 1667 750
rect 1518 747 1524 748
rect 1518 743 1519 747
rect 1523 743 1524 747
rect 1518 742 1524 743
rect 1582 747 1588 748
rect 1582 743 1583 747
rect 1587 743 1588 747
rect 1582 742 1588 743
rect 1622 747 1628 748
rect 1622 743 1623 747
rect 1627 743 1628 747
rect 1664 746 1666 749
rect 1622 742 1628 743
rect 1662 745 1668 746
rect 1662 741 1663 745
rect 1667 741 1668 745
rect 1662 740 1668 741
rect 1638 739 1644 740
rect 1638 735 1639 739
rect 1643 735 1644 739
rect 1638 734 1644 735
rect 1518 730 1524 731
rect 1518 726 1519 730
rect 1523 726 1524 730
rect 1518 725 1524 726
rect 1582 730 1588 731
rect 1582 726 1583 730
rect 1587 726 1588 730
rect 1582 725 1588 726
rect 1622 730 1628 731
rect 1622 726 1623 730
rect 1627 726 1628 730
rect 1622 725 1628 726
rect 1510 723 1516 724
rect 1510 719 1511 723
rect 1515 719 1516 723
rect 1510 718 1516 719
rect 1520 711 1522 725
rect 1546 723 1552 724
rect 1546 719 1547 723
rect 1551 719 1552 723
rect 1546 718 1552 719
rect 991 710 995 711
rect 991 705 995 706
rect 1023 710 1027 711
rect 1023 705 1027 706
rect 1055 710 1059 711
rect 1055 705 1059 706
rect 1087 710 1091 711
rect 1102 707 1103 711
rect 1107 707 1108 711
rect 1102 706 1108 707
rect 1119 710 1123 711
rect 1087 705 1091 706
rect 1024 695 1026 705
rect 1030 699 1036 700
rect 1030 695 1031 699
rect 1035 695 1036 699
rect 1088 695 1090 705
rect 1022 694 1028 695
rect 1030 694 1036 695
rect 1086 694 1092 695
rect 1022 690 1023 694
rect 1027 690 1028 694
rect 1022 689 1028 690
rect 364 680 370 682
rect 390 683 396 684
rect 364 679 365 680
rect 359 678 365 679
rect 390 679 391 683
rect 395 679 396 683
rect 390 678 396 679
rect 926 683 932 684
rect 926 679 927 683
rect 931 679 932 683
rect 926 678 932 679
rect 974 683 980 684
rect 974 679 975 683
rect 979 679 980 683
rect 974 678 980 679
rect 110 674 116 675
rect 278 677 284 678
rect 112 671 114 674
rect 278 673 279 677
rect 283 673 284 677
rect 278 672 284 673
rect 310 677 316 678
rect 310 673 311 677
rect 315 673 316 677
rect 310 672 316 673
rect 342 677 348 678
rect 342 673 343 677
rect 347 673 348 677
rect 342 672 348 673
rect 374 677 380 678
rect 374 673 375 677
rect 379 673 380 677
rect 374 672 380 673
rect 406 677 412 678
rect 406 673 407 677
rect 411 673 412 677
rect 406 672 412 673
rect 438 677 444 678
rect 438 673 439 677
rect 443 673 444 677
rect 438 672 444 673
rect 470 677 476 678
rect 470 673 471 677
rect 475 673 476 677
rect 470 672 476 673
rect 502 677 508 678
rect 502 673 503 677
rect 507 673 508 677
rect 502 672 508 673
rect 542 677 548 678
rect 542 673 543 677
rect 547 673 548 677
rect 542 672 548 673
rect 590 677 596 678
rect 590 673 591 677
rect 595 673 596 677
rect 590 672 596 673
rect 646 677 652 678
rect 646 673 647 677
rect 651 673 652 677
rect 646 672 652 673
rect 702 677 708 678
rect 702 673 703 677
rect 707 673 708 677
rect 702 672 708 673
rect 758 677 764 678
rect 758 673 759 677
rect 763 673 764 677
rect 758 672 764 673
rect 822 677 828 678
rect 822 673 823 677
rect 827 673 828 677
rect 822 672 828 673
rect 886 677 892 678
rect 886 673 887 677
rect 891 673 892 677
rect 886 672 892 673
rect 111 670 115 671
rect 111 665 115 666
rect 279 670 283 672
rect 279 665 283 666
rect 295 670 299 671
rect 112 662 114 665
rect 295 664 299 666
rect 311 670 315 672
rect 311 665 315 666
rect 327 670 331 671
rect 327 664 331 666
rect 343 670 347 672
rect 343 665 347 666
rect 359 670 363 671
rect 359 664 363 666
rect 375 670 379 672
rect 375 665 379 666
rect 391 670 395 671
rect 391 664 395 666
rect 407 670 411 672
rect 407 665 411 666
rect 423 670 427 671
rect 423 664 427 666
rect 439 670 443 672
rect 439 665 443 666
rect 455 670 459 671
rect 455 664 459 666
rect 471 670 475 672
rect 471 665 475 666
rect 487 670 491 671
rect 487 664 491 666
rect 503 670 507 672
rect 534 671 540 672
rect 503 665 507 666
rect 519 670 523 671
rect 534 667 535 671
rect 539 667 540 671
rect 534 666 540 667
rect 543 670 547 672
rect 519 664 523 666
rect 294 663 300 664
rect 110 661 116 662
rect 110 657 111 661
rect 115 657 116 661
rect 294 659 295 663
rect 299 659 300 663
rect 294 658 300 659
rect 326 663 332 664
rect 326 659 327 663
rect 331 659 332 663
rect 326 658 332 659
rect 358 663 364 664
rect 358 659 359 663
rect 363 659 364 663
rect 358 658 364 659
rect 390 663 396 664
rect 390 659 391 663
rect 395 659 396 663
rect 390 658 396 659
rect 422 663 428 664
rect 422 659 423 663
rect 427 659 428 663
rect 422 658 428 659
rect 454 663 460 664
rect 454 659 455 663
rect 459 659 460 663
rect 454 658 460 659
rect 486 663 492 664
rect 486 659 487 663
rect 491 659 492 663
rect 486 658 492 659
rect 518 663 524 664
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 110 656 116 657
rect 294 646 300 647
rect 110 644 116 645
rect 110 640 111 644
rect 115 640 116 644
rect 294 642 295 646
rect 299 642 300 646
rect 294 641 300 642
rect 326 646 332 647
rect 326 642 327 646
rect 331 642 332 646
rect 326 641 332 642
rect 358 646 364 647
rect 358 642 359 646
rect 363 642 364 646
rect 358 641 364 642
rect 390 646 396 647
rect 390 642 391 646
rect 395 642 396 646
rect 390 641 396 642
rect 422 646 428 647
rect 422 642 423 646
rect 427 642 428 646
rect 422 641 428 642
rect 454 646 460 647
rect 454 642 455 646
rect 459 642 460 646
rect 454 641 460 642
rect 486 646 492 647
rect 486 642 487 646
rect 491 642 492 646
rect 486 641 492 642
rect 518 646 524 647
rect 518 642 519 646
rect 523 642 524 646
rect 518 641 524 642
rect 110 639 116 640
rect 112 631 114 639
rect 296 631 298 641
rect 328 631 330 641
rect 360 631 362 641
rect 392 631 394 641
rect 424 631 426 641
rect 456 631 458 641
rect 478 631 484 632
rect 488 631 490 641
rect 520 631 522 641
rect 536 640 538 666
rect 543 665 547 666
rect 551 670 555 671
rect 551 664 555 666
rect 591 670 595 672
rect 591 664 595 666
rect 639 670 643 671
rect 639 664 643 666
rect 647 670 651 672
rect 647 665 651 666
rect 687 670 691 671
rect 687 664 691 666
rect 703 670 707 672
rect 703 665 707 666
rect 735 670 739 671
rect 735 664 739 666
rect 759 670 763 672
rect 759 665 763 666
rect 791 670 795 671
rect 791 664 795 666
rect 823 670 827 672
rect 823 665 827 666
rect 847 670 851 671
rect 847 664 851 666
rect 887 670 891 672
rect 887 665 891 666
rect 911 670 915 671
rect 911 664 915 666
rect 550 663 556 664
rect 550 659 551 663
rect 555 659 556 663
rect 550 658 556 659
rect 590 663 596 664
rect 590 659 591 663
rect 595 659 596 663
rect 590 658 596 659
rect 638 663 644 664
rect 638 659 639 663
rect 643 659 644 663
rect 638 658 644 659
rect 686 663 692 664
rect 686 659 687 663
rect 691 659 692 663
rect 686 658 692 659
rect 734 663 740 664
rect 734 659 735 663
rect 739 659 740 663
rect 734 658 740 659
rect 790 663 796 664
rect 790 659 791 663
rect 795 659 796 663
rect 790 658 796 659
rect 846 663 852 664
rect 846 659 847 663
rect 851 659 852 663
rect 846 658 852 659
rect 910 663 916 664
rect 910 659 911 663
rect 915 659 916 663
rect 910 658 916 659
rect 750 655 756 656
rect 750 651 751 655
rect 755 651 756 655
rect 750 650 756 651
rect 838 655 844 656
rect 838 651 839 655
rect 843 651 844 655
rect 838 650 844 651
rect 550 646 556 647
rect 550 642 551 646
rect 555 642 556 646
rect 550 641 556 642
rect 590 646 596 647
rect 590 642 591 646
rect 595 642 596 646
rect 590 641 596 642
rect 638 646 644 647
rect 638 642 639 646
rect 643 642 644 646
rect 638 641 644 642
rect 686 646 692 647
rect 686 642 687 646
rect 691 642 692 646
rect 686 641 692 642
rect 734 646 740 647
rect 734 642 735 646
rect 739 642 740 646
rect 734 641 740 642
rect 534 639 540 640
rect 534 635 535 639
rect 539 635 540 639
rect 534 634 540 635
rect 552 631 554 641
rect 592 631 594 641
rect 640 631 642 641
rect 688 631 690 641
rect 736 631 738 641
rect 752 632 754 650
rect 790 646 796 647
rect 790 642 791 646
rect 795 642 796 646
rect 790 641 796 642
rect 750 631 756 632
rect 792 631 794 641
rect 111 630 115 631
rect 111 625 115 626
rect 247 630 251 631
rect 247 625 251 626
rect 279 630 283 631
rect 279 625 283 626
rect 295 630 299 631
rect 295 625 299 626
rect 319 630 323 631
rect 319 625 323 626
rect 327 630 331 631
rect 327 625 331 626
rect 359 630 363 631
rect 359 625 363 626
rect 367 630 371 631
rect 367 625 371 626
rect 391 630 395 631
rect 391 625 395 626
rect 423 630 427 631
rect 423 625 427 626
rect 455 630 459 631
rect 455 625 459 626
rect 471 630 475 631
rect 478 627 479 631
rect 483 627 484 631
rect 478 626 484 627
rect 487 630 491 631
rect 471 625 475 626
rect 112 617 114 625
rect 110 616 116 617
rect 110 612 111 616
rect 115 612 116 616
rect 248 615 250 625
rect 262 619 268 620
rect 262 615 263 619
rect 267 615 268 619
rect 280 615 282 625
rect 320 615 322 625
rect 368 615 370 625
rect 424 615 426 625
rect 472 615 474 625
rect 110 611 116 612
rect 246 614 252 615
rect 262 614 268 615
rect 278 614 284 615
rect 246 610 247 614
rect 251 610 252 614
rect 246 609 252 610
rect 110 599 116 600
rect 110 595 111 599
rect 115 595 116 599
rect 110 594 116 595
rect 246 597 252 598
rect 112 591 114 594
rect 246 593 247 597
rect 251 593 252 597
rect 246 592 252 593
rect 264 592 266 614
rect 278 610 279 614
rect 283 610 284 614
rect 278 609 284 610
rect 318 614 324 615
rect 318 610 319 614
rect 323 610 324 614
rect 318 609 324 610
rect 366 614 372 615
rect 366 610 367 614
rect 371 610 372 614
rect 366 609 372 610
rect 422 614 428 615
rect 422 610 423 614
rect 427 610 428 614
rect 422 609 428 610
rect 470 614 476 615
rect 470 610 471 614
rect 475 610 476 614
rect 470 609 476 610
rect 480 604 482 626
rect 487 625 491 626
rect 519 630 523 631
rect 519 625 523 626
rect 551 630 555 631
rect 551 625 555 626
rect 567 630 571 631
rect 567 625 571 626
rect 591 630 595 631
rect 591 625 595 626
rect 615 630 619 631
rect 615 625 619 626
rect 639 630 643 631
rect 639 625 643 626
rect 663 630 667 631
rect 663 625 667 626
rect 687 630 691 631
rect 687 625 691 626
rect 719 630 723 631
rect 719 625 723 626
rect 735 630 739 631
rect 750 627 751 631
rect 755 627 756 631
rect 750 626 756 627
rect 775 630 779 631
rect 735 625 739 626
rect 775 625 779 626
rect 791 630 795 631
rect 791 625 795 626
rect 831 630 835 631
rect 831 625 835 626
rect 520 615 522 625
rect 568 615 570 625
rect 616 615 618 625
rect 664 615 666 625
rect 720 615 722 625
rect 776 615 778 625
rect 832 615 834 625
rect 840 620 842 650
rect 846 646 852 647
rect 846 642 847 646
rect 851 642 852 646
rect 846 641 852 642
rect 910 646 916 647
rect 910 642 911 646
rect 915 642 916 646
rect 910 641 916 642
rect 848 631 850 641
rect 912 631 914 641
rect 928 640 930 678
rect 958 677 964 678
rect 958 673 959 677
rect 963 673 964 677
rect 958 672 964 673
rect 1022 677 1028 678
rect 1022 673 1023 677
rect 1027 673 1028 677
rect 1022 672 1028 673
rect 959 670 963 672
rect 959 665 963 666
rect 975 670 979 671
rect 975 664 979 666
rect 1023 670 1027 672
rect 1023 665 1027 666
rect 974 663 980 664
rect 974 659 975 663
rect 979 659 980 663
rect 974 658 980 659
rect 1032 656 1034 694
rect 1086 690 1087 694
rect 1091 690 1092 694
rect 1086 689 1092 690
rect 1104 684 1106 706
rect 1119 705 1123 706
rect 1159 710 1163 711
rect 1159 705 1163 706
rect 1183 710 1187 711
rect 1183 705 1187 706
rect 1223 710 1227 711
rect 1223 705 1227 706
rect 1239 710 1243 711
rect 1239 705 1243 706
rect 1287 710 1291 711
rect 1287 705 1291 706
rect 1295 710 1299 711
rect 1295 705 1299 706
rect 1351 710 1355 711
rect 1351 705 1355 706
rect 1407 710 1411 711
rect 1407 705 1411 706
rect 1415 710 1419 711
rect 1415 705 1419 706
rect 1463 710 1467 711
rect 1463 705 1467 706
rect 1471 710 1475 711
rect 1471 705 1475 706
rect 1519 710 1523 711
rect 1519 705 1523 706
rect 1527 710 1531 711
rect 1527 705 1531 706
rect 1160 695 1162 705
rect 1224 695 1226 705
rect 1288 695 1290 705
rect 1352 695 1354 705
rect 1416 695 1418 705
rect 1472 695 1474 705
rect 1486 699 1492 700
rect 1486 695 1487 699
rect 1491 695 1492 699
rect 1528 695 1530 705
rect 1158 694 1164 695
rect 1158 690 1159 694
rect 1163 690 1164 694
rect 1158 689 1164 690
rect 1222 694 1228 695
rect 1222 690 1223 694
rect 1227 690 1228 694
rect 1222 689 1228 690
rect 1286 694 1292 695
rect 1286 690 1287 694
rect 1291 690 1292 694
rect 1286 689 1292 690
rect 1350 694 1356 695
rect 1350 690 1351 694
rect 1355 690 1356 694
rect 1350 689 1356 690
rect 1414 694 1420 695
rect 1414 690 1415 694
rect 1419 690 1420 694
rect 1414 689 1420 690
rect 1470 694 1476 695
rect 1486 694 1492 695
rect 1526 694 1532 695
rect 1470 690 1471 694
rect 1475 690 1476 694
rect 1470 689 1476 690
rect 1102 683 1108 684
rect 1102 679 1103 683
rect 1107 679 1108 683
rect 1102 678 1108 679
rect 1426 683 1432 684
rect 1426 679 1427 683
rect 1431 679 1432 683
rect 1426 678 1432 679
rect 1086 677 1092 678
rect 1086 673 1087 677
rect 1091 673 1092 677
rect 1086 672 1092 673
rect 1158 677 1164 678
rect 1158 673 1159 677
rect 1163 673 1164 677
rect 1158 672 1164 673
rect 1222 677 1228 678
rect 1222 673 1223 677
rect 1227 673 1228 677
rect 1222 672 1228 673
rect 1286 677 1292 678
rect 1286 673 1287 677
rect 1291 673 1292 677
rect 1286 672 1292 673
rect 1350 677 1356 678
rect 1350 673 1351 677
rect 1355 673 1356 677
rect 1350 672 1356 673
rect 1414 677 1420 678
rect 1414 673 1415 677
rect 1419 673 1420 677
rect 1414 672 1420 673
rect 1047 670 1051 671
rect 1047 664 1051 666
rect 1087 670 1091 672
rect 1087 665 1091 666
rect 1127 670 1131 671
rect 1127 664 1131 666
rect 1159 670 1163 672
rect 1159 665 1163 666
rect 1215 670 1219 671
rect 1215 664 1219 666
rect 1223 670 1227 672
rect 1223 665 1227 666
rect 1287 670 1291 672
rect 1287 665 1291 666
rect 1295 670 1299 671
rect 1295 664 1299 666
rect 1351 670 1355 672
rect 1351 665 1355 666
rect 1383 670 1387 671
rect 1383 664 1387 666
rect 1415 670 1419 672
rect 1415 665 1419 666
rect 1046 663 1052 664
rect 1046 659 1047 663
rect 1051 659 1052 663
rect 1046 658 1052 659
rect 1126 663 1132 664
rect 1126 659 1127 663
rect 1131 659 1132 663
rect 1126 658 1132 659
rect 1214 663 1220 664
rect 1214 659 1215 663
rect 1219 659 1220 663
rect 1214 658 1220 659
rect 1294 663 1300 664
rect 1294 659 1295 663
rect 1299 659 1300 663
rect 1294 658 1300 659
rect 1382 663 1388 664
rect 1382 659 1383 663
rect 1387 659 1388 663
rect 1382 658 1388 659
rect 1030 655 1036 656
rect 1030 651 1031 655
rect 1035 651 1036 655
rect 1030 650 1036 651
rect 1226 655 1232 656
rect 1226 651 1227 655
rect 1231 651 1232 655
rect 1226 650 1232 651
rect 974 646 980 647
rect 974 642 975 646
rect 979 642 980 646
rect 974 641 980 642
rect 1046 646 1052 647
rect 1046 642 1047 646
rect 1051 642 1052 646
rect 1046 641 1052 642
rect 1126 646 1132 647
rect 1126 642 1127 646
rect 1131 642 1132 646
rect 1126 641 1132 642
rect 1214 646 1220 647
rect 1214 642 1215 646
rect 1219 642 1220 646
rect 1214 641 1220 642
rect 926 639 932 640
rect 926 635 927 639
rect 931 635 932 639
rect 926 634 932 635
rect 976 631 978 641
rect 1048 631 1050 641
rect 1128 631 1130 641
rect 1142 639 1148 640
rect 1142 635 1143 639
rect 1147 635 1148 639
rect 1142 634 1148 635
rect 847 630 851 631
rect 847 625 851 626
rect 895 630 899 631
rect 895 625 899 626
rect 911 630 915 631
rect 911 625 915 626
rect 967 630 971 631
rect 967 625 971 626
rect 975 630 979 631
rect 975 625 979 626
rect 1047 630 1051 631
rect 1047 625 1051 626
rect 1127 630 1131 631
rect 1127 625 1131 626
rect 838 619 844 620
rect 838 615 839 619
rect 843 615 844 619
rect 896 615 898 625
rect 968 615 970 625
rect 1048 615 1050 625
rect 1118 615 1124 616
rect 1128 615 1130 625
rect 518 614 524 615
rect 518 610 519 614
rect 523 610 524 614
rect 518 609 524 610
rect 566 614 572 615
rect 566 610 567 614
rect 571 610 572 614
rect 566 609 572 610
rect 614 614 620 615
rect 614 610 615 614
rect 619 610 620 614
rect 614 609 620 610
rect 662 614 668 615
rect 662 610 663 614
rect 667 610 668 614
rect 662 609 668 610
rect 718 614 724 615
rect 718 610 719 614
rect 723 610 724 614
rect 718 609 724 610
rect 774 614 780 615
rect 774 610 775 614
rect 779 610 780 614
rect 774 609 780 610
rect 830 614 836 615
rect 838 614 844 615
rect 894 614 900 615
rect 830 610 831 614
rect 835 610 836 614
rect 830 609 836 610
rect 894 610 895 614
rect 899 610 900 614
rect 894 609 900 610
rect 966 614 972 615
rect 966 610 967 614
rect 971 610 972 614
rect 966 609 972 610
rect 1046 614 1052 615
rect 1046 610 1047 614
rect 1051 610 1052 614
rect 1118 611 1119 615
rect 1123 611 1124 615
rect 1118 610 1124 611
rect 1126 614 1132 615
rect 1126 610 1127 614
rect 1131 610 1132 614
rect 1046 609 1052 610
rect 480 603 488 604
rect 480 601 483 603
rect 482 599 483 601
rect 487 599 488 603
rect 482 598 488 599
rect 978 603 984 604
rect 978 599 979 603
rect 983 599 984 603
rect 978 598 984 599
rect 278 597 284 598
rect 278 593 279 597
rect 283 593 284 597
rect 278 592 284 593
rect 318 597 324 598
rect 318 593 319 597
rect 323 593 324 597
rect 318 592 324 593
rect 366 597 372 598
rect 366 593 367 597
rect 371 593 372 597
rect 366 592 372 593
rect 422 597 428 598
rect 422 593 423 597
rect 427 593 428 597
rect 422 592 428 593
rect 470 597 476 598
rect 470 593 471 597
rect 475 593 476 597
rect 470 592 476 593
rect 518 597 524 598
rect 518 593 519 597
rect 523 593 524 597
rect 518 592 524 593
rect 566 597 572 598
rect 566 593 567 597
rect 571 593 572 597
rect 566 592 572 593
rect 614 597 620 598
rect 614 593 615 597
rect 619 593 620 597
rect 614 592 620 593
rect 662 597 668 598
rect 662 593 663 597
rect 667 593 668 597
rect 662 592 668 593
rect 718 597 724 598
rect 718 593 719 597
rect 723 593 724 597
rect 718 592 724 593
rect 774 597 780 598
rect 774 593 775 597
rect 779 593 780 597
rect 774 592 780 593
rect 830 597 836 598
rect 830 593 831 597
rect 835 593 836 597
rect 830 592 836 593
rect 894 597 900 598
rect 894 593 895 597
rect 899 593 900 597
rect 894 592 900 593
rect 966 597 972 598
rect 966 593 967 597
rect 971 593 972 597
rect 966 592 972 593
rect 111 590 115 591
rect 111 585 115 586
rect 167 590 171 591
rect 112 582 114 585
rect 167 584 171 586
rect 215 590 219 591
rect 215 584 219 586
rect 247 590 251 592
rect 262 591 268 592
rect 262 587 263 591
rect 267 587 268 591
rect 262 586 268 587
rect 271 590 275 591
rect 247 585 251 586
rect 271 584 275 586
rect 279 590 283 592
rect 279 585 283 586
rect 319 590 323 592
rect 319 585 323 586
rect 335 590 339 591
rect 335 584 339 586
rect 367 590 371 592
rect 367 585 371 586
rect 407 590 411 591
rect 407 584 411 586
rect 423 590 427 592
rect 423 585 427 586
rect 471 590 475 592
rect 471 585 475 586
rect 487 590 491 591
rect 487 584 491 586
rect 519 590 523 592
rect 519 585 523 586
rect 559 590 563 591
rect 559 584 563 586
rect 567 590 571 592
rect 578 591 584 592
rect 578 587 579 591
rect 583 587 584 591
rect 578 586 584 587
rect 615 590 619 592
rect 567 585 571 586
rect 166 583 172 584
rect 110 581 116 582
rect 110 577 111 581
rect 115 577 116 581
rect 166 579 167 583
rect 171 579 172 583
rect 166 578 172 579
rect 214 583 220 584
rect 214 579 215 583
rect 219 579 220 583
rect 214 578 220 579
rect 270 583 276 584
rect 270 579 271 583
rect 275 579 276 583
rect 270 578 276 579
rect 334 583 340 584
rect 334 579 335 583
rect 339 579 340 583
rect 334 578 340 579
rect 406 583 412 584
rect 406 579 407 583
rect 411 579 412 583
rect 406 578 412 579
rect 486 583 492 584
rect 486 579 487 583
rect 491 579 492 583
rect 486 578 492 579
rect 558 583 564 584
rect 558 579 559 583
rect 563 579 564 583
rect 558 578 564 579
rect 110 576 116 577
rect 166 566 172 567
rect 110 564 116 565
rect 110 560 111 564
rect 115 560 116 564
rect 166 562 167 566
rect 171 562 172 566
rect 166 561 172 562
rect 214 566 220 567
rect 214 562 215 566
rect 219 562 220 566
rect 214 561 220 562
rect 270 566 276 567
rect 270 562 271 566
rect 275 562 276 566
rect 270 561 276 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 406 566 412 567
rect 406 562 407 566
rect 411 562 412 566
rect 406 561 412 562
rect 486 566 492 567
rect 486 562 487 566
rect 491 562 492 566
rect 486 561 492 562
rect 558 566 564 567
rect 558 562 559 566
rect 563 562 564 566
rect 558 561 564 562
rect 110 559 116 560
rect 112 547 114 559
rect 168 547 170 561
rect 216 547 218 561
rect 272 547 274 561
rect 336 547 338 561
rect 342 551 348 552
rect 342 547 343 551
rect 347 547 348 551
rect 408 547 410 561
rect 488 547 490 561
rect 510 547 516 548
rect 560 547 562 561
rect 580 560 582 586
rect 615 585 619 586
rect 631 590 635 591
rect 631 584 635 586
rect 663 590 667 592
rect 663 585 667 586
rect 703 590 707 591
rect 703 584 707 586
rect 719 590 723 592
rect 719 585 723 586
rect 767 590 771 591
rect 767 584 771 586
rect 775 590 779 592
rect 775 585 779 586
rect 823 590 827 591
rect 823 584 827 586
rect 831 590 835 592
rect 831 585 835 586
rect 879 590 883 591
rect 879 584 883 586
rect 895 590 899 592
rect 895 585 899 586
rect 935 590 939 591
rect 935 584 939 586
rect 967 590 971 592
rect 967 585 971 586
rect 630 583 636 584
rect 630 579 631 583
rect 635 579 636 583
rect 630 578 636 579
rect 702 583 708 584
rect 702 579 703 583
rect 707 579 708 583
rect 702 578 708 579
rect 766 583 772 584
rect 766 579 767 583
rect 771 579 772 583
rect 766 578 772 579
rect 822 583 828 584
rect 822 579 823 583
rect 827 579 828 583
rect 822 578 828 579
rect 878 583 884 584
rect 878 579 879 583
rect 883 579 884 583
rect 878 578 884 579
rect 934 583 940 584
rect 934 579 935 583
rect 939 579 940 583
rect 934 578 940 579
rect 806 575 812 576
rect 806 571 807 575
rect 811 571 812 575
rect 806 570 812 571
rect 894 575 900 576
rect 894 571 895 575
rect 899 571 900 575
rect 894 570 900 571
rect 630 566 636 567
rect 630 562 631 566
rect 635 562 636 566
rect 630 561 636 562
rect 702 566 708 567
rect 702 562 703 566
rect 707 562 708 566
rect 702 561 708 562
rect 766 566 772 567
rect 766 562 767 566
rect 771 562 772 566
rect 766 561 772 562
rect 578 559 584 560
rect 578 555 579 559
rect 583 555 584 559
rect 578 554 584 555
rect 632 547 634 561
rect 704 547 706 561
rect 768 547 770 561
rect 111 546 115 547
rect 111 541 115 542
rect 135 546 139 547
rect 135 541 139 542
rect 167 546 171 547
rect 167 541 171 542
rect 199 546 203 547
rect 199 541 203 542
rect 215 546 219 547
rect 215 541 219 542
rect 231 546 235 547
rect 231 541 235 542
rect 271 546 275 547
rect 271 541 275 542
rect 279 546 283 547
rect 279 541 283 542
rect 327 546 331 547
rect 327 541 331 542
rect 335 546 339 547
rect 342 546 348 547
rect 375 546 379 547
rect 335 541 339 542
rect 112 533 114 541
rect 110 532 116 533
rect 110 528 111 532
rect 115 528 116 532
rect 136 531 138 541
rect 150 535 156 536
rect 150 531 151 535
rect 155 531 156 535
rect 168 531 170 541
rect 200 531 202 541
rect 232 531 234 541
rect 280 531 282 541
rect 328 531 330 541
rect 110 527 116 528
rect 134 530 140 531
rect 150 530 156 531
rect 166 530 172 531
rect 134 526 135 530
rect 139 526 140 530
rect 134 525 140 526
rect 110 515 116 516
rect 110 511 111 515
rect 115 511 116 515
rect 110 510 116 511
rect 134 513 140 514
rect 112 507 114 510
rect 134 509 135 513
rect 139 509 140 513
rect 134 508 140 509
rect 152 508 154 530
rect 166 526 167 530
rect 171 526 172 530
rect 166 525 172 526
rect 198 530 204 531
rect 198 526 199 530
rect 203 526 204 530
rect 198 525 204 526
rect 230 530 236 531
rect 230 526 231 530
rect 235 526 236 530
rect 230 525 236 526
rect 278 530 284 531
rect 278 526 279 530
rect 283 526 284 530
rect 278 525 284 526
rect 326 530 332 531
rect 326 526 327 530
rect 331 526 332 530
rect 326 525 332 526
rect 344 520 346 546
rect 375 541 379 542
rect 407 546 411 547
rect 407 541 411 542
rect 431 546 435 547
rect 431 541 435 542
rect 487 546 491 547
rect 487 541 491 542
rect 495 546 499 547
rect 510 543 511 547
rect 515 543 516 547
rect 510 542 516 543
rect 559 546 563 547
rect 495 541 499 542
rect 376 531 378 541
rect 432 531 434 541
rect 496 531 498 541
rect 374 530 380 531
rect 374 526 375 530
rect 379 526 380 530
rect 374 525 380 526
rect 430 530 436 531
rect 430 526 431 530
rect 435 526 436 530
rect 430 525 436 526
rect 494 530 500 531
rect 494 526 495 530
rect 499 526 500 530
rect 494 525 500 526
rect 512 520 514 542
rect 559 541 563 542
rect 623 546 627 547
rect 623 541 627 542
rect 631 546 635 547
rect 687 546 691 547
rect 631 541 635 542
rect 638 543 644 544
rect 560 531 562 541
rect 624 531 626 541
rect 638 539 639 543
rect 643 539 644 543
rect 687 541 691 542
rect 703 546 707 547
rect 703 541 707 542
rect 751 546 755 547
rect 751 541 755 542
rect 767 546 771 547
rect 767 541 771 542
rect 638 538 644 539
rect 630 535 636 536
rect 630 531 631 535
rect 635 531 636 535
rect 558 530 564 531
rect 558 526 559 530
rect 563 526 564 530
rect 558 525 564 526
rect 622 530 628 531
rect 630 530 636 531
rect 622 526 623 530
rect 627 526 628 530
rect 622 525 628 526
rect 342 519 348 520
rect 342 515 343 519
rect 347 515 348 519
rect 342 514 348 515
rect 486 519 492 520
rect 486 515 487 519
rect 491 515 492 519
rect 486 514 492 515
rect 510 519 516 520
rect 510 515 511 519
rect 515 515 516 519
rect 510 514 516 515
rect 166 513 172 514
rect 166 509 167 513
rect 171 509 172 513
rect 166 508 172 509
rect 198 513 204 514
rect 198 509 199 513
rect 203 509 204 513
rect 198 508 204 509
rect 230 513 236 514
rect 230 509 231 513
rect 235 509 236 513
rect 230 508 236 509
rect 278 513 284 514
rect 278 509 279 513
rect 283 509 284 513
rect 278 508 284 509
rect 326 513 332 514
rect 326 509 327 513
rect 331 509 332 513
rect 326 508 332 509
rect 374 513 380 514
rect 374 509 375 513
rect 379 509 380 513
rect 374 508 380 509
rect 430 513 436 514
rect 430 509 431 513
rect 435 509 436 513
rect 430 508 436 509
rect 111 506 115 507
rect 111 501 115 502
rect 135 506 139 508
rect 150 507 156 508
rect 150 503 151 507
rect 155 503 156 507
rect 150 502 156 503
rect 167 506 171 508
rect 112 498 114 501
rect 135 500 139 502
rect 167 500 171 502
rect 199 506 203 508
rect 199 500 203 502
rect 231 506 235 508
rect 231 501 235 502
rect 239 506 243 507
rect 239 500 243 502
rect 279 506 283 508
rect 279 501 283 502
rect 287 506 291 507
rect 287 500 291 502
rect 327 506 331 508
rect 327 500 331 502
rect 375 506 379 508
rect 375 500 379 502
rect 423 506 427 507
rect 423 500 427 502
rect 431 506 435 508
rect 431 501 435 502
rect 479 506 483 507
rect 479 500 483 502
rect 134 499 140 500
rect 110 497 116 498
rect 110 493 111 497
rect 115 493 116 497
rect 134 495 135 499
rect 139 495 140 499
rect 134 494 140 495
rect 166 499 172 500
rect 166 495 167 499
rect 171 495 172 499
rect 166 494 172 495
rect 198 499 204 500
rect 198 495 199 499
rect 203 495 204 499
rect 198 494 204 495
rect 238 499 244 500
rect 238 495 239 499
rect 243 495 244 499
rect 238 494 244 495
rect 286 499 292 500
rect 286 495 287 499
rect 291 495 292 499
rect 286 494 292 495
rect 326 499 332 500
rect 326 495 327 499
rect 331 495 332 499
rect 326 494 332 495
rect 374 499 380 500
rect 374 495 375 499
rect 379 495 380 499
rect 374 494 380 495
rect 422 499 428 500
rect 422 495 423 499
rect 427 495 428 499
rect 422 494 428 495
rect 478 499 484 500
rect 478 495 479 499
rect 483 495 484 499
rect 478 494 484 495
rect 110 492 116 493
rect 134 482 140 483
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 134 478 135 482
rect 139 478 140 482
rect 134 477 140 478
rect 166 482 172 483
rect 166 478 167 482
rect 171 478 172 482
rect 166 477 172 478
rect 198 482 204 483
rect 198 478 199 482
rect 203 478 204 482
rect 198 477 204 478
rect 238 482 244 483
rect 238 478 239 482
rect 243 478 244 482
rect 238 477 244 478
rect 286 482 292 483
rect 286 478 287 482
rect 291 478 292 482
rect 286 477 292 478
rect 326 482 332 483
rect 326 478 327 482
rect 331 478 332 482
rect 326 477 332 478
rect 374 482 380 483
rect 374 478 375 482
rect 379 478 380 482
rect 374 477 380 478
rect 422 482 428 483
rect 422 478 423 482
rect 427 478 428 482
rect 422 477 428 478
rect 478 482 484 483
rect 478 478 479 482
rect 483 478 484 482
rect 478 477 484 478
rect 110 475 116 476
rect 112 467 114 475
rect 136 467 138 477
rect 168 467 170 477
rect 200 467 202 477
rect 240 467 242 477
rect 274 475 280 476
rect 274 471 275 475
rect 279 471 280 475
rect 274 470 280 471
rect 111 466 115 467
rect 111 461 115 462
rect 135 466 139 467
rect 135 461 139 462
rect 151 466 155 467
rect 151 461 155 462
rect 167 466 171 467
rect 167 461 171 462
rect 199 466 203 467
rect 199 461 203 462
rect 207 466 211 467
rect 207 461 211 462
rect 239 466 243 467
rect 239 461 243 462
rect 255 466 259 467
rect 255 461 259 462
rect 112 453 114 461
rect 110 452 116 453
rect 110 448 111 452
rect 115 448 116 452
rect 152 451 154 461
rect 190 455 196 456
rect 190 451 191 455
rect 195 451 196 455
rect 208 451 210 461
rect 256 451 258 461
rect 110 447 116 448
rect 150 450 156 451
rect 190 450 196 451
rect 206 450 212 451
rect 150 446 151 450
rect 155 446 156 450
rect 150 445 156 446
rect 110 435 116 436
rect 110 431 111 435
rect 115 431 116 435
rect 110 430 116 431
rect 150 433 156 434
rect 112 427 114 430
rect 150 429 151 433
rect 155 429 156 433
rect 150 428 156 429
rect 111 426 115 427
rect 111 421 115 422
rect 151 426 155 428
rect 151 421 155 422
rect 175 426 179 427
rect 112 418 114 421
rect 175 420 179 422
rect 174 419 180 420
rect 110 417 116 418
rect 110 413 111 417
rect 115 413 116 417
rect 174 415 175 419
rect 179 415 180 419
rect 174 414 180 415
rect 110 412 116 413
rect 192 412 194 450
rect 206 446 207 450
rect 211 446 212 450
rect 206 445 212 446
rect 254 450 260 451
rect 254 446 255 450
rect 259 446 260 450
rect 254 445 260 446
rect 276 440 278 470
rect 288 467 290 477
rect 328 467 330 477
rect 376 467 378 477
rect 424 467 426 477
rect 480 467 482 477
rect 488 476 490 514
rect 494 513 500 514
rect 494 509 495 513
rect 499 509 500 513
rect 494 508 500 509
rect 558 513 564 514
rect 558 509 559 513
rect 563 509 564 513
rect 558 508 564 509
rect 622 513 628 514
rect 622 509 623 513
rect 627 509 628 513
rect 622 508 628 509
rect 495 506 499 508
rect 495 501 499 502
rect 543 506 547 507
rect 543 500 547 502
rect 559 506 563 508
rect 559 501 563 502
rect 615 506 619 507
rect 615 500 619 502
rect 623 506 627 508
rect 623 501 627 502
rect 542 499 548 500
rect 542 495 543 499
rect 547 495 548 499
rect 542 494 548 495
rect 614 499 620 500
rect 614 495 615 499
rect 619 495 620 499
rect 614 494 620 495
rect 632 492 634 530
rect 640 520 642 538
rect 688 531 690 541
rect 752 531 754 541
rect 808 540 810 570
rect 822 566 828 567
rect 822 562 823 566
rect 827 562 828 566
rect 822 561 828 562
rect 878 566 884 567
rect 878 562 879 566
rect 883 562 884 566
rect 878 561 884 562
rect 824 547 826 561
rect 830 547 836 548
rect 880 547 882 561
rect 815 546 819 547
rect 815 541 819 542
rect 823 546 827 547
rect 830 543 831 547
rect 835 543 836 547
rect 830 542 836 543
rect 879 546 883 547
rect 823 541 827 542
rect 806 539 812 540
rect 806 535 807 539
rect 811 535 812 539
rect 806 534 812 535
rect 816 531 818 541
rect 686 530 692 531
rect 686 526 687 530
rect 691 526 692 530
rect 686 525 692 526
rect 750 530 756 531
rect 750 526 751 530
rect 755 526 756 530
rect 750 525 756 526
rect 814 530 820 531
rect 814 526 815 530
rect 819 526 820 530
rect 814 525 820 526
rect 832 520 834 542
rect 879 541 883 542
rect 880 531 882 541
rect 896 536 898 570
rect 934 566 940 567
rect 934 562 935 566
rect 939 562 940 566
rect 934 561 940 562
rect 936 547 938 561
rect 980 560 982 598
rect 1046 597 1052 598
rect 1046 593 1047 597
rect 1051 593 1052 597
rect 1046 592 1052 593
rect 991 590 995 591
rect 991 584 995 586
rect 1047 590 1051 592
rect 1047 584 1051 586
rect 1103 590 1107 591
rect 1103 584 1107 586
rect 990 583 996 584
rect 990 579 991 583
rect 995 579 996 583
rect 990 578 996 579
rect 1046 583 1052 584
rect 1046 579 1047 583
rect 1051 579 1052 583
rect 1046 578 1052 579
rect 1102 583 1108 584
rect 1102 579 1103 583
rect 1107 579 1108 583
rect 1102 578 1108 579
rect 1120 576 1122 610
rect 1126 609 1132 610
rect 1144 604 1146 634
rect 1216 631 1218 641
rect 1207 630 1211 631
rect 1207 625 1211 626
rect 1215 630 1219 631
rect 1215 625 1219 626
rect 1208 615 1210 625
rect 1228 620 1230 650
rect 1294 646 1300 647
rect 1294 642 1295 646
rect 1299 642 1300 646
rect 1294 641 1300 642
rect 1382 646 1388 647
rect 1382 642 1383 646
rect 1387 642 1388 646
rect 1382 641 1388 642
rect 1296 631 1298 641
rect 1384 631 1386 641
rect 1428 640 1430 678
rect 1470 677 1476 678
rect 1470 673 1471 677
rect 1475 673 1476 677
rect 1470 672 1476 673
rect 1471 670 1475 672
rect 1471 664 1475 666
rect 1470 663 1476 664
rect 1470 659 1471 663
rect 1475 659 1476 663
rect 1470 658 1476 659
rect 1488 656 1490 694
rect 1526 690 1527 694
rect 1531 690 1532 694
rect 1526 689 1532 690
rect 1548 684 1550 718
rect 1584 711 1586 725
rect 1624 711 1626 725
rect 1640 712 1642 734
rect 1662 728 1668 729
rect 1662 724 1663 728
rect 1667 724 1668 728
rect 1662 723 1668 724
rect 1638 711 1644 712
rect 1664 711 1666 723
rect 1583 710 1587 711
rect 1583 705 1587 706
rect 1623 710 1627 711
rect 1638 707 1639 711
rect 1643 707 1644 711
rect 1638 706 1644 707
rect 1663 710 1667 711
rect 1623 705 1627 706
rect 1663 705 1667 706
rect 1584 695 1586 705
rect 1624 695 1626 705
rect 1664 697 1666 705
rect 1662 696 1668 697
rect 1582 694 1588 695
rect 1582 690 1583 694
rect 1587 690 1588 694
rect 1582 689 1588 690
rect 1622 694 1628 695
rect 1622 690 1623 694
rect 1627 690 1628 694
rect 1662 692 1663 696
rect 1667 692 1668 696
rect 1662 691 1668 692
rect 1622 689 1628 690
rect 1546 683 1552 684
rect 1546 679 1547 683
rect 1551 679 1552 683
rect 1546 678 1552 679
rect 1638 683 1644 684
rect 1638 679 1639 683
rect 1643 679 1644 683
rect 1638 678 1644 679
rect 1662 679 1668 680
rect 1526 677 1532 678
rect 1526 673 1527 677
rect 1531 673 1532 677
rect 1526 672 1532 673
rect 1582 677 1588 678
rect 1582 673 1583 677
rect 1587 673 1588 677
rect 1582 672 1588 673
rect 1622 677 1628 678
rect 1622 673 1623 677
rect 1627 673 1628 677
rect 1622 672 1628 673
rect 1527 670 1531 672
rect 1527 665 1531 666
rect 1559 670 1563 671
rect 1559 664 1563 666
rect 1583 670 1587 672
rect 1583 665 1587 666
rect 1623 670 1627 672
rect 1623 664 1627 666
rect 1558 663 1564 664
rect 1558 659 1559 663
rect 1563 659 1564 663
rect 1558 658 1564 659
rect 1622 663 1628 664
rect 1622 659 1623 663
rect 1627 659 1628 663
rect 1622 658 1628 659
rect 1486 655 1492 656
rect 1486 651 1487 655
rect 1491 651 1492 655
rect 1486 650 1492 651
rect 1470 646 1476 647
rect 1470 642 1471 646
rect 1475 642 1476 646
rect 1470 641 1476 642
rect 1558 646 1564 647
rect 1558 642 1559 646
rect 1563 642 1564 646
rect 1558 641 1564 642
rect 1622 646 1628 647
rect 1622 642 1623 646
rect 1627 642 1628 646
rect 1622 641 1628 642
rect 1426 639 1432 640
rect 1426 635 1427 639
rect 1431 635 1432 639
rect 1426 634 1432 635
rect 1472 631 1474 641
rect 1560 631 1562 641
rect 1590 639 1596 640
rect 1590 635 1591 639
rect 1595 635 1596 639
rect 1590 634 1596 635
rect 1287 630 1291 631
rect 1287 625 1291 626
rect 1295 630 1299 631
rect 1295 625 1299 626
rect 1359 630 1363 631
rect 1359 625 1363 626
rect 1383 630 1387 631
rect 1383 625 1387 626
rect 1431 630 1435 631
rect 1431 625 1435 626
rect 1471 630 1475 631
rect 1471 625 1475 626
rect 1503 630 1507 631
rect 1503 625 1507 626
rect 1559 630 1563 631
rect 1559 625 1563 626
rect 1575 630 1579 631
rect 1575 625 1579 626
rect 1234 623 1240 624
rect 1226 619 1232 620
rect 1226 615 1227 619
rect 1231 615 1232 619
rect 1234 619 1235 623
rect 1239 619 1240 623
rect 1234 618 1240 619
rect 1206 614 1212 615
rect 1226 614 1232 615
rect 1206 610 1207 614
rect 1211 610 1212 614
rect 1206 609 1212 610
rect 1236 604 1238 618
rect 1288 615 1290 625
rect 1360 615 1362 625
rect 1374 619 1380 620
rect 1374 615 1375 619
rect 1379 615 1380 619
rect 1432 615 1434 625
rect 1504 615 1506 625
rect 1576 615 1578 625
rect 1286 614 1292 615
rect 1286 610 1287 614
rect 1291 610 1292 614
rect 1286 609 1292 610
rect 1358 614 1364 615
rect 1374 614 1380 615
rect 1430 614 1436 615
rect 1358 610 1359 614
rect 1363 610 1364 614
rect 1358 609 1364 610
rect 1142 603 1148 604
rect 1142 599 1143 603
rect 1147 599 1148 603
rect 1142 598 1148 599
rect 1234 603 1240 604
rect 1234 599 1235 603
rect 1239 599 1240 603
rect 1234 598 1240 599
rect 1298 603 1304 604
rect 1298 599 1299 603
rect 1303 599 1304 603
rect 1298 598 1304 599
rect 1126 597 1132 598
rect 1126 593 1127 597
rect 1131 593 1132 597
rect 1126 592 1132 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1286 597 1292 598
rect 1286 593 1287 597
rect 1291 593 1292 597
rect 1286 592 1292 593
rect 1127 590 1131 592
rect 1127 585 1131 586
rect 1159 590 1163 591
rect 1159 584 1163 586
rect 1207 590 1211 592
rect 1207 585 1211 586
rect 1215 590 1219 591
rect 1215 584 1219 586
rect 1271 590 1275 591
rect 1271 584 1275 586
rect 1287 590 1291 592
rect 1287 585 1291 586
rect 1158 583 1164 584
rect 1158 579 1159 583
rect 1163 579 1164 583
rect 1158 578 1164 579
rect 1214 583 1220 584
rect 1214 579 1215 583
rect 1219 579 1220 583
rect 1214 578 1220 579
rect 1270 583 1276 584
rect 1270 579 1271 583
rect 1275 579 1276 583
rect 1270 578 1276 579
rect 1118 575 1124 576
rect 1118 571 1119 575
rect 1123 571 1124 575
rect 1118 570 1124 571
rect 1198 575 1204 576
rect 1198 571 1199 575
rect 1203 571 1204 575
rect 1198 570 1204 571
rect 990 566 996 567
rect 990 562 991 566
rect 995 562 996 566
rect 990 561 996 562
rect 1046 566 1052 567
rect 1046 562 1047 566
rect 1051 562 1052 566
rect 1046 561 1052 562
rect 1102 566 1108 567
rect 1102 562 1103 566
rect 1107 562 1108 566
rect 1102 561 1108 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 978 559 984 560
rect 978 555 979 559
rect 983 555 984 559
rect 978 554 984 555
rect 992 547 994 561
rect 1022 559 1028 560
rect 1022 555 1023 559
rect 1027 555 1028 559
rect 1022 554 1028 555
rect 935 546 939 547
rect 935 541 939 542
rect 943 546 947 547
rect 943 541 947 542
rect 991 546 995 547
rect 991 541 995 542
rect 1007 546 1011 547
rect 1007 541 1011 542
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 944 531 946 541
rect 1008 531 1010 541
rect 878 530 884 531
rect 894 530 900 531
rect 942 530 948 531
rect 878 526 879 530
rect 883 526 884 530
rect 878 525 884 526
rect 942 526 943 530
rect 947 526 948 530
rect 942 525 948 526
rect 1006 530 1012 531
rect 1006 526 1007 530
rect 1011 526 1012 530
rect 1006 525 1012 526
rect 1024 520 1026 554
rect 1048 547 1050 561
rect 1104 547 1106 561
rect 1160 547 1162 561
rect 1047 546 1051 547
rect 1047 541 1051 542
rect 1071 546 1075 547
rect 1071 541 1075 542
rect 1103 546 1107 547
rect 1103 541 1107 542
rect 1127 546 1131 547
rect 1127 541 1131 542
rect 1159 546 1163 547
rect 1159 541 1163 542
rect 1183 546 1187 547
rect 1183 541 1187 542
rect 1072 531 1074 541
rect 1128 531 1130 541
rect 1184 531 1186 541
rect 1200 536 1202 570
rect 1214 566 1220 567
rect 1214 562 1215 566
rect 1219 562 1220 566
rect 1214 561 1220 562
rect 1270 566 1276 567
rect 1270 562 1271 566
rect 1275 562 1276 566
rect 1270 561 1276 562
rect 1216 547 1218 561
rect 1272 547 1274 561
rect 1300 560 1302 598
rect 1358 597 1364 598
rect 1358 593 1359 597
rect 1363 593 1364 597
rect 1358 592 1364 593
rect 1376 592 1378 614
rect 1430 610 1431 614
rect 1435 610 1436 614
rect 1430 609 1436 610
rect 1502 614 1508 615
rect 1502 610 1503 614
rect 1507 610 1508 614
rect 1502 609 1508 610
rect 1574 614 1580 615
rect 1574 610 1575 614
rect 1579 610 1580 614
rect 1574 609 1580 610
rect 1592 604 1594 634
rect 1624 631 1626 641
rect 1640 640 1642 678
rect 1662 675 1663 679
rect 1667 675 1668 679
rect 1662 674 1668 675
rect 1664 671 1666 674
rect 1663 670 1667 671
rect 1663 665 1667 666
rect 1664 662 1666 665
rect 1662 661 1668 662
rect 1662 657 1663 661
rect 1667 657 1668 661
rect 1662 656 1668 657
rect 1662 644 1668 645
rect 1662 640 1663 644
rect 1667 640 1668 644
rect 1638 639 1644 640
rect 1662 639 1668 640
rect 1638 635 1639 639
rect 1643 635 1644 639
rect 1638 634 1644 635
rect 1664 631 1666 639
rect 1623 630 1627 631
rect 1623 625 1627 626
rect 1663 630 1667 631
rect 1663 625 1667 626
rect 1624 615 1626 625
rect 1664 617 1666 625
rect 1662 616 1668 617
rect 1622 614 1628 615
rect 1622 610 1623 614
rect 1627 610 1628 614
rect 1662 612 1663 616
rect 1667 612 1668 616
rect 1662 611 1668 612
rect 1622 609 1628 610
rect 1590 603 1596 604
rect 1590 599 1591 603
rect 1595 599 1596 603
rect 1590 598 1596 599
rect 1638 603 1644 604
rect 1638 599 1639 603
rect 1643 599 1644 603
rect 1638 598 1644 599
rect 1662 599 1668 600
rect 1430 597 1436 598
rect 1430 593 1431 597
rect 1435 593 1436 597
rect 1430 592 1436 593
rect 1502 597 1508 598
rect 1502 593 1503 597
rect 1507 593 1508 597
rect 1502 592 1508 593
rect 1574 597 1580 598
rect 1574 593 1575 597
rect 1579 593 1580 597
rect 1574 592 1580 593
rect 1622 597 1628 598
rect 1622 593 1623 597
rect 1627 593 1628 597
rect 1622 592 1628 593
rect 1327 590 1331 591
rect 1327 584 1331 586
rect 1359 590 1363 592
rect 1374 591 1380 592
rect 1374 587 1375 591
rect 1379 587 1380 591
rect 1374 586 1380 587
rect 1383 590 1387 591
rect 1359 585 1363 586
rect 1383 584 1387 586
rect 1431 590 1435 592
rect 1431 585 1435 586
rect 1447 590 1451 591
rect 1447 584 1451 586
rect 1503 590 1507 592
rect 1503 585 1507 586
rect 1511 590 1515 591
rect 1511 584 1515 586
rect 1575 590 1579 592
rect 1575 584 1579 586
rect 1623 590 1627 592
rect 1623 584 1627 586
rect 1326 583 1332 584
rect 1326 579 1327 583
rect 1331 579 1332 583
rect 1326 578 1332 579
rect 1382 583 1388 584
rect 1382 579 1383 583
rect 1387 579 1388 583
rect 1382 578 1388 579
rect 1446 583 1452 584
rect 1446 579 1447 583
rect 1451 579 1452 583
rect 1446 578 1452 579
rect 1510 583 1516 584
rect 1510 579 1511 583
rect 1515 579 1516 583
rect 1510 578 1516 579
rect 1574 583 1580 584
rect 1574 579 1575 583
rect 1579 579 1580 583
rect 1574 578 1580 579
rect 1622 583 1628 584
rect 1622 579 1623 583
rect 1627 579 1628 583
rect 1622 578 1628 579
rect 1326 566 1332 567
rect 1326 562 1327 566
rect 1331 562 1332 566
rect 1326 561 1332 562
rect 1382 566 1388 567
rect 1382 562 1383 566
rect 1387 562 1388 566
rect 1382 561 1388 562
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1510 566 1516 567
rect 1510 562 1511 566
rect 1515 562 1516 566
rect 1510 561 1516 562
rect 1574 566 1580 567
rect 1574 562 1575 566
rect 1579 562 1580 566
rect 1574 561 1580 562
rect 1622 566 1628 567
rect 1622 562 1623 566
rect 1627 562 1628 566
rect 1622 561 1628 562
rect 1298 559 1304 560
rect 1298 555 1299 559
rect 1303 555 1304 559
rect 1298 554 1304 555
rect 1328 547 1330 561
rect 1384 547 1386 561
rect 1448 547 1450 561
rect 1512 547 1514 561
rect 1526 551 1532 552
rect 1526 547 1527 551
rect 1531 547 1532 551
rect 1576 547 1578 561
rect 1624 547 1626 561
rect 1640 560 1642 598
rect 1662 595 1663 599
rect 1667 595 1668 599
rect 1662 594 1668 595
rect 1664 591 1666 594
rect 1663 590 1667 591
rect 1663 585 1667 586
rect 1664 582 1666 585
rect 1662 581 1668 582
rect 1662 577 1663 581
rect 1667 577 1668 581
rect 1662 576 1668 577
rect 1662 564 1668 565
rect 1662 560 1663 564
rect 1667 560 1668 564
rect 1638 559 1644 560
rect 1662 559 1668 560
rect 1638 555 1639 559
rect 1643 555 1644 559
rect 1638 554 1644 555
rect 1664 547 1666 559
rect 1215 546 1219 547
rect 1215 541 1219 542
rect 1231 546 1235 547
rect 1231 541 1235 542
rect 1271 546 1275 547
rect 1271 541 1275 542
rect 1279 546 1283 547
rect 1279 541 1283 542
rect 1327 546 1331 547
rect 1327 541 1331 542
rect 1335 546 1339 547
rect 1335 541 1339 542
rect 1383 546 1387 547
rect 1383 541 1387 542
rect 1391 546 1395 547
rect 1391 541 1395 542
rect 1447 546 1451 547
rect 1447 541 1451 542
rect 1511 546 1515 547
rect 1526 546 1532 547
rect 1575 546 1579 547
rect 1511 541 1515 542
rect 1198 535 1204 536
rect 1198 531 1199 535
rect 1203 531 1204 535
rect 1232 531 1234 541
rect 1246 535 1252 536
rect 1246 531 1247 535
rect 1251 531 1252 535
rect 1280 531 1282 541
rect 1336 531 1338 541
rect 1392 531 1394 541
rect 1448 531 1450 541
rect 1512 531 1514 541
rect 1070 530 1076 531
rect 1070 526 1071 530
rect 1075 526 1076 530
rect 1070 525 1076 526
rect 1126 530 1132 531
rect 1126 526 1127 530
rect 1131 526 1132 530
rect 1126 525 1132 526
rect 1182 530 1188 531
rect 1198 530 1204 531
rect 1230 530 1236 531
rect 1246 530 1252 531
rect 1278 530 1284 531
rect 1182 526 1183 530
rect 1187 526 1188 530
rect 1182 525 1188 526
rect 1230 526 1231 530
rect 1235 526 1236 530
rect 1230 525 1236 526
rect 638 519 644 520
rect 638 515 639 519
rect 643 515 644 519
rect 638 514 644 515
rect 790 519 796 520
rect 790 515 791 519
rect 795 515 796 519
rect 790 514 796 515
rect 830 519 836 520
rect 830 515 831 519
rect 835 515 836 519
rect 830 514 836 515
rect 1022 519 1028 520
rect 1022 515 1023 519
rect 1027 515 1028 519
rect 1022 514 1028 515
rect 686 513 692 514
rect 686 509 687 513
rect 691 509 692 513
rect 686 508 692 509
rect 750 513 756 514
rect 750 509 751 513
rect 755 509 756 513
rect 750 508 756 509
rect 687 506 691 508
rect 687 501 691 502
rect 695 506 699 507
rect 695 500 699 502
rect 751 506 755 508
rect 751 501 755 502
rect 775 506 779 507
rect 775 500 779 502
rect 694 499 700 500
rect 694 495 695 499
rect 699 495 700 499
rect 694 494 700 495
rect 774 499 780 500
rect 774 495 775 499
rect 779 495 780 499
rect 774 494 780 495
rect 630 491 636 492
rect 630 487 631 491
rect 635 487 636 491
rect 630 486 636 487
rect 542 482 548 483
rect 542 478 543 482
rect 547 478 548 482
rect 542 477 548 478
rect 614 482 620 483
rect 614 478 615 482
rect 619 478 620 482
rect 614 477 620 478
rect 694 482 700 483
rect 694 478 695 482
rect 699 478 700 482
rect 694 477 700 478
rect 774 482 780 483
rect 774 478 775 482
rect 779 478 780 482
rect 774 477 780 478
rect 486 475 492 476
rect 486 471 487 475
rect 491 471 492 475
rect 486 470 492 471
rect 544 467 546 477
rect 616 467 618 477
rect 696 467 698 477
rect 702 475 708 476
rect 702 471 703 475
rect 707 471 708 475
rect 702 470 708 471
rect 287 466 291 467
rect 287 461 291 462
rect 311 466 315 467
rect 311 461 315 462
rect 327 466 331 467
rect 327 461 331 462
rect 367 466 371 467
rect 367 461 371 462
rect 375 466 379 467
rect 375 461 379 462
rect 423 466 427 467
rect 423 461 427 462
rect 439 466 443 467
rect 439 461 443 462
rect 479 466 483 467
rect 479 461 483 462
rect 519 466 523 467
rect 519 461 523 462
rect 543 466 547 467
rect 543 461 547 462
rect 599 466 603 467
rect 599 461 603 462
rect 615 466 619 467
rect 615 461 619 462
rect 679 466 683 467
rect 679 461 683 462
rect 695 466 699 467
rect 695 461 699 462
rect 312 451 314 461
rect 368 451 370 461
rect 440 451 442 461
rect 520 451 522 461
rect 600 451 602 461
rect 680 451 682 461
rect 310 450 316 451
rect 310 446 311 450
rect 315 446 316 450
rect 310 445 316 446
rect 366 450 372 451
rect 366 446 367 450
rect 371 446 372 450
rect 366 445 372 446
rect 438 450 444 451
rect 438 446 439 450
rect 443 446 444 450
rect 438 445 444 446
rect 518 450 524 451
rect 518 446 519 450
rect 523 446 524 450
rect 518 445 524 446
rect 598 450 604 451
rect 598 446 599 450
rect 603 446 604 450
rect 598 445 604 446
rect 678 450 684 451
rect 678 446 679 450
rect 683 446 684 450
rect 678 445 684 446
rect 274 439 280 440
rect 274 435 275 439
rect 279 435 280 439
rect 274 434 280 435
rect 326 439 332 440
rect 326 435 327 439
rect 331 435 332 439
rect 326 434 332 435
rect 695 439 701 440
rect 695 435 696 439
rect 700 438 701 439
rect 704 438 706 470
rect 776 467 778 477
rect 792 476 794 514
rect 814 513 820 514
rect 814 509 815 513
rect 819 509 820 513
rect 814 508 820 509
rect 878 513 884 514
rect 878 509 879 513
rect 883 509 884 513
rect 878 508 884 509
rect 942 513 948 514
rect 942 509 943 513
rect 947 509 948 513
rect 942 508 948 509
rect 1006 513 1012 514
rect 1006 509 1007 513
rect 1011 509 1012 513
rect 1006 508 1012 509
rect 1070 513 1076 514
rect 1070 509 1071 513
rect 1075 509 1076 513
rect 1070 508 1076 509
rect 1126 513 1132 514
rect 1126 509 1127 513
rect 1131 509 1132 513
rect 1126 508 1132 509
rect 1182 513 1188 514
rect 1182 509 1183 513
rect 1187 509 1188 513
rect 1182 508 1188 509
rect 1230 513 1236 514
rect 1230 509 1231 513
rect 1235 509 1236 513
rect 1230 508 1236 509
rect 1248 508 1250 530
rect 1278 526 1279 530
rect 1283 526 1284 530
rect 1278 525 1284 526
rect 1334 530 1340 531
rect 1334 526 1335 530
rect 1339 526 1340 530
rect 1334 525 1340 526
rect 1390 530 1396 531
rect 1390 526 1391 530
rect 1395 526 1396 530
rect 1390 525 1396 526
rect 1446 530 1452 531
rect 1446 526 1447 530
rect 1451 526 1452 530
rect 1446 525 1452 526
rect 1510 530 1516 531
rect 1510 526 1511 530
rect 1515 526 1516 530
rect 1510 525 1516 526
rect 1528 520 1530 546
rect 1575 541 1579 542
rect 1623 546 1627 547
rect 1623 541 1627 542
rect 1663 546 1667 547
rect 1663 541 1667 542
rect 1576 531 1578 541
rect 1624 531 1626 541
rect 1664 533 1666 541
rect 1662 532 1668 533
rect 1574 530 1580 531
rect 1574 526 1575 530
rect 1579 526 1580 530
rect 1574 525 1580 526
rect 1622 530 1628 531
rect 1622 526 1623 530
rect 1627 526 1628 530
rect 1662 528 1663 532
rect 1667 528 1668 532
rect 1662 527 1668 528
rect 1622 525 1628 526
rect 1526 519 1532 520
rect 1526 515 1527 519
rect 1531 515 1532 519
rect 1526 514 1532 515
rect 1606 519 1612 520
rect 1606 515 1607 519
rect 1611 515 1612 519
rect 1606 514 1612 515
rect 1662 515 1668 516
rect 1278 513 1284 514
rect 1278 509 1279 513
rect 1283 509 1284 513
rect 1278 508 1284 509
rect 1334 513 1340 514
rect 1334 509 1335 513
rect 1339 509 1340 513
rect 1334 508 1340 509
rect 1390 513 1396 514
rect 1390 509 1391 513
rect 1395 509 1396 513
rect 1390 508 1396 509
rect 1446 513 1452 514
rect 1446 509 1447 513
rect 1451 509 1452 513
rect 1446 508 1452 509
rect 1510 513 1516 514
rect 1510 509 1511 513
rect 1515 509 1516 513
rect 1510 508 1516 509
rect 1574 513 1580 514
rect 1574 509 1575 513
rect 1579 509 1580 513
rect 1574 508 1580 509
rect 815 506 819 508
rect 815 501 819 502
rect 847 506 851 507
rect 847 500 851 502
rect 879 506 883 508
rect 879 501 883 502
rect 919 506 923 507
rect 919 500 923 502
rect 943 506 947 508
rect 950 507 956 508
rect 950 503 951 507
rect 955 503 956 507
rect 950 502 956 503
rect 983 506 987 507
rect 943 501 947 502
rect 846 499 852 500
rect 846 495 847 499
rect 851 495 852 499
rect 846 494 852 495
rect 918 499 924 500
rect 918 495 919 499
rect 923 495 924 499
rect 918 494 924 495
rect 834 491 840 492
rect 834 487 835 491
rect 839 487 840 491
rect 834 486 840 487
rect 790 475 796 476
rect 836 475 838 486
rect 846 482 852 483
rect 846 478 847 482
rect 851 478 852 482
rect 846 477 852 478
rect 918 482 924 483
rect 918 478 919 482
rect 923 478 924 482
rect 918 477 924 478
rect 790 471 791 475
rect 795 471 796 475
rect 790 470 796 471
rect 832 473 838 475
rect 759 466 763 467
rect 759 461 763 462
rect 775 466 779 467
rect 775 461 779 462
rect 760 451 762 461
rect 832 456 834 473
rect 848 467 850 477
rect 920 467 922 477
rect 952 476 954 502
rect 983 500 987 502
rect 1007 506 1011 508
rect 1007 501 1011 502
rect 1039 506 1043 507
rect 1039 500 1043 502
rect 1071 506 1075 508
rect 1071 501 1075 502
rect 1095 506 1099 507
rect 1095 500 1099 502
rect 1127 506 1131 508
rect 1127 501 1131 502
rect 1143 506 1147 507
rect 1143 500 1147 502
rect 1183 506 1187 508
rect 1183 501 1187 502
rect 1191 506 1195 507
rect 1191 500 1195 502
rect 1231 506 1235 508
rect 1246 507 1252 508
rect 1231 501 1235 502
rect 1239 506 1243 507
rect 1246 503 1247 507
rect 1251 503 1252 507
rect 1246 502 1252 503
rect 1279 506 1283 508
rect 1239 500 1243 502
rect 1279 501 1283 502
rect 1287 506 1291 507
rect 1287 500 1291 502
rect 1335 506 1339 508
rect 1335 500 1339 502
rect 1383 506 1387 507
rect 1383 500 1387 502
rect 1391 506 1395 508
rect 1391 501 1395 502
rect 1431 506 1435 507
rect 1431 500 1435 502
rect 1447 506 1451 508
rect 1447 501 1451 502
rect 1479 506 1483 507
rect 1479 500 1483 502
rect 1511 506 1515 508
rect 1511 501 1515 502
rect 1535 506 1539 507
rect 1535 500 1539 502
rect 1575 506 1579 508
rect 1575 501 1579 502
rect 1591 506 1595 507
rect 1591 500 1595 502
rect 982 499 988 500
rect 982 495 983 499
rect 987 495 988 499
rect 982 494 988 495
rect 1038 499 1044 500
rect 1038 495 1039 499
rect 1043 495 1044 499
rect 1038 494 1044 495
rect 1094 499 1100 500
rect 1094 495 1095 499
rect 1099 495 1100 499
rect 1094 494 1100 495
rect 1142 499 1148 500
rect 1142 495 1143 499
rect 1147 495 1148 499
rect 1142 494 1148 495
rect 1190 499 1196 500
rect 1190 495 1191 499
rect 1195 495 1196 499
rect 1190 494 1196 495
rect 1238 499 1244 500
rect 1238 495 1239 499
rect 1243 495 1244 499
rect 1238 494 1244 495
rect 1286 499 1292 500
rect 1286 495 1287 499
rect 1291 495 1292 499
rect 1286 494 1292 495
rect 1334 499 1340 500
rect 1334 495 1335 499
rect 1339 495 1340 499
rect 1334 494 1340 495
rect 1382 499 1388 500
rect 1382 495 1383 499
rect 1387 495 1388 499
rect 1382 494 1388 495
rect 1430 499 1436 500
rect 1430 495 1431 499
rect 1435 495 1436 499
rect 1430 494 1436 495
rect 1478 499 1484 500
rect 1478 495 1479 499
rect 1483 495 1484 499
rect 1478 494 1484 495
rect 1534 499 1540 500
rect 1534 495 1535 499
rect 1539 495 1540 499
rect 1534 494 1540 495
rect 1590 499 1596 500
rect 1590 495 1591 499
rect 1595 495 1596 499
rect 1590 494 1596 495
rect 1510 491 1516 492
rect 1510 487 1511 491
rect 1515 487 1516 491
rect 1510 486 1516 487
rect 1518 491 1524 492
rect 1518 487 1519 491
rect 1523 487 1524 491
rect 1518 486 1524 487
rect 982 482 988 483
rect 982 478 983 482
rect 987 478 988 482
rect 982 477 988 478
rect 1038 482 1044 483
rect 1038 478 1039 482
rect 1043 478 1044 482
rect 1038 477 1044 478
rect 1094 482 1100 483
rect 1094 478 1095 482
rect 1099 478 1100 482
rect 1094 477 1100 478
rect 1142 482 1148 483
rect 1142 478 1143 482
rect 1147 478 1148 482
rect 1142 477 1148 478
rect 1190 482 1196 483
rect 1190 478 1191 482
rect 1195 478 1196 482
rect 1190 477 1196 478
rect 1238 482 1244 483
rect 1238 478 1239 482
rect 1243 478 1244 482
rect 1238 477 1244 478
rect 1286 482 1292 483
rect 1286 478 1287 482
rect 1291 478 1292 482
rect 1286 477 1292 478
rect 1334 482 1340 483
rect 1334 478 1335 482
rect 1339 478 1340 482
rect 1334 477 1340 478
rect 1382 482 1388 483
rect 1382 478 1383 482
rect 1387 478 1388 482
rect 1382 477 1388 478
rect 1430 482 1436 483
rect 1430 478 1431 482
rect 1435 478 1436 482
rect 1430 477 1436 478
rect 1478 482 1484 483
rect 1478 478 1479 482
rect 1483 478 1484 482
rect 1478 477 1484 478
rect 950 475 956 476
rect 950 471 951 475
rect 955 471 956 475
rect 950 470 956 471
rect 984 467 986 477
rect 998 467 1004 468
rect 1040 467 1042 477
rect 1096 467 1098 477
rect 1144 467 1146 477
rect 1192 467 1194 477
rect 1240 467 1242 477
rect 1288 467 1290 477
rect 1336 467 1338 477
rect 1384 467 1386 477
rect 1390 467 1396 468
rect 1432 467 1434 477
rect 1480 467 1482 477
rect 839 466 843 467
rect 839 461 843 462
rect 847 466 851 467
rect 847 461 851 462
rect 911 466 915 467
rect 911 461 915 462
rect 919 466 923 467
rect 919 461 923 462
rect 983 466 987 467
rect 998 463 999 467
rect 1003 463 1004 467
rect 998 462 1004 463
rect 1039 466 1043 467
rect 983 461 987 462
rect 830 455 836 456
rect 830 451 831 455
rect 835 451 836 455
rect 840 451 842 461
rect 912 451 914 461
rect 984 451 986 461
rect 758 450 764 451
rect 830 450 836 451
rect 838 450 844 451
rect 758 446 759 450
rect 763 446 764 450
rect 758 445 764 446
rect 838 446 839 450
rect 843 446 844 450
rect 838 445 844 446
rect 910 450 916 451
rect 910 446 911 450
rect 915 446 916 450
rect 910 445 916 446
rect 982 450 988 451
rect 982 446 983 450
rect 987 446 988 450
rect 982 445 988 446
rect 1000 440 1002 462
rect 1039 461 1043 462
rect 1055 466 1059 467
rect 1055 461 1059 462
rect 1095 466 1099 467
rect 1095 461 1099 462
rect 1127 466 1131 467
rect 1127 461 1131 462
rect 1143 466 1147 467
rect 1143 461 1147 462
rect 1191 466 1195 467
rect 1191 461 1195 462
rect 1199 466 1203 467
rect 1199 461 1203 462
rect 1239 466 1243 467
rect 1239 461 1243 462
rect 1263 466 1267 467
rect 1263 461 1267 462
rect 1287 466 1291 467
rect 1287 461 1291 462
rect 1319 466 1323 467
rect 1319 461 1323 462
rect 1335 466 1339 467
rect 1335 461 1339 462
rect 1375 466 1379 467
rect 1375 461 1379 462
rect 1383 466 1387 467
rect 1390 463 1391 467
rect 1395 463 1396 467
rect 1390 462 1396 463
rect 1431 466 1435 467
rect 1383 461 1387 462
rect 1056 451 1058 461
rect 1128 451 1130 461
rect 1200 451 1202 461
rect 1214 455 1220 456
rect 1214 451 1215 455
rect 1219 451 1220 455
rect 1264 451 1266 461
rect 1320 451 1322 461
rect 1376 451 1378 461
rect 1054 450 1060 451
rect 1054 446 1055 450
rect 1059 446 1060 450
rect 1054 445 1060 446
rect 1126 450 1132 451
rect 1126 446 1127 450
rect 1131 446 1132 450
rect 1126 445 1132 446
rect 1198 450 1204 451
rect 1214 450 1220 451
rect 1262 450 1268 451
rect 1198 446 1199 450
rect 1203 446 1204 450
rect 1198 445 1204 446
rect 700 436 706 438
rect 822 439 828 440
rect 700 435 701 436
rect 695 434 701 435
rect 822 435 823 439
rect 827 435 828 439
rect 822 434 828 435
rect 950 439 956 440
rect 950 435 951 439
rect 955 435 956 439
rect 950 434 956 435
rect 998 439 1004 440
rect 998 435 999 439
rect 1003 435 1004 439
rect 998 434 1004 435
rect 206 433 212 434
rect 206 429 207 433
rect 211 429 212 433
rect 206 428 212 429
rect 254 433 260 434
rect 254 429 255 433
rect 259 429 260 433
rect 254 428 260 429
rect 310 433 316 434
rect 310 429 311 433
rect 315 429 316 433
rect 310 428 316 429
rect 207 426 211 428
rect 207 421 211 422
rect 223 426 227 427
rect 223 420 227 422
rect 255 426 259 428
rect 255 421 259 422
rect 271 426 275 427
rect 271 420 275 422
rect 311 426 315 428
rect 311 421 315 422
rect 319 426 323 427
rect 319 420 323 422
rect 222 419 228 420
rect 222 415 223 419
rect 227 415 228 419
rect 222 414 228 415
rect 270 419 276 420
rect 270 415 271 419
rect 275 415 276 419
rect 270 414 276 415
rect 318 419 324 420
rect 318 415 319 419
rect 323 415 324 419
rect 318 414 324 415
rect 190 411 196 412
rect 190 407 191 411
rect 195 407 196 411
rect 190 406 196 407
rect 174 402 180 403
rect 110 400 116 401
rect 110 396 111 400
rect 115 396 116 400
rect 174 398 175 402
rect 179 398 180 402
rect 174 397 180 398
rect 222 402 228 403
rect 222 398 223 402
rect 227 398 228 402
rect 222 397 228 398
rect 270 402 276 403
rect 270 398 271 402
rect 275 398 276 402
rect 270 397 276 398
rect 318 402 324 403
rect 318 398 319 402
rect 323 398 324 402
rect 318 397 324 398
rect 110 395 116 396
rect 112 383 114 395
rect 176 383 178 397
rect 224 383 226 397
rect 230 395 236 396
rect 230 391 231 395
rect 235 391 236 395
rect 230 390 236 391
rect 111 382 115 383
rect 111 377 115 378
rect 135 382 139 383
rect 135 377 139 378
rect 167 382 171 383
rect 167 377 171 378
rect 175 382 179 383
rect 175 377 179 378
rect 199 382 203 383
rect 199 377 203 378
rect 223 382 227 383
rect 223 377 227 378
rect 112 369 114 377
rect 110 368 116 369
rect 110 364 111 368
rect 115 364 116 368
rect 136 367 138 377
rect 150 371 156 372
rect 150 367 151 371
rect 155 367 156 371
rect 168 367 170 377
rect 200 367 202 377
rect 110 363 116 364
rect 134 366 140 367
rect 150 366 156 367
rect 166 366 172 367
rect 134 362 135 366
rect 139 362 140 366
rect 134 361 140 362
rect 110 351 116 352
rect 110 347 111 351
rect 115 347 116 351
rect 110 346 116 347
rect 134 349 140 350
rect 112 343 114 346
rect 134 345 135 349
rect 139 345 140 349
rect 134 344 140 345
rect 152 344 154 366
rect 166 362 167 366
rect 171 362 172 366
rect 166 361 172 362
rect 198 366 204 367
rect 198 362 199 366
rect 203 362 204 366
rect 198 361 204 362
rect 232 356 234 390
rect 272 383 274 397
rect 320 383 322 397
rect 328 396 330 434
rect 366 433 372 434
rect 366 429 367 433
rect 371 429 372 433
rect 366 428 372 429
rect 438 433 444 434
rect 438 429 439 433
rect 443 429 444 433
rect 438 428 444 429
rect 518 433 524 434
rect 518 429 519 433
rect 523 429 524 433
rect 518 428 524 429
rect 598 433 604 434
rect 598 429 599 433
rect 603 429 604 433
rect 598 428 604 429
rect 678 433 684 434
rect 678 429 679 433
rect 683 429 684 433
rect 678 428 684 429
rect 758 433 764 434
rect 758 429 759 433
rect 763 429 764 433
rect 758 428 764 429
rect 367 426 371 428
rect 367 420 371 422
rect 415 426 419 427
rect 415 420 419 422
rect 439 426 443 428
rect 439 421 443 422
rect 471 426 475 427
rect 471 420 475 422
rect 519 426 523 428
rect 519 421 523 422
rect 527 426 531 427
rect 527 420 531 422
rect 591 426 595 427
rect 591 420 595 422
rect 599 426 603 428
rect 599 421 603 422
rect 663 426 667 427
rect 663 420 667 422
rect 679 426 683 428
rect 679 421 683 422
rect 735 426 739 427
rect 735 420 739 422
rect 759 426 763 428
rect 759 421 763 422
rect 807 426 811 427
rect 807 420 811 422
rect 366 419 372 420
rect 366 415 367 419
rect 371 415 372 419
rect 366 414 372 415
rect 414 419 420 420
rect 414 415 415 419
rect 419 415 420 419
rect 414 414 420 415
rect 470 419 476 420
rect 470 415 471 419
rect 475 415 476 419
rect 470 414 476 415
rect 526 419 532 420
rect 526 415 527 419
rect 531 415 532 419
rect 526 414 532 415
rect 590 419 596 420
rect 590 415 591 419
rect 595 415 596 419
rect 590 414 596 415
rect 662 419 668 420
rect 662 415 663 419
rect 667 415 668 419
rect 662 414 668 415
rect 734 419 740 420
rect 734 415 735 419
rect 739 415 740 419
rect 734 414 740 415
rect 806 419 812 420
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 426 411 432 412
rect 426 407 427 411
rect 431 407 432 411
rect 426 406 432 407
rect 754 411 760 412
rect 754 407 755 411
rect 759 407 760 411
rect 754 406 760 407
rect 366 402 372 403
rect 366 398 367 402
rect 371 398 372 402
rect 366 397 372 398
rect 414 402 420 403
rect 414 398 415 402
rect 419 398 420 402
rect 414 397 420 398
rect 326 395 332 396
rect 326 391 327 395
rect 331 391 332 395
rect 326 390 332 391
rect 368 383 370 397
rect 416 383 418 397
rect 239 382 243 383
rect 239 377 243 378
rect 271 382 275 383
rect 271 377 275 378
rect 295 382 299 383
rect 295 377 299 378
rect 319 382 323 383
rect 319 377 323 378
rect 351 382 355 383
rect 351 377 355 378
rect 367 382 371 383
rect 367 377 371 378
rect 407 382 411 383
rect 407 377 411 378
rect 415 382 419 383
rect 415 377 419 378
rect 240 367 242 377
rect 296 367 298 377
rect 352 367 354 377
rect 408 367 410 377
rect 428 372 430 406
rect 470 402 476 403
rect 470 398 471 402
rect 475 398 476 402
rect 470 397 476 398
rect 526 402 532 403
rect 526 398 527 402
rect 531 398 532 402
rect 526 397 532 398
rect 590 402 596 403
rect 590 398 591 402
rect 595 398 596 402
rect 590 397 596 398
rect 662 402 668 403
rect 662 398 663 402
rect 667 398 668 402
rect 662 397 668 398
rect 734 402 740 403
rect 734 398 735 402
rect 739 398 740 402
rect 734 397 740 398
rect 472 383 474 397
rect 528 383 530 397
rect 592 383 594 397
rect 664 383 666 397
rect 670 395 676 396
rect 670 391 671 395
rect 675 391 676 395
rect 670 390 676 391
rect 463 382 467 383
rect 463 377 467 378
rect 471 382 475 383
rect 471 377 475 378
rect 519 382 523 383
rect 519 377 523 378
rect 527 382 531 383
rect 527 377 531 378
rect 575 382 579 383
rect 575 377 579 378
rect 591 382 595 383
rect 591 377 595 378
rect 631 382 635 383
rect 631 377 635 378
rect 663 382 667 383
rect 663 377 667 378
rect 426 371 432 372
rect 426 367 427 371
rect 431 367 432 371
rect 464 367 466 377
rect 474 371 480 372
rect 474 367 475 371
rect 479 367 480 371
rect 520 367 522 377
rect 576 367 578 377
rect 632 367 634 377
rect 238 366 244 367
rect 238 362 239 366
rect 243 362 244 366
rect 238 361 244 362
rect 294 366 300 367
rect 294 362 295 366
rect 299 362 300 366
rect 294 361 300 362
rect 350 366 356 367
rect 350 362 351 366
rect 355 362 356 366
rect 350 361 356 362
rect 406 366 412 367
rect 426 366 432 367
rect 462 366 468 367
rect 474 366 480 367
rect 518 366 524 367
rect 406 362 407 366
rect 411 362 412 366
rect 406 361 412 362
rect 462 362 463 366
rect 467 362 468 366
rect 462 361 468 362
rect 230 355 236 356
rect 230 351 231 355
rect 235 351 236 355
rect 230 350 236 351
rect 250 355 256 356
rect 250 351 251 355
rect 255 351 256 355
rect 250 350 256 351
rect 166 349 172 350
rect 166 345 167 349
rect 171 345 172 349
rect 166 344 172 345
rect 198 349 204 350
rect 198 345 199 349
rect 203 345 204 349
rect 198 344 204 345
rect 238 349 244 350
rect 238 345 239 349
rect 243 345 244 349
rect 238 344 244 345
rect 111 342 115 343
rect 111 337 115 338
rect 135 342 139 344
rect 150 343 156 344
rect 150 339 151 343
rect 155 339 156 343
rect 150 338 156 339
rect 167 342 171 344
rect 112 334 114 337
rect 135 336 139 338
rect 167 336 171 338
rect 199 342 203 344
rect 199 337 203 338
rect 207 342 211 343
rect 207 336 211 338
rect 239 342 243 344
rect 239 337 243 338
rect 134 335 140 336
rect 110 333 116 334
rect 110 329 111 333
rect 115 329 116 333
rect 134 331 135 335
rect 139 331 140 335
rect 134 330 140 331
rect 166 335 172 336
rect 166 331 167 335
rect 171 331 172 335
rect 166 330 172 331
rect 206 335 212 336
rect 206 331 207 335
rect 211 331 212 335
rect 206 330 212 331
rect 110 328 116 329
rect 134 318 140 319
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 134 314 135 318
rect 139 314 140 318
rect 134 313 140 314
rect 166 318 172 319
rect 166 314 167 318
rect 171 314 172 318
rect 166 313 172 314
rect 206 318 212 319
rect 206 314 207 318
rect 211 314 212 318
rect 206 313 212 314
rect 110 311 116 312
rect 112 303 114 311
rect 136 303 138 313
rect 150 311 156 312
rect 150 307 151 311
rect 155 307 156 311
rect 150 306 156 307
rect 111 302 115 303
rect 111 297 115 298
rect 135 302 139 303
rect 135 297 139 298
rect 112 289 114 297
rect 110 288 116 289
rect 110 284 111 288
rect 115 284 116 288
rect 136 287 138 297
rect 110 283 116 284
rect 134 286 140 287
rect 134 282 135 286
rect 139 282 140 286
rect 134 281 140 282
rect 152 276 154 306
rect 168 303 170 313
rect 208 303 210 313
rect 252 312 254 350
rect 294 349 300 350
rect 294 345 295 349
rect 299 345 300 349
rect 294 344 300 345
rect 350 349 356 350
rect 350 345 351 349
rect 355 345 356 349
rect 350 344 356 345
rect 406 349 412 350
rect 406 345 407 349
rect 411 345 412 349
rect 406 344 412 345
rect 462 349 468 350
rect 462 345 463 349
rect 467 345 468 349
rect 462 344 468 345
rect 263 342 267 343
rect 263 336 267 338
rect 295 342 299 344
rect 295 337 299 338
rect 327 342 331 343
rect 327 336 331 338
rect 351 342 355 344
rect 351 337 355 338
rect 391 342 395 343
rect 391 336 395 338
rect 407 342 411 344
rect 407 337 411 338
rect 455 342 459 343
rect 455 336 459 338
rect 463 342 467 344
rect 463 337 467 338
rect 262 335 268 336
rect 262 331 263 335
rect 267 331 268 335
rect 262 330 268 331
rect 326 335 332 336
rect 326 331 327 335
rect 331 331 332 335
rect 326 330 332 331
rect 390 335 396 336
rect 390 331 391 335
rect 395 331 396 335
rect 390 330 396 331
rect 454 335 460 336
rect 454 331 455 335
rect 459 331 460 335
rect 454 330 460 331
rect 476 328 478 366
rect 518 362 519 366
rect 523 362 524 366
rect 518 361 524 362
rect 574 366 580 367
rect 574 362 575 366
rect 579 362 580 366
rect 574 361 580 362
rect 630 366 636 367
rect 630 362 631 366
rect 635 362 636 366
rect 630 361 636 362
rect 672 356 674 390
rect 736 383 738 397
rect 687 382 691 383
rect 687 377 691 378
rect 735 382 739 383
rect 735 377 739 378
rect 743 382 747 383
rect 743 377 747 378
rect 688 367 690 377
rect 744 367 746 377
rect 756 372 758 406
rect 806 402 812 403
rect 806 398 807 402
rect 811 398 812 402
rect 806 397 812 398
rect 808 383 810 397
rect 824 396 826 434
rect 838 433 844 434
rect 838 429 839 433
rect 843 429 844 433
rect 838 428 844 429
rect 910 433 916 434
rect 910 429 911 433
rect 915 429 916 433
rect 910 428 916 429
rect 839 426 843 428
rect 839 421 843 422
rect 871 426 875 427
rect 871 420 875 422
rect 911 426 915 428
rect 911 421 915 422
rect 935 426 939 427
rect 935 420 939 422
rect 870 419 876 420
rect 870 415 871 419
rect 875 415 876 419
rect 870 414 876 415
rect 934 419 940 420
rect 934 415 935 419
rect 939 415 940 419
rect 934 414 940 415
rect 882 411 888 412
rect 882 407 883 411
rect 887 407 888 411
rect 882 406 888 407
rect 870 402 876 403
rect 870 398 871 402
rect 875 398 876 402
rect 870 397 876 398
rect 822 395 828 396
rect 822 391 823 395
rect 827 391 828 395
rect 822 390 828 391
rect 814 383 820 384
rect 872 383 874 397
rect 799 382 803 383
rect 799 377 803 378
rect 807 382 811 383
rect 814 379 815 383
rect 819 379 820 383
rect 814 378 820 379
rect 855 382 859 383
rect 807 377 811 378
rect 754 371 760 372
rect 754 367 755 371
rect 759 367 760 371
rect 800 367 802 377
rect 686 366 692 367
rect 686 362 687 366
rect 691 362 692 366
rect 686 361 692 362
rect 742 366 748 367
rect 754 366 760 367
rect 798 366 804 367
rect 742 362 743 366
rect 747 362 748 366
rect 742 361 748 362
rect 798 362 799 366
rect 803 362 804 366
rect 798 361 804 362
rect 816 356 818 378
rect 855 377 859 378
rect 871 382 875 383
rect 871 377 875 378
rect 856 367 858 377
rect 884 372 886 406
rect 934 402 940 403
rect 934 398 935 402
rect 939 398 940 402
rect 934 397 940 398
rect 936 383 938 397
rect 952 396 954 434
rect 982 433 988 434
rect 982 429 983 433
rect 987 429 988 433
rect 982 428 988 429
rect 1054 433 1060 434
rect 1054 429 1055 433
rect 1059 429 1060 433
rect 1054 428 1060 429
rect 1126 433 1132 434
rect 1126 429 1127 433
rect 1131 429 1132 433
rect 1126 428 1132 429
rect 1198 433 1204 434
rect 1198 429 1199 433
rect 1203 429 1204 433
rect 1198 428 1204 429
rect 1216 428 1218 450
rect 1262 446 1263 450
rect 1267 446 1268 450
rect 1262 445 1268 446
rect 1318 450 1324 451
rect 1318 446 1319 450
rect 1323 446 1324 450
rect 1318 445 1324 446
rect 1374 450 1380 451
rect 1374 446 1375 450
rect 1379 446 1380 450
rect 1374 445 1380 446
rect 1392 440 1394 462
rect 1431 461 1435 462
rect 1479 466 1483 467
rect 1479 461 1483 462
rect 1495 466 1499 467
rect 1495 461 1499 462
rect 1432 451 1434 461
rect 1496 451 1498 461
rect 1512 456 1514 486
rect 1520 468 1522 486
rect 1534 482 1540 483
rect 1534 478 1535 482
rect 1539 478 1540 482
rect 1534 477 1540 478
rect 1590 482 1596 483
rect 1590 478 1591 482
rect 1595 478 1596 482
rect 1590 477 1596 478
rect 1518 467 1524 468
rect 1536 467 1538 477
rect 1592 467 1594 477
rect 1608 476 1610 514
rect 1622 513 1628 514
rect 1622 509 1623 513
rect 1627 509 1628 513
rect 1662 511 1663 515
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1622 508 1628 509
rect 1623 506 1627 508
rect 1664 507 1666 510
rect 1623 500 1627 502
rect 1663 506 1667 507
rect 1663 501 1667 502
rect 1622 499 1628 500
rect 1622 495 1623 499
rect 1627 495 1628 499
rect 1664 498 1666 501
rect 1622 494 1628 495
rect 1662 497 1668 498
rect 1662 493 1663 497
rect 1667 493 1668 497
rect 1662 492 1668 493
rect 1638 491 1644 492
rect 1638 487 1639 491
rect 1643 487 1644 491
rect 1638 486 1644 487
rect 1622 482 1628 483
rect 1622 478 1623 482
rect 1627 478 1628 482
rect 1622 477 1628 478
rect 1606 475 1612 476
rect 1606 471 1607 475
rect 1611 471 1612 475
rect 1606 470 1612 471
rect 1624 467 1626 477
rect 1640 468 1642 486
rect 1662 480 1668 481
rect 1662 476 1663 480
rect 1667 476 1668 480
rect 1662 475 1668 476
rect 1638 467 1644 468
rect 1664 467 1666 475
rect 1518 463 1519 467
rect 1523 463 1524 467
rect 1518 462 1524 463
rect 1535 466 1539 467
rect 1535 461 1539 462
rect 1591 466 1595 467
rect 1591 461 1595 462
rect 1623 466 1627 467
rect 1638 463 1639 467
rect 1643 463 1644 467
rect 1638 462 1644 463
rect 1663 466 1667 467
rect 1623 461 1627 462
rect 1663 461 1667 462
rect 1510 455 1516 456
rect 1510 451 1511 455
rect 1515 451 1516 455
rect 1664 453 1666 461
rect 1430 450 1436 451
rect 1430 446 1431 450
rect 1435 446 1436 450
rect 1430 445 1436 446
rect 1494 450 1500 451
rect 1510 450 1516 451
rect 1662 452 1668 453
rect 1494 446 1495 450
rect 1499 446 1500 450
rect 1662 448 1663 452
rect 1667 448 1668 452
rect 1662 447 1668 448
rect 1494 445 1500 446
rect 1350 439 1356 440
rect 1350 435 1351 439
rect 1355 435 1356 439
rect 1350 434 1356 435
rect 1390 439 1396 440
rect 1390 435 1391 439
rect 1395 435 1396 439
rect 1390 434 1396 435
rect 1662 435 1668 436
rect 1262 433 1268 434
rect 1262 429 1263 433
rect 1267 429 1268 433
rect 1262 428 1268 429
rect 1318 433 1324 434
rect 1318 429 1319 433
rect 1323 429 1324 433
rect 1318 428 1324 429
rect 983 426 987 428
rect 983 421 987 422
rect 991 426 995 427
rect 991 420 995 422
rect 1039 426 1043 427
rect 1039 420 1043 422
rect 1055 426 1059 428
rect 1055 421 1059 422
rect 1087 426 1091 427
rect 1087 420 1091 422
rect 1127 426 1131 428
rect 1127 420 1131 422
rect 1167 426 1171 427
rect 1167 420 1171 422
rect 1199 426 1203 428
rect 1214 427 1220 428
rect 1199 421 1203 422
rect 1207 426 1211 427
rect 1214 423 1215 427
rect 1219 423 1220 427
rect 1214 422 1220 423
rect 1247 426 1251 427
rect 1207 420 1211 422
rect 1247 420 1251 422
rect 1263 426 1267 428
rect 1263 421 1267 422
rect 1287 426 1291 427
rect 1287 420 1291 422
rect 1319 426 1323 428
rect 1319 421 1323 422
rect 1335 426 1339 427
rect 1335 420 1339 422
rect 990 419 996 420
rect 990 415 991 419
rect 995 415 996 419
rect 990 414 996 415
rect 1038 419 1044 420
rect 1038 415 1039 419
rect 1043 415 1044 419
rect 1038 414 1044 415
rect 1086 419 1092 420
rect 1086 415 1087 419
rect 1091 415 1092 419
rect 1086 414 1092 415
rect 1126 419 1132 420
rect 1126 415 1127 419
rect 1131 415 1132 419
rect 1126 414 1132 415
rect 1166 419 1172 420
rect 1166 415 1167 419
rect 1171 415 1172 419
rect 1166 414 1172 415
rect 1206 419 1212 420
rect 1206 415 1207 419
rect 1211 415 1212 419
rect 1206 414 1212 415
rect 1246 419 1252 420
rect 1246 415 1247 419
rect 1251 415 1252 419
rect 1246 414 1252 415
rect 1286 419 1292 420
rect 1286 415 1287 419
rect 1291 415 1292 419
rect 1286 414 1292 415
rect 1334 419 1340 420
rect 1334 415 1335 419
rect 1339 415 1340 419
rect 1334 414 1340 415
rect 1002 411 1008 412
rect 1002 407 1003 411
rect 1007 407 1008 411
rect 1002 406 1008 407
rect 990 402 996 403
rect 990 398 991 402
rect 995 398 996 402
rect 990 397 996 398
rect 950 395 956 396
rect 950 391 951 395
rect 955 391 956 395
rect 950 390 956 391
rect 992 383 994 397
rect 1004 388 1006 406
rect 1038 402 1044 403
rect 1038 398 1039 402
rect 1043 398 1044 402
rect 1038 397 1044 398
rect 1086 402 1092 403
rect 1086 398 1087 402
rect 1091 398 1092 402
rect 1086 397 1092 398
rect 1126 402 1132 403
rect 1126 398 1127 402
rect 1131 398 1132 402
rect 1126 397 1132 398
rect 1166 402 1172 403
rect 1166 398 1167 402
rect 1171 398 1172 402
rect 1166 397 1172 398
rect 1206 402 1212 403
rect 1206 398 1207 402
rect 1211 398 1212 402
rect 1206 397 1212 398
rect 1246 402 1252 403
rect 1246 398 1247 402
rect 1251 398 1252 402
rect 1246 397 1252 398
rect 1286 402 1292 403
rect 1286 398 1287 402
rect 1291 398 1292 402
rect 1286 397 1292 398
rect 1334 402 1340 403
rect 1334 398 1335 402
rect 1339 398 1340 402
rect 1334 397 1340 398
rect 1002 387 1008 388
rect 1002 383 1003 387
rect 1007 383 1008 387
rect 1040 383 1042 397
rect 1088 383 1090 397
rect 1110 387 1116 388
rect 1110 383 1111 387
rect 1115 383 1116 387
rect 1128 383 1130 397
rect 1168 383 1170 397
rect 1208 383 1210 397
rect 1248 383 1250 397
rect 1288 383 1290 397
rect 1336 383 1338 397
rect 1352 396 1354 434
rect 1374 433 1380 434
rect 1374 429 1375 433
rect 1379 429 1380 433
rect 1374 428 1380 429
rect 1430 433 1436 434
rect 1430 429 1431 433
rect 1435 429 1436 433
rect 1430 428 1436 429
rect 1494 433 1500 434
rect 1494 429 1495 433
rect 1499 429 1500 433
rect 1662 431 1663 435
rect 1667 431 1668 435
rect 1662 430 1668 431
rect 1494 428 1500 429
rect 1375 426 1379 428
rect 1375 421 1379 422
rect 1383 426 1387 427
rect 1383 420 1387 422
rect 1431 426 1435 428
rect 1431 421 1435 422
rect 1495 426 1499 428
rect 1664 427 1666 430
rect 1495 421 1499 422
rect 1663 426 1667 427
rect 1663 421 1667 422
rect 1382 419 1388 420
rect 1382 415 1383 419
rect 1387 415 1388 419
rect 1664 418 1666 421
rect 1382 414 1388 415
rect 1662 417 1668 418
rect 1662 413 1663 417
rect 1667 413 1668 417
rect 1662 412 1668 413
rect 1382 402 1388 403
rect 1382 398 1383 402
rect 1387 398 1388 402
rect 1382 397 1388 398
rect 1662 400 1668 401
rect 1350 395 1356 396
rect 1350 391 1351 395
rect 1355 391 1356 395
rect 1350 390 1356 391
rect 1384 383 1386 397
rect 1662 396 1663 400
rect 1667 396 1668 400
rect 1662 395 1668 396
rect 1664 383 1666 395
rect 919 382 923 383
rect 919 377 923 378
rect 935 382 939 383
rect 935 377 939 378
rect 983 382 987 383
rect 983 377 987 378
rect 991 382 995 383
rect 1002 382 1008 383
rect 1039 382 1043 383
rect 991 377 995 378
rect 1039 377 1043 378
rect 1087 382 1091 383
rect 1087 377 1091 378
rect 1095 382 1099 383
rect 1110 382 1116 383
rect 1127 382 1131 383
rect 1095 377 1099 378
rect 890 375 896 376
rect 882 371 888 372
rect 882 367 883 371
rect 887 367 888 371
rect 890 371 891 375
rect 895 371 896 375
rect 890 370 896 371
rect 854 366 860 367
rect 882 366 888 367
rect 854 362 855 366
rect 859 362 860 366
rect 854 361 860 362
rect 892 356 894 370
rect 920 367 922 377
rect 984 367 986 377
rect 1040 367 1042 377
rect 1096 367 1098 377
rect 918 366 924 367
rect 918 362 919 366
rect 923 362 924 366
rect 918 361 924 362
rect 982 366 988 367
rect 982 362 983 366
rect 987 362 988 366
rect 982 361 988 362
rect 1038 366 1044 367
rect 1038 362 1039 366
rect 1043 362 1044 366
rect 1038 361 1044 362
rect 1094 366 1100 367
rect 1094 362 1095 366
rect 1099 362 1100 366
rect 1094 361 1100 362
rect 1112 356 1114 382
rect 1127 377 1131 378
rect 1151 382 1155 383
rect 1151 377 1155 378
rect 1167 382 1171 383
rect 1167 377 1171 378
rect 1207 382 1211 383
rect 1207 377 1211 378
rect 1247 382 1251 383
rect 1247 377 1251 378
rect 1255 382 1259 383
rect 1255 377 1259 378
rect 1287 382 1291 383
rect 1287 377 1291 378
rect 1303 382 1307 383
rect 1303 377 1307 378
rect 1335 382 1339 383
rect 1335 377 1339 378
rect 1351 382 1355 383
rect 1351 377 1355 378
rect 1383 382 1387 383
rect 1383 377 1387 378
rect 1399 382 1403 383
rect 1399 377 1403 378
rect 1447 382 1451 383
rect 1447 377 1451 378
rect 1495 382 1499 383
rect 1495 377 1499 378
rect 1543 382 1547 383
rect 1543 377 1547 378
rect 1591 382 1595 383
rect 1591 377 1595 378
rect 1623 382 1627 383
rect 1623 377 1627 378
rect 1663 382 1667 383
rect 1663 377 1667 378
rect 1152 367 1154 377
rect 1158 371 1164 372
rect 1158 367 1159 371
rect 1163 367 1164 371
rect 1208 367 1210 377
rect 1238 375 1244 376
rect 1238 371 1239 375
rect 1243 371 1244 375
rect 1238 370 1244 371
rect 1150 366 1156 367
rect 1158 366 1164 367
rect 1206 366 1212 367
rect 1150 362 1151 366
rect 1155 362 1156 366
rect 1150 361 1156 362
rect 670 355 676 356
rect 670 351 671 355
rect 675 351 676 355
rect 670 350 676 351
rect 698 355 704 356
rect 698 351 699 355
rect 703 351 704 355
rect 698 350 704 351
rect 814 355 820 356
rect 814 351 815 355
rect 819 351 820 355
rect 814 350 820 351
rect 890 355 896 356
rect 890 351 891 355
rect 895 351 896 355
rect 890 350 896 351
rect 1050 355 1056 356
rect 1050 351 1051 355
rect 1055 351 1056 355
rect 1050 350 1056 351
rect 1110 355 1116 356
rect 1110 351 1111 355
rect 1115 351 1116 355
rect 1110 350 1116 351
rect 518 349 524 350
rect 518 345 519 349
rect 523 345 524 349
rect 518 344 524 345
rect 574 349 580 350
rect 574 345 575 349
rect 579 345 580 349
rect 574 344 580 345
rect 630 349 636 350
rect 630 345 631 349
rect 635 345 636 349
rect 630 344 636 345
rect 686 349 692 350
rect 686 345 687 349
rect 691 345 692 349
rect 686 344 692 345
rect 519 342 523 344
rect 519 336 523 338
rect 575 342 579 344
rect 575 336 579 338
rect 631 342 635 344
rect 631 336 635 338
rect 687 342 691 344
rect 687 336 691 338
rect 518 335 524 336
rect 518 331 519 335
rect 523 331 524 335
rect 518 330 524 331
rect 574 335 580 336
rect 574 331 575 335
rect 579 331 580 335
rect 574 330 580 331
rect 630 335 636 336
rect 630 331 631 335
rect 635 331 636 335
rect 630 330 636 331
rect 686 335 692 336
rect 686 331 687 335
rect 691 331 692 335
rect 686 330 692 331
rect 446 327 452 328
rect 446 323 447 327
rect 451 323 452 327
rect 446 322 452 323
rect 474 327 480 328
rect 474 323 475 327
rect 479 323 480 327
rect 474 322 480 323
rect 586 327 592 328
rect 586 323 587 327
rect 591 323 592 327
rect 586 322 592 323
rect 262 318 268 319
rect 262 314 263 318
rect 267 314 268 318
rect 262 313 268 314
rect 326 318 332 319
rect 326 314 327 318
rect 331 314 332 318
rect 326 313 332 314
rect 390 318 396 319
rect 390 314 391 318
rect 395 314 396 318
rect 390 313 396 314
rect 250 311 256 312
rect 250 307 251 311
rect 255 307 256 311
rect 250 306 256 307
rect 264 303 266 313
rect 328 303 330 313
rect 392 303 394 313
rect 167 302 171 303
rect 167 297 171 298
rect 207 302 211 303
rect 207 297 211 298
rect 231 302 235 303
rect 263 302 267 303
rect 231 297 235 298
rect 246 299 252 300
rect 168 287 170 297
rect 232 287 234 297
rect 246 295 247 299
rect 251 295 252 299
rect 263 297 267 298
rect 295 302 299 303
rect 295 297 299 298
rect 327 302 331 303
rect 327 297 331 298
rect 367 302 371 303
rect 367 297 371 298
rect 391 302 395 303
rect 391 297 395 298
rect 439 302 443 303
rect 439 297 443 298
rect 246 294 252 295
rect 238 291 244 292
rect 238 287 239 291
rect 243 287 244 291
rect 166 286 172 287
rect 166 282 167 286
rect 171 282 172 286
rect 166 281 172 282
rect 230 286 236 287
rect 238 286 244 287
rect 230 282 231 286
rect 235 282 236 286
rect 230 281 236 282
rect 150 275 156 276
rect 110 271 116 272
rect 110 267 111 271
rect 115 267 116 271
rect 150 271 151 275
rect 155 271 156 275
rect 150 270 156 271
rect 110 266 116 267
rect 134 269 140 270
rect 112 259 114 266
rect 134 265 135 269
rect 139 265 140 269
rect 134 264 140 265
rect 166 269 172 270
rect 166 265 167 269
rect 171 265 172 269
rect 166 264 172 265
rect 230 269 236 270
rect 230 265 231 269
rect 235 265 236 269
rect 230 264 236 265
rect 136 259 138 264
rect 168 259 170 264
rect 232 259 234 264
rect 111 258 115 259
rect 111 253 115 254
rect 135 258 139 259
rect 112 250 114 253
rect 135 252 139 254
rect 167 258 171 259
rect 167 253 171 254
rect 175 258 179 259
rect 175 252 179 254
rect 231 258 235 259
rect 231 253 235 254
rect 134 251 140 252
rect 110 249 116 250
rect 110 245 111 249
rect 115 245 116 249
rect 134 247 135 251
rect 139 247 140 251
rect 134 246 140 247
rect 174 251 180 252
rect 174 247 175 251
rect 179 247 180 251
rect 174 246 180 247
rect 110 244 116 245
rect 240 244 242 286
rect 248 276 250 294
rect 296 287 298 297
rect 368 287 370 297
rect 440 287 442 297
rect 448 292 450 322
rect 454 318 460 319
rect 454 314 455 318
rect 459 314 460 318
rect 454 313 460 314
rect 518 318 524 319
rect 518 314 519 318
rect 523 314 524 318
rect 518 313 524 314
rect 574 318 580 319
rect 574 314 575 318
rect 579 314 580 318
rect 574 313 580 314
rect 456 303 458 313
rect 520 303 522 313
rect 576 303 578 313
rect 455 302 459 303
rect 455 297 459 298
rect 503 302 507 303
rect 503 297 507 298
rect 519 302 523 303
rect 519 297 523 298
rect 567 302 571 303
rect 567 297 571 298
rect 575 302 579 303
rect 575 297 579 298
rect 446 291 452 292
rect 446 287 447 291
rect 451 287 452 291
rect 504 287 506 297
rect 568 287 570 297
rect 588 292 590 322
rect 630 318 636 319
rect 630 314 631 318
rect 635 314 636 318
rect 630 313 636 314
rect 686 318 692 319
rect 686 314 687 318
rect 691 314 692 318
rect 686 313 692 314
rect 700 313 702 350
rect 742 349 748 350
rect 742 345 743 349
rect 747 345 748 349
rect 742 344 748 345
rect 798 349 804 350
rect 798 345 799 349
rect 803 345 804 349
rect 798 344 804 345
rect 854 349 860 350
rect 854 345 855 349
rect 859 345 860 349
rect 854 344 860 345
rect 918 349 924 350
rect 918 345 919 349
rect 923 345 924 349
rect 918 344 924 345
rect 982 349 988 350
rect 982 345 983 349
rect 987 345 988 349
rect 982 344 988 345
rect 1038 349 1044 350
rect 1038 345 1039 349
rect 1043 345 1044 349
rect 1038 344 1044 345
rect 743 342 747 344
rect 743 337 747 338
rect 751 342 755 343
rect 751 336 755 338
rect 799 342 803 344
rect 799 337 803 338
rect 815 342 819 343
rect 815 336 819 338
rect 855 342 859 344
rect 855 337 859 338
rect 879 342 883 343
rect 879 336 883 338
rect 919 342 923 344
rect 919 337 923 338
rect 951 342 955 343
rect 951 336 955 338
rect 983 342 987 344
rect 983 337 987 338
rect 1031 342 1035 343
rect 1031 336 1035 338
rect 1039 342 1043 344
rect 1039 337 1043 338
rect 750 335 756 336
rect 750 331 751 335
rect 755 331 756 335
rect 750 330 756 331
rect 814 335 820 336
rect 814 331 815 335
rect 819 331 820 335
rect 814 330 820 331
rect 878 335 884 336
rect 878 331 879 335
rect 883 331 884 335
rect 878 330 884 331
rect 950 335 956 336
rect 950 331 951 335
rect 955 331 956 335
rect 950 330 956 331
rect 1030 335 1036 336
rect 1030 331 1031 335
rect 1035 331 1036 335
rect 1030 330 1036 331
rect 750 318 756 319
rect 750 314 751 318
rect 755 314 756 318
rect 750 313 756 314
rect 814 318 820 319
rect 814 314 815 318
rect 819 314 820 318
rect 814 313 820 314
rect 878 318 884 319
rect 878 314 879 318
rect 883 314 884 318
rect 878 313 884 314
rect 950 318 956 319
rect 950 314 951 318
rect 955 314 956 318
rect 950 313 956 314
rect 1030 318 1036 319
rect 1030 314 1031 318
rect 1035 314 1036 318
rect 1030 313 1036 314
rect 632 303 634 313
rect 688 303 690 313
rect 696 312 702 313
rect 694 311 702 312
rect 694 307 695 311
rect 699 307 700 311
rect 694 306 700 307
rect 706 303 712 304
rect 752 303 754 313
rect 816 303 818 313
rect 880 303 882 313
rect 952 303 954 313
rect 1032 303 1034 313
rect 1052 312 1054 350
rect 1094 349 1100 350
rect 1094 345 1095 349
rect 1099 345 1100 349
rect 1094 344 1100 345
rect 1150 349 1156 350
rect 1150 345 1151 349
rect 1155 345 1156 349
rect 1150 344 1156 345
rect 1095 342 1099 344
rect 1095 337 1099 338
rect 1111 342 1115 343
rect 1111 336 1115 338
rect 1151 342 1155 344
rect 1151 337 1155 338
rect 1110 335 1116 336
rect 1110 331 1111 335
rect 1115 331 1116 335
rect 1110 330 1116 331
rect 1160 328 1162 366
rect 1206 362 1207 366
rect 1211 362 1212 366
rect 1206 361 1212 362
rect 1240 356 1242 370
rect 1256 367 1258 377
rect 1304 367 1306 377
rect 1352 367 1354 377
rect 1400 367 1402 377
rect 1438 375 1444 376
rect 1438 371 1439 375
rect 1443 371 1444 375
rect 1438 370 1444 371
rect 1254 366 1260 367
rect 1254 362 1255 366
rect 1259 362 1260 366
rect 1254 361 1260 362
rect 1302 366 1308 367
rect 1302 362 1303 366
rect 1307 362 1308 366
rect 1302 361 1308 362
rect 1350 366 1356 367
rect 1350 362 1351 366
rect 1355 362 1356 366
rect 1350 361 1356 362
rect 1398 366 1404 367
rect 1398 362 1399 366
rect 1403 362 1404 366
rect 1398 361 1404 362
rect 1440 356 1442 370
rect 1448 367 1450 377
rect 1496 367 1498 377
rect 1534 367 1540 368
rect 1544 367 1546 377
rect 1592 367 1594 377
rect 1624 367 1626 377
rect 1664 369 1666 377
rect 1662 368 1668 369
rect 1446 366 1452 367
rect 1446 362 1447 366
rect 1451 362 1452 366
rect 1446 361 1452 362
rect 1494 366 1500 367
rect 1494 362 1495 366
rect 1499 362 1500 366
rect 1534 363 1535 367
rect 1539 363 1540 367
rect 1534 362 1540 363
rect 1542 366 1548 367
rect 1542 362 1543 366
rect 1547 362 1548 366
rect 1494 361 1500 362
rect 1238 355 1244 356
rect 1238 351 1239 355
rect 1243 351 1244 355
rect 1238 350 1244 351
rect 1438 355 1444 356
rect 1438 351 1439 355
rect 1443 351 1444 355
rect 1438 350 1444 351
rect 1206 349 1212 350
rect 1206 345 1207 349
rect 1211 345 1212 349
rect 1206 344 1212 345
rect 1254 349 1260 350
rect 1254 345 1255 349
rect 1259 345 1260 349
rect 1254 344 1260 345
rect 1302 349 1308 350
rect 1302 345 1303 349
rect 1307 345 1308 349
rect 1302 344 1308 345
rect 1350 349 1356 350
rect 1350 345 1351 349
rect 1355 345 1356 349
rect 1350 344 1356 345
rect 1398 349 1404 350
rect 1398 345 1399 349
rect 1403 345 1404 349
rect 1398 344 1404 345
rect 1446 349 1452 350
rect 1446 345 1447 349
rect 1451 345 1452 349
rect 1446 344 1452 345
rect 1494 349 1500 350
rect 1494 345 1495 349
rect 1499 345 1500 349
rect 1494 344 1500 345
rect 1191 342 1195 343
rect 1191 336 1195 338
rect 1207 342 1211 344
rect 1207 337 1211 338
rect 1255 342 1259 344
rect 1255 337 1259 338
rect 1271 342 1275 343
rect 1271 336 1275 338
rect 1303 342 1307 344
rect 1303 337 1307 338
rect 1343 342 1347 343
rect 1343 336 1347 338
rect 1351 342 1355 344
rect 1351 337 1355 338
rect 1399 342 1403 344
rect 1399 337 1403 338
rect 1407 342 1411 343
rect 1407 336 1411 338
rect 1447 342 1451 344
rect 1447 337 1451 338
rect 1463 342 1467 343
rect 1463 336 1467 338
rect 1495 342 1499 344
rect 1495 337 1499 338
rect 1519 342 1523 343
rect 1519 336 1523 338
rect 1536 336 1538 362
rect 1542 361 1548 362
rect 1590 366 1596 367
rect 1590 362 1591 366
rect 1595 362 1596 366
rect 1590 361 1596 362
rect 1622 366 1628 367
rect 1622 362 1623 366
rect 1627 362 1628 366
rect 1662 364 1663 368
rect 1667 364 1668 368
rect 1662 363 1668 364
rect 1622 361 1628 362
rect 1638 355 1644 356
rect 1638 351 1639 355
rect 1643 351 1644 355
rect 1638 350 1644 351
rect 1662 351 1668 352
rect 1542 349 1548 350
rect 1542 345 1543 349
rect 1547 345 1548 349
rect 1542 344 1548 345
rect 1590 349 1596 350
rect 1590 345 1591 349
rect 1595 345 1596 349
rect 1590 344 1596 345
rect 1622 349 1628 350
rect 1622 345 1623 349
rect 1627 345 1628 349
rect 1622 344 1628 345
rect 1543 342 1547 344
rect 1543 337 1547 338
rect 1583 342 1587 343
rect 1583 336 1587 338
rect 1591 342 1595 344
rect 1591 337 1595 338
rect 1623 342 1627 344
rect 1623 336 1627 338
rect 1190 335 1196 336
rect 1190 331 1191 335
rect 1195 331 1196 335
rect 1190 330 1196 331
rect 1270 335 1276 336
rect 1270 331 1271 335
rect 1275 331 1276 335
rect 1270 330 1276 331
rect 1342 335 1348 336
rect 1342 331 1343 335
rect 1347 331 1348 335
rect 1342 330 1348 331
rect 1406 335 1412 336
rect 1406 331 1407 335
rect 1411 331 1412 335
rect 1406 330 1412 331
rect 1462 335 1468 336
rect 1462 331 1463 335
rect 1467 331 1468 335
rect 1462 330 1468 331
rect 1518 335 1524 336
rect 1518 331 1519 335
rect 1523 331 1524 335
rect 1518 330 1524 331
rect 1534 335 1540 336
rect 1534 331 1535 335
rect 1539 331 1540 335
rect 1534 330 1540 331
rect 1582 335 1588 336
rect 1582 331 1583 335
rect 1587 331 1588 335
rect 1582 330 1588 331
rect 1622 335 1628 336
rect 1622 331 1623 335
rect 1627 331 1628 335
rect 1622 330 1628 331
rect 1158 327 1164 328
rect 1158 323 1159 327
rect 1163 323 1164 327
rect 1158 322 1164 323
rect 1110 318 1116 319
rect 1110 314 1111 318
rect 1115 314 1116 318
rect 1110 313 1116 314
rect 1190 318 1196 319
rect 1190 314 1191 318
rect 1195 314 1196 318
rect 1190 313 1196 314
rect 1270 318 1276 319
rect 1270 314 1271 318
rect 1275 314 1276 318
rect 1270 313 1276 314
rect 1342 318 1348 319
rect 1342 314 1343 318
rect 1347 314 1348 318
rect 1342 313 1348 314
rect 1406 318 1412 319
rect 1406 314 1407 318
rect 1411 314 1412 318
rect 1406 313 1412 314
rect 1462 318 1468 319
rect 1462 314 1463 318
rect 1467 314 1468 318
rect 1462 313 1468 314
rect 1518 318 1524 319
rect 1518 314 1519 318
rect 1523 314 1524 318
rect 1518 313 1524 314
rect 1582 318 1588 319
rect 1582 314 1583 318
rect 1587 314 1588 318
rect 1582 313 1588 314
rect 1622 318 1628 319
rect 1622 314 1623 318
rect 1627 314 1628 318
rect 1622 313 1628 314
rect 1050 311 1056 312
rect 1050 307 1051 311
rect 1055 307 1056 311
rect 1050 306 1056 307
rect 1112 303 1114 313
rect 1192 303 1194 313
rect 1272 303 1274 313
rect 1282 311 1288 312
rect 1282 307 1283 311
rect 1287 307 1288 311
rect 1282 306 1288 307
rect 631 302 635 303
rect 631 297 635 298
rect 687 302 691 303
rect 706 299 707 303
rect 711 299 712 303
rect 706 298 712 299
rect 743 302 747 303
rect 687 297 691 298
rect 586 291 592 292
rect 586 287 587 291
rect 591 287 592 291
rect 632 287 634 297
rect 678 291 684 292
rect 678 287 679 291
rect 683 287 684 291
rect 688 287 690 297
rect 294 286 300 287
rect 294 282 295 286
rect 299 282 300 286
rect 294 281 300 282
rect 366 286 372 287
rect 366 282 367 286
rect 371 282 372 286
rect 366 281 372 282
rect 438 286 444 287
rect 446 286 452 287
rect 502 286 508 287
rect 438 282 439 286
rect 443 282 444 286
rect 438 281 444 282
rect 502 282 503 286
rect 507 282 508 286
rect 502 281 508 282
rect 566 286 572 287
rect 586 286 592 287
rect 630 286 636 287
rect 678 286 684 287
rect 686 286 692 287
rect 566 282 567 286
rect 571 282 572 286
rect 566 281 572 282
rect 630 282 631 286
rect 635 282 636 286
rect 630 281 636 282
rect 246 275 252 276
rect 246 271 247 275
rect 251 271 252 275
rect 246 270 252 271
rect 306 275 312 276
rect 306 271 307 275
rect 311 271 312 275
rect 306 270 312 271
rect 534 275 540 276
rect 534 271 535 275
rect 539 271 540 275
rect 534 270 540 271
rect 294 269 300 270
rect 294 265 295 269
rect 299 265 300 269
rect 294 264 300 265
rect 296 259 298 264
rect 247 258 251 259
rect 247 252 251 254
rect 295 258 299 259
rect 295 253 299 254
rect 246 251 252 252
rect 246 247 247 251
rect 251 247 252 251
rect 246 246 252 247
rect 238 243 244 244
rect 238 239 239 243
rect 243 239 244 243
rect 238 238 244 239
rect 134 234 140 235
rect 110 232 116 233
rect 110 228 111 232
rect 115 228 116 232
rect 134 230 135 234
rect 139 230 140 234
rect 134 229 140 230
rect 174 234 180 235
rect 174 230 175 234
rect 179 230 180 234
rect 174 229 180 230
rect 246 234 252 235
rect 246 230 247 234
rect 251 230 252 234
rect 246 229 252 230
rect 110 227 116 228
rect 112 219 114 227
rect 136 219 138 229
rect 150 227 156 228
rect 150 223 151 227
rect 155 223 156 227
rect 150 222 156 223
rect 111 218 115 219
rect 111 213 115 214
rect 135 218 139 219
rect 135 213 139 214
rect 112 205 114 213
rect 110 204 116 205
rect 110 200 111 204
rect 115 200 116 204
rect 136 203 138 213
rect 110 199 116 200
rect 134 202 140 203
rect 134 198 135 202
rect 139 198 140 202
rect 134 197 140 198
rect 152 192 154 222
rect 176 219 178 229
rect 248 219 250 229
rect 308 228 310 270
rect 366 269 372 270
rect 366 265 367 269
rect 371 265 372 269
rect 366 264 372 265
rect 438 269 444 270
rect 438 265 439 269
rect 443 265 444 269
rect 438 264 444 265
rect 502 269 508 270
rect 502 265 503 269
rect 507 265 508 269
rect 502 264 508 265
rect 368 259 370 264
rect 440 259 442 264
rect 504 259 506 264
rect 319 258 323 259
rect 319 252 323 254
rect 367 258 371 259
rect 367 253 371 254
rect 383 258 387 259
rect 383 252 387 254
rect 439 258 443 259
rect 439 253 443 254
rect 447 258 451 259
rect 447 252 451 254
rect 503 258 507 259
rect 503 253 507 254
rect 519 258 523 259
rect 519 252 523 254
rect 318 251 324 252
rect 318 247 319 251
rect 323 247 324 251
rect 318 246 324 247
rect 382 251 388 252
rect 382 247 383 251
rect 387 247 388 251
rect 382 246 388 247
rect 446 251 452 252
rect 446 247 447 251
rect 451 247 452 251
rect 446 246 452 247
rect 518 251 524 252
rect 518 247 519 251
rect 523 247 524 251
rect 518 246 524 247
rect 438 243 444 244
rect 438 239 439 243
rect 443 239 444 243
rect 438 238 444 239
rect 318 234 324 235
rect 318 230 319 234
rect 323 230 324 234
rect 318 229 324 230
rect 382 234 388 235
rect 382 230 383 234
rect 387 230 388 234
rect 382 229 388 230
rect 306 227 312 228
rect 306 223 307 227
rect 311 223 312 227
rect 306 222 312 223
rect 320 219 322 229
rect 384 219 386 229
rect 440 220 442 238
rect 446 234 452 235
rect 446 230 447 234
rect 451 230 452 234
rect 446 229 452 230
rect 518 234 524 235
rect 518 230 519 234
rect 523 230 524 234
rect 518 229 524 230
rect 438 219 444 220
rect 448 219 450 229
rect 520 219 522 229
rect 536 228 538 270
rect 566 269 572 270
rect 566 265 567 269
rect 571 265 572 269
rect 566 264 572 265
rect 630 269 636 270
rect 630 265 631 269
rect 635 265 636 269
rect 630 264 636 265
rect 568 259 570 264
rect 632 259 634 264
rect 567 258 571 259
rect 567 253 571 254
rect 591 258 595 259
rect 591 252 595 254
rect 631 258 635 259
rect 631 253 635 254
rect 663 258 667 259
rect 663 252 667 254
rect 590 251 596 252
rect 590 247 591 251
rect 595 247 596 251
rect 590 246 596 247
rect 662 251 668 252
rect 662 247 663 251
rect 667 247 668 251
rect 662 246 668 247
rect 680 244 682 286
rect 686 282 687 286
rect 691 282 692 286
rect 686 281 692 282
rect 708 276 710 298
rect 743 297 747 298
rect 751 302 755 303
rect 751 297 755 298
rect 807 302 811 303
rect 807 297 811 298
rect 815 302 819 303
rect 815 297 819 298
rect 879 302 883 303
rect 879 297 883 298
rect 951 302 955 303
rect 951 297 955 298
rect 1031 302 1035 303
rect 1031 297 1035 298
rect 1111 302 1115 303
rect 1111 297 1115 298
rect 1191 302 1195 303
rect 1191 297 1195 298
rect 1263 302 1267 303
rect 1263 297 1267 298
rect 1271 302 1275 303
rect 1271 297 1275 298
rect 744 287 746 297
rect 808 287 810 297
rect 880 287 882 297
rect 952 287 954 297
rect 1032 287 1034 297
rect 1112 287 1114 297
rect 1126 291 1132 292
rect 1126 287 1127 291
rect 1131 287 1132 291
rect 1192 287 1194 297
rect 1264 287 1266 297
rect 742 286 748 287
rect 742 282 743 286
rect 747 282 748 286
rect 742 281 748 282
rect 806 286 812 287
rect 806 282 807 286
rect 811 282 812 286
rect 806 281 812 282
rect 878 286 884 287
rect 878 282 879 286
rect 883 282 884 286
rect 878 281 884 282
rect 950 286 956 287
rect 950 282 951 286
rect 955 282 956 286
rect 950 281 956 282
rect 1030 286 1036 287
rect 1030 282 1031 286
rect 1035 282 1036 286
rect 1030 281 1036 282
rect 1110 286 1116 287
rect 1126 286 1132 287
rect 1190 286 1196 287
rect 1110 282 1111 286
rect 1115 282 1116 286
rect 1110 281 1116 282
rect 706 275 712 276
rect 706 271 707 275
rect 711 271 712 275
rect 706 270 712 271
rect 686 269 692 270
rect 686 265 687 269
rect 691 265 692 269
rect 686 264 692 265
rect 742 269 748 270
rect 742 265 743 269
rect 747 265 748 269
rect 742 264 748 265
rect 806 269 812 270
rect 806 265 807 269
rect 811 265 812 269
rect 806 264 812 265
rect 878 269 884 270
rect 878 265 879 269
rect 883 265 884 269
rect 878 264 884 265
rect 950 269 956 270
rect 950 265 951 269
rect 955 265 956 269
rect 950 264 956 265
rect 1030 269 1036 270
rect 1030 265 1031 269
rect 1035 265 1036 269
rect 1030 264 1036 265
rect 1110 269 1116 270
rect 1110 265 1111 269
rect 1115 265 1116 269
rect 1110 264 1116 265
rect 688 259 690 264
rect 744 259 746 264
rect 808 259 810 264
rect 880 259 882 264
rect 914 263 920 264
rect 914 259 915 263
rect 919 259 920 263
rect 952 259 954 264
rect 1032 259 1034 264
rect 1112 259 1114 264
rect 1128 260 1130 286
rect 1190 282 1191 286
rect 1195 282 1196 286
rect 1190 281 1196 282
rect 1262 286 1268 287
rect 1262 282 1263 286
rect 1267 282 1268 286
rect 1262 281 1268 282
rect 1284 276 1286 306
rect 1344 303 1346 313
rect 1408 303 1410 313
rect 1464 303 1466 313
rect 1520 303 1522 313
rect 1584 303 1586 313
rect 1624 303 1626 313
rect 1640 312 1642 350
rect 1662 347 1663 351
rect 1667 347 1668 351
rect 1662 346 1668 347
rect 1664 343 1666 346
rect 1663 342 1667 343
rect 1663 337 1667 338
rect 1664 334 1666 337
rect 1662 333 1668 334
rect 1662 329 1663 333
rect 1667 329 1668 333
rect 1662 328 1668 329
rect 1662 316 1668 317
rect 1662 312 1663 316
rect 1667 312 1668 316
rect 1638 311 1644 312
rect 1662 311 1668 312
rect 1638 307 1639 311
rect 1643 307 1644 311
rect 1638 306 1644 307
rect 1664 303 1666 311
rect 1327 302 1331 303
rect 1327 297 1331 298
rect 1343 302 1347 303
rect 1343 297 1347 298
rect 1391 302 1395 303
rect 1391 297 1395 298
rect 1407 302 1411 303
rect 1407 297 1411 298
rect 1447 302 1451 303
rect 1447 297 1451 298
rect 1463 302 1467 303
rect 1463 297 1467 298
rect 1495 302 1499 303
rect 1495 297 1499 298
rect 1519 302 1523 303
rect 1519 297 1523 298
rect 1543 302 1547 303
rect 1543 297 1547 298
rect 1583 302 1587 303
rect 1583 297 1587 298
rect 1591 302 1595 303
rect 1591 297 1595 298
rect 1623 302 1627 303
rect 1623 297 1627 298
rect 1663 302 1667 303
rect 1663 297 1667 298
rect 1328 287 1330 297
rect 1342 291 1348 292
rect 1342 287 1343 291
rect 1347 287 1348 291
rect 1392 287 1394 297
rect 1448 287 1450 297
rect 1496 287 1498 297
rect 1544 287 1546 297
rect 1592 287 1594 297
rect 1624 287 1626 297
rect 1664 289 1666 297
rect 1662 288 1668 289
rect 1326 286 1332 287
rect 1342 286 1348 287
rect 1390 286 1396 287
rect 1326 282 1327 286
rect 1331 282 1332 286
rect 1326 281 1332 282
rect 1282 275 1288 276
rect 1282 271 1283 275
rect 1287 271 1288 275
rect 1282 270 1288 271
rect 1190 269 1196 270
rect 1190 265 1191 269
rect 1195 265 1196 269
rect 1190 264 1196 265
rect 1262 269 1268 270
rect 1262 265 1263 269
rect 1267 265 1268 269
rect 1262 264 1268 265
rect 1326 269 1332 270
rect 1326 265 1327 269
rect 1331 265 1332 269
rect 1326 264 1332 265
rect 1344 264 1346 286
rect 1390 282 1391 286
rect 1395 282 1396 286
rect 1390 281 1396 282
rect 1446 286 1452 287
rect 1446 282 1447 286
rect 1451 282 1452 286
rect 1446 281 1452 282
rect 1494 286 1500 287
rect 1494 282 1495 286
rect 1499 282 1500 286
rect 1494 281 1500 282
rect 1542 286 1548 287
rect 1542 282 1543 286
rect 1547 282 1548 286
rect 1542 281 1548 282
rect 1590 286 1596 287
rect 1590 282 1591 286
rect 1595 282 1596 286
rect 1590 281 1596 282
rect 1622 286 1628 287
rect 1622 282 1623 286
rect 1627 282 1628 286
rect 1662 284 1663 288
rect 1667 284 1668 288
rect 1662 283 1668 284
rect 1622 281 1628 282
rect 1430 275 1436 276
rect 1430 271 1431 275
rect 1435 271 1436 275
rect 1430 270 1436 271
rect 1662 271 1668 272
rect 1390 269 1396 270
rect 1390 265 1391 269
rect 1395 265 1396 269
rect 1390 264 1396 265
rect 1126 259 1132 260
rect 1192 259 1194 264
rect 1264 259 1266 264
rect 1328 259 1330 264
rect 1342 263 1348 264
rect 1342 259 1343 263
rect 1347 259 1348 263
rect 1392 259 1394 264
rect 687 258 691 259
rect 687 253 691 254
rect 743 258 747 259
rect 743 252 747 254
rect 807 258 811 259
rect 807 253 811 254
rect 823 258 827 259
rect 823 252 827 254
rect 879 258 883 259
rect 879 253 883 254
rect 895 258 899 259
rect 914 258 920 259
rect 951 258 955 259
rect 895 252 899 254
rect 742 251 748 252
rect 742 247 743 251
rect 747 247 748 251
rect 742 246 748 247
rect 822 251 828 252
rect 822 247 823 251
rect 827 247 828 251
rect 822 246 828 247
rect 894 251 900 252
rect 894 247 895 251
rect 899 247 900 251
rect 894 246 900 247
rect 574 243 580 244
rect 574 239 575 243
rect 579 239 580 243
rect 574 238 580 239
rect 678 243 684 244
rect 678 239 679 243
rect 683 239 684 243
rect 678 238 684 239
rect 534 227 540 228
rect 534 223 535 227
rect 539 223 540 227
rect 534 222 540 223
rect 167 218 171 219
rect 167 213 171 214
rect 175 218 179 219
rect 175 213 179 214
rect 207 218 211 219
rect 207 213 211 214
rect 247 218 251 219
rect 247 213 251 214
rect 255 218 259 219
rect 255 213 259 214
rect 303 218 307 219
rect 303 213 307 214
rect 319 218 323 219
rect 319 213 323 214
rect 343 218 347 219
rect 343 213 347 214
rect 375 218 379 219
rect 375 213 379 214
rect 383 218 387 219
rect 383 213 387 214
rect 415 218 419 219
rect 438 215 439 219
rect 443 215 444 219
rect 438 214 444 215
rect 447 218 451 219
rect 415 213 419 214
rect 447 213 451 214
rect 471 218 475 219
rect 519 218 523 219
rect 471 213 475 214
rect 490 215 496 216
rect 168 203 170 213
rect 208 203 210 213
rect 246 207 252 208
rect 246 203 247 207
rect 251 203 252 207
rect 256 203 258 213
rect 304 203 306 213
rect 344 203 346 213
rect 376 203 378 213
rect 390 207 396 208
rect 390 203 391 207
rect 395 203 396 207
rect 416 203 418 213
rect 472 203 474 213
rect 490 211 491 215
rect 495 211 496 215
rect 519 213 523 214
rect 535 218 539 219
rect 535 213 539 214
rect 490 210 496 211
rect 166 202 172 203
rect 166 198 167 202
rect 171 198 172 202
rect 166 197 172 198
rect 206 202 212 203
rect 246 202 252 203
rect 254 202 260 203
rect 206 198 207 202
rect 211 198 212 202
rect 206 197 212 198
rect 150 191 156 192
rect 110 187 116 188
rect 110 183 111 187
rect 115 183 116 187
rect 150 187 151 191
rect 155 187 156 191
rect 150 186 156 187
rect 110 182 116 183
rect 134 185 140 186
rect 112 179 114 182
rect 134 181 135 185
rect 139 181 140 185
rect 134 180 140 181
rect 166 185 172 186
rect 166 181 167 185
rect 171 181 172 185
rect 166 180 172 181
rect 206 185 212 186
rect 206 181 207 185
rect 211 181 212 185
rect 206 180 212 181
rect 111 178 115 179
rect 111 173 115 174
rect 135 178 139 180
rect 112 170 114 173
rect 135 172 139 174
rect 167 178 171 180
rect 167 173 171 174
rect 175 178 179 179
rect 175 172 179 174
rect 207 178 211 180
rect 207 173 211 174
rect 231 178 235 179
rect 231 172 235 174
rect 134 171 140 172
rect 110 169 116 170
rect 110 165 111 169
rect 115 165 116 169
rect 134 167 135 171
rect 139 167 140 171
rect 134 166 140 167
rect 174 171 180 172
rect 174 167 175 171
rect 179 167 180 171
rect 174 166 180 167
rect 230 171 236 172
rect 230 167 231 171
rect 235 167 236 171
rect 230 166 236 167
rect 110 164 116 165
rect 248 164 250 202
rect 254 198 255 202
rect 259 198 260 202
rect 254 197 260 198
rect 302 202 308 203
rect 302 198 303 202
rect 307 198 308 202
rect 302 197 308 198
rect 342 202 348 203
rect 342 198 343 202
rect 347 198 348 202
rect 342 197 348 198
rect 374 202 380 203
rect 390 202 396 203
rect 414 202 420 203
rect 374 198 375 202
rect 379 198 380 202
rect 374 197 380 198
rect 294 191 300 192
rect 294 187 295 191
rect 299 187 300 191
rect 294 186 300 187
rect 254 185 260 186
rect 254 181 255 185
rect 259 181 260 185
rect 254 180 260 181
rect 255 178 259 180
rect 255 173 259 174
rect 287 178 291 179
rect 287 172 291 174
rect 286 171 292 172
rect 286 167 287 171
rect 291 167 292 171
rect 286 166 292 167
rect 246 163 252 164
rect 246 159 247 163
rect 251 159 252 163
rect 246 158 252 159
rect 134 154 140 155
rect 110 152 116 153
rect 110 148 111 152
rect 115 148 116 152
rect 134 150 135 154
rect 139 150 140 154
rect 134 149 140 150
rect 174 154 180 155
rect 174 150 175 154
rect 179 150 180 154
rect 174 149 180 150
rect 230 154 236 155
rect 230 150 231 154
rect 235 150 236 154
rect 230 149 236 150
rect 286 154 292 155
rect 286 150 287 154
rect 291 150 292 154
rect 286 149 292 150
rect 110 147 116 148
rect 112 123 114 147
rect 136 123 138 149
rect 150 147 156 148
rect 150 143 151 147
rect 155 143 156 147
rect 150 142 156 143
rect 111 122 115 123
rect 111 117 115 118
rect 135 122 139 123
rect 135 117 139 118
rect 112 109 114 117
rect 110 108 116 109
rect 110 104 111 108
rect 115 104 116 108
rect 136 107 138 117
rect 110 103 116 104
rect 134 106 140 107
rect 134 102 135 106
rect 139 102 140 106
rect 134 101 140 102
rect 152 96 154 142
rect 176 123 178 149
rect 232 123 234 149
rect 288 123 290 149
rect 296 148 298 186
rect 302 185 308 186
rect 302 181 303 185
rect 307 181 308 185
rect 302 180 308 181
rect 342 185 348 186
rect 342 181 343 185
rect 347 181 348 185
rect 342 180 348 181
rect 374 185 380 186
rect 374 181 375 185
rect 379 181 380 185
rect 374 180 380 181
rect 392 180 394 202
rect 414 198 415 202
rect 419 198 420 202
rect 414 197 420 198
rect 470 202 476 203
rect 470 198 471 202
rect 475 198 476 202
rect 470 197 476 198
rect 492 192 494 210
rect 536 203 538 213
rect 576 208 578 238
rect 590 234 596 235
rect 590 230 591 234
rect 595 230 596 234
rect 590 229 596 230
rect 662 234 668 235
rect 662 230 663 234
rect 667 230 668 234
rect 662 229 668 230
rect 742 234 748 235
rect 742 230 743 234
rect 747 230 748 234
rect 742 229 748 230
rect 822 234 828 235
rect 822 230 823 234
rect 827 230 828 234
rect 822 229 828 230
rect 894 234 900 235
rect 894 230 895 234
rect 899 230 900 234
rect 894 229 900 230
rect 592 219 594 229
rect 664 219 666 229
rect 744 219 746 229
rect 824 219 826 229
rect 896 219 898 229
rect 916 228 918 258
rect 951 253 955 254
rect 967 258 971 259
rect 967 252 971 254
rect 1031 258 1035 259
rect 1031 252 1035 254
rect 1087 258 1091 259
rect 1087 252 1091 254
rect 1111 258 1115 259
rect 1126 255 1127 259
rect 1131 255 1132 259
rect 1126 254 1132 255
rect 1143 258 1147 259
rect 1111 253 1115 254
rect 1143 252 1147 254
rect 1191 258 1195 259
rect 1191 253 1195 254
rect 1199 258 1203 259
rect 1199 252 1203 254
rect 1255 258 1259 259
rect 1255 252 1259 254
rect 1263 258 1267 259
rect 1263 253 1267 254
rect 1311 258 1315 259
rect 1311 252 1315 254
rect 1327 258 1331 259
rect 1342 258 1348 259
rect 1367 258 1371 259
rect 1327 253 1331 254
rect 1367 252 1371 254
rect 1391 258 1395 259
rect 1391 253 1395 254
rect 1415 258 1419 259
rect 1415 252 1419 254
rect 966 251 972 252
rect 966 247 967 251
rect 971 247 972 251
rect 966 246 972 247
rect 1030 251 1036 252
rect 1030 247 1031 251
rect 1035 247 1036 251
rect 1030 246 1036 247
rect 1086 251 1092 252
rect 1086 247 1087 251
rect 1091 247 1092 251
rect 1086 246 1092 247
rect 1142 251 1148 252
rect 1142 247 1143 251
rect 1147 247 1148 251
rect 1142 246 1148 247
rect 1198 251 1204 252
rect 1198 247 1199 251
rect 1203 247 1204 251
rect 1198 246 1204 247
rect 1254 251 1260 252
rect 1254 247 1255 251
rect 1259 247 1260 251
rect 1254 246 1260 247
rect 1310 251 1316 252
rect 1310 247 1311 251
rect 1315 247 1316 251
rect 1310 246 1316 247
rect 1366 251 1372 252
rect 1366 247 1367 251
rect 1371 247 1372 251
rect 1366 246 1372 247
rect 1414 251 1420 252
rect 1414 247 1415 251
rect 1419 247 1420 251
rect 1414 246 1420 247
rect 1322 243 1328 244
rect 1322 239 1323 243
rect 1327 239 1328 243
rect 1322 238 1328 239
rect 966 234 972 235
rect 966 230 967 234
rect 971 230 972 234
rect 966 229 972 230
rect 1030 234 1036 235
rect 1030 230 1031 234
rect 1035 230 1036 234
rect 1030 229 1036 230
rect 1086 234 1092 235
rect 1086 230 1087 234
rect 1091 230 1092 234
rect 1086 229 1092 230
rect 1142 234 1148 235
rect 1142 230 1143 234
rect 1147 230 1148 234
rect 1142 229 1148 230
rect 1198 234 1204 235
rect 1198 230 1199 234
rect 1203 230 1204 234
rect 1198 229 1204 230
rect 1254 234 1260 235
rect 1254 230 1255 234
rect 1259 230 1260 234
rect 1254 229 1260 230
rect 1310 234 1316 235
rect 1310 230 1311 234
rect 1315 230 1316 234
rect 1310 229 1316 230
rect 914 227 920 228
rect 914 223 915 227
rect 919 223 920 227
rect 914 222 920 223
rect 968 219 970 229
rect 1032 219 1034 229
rect 1088 219 1090 229
rect 1144 219 1146 229
rect 1200 219 1202 229
rect 1230 219 1236 220
rect 1256 219 1258 229
rect 1312 219 1314 229
rect 591 218 595 219
rect 591 213 595 214
rect 615 218 619 219
rect 615 213 619 214
rect 663 218 667 219
rect 663 213 667 214
rect 695 218 699 219
rect 695 213 699 214
rect 743 218 747 219
rect 743 213 747 214
rect 775 218 779 219
rect 775 213 779 214
rect 823 218 827 219
rect 823 213 827 214
rect 855 218 859 219
rect 855 213 859 214
rect 895 218 899 219
rect 895 213 899 214
rect 927 218 931 219
rect 927 213 931 214
rect 967 218 971 219
rect 967 213 971 214
rect 999 218 1003 219
rect 999 213 1003 214
rect 1031 218 1035 219
rect 1031 213 1035 214
rect 1071 218 1075 219
rect 1071 213 1075 214
rect 1087 218 1091 219
rect 1087 213 1091 214
rect 1143 218 1147 219
rect 1143 213 1147 214
rect 1199 218 1203 219
rect 1199 213 1203 214
rect 1215 218 1219 219
rect 1230 215 1231 219
rect 1235 215 1236 219
rect 1230 214 1236 215
rect 1255 218 1259 219
rect 1215 213 1219 214
rect 574 207 580 208
rect 574 203 575 207
rect 579 203 580 207
rect 616 203 618 213
rect 696 203 698 213
rect 776 203 778 213
rect 856 203 858 213
rect 870 207 876 208
rect 870 203 871 207
rect 875 203 876 207
rect 928 203 930 213
rect 1000 203 1002 213
rect 1072 203 1074 213
rect 1144 203 1146 213
rect 1216 203 1218 213
rect 534 202 540 203
rect 574 202 580 203
rect 614 202 620 203
rect 534 198 535 202
rect 539 198 540 202
rect 534 197 540 198
rect 614 198 615 202
rect 619 198 620 202
rect 614 197 620 198
rect 694 202 700 203
rect 694 198 695 202
rect 699 198 700 202
rect 694 197 700 198
rect 774 202 780 203
rect 774 198 775 202
rect 779 198 780 202
rect 774 197 780 198
rect 854 202 860 203
rect 870 202 876 203
rect 926 202 932 203
rect 854 198 855 202
rect 859 198 860 202
rect 854 197 860 198
rect 490 191 496 192
rect 490 187 491 191
rect 495 187 496 191
rect 490 186 496 187
rect 786 191 792 192
rect 786 187 787 191
rect 791 187 792 191
rect 786 186 792 187
rect 414 185 420 186
rect 414 181 415 185
rect 419 181 420 185
rect 414 180 420 181
rect 470 185 476 186
rect 470 181 471 185
rect 475 181 476 185
rect 470 180 476 181
rect 534 185 540 186
rect 534 181 535 185
rect 539 181 540 185
rect 534 180 540 181
rect 614 185 620 186
rect 614 181 615 185
rect 619 181 620 185
rect 614 180 620 181
rect 694 185 700 186
rect 694 181 695 185
rect 699 181 700 185
rect 694 180 700 181
rect 774 185 780 186
rect 774 181 775 185
rect 779 181 780 185
rect 774 180 780 181
rect 303 178 307 180
rect 303 173 307 174
rect 343 178 347 180
rect 343 172 347 174
rect 375 178 379 180
rect 390 179 396 180
rect 390 175 391 179
rect 395 175 396 179
rect 390 174 396 175
rect 399 178 403 179
rect 375 173 379 174
rect 399 172 403 174
rect 415 178 419 180
rect 415 173 419 174
rect 455 178 459 179
rect 455 172 459 174
rect 471 178 475 180
rect 471 173 475 174
rect 511 178 515 179
rect 511 172 515 174
rect 535 178 539 180
rect 535 173 539 174
rect 575 178 579 179
rect 575 172 579 174
rect 615 178 619 180
rect 615 173 619 174
rect 639 178 643 179
rect 639 172 643 174
rect 695 178 699 180
rect 695 173 699 174
rect 703 178 707 179
rect 703 172 707 174
rect 767 178 771 179
rect 767 172 771 174
rect 775 178 779 180
rect 775 173 779 174
rect 342 171 348 172
rect 342 167 343 171
rect 347 167 348 171
rect 342 166 348 167
rect 398 171 404 172
rect 398 167 399 171
rect 403 167 404 171
rect 398 166 404 167
rect 454 171 460 172
rect 454 167 455 171
rect 459 167 460 171
rect 454 166 460 167
rect 510 171 516 172
rect 510 167 511 171
rect 515 167 516 171
rect 510 166 516 167
rect 574 171 580 172
rect 574 167 575 171
rect 579 167 580 171
rect 574 166 580 167
rect 638 171 644 172
rect 638 167 639 171
rect 643 167 644 171
rect 638 166 644 167
rect 702 171 708 172
rect 702 167 703 171
rect 707 167 708 171
rect 702 166 708 167
rect 766 171 772 172
rect 766 167 767 171
rect 771 167 772 171
rect 766 166 772 167
rect 438 163 444 164
rect 438 159 439 163
rect 443 159 444 163
rect 438 158 444 159
rect 758 163 764 164
rect 758 159 759 163
rect 763 159 764 163
rect 758 158 764 159
rect 342 154 348 155
rect 342 150 343 154
rect 347 150 348 154
rect 342 149 348 150
rect 398 154 404 155
rect 398 150 399 154
rect 403 150 404 154
rect 398 149 404 150
rect 294 147 300 148
rect 294 143 295 147
rect 299 143 300 147
rect 294 142 300 143
rect 344 123 346 149
rect 400 123 402 149
rect 167 122 171 123
rect 167 117 171 118
rect 175 122 179 123
rect 175 117 179 118
rect 199 122 203 123
rect 199 117 203 118
rect 231 122 235 123
rect 231 117 235 118
rect 263 122 267 123
rect 263 117 267 118
rect 287 122 291 123
rect 287 117 291 118
rect 295 122 299 123
rect 295 117 299 118
rect 327 122 331 123
rect 327 117 331 118
rect 343 122 347 123
rect 343 117 347 118
rect 359 122 363 123
rect 359 117 363 118
rect 391 122 395 123
rect 391 117 395 118
rect 399 122 403 123
rect 399 117 403 118
rect 423 122 427 123
rect 423 117 427 118
rect 168 107 170 117
rect 200 107 202 117
rect 232 107 234 117
rect 264 107 266 117
rect 296 107 298 117
rect 328 107 330 117
rect 360 107 362 117
rect 392 107 394 117
rect 424 107 426 117
rect 440 112 442 158
rect 454 154 460 155
rect 454 150 455 154
rect 459 150 460 154
rect 454 149 460 150
rect 510 154 516 155
rect 510 150 511 154
rect 515 150 516 154
rect 510 149 516 150
rect 574 154 580 155
rect 574 150 575 154
rect 579 150 580 154
rect 574 149 580 150
rect 638 154 644 155
rect 638 150 639 154
rect 643 150 644 154
rect 638 149 644 150
rect 702 154 708 155
rect 702 150 703 154
rect 707 150 708 154
rect 702 149 708 150
rect 456 123 458 149
rect 478 131 484 132
rect 478 127 479 131
rect 483 127 484 131
rect 478 126 484 127
rect 455 122 459 123
rect 455 117 459 118
rect 463 122 467 123
rect 463 117 467 118
rect 438 111 444 112
rect 438 107 439 111
rect 443 107 444 111
rect 464 107 466 117
rect 480 112 482 126
rect 512 123 514 149
rect 576 123 578 149
rect 640 123 642 149
rect 704 123 706 149
rect 760 132 762 158
rect 766 154 772 155
rect 766 150 767 154
rect 771 150 772 154
rect 766 149 772 150
rect 758 131 764 132
rect 758 127 759 131
rect 763 127 764 131
rect 758 126 764 127
rect 768 123 770 149
rect 788 140 790 186
rect 854 185 860 186
rect 854 181 855 185
rect 859 181 860 185
rect 854 180 860 181
rect 872 180 874 202
rect 926 198 927 202
rect 931 198 932 202
rect 926 197 932 198
rect 998 202 1004 203
rect 998 198 999 202
rect 1003 198 1004 202
rect 998 197 1004 198
rect 1070 202 1076 203
rect 1070 198 1071 202
rect 1075 198 1076 202
rect 1070 197 1076 198
rect 1142 202 1148 203
rect 1142 198 1143 202
rect 1147 198 1148 202
rect 1142 197 1148 198
rect 1214 202 1220 203
rect 1214 198 1215 202
rect 1219 198 1220 202
rect 1214 197 1220 198
rect 1232 192 1234 214
rect 1255 213 1259 214
rect 1287 218 1291 219
rect 1287 213 1291 214
rect 1311 218 1315 219
rect 1311 213 1315 214
rect 1288 203 1290 213
rect 1324 208 1326 238
rect 1366 234 1372 235
rect 1366 230 1367 234
rect 1371 230 1372 234
rect 1366 229 1372 230
rect 1414 234 1420 235
rect 1414 230 1415 234
rect 1419 230 1420 234
rect 1414 229 1420 230
rect 1368 219 1370 229
rect 1416 219 1418 229
rect 1432 228 1434 270
rect 1446 269 1452 270
rect 1446 265 1447 269
rect 1451 265 1452 269
rect 1446 264 1452 265
rect 1494 269 1500 270
rect 1494 265 1495 269
rect 1499 265 1500 269
rect 1494 264 1500 265
rect 1542 269 1548 270
rect 1542 265 1543 269
rect 1547 265 1548 269
rect 1542 264 1548 265
rect 1590 269 1596 270
rect 1590 265 1591 269
rect 1595 265 1596 269
rect 1590 264 1596 265
rect 1622 269 1628 270
rect 1622 265 1623 269
rect 1627 265 1628 269
rect 1662 267 1663 271
rect 1667 267 1668 271
rect 1662 266 1668 267
rect 1622 264 1628 265
rect 1448 259 1450 264
rect 1496 259 1498 264
rect 1544 259 1546 264
rect 1592 259 1594 264
rect 1624 259 1626 264
rect 1664 259 1666 266
rect 1447 258 1451 259
rect 1447 253 1451 254
rect 1463 258 1467 259
rect 1463 252 1467 254
rect 1495 258 1499 259
rect 1495 253 1499 254
rect 1519 258 1523 259
rect 1519 252 1523 254
rect 1543 258 1547 259
rect 1543 253 1547 254
rect 1575 258 1579 259
rect 1575 252 1579 254
rect 1591 258 1595 259
rect 1591 253 1595 254
rect 1623 258 1627 259
rect 1623 252 1627 254
rect 1663 258 1667 259
rect 1663 253 1667 254
rect 1462 251 1468 252
rect 1462 247 1463 251
rect 1467 247 1468 251
rect 1462 246 1468 247
rect 1518 251 1524 252
rect 1518 247 1519 251
rect 1523 247 1524 251
rect 1518 246 1524 247
rect 1574 251 1580 252
rect 1574 247 1575 251
rect 1579 247 1580 251
rect 1574 246 1580 247
rect 1622 251 1628 252
rect 1622 247 1623 251
rect 1627 247 1628 251
rect 1664 250 1666 253
rect 1622 246 1628 247
rect 1662 249 1668 250
rect 1662 245 1663 249
rect 1667 245 1668 249
rect 1662 244 1668 245
rect 1634 243 1640 244
rect 1634 239 1635 243
rect 1639 239 1640 243
rect 1634 238 1640 239
rect 1462 234 1468 235
rect 1462 230 1463 234
rect 1467 230 1468 234
rect 1462 229 1468 230
rect 1518 234 1524 235
rect 1518 230 1519 234
rect 1523 230 1524 234
rect 1518 229 1524 230
rect 1574 234 1580 235
rect 1574 230 1575 234
rect 1579 230 1580 234
rect 1574 229 1580 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1430 227 1436 228
rect 1430 223 1431 227
rect 1435 223 1436 227
rect 1430 222 1436 223
rect 1464 219 1466 229
rect 1482 227 1488 228
rect 1482 223 1483 227
rect 1487 223 1488 227
rect 1482 222 1488 223
rect 1351 218 1355 219
rect 1351 213 1355 214
rect 1367 218 1371 219
rect 1367 213 1371 214
rect 1415 218 1419 219
rect 1415 213 1419 214
rect 1463 218 1467 219
rect 1463 213 1467 214
rect 1471 218 1475 219
rect 1471 213 1475 214
rect 1330 211 1336 212
rect 1322 207 1328 208
rect 1322 203 1323 207
rect 1327 203 1328 207
rect 1330 207 1331 211
rect 1335 207 1336 211
rect 1330 206 1336 207
rect 1286 202 1292 203
rect 1322 202 1328 203
rect 1286 198 1287 202
rect 1291 198 1292 202
rect 1286 197 1292 198
rect 1332 192 1334 206
rect 1352 203 1354 213
rect 1416 203 1418 213
rect 1454 211 1460 212
rect 1434 207 1440 208
rect 1434 203 1435 207
rect 1439 203 1440 207
rect 1454 207 1455 211
rect 1459 207 1460 211
rect 1454 206 1460 207
rect 1350 202 1356 203
rect 1350 198 1351 202
rect 1355 198 1356 202
rect 1350 197 1356 198
rect 1414 202 1420 203
rect 1434 202 1440 203
rect 1414 198 1415 202
rect 1419 198 1420 202
rect 1414 197 1420 198
rect 1230 191 1236 192
rect 1230 187 1231 191
rect 1235 187 1236 191
rect 1230 186 1236 187
rect 1330 191 1336 192
rect 1330 187 1331 191
rect 1335 187 1336 191
rect 1330 186 1336 187
rect 1366 191 1372 192
rect 1366 187 1367 191
rect 1371 187 1372 191
rect 1366 186 1372 187
rect 926 185 932 186
rect 926 181 927 185
rect 931 181 932 185
rect 926 180 932 181
rect 998 185 1004 186
rect 998 181 999 185
rect 1003 181 1004 185
rect 998 180 1004 181
rect 1070 185 1076 186
rect 1070 181 1071 185
rect 1075 181 1076 185
rect 1070 180 1076 181
rect 1142 185 1148 186
rect 1142 181 1143 185
rect 1147 181 1148 185
rect 1142 180 1148 181
rect 1214 185 1220 186
rect 1214 181 1215 185
rect 1219 181 1220 185
rect 1214 180 1220 181
rect 1286 185 1292 186
rect 1286 181 1287 185
rect 1291 181 1292 185
rect 1286 180 1292 181
rect 1350 185 1356 186
rect 1350 181 1351 185
rect 1355 181 1356 185
rect 1350 180 1356 181
rect 831 178 835 179
rect 831 172 835 174
rect 855 178 859 180
rect 870 179 876 180
rect 870 175 871 179
rect 875 175 876 179
rect 870 174 876 175
rect 895 178 899 179
rect 855 173 859 174
rect 895 172 899 174
rect 927 178 931 180
rect 927 173 931 174
rect 951 178 955 179
rect 951 172 955 174
rect 999 178 1003 180
rect 999 173 1003 174
rect 1015 178 1019 179
rect 1015 172 1019 174
rect 1071 178 1075 180
rect 1071 173 1075 174
rect 1079 178 1083 179
rect 1079 172 1083 174
rect 1143 178 1147 180
rect 1143 172 1147 174
rect 1207 178 1211 179
rect 1207 172 1211 174
rect 1215 178 1219 180
rect 1215 173 1219 174
rect 1279 178 1283 179
rect 1279 172 1283 174
rect 1287 178 1291 180
rect 1287 173 1291 174
rect 1351 178 1355 180
rect 1351 172 1355 174
rect 830 171 836 172
rect 830 167 831 171
rect 835 167 836 171
rect 830 166 836 167
rect 894 171 900 172
rect 894 167 895 171
rect 899 167 900 171
rect 894 166 900 167
rect 950 171 956 172
rect 950 167 951 171
rect 955 167 956 171
rect 950 166 956 167
rect 1014 171 1020 172
rect 1014 167 1015 171
rect 1019 167 1020 171
rect 1014 166 1020 167
rect 1078 171 1084 172
rect 1078 167 1079 171
rect 1083 167 1084 171
rect 1078 166 1084 167
rect 1142 171 1148 172
rect 1142 167 1143 171
rect 1147 167 1148 171
rect 1142 166 1148 167
rect 1206 171 1212 172
rect 1206 167 1207 171
rect 1211 167 1212 171
rect 1206 166 1212 167
rect 1278 171 1284 172
rect 1278 167 1279 171
rect 1283 167 1284 171
rect 1278 166 1284 167
rect 1350 171 1356 172
rect 1350 167 1351 171
rect 1355 167 1356 171
rect 1350 166 1356 167
rect 1198 163 1204 164
rect 1198 159 1199 163
rect 1203 159 1204 163
rect 1198 158 1204 159
rect 830 154 836 155
rect 830 150 831 154
rect 835 150 836 154
rect 830 149 836 150
rect 894 154 900 155
rect 894 150 895 154
rect 899 150 900 154
rect 894 149 900 150
rect 950 154 956 155
rect 950 150 951 154
rect 955 150 956 154
rect 950 149 956 150
rect 1014 154 1020 155
rect 1014 150 1015 154
rect 1019 150 1020 154
rect 1014 149 1020 150
rect 1078 154 1084 155
rect 1078 150 1079 154
rect 1083 150 1084 154
rect 1078 149 1084 150
rect 1142 154 1148 155
rect 1142 150 1143 154
rect 1147 150 1148 154
rect 1142 149 1148 150
rect 786 139 792 140
rect 786 135 787 139
rect 791 135 792 139
rect 786 134 792 135
rect 832 123 834 149
rect 896 123 898 149
rect 952 123 954 149
rect 1016 123 1018 149
rect 1080 123 1082 149
rect 1144 123 1146 149
rect 1158 139 1164 140
rect 1158 135 1159 139
rect 1163 135 1164 139
rect 1158 134 1164 135
rect 503 122 507 123
rect 503 117 507 118
rect 511 122 515 123
rect 511 117 515 118
rect 543 122 547 123
rect 543 117 547 118
rect 575 122 579 123
rect 575 117 579 118
rect 607 122 611 123
rect 607 117 611 118
rect 639 122 643 123
rect 639 117 643 118
rect 671 122 675 123
rect 671 117 675 118
rect 703 122 707 123
rect 703 117 707 118
rect 735 122 739 123
rect 735 117 739 118
rect 767 122 771 123
rect 767 117 771 118
rect 799 122 803 123
rect 799 117 803 118
rect 831 122 835 123
rect 831 117 835 118
rect 863 122 867 123
rect 863 117 867 118
rect 895 122 899 123
rect 895 117 899 118
rect 935 122 939 123
rect 935 117 939 118
rect 951 122 955 123
rect 951 117 955 118
rect 975 122 979 123
rect 975 117 979 118
rect 1015 122 1019 123
rect 1015 117 1019 118
rect 1063 122 1067 123
rect 1063 117 1067 118
rect 1079 122 1083 123
rect 1079 117 1083 118
rect 1103 122 1107 123
rect 1103 117 1107 118
rect 1143 122 1147 123
rect 1143 117 1147 118
rect 478 111 484 112
rect 478 107 479 111
rect 483 107 484 111
rect 504 107 506 117
rect 544 107 546 117
rect 576 107 578 117
rect 608 107 610 117
rect 640 107 642 117
rect 672 107 674 117
rect 704 107 706 117
rect 736 107 738 117
rect 768 107 770 117
rect 800 107 802 117
rect 832 107 834 117
rect 864 107 866 117
rect 896 107 898 117
rect 936 107 938 117
rect 976 107 978 117
rect 1016 107 1018 117
rect 1064 107 1066 117
rect 1104 107 1106 117
rect 1144 107 1146 117
rect 166 106 172 107
rect 166 102 167 106
rect 171 102 172 106
rect 166 101 172 102
rect 198 106 204 107
rect 198 102 199 106
rect 203 102 204 106
rect 198 101 204 102
rect 230 106 236 107
rect 230 102 231 106
rect 235 102 236 106
rect 230 101 236 102
rect 262 106 268 107
rect 262 102 263 106
rect 267 102 268 106
rect 262 101 268 102
rect 294 106 300 107
rect 294 102 295 106
rect 299 102 300 106
rect 294 101 300 102
rect 326 106 332 107
rect 326 102 327 106
rect 331 102 332 106
rect 326 101 332 102
rect 358 106 364 107
rect 358 102 359 106
rect 363 102 364 106
rect 358 101 364 102
rect 390 106 396 107
rect 390 102 391 106
rect 395 102 396 106
rect 390 101 396 102
rect 422 106 428 107
rect 438 106 444 107
rect 462 106 468 107
rect 478 106 484 107
rect 502 106 508 107
rect 422 102 423 106
rect 427 102 428 106
rect 422 101 428 102
rect 462 102 463 106
rect 467 102 468 106
rect 462 101 468 102
rect 502 102 503 106
rect 507 102 508 106
rect 502 101 508 102
rect 542 106 548 107
rect 542 102 543 106
rect 547 102 548 106
rect 542 101 548 102
rect 574 106 580 107
rect 574 102 575 106
rect 579 102 580 106
rect 574 101 580 102
rect 606 106 612 107
rect 606 102 607 106
rect 611 102 612 106
rect 606 101 612 102
rect 638 106 644 107
rect 638 102 639 106
rect 643 102 644 106
rect 638 101 644 102
rect 670 106 676 107
rect 670 102 671 106
rect 675 102 676 106
rect 670 101 676 102
rect 702 106 708 107
rect 702 102 703 106
rect 707 102 708 106
rect 702 101 708 102
rect 734 106 740 107
rect 734 102 735 106
rect 739 102 740 106
rect 734 101 740 102
rect 766 106 772 107
rect 766 102 767 106
rect 771 102 772 106
rect 766 101 772 102
rect 798 106 804 107
rect 798 102 799 106
rect 803 102 804 106
rect 798 101 804 102
rect 830 106 836 107
rect 830 102 831 106
rect 835 102 836 106
rect 830 101 836 102
rect 862 106 868 107
rect 862 102 863 106
rect 867 102 868 106
rect 862 101 868 102
rect 894 106 900 107
rect 894 102 895 106
rect 899 102 900 106
rect 894 101 900 102
rect 934 106 940 107
rect 934 102 935 106
rect 939 102 940 106
rect 934 101 940 102
rect 974 106 980 107
rect 974 102 975 106
rect 979 102 980 106
rect 974 101 980 102
rect 1014 106 1020 107
rect 1014 102 1015 106
rect 1019 102 1020 106
rect 1014 101 1020 102
rect 1062 106 1068 107
rect 1062 102 1063 106
rect 1067 102 1068 106
rect 1062 101 1068 102
rect 1102 106 1108 107
rect 1102 102 1103 106
rect 1107 102 1108 106
rect 1102 101 1108 102
rect 1142 106 1148 107
rect 1142 102 1143 106
rect 1147 102 1148 106
rect 1142 101 1148 102
rect 1160 96 1162 134
rect 1183 122 1187 123
rect 1183 117 1187 118
rect 1184 107 1186 117
rect 1200 112 1202 158
rect 1206 154 1212 155
rect 1206 150 1207 154
rect 1211 150 1212 154
rect 1206 149 1212 150
rect 1278 154 1284 155
rect 1278 150 1279 154
rect 1283 150 1284 154
rect 1278 149 1284 150
rect 1350 154 1356 155
rect 1350 150 1351 154
rect 1355 150 1356 154
rect 1350 149 1356 150
rect 1208 123 1210 149
rect 1280 123 1282 149
rect 1352 123 1354 149
rect 1368 148 1370 186
rect 1414 185 1420 186
rect 1414 181 1415 185
rect 1419 181 1420 185
rect 1414 180 1420 181
rect 1415 178 1419 180
rect 1415 173 1419 174
rect 1423 178 1427 179
rect 1423 172 1427 174
rect 1422 171 1428 172
rect 1422 167 1423 171
rect 1427 167 1428 171
rect 1422 166 1428 167
rect 1436 164 1438 202
rect 1456 192 1458 206
rect 1472 203 1474 213
rect 1470 202 1476 203
rect 1470 198 1471 202
rect 1475 198 1476 202
rect 1470 197 1476 198
rect 1484 192 1486 222
rect 1520 219 1522 229
rect 1576 219 1578 229
rect 1624 219 1626 229
rect 1636 220 1638 238
rect 1662 232 1668 233
rect 1662 228 1663 232
rect 1667 228 1668 232
rect 1662 227 1668 228
rect 1634 219 1640 220
rect 1664 219 1666 227
rect 1519 218 1523 219
rect 1519 213 1523 214
rect 1527 218 1531 219
rect 1527 213 1531 214
rect 1575 218 1579 219
rect 1575 213 1579 214
rect 1583 218 1587 219
rect 1583 213 1587 214
rect 1623 218 1627 219
rect 1634 215 1635 219
rect 1639 215 1640 219
rect 1634 214 1640 215
rect 1663 218 1667 219
rect 1623 213 1627 214
rect 1663 213 1667 214
rect 1528 203 1530 213
rect 1584 203 1586 213
rect 1624 203 1626 213
rect 1664 205 1666 213
rect 1662 204 1668 205
rect 1526 202 1532 203
rect 1526 198 1527 202
rect 1531 198 1532 202
rect 1526 197 1532 198
rect 1582 202 1588 203
rect 1582 198 1583 202
rect 1587 198 1588 202
rect 1582 197 1588 198
rect 1622 202 1628 203
rect 1622 198 1623 202
rect 1627 198 1628 202
rect 1662 200 1663 204
rect 1667 200 1668 204
rect 1662 199 1668 200
rect 1622 197 1628 198
rect 1454 191 1460 192
rect 1454 187 1455 191
rect 1459 187 1460 191
rect 1454 186 1460 187
rect 1482 191 1488 192
rect 1482 187 1483 191
rect 1487 187 1488 191
rect 1482 186 1488 187
rect 1638 191 1644 192
rect 1638 187 1639 191
rect 1643 187 1644 191
rect 1638 186 1644 187
rect 1662 187 1668 188
rect 1470 185 1476 186
rect 1470 181 1471 185
rect 1475 181 1476 185
rect 1470 180 1476 181
rect 1526 185 1532 186
rect 1526 181 1527 185
rect 1531 181 1532 185
rect 1526 180 1532 181
rect 1582 185 1588 186
rect 1582 181 1583 185
rect 1587 181 1588 185
rect 1582 180 1588 181
rect 1622 185 1628 186
rect 1622 181 1623 185
rect 1627 181 1628 185
rect 1622 180 1628 181
rect 1471 178 1475 180
rect 1471 173 1475 174
rect 1495 178 1499 179
rect 1495 172 1499 174
rect 1527 178 1531 180
rect 1527 173 1531 174
rect 1567 178 1571 179
rect 1567 172 1571 174
rect 1583 178 1587 180
rect 1583 173 1587 174
rect 1623 178 1627 180
rect 1623 172 1627 174
rect 1494 171 1500 172
rect 1494 167 1495 171
rect 1499 167 1500 171
rect 1494 166 1500 167
rect 1566 171 1572 172
rect 1566 167 1567 171
rect 1571 167 1572 171
rect 1566 166 1572 167
rect 1622 171 1628 172
rect 1622 167 1623 171
rect 1627 167 1628 171
rect 1622 166 1628 167
rect 1434 163 1440 164
rect 1434 159 1435 163
rect 1439 159 1440 163
rect 1434 158 1440 159
rect 1422 154 1428 155
rect 1422 150 1423 154
rect 1427 150 1428 154
rect 1422 149 1428 150
rect 1494 154 1500 155
rect 1494 150 1495 154
rect 1499 150 1500 154
rect 1494 149 1500 150
rect 1566 154 1572 155
rect 1566 150 1567 154
rect 1571 150 1572 154
rect 1566 149 1572 150
rect 1622 154 1628 155
rect 1622 150 1623 154
rect 1627 150 1628 154
rect 1622 149 1628 150
rect 1366 147 1372 148
rect 1366 143 1367 147
rect 1371 143 1372 147
rect 1366 142 1372 143
rect 1424 123 1426 149
rect 1496 123 1498 149
rect 1568 123 1570 149
rect 1574 147 1580 148
rect 1574 143 1575 147
rect 1579 143 1580 147
rect 1574 142 1580 143
rect 1207 122 1211 123
rect 1207 117 1211 118
rect 1223 122 1227 123
rect 1223 117 1227 118
rect 1263 122 1267 123
rect 1263 117 1267 118
rect 1279 122 1283 123
rect 1279 117 1283 118
rect 1295 122 1299 123
rect 1295 117 1299 118
rect 1335 122 1339 123
rect 1335 117 1339 118
rect 1351 122 1355 123
rect 1351 117 1355 118
rect 1375 122 1379 123
rect 1375 117 1379 118
rect 1415 122 1419 123
rect 1415 117 1419 118
rect 1423 122 1427 123
rect 1423 117 1427 118
rect 1455 122 1459 123
rect 1455 117 1459 118
rect 1495 122 1499 123
rect 1495 117 1499 118
rect 1503 122 1507 123
rect 1503 117 1507 118
rect 1551 122 1555 123
rect 1551 117 1555 118
rect 1567 122 1571 123
rect 1567 117 1571 118
rect 1198 111 1204 112
rect 1198 107 1199 111
rect 1203 107 1204 111
rect 1224 107 1226 117
rect 1264 107 1266 117
rect 1296 107 1298 117
rect 1336 107 1338 117
rect 1376 107 1378 117
rect 1416 107 1418 117
rect 1456 107 1458 117
rect 1504 107 1506 117
rect 1552 107 1554 117
rect 1182 106 1188 107
rect 1198 106 1204 107
rect 1222 106 1228 107
rect 1182 102 1183 106
rect 1187 102 1188 106
rect 1182 101 1188 102
rect 1222 102 1223 106
rect 1227 102 1228 106
rect 1222 101 1228 102
rect 1262 106 1268 107
rect 1262 102 1263 106
rect 1267 102 1268 106
rect 1262 101 1268 102
rect 1294 106 1300 107
rect 1294 102 1295 106
rect 1299 102 1300 106
rect 1294 101 1300 102
rect 1334 106 1340 107
rect 1334 102 1335 106
rect 1339 102 1340 106
rect 1334 101 1340 102
rect 1374 106 1380 107
rect 1374 102 1375 106
rect 1379 102 1380 106
rect 1374 101 1380 102
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1454 106 1460 107
rect 1454 102 1455 106
rect 1459 102 1460 106
rect 1454 101 1460 102
rect 1502 106 1508 107
rect 1502 102 1503 106
rect 1507 102 1508 106
rect 1502 101 1508 102
rect 1550 106 1556 107
rect 1550 102 1551 106
rect 1555 102 1556 106
rect 1550 101 1556 102
rect 150 95 156 96
rect 110 91 116 92
rect 110 87 111 91
rect 115 87 116 91
rect 150 91 151 95
rect 155 91 156 95
rect 150 90 156 91
rect 1158 95 1164 96
rect 1158 91 1159 95
rect 1163 91 1164 95
rect 1158 90 1164 91
rect 1567 95 1573 96
rect 1567 91 1568 95
rect 1572 94 1573 95
rect 1576 94 1578 142
rect 1624 123 1626 149
rect 1640 148 1642 186
rect 1662 183 1663 187
rect 1667 183 1668 187
rect 1662 182 1668 183
rect 1664 179 1666 182
rect 1663 178 1667 179
rect 1663 173 1667 174
rect 1664 170 1666 173
rect 1662 169 1668 170
rect 1662 165 1663 169
rect 1667 165 1668 169
rect 1662 164 1668 165
rect 1662 152 1668 153
rect 1662 148 1663 152
rect 1667 148 1668 152
rect 1638 147 1644 148
rect 1662 147 1668 148
rect 1638 143 1639 147
rect 1643 143 1644 147
rect 1638 142 1644 143
rect 1664 123 1666 147
rect 1591 122 1595 123
rect 1591 117 1595 118
rect 1623 122 1627 123
rect 1623 117 1627 118
rect 1663 122 1667 123
rect 1663 117 1667 118
rect 1592 107 1594 117
rect 1624 107 1626 117
rect 1664 109 1666 117
rect 1662 108 1668 109
rect 1590 106 1596 107
rect 1590 102 1591 106
rect 1595 102 1596 106
rect 1590 101 1596 102
rect 1622 106 1628 107
rect 1622 102 1623 106
rect 1627 102 1628 106
rect 1662 104 1663 108
rect 1667 104 1668 108
rect 1662 103 1668 104
rect 1622 101 1628 102
rect 1572 92 1578 94
rect 1572 91 1573 92
rect 1567 90 1573 91
rect 1662 91 1668 92
rect 110 86 116 87
rect 134 89 140 90
rect 112 83 114 86
rect 134 85 135 89
rect 139 85 140 89
rect 134 84 140 85
rect 166 89 172 90
rect 166 85 167 89
rect 171 85 172 89
rect 166 84 172 85
rect 198 89 204 90
rect 198 85 199 89
rect 203 85 204 89
rect 198 84 204 85
rect 230 89 236 90
rect 230 85 231 89
rect 235 85 236 89
rect 230 84 236 85
rect 262 89 268 90
rect 262 85 263 89
rect 267 85 268 89
rect 262 84 268 85
rect 294 89 300 90
rect 294 85 295 89
rect 299 85 300 89
rect 294 84 300 85
rect 326 89 332 90
rect 326 85 327 89
rect 331 85 332 89
rect 326 84 332 85
rect 358 89 364 90
rect 358 85 359 89
rect 363 85 364 89
rect 358 84 364 85
rect 390 89 396 90
rect 390 85 391 89
rect 395 85 396 89
rect 390 84 396 85
rect 422 89 428 90
rect 422 85 423 89
rect 427 85 428 89
rect 422 84 428 85
rect 462 89 468 90
rect 462 85 463 89
rect 467 85 468 89
rect 462 84 468 85
rect 502 89 508 90
rect 502 85 503 89
rect 507 85 508 89
rect 502 84 508 85
rect 542 89 548 90
rect 542 85 543 89
rect 547 85 548 89
rect 542 84 548 85
rect 574 89 580 90
rect 574 85 575 89
rect 579 85 580 89
rect 574 84 580 85
rect 606 89 612 90
rect 606 85 607 89
rect 611 85 612 89
rect 606 84 612 85
rect 638 89 644 90
rect 638 85 639 89
rect 643 85 644 89
rect 638 84 644 85
rect 670 89 676 90
rect 670 85 671 89
rect 675 85 676 89
rect 670 84 676 85
rect 702 89 708 90
rect 702 85 703 89
rect 707 85 708 89
rect 702 84 708 85
rect 734 89 740 90
rect 734 85 735 89
rect 739 85 740 89
rect 734 84 740 85
rect 766 89 772 90
rect 766 85 767 89
rect 771 85 772 89
rect 766 84 772 85
rect 798 89 804 90
rect 798 85 799 89
rect 803 85 804 89
rect 798 84 804 85
rect 830 89 836 90
rect 830 85 831 89
rect 835 85 836 89
rect 830 84 836 85
rect 862 89 868 90
rect 862 85 863 89
rect 867 85 868 89
rect 862 84 868 85
rect 894 89 900 90
rect 894 85 895 89
rect 899 85 900 89
rect 894 84 900 85
rect 934 89 940 90
rect 934 85 935 89
rect 939 85 940 89
rect 934 84 940 85
rect 974 89 980 90
rect 974 85 975 89
rect 979 85 980 89
rect 974 84 980 85
rect 1014 89 1020 90
rect 1014 85 1015 89
rect 1019 85 1020 89
rect 1014 84 1020 85
rect 1062 89 1068 90
rect 1062 85 1063 89
rect 1067 85 1068 89
rect 1062 84 1068 85
rect 1102 89 1108 90
rect 1102 85 1103 89
rect 1107 85 1108 89
rect 1102 84 1108 85
rect 1142 89 1148 90
rect 1142 85 1143 89
rect 1147 85 1148 89
rect 1142 84 1148 85
rect 1182 89 1188 90
rect 1182 85 1183 89
rect 1187 85 1188 89
rect 1182 84 1188 85
rect 1222 89 1228 90
rect 1222 85 1223 89
rect 1227 85 1228 89
rect 1222 84 1228 85
rect 1262 89 1268 90
rect 1262 85 1263 89
rect 1267 85 1268 89
rect 1262 84 1268 85
rect 1294 89 1300 90
rect 1294 85 1295 89
rect 1299 85 1300 89
rect 1294 84 1300 85
rect 1334 89 1340 90
rect 1334 85 1335 89
rect 1339 85 1340 89
rect 1334 84 1340 85
rect 1374 89 1380 90
rect 1374 85 1375 89
rect 1379 85 1380 89
rect 1374 84 1380 85
rect 1414 89 1420 90
rect 1414 85 1415 89
rect 1419 85 1420 89
rect 1414 84 1420 85
rect 1454 89 1460 90
rect 1454 85 1455 89
rect 1459 85 1460 89
rect 1454 84 1460 85
rect 1502 89 1508 90
rect 1502 85 1503 89
rect 1507 85 1508 89
rect 1502 84 1508 85
rect 1550 89 1556 90
rect 1550 85 1551 89
rect 1555 85 1556 89
rect 1550 84 1556 85
rect 1590 89 1596 90
rect 1590 85 1591 89
rect 1595 85 1596 89
rect 1590 84 1596 85
rect 1622 89 1628 90
rect 1622 85 1623 89
rect 1627 85 1628 89
rect 1662 87 1663 91
rect 1667 87 1668 91
rect 1662 86 1668 87
rect 1622 84 1628 85
rect 111 82 115 83
rect 111 77 115 78
rect 135 82 139 84
rect 135 77 139 78
rect 167 82 171 84
rect 167 77 171 78
rect 199 82 203 84
rect 199 77 203 78
rect 231 82 235 84
rect 231 77 235 78
rect 263 82 267 84
rect 263 77 267 78
rect 295 82 299 84
rect 295 77 299 78
rect 327 82 331 84
rect 327 77 331 78
rect 359 82 363 84
rect 359 77 363 78
rect 391 82 395 84
rect 391 77 395 78
rect 423 82 427 84
rect 423 77 427 78
rect 463 82 467 84
rect 463 77 467 78
rect 503 82 507 84
rect 503 77 507 78
rect 543 82 547 84
rect 543 77 547 78
rect 575 82 579 84
rect 575 77 579 78
rect 607 82 611 84
rect 607 77 611 78
rect 639 82 643 84
rect 639 77 643 78
rect 671 82 675 84
rect 671 77 675 78
rect 703 82 707 84
rect 703 77 707 78
rect 735 82 739 84
rect 735 77 739 78
rect 767 82 771 84
rect 767 77 771 78
rect 799 82 803 84
rect 799 77 803 78
rect 831 82 835 84
rect 831 77 835 78
rect 863 82 867 84
rect 863 77 867 78
rect 895 82 899 84
rect 895 77 899 78
rect 935 82 939 84
rect 935 77 939 78
rect 975 82 979 84
rect 975 77 979 78
rect 1015 82 1019 84
rect 1015 77 1019 78
rect 1063 82 1067 84
rect 1063 77 1067 78
rect 1103 82 1107 84
rect 1103 77 1107 78
rect 1143 82 1147 84
rect 1143 77 1147 78
rect 1183 82 1187 84
rect 1183 77 1187 78
rect 1223 82 1227 84
rect 1223 77 1227 78
rect 1263 82 1267 84
rect 1263 77 1267 78
rect 1295 82 1299 84
rect 1295 77 1299 78
rect 1335 82 1339 84
rect 1335 77 1339 78
rect 1375 82 1379 84
rect 1375 77 1379 78
rect 1415 82 1419 84
rect 1415 77 1419 78
rect 1455 82 1459 84
rect 1455 77 1459 78
rect 1503 82 1507 84
rect 1503 77 1507 78
rect 1551 82 1555 84
rect 1551 77 1555 78
rect 1591 82 1595 84
rect 1591 77 1595 78
rect 1623 82 1627 84
rect 1664 83 1666 86
rect 1623 77 1627 78
rect 1663 82 1667 83
rect 1663 77 1667 78
<< m4c >>
rect 111 1714 115 1718
rect 255 1714 259 1718
rect 287 1714 291 1718
rect 319 1714 323 1718
rect 359 1714 363 1718
rect 407 1714 411 1718
rect 455 1714 459 1718
rect 503 1714 507 1718
rect 551 1714 555 1718
rect 607 1714 611 1718
rect 663 1714 667 1718
rect 727 1714 731 1718
rect 783 1714 787 1718
rect 839 1714 843 1718
rect 895 1714 899 1718
rect 951 1714 955 1718
rect 1007 1714 1011 1718
rect 1063 1714 1067 1718
rect 1119 1714 1123 1718
rect 111 1674 115 1678
rect 135 1674 139 1678
rect 167 1674 171 1678
rect 215 1674 219 1678
rect 255 1674 259 1678
rect 279 1674 283 1678
rect 287 1674 291 1678
rect 319 1674 323 1678
rect 343 1674 347 1678
rect 111 1634 115 1638
rect 135 1634 139 1638
rect 359 1674 363 1678
rect 407 1674 411 1678
rect 415 1674 419 1678
rect 455 1674 459 1678
rect 487 1674 491 1678
rect 503 1674 507 1678
rect 551 1674 555 1678
rect 559 1674 563 1678
rect 607 1674 611 1678
rect 631 1674 635 1678
rect 663 1674 667 1678
rect 711 1674 715 1678
rect 727 1674 731 1678
rect 783 1674 787 1678
rect 791 1674 795 1678
rect 167 1634 171 1638
rect 183 1634 187 1638
rect 215 1634 219 1638
rect 247 1634 251 1638
rect 279 1634 283 1638
rect 303 1634 307 1638
rect 343 1634 347 1638
rect 359 1634 363 1638
rect 415 1634 419 1638
rect 471 1634 475 1638
rect 487 1634 491 1638
rect 535 1634 539 1638
rect 559 1634 563 1638
rect 599 1634 603 1638
rect 111 1594 115 1598
rect 135 1594 139 1598
rect 167 1594 171 1598
rect 183 1594 187 1598
rect 223 1594 227 1598
rect 247 1594 251 1598
rect 279 1594 283 1598
rect 303 1594 307 1598
rect 335 1594 339 1598
rect 359 1594 363 1598
rect 383 1594 387 1598
rect 415 1594 419 1598
rect 431 1594 435 1598
rect 111 1554 115 1558
rect 135 1554 139 1558
rect 167 1554 171 1558
rect 215 1554 219 1558
rect 223 1554 227 1558
rect 263 1554 267 1558
rect 279 1554 283 1558
rect 311 1554 315 1558
rect 335 1554 339 1558
rect 359 1554 363 1558
rect 471 1594 475 1598
rect 479 1594 483 1598
rect 631 1634 635 1638
rect 663 1634 667 1638
rect 839 1674 843 1678
rect 871 1674 875 1678
rect 1175 1714 1179 1718
rect 1231 1714 1235 1718
rect 1287 1714 1291 1718
rect 1335 1714 1339 1718
rect 1375 1714 1379 1718
rect 1423 1714 1427 1718
rect 1471 1714 1475 1718
rect 1519 1714 1523 1718
rect 1663 1714 1667 1718
rect 895 1674 899 1678
rect 951 1674 955 1678
rect 1007 1674 1011 1678
rect 1031 1674 1035 1678
rect 1063 1674 1067 1678
rect 1103 1674 1107 1678
rect 1119 1674 1123 1678
rect 1175 1674 1179 1678
rect 711 1634 715 1638
rect 727 1634 731 1638
rect 791 1634 795 1638
rect 799 1634 803 1638
rect 871 1634 875 1638
rect 943 1634 947 1638
rect 951 1634 955 1638
rect 535 1594 539 1598
rect 599 1594 603 1598
rect 663 1594 667 1598
rect 727 1594 731 1598
rect 383 1554 387 1558
rect 407 1554 411 1558
rect 431 1554 435 1558
rect 455 1554 459 1558
rect 479 1554 483 1558
rect 511 1554 515 1558
rect 535 1554 539 1558
rect 567 1554 571 1558
rect 111 1510 115 1514
rect 135 1510 139 1514
rect 799 1594 803 1598
rect 1023 1634 1027 1638
rect 1031 1634 1035 1638
rect 1103 1634 1107 1638
rect 1231 1674 1235 1678
rect 1247 1674 1251 1678
rect 1287 1674 1291 1678
rect 1319 1674 1323 1678
rect 1335 1674 1339 1678
rect 1375 1674 1379 1678
rect 1391 1674 1395 1678
rect 1423 1674 1427 1678
rect 1175 1634 1179 1638
rect 1247 1634 1251 1638
rect 1319 1634 1323 1638
rect 871 1594 875 1598
rect 943 1594 947 1598
rect 951 1594 955 1598
rect 1023 1594 1027 1598
rect 599 1554 603 1558
rect 631 1554 635 1558
rect 663 1554 667 1558
rect 695 1554 699 1558
rect 727 1554 731 1558
rect 759 1554 763 1558
rect 799 1554 803 1558
rect 831 1554 835 1558
rect 1039 1594 1043 1598
rect 1103 1594 1107 1598
rect 1119 1594 1123 1598
rect 1175 1594 1179 1598
rect 1199 1594 1203 1598
rect 1247 1594 1251 1598
rect 1279 1594 1283 1598
rect 1455 1674 1459 1678
rect 1471 1674 1475 1678
rect 1519 1674 1523 1678
rect 1583 1674 1587 1678
rect 1623 1674 1627 1678
rect 1663 1674 1667 1678
rect 1391 1634 1395 1638
rect 1399 1634 1403 1638
rect 1455 1634 1459 1638
rect 1479 1634 1483 1638
rect 1519 1634 1523 1638
rect 1319 1594 1323 1598
rect 1351 1594 1355 1598
rect 1399 1594 1403 1598
rect 1415 1594 1419 1598
rect 871 1554 875 1558
rect 919 1554 923 1558
rect 951 1554 955 1558
rect 1007 1554 1011 1558
rect 1039 1554 1043 1558
rect 1095 1554 1099 1558
rect 1119 1554 1123 1558
rect 1183 1554 1187 1558
rect 1199 1554 1203 1558
rect 1263 1554 1267 1558
rect 1279 1554 1283 1558
rect 167 1510 171 1514
rect 215 1510 219 1514
rect 223 1510 227 1514
rect 263 1510 267 1514
rect 295 1510 299 1514
rect 311 1510 315 1514
rect 359 1510 363 1514
rect 375 1510 379 1514
rect 407 1510 411 1514
rect 455 1510 459 1514
rect 511 1510 515 1514
rect 527 1510 531 1514
rect 567 1510 571 1514
rect 599 1510 603 1514
rect 631 1510 635 1514
rect 671 1510 675 1514
rect 695 1510 699 1514
rect 743 1510 747 1514
rect 759 1510 763 1514
rect 111 1470 115 1474
rect 135 1470 139 1474
rect 167 1470 171 1474
rect 223 1470 227 1474
rect 295 1470 299 1474
rect 375 1470 379 1474
rect 455 1470 459 1474
rect 527 1470 531 1474
rect 815 1510 819 1514
rect 831 1510 835 1514
rect 879 1510 883 1514
rect 1335 1554 1339 1558
rect 1351 1554 1355 1558
rect 1471 1594 1475 1598
rect 1479 1594 1483 1598
rect 1527 1594 1531 1598
rect 1559 1634 1563 1638
rect 1583 1634 1587 1638
rect 1623 1634 1627 1638
rect 1663 1634 1667 1638
rect 1559 1594 1563 1598
rect 1583 1594 1587 1598
rect 1623 1594 1627 1598
rect 1407 1554 1411 1558
rect 1415 1554 1419 1558
rect 1471 1554 1475 1558
rect 1527 1554 1531 1558
rect 1583 1554 1587 1558
rect 919 1510 923 1514
rect 943 1510 947 1514
rect 599 1470 603 1474
rect 663 1470 667 1474
rect 671 1470 675 1474
rect 719 1470 723 1474
rect 743 1470 747 1474
rect 783 1470 787 1474
rect 111 1426 115 1430
rect 135 1426 139 1430
rect 167 1426 171 1430
rect 215 1426 219 1430
rect 223 1426 227 1430
rect 287 1426 291 1430
rect 295 1426 299 1430
rect 359 1426 363 1430
rect 375 1426 379 1430
rect 439 1426 443 1430
rect 455 1426 459 1430
rect 1663 1594 1667 1598
rect 1623 1554 1627 1558
rect 1663 1554 1667 1558
rect 1007 1510 1011 1514
rect 1063 1510 1067 1514
rect 1095 1510 1099 1514
rect 1111 1510 1115 1514
rect 1151 1510 1155 1514
rect 1183 1510 1187 1514
rect 1215 1510 1219 1514
rect 1255 1510 1259 1514
rect 1263 1510 1267 1514
rect 1295 1510 1299 1514
rect 1335 1510 1339 1514
rect 1351 1510 1355 1514
rect 1407 1510 1411 1514
rect 1415 1510 1419 1514
rect 1471 1510 1475 1514
rect 1487 1510 1491 1514
rect 1527 1510 1531 1514
rect 1567 1510 1571 1514
rect 1583 1510 1587 1514
rect 1623 1510 1627 1514
rect 815 1470 819 1474
rect 847 1470 851 1474
rect 879 1470 883 1474
rect 903 1470 907 1474
rect 943 1470 947 1474
rect 959 1470 963 1474
rect 1007 1470 1011 1474
rect 1015 1470 1019 1474
rect 1663 1510 1667 1514
rect 1063 1470 1067 1474
rect 1071 1470 1075 1474
rect 1111 1470 1115 1474
rect 1119 1470 1123 1474
rect 1151 1470 1155 1474
rect 1159 1470 1163 1474
rect 1183 1470 1187 1474
rect 1207 1470 1211 1474
rect 1215 1470 1219 1474
rect 1255 1470 1259 1474
rect 1263 1470 1267 1474
rect 1295 1470 1299 1474
rect 1327 1470 1331 1474
rect 1351 1470 1355 1474
rect 1399 1470 1403 1474
rect 1415 1470 1419 1474
rect 1479 1470 1483 1474
rect 1487 1470 1491 1474
rect 1559 1470 1563 1474
rect 519 1426 523 1430
rect 527 1426 531 1430
rect 599 1426 603 1430
rect 663 1426 667 1430
rect 679 1426 683 1430
rect 719 1426 723 1430
rect 759 1426 763 1430
rect 783 1426 787 1430
rect 831 1426 835 1430
rect 847 1426 851 1430
rect 111 1386 115 1390
rect 135 1386 139 1390
rect 167 1386 171 1390
rect 215 1386 219 1390
rect 223 1386 227 1390
rect 287 1386 291 1390
rect 359 1386 363 1390
rect 431 1386 435 1390
rect 439 1386 443 1390
rect 503 1386 507 1390
rect 519 1386 523 1390
rect 583 1386 587 1390
rect 599 1386 603 1390
rect 663 1386 667 1390
rect 679 1386 683 1390
rect 743 1386 747 1390
rect 1567 1470 1571 1474
rect 1623 1470 1627 1474
rect 1663 1470 1667 1474
rect 903 1426 907 1430
rect 959 1426 963 1430
rect 967 1426 971 1430
rect 1015 1426 1019 1430
rect 1031 1426 1035 1430
rect 1071 1426 1075 1430
rect 1103 1426 1107 1430
rect 1119 1426 1123 1430
rect 1159 1426 1163 1430
rect 1167 1426 1171 1430
rect 1207 1426 1211 1430
rect 1231 1426 1235 1430
rect 1263 1426 1267 1430
rect 1295 1426 1299 1430
rect 1327 1426 1331 1430
rect 1359 1426 1363 1430
rect 1399 1426 1403 1430
rect 1415 1426 1419 1430
rect 1463 1426 1467 1430
rect 1479 1426 1483 1430
rect 1503 1426 1507 1430
rect 1551 1426 1555 1430
rect 1559 1426 1563 1430
rect 1591 1426 1595 1430
rect 1623 1426 1627 1430
rect 1663 1426 1667 1430
rect 759 1386 763 1390
rect 815 1386 819 1390
rect 831 1386 835 1390
rect 887 1386 891 1390
rect 903 1386 907 1390
rect 959 1386 963 1390
rect 967 1386 971 1390
rect 1031 1386 1035 1390
rect 1103 1386 1107 1390
rect 1167 1386 1171 1390
rect 1175 1386 1179 1390
rect 1231 1386 1235 1390
rect 1239 1386 1243 1390
rect 1295 1386 1299 1390
rect 111 1346 115 1350
rect 135 1346 139 1350
rect 167 1346 171 1350
rect 183 1346 187 1350
rect 111 1302 115 1306
rect 135 1302 139 1306
rect 223 1346 227 1350
rect 239 1346 243 1350
rect 287 1346 291 1350
rect 295 1346 299 1350
rect 351 1346 355 1350
rect 359 1346 363 1350
rect 399 1346 403 1350
rect 431 1346 435 1350
rect 455 1346 459 1350
rect 503 1346 507 1350
rect 511 1346 515 1350
rect 567 1346 571 1350
rect 583 1346 587 1350
rect 631 1346 635 1350
rect 663 1346 667 1350
rect 695 1346 699 1350
rect 183 1302 187 1306
rect 231 1302 235 1306
rect 239 1302 243 1306
rect 279 1302 283 1306
rect 295 1302 299 1306
rect 327 1302 331 1306
rect 351 1302 355 1306
rect 375 1302 379 1306
rect 111 1262 115 1266
rect 135 1262 139 1266
rect 167 1262 171 1266
rect 183 1262 187 1266
rect 223 1262 227 1266
rect 231 1262 235 1266
rect 111 1218 115 1222
rect 135 1218 139 1222
rect 279 1262 283 1266
rect 399 1302 403 1306
rect 431 1302 435 1306
rect 455 1302 459 1306
rect 487 1302 491 1306
rect 511 1302 515 1306
rect 543 1302 547 1306
rect 567 1302 571 1306
rect 607 1302 611 1306
rect 1303 1386 1307 1390
rect 1359 1386 1363 1390
rect 1367 1386 1371 1390
rect 1415 1386 1419 1390
rect 1431 1386 1435 1390
rect 1463 1386 1467 1390
rect 1495 1386 1499 1390
rect 1503 1386 1507 1390
rect 1551 1386 1555 1390
rect 1567 1386 1571 1390
rect 1591 1386 1595 1390
rect 1623 1386 1627 1390
rect 1663 1386 1667 1390
rect 743 1346 747 1350
rect 759 1346 763 1350
rect 815 1346 819 1350
rect 823 1346 827 1350
rect 887 1346 891 1350
rect 959 1346 963 1350
rect 1023 1346 1027 1350
rect 1031 1346 1035 1350
rect 1087 1346 1091 1350
rect 1103 1346 1107 1350
rect 1151 1346 1155 1350
rect 1175 1346 1179 1350
rect 1215 1346 1219 1350
rect 1239 1346 1243 1350
rect 1279 1346 1283 1350
rect 1303 1346 1307 1350
rect 1343 1346 1347 1350
rect 1367 1346 1371 1350
rect 1407 1346 1411 1350
rect 1431 1346 1435 1350
rect 1479 1346 1483 1350
rect 631 1302 635 1306
rect 663 1302 667 1306
rect 695 1302 699 1306
rect 719 1302 723 1306
rect 759 1302 763 1306
rect 775 1302 779 1306
rect 823 1302 827 1306
rect 831 1302 835 1306
rect 887 1302 891 1306
rect 895 1302 899 1306
rect 959 1302 963 1306
rect 1023 1302 1027 1306
rect 1079 1302 1083 1306
rect 1087 1302 1091 1306
rect 327 1262 331 1266
rect 375 1262 379 1266
rect 383 1262 387 1266
rect 431 1262 435 1266
rect 439 1262 443 1266
rect 167 1218 171 1222
rect 223 1218 227 1222
rect 279 1218 283 1222
rect 327 1218 331 1222
rect 335 1218 339 1222
rect 383 1218 387 1222
rect 111 1174 115 1178
rect 135 1174 139 1178
rect 167 1174 171 1178
rect 223 1174 227 1178
rect 111 1130 115 1134
rect 135 1130 139 1134
rect 143 1130 147 1134
rect 279 1174 283 1178
rect 287 1174 291 1178
rect 487 1262 491 1266
rect 495 1262 499 1266
rect 543 1262 547 1266
rect 551 1262 555 1266
rect 607 1262 611 1266
rect 663 1262 667 1266
rect 719 1262 723 1266
rect 767 1262 771 1266
rect 775 1262 779 1266
rect 1143 1302 1147 1306
rect 1151 1302 1155 1306
rect 1207 1302 1211 1306
rect 1215 1302 1219 1306
rect 1279 1302 1283 1306
rect 1343 1302 1347 1306
rect 1359 1302 1363 1306
rect 1495 1346 1499 1350
rect 1559 1346 1563 1350
rect 1567 1346 1571 1350
rect 1623 1346 1627 1350
rect 1407 1302 1411 1306
rect 1447 1302 1451 1306
rect 1479 1302 1483 1306
rect 1543 1302 1547 1306
rect 1559 1302 1563 1306
rect 1623 1302 1627 1306
rect 815 1262 819 1266
rect 831 1262 835 1266
rect 871 1262 875 1266
rect 895 1262 899 1266
rect 927 1262 931 1266
rect 959 1262 963 1266
rect 983 1262 987 1266
rect 1023 1262 1027 1266
rect 1039 1262 1043 1266
rect 1079 1262 1083 1266
rect 1095 1262 1099 1266
rect 1143 1262 1147 1266
rect 431 1218 435 1222
rect 439 1218 443 1222
rect 487 1218 491 1222
rect 495 1218 499 1222
rect 543 1218 547 1222
rect 551 1218 555 1222
rect 599 1218 603 1222
rect 607 1218 611 1222
rect 655 1218 659 1222
rect 663 1218 667 1222
rect 711 1218 715 1222
rect 719 1218 723 1222
rect 767 1218 771 1222
rect 815 1218 819 1222
rect 823 1218 827 1222
rect 871 1218 875 1222
rect 887 1218 891 1222
rect 1663 1346 1667 1350
rect 1159 1262 1163 1266
rect 1207 1262 1211 1266
rect 1231 1262 1235 1266
rect 1279 1262 1283 1266
rect 1319 1262 1323 1266
rect 1359 1262 1363 1266
rect 1423 1262 1427 1266
rect 1447 1262 1451 1266
rect 1535 1262 1539 1266
rect 1543 1262 1547 1266
rect 1623 1262 1627 1266
rect 927 1218 931 1222
rect 951 1218 955 1222
rect 983 1218 987 1222
rect 1015 1218 1019 1222
rect 1039 1218 1043 1222
rect 1079 1218 1083 1222
rect 1095 1218 1099 1222
rect 1143 1218 1147 1222
rect 1159 1218 1163 1222
rect 1207 1218 1211 1222
rect 1231 1218 1235 1222
rect 1279 1218 1283 1222
rect 1319 1218 1323 1222
rect 1359 1218 1363 1222
rect 1423 1218 1427 1222
rect 1447 1218 1451 1222
rect 1535 1218 1539 1222
rect 1543 1218 1547 1222
rect 1623 1218 1627 1222
rect 1663 1302 1667 1306
rect 1663 1262 1667 1266
rect 1663 1218 1667 1222
rect 335 1174 339 1178
rect 351 1174 355 1178
rect 383 1174 387 1178
rect 415 1174 419 1178
rect 431 1174 435 1178
rect 471 1174 475 1178
rect 487 1174 491 1178
rect 535 1174 539 1178
rect 543 1174 547 1178
rect 599 1174 603 1178
rect 655 1174 659 1178
rect 663 1174 667 1178
rect 711 1174 715 1178
rect 727 1174 731 1178
rect 767 1174 771 1178
rect 783 1174 787 1178
rect 823 1174 827 1178
rect 839 1174 843 1178
rect 887 1174 891 1178
rect 903 1174 907 1178
rect 951 1174 955 1178
rect 967 1174 971 1178
rect 1015 1174 1019 1178
rect 167 1130 171 1134
rect 175 1130 179 1134
rect 215 1130 219 1134
rect 223 1130 227 1134
rect 271 1130 275 1134
rect 287 1130 291 1134
rect 335 1130 339 1134
rect 351 1130 355 1134
rect 399 1130 403 1134
rect 415 1130 419 1134
rect 463 1130 467 1134
rect 471 1130 475 1134
rect 111 1086 115 1090
rect 143 1086 147 1090
rect 175 1086 179 1090
rect 215 1086 219 1090
rect 247 1086 251 1090
rect 271 1086 275 1090
rect 279 1086 283 1090
rect 1031 1174 1035 1178
rect 1079 1174 1083 1178
rect 1095 1174 1099 1178
rect 1143 1174 1147 1178
rect 1159 1174 1163 1178
rect 1207 1174 1211 1178
rect 1215 1174 1219 1178
rect 527 1130 531 1134
rect 535 1130 539 1134
rect 599 1130 603 1134
rect 663 1130 667 1134
rect 727 1130 731 1134
rect 783 1130 787 1134
rect 791 1130 795 1134
rect 839 1130 843 1134
rect 855 1130 859 1134
rect 903 1130 907 1134
rect 911 1130 915 1134
rect 967 1130 971 1134
rect 1023 1130 1027 1134
rect 1031 1130 1035 1134
rect 1279 1174 1283 1178
rect 1343 1174 1347 1178
rect 1359 1174 1363 1178
rect 1407 1174 1411 1178
rect 1447 1174 1451 1178
rect 1479 1174 1483 1178
rect 1543 1174 1547 1178
rect 1559 1174 1563 1178
rect 1623 1174 1627 1178
rect 1663 1174 1667 1178
rect 1087 1130 1091 1134
rect 1095 1130 1099 1134
rect 1151 1130 1155 1134
rect 1159 1130 1163 1134
rect 1215 1130 1219 1134
rect 1279 1130 1283 1134
rect 1335 1130 1339 1134
rect 1343 1130 1347 1134
rect 1391 1130 1395 1134
rect 1407 1130 1411 1134
rect 1447 1130 1451 1134
rect 1479 1130 1483 1134
rect 1495 1130 1499 1134
rect 1543 1130 1547 1134
rect 1559 1130 1563 1134
rect 1591 1130 1595 1134
rect 1623 1130 1627 1134
rect 1663 1130 1667 1134
rect 311 1086 315 1090
rect 335 1086 339 1090
rect 351 1086 355 1090
rect 391 1086 395 1090
rect 399 1086 403 1090
rect 439 1086 443 1090
rect 463 1086 467 1090
rect 503 1086 507 1090
rect 527 1086 531 1090
rect 575 1086 579 1090
rect 599 1086 603 1090
rect 655 1086 659 1090
rect 663 1086 667 1090
rect 727 1086 731 1090
rect 735 1086 739 1090
rect 791 1086 795 1090
rect 815 1086 819 1090
rect 855 1086 859 1090
rect 895 1086 899 1090
rect 111 1042 115 1046
rect 215 1042 219 1046
rect 247 1042 251 1046
rect 279 1042 283 1046
rect 295 1042 299 1046
rect 311 1042 315 1046
rect 327 1042 331 1046
rect 351 1042 355 1046
rect 359 1042 363 1046
rect 391 1042 395 1046
rect 423 1042 427 1046
rect 439 1042 443 1046
rect 455 1042 459 1046
rect 503 1042 507 1046
rect 559 1042 563 1046
rect 575 1042 579 1046
rect 631 1042 635 1046
rect 655 1042 659 1046
rect 711 1042 715 1046
rect 735 1042 739 1046
rect 799 1042 803 1046
rect 911 1086 915 1090
rect 967 1086 971 1090
rect 1023 1086 1027 1090
rect 1039 1086 1043 1090
rect 1087 1086 1091 1090
rect 1111 1086 1115 1090
rect 1151 1086 1155 1090
rect 1175 1086 1179 1090
rect 1215 1086 1219 1090
rect 1239 1086 1243 1090
rect 1279 1086 1283 1090
rect 1303 1086 1307 1090
rect 1335 1086 1339 1090
rect 1359 1086 1363 1090
rect 815 1042 819 1046
rect 879 1042 883 1046
rect 895 1042 899 1046
rect 959 1042 963 1046
rect 967 1042 971 1046
rect 1031 1042 1035 1046
rect 1039 1042 1043 1046
rect 1095 1042 1099 1046
rect 1111 1042 1115 1046
rect 1159 1042 1163 1046
rect 1175 1042 1179 1046
rect 1223 1042 1227 1046
rect 1239 1042 1243 1046
rect 1279 1042 1283 1046
rect 1303 1042 1307 1046
rect 111 1002 115 1006
rect 247 1002 251 1006
rect 279 1002 283 1006
rect 295 1002 299 1006
rect 311 1002 315 1006
rect 327 1002 331 1006
rect 343 1002 347 1006
rect 359 1002 363 1006
rect 383 1002 387 1006
rect 391 1002 395 1006
rect 423 1002 427 1006
rect 455 1002 459 1006
rect 479 1002 483 1006
rect 503 1002 507 1006
rect 543 1002 547 1006
rect 559 1002 563 1006
rect 615 1002 619 1006
rect 631 1002 635 1006
rect 687 1002 691 1006
rect 711 1002 715 1006
rect 759 1002 763 1006
rect 799 1002 803 1006
rect 831 1002 835 1006
rect 879 1002 883 1006
rect 111 962 115 966
rect 167 962 171 966
rect 199 962 203 966
rect 239 962 243 966
rect 247 962 251 966
rect 279 962 283 966
rect 287 962 291 966
rect 311 962 315 966
rect 343 962 347 966
rect 383 962 387 966
rect 407 962 411 966
rect 423 962 427 966
rect 471 962 475 966
rect 479 962 483 966
rect 535 962 539 966
rect 543 962 547 966
rect 599 962 603 966
rect 615 962 619 966
rect 663 962 667 966
rect 687 962 691 966
rect 727 962 731 966
rect 759 962 763 966
rect 791 962 795 966
rect 1391 1086 1395 1090
rect 1415 1086 1419 1090
rect 1447 1086 1451 1090
rect 1463 1086 1467 1090
rect 1495 1086 1499 1090
rect 1503 1086 1507 1090
rect 1543 1086 1547 1090
rect 1551 1086 1555 1090
rect 1591 1086 1595 1090
rect 1623 1086 1627 1090
rect 1335 1042 1339 1046
rect 1359 1042 1363 1046
rect 1383 1042 1387 1046
rect 1415 1042 1419 1046
rect 1431 1042 1435 1046
rect 1463 1042 1467 1046
rect 1479 1042 1483 1046
rect 1503 1042 1507 1046
rect 1535 1042 1539 1046
rect 1551 1042 1555 1046
rect 1591 1042 1595 1046
rect 1663 1086 1667 1090
rect 1623 1042 1627 1046
rect 1663 1042 1667 1046
rect 903 1002 907 1006
rect 959 1002 963 1006
rect 967 1002 971 1006
rect 1031 1002 1035 1006
rect 1095 1002 1099 1006
rect 1159 1002 1163 1006
rect 1223 1002 1227 1006
rect 1279 1002 1283 1006
rect 1287 1002 1291 1006
rect 1335 1002 1339 1006
rect 1343 1002 1347 1006
rect 1383 1002 1387 1006
rect 1399 1002 1403 1006
rect 831 962 835 966
rect 847 962 851 966
rect 903 962 907 966
rect 911 962 915 966
rect 967 962 971 966
rect 975 962 979 966
rect 1031 962 1035 966
rect 1039 962 1043 966
rect 1095 962 1099 966
rect 1103 962 1107 966
rect 1159 962 1163 966
rect 1167 962 1171 966
rect 1223 962 1227 966
rect 111 918 115 922
rect 135 918 139 922
rect 167 918 171 922
rect 199 918 203 922
rect 207 918 211 922
rect 239 918 243 922
rect 271 918 275 922
rect 287 918 291 922
rect 335 918 339 922
rect 343 918 347 922
rect 407 918 411 922
rect 471 918 475 922
rect 535 918 539 922
rect 591 918 595 922
rect 599 918 603 922
rect 647 918 651 922
rect 663 918 667 922
rect 111 874 115 878
rect 135 874 139 878
rect 167 874 171 878
rect 207 874 211 878
rect 271 874 275 878
rect 335 874 339 878
rect 407 874 411 878
rect 111 834 115 838
rect 135 834 139 838
rect 471 874 475 878
rect 535 874 539 878
rect 591 874 595 878
rect 599 874 603 878
rect 647 874 651 878
rect 655 874 659 878
rect 703 918 707 922
rect 727 918 731 922
rect 751 918 755 922
rect 1231 962 1235 966
rect 1287 962 1291 966
rect 1431 1002 1435 1006
rect 1447 1002 1451 1006
rect 1479 1002 1483 1006
rect 1495 1002 1499 1006
rect 1535 1002 1539 1006
rect 1543 1002 1547 1006
rect 1591 1002 1595 1006
rect 1623 1002 1627 1006
rect 1343 962 1347 966
rect 1391 962 1395 966
rect 1399 962 1403 966
rect 1431 962 1435 966
rect 1447 962 1451 966
rect 1471 962 1475 966
rect 1495 962 1499 966
rect 1511 962 1515 966
rect 1543 962 1547 966
rect 1551 962 1555 966
rect 1591 962 1595 966
rect 1663 1002 1667 1006
rect 1623 962 1627 966
rect 1663 962 1667 966
rect 791 918 795 922
rect 799 918 803 922
rect 847 918 851 922
rect 903 918 907 922
rect 911 918 915 922
rect 959 918 963 922
rect 975 918 979 922
rect 1023 918 1027 922
rect 1039 918 1043 922
rect 1087 918 1091 922
rect 1103 918 1107 922
rect 1143 918 1147 922
rect 1167 918 1171 922
rect 703 874 707 878
rect 751 874 755 878
rect 799 874 803 878
rect 1199 918 1203 922
rect 1231 918 1235 922
rect 1255 918 1259 922
rect 1287 918 1291 922
rect 1319 918 1323 922
rect 1343 918 1347 922
rect 1383 918 1387 922
rect 1391 918 1395 922
rect 1431 918 1435 922
rect 1471 918 1475 922
rect 1511 918 1515 922
rect 1551 918 1555 922
rect 1591 918 1595 922
rect 1623 918 1627 922
rect 1663 918 1667 922
rect 847 874 851 878
rect 903 874 907 878
rect 959 874 963 878
rect 967 874 971 878
rect 1023 874 1027 878
rect 1039 874 1043 878
rect 1087 874 1091 878
rect 1103 874 1107 878
rect 1143 874 1147 878
rect 167 834 171 838
rect 207 834 211 838
rect 215 834 219 838
rect 271 834 275 838
rect 279 834 283 838
rect 335 834 339 838
rect 343 834 347 838
rect 407 834 411 838
rect 415 834 419 838
rect 471 834 475 838
rect 479 834 483 838
rect 535 834 539 838
rect 543 834 547 838
rect 599 834 603 838
rect 607 834 611 838
rect 111 790 115 794
rect 135 790 139 794
rect 167 790 171 794
rect 175 790 179 794
rect 215 790 219 794
rect 231 790 235 794
rect 279 790 283 794
rect 295 790 299 794
rect 343 790 347 794
rect 367 790 371 794
rect 415 790 419 794
rect 447 790 451 794
rect 479 790 483 794
rect 527 790 531 794
rect 111 750 115 754
rect 135 750 139 754
rect 175 750 179 754
rect 215 750 219 754
rect 231 750 235 754
rect 247 750 251 754
rect 279 750 283 754
rect 295 750 299 754
rect 655 834 659 838
rect 671 834 675 838
rect 703 834 707 838
rect 735 834 739 838
rect 751 834 755 838
rect 791 834 795 838
rect 799 834 803 838
rect 847 834 851 838
rect 903 834 907 838
rect 911 834 915 838
rect 967 834 971 838
rect 975 834 979 838
rect 1039 834 1043 838
rect 1167 874 1171 878
rect 1199 874 1203 878
rect 1231 874 1235 878
rect 1255 874 1259 878
rect 1287 874 1291 878
rect 1319 874 1323 878
rect 1343 874 1347 878
rect 1383 874 1387 878
rect 1399 874 1403 878
rect 1463 874 1467 878
rect 1663 874 1667 878
rect 1103 834 1107 838
rect 1111 834 1115 838
rect 1167 834 1171 838
rect 1183 834 1187 838
rect 1231 834 1235 838
rect 1247 834 1251 838
rect 1287 834 1291 838
rect 1311 834 1315 838
rect 1343 834 1347 838
rect 543 790 547 794
rect 607 790 611 794
rect 615 790 619 794
rect 671 790 675 794
rect 703 790 707 794
rect 735 790 739 794
rect 791 790 795 794
rect 847 790 851 794
rect 871 790 875 794
rect 911 790 915 794
rect 951 790 955 794
rect 975 790 979 794
rect 1023 790 1027 794
rect 1039 790 1043 794
rect 1095 790 1099 794
rect 1111 790 1115 794
rect 1167 790 1171 794
rect 1183 790 1187 794
rect 1231 790 1235 794
rect 1247 790 1251 794
rect 1295 790 1299 794
rect 319 750 323 754
rect 359 750 363 754
rect 367 750 371 754
rect 399 750 403 754
rect 439 750 443 754
rect 447 750 451 754
rect 487 750 491 754
rect 527 750 531 754
rect 543 750 547 754
rect 607 750 611 754
rect 615 750 619 754
rect 671 750 675 754
rect 111 706 115 710
rect 215 706 219 710
rect 247 706 251 710
rect 279 706 283 710
rect 311 706 315 710
rect 319 706 323 710
rect 343 706 347 710
rect 359 706 363 710
rect 703 750 707 754
rect 735 750 739 754
rect 791 750 795 754
rect 799 750 803 754
rect 863 750 867 754
rect 871 750 875 754
rect 375 706 379 710
rect 399 706 403 710
rect 407 706 411 710
rect 439 706 443 710
rect 471 706 475 710
rect 487 706 491 710
rect 503 706 507 710
rect 543 706 547 710
rect 591 706 595 710
rect 607 706 611 710
rect 647 706 651 710
rect 671 706 675 710
rect 703 706 707 710
rect 735 706 739 710
rect 759 706 763 710
rect 1367 834 1371 838
rect 1399 834 1403 838
rect 1423 834 1427 838
rect 1463 834 1467 838
rect 1479 834 1483 838
rect 1535 834 1539 838
rect 1591 834 1595 838
rect 1663 834 1667 838
rect 1311 790 1315 794
rect 1359 790 1363 794
rect 1367 790 1371 794
rect 1415 790 1419 794
rect 1423 790 1427 794
rect 1471 790 1475 794
rect 1479 790 1483 794
rect 1527 790 1531 794
rect 1535 790 1539 794
rect 1591 790 1595 794
rect 1663 790 1667 794
rect 927 750 931 754
rect 951 750 955 754
rect 991 750 995 754
rect 1023 750 1027 754
rect 1055 750 1059 754
rect 1095 750 1099 754
rect 1119 750 1123 754
rect 1167 750 1171 754
rect 1183 750 1187 754
rect 1231 750 1235 754
rect 1239 750 1243 754
rect 1295 750 1299 754
rect 1351 750 1355 754
rect 1359 750 1363 754
rect 1407 750 1411 754
rect 1415 750 1419 754
rect 1463 750 1467 754
rect 1471 750 1475 754
rect 799 706 803 710
rect 823 706 827 710
rect 863 706 867 710
rect 887 706 891 710
rect 927 706 931 710
rect 959 706 963 710
rect 1519 750 1523 754
rect 1527 750 1531 754
rect 1583 750 1587 754
rect 1591 750 1595 754
rect 1623 750 1627 754
rect 1663 750 1667 754
rect 991 706 995 710
rect 1023 706 1027 710
rect 1055 706 1059 710
rect 1087 706 1091 710
rect 1119 706 1123 710
rect 111 666 115 670
rect 279 666 283 670
rect 295 666 299 670
rect 311 666 315 670
rect 327 666 331 670
rect 343 666 347 670
rect 359 666 363 670
rect 375 666 379 670
rect 391 666 395 670
rect 407 666 411 670
rect 423 666 427 670
rect 439 666 443 670
rect 455 666 459 670
rect 471 666 475 670
rect 487 666 491 670
rect 503 666 507 670
rect 519 666 523 670
rect 543 666 547 670
rect 551 666 555 670
rect 591 666 595 670
rect 639 666 643 670
rect 647 666 651 670
rect 687 666 691 670
rect 703 666 707 670
rect 735 666 739 670
rect 759 666 763 670
rect 791 666 795 670
rect 823 666 827 670
rect 847 666 851 670
rect 887 666 891 670
rect 911 666 915 670
rect 111 626 115 630
rect 247 626 251 630
rect 279 626 283 630
rect 295 626 299 630
rect 319 626 323 630
rect 327 626 331 630
rect 359 626 363 630
rect 367 626 371 630
rect 391 626 395 630
rect 423 626 427 630
rect 455 626 459 630
rect 471 626 475 630
rect 487 626 491 630
rect 519 626 523 630
rect 551 626 555 630
rect 567 626 571 630
rect 591 626 595 630
rect 615 626 619 630
rect 639 626 643 630
rect 663 626 667 630
rect 687 626 691 630
rect 719 626 723 630
rect 735 626 739 630
rect 775 626 779 630
rect 791 626 795 630
rect 831 626 835 630
rect 959 666 963 670
rect 975 666 979 670
rect 1023 666 1027 670
rect 1159 706 1163 710
rect 1183 706 1187 710
rect 1223 706 1227 710
rect 1239 706 1243 710
rect 1287 706 1291 710
rect 1295 706 1299 710
rect 1351 706 1355 710
rect 1407 706 1411 710
rect 1415 706 1419 710
rect 1463 706 1467 710
rect 1471 706 1475 710
rect 1519 706 1523 710
rect 1527 706 1531 710
rect 1047 666 1051 670
rect 1087 666 1091 670
rect 1127 666 1131 670
rect 1159 666 1163 670
rect 1215 666 1219 670
rect 1223 666 1227 670
rect 1287 666 1291 670
rect 1295 666 1299 670
rect 1351 666 1355 670
rect 1383 666 1387 670
rect 1415 666 1419 670
rect 847 626 851 630
rect 895 626 899 630
rect 911 626 915 630
rect 967 626 971 630
rect 975 626 979 630
rect 1047 626 1051 630
rect 1127 626 1131 630
rect 111 586 115 590
rect 167 586 171 590
rect 215 586 219 590
rect 247 586 251 590
rect 271 586 275 590
rect 279 586 283 590
rect 319 586 323 590
rect 335 586 339 590
rect 367 586 371 590
rect 407 586 411 590
rect 423 586 427 590
rect 471 586 475 590
rect 487 586 491 590
rect 519 586 523 590
rect 559 586 563 590
rect 567 586 571 590
rect 615 586 619 590
rect 631 586 635 590
rect 663 586 667 590
rect 703 586 707 590
rect 719 586 723 590
rect 767 586 771 590
rect 775 586 779 590
rect 823 586 827 590
rect 831 586 835 590
rect 879 586 883 590
rect 895 586 899 590
rect 935 586 939 590
rect 967 586 971 590
rect 111 542 115 546
rect 135 542 139 546
rect 167 542 171 546
rect 199 542 203 546
rect 215 542 219 546
rect 231 542 235 546
rect 271 542 275 546
rect 279 542 283 546
rect 327 542 331 546
rect 335 542 339 546
rect 375 542 379 546
rect 407 542 411 546
rect 431 542 435 546
rect 487 542 491 546
rect 495 542 499 546
rect 559 542 563 546
rect 623 542 627 546
rect 631 542 635 546
rect 687 542 691 546
rect 703 542 707 546
rect 751 542 755 546
rect 767 542 771 546
rect 111 502 115 506
rect 135 502 139 506
rect 167 502 171 506
rect 199 502 203 506
rect 231 502 235 506
rect 239 502 243 506
rect 279 502 283 506
rect 287 502 291 506
rect 327 502 331 506
rect 375 502 379 506
rect 423 502 427 506
rect 431 502 435 506
rect 479 502 483 506
rect 111 462 115 466
rect 135 462 139 466
rect 151 462 155 466
rect 167 462 171 466
rect 199 462 203 466
rect 207 462 211 466
rect 239 462 243 466
rect 255 462 259 466
rect 111 422 115 426
rect 151 422 155 426
rect 175 422 179 426
rect 495 502 499 506
rect 543 502 547 506
rect 559 502 563 506
rect 615 502 619 506
rect 623 502 627 506
rect 815 542 819 546
rect 823 542 827 546
rect 879 542 883 546
rect 991 586 995 590
rect 1047 586 1051 590
rect 1103 586 1107 590
rect 1207 626 1211 630
rect 1215 626 1219 630
rect 1471 666 1475 670
rect 1583 706 1587 710
rect 1623 706 1627 710
rect 1663 706 1667 710
rect 1527 666 1531 670
rect 1559 666 1563 670
rect 1583 666 1587 670
rect 1623 666 1627 670
rect 1287 626 1291 630
rect 1295 626 1299 630
rect 1359 626 1363 630
rect 1383 626 1387 630
rect 1431 626 1435 630
rect 1471 626 1475 630
rect 1503 626 1507 630
rect 1559 626 1563 630
rect 1575 626 1579 630
rect 1127 586 1131 590
rect 1159 586 1163 590
rect 1207 586 1211 590
rect 1215 586 1219 590
rect 1271 586 1275 590
rect 1287 586 1291 590
rect 935 542 939 546
rect 943 542 947 546
rect 991 542 995 546
rect 1007 542 1011 546
rect 1047 542 1051 546
rect 1071 542 1075 546
rect 1103 542 1107 546
rect 1127 542 1131 546
rect 1159 542 1163 546
rect 1183 542 1187 546
rect 1663 666 1667 670
rect 1623 626 1627 630
rect 1663 626 1667 630
rect 1327 586 1331 590
rect 1359 586 1363 590
rect 1383 586 1387 590
rect 1431 586 1435 590
rect 1447 586 1451 590
rect 1503 586 1507 590
rect 1511 586 1515 590
rect 1575 586 1579 590
rect 1623 586 1627 590
rect 1663 586 1667 590
rect 1215 542 1219 546
rect 1231 542 1235 546
rect 1271 542 1275 546
rect 1279 542 1283 546
rect 1327 542 1331 546
rect 1335 542 1339 546
rect 1383 542 1387 546
rect 1391 542 1395 546
rect 1447 542 1451 546
rect 1511 542 1515 546
rect 687 502 691 506
rect 695 502 699 506
rect 751 502 755 506
rect 775 502 779 506
rect 287 462 291 466
rect 311 462 315 466
rect 327 462 331 466
rect 367 462 371 466
rect 375 462 379 466
rect 423 462 427 466
rect 439 462 443 466
rect 479 462 483 466
rect 519 462 523 466
rect 543 462 547 466
rect 599 462 603 466
rect 615 462 619 466
rect 679 462 683 466
rect 695 462 699 466
rect 1575 542 1579 546
rect 1623 542 1627 546
rect 1663 542 1667 546
rect 815 502 819 506
rect 847 502 851 506
rect 879 502 883 506
rect 919 502 923 506
rect 943 502 947 506
rect 983 502 987 506
rect 759 462 763 466
rect 775 462 779 466
rect 1007 502 1011 506
rect 1039 502 1043 506
rect 1071 502 1075 506
rect 1095 502 1099 506
rect 1127 502 1131 506
rect 1143 502 1147 506
rect 1183 502 1187 506
rect 1191 502 1195 506
rect 1231 502 1235 506
rect 1239 502 1243 506
rect 1279 502 1283 506
rect 1287 502 1291 506
rect 1335 502 1339 506
rect 1383 502 1387 506
rect 1391 502 1395 506
rect 1431 502 1435 506
rect 1447 502 1451 506
rect 1479 502 1483 506
rect 1511 502 1515 506
rect 1535 502 1539 506
rect 1575 502 1579 506
rect 1591 502 1595 506
rect 839 462 843 466
rect 847 462 851 466
rect 911 462 915 466
rect 919 462 923 466
rect 983 462 987 466
rect 1039 462 1043 466
rect 1055 462 1059 466
rect 1095 462 1099 466
rect 1127 462 1131 466
rect 1143 462 1147 466
rect 1191 462 1195 466
rect 1199 462 1203 466
rect 1239 462 1243 466
rect 1263 462 1267 466
rect 1287 462 1291 466
rect 1319 462 1323 466
rect 1335 462 1339 466
rect 1375 462 1379 466
rect 1383 462 1387 466
rect 1431 462 1435 466
rect 207 422 211 426
rect 223 422 227 426
rect 255 422 259 426
rect 271 422 275 426
rect 311 422 315 426
rect 319 422 323 426
rect 111 378 115 382
rect 135 378 139 382
rect 167 378 171 382
rect 175 378 179 382
rect 199 378 203 382
rect 223 378 227 382
rect 367 422 371 426
rect 415 422 419 426
rect 439 422 443 426
rect 471 422 475 426
rect 519 422 523 426
rect 527 422 531 426
rect 591 422 595 426
rect 599 422 603 426
rect 663 422 667 426
rect 679 422 683 426
rect 735 422 739 426
rect 759 422 763 426
rect 807 422 811 426
rect 239 378 243 382
rect 271 378 275 382
rect 295 378 299 382
rect 319 378 323 382
rect 351 378 355 382
rect 367 378 371 382
rect 407 378 411 382
rect 415 378 419 382
rect 463 378 467 382
rect 471 378 475 382
rect 519 378 523 382
rect 527 378 531 382
rect 575 378 579 382
rect 591 378 595 382
rect 631 378 635 382
rect 663 378 667 382
rect 111 338 115 342
rect 135 338 139 342
rect 167 338 171 342
rect 199 338 203 342
rect 207 338 211 342
rect 239 338 243 342
rect 111 298 115 302
rect 135 298 139 302
rect 263 338 267 342
rect 295 338 299 342
rect 327 338 331 342
rect 351 338 355 342
rect 391 338 395 342
rect 407 338 411 342
rect 455 338 459 342
rect 463 338 467 342
rect 687 378 691 382
rect 735 378 739 382
rect 743 378 747 382
rect 839 422 843 426
rect 871 422 875 426
rect 911 422 915 426
rect 935 422 939 426
rect 799 378 803 382
rect 807 378 811 382
rect 855 378 859 382
rect 871 378 875 382
rect 1479 462 1483 466
rect 1495 462 1499 466
rect 1623 502 1627 506
rect 1663 502 1667 506
rect 1535 462 1539 466
rect 1591 462 1595 466
rect 1623 462 1627 466
rect 1663 462 1667 466
rect 983 422 987 426
rect 991 422 995 426
rect 1039 422 1043 426
rect 1055 422 1059 426
rect 1087 422 1091 426
rect 1127 422 1131 426
rect 1167 422 1171 426
rect 1199 422 1203 426
rect 1207 422 1211 426
rect 1247 422 1251 426
rect 1263 422 1267 426
rect 1287 422 1291 426
rect 1319 422 1323 426
rect 1335 422 1339 426
rect 1375 422 1379 426
rect 1383 422 1387 426
rect 1431 422 1435 426
rect 1495 422 1499 426
rect 1663 422 1667 426
rect 919 378 923 382
rect 935 378 939 382
rect 983 378 987 382
rect 991 378 995 382
rect 1039 378 1043 382
rect 1087 378 1091 382
rect 1095 378 1099 382
rect 1127 378 1131 382
rect 1151 378 1155 382
rect 1167 378 1171 382
rect 1207 378 1211 382
rect 1247 378 1251 382
rect 1255 378 1259 382
rect 1287 378 1291 382
rect 1303 378 1307 382
rect 1335 378 1339 382
rect 1351 378 1355 382
rect 1383 378 1387 382
rect 1399 378 1403 382
rect 1447 378 1451 382
rect 1495 378 1499 382
rect 1543 378 1547 382
rect 1591 378 1595 382
rect 1623 378 1627 382
rect 1663 378 1667 382
rect 519 338 523 342
rect 575 338 579 342
rect 631 338 635 342
rect 687 338 691 342
rect 167 298 171 302
rect 207 298 211 302
rect 231 298 235 302
rect 263 298 267 302
rect 295 298 299 302
rect 327 298 331 302
rect 367 298 371 302
rect 391 298 395 302
rect 439 298 443 302
rect 111 254 115 258
rect 135 254 139 258
rect 167 254 171 258
rect 175 254 179 258
rect 231 254 235 258
rect 455 298 459 302
rect 503 298 507 302
rect 519 298 523 302
rect 567 298 571 302
rect 575 298 579 302
rect 743 338 747 342
rect 751 338 755 342
rect 799 338 803 342
rect 815 338 819 342
rect 855 338 859 342
rect 879 338 883 342
rect 919 338 923 342
rect 951 338 955 342
rect 983 338 987 342
rect 1031 338 1035 342
rect 1039 338 1043 342
rect 1095 338 1099 342
rect 1111 338 1115 342
rect 1151 338 1155 342
rect 1191 338 1195 342
rect 1207 338 1211 342
rect 1255 338 1259 342
rect 1271 338 1275 342
rect 1303 338 1307 342
rect 1343 338 1347 342
rect 1351 338 1355 342
rect 1399 338 1403 342
rect 1407 338 1411 342
rect 1447 338 1451 342
rect 1463 338 1467 342
rect 1495 338 1499 342
rect 1519 338 1523 342
rect 1543 338 1547 342
rect 1583 338 1587 342
rect 1591 338 1595 342
rect 1623 338 1627 342
rect 631 298 635 302
rect 687 298 691 302
rect 743 298 747 302
rect 247 254 251 258
rect 295 254 299 258
rect 111 214 115 218
rect 135 214 139 218
rect 319 254 323 258
rect 367 254 371 258
rect 383 254 387 258
rect 439 254 443 258
rect 447 254 451 258
rect 503 254 507 258
rect 519 254 523 258
rect 567 254 571 258
rect 591 254 595 258
rect 631 254 635 258
rect 663 254 667 258
rect 751 298 755 302
rect 807 298 811 302
rect 815 298 819 302
rect 879 298 883 302
rect 951 298 955 302
rect 1031 298 1035 302
rect 1111 298 1115 302
rect 1191 298 1195 302
rect 1263 298 1267 302
rect 1271 298 1275 302
rect 1663 338 1667 342
rect 1327 298 1331 302
rect 1343 298 1347 302
rect 1391 298 1395 302
rect 1407 298 1411 302
rect 1447 298 1451 302
rect 1463 298 1467 302
rect 1495 298 1499 302
rect 1519 298 1523 302
rect 1543 298 1547 302
rect 1583 298 1587 302
rect 1591 298 1595 302
rect 1623 298 1627 302
rect 1663 298 1667 302
rect 687 254 691 258
rect 743 254 747 258
rect 807 254 811 258
rect 823 254 827 258
rect 879 254 883 258
rect 895 254 899 258
rect 167 214 171 218
rect 175 214 179 218
rect 207 214 211 218
rect 247 214 251 218
rect 255 214 259 218
rect 303 214 307 218
rect 319 214 323 218
rect 343 214 347 218
rect 375 214 379 218
rect 383 214 387 218
rect 415 214 419 218
rect 447 214 451 218
rect 471 214 475 218
rect 519 214 523 218
rect 535 214 539 218
rect 111 174 115 178
rect 135 174 139 178
rect 167 174 171 178
rect 175 174 179 178
rect 207 174 211 178
rect 231 174 235 178
rect 255 174 259 178
rect 287 174 291 178
rect 111 118 115 122
rect 135 118 139 122
rect 951 254 955 258
rect 967 254 971 258
rect 1031 254 1035 258
rect 1087 254 1091 258
rect 1111 254 1115 258
rect 1143 254 1147 258
rect 1191 254 1195 258
rect 1199 254 1203 258
rect 1255 254 1259 258
rect 1263 254 1267 258
rect 1311 254 1315 258
rect 1327 254 1331 258
rect 1367 254 1371 258
rect 1391 254 1395 258
rect 1415 254 1419 258
rect 591 214 595 218
rect 615 214 619 218
rect 663 214 667 218
rect 695 214 699 218
rect 743 214 747 218
rect 775 214 779 218
rect 823 214 827 218
rect 855 214 859 218
rect 895 214 899 218
rect 927 214 931 218
rect 967 214 971 218
rect 999 214 1003 218
rect 1031 214 1035 218
rect 1071 214 1075 218
rect 1087 214 1091 218
rect 1143 214 1147 218
rect 1199 214 1203 218
rect 1215 214 1219 218
rect 1255 214 1259 218
rect 303 174 307 178
rect 343 174 347 178
rect 375 174 379 178
rect 399 174 403 178
rect 415 174 419 178
rect 455 174 459 178
rect 471 174 475 178
rect 511 174 515 178
rect 535 174 539 178
rect 575 174 579 178
rect 615 174 619 178
rect 639 174 643 178
rect 695 174 699 178
rect 703 174 707 178
rect 767 174 771 178
rect 775 174 779 178
rect 167 118 171 122
rect 175 118 179 122
rect 199 118 203 122
rect 231 118 235 122
rect 263 118 267 122
rect 287 118 291 122
rect 295 118 299 122
rect 327 118 331 122
rect 343 118 347 122
rect 359 118 363 122
rect 391 118 395 122
rect 399 118 403 122
rect 423 118 427 122
rect 455 118 459 122
rect 463 118 467 122
rect 1287 214 1291 218
rect 1311 214 1315 218
rect 1447 254 1451 258
rect 1463 254 1467 258
rect 1495 254 1499 258
rect 1519 254 1523 258
rect 1543 254 1547 258
rect 1575 254 1579 258
rect 1591 254 1595 258
rect 1623 254 1627 258
rect 1663 254 1667 258
rect 1351 214 1355 218
rect 1367 214 1371 218
rect 1415 214 1419 218
rect 1463 214 1467 218
rect 1471 214 1475 218
rect 831 174 835 178
rect 855 174 859 178
rect 895 174 899 178
rect 927 174 931 178
rect 951 174 955 178
rect 999 174 1003 178
rect 1015 174 1019 178
rect 1071 174 1075 178
rect 1079 174 1083 178
rect 1143 174 1147 178
rect 1207 174 1211 178
rect 1215 174 1219 178
rect 1279 174 1283 178
rect 1287 174 1291 178
rect 1351 174 1355 178
rect 503 118 507 122
rect 511 118 515 122
rect 543 118 547 122
rect 575 118 579 122
rect 607 118 611 122
rect 639 118 643 122
rect 671 118 675 122
rect 703 118 707 122
rect 735 118 739 122
rect 767 118 771 122
rect 799 118 803 122
rect 831 118 835 122
rect 863 118 867 122
rect 895 118 899 122
rect 935 118 939 122
rect 951 118 955 122
rect 975 118 979 122
rect 1015 118 1019 122
rect 1063 118 1067 122
rect 1079 118 1083 122
rect 1103 118 1107 122
rect 1143 118 1147 122
rect 1183 118 1187 122
rect 1415 174 1419 178
rect 1423 174 1427 178
rect 1519 214 1523 218
rect 1527 214 1531 218
rect 1575 214 1579 218
rect 1583 214 1587 218
rect 1623 214 1627 218
rect 1663 214 1667 218
rect 1471 174 1475 178
rect 1495 174 1499 178
rect 1527 174 1531 178
rect 1567 174 1571 178
rect 1583 174 1587 178
rect 1623 174 1627 178
rect 1207 118 1211 122
rect 1223 118 1227 122
rect 1263 118 1267 122
rect 1279 118 1283 122
rect 1295 118 1299 122
rect 1335 118 1339 122
rect 1351 118 1355 122
rect 1375 118 1379 122
rect 1415 118 1419 122
rect 1423 118 1427 122
rect 1455 118 1459 122
rect 1495 118 1499 122
rect 1503 118 1507 122
rect 1551 118 1555 122
rect 1567 118 1571 122
rect 1663 174 1667 178
rect 1591 118 1595 122
rect 1623 118 1627 122
rect 1663 118 1667 122
rect 111 78 115 82
rect 135 78 139 82
rect 167 78 171 82
rect 199 78 203 82
rect 231 78 235 82
rect 263 78 267 82
rect 295 78 299 82
rect 327 78 331 82
rect 359 78 363 82
rect 391 78 395 82
rect 423 78 427 82
rect 463 78 467 82
rect 503 78 507 82
rect 543 78 547 82
rect 575 78 579 82
rect 607 78 611 82
rect 639 78 643 82
rect 671 78 675 82
rect 703 78 707 82
rect 735 78 739 82
rect 767 78 771 82
rect 799 78 803 82
rect 831 78 835 82
rect 863 78 867 82
rect 895 78 899 82
rect 935 78 939 82
rect 975 78 979 82
rect 1015 78 1019 82
rect 1063 78 1067 82
rect 1103 78 1107 82
rect 1143 78 1147 82
rect 1183 78 1187 82
rect 1223 78 1227 82
rect 1263 78 1267 82
rect 1295 78 1299 82
rect 1335 78 1339 82
rect 1375 78 1379 82
rect 1415 78 1419 82
rect 1455 78 1459 82
rect 1503 78 1507 82
rect 1551 78 1555 82
rect 1591 78 1595 82
rect 1623 78 1627 82
rect 1663 78 1667 82
<< m4 >>
rect 96 1713 97 1719
rect 103 1718 1699 1719
rect 103 1714 111 1718
rect 115 1714 255 1718
rect 259 1714 287 1718
rect 291 1714 319 1718
rect 323 1714 359 1718
rect 363 1714 407 1718
rect 411 1714 455 1718
rect 459 1714 503 1718
rect 507 1714 551 1718
rect 555 1714 607 1718
rect 611 1714 663 1718
rect 667 1714 727 1718
rect 731 1714 783 1718
rect 787 1714 839 1718
rect 843 1714 895 1718
rect 899 1714 951 1718
rect 955 1714 1007 1718
rect 1011 1714 1063 1718
rect 1067 1714 1119 1718
rect 1123 1714 1175 1718
rect 1179 1714 1231 1718
rect 1235 1714 1287 1718
rect 1291 1714 1335 1718
rect 1339 1714 1375 1718
rect 1379 1714 1423 1718
rect 1427 1714 1471 1718
rect 1475 1714 1519 1718
rect 1523 1714 1663 1718
rect 1667 1714 1699 1718
rect 103 1713 1699 1714
rect 1705 1713 1706 1719
rect 84 1673 85 1679
rect 91 1678 1687 1679
rect 91 1674 111 1678
rect 115 1674 135 1678
rect 139 1674 167 1678
rect 171 1674 215 1678
rect 219 1674 255 1678
rect 259 1674 279 1678
rect 283 1674 287 1678
rect 291 1674 319 1678
rect 323 1674 343 1678
rect 347 1674 359 1678
rect 363 1674 407 1678
rect 411 1674 415 1678
rect 419 1674 455 1678
rect 459 1674 487 1678
rect 491 1674 503 1678
rect 507 1674 551 1678
rect 555 1674 559 1678
rect 563 1674 607 1678
rect 611 1674 631 1678
rect 635 1674 663 1678
rect 667 1674 711 1678
rect 715 1674 727 1678
rect 731 1674 783 1678
rect 787 1674 791 1678
rect 795 1674 839 1678
rect 843 1674 871 1678
rect 875 1674 895 1678
rect 899 1674 951 1678
rect 955 1674 1007 1678
rect 1011 1674 1031 1678
rect 1035 1674 1063 1678
rect 1067 1674 1103 1678
rect 1107 1674 1119 1678
rect 1123 1674 1175 1678
rect 1179 1674 1231 1678
rect 1235 1674 1247 1678
rect 1251 1674 1287 1678
rect 1291 1674 1319 1678
rect 1323 1674 1335 1678
rect 1339 1674 1375 1678
rect 1379 1674 1391 1678
rect 1395 1674 1423 1678
rect 1427 1674 1455 1678
rect 1459 1674 1471 1678
rect 1475 1674 1519 1678
rect 1523 1674 1583 1678
rect 1587 1674 1623 1678
rect 1627 1674 1663 1678
rect 1667 1674 1687 1678
rect 91 1673 1687 1674
rect 1693 1673 1694 1679
rect 96 1633 97 1639
rect 103 1638 1699 1639
rect 103 1634 111 1638
rect 115 1634 135 1638
rect 139 1634 167 1638
rect 171 1634 183 1638
rect 187 1634 215 1638
rect 219 1634 247 1638
rect 251 1634 279 1638
rect 283 1634 303 1638
rect 307 1634 343 1638
rect 347 1634 359 1638
rect 363 1634 415 1638
rect 419 1634 471 1638
rect 475 1634 487 1638
rect 491 1634 535 1638
rect 539 1634 559 1638
rect 563 1634 599 1638
rect 603 1634 631 1638
rect 635 1634 663 1638
rect 667 1634 711 1638
rect 715 1634 727 1638
rect 731 1634 791 1638
rect 795 1634 799 1638
rect 803 1634 871 1638
rect 875 1634 943 1638
rect 947 1634 951 1638
rect 955 1634 1023 1638
rect 1027 1634 1031 1638
rect 1035 1634 1103 1638
rect 1107 1634 1175 1638
rect 1179 1634 1247 1638
rect 1251 1634 1319 1638
rect 1323 1634 1391 1638
rect 1395 1634 1399 1638
rect 1403 1634 1455 1638
rect 1459 1634 1479 1638
rect 1483 1634 1519 1638
rect 1523 1634 1559 1638
rect 1563 1634 1583 1638
rect 1587 1634 1623 1638
rect 1627 1634 1663 1638
rect 1667 1634 1699 1638
rect 103 1633 1699 1634
rect 1705 1633 1706 1639
rect 84 1593 85 1599
rect 91 1598 1687 1599
rect 91 1594 111 1598
rect 115 1594 135 1598
rect 139 1594 167 1598
rect 171 1594 183 1598
rect 187 1594 223 1598
rect 227 1594 247 1598
rect 251 1594 279 1598
rect 283 1594 303 1598
rect 307 1594 335 1598
rect 339 1594 359 1598
rect 363 1594 383 1598
rect 387 1594 415 1598
rect 419 1594 431 1598
rect 435 1594 471 1598
rect 475 1594 479 1598
rect 483 1594 535 1598
rect 539 1594 599 1598
rect 603 1594 663 1598
rect 667 1594 727 1598
rect 731 1594 799 1598
rect 803 1594 871 1598
rect 875 1594 943 1598
rect 947 1594 951 1598
rect 955 1594 1023 1598
rect 1027 1594 1039 1598
rect 1043 1594 1103 1598
rect 1107 1594 1119 1598
rect 1123 1594 1175 1598
rect 1179 1594 1199 1598
rect 1203 1594 1247 1598
rect 1251 1594 1279 1598
rect 1283 1594 1319 1598
rect 1323 1594 1351 1598
rect 1355 1594 1399 1598
rect 1403 1594 1415 1598
rect 1419 1594 1471 1598
rect 1475 1594 1479 1598
rect 1483 1594 1527 1598
rect 1531 1594 1559 1598
rect 1563 1594 1583 1598
rect 1587 1594 1623 1598
rect 1627 1594 1663 1598
rect 1667 1594 1687 1598
rect 91 1593 1687 1594
rect 1693 1593 1694 1599
rect 96 1553 97 1559
rect 103 1558 1699 1559
rect 103 1554 111 1558
rect 115 1554 135 1558
rect 139 1554 167 1558
rect 171 1554 215 1558
rect 219 1554 223 1558
rect 227 1554 263 1558
rect 267 1554 279 1558
rect 283 1554 311 1558
rect 315 1554 335 1558
rect 339 1554 359 1558
rect 363 1554 383 1558
rect 387 1554 407 1558
rect 411 1554 431 1558
rect 435 1554 455 1558
rect 459 1554 479 1558
rect 483 1554 511 1558
rect 515 1554 535 1558
rect 539 1554 567 1558
rect 571 1554 599 1558
rect 603 1554 631 1558
rect 635 1554 663 1558
rect 667 1554 695 1558
rect 699 1554 727 1558
rect 731 1554 759 1558
rect 763 1554 799 1558
rect 803 1554 831 1558
rect 835 1554 871 1558
rect 875 1554 919 1558
rect 923 1554 951 1558
rect 955 1554 1007 1558
rect 1011 1554 1039 1558
rect 1043 1554 1095 1558
rect 1099 1554 1119 1558
rect 1123 1554 1183 1558
rect 1187 1554 1199 1558
rect 1203 1554 1263 1558
rect 1267 1554 1279 1558
rect 1283 1554 1335 1558
rect 1339 1554 1351 1558
rect 1355 1554 1407 1558
rect 1411 1554 1415 1558
rect 1419 1554 1471 1558
rect 1475 1554 1527 1558
rect 1531 1554 1583 1558
rect 1587 1554 1623 1558
rect 1627 1554 1663 1558
rect 1667 1554 1699 1558
rect 103 1553 1699 1554
rect 1705 1553 1706 1559
rect 84 1509 85 1515
rect 91 1514 1687 1515
rect 91 1510 111 1514
rect 115 1510 135 1514
rect 139 1510 167 1514
rect 171 1510 215 1514
rect 219 1510 223 1514
rect 227 1510 263 1514
rect 267 1510 295 1514
rect 299 1510 311 1514
rect 315 1510 359 1514
rect 363 1510 375 1514
rect 379 1510 407 1514
rect 411 1510 455 1514
rect 459 1510 511 1514
rect 515 1510 527 1514
rect 531 1510 567 1514
rect 571 1510 599 1514
rect 603 1510 631 1514
rect 635 1510 671 1514
rect 675 1510 695 1514
rect 699 1510 743 1514
rect 747 1510 759 1514
rect 763 1510 815 1514
rect 819 1510 831 1514
rect 835 1510 879 1514
rect 883 1510 919 1514
rect 923 1510 943 1514
rect 947 1510 1007 1514
rect 1011 1510 1063 1514
rect 1067 1510 1095 1514
rect 1099 1510 1111 1514
rect 1115 1510 1151 1514
rect 1155 1510 1183 1514
rect 1187 1510 1215 1514
rect 1219 1510 1255 1514
rect 1259 1510 1263 1514
rect 1267 1510 1295 1514
rect 1299 1510 1335 1514
rect 1339 1510 1351 1514
rect 1355 1510 1407 1514
rect 1411 1510 1415 1514
rect 1419 1510 1471 1514
rect 1475 1510 1487 1514
rect 1491 1510 1527 1514
rect 1531 1510 1567 1514
rect 1571 1510 1583 1514
rect 1587 1510 1623 1514
rect 1627 1510 1663 1514
rect 1667 1510 1687 1514
rect 91 1509 1687 1510
rect 1693 1509 1694 1515
rect 96 1469 97 1475
rect 103 1474 1699 1475
rect 103 1470 111 1474
rect 115 1470 135 1474
rect 139 1470 167 1474
rect 171 1470 223 1474
rect 227 1470 295 1474
rect 299 1470 375 1474
rect 379 1470 455 1474
rect 459 1470 527 1474
rect 531 1470 599 1474
rect 603 1470 663 1474
rect 667 1470 671 1474
rect 675 1470 719 1474
rect 723 1470 743 1474
rect 747 1470 783 1474
rect 787 1470 815 1474
rect 819 1470 847 1474
rect 851 1470 879 1474
rect 883 1470 903 1474
rect 907 1470 943 1474
rect 947 1470 959 1474
rect 963 1470 1007 1474
rect 1011 1470 1015 1474
rect 1019 1470 1063 1474
rect 1067 1470 1071 1474
rect 1075 1470 1111 1474
rect 1115 1470 1119 1474
rect 1123 1470 1151 1474
rect 1155 1470 1159 1474
rect 1163 1470 1183 1474
rect 1187 1470 1207 1474
rect 1211 1470 1215 1474
rect 1219 1470 1255 1474
rect 1259 1470 1263 1474
rect 1267 1470 1295 1474
rect 1299 1470 1327 1474
rect 1331 1470 1351 1474
rect 1355 1470 1399 1474
rect 1403 1470 1415 1474
rect 1419 1470 1479 1474
rect 1483 1470 1487 1474
rect 1491 1470 1559 1474
rect 1563 1470 1567 1474
rect 1571 1470 1623 1474
rect 1627 1470 1663 1474
rect 1667 1470 1699 1474
rect 103 1469 1699 1470
rect 1705 1469 1706 1475
rect 84 1425 85 1431
rect 91 1430 1687 1431
rect 91 1426 111 1430
rect 115 1426 135 1430
rect 139 1426 167 1430
rect 171 1426 215 1430
rect 219 1426 223 1430
rect 227 1426 287 1430
rect 291 1426 295 1430
rect 299 1426 359 1430
rect 363 1426 375 1430
rect 379 1426 439 1430
rect 443 1426 455 1430
rect 459 1426 519 1430
rect 523 1426 527 1430
rect 531 1426 599 1430
rect 603 1426 663 1430
rect 667 1426 679 1430
rect 683 1426 719 1430
rect 723 1426 759 1430
rect 763 1426 783 1430
rect 787 1426 831 1430
rect 835 1426 847 1430
rect 851 1426 903 1430
rect 907 1426 959 1430
rect 963 1426 967 1430
rect 971 1426 1015 1430
rect 1019 1426 1031 1430
rect 1035 1426 1071 1430
rect 1075 1426 1103 1430
rect 1107 1426 1119 1430
rect 1123 1426 1159 1430
rect 1163 1426 1167 1430
rect 1171 1426 1207 1430
rect 1211 1426 1231 1430
rect 1235 1426 1263 1430
rect 1267 1426 1295 1430
rect 1299 1426 1327 1430
rect 1331 1426 1359 1430
rect 1363 1426 1399 1430
rect 1403 1426 1415 1430
rect 1419 1426 1463 1430
rect 1467 1426 1479 1430
rect 1483 1426 1503 1430
rect 1507 1426 1551 1430
rect 1555 1426 1559 1430
rect 1563 1426 1591 1430
rect 1595 1426 1623 1430
rect 1627 1426 1663 1430
rect 1667 1426 1687 1430
rect 91 1425 1687 1426
rect 1693 1425 1694 1431
rect 96 1385 97 1391
rect 103 1390 1699 1391
rect 103 1386 111 1390
rect 115 1386 135 1390
rect 139 1386 167 1390
rect 171 1386 215 1390
rect 219 1386 223 1390
rect 227 1386 287 1390
rect 291 1386 359 1390
rect 363 1386 431 1390
rect 435 1386 439 1390
rect 443 1386 503 1390
rect 507 1386 519 1390
rect 523 1386 583 1390
rect 587 1386 599 1390
rect 603 1386 663 1390
rect 667 1386 679 1390
rect 683 1386 743 1390
rect 747 1386 759 1390
rect 763 1386 815 1390
rect 819 1386 831 1390
rect 835 1386 887 1390
rect 891 1386 903 1390
rect 907 1386 959 1390
rect 963 1386 967 1390
rect 971 1386 1031 1390
rect 1035 1386 1103 1390
rect 1107 1386 1167 1390
rect 1171 1386 1175 1390
rect 1179 1386 1231 1390
rect 1235 1386 1239 1390
rect 1243 1386 1295 1390
rect 1299 1386 1303 1390
rect 1307 1386 1359 1390
rect 1363 1386 1367 1390
rect 1371 1386 1415 1390
rect 1419 1386 1431 1390
rect 1435 1386 1463 1390
rect 1467 1386 1495 1390
rect 1499 1386 1503 1390
rect 1507 1386 1551 1390
rect 1555 1386 1567 1390
rect 1571 1386 1591 1390
rect 1595 1386 1623 1390
rect 1627 1386 1663 1390
rect 1667 1386 1699 1390
rect 103 1385 1699 1386
rect 1705 1385 1706 1391
rect 84 1345 85 1351
rect 91 1350 1687 1351
rect 91 1346 111 1350
rect 115 1346 135 1350
rect 139 1346 167 1350
rect 171 1346 183 1350
rect 187 1346 223 1350
rect 227 1346 239 1350
rect 243 1346 287 1350
rect 291 1346 295 1350
rect 299 1346 351 1350
rect 355 1346 359 1350
rect 363 1346 399 1350
rect 403 1346 431 1350
rect 435 1346 455 1350
rect 459 1346 503 1350
rect 507 1346 511 1350
rect 515 1346 567 1350
rect 571 1346 583 1350
rect 587 1346 631 1350
rect 635 1346 663 1350
rect 667 1346 695 1350
rect 699 1346 743 1350
rect 747 1346 759 1350
rect 763 1346 815 1350
rect 819 1346 823 1350
rect 827 1346 887 1350
rect 891 1346 959 1350
rect 963 1346 1023 1350
rect 1027 1346 1031 1350
rect 1035 1346 1087 1350
rect 1091 1346 1103 1350
rect 1107 1346 1151 1350
rect 1155 1346 1175 1350
rect 1179 1346 1215 1350
rect 1219 1346 1239 1350
rect 1243 1346 1279 1350
rect 1283 1346 1303 1350
rect 1307 1346 1343 1350
rect 1347 1346 1367 1350
rect 1371 1346 1407 1350
rect 1411 1346 1431 1350
rect 1435 1346 1479 1350
rect 1483 1346 1495 1350
rect 1499 1346 1559 1350
rect 1563 1346 1567 1350
rect 1571 1346 1623 1350
rect 1627 1346 1663 1350
rect 1667 1346 1687 1350
rect 91 1345 1687 1346
rect 1693 1345 1694 1351
rect 96 1301 97 1307
rect 103 1306 1699 1307
rect 103 1302 111 1306
rect 115 1302 135 1306
rect 139 1302 183 1306
rect 187 1302 231 1306
rect 235 1302 239 1306
rect 243 1302 279 1306
rect 283 1302 295 1306
rect 299 1302 327 1306
rect 331 1302 351 1306
rect 355 1302 375 1306
rect 379 1302 399 1306
rect 403 1302 431 1306
rect 435 1302 455 1306
rect 459 1302 487 1306
rect 491 1302 511 1306
rect 515 1302 543 1306
rect 547 1302 567 1306
rect 571 1302 607 1306
rect 611 1302 631 1306
rect 635 1302 663 1306
rect 667 1302 695 1306
rect 699 1302 719 1306
rect 723 1302 759 1306
rect 763 1302 775 1306
rect 779 1302 823 1306
rect 827 1302 831 1306
rect 835 1302 887 1306
rect 891 1302 895 1306
rect 899 1302 959 1306
rect 963 1302 1023 1306
rect 1027 1302 1079 1306
rect 1083 1302 1087 1306
rect 1091 1302 1143 1306
rect 1147 1302 1151 1306
rect 1155 1302 1207 1306
rect 1211 1302 1215 1306
rect 1219 1302 1279 1306
rect 1283 1302 1343 1306
rect 1347 1302 1359 1306
rect 1363 1302 1407 1306
rect 1411 1302 1447 1306
rect 1451 1302 1479 1306
rect 1483 1302 1543 1306
rect 1547 1302 1559 1306
rect 1563 1302 1623 1306
rect 1627 1302 1663 1306
rect 1667 1302 1699 1306
rect 103 1301 1699 1302
rect 1705 1301 1706 1307
rect 84 1261 85 1267
rect 91 1266 1687 1267
rect 91 1262 111 1266
rect 115 1262 135 1266
rect 139 1262 167 1266
rect 171 1262 183 1266
rect 187 1262 223 1266
rect 227 1262 231 1266
rect 235 1262 279 1266
rect 283 1262 327 1266
rect 331 1262 375 1266
rect 379 1262 383 1266
rect 387 1262 431 1266
rect 435 1262 439 1266
rect 443 1262 487 1266
rect 491 1262 495 1266
rect 499 1262 543 1266
rect 547 1262 551 1266
rect 555 1262 607 1266
rect 611 1262 663 1266
rect 667 1262 719 1266
rect 723 1262 767 1266
rect 771 1262 775 1266
rect 779 1262 815 1266
rect 819 1262 831 1266
rect 835 1262 871 1266
rect 875 1262 895 1266
rect 899 1262 927 1266
rect 931 1262 959 1266
rect 963 1262 983 1266
rect 987 1262 1023 1266
rect 1027 1262 1039 1266
rect 1043 1262 1079 1266
rect 1083 1262 1095 1266
rect 1099 1262 1143 1266
rect 1147 1262 1159 1266
rect 1163 1262 1207 1266
rect 1211 1262 1231 1266
rect 1235 1262 1279 1266
rect 1283 1262 1319 1266
rect 1323 1262 1359 1266
rect 1363 1262 1423 1266
rect 1427 1262 1447 1266
rect 1451 1262 1535 1266
rect 1539 1262 1543 1266
rect 1547 1262 1623 1266
rect 1627 1262 1663 1266
rect 1667 1262 1687 1266
rect 91 1261 1687 1262
rect 1693 1261 1694 1267
rect 96 1217 97 1223
rect 103 1222 1699 1223
rect 103 1218 111 1222
rect 115 1218 135 1222
rect 139 1218 167 1222
rect 171 1218 223 1222
rect 227 1218 279 1222
rect 283 1218 327 1222
rect 331 1218 335 1222
rect 339 1218 383 1222
rect 387 1218 431 1222
rect 435 1218 439 1222
rect 443 1218 487 1222
rect 491 1218 495 1222
rect 499 1218 543 1222
rect 547 1218 551 1222
rect 555 1218 599 1222
rect 603 1218 607 1222
rect 611 1218 655 1222
rect 659 1218 663 1222
rect 667 1218 711 1222
rect 715 1218 719 1222
rect 723 1218 767 1222
rect 771 1218 815 1222
rect 819 1218 823 1222
rect 827 1218 871 1222
rect 875 1218 887 1222
rect 891 1218 927 1222
rect 931 1218 951 1222
rect 955 1218 983 1222
rect 987 1218 1015 1222
rect 1019 1218 1039 1222
rect 1043 1218 1079 1222
rect 1083 1218 1095 1222
rect 1099 1218 1143 1222
rect 1147 1218 1159 1222
rect 1163 1218 1207 1222
rect 1211 1218 1231 1222
rect 1235 1218 1279 1222
rect 1283 1218 1319 1222
rect 1323 1218 1359 1222
rect 1363 1218 1423 1222
rect 1427 1218 1447 1222
rect 1451 1218 1535 1222
rect 1539 1218 1543 1222
rect 1547 1218 1623 1222
rect 1627 1218 1663 1222
rect 1667 1218 1699 1222
rect 103 1217 1699 1218
rect 1705 1217 1706 1223
rect 84 1173 85 1179
rect 91 1178 1687 1179
rect 91 1174 111 1178
rect 115 1174 135 1178
rect 139 1174 167 1178
rect 171 1174 223 1178
rect 227 1174 279 1178
rect 283 1174 287 1178
rect 291 1174 335 1178
rect 339 1174 351 1178
rect 355 1174 383 1178
rect 387 1174 415 1178
rect 419 1174 431 1178
rect 435 1174 471 1178
rect 475 1174 487 1178
rect 491 1174 535 1178
rect 539 1174 543 1178
rect 547 1174 599 1178
rect 603 1174 655 1178
rect 659 1174 663 1178
rect 667 1174 711 1178
rect 715 1174 727 1178
rect 731 1174 767 1178
rect 771 1174 783 1178
rect 787 1174 823 1178
rect 827 1174 839 1178
rect 843 1174 887 1178
rect 891 1174 903 1178
rect 907 1174 951 1178
rect 955 1174 967 1178
rect 971 1174 1015 1178
rect 1019 1174 1031 1178
rect 1035 1174 1079 1178
rect 1083 1174 1095 1178
rect 1099 1174 1143 1178
rect 1147 1174 1159 1178
rect 1163 1174 1207 1178
rect 1211 1174 1215 1178
rect 1219 1174 1279 1178
rect 1283 1174 1343 1178
rect 1347 1174 1359 1178
rect 1363 1174 1407 1178
rect 1411 1174 1447 1178
rect 1451 1174 1479 1178
rect 1483 1174 1543 1178
rect 1547 1174 1559 1178
rect 1563 1174 1623 1178
rect 1627 1174 1663 1178
rect 1667 1174 1687 1178
rect 91 1173 1687 1174
rect 1693 1173 1694 1179
rect 96 1129 97 1135
rect 103 1134 1699 1135
rect 103 1130 111 1134
rect 115 1130 135 1134
rect 139 1130 143 1134
rect 147 1130 167 1134
rect 171 1130 175 1134
rect 179 1130 215 1134
rect 219 1130 223 1134
rect 227 1130 271 1134
rect 275 1130 287 1134
rect 291 1130 335 1134
rect 339 1130 351 1134
rect 355 1130 399 1134
rect 403 1130 415 1134
rect 419 1130 463 1134
rect 467 1130 471 1134
rect 475 1130 527 1134
rect 531 1130 535 1134
rect 539 1130 599 1134
rect 603 1130 663 1134
rect 667 1130 727 1134
rect 731 1130 783 1134
rect 787 1130 791 1134
rect 795 1130 839 1134
rect 843 1130 855 1134
rect 859 1130 903 1134
rect 907 1130 911 1134
rect 915 1130 967 1134
rect 971 1130 1023 1134
rect 1027 1130 1031 1134
rect 1035 1130 1087 1134
rect 1091 1130 1095 1134
rect 1099 1130 1151 1134
rect 1155 1130 1159 1134
rect 1163 1130 1215 1134
rect 1219 1130 1279 1134
rect 1283 1130 1335 1134
rect 1339 1130 1343 1134
rect 1347 1130 1391 1134
rect 1395 1130 1407 1134
rect 1411 1130 1447 1134
rect 1451 1130 1479 1134
rect 1483 1130 1495 1134
rect 1499 1130 1543 1134
rect 1547 1130 1559 1134
rect 1563 1130 1591 1134
rect 1595 1130 1623 1134
rect 1627 1130 1663 1134
rect 1667 1130 1699 1134
rect 103 1129 1699 1130
rect 1705 1129 1706 1135
rect 84 1085 85 1091
rect 91 1090 1687 1091
rect 91 1086 111 1090
rect 115 1086 143 1090
rect 147 1086 175 1090
rect 179 1086 215 1090
rect 219 1086 247 1090
rect 251 1086 271 1090
rect 275 1086 279 1090
rect 283 1086 311 1090
rect 315 1086 335 1090
rect 339 1086 351 1090
rect 355 1086 391 1090
rect 395 1086 399 1090
rect 403 1086 439 1090
rect 443 1086 463 1090
rect 467 1086 503 1090
rect 507 1086 527 1090
rect 531 1086 575 1090
rect 579 1086 599 1090
rect 603 1086 655 1090
rect 659 1086 663 1090
rect 667 1086 727 1090
rect 731 1086 735 1090
rect 739 1086 791 1090
rect 795 1086 815 1090
rect 819 1086 855 1090
rect 859 1086 895 1090
rect 899 1086 911 1090
rect 915 1086 967 1090
rect 971 1086 1023 1090
rect 1027 1086 1039 1090
rect 1043 1086 1087 1090
rect 1091 1086 1111 1090
rect 1115 1086 1151 1090
rect 1155 1086 1175 1090
rect 1179 1086 1215 1090
rect 1219 1086 1239 1090
rect 1243 1086 1279 1090
rect 1283 1086 1303 1090
rect 1307 1086 1335 1090
rect 1339 1086 1359 1090
rect 1363 1086 1391 1090
rect 1395 1086 1415 1090
rect 1419 1086 1447 1090
rect 1451 1086 1463 1090
rect 1467 1086 1495 1090
rect 1499 1086 1503 1090
rect 1507 1086 1543 1090
rect 1547 1086 1551 1090
rect 1555 1086 1591 1090
rect 1595 1086 1623 1090
rect 1627 1086 1663 1090
rect 1667 1086 1687 1090
rect 91 1085 1687 1086
rect 1693 1085 1694 1091
rect 96 1041 97 1047
rect 103 1046 1699 1047
rect 103 1042 111 1046
rect 115 1042 215 1046
rect 219 1042 247 1046
rect 251 1042 279 1046
rect 283 1042 295 1046
rect 299 1042 311 1046
rect 315 1042 327 1046
rect 331 1042 351 1046
rect 355 1042 359 1046
rect 363 1042 391 1046
rect 395 1042 423 1046
rect 427 1042 439 1046
rect 443 1042 455 1046
rect 459 1042 503 1046
rect 507 1042 559 1046
rect 563 1042 575 1046
rect 579 1042 631 1046
rect 635 1042 655 1046
rect 659 1042 711 1046
rect 715 1042 735 1046
rect 739 1042 799 1046
rect 803 1042 815 1046
rect 819 1042 879 1046
rect 883 1042 895 1046
rect 899 1042 959 1046
rect 963 1042 967 1046
rect 971 1042 1031 1046
rect 1035 1042 1039 1046
rect 1043 1042 1095 1046
rect 1099 1042 1111 1046
rect 1115 1042 1159 1046
rect 1163 1042 1175 1046
rect 1179 1042 1223 1046
rect 1227 1042 1239 1046
rect 1243 1042 1279 1046
rect 1283 1042 1303 1046
rect 1307 1042 1335 1046
rect 1339 1042 1359 1046
rect 1363 1042 1383 1046
rect 1387 1042 1415 1046
rect 1419 1042 1431 1046
rect 1435 1042 1463 1046
rect 1467 1042 1479 1046
rect 1483 1042 1503 1046
rect 1507 1042 1535 1046
rect 1539 1042 1551 1046
rect 1555 1042 1591 1046
rect 1595 1042 1623 1046
rect 1627 1042 1663 1046
rect 1667 1042 1699 1046
rect 103 1041 1699 1042
rect 1705 1041 1706 1047
rect 84 1001 85 1007
rect 91 1006 1687 1007
rect 91 1002 111 1006
rect 115 1002 247 1006
rect 251 1002 279 1006
rect 283 1002 295 1006
rect 299 1002 311 1006
rect 315 1002 327 1006
rect 331 1002 343 1006
rect 347 1002 359 1006
rect 363 1002 383 1006
rect 387 1002 391 1006
rect 395 1002 423 1006
rect 427 1002 455 1006
rect 459 1002 479 1006
rect 483 1002 503 1006
rect 507 1002 543 1006
rect 547 1002 559 1006
rect 563 1002 615 1006
rect 619 1002 631 1006
rect 635 1002 687 1006
rect 691 1002 711 1006
rect 715 1002 759 1006
rect 763 1002 799 1006
rect 803 1002 831 1006
rect 835 1002 879 1006
rect 883 1002 903 1006
rect 907 1002 959 1006
rect 963 1002 967 1006
rect 971 1002 1031 1006
rect 1035 1002 1095 1006
rect 1099 1002 1159 1006
rect 1163 1002 1223 1006
rect 1227 1002 1279 1006
rect 1283 1002 1287 1006
rect 1291 1002 1335 1006
rect 1339 1002 1343 1006
rect 1347 1002 1383 1006
rect 1387 1002 1399 1006
rect 1403 1002 1431 1006
rect 1435 1002 1447 1006
rect 1451 1002 1479 1006
rect 1483 1002 1495 1006
rect 1499 1002 1535 1006
rect 1539 1002 1543 1006
rect 1547 1002 1591 1006
rect 1595 1002 1623 1006
rect 1627 1002 1663 1006
rect 1667 1002 1687 1006
rect 91 1001 1687 1002
rect 1693 1001 1694 1007
rect 96 961 97 967
rect 103 966 1699 967
rect 103 962 111 966
rect 115 962 167 966
rect 171 962 199 966
rect 203 962 239 966
rect 243 962 247 966
rect 251 962 279 966
rect 283 962 287 966
rect 291 962 311 966
rect 315 962 343 966
rect 347 962 383 966
rect 387 962 407 966
rect 411 962 423 966
rect 427 962 471 966
rect 475 962 479 966
rect 483 962 535 966
rect 539 962 543 966
rect 547 962 599 966
rect 603 962 615 966
rect 619 962 663 966
rect 667 962 687 966
rect 691 962 727 966
rect 731 962 759 966
rect 763 962 791 966
rect 795 962 831 966
rect 835 962 847 966
rect 851 962 903 966
rect 907 962 911 966
rect 915 962 967 966
rect 971 962 975 966
rect 979 962 1031 966
rect 1035 962 1039 966
rect 1043 962 1095 966
rect 1099 962 1103 966
rect 1107 962 1159 966
rect 1163 962 1167 966
rect 1171 962 1223 966
rect 1227 962 1231 966
rect 1235 962 1287 966
rect 1291 962 1343 966
rect 1347 962 1391 966
rect 1395 962 1399 966
rect 1403 962 1431 966
rect 1435 962 1447 966
rect 1451 962 1471 966
rect 1475 962 1495 966
rect 1499 962 1511 966
rect 1515 962 1543 966
rect 1547 962 1551 966
rect 1555 962 1591 966
rect 1595 962 1623 966
rect 1627 962 1663 966
rect 1667 962 1699 966
rect 103 961 1699 962
rect 1705 961 1706 967
rect 84 917 85 923
rect 91 922 1687 923
rect 91 918 111 922
rect 115 918 135 922
rect 139 918 167 922
rect 171 918 199 922
rect 203 918 207 922
rect 211 918 239 922
rect 243 918 271 922
rect 275 918 287 922
rect 291 918 335 922
rect 339 918 343 922
rect 347 918 407 922
rect 411 918 471 922
rect 475 918 535 922
rect 539 918 591 922
rect 595 918 599 922
rect 603 918 647 922
rect 651 918 663 922
rect 667 918 703 922
rect 707 918 727 922
rect 731 918 751 922
rect 755 918 791 922
rect 795 918 799 922
rect 803 918 847 922
rect 851 918 903 922
rect 907 918 911 922
rect 915 918 959 922
rect 963 918 975 922
rect 979 918 1023 922
rect 1027 918 1039 922
rect 1043 918 1087 922
rect 1091 918 1103 922
rect 1107 918 1143 922
rect 1147 918 1167 922
rect 1171 918 1199 922
rect 1203 918 1231 922
rect 1235 918 1255 922
rect 1259 918 1287 922
rect 1291 918 1319 922
rect 1323 918 1343 922
rect 1347 918 1383 922
rect 1387 918 1391 922
rect 1395 918 1431 922
rect 1435 918 1471 922
rect 1475 918 1511 922
rect 1515 918 1551 922
rect 1555 918 1591 922
rect 1595 918 1623 922
rect 1627 918 1663 922
rect 1667 918 1687 922
rect 91 917 1687 918
rect 1693 917 1694 923
rect 96 873 97 879
rect 103 878 1699 879
rect 103 874 111 878
rect 115 874 135 878
rect 139 874 167 878
rect 171 874 207 878
rect 211 874 271 878
rect 275 874 335 878
rect 339 874 407 878
rect 411 874 471 878
rect 475 874 535 878
rect 539 874 591 878
rect 595 874 599 878
rect 603 874 647 878
rect 651 874 655 878
rect 659 874 703 878
rect 707 874 751 878
rect 755 874 799 878
rect 803 874 847 878
rect 851 874 903 878
rect 907 874 959 878
rect 963 874 967 878
rect 971 874 1023 878
rect 1027 874 1039 878
rect 1043 874 1087 878
rect 1091 874 1103 878
rect 1107 874 1143 878
rect 1147 874 1167 878
rect 1171 874 1199 878
rect 1203 874 1231 878
rect 1235 874 1255 878
rect 1259 874 1287 878
rect 1291 874 1319 878
rect 1323 874 1343 878
rect 1347 874 1383 878
rect 1387 874 1399 878
rect 1403 874 1463 878
rect 1467 874 1663 878
rect 1667 874 1699 878
rect 103 873 1699 874
rect 1705 873 1706 879
rect 84 833 85 839
rect 91 838 1687 839
rect 91 834 111 838
rect 115 834 135 838
rect 139 834 167 838
rect 171 834 207 838
rect 211 834 215 838
rect 219 834 271 838
rect 275 834 279 838
rect 283 834 335 838
rect 339 834 343 838
rect 347 834 407 838
rect 411 834 415 838
rect 419 834 471 838
rect 475 834 479 838
rect 483 834 535 838
rect 539 834 543 838
rect 547 834 599 838
rect 603 834 607 838
rect 611 834 655 838
rect 659 834 671 838
rect 675 834 703 838
rect 707 834 735 838
rect 739 834 751 838
rect 755 834 791 838
rect 795 834 799 838
rect 803 834 847 838
rect 851 834 903 838
rect 907 834 911 838
rect 915 834 967 838
rect 971 834 975 838
rect 979 834 1039 838
rect 1043 834 1103 838
rect 1107 834 1111 838
rect 1115 834 1167 838
rect 1171 834 1183 838
rect 1187 834 1231 838
rect 1235 834 1247 838
rect 1251 834 1287 838
rect 1291 834 1311 838
rect 1315 834 1343 838
rect 1347 834 1367 838
rect 1371 834 1399 838
rect 1403 834 1423 838
rect 1427 834 1463 838
rect 1467 834 1479 838
rect 1483 834 1535 838
rect 1539 834 1591 838
rect 1595 834 1663 838
rect 1667 834 1687 838
rect 91 833 1687 834
rect 1693 833 1694 839
rect 96 789 97 795
rect 103 794 1699 795
rect 103 790 111 794
rect 115 790 135 794
rect 139 790 167 794
rect 171 790 175 794
rect 179 790 215 794
rect 219 790 231 794
rect 235 790 279 794
rect 283 790 295 794
rect 299 790 343 794
rect 347 790 367 794
rect 371 790 415 794
rect 419 790 447 794
rect 451 790 479 794
rect 483 790 527 794
rect 531 790 543 794
rect 547 790 607 794
rect 611 790 615 794
rect 619 790 671 794
rect 675 790 703 794
rect 707 790 735 794
rect 739 790 791 794
rect 795 790 847 794
rect 851 790 871 794
rect 875 790 911 794
rect 915 790 951 794
rect 955 790 975 794
rect 979 790 1023 794
rect 1027 790 1039 794
rect 1043 790 1095 794
rect 1099 790 1111 794
rect 1115 790 1167 794
rect 1171 790 1183 794
rect 1187 790 1231 794
rect 1235 790 1247 794
rect 1251 790 1295 794
rect 1299 790 1311 794
rect 1315 790 1359 794
rect 1363 790 1367 794
rect 1371 790 1415 794
rect 1419 790 1423 794
rect 1427 790 1471 794
rect 1475 790 1479 794
rect 1483 790 1527 794
rect 1531 790 1535 794
rect 1539 790 1591 794
rect 1595 790 1663 794
rect 1667 790 1699 794
rect 103 789 1699 790
rect 1705 789 1706 795
rect 84 749 85 755
rect 91 754 1687 755
rect 91 750 111 754
rect 115 750 135 754
rect 139 750 175 754
rect 179 750 215 754
rect 219 750 231 754
rect 235 750 247 754
rect 251 750 279 754
rect 283 750 295 754
rect 299 750 319 754
rect 323 750 359 754
rect 363 750 367 754
rect 371 750 399 754
rect 403 750 439 754
rect 443 750 447 754
rect 451 750 487 754
rect 491 750 527 754
rect 531 750 543 754
rect 547 750 607 754
rect 611 750 615 754
rect 619 750 671 754
rect 675 750 703 754
rect 707 750 735 754
rect 739 750 791 754
rect 795 750 799 754
rect 803 750 863 754
rect 867 750 871 754
rect 875 750 927 754
rect 931 750 951 754
rect 955 750 991 754
rect 995 750 1023 754
rect 1027 750 1055 754
rect 1059 750 1095 754
rect 1099 750 1119 754
rect 1123 750 1167 754
rect 1171 750 1183 754
rect 1187 750 1231 754
rect 1235 750 1239 754
rect 1243 750 1295 754
rect 1299 750 1351 754
rect 1355 750 1359 754
rect 1363 750 1407 754
rect 1411 750 1415 754
rect 1419 750 1463 754
rect 1467 750 1471 754
rect 1475 750 1519 754
rect 1523 750 1527 754
rect 1531 750 1583 754
rect 1587 750 1591 754
rect 1595 750 1623 754
rect 1627 750 1663 754
rect 1667 750 1687 754
rect 91 749 1687 750
rect 1693 749 1694 755
rect 96 705 97 711
rect 103 710 1699 711
rect 103 706 111 710
rect 115 706 215 710
rect 219 706 247 710
rect 251 706 279 710
rect 283 706 311 710
rect 315 706 319 710
rect 323 706 343 710
rect 347 706 359 710
rect 363 706 375 710
rect 379 706 399 710
rect 403 706 407 710
rect 411 706 439 710
rect 443 706 471 710
rect 475 706 487 710
rect 491 706 503 710
rect 507 706 543 710
rect 547 706 591 710
rect 595 706 607 710
rect 611 706 647 710
rect 651 706 671 710
rect 675 706 703 710
rect 707 706 735 710
rect 739 706 759 710
rect 763 706 799 710
rect 803 706 823 710
rect 827 706 863 710
rect 867 706 887 710
rect 891 706 927 710
rect 931 706 959 710
rect 963 706 991 710
rect 995 706 1023 710
rect 1027 706 1055 710
rect 1059 706 1087 710
rect 1091 706 1119 710
rect 1123 706 1159 710
rect 1163 706 1183 710
rect 1187 706 1223 710
rect 1227 706 1239 710
rect 1243 706 1287 710
rect 1291 706 1295 710
rect 1299 706 1351 710
rect 1355 706 1407 710
rect 1411 706 1415 710
rect 1419 706 1463 710
rect 1467 706 1471 710
rect 1475 706 1519 710
rect 1523 706 1527 710
rect 1531 706 1583 710
rect 1587 706 1623 710
rect 1627 706 1663 710
rect 1667 706 1699 710
rect 103 705 1699 706
rect 1705 705 1706 711
rect 84 665 85 671
rect 91 670 1687 671
rect 91 666 111 670
rect 115 666 279 670
rect 283 666 295 670
rect 299 666 311 670
rect 315 666 327 670
rect 331 666 343 670
rect 347 666 359 670
rect 363 666 375 670
rect 379 666 391 670
rect 395 666 407 670
rect 411 666 423 670
rect 427 666 439 670
rect 443 666 455 670
rect 459 666 471 670
rect 475 666 487 670
rect 491 666 503 670
rect 507 666 519 670
rect 523 666 543 670
rect 547 666 551 670
rect 555 666 591 670
rect 595 666 639 670
rect 643 666 647 670
rect 651 666 687 670
rect 691 666 703 670
rect 707 666 735 670
rect 739 666 759 670
rect 763 666 791 670
rect 795 666 823 670
rect 827 666 847 670
rect 851 666 887 670
rect 891 666 911 670
rect 915 666 959 670
rect 963 666 975 670
rect 979 666 1023 670
rect 1027 666 1047 670
rect 1051 666 1087 670
rect 1091 666 1127 670
rect 1131 666 1159 670
rect 1163 666 1215 670
rect 1219 666 1223 670
rect 1227 666 1287 670
rect 1291 666 1295 670
rect 1299 666 1351 670
rect 1355 666 1383 670
rect 1387 666 1415 670
rect 1419 666 1471 670
rect 1475 666 1527 670
rect 1531 666 1559 670
rect 1563 666 1583 670
rect 1587 666 1623 670
rect 1627 666 1663 670
rect 1667 666 1687 670
rect 91 665 1687 666
rect 1693 665 1694 671
rect 96 625 97 631
rect 103 630 1699 631
rect 103 626 111 630
rect 115 626 247 630
rect 251 626 279 630
rect 283 626 295 630
rect 299 626 319 630
rect 323 626 327 630
rect 331 626 359 630
rect 363 626 367 630
rect 371 626 391 630
rect 395 626 423 630
rect 427 626 455 630
rect 459 626 471 630
rect 475 626 487 630
rect 491 626 519 630
rect 523 626 551 630
rect 555 626 567 630
rect 571 626 591 630
rect 595 626 615 630
rect 619 626 639 630
rect 643 626 663 630
rect 667 626 687 630
rect 691 626 719 630
rect 723 626 735 630
rect 739 626 775 630
rect 779 626 791 630
rect 795 626 831 630
rect 835 626 847 630
rect 851 626 895 630
rect 899 626 911 630
rect 915 626 967 630
rect 971 626 975 630
rect 979 626 1047 630
rect 1051 626 1127 630
rect 1131 626 1207 630
rect 1211 626 1215 630
rect 1219 626 1287 630
rect 1291 626 1295 630
rect 1299 626 1359 630
rect 1363 626 1383 630
rect 1387 626 1431 630
rect 1435 626 1471 630
rect 1475 626 1503 630
rect 1507 626 1559 630
rect 1563 626 1575 630
rect 1579 626 1623 630
rect 1627 626 1663 630
rect 1667 626 1699 630
rect 103 625 1699 626
rect 1705 625 1706 631
rect 84 585 85 591
rect 91 590 1687 591
rect 91 586 111 590
rect 115 586 167 590
rect 171 586 215 590
rect 219 586 247 590
rect 251 586 271 590
rect 275 586 279 590
rect 283 586 319 590
rect 323 586 335 590
rect 339 586 367 590
rect 371 586 407 590
rect 411 586 423 590
rect 427 586 471 590
rect 475 586 487 590
rect 491 586 519 590
rect 523 586 559 590
rect 563 586 567 590
rect 571 586 615 590
rect 619 586 631 590
rect 635 586 663 590
rect 667 586 703 590
rect 707 586 719 590
rect 723 586 767 590
rect 771 586 775 590
rect 779 586 823 590
rect 827 586 831 590
rect 835 586 879 590
rect 883 586 895 590
rect 899 586 935 590
rect 939 586 967 590
rect 971 586 991 590
rect 995 586 1047 590
rect 1051 586 1103 590
rect 1107 586 1127 590
rect 1131 586 1159 590
rect 1163 586 1207 590
rect 1211 586 1215 590
rect 1219 586 1271 590
rect 1275 586 1287 590
rect 1291 586 1327 590
rect 1331 586 1359 590
rect 1363 586 1383 590
rect 1387 586 1431 590
rect 1435 586 1447 590
rect 1451 586 1503 590
rect 1507 586 1511 590
rect 1515 586 1575 590
rect 1579 586 1623 590
rect 1627 586 1663 590
rect 1667 586 1687 590
rect 91 585 1687 586
rect 1693 585 1694 591
rect 96 541 97 547
rect 103 546 1699 547
rect 103 542 111 546
rect 115 542 135 546
rect 139 542 167 546
rect 171 542 199 546
rect 203 542 215 546
rect 219 542 231 546
rect 235 542 271 546
rect 275 542 279 546
rect 283 542 327 546
rect 331 542 335 546
rect 339 542 375 546
rect 379 542 407 546
rect 411 542 431 546
rect 435 542 487 546
rect 491 542 495 546
rect 499 542 559 546
rect 563 542 623 546
rect 627 542 631 546
rect 635 542 687 546
rect 691 542 703 546
rect 707 542 751 546
rect 755 542 767 546
rect 771 542 815 546
rect 819 542 823 546
rect 827 542 879 546
rect 883 542 935 546
rect 939 542 943 546
rect 947 542 991 546
rect 995 542 1007 546
rect 1011 542 1047 546
rect 1051 542 1071 546
rect 1075 542 1103 546
rect 1107 542 1127 546
rect 1131 542 1159 546
rect 1163 542 1183 546
rect 1187 542 1215 546
rect 1219 542 1231 546
rect 1235 542 1271 546
rect 1275 542 1279 546
rect 1283 542 1327 546
rect 1331 542 1335 546
rect 1339 542 1383 546
rect 1387 542 1391 546
rect 1395 542 1447 546
rect 1451 542 1511 546
rect 1515 542 1575 546
rect 1579 542 1623 546
rect 1627 542 1663 546
rect 1667 542 1699 546
rect 103 541 1699 542
rect 1705 541 1706 547
rect 84 501 85 507
rect 91 506 1687 507
rect 91 502 111 506
rect 115 502 135 506
rect 139 502 167 506
rect 171 502 199 506
rect 203 502 231 506
rect 235 502 239 506
rect 243 502 279 506
rect 283 502 287 506
rect 291 502 327 506
rect 331 502 375 506
rect 379 502 423 506
rect 427 502 431 506
rect 435 502 479 506
rect 483 502 495 506
rect 499 502 543 506
rect 547 502 559 506
rect 563 502 615 506
rect 619 502 623 506
rect 627 502 687 506
rect 691 502 695 506
rect 699 502 751 506
rect 755 502 775 506
rect 779 502 815 506
rect 819 502 847 506
rect 851 502 879 506
rect 883 502 919 506
rect 923 502 943 506
rect 947 502 983 506
rect 987 502 1007 506
rect 1011 502 1039 506
rect 1043 502 1071 506
rect 1075 502 1095 506
rect 1099 502 1127 506
rect 1131 502 1143 506
rect 1147 502 1183 506
rect 1187 502 1191 506
rect 1195 502 1231 506
rect 1235 502 1239 506
rect 1243 502 1279 506
rect 1283 502 1287 506
rect 1291 502 1335 506
rect 1339 502 1383 506
rect 1387 502 1391 506
rect 1395 502 1431 506
rect 1435 502 1447 506
rect 1451 502 1479 506
rect 1483 502 1511 506
rect 1515 502 1535 506
rect 1539 502 1575 506
rect 1579 502 1591 506
rect 1595 502 1623 506
rect 1627 502 1663 506
rect 1667 502 1687 506
rect 91 501 1687 502
rect 1693 501 1694 507
rect 96 461 97 467
rect 103 466 1699 467
rect 103 462 111 466
rect 115 462 135 466
rect 139 462 151 466
rect 155 462 167 466
rect 171 462 199 466
rect 203 462 207 466
rect 211 462 239 466
rect 243 462 255 466
rect 259 462 287 466
rect 291 462 311 466
rect 315 462 327 466
rect 331 462 367 466
rect 371 462 375 466
rect 379 462 423 466
rect 427 462 439 466
rect 443 462 479 466
rect 483 462 519 466
rect 523 462 543 466
rect 547 462 599 466
rect 603 462 615 466
rect 619 462 679 466
rect 683 462 695 466
rect 699 462 759 466
rect 763 462 775 466
rect 779 462 839 466
rect 843 462 847 466
rect 851 462 911 466
rect 915 462 919 466
rect 923 462 983 466
rect 987 462 1039 466
rect 1043 462 1055 466
rect 1059 462 1095 466
rect 1099 462 1127 466
rect 1131 462 1143 466
rect 1147 462 1191 466
rect 1195 462 1199 466
rect 1203 462 1239 466
rect 1243 462 1263 466
rect 1267 462 1287 466
rect 1291 462 1319 466
rect 1323 462 1335 466
rect 1339 462 1375 466
rect 1379 462 1383 466
rect 1387 462 1431 466
rect 1435 462 1479 466
rect 1483 462 1495 466
rect 1499 462 1535 466
rect 1539 462 1591 466
rect 1595 462 1623 466
rect 1627 462 1663 466
rect 1667 462 1699 466
rect 103 461 1699 462
rect 1705 461 1706 467
rect 84 421 85 427
rect 91 426 1687 427
rect 91 422 111 426
rect 115 422 151 426
rect 155 422 175 426
rect 179 422 207 426
rect 211 422 223 426
rect 227 422 255 426
rect 259 422 271 426
rect 275 422 311 426
rect 315 422 319 426
rect 323 422 367 426
rect 371 422 415 426
rect 419 422 439 426
rect 443 422 471 426
rect 475 422 519 426
rect 523 422 527 426
rect 531 422 591 426
rect 595 422 599 426
rect 603 422 663 426
rect 667 422 679 426
rect 683 422 735 426
rect 739 422 759 426
rect 763 422 807 426
rect 811 422 839 426
rect 843 422 871 426
rect 875 422 911 426
rect 915 422 935 426
rect 939 422 983 426
rect 987 422 991 426
rect 995 422 1039 426
rect 1043 422 1055 426
rect 1059 422 1087 426
rect 1091 422 1127 426
rect 1131 422 1167 426
rect 1171 422 1199 426
rect 1203 422 1207 426
rect 1211 422 1247 426
rect 1251 422 1263 426
rect 1267 422 1287 426
rect 1291 422 1319 426
rect 1323 422 1335 426
rect 1339 422 1375 426
rect 1379 422 1383 426
rect 1387 422 1431 426
rect 1435 422 1495 426
rect 1499 422 1663 426
rect 1667 422 1687 426
rect 91 421 1687 422
rect 1693 421 1694 427
rect 96 377 97 383
rect 103 382 1699 383
rect 103 378 111 382
rect 115 378 135 382
rect 139 378 167 382
rect 171 378 175 382
rect 179 378 199 382
rect 203 378 223 382
rect 227 378 239 382
rect 243 378 271 382
rect 275 378 295 382
rect 299 378 319 382
rect 323 378 351 382
rect 355 378 367 382
rect 371 378 407 382
rect 411 378 415 382
rect 419 378 463 382
rect 467 378 471 382
rect 475 378 519 382
rect 523 378 527 382
rect 531 378 575 382
rect 579 378 591 382
rect 595 378 631 382
rect 635 378 663 382
rect 667 378 687 382
rect 691 378 735 382
rect 739 378 743 382
rect 747 378 799 382
rect 803 378 807 382
rect 811 378 855 382
rect 859 378 871 382
rect 875 378 919 382
rect 923 378 935 382
rect 939 378 983 382
rect 987 378 991 382
rect 995 378 1039 382
rect 1043 378 1087 382
rect 1091 378 1095 382
rect 1099 378 1127 382
rect 1131 378 1151 382
rect 1155 378 1167 382
rect 1171 378 1207 382
rect 1211 378 1247 382
rect 1251 378 1255 382
rect 1259 378 1287 382
rect 1291 378 1303 382
rect 1307 378 1335 382
rect 1339 378 1351 382
rect 1355 378 1383 382
rect 1387 378 1399 382
rect 1403 378 1447 382
rect 1451 378 1495 382
rect 1499 378 1543 382
rect 1547 378 1591 382
rect 1595 378 1623 382
rect 1627 378 1663 382
rect 1667 378 1699 382
rect 103 377 1699 378
rect 1705 377 1706 383
rect 84 337 85 343
rect 91 342 1687 343
rect 91 338 111 342
rect 115 338 135 342
rect 139 338 167 342
rect 171 338 199 342
rect 203 338 207 342
rect 211 338 239 342
rect 243 338 263 342
rect 267 338 295 342
rect 299 338 327 342
rect 331 338 351 342
rect 355 338 391 342
rect 395 338 407 342
rect 411 338 455 342
rect 459 338 463 342
rect 467 338 519 342
rect 523 338 575 342
rect 579 338 631 342
rect 635 338 687 342
rect 691 338 743 342
rect 747 338 751 342
rect 755 338 799 342
rect 803 338 815 342
rect 819 338 855 342
rect 859 338 879 342
rect 883 338 919 342
rect 923 338 951 342
rect 955 338 983 342
rect 987 338 1031 342
rect 1035 338 1039 342
rect 1043 338 1095 342
rect 1099 338 1111 342
rect 1115 338 1151 342
rect 1155 338 1191 342
rect 1195 338 1207 342
rect 1211 338 1255 342
rect 1259 338 1271 342
rect 1275 338 1303 342
rect 1307 338 1343 342
rect 1347 338 1351 342
rect 1355 338 1399 342
rect 1403 338 1407 342
rect 1411 338 1447 342
rect 1451 338 1463 342
rect 1467 338 1495 342
rect 1499 338 1519 342
rect 1523 338 1543 342
rect 1547 338 1583 342
rect 1587 338 1591 342
rect 1595 338 1623 342
rect 1627 338 1663 342
rect 1667 338 1687 342
rect 91 337 1687 338
rect 1693 337 1694 343
rect 96 297 97 303
rect 103 302 1699 303
rect 103 298 111 302
rect 115 298 135 302
rect 139 298 167 302
rect 171 298 207 302
rect 211 298 231 302
rect 235 298 263 302
rect 267 298 295 302
rect 299 298 327 302
rect 331 298 367 302
rect 371 298 391 302
rect 395 298 439 302
rect 443 298 455 302
rect 459 298 503 302
rect 507 298 519 302
rect 523 298 567 302
rect 571 298 575 302
rect 579 298 631 302
rect 635 298 687 302
rect 691 298 743 302
rect 747 298 751 302
rect 755 298 807 302
rect 811 298 815 302
rect 819 298 879 302
rect 883 298 951 302
rect 955 298 1031 302
rect 1035 298 1111 302
rect 1115 298 1191 302
rect 1195 298 1263 302
rect 1267 298 1271 302
rect 1275 298 1327 302
rect 1331 298 1343 302
rect 1347 298 1391 302
rect 1395 298 1407 302
rect 1411 298 1447 302
rect 1451 298 1463 302
rect 1467 298 1495 302
rect 1499 298 1519 302
rect 1523 298 1543 302
rect 1547 298 1583 302
rect 1587 298 1591 302
rect 1595 298 1623 302
rect 1627 298 1663 302
rect 1667 298 1699 302
rect 103 297 1699 298
rect 1705 297 1706 303
rect 84 253 85 259
rect 91 258 1687 259
rect 91 254 111 258
rect 115 254 135 258
rect 139 254 167 258
rect 171 254 175 258
rect 179 254 231 258
rect 235 254 247 258
rect 251 254 295 258
rect 299 254 319 258
rect 323 254 367 258
rect 371 254 383 258
rect 387 254 439 258
rect 443 254 447 258
rect 451 254 503 258
rect 507 254 519 258
rect 523 254 567 258
rect 571 254 591 258
rect 595 254 631 258
rect 635 254 663 258
rect 667 254 687 258
rect 691 254 743 258
rect 747 254 807 258
rect 811 254 823 258
rect 827 254 879 258
rect 883 254 895 258
rect 899 254 951 258
rect 955 254 967 258
rect 971 254 1031 258
rect 1035 254 1087 258
rect 1091 254 1111 258
rect 1115 254 1143 258
rect 1147 254 1191 258
rect 1195 254 1199 258
rect 1203 254 1255 258
rect 1259 254 1263 258
rect 1267 254 1311 258
rect 1315 254 1327 258
rect 1331 254 1367 258
rect 1371 254 1391 258
rect 1395 254 1415 258
rect 1419 254 1447 258
rect 1451 254 1463 258
rect 1467 254 1495 258
rect 1499 254 1519 258
rect 1523 254 1543 258
rect 1547 254 1575 258
rect 1579 254 1591 258
rect 1595 254 1623 258
rect 1627 254 1663 258
rect 1667 254 1687 258
rect 91 253 1687 254
rect 1693 253 1694 259
rect 96 213 97 219
rect 103 218 1699 219
rect 103 214 111 218
rect 115 214 135 218
rect 139 214 167 218
rect 171 214 175 218
rect 179 214 207 218
rect 211 214 247 218
rect 251 214 255 218
rect 259 214 303 218
rect 307 214 319 218
rect 323 214 343 218
rect 347 214 375 218
rect 379 214 383 218
rect 387 214 415 218
rect 419 214 447 218
rect 451 214 471 218
rect 475 214 519 218
rect 523 214 535 218
rect 539 214 591 218
rect 595 214 615 218
rect 619 214 663 218
rect 667 214 695 218
rect 699 214 743 218
rect 747 214 775 218
rect 779 214 823 218
rect 827 214 855 218
rect 859 214 895 218
rect 899 214 927 218
rect 931 214 967 218
rect 971 214 999 218
rect 1003 214 1031 218
rect 1035 214 1071 218
rect 1075 214 1087 218
rect 1091 214 1143 218
rect 1147 214 1199 218
rect 1203 214 1215 218
rect 1219 214 1255 218
rect 1259 214 1287 218
rect 1291 214 1311 218
rect 1315 214 1351 218
rect 1355 214 1367 218
rect 1371 214 1415 218
rect 1419 214 1463 218
rect 1467 214 1471 218
rect 1475 214 1519 218
rect 1523 214 1527 218
rect 1531 214 1575 218
rect 1579 214 1583 218
rect 1587 214 1623 218
rect 1627 214 1663 218
rect 1667 214 1699 218
rect 103 213 1699 214
rect 1705 213 1706 219
rect 84 173 85 179
rect 91 178 1687 179
rect 91 174 111 178
rect 115 174 135 178
rect 139 174 167 178
rect 171 174 175 178
rect 179 174 207 178
rect 211 174 231 178
rect 235 174 255 178
rect 259 174 287 178
rect 291 174 303 178
rect 307 174 343 178
rect 347 174 375 178
rect 379 174 399 178
rect 403 174 415 178
rect 419 174 455 178
rect 459 174 471 178
rect 475 174 511 178
rect 515 174 535 178
rect 539 174 575 178
rect 579 174 615 178
rect 619 174 639 178
rect 643 174 695 178
rect 699 174 703 178
rect 707 174 767 178
rect 771 174 775 178
rect 779 174 831 178
rect 835 174 855 178
rect 859 174 895 178
rect 899 174 927 178
rect 931 174 951 178
rect 955 174 999 178
rect 1003 174 1015 178
rect 1019 174 1071 178
rect 1075 174 1079 178
rect 1083 174 1143 178
rect 1147 174 1207 178
rect 1211 174 1215 178
rect 1219 174 1279 178
rect 1283 174 1287 178
rect 1291 174 1351 178
rect 1355 174 1415 178
rect 1419 174 1423 178
rect 1427 174 1471 178
rect 1475 174 1495 178
rect 1499 174 1527 178
rect 1531 174 1567 178
rect 1571 174 1583 178
rect 1587 174 1623 178
rect 1627 174 1663 178
rect 1667 174 1687 178
rect 91 173 1687 174
rect 1693 173 1694 179
rect 96 117 97 123
rect 103 122 1699 123
rect 103 118 111 122
rect 115 118 135 122
rect 139 118 167 122
rect 171 118 175 122
rect 179 118 199 122
rect 203 118 231 122
rect 235 118 263 122
rect 267 118 287 122
rect 291 118 295 122
rect 299 118 327 122
rect 331 118 343 122
rect 347 118 359 122
rect 363 118 391 122
rect 395 118 399 122
rect 403 118 423 122
rect 427 118 455 122
rect 459 118 463 122
rect 467 118 503 122
rect 507 118 511 122
rect 515 118 543 122
rect 547 118 575 122
rect 579 118 607 122
rect 611 118 639 122
rect 643 118 671 122
rect 675 118 703 122
rect 707 118 735 122
rect 739 118 767 122
rect 771 118 799 122
rect 803 118 831 122
rect 835 118 863 122
rect 867 118 895 122
rect 899 118 935 122
rect 939 118 951 122
rect 955 118 975 122
rect 979 118 1015 122
rect 1019 118 1063 122
rect 1067 118 1079 122
rect 1083 118 1103 122
rect 1107 118 1143 122
rect 1147 118 1183 122
rect 1187 118 1207 122
rect 1211 118 1223 122
rect 1227 118 1263 122
rect 1267 118 1279 122
rect 1283 118 1295 122
rect 1299 118 1335 122
rect 1339 118 1351 122
rect 1355 118 1375 122
rect 1379 118 1415 122
rect 1419 118 1423 122
rect 1427 118 1455 122
rect 1459 118 1495 122
rect 1499 118 1503 122
rect 1507 118 1551 122
rect 1555 118 1567 122
rect 1571 118 1591 122
rect 1595 118 1623 122
rect 1627 118 1663 122
rect 1667 118 1699 122
rect 103 117 1699 118
rect 1705 117 1706 123
rect 84 77 85 83
rect 91 82 1687 83
rect 91 78 111 82
rect 115 78 135 82
rect 139 78 167 82
rect 171 78 199 82
rect 203 78 231 82
rect 235 78 263 82
rect 267 78 295 82
rect 299 78 327 82
rect 331 78 359 82
rect 363 78 391 82
rect 395 78 423 82
rect 427 78 463 82
rect 467 78 503 82
rect 507 78 543 82
rect 547 78 575 82
rect 579 78 607 82
rect 611 78 639 82
rect 643 78 671 82
rect 675 78 703 82
rect 707 78 735 82
rect 739 78 767 82
rect 771 78 799 82
rect 803 78 831 82
rect 835 78 863 82
rect 867 78 895 82
rect 899 78 935 82
rect 939 78 975 82
rect 979 78 1015 82
rect 1019 78 1063 82
rect 1067 78 1103 82
rect 1107 78 1143 82
rect 1147 78 1183 82
rect 1187 78 1223 82
rect 1227 78 1263 82
rect 1267 78 1295 82
rect 1299 78 1335 82
rect 1339 78 1375 82
rect 1379 78 1415 82
rect 1419 78 1455 82
rect 1459 78 1503 82
rect 1507 78 1551 82
rect 1555 78 1591 82
rect 1595 78 1623 82
rect 1627 78 1663 82
rect 1667 78 1687 82
rect 91 77 1687 78
rect 1693 77 1694 83
<< m5c >>
rect 97 1713 103 1719
rect 1699 1713 1705 1719
rect 85 1673 91 1679
rect 1687 1673 1693 1679
rect 97 1633 103 1639
rect 1699 1633 1705 1639
rect 85 1593 91 1599
rect 1687 1593 1693 1599
rect 97 1553 103 1559
rect 1699 1553 1705 1559
rect 85 1509 91 1515
rect 1687 1509 1693 1515
rect 97 1469 103 1475
rect 1699 1469 1705 1475
rect 85 1425 91 1431
rect 1687 1425 1693 1431
rect 97 1385 103 1391
rect 1699 1385 1705 1391
rect 85 1345 91 1351
rect 1687 1345 1693 1351
rect 97 1301 103 1307
rect 1699 1301 1705 1307
rect 85 1261 91 1267
rect 1687 1261 1693 1267
rect 97 1217 103 1223
rect 1699 1217 1705 1223
rect 85 1173 91 1179
rect 1687 1173 1693 1179
rect 97 1129 103 1135
rect 1699 1129 1705 1135
rect 85 1085 91 1091
rect 1687 1085 1693 1091
rect 97 1041 103 1047
rect 1699 1041 1705 1047
rect 85 1001 91 1007
rect 1687 1001 1693 1007
rect 97 961 103 967
rect 1699 961 1705 967
rect 85 917 91 923
rect 1687 917 1693 923
rect 97 873 103 879
rect 1699 873 1705 879
rect 85 833 91 839
rect 1687 833 1693 839
rect 97 789 103 795
rect 1699 789 1705 795
rect 85 749 91 755
rect 1687 749 1693 755
rect 97 705 103 711
rect 1699 705 1705 711
rect 85 665 91 671
rect 1687 665 1693 671
rect 97 625 103 631
rect 1699 625 1705 631
rect 85 585 91 591
rect 1687 585 1693 591
rect 97 541 103 547
rect 1699 541 1705 547
rect 85 501 91 507
rect 1687 501 1693 507
rect 97 461 103 467
rect 1699 461 1705 467
rect 85 421 91 427
rect 1687 421 1693 427
rect 97 377 103 383
rect 1699 377 1705 383
rect 85 337 91 343
rect 1687 337 1693 343
rect 97 297 103 303
rect 1699 297 1705 303
rect 85 253 91 259
rect 1687 253 1693 259
rect 97 213 103 219
rect 1699 213 1705 219
rect 85 173 91 179
rect 1687 173 1693 179
rect 97 117 103 123
rect 1699 117 1705 123
rect 85 77 91 83
rect 1687 77 1693 83
<< m5 >>
rect 84 1679 92 1728
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1599 92 1673
rect 84 1593 85 1599
rect 91 1593 92 1599
rect 84 1515 92 1593
rect 84 1509 85 1515
rect 91 1509 92 1515
rect 84 1431 92 1509
rect 84 1425 85 1431
rect 91 1425 92 1431
rect 84 1351 92 1425
rect 84 1345 85 1351
rect 91 1345 92 1351
rect 84 1267 92 1345
rect 84 1261 85 1267
rect 91 1261 92 1267
rect 84 1179 92 1261
rect 84 1173 85 1179
rect 91 1173 92 1179
rect 84 1091 92 1173
rect 84 1085 85 1091
rect 91 1085 92 1091
rect 84 1007 92 1085
rect 84 1001 85 1007
rect 91 1001 92 1007
rect 84 923 92 1001
rect 84 917 85 923
rect 91 917 92 923
rect 84 839 92 917
rect 84 833 85 839
rect 91 833 92 839
rect 84 755 92 833
rect 84 749 85 755
rect 91 749 92 755
rect 84 671 92 749
rect 84 665 85 671
rect 91 665 92 671
rect 84 591 92 665
rect 84 585 85 591
rect 91 585 92 591
rect 84 507 92 585
rect 84 501 85 507
rect 91 501 92 507
rect 84 427 92 501
rect 84 421 85 427
rect 91 421 92 427
rect 84 343 92 421
rect 84 337 85 343
rect 91 337 92 343
rect 84 259 92 337
rect 84 253 85 259
rect 91 253 92 259
rect 84 179 92 253
rect 84 173 85 179
rect 91 173 92 179
rect 84 83 92 173
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 1719 104 1728
rect 96 1713 97 1719
rect 103 1713 104 1719
rect 96 1639 104 1713
rect 96 1633 97 1639
rect 103 1633 104 1639
rect 96 1559 104 1633
rect 96 1553 97 1559
rect 103 1553 104 1559
rect 96 1475 104 1553
rect 96 1469 97 1475
rect 103 1469 104 1475
rect 96 1391 104 1469
rect 96 1385 97 1391
rect 103 1385 104 1391
rect 96 1307 104 1385
rect 96 1301 97 1307
rect 103 1301 104 1307
rect 96 1223 104 1301
rect 96 1217 97 1223
rect 103 1217 104 1223
rect 96 1135 104 1217
rect 96 1129 97 1135
rect 103 1129 104 1135
rect 96 1047 104 1129
rect 96 1041 97 1047
rect 103 1041 104 1047
rect 96 967 104 1041
rect 96 961 97 967
rect 103 961 104 967
rect 96 879 104 961
rect 96 873 97 879
rect 103 873 104 879
rect 96 795 104 873
rect 96 789 97 795
rect 103 789 104 795
rect 96 711 104 789
rect 96 705 97 711
rect 103 705 104 711
rect 96 631 104 705
rect 96 625 97 631
rect 103 625 104 631
rect 96 547 104 625
rect 96 541 97 547
rect 103 541 104 547
rect 96 467 104 541
rect 96 461 97 467
rect 103 461 104 467
rect 96 383 104 461
rect 96 377 97 383
rect 103 377 104 383
rect 96 303 104 377
rect 96 297 97 303
rect 103 297 104 303
rect 96 219 104 297
rect 96 213 97 219
rect 103 213 104 219
rect 96 123 104 213
rect 96 117 97 123
rect 103 117 104 123
rect 96 72 104 117
rect 1686 1679 1694 1728
rect 1686 1673 1687 1679
rect 1693 1673 1694 1679
rect 1686 1599 1694 1673
rect 1686 1593 1687 1599
rect 1693 1593 1694 1599
rect 1686 1515 1694 1593
rect 1686 1509 1687 1515
rect 1693 1509 1694 1515
rect 1686 1431 1694 1509
rect 1686 1425 1687 1431
rect 1693 1425 1694 1431
rect 1686 1351 1694 1425
rect 1686 1345 1687 1351
rect 1693 1345 1694 1351
rect 1686 1267 1694 1345
rect 1686 1261 1687 1267
rect 1693 1261 1694 1267
rect 1686 1179 1694 1261
rect 1686 1173 1687 1179
rect 1693 1173 1694 1179
rect 1686 1091 1694 1173
rect 1686 1085 1687 1091
rect 1693 1085 1694 1091
rect 1686 1007 1694 1085
rect 1686 1001 1687 1007
rect 1693 1001 1694 1007
rect 1686 923 1694 1001
rect 1686 917 1687 923
rect 1693 917 1694 923
rect 1686 839 1694 917
rect 1686 833 1687 839
rect 1693 833 1694 839
rect 1686 755 1694 833
rect 1686 749 1687 755
rect 1693 749 1694 755
rect 1686 671 1694 749
rect 1686 665 1687 671
rect 1693 665 1694 671
rect 1686 591 1694 665
rect 1686 585 1687 591
rect 1693 585 1694 591
rect 1686 507 1694 585
rect 1686 501 1687 507
rect 1693 501 1694 507
rect 1686 427 1694 501
rect 1686 421 1687 427
rect 1693 421 1694 427
rect 1686 343 1694 421
rect 1686 337 1687 343
rect 1693 337 1694 343
rect 1686 259 1694 337
rect 1686 253 1687 259
rect 1693 253 1694 259
rect 1686 179 1694 253
rect 1686 173 1687 179
rect 1693 173 1694 179
rect 1686 83 1694 173
rect 1686 77 1687 83
rect 1693 77 1694 83
rect 1686 72 1694 77
rect 1698 1719 1706 1728
rect 1698 1713 1699 1719
rect 1705 1713 1706 1719
rect 1698 1639 1706 1713
rect 1698 1633 1699 1639
rect 1705 1633 1706 1639
rect 1698 1559 1706 1633
rect 1698 1553 1699 1559
rect 1705 1553 1706 1559
rect 1698 1475 1706 1553
rect 1698 1469 1699 1475
rect 1705 1469 1706 1475
rect 1698 1391 1706 1469
rect 1698 1385 1699 1391
rect 1705 1385 1706 1391
rect 1698 1307 1706 1385
rect 1698 1301 1699 1307
rect 1705 1301 1706 1307
rect 1698 1223 1706 1301
rect 1698 1217 1699 1223
rect 1705 1217 1706 1223
rect 1698 1135 1706 1217
rect 1698 1129 1699 1135
rect 1705 1129 1706 1135
rect 1698 1047 1706 1129
rect 1698 1041 1699 1047
rect 1705 1041 1706 1047
rect 1698 967 1706 1041
rect 1698 961 1699 967
rect 1705 961 1706 967
rect 1698 879 1706 961
rect 1698 873 1699 879
rect 1705 873 1706 879
rect 1698 795 1706 873
rect 1698 789 1699 795
rect 1705 789 1706 795
rect 1698 711 1706 789
rect 1698 705 1699 711
rect 1705 705 1706 711
rect 1698 631 1706 705
rect 1698 625 1699 631
rect 1705 625 1706 631
rect 1698 547 1706 625
rect 1698 541 1699 547
rect 1705 541 1706 547
rect 1698 467 1706 541
rect 1698 461 1699 467
rect 1705 461 1706 467
rect 1698 383 1706 461
rect 1698 377 1699 383
rect 1705 377 1706 383
rect 1698 303 1706 377
rect 1698 297 1699 303
rect 1705 297 1706 303
rect 1698 219 1706 297
rect 1698 213 1699 219
rect 1705 213 1706 219
rect 1698 123 1706 213
rect 1698 117 1699 123
rect 1705 117 1706 123
rect 1698 72 1706 117
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__77
timestamp 1731220534
transform 1 0 1656 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220534
transform 1 0 104 0 1 1680
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220534
transform 1 0 1656 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220534
transform 1 0 104 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220534
transform 1 0 1656 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220534
transform 1 0 104 0 1 1600
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220534
transform 1 0 1656 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220534
transform 1 0 104 0 -1 1592
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220534
transform 1 0 1656 0 1 1520
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220534
transform 1 0 104 0 1 1520
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220534
transform 1 0 1656 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220534
transform 1 0 104 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220534
transform 1 0 1656 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220534
transform 1 0 104 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220534
transform 1 0 1656 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220534
transform 1 0 104 0 -1 1424
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220534
transform 1 0 1656 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220534
transform 1 0 104 0 1 1352
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220534
transform 1 0 1656 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220534
transform 1 0 104 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220534
transform 1 0 1656 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220534
transform 1 0 104 0 1 1268
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220534
transform 1 0 1656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220534
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220534
transform 1 0 1656 0 1 1184
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220534
transform 1 0 104 0 1 1184
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220534
transform 1 0 1656 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220534
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220534
transform 1 0 1656 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220534
transform 1 0 104 0 1 1096
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220534
transform 1 0 1656 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220534
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220534
transform 1 0 1656 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220534
transform 1 0 104 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220534
transform 1 0 1656 0 -1 1000
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220534
transform 1 0 104 0 -1 1000
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220534
transform 1 0 1656 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220534
transform 1 0 104 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220534
transform 1 0 1656 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220534
transform 1 0 104 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220534
transform 1 0 1656 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220534
transform 1 0 104 0 1 840
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220534
transform 1 0 1656 0 -1 832
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220534
transform 1 0 104 0 -1 832
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220534
transform 1 0 1656 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220534
transform 1 0 104 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220534
transform 1 0 1656 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220534
transform 1 0 104 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220534
transform 1 0 1656 0 1 672
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220534
transform 1 0 104 0 1 672
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220534
transform 1 0 1656 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220534
transform 1 0 104 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220534
transform 1 0 1656 0 1 592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220534
transform 1 0 104 0 1 592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220534
transform 1 0 1656 0 -1 584
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220534
transform 1 0 104 0 -1 584
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220534
transform 1 0 1656 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220534
transform 1 0 104 0 1 508
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220534
transform 1 0 1656 0 -1 500
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220534
transform 1 0 104 0 -1 500
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220534
transform 1 0 1656 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220534
transform 1 0 104 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220534
transform 1 0 1656 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220534
transform 1 0 104 0 -1 420
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220534
transform 1 0 1656 0 1 344
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220534
transform 1 0 104 0 1 344
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220534
transform 1 0 1656 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220534
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220534
transform 1 0 1656 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220534
transform 1 0 104 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220534
transform 1 0 1656 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220534
transform 1 0 104 0 -1 252
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220534
transform 1 0 1656 0 1 180
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220534
transform 1 0 104 0 1 180
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220534
transform 1 0 1656 0 -1 172
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220534
transform 1 0 104 0 -1 172
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220534
transform 1 0 1656 0 1 84
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220534
transform 1 0 104 0 1 84
box 7 3 12 24
use _0_0std_0_0cells_0_0INVX1  tst_5999_6
timestamp 1731220534
transform 1 0 1584 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5998_6
timestamp 1731220534
transform 1 0 1616 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5997_6
timestamp 1731220534
transform 1 0 1616 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5996_6
timestamp 1731220534
transform 1 0 1616 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5995_6
timestamp 1731220534
transform 1 0 1576 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5994_6
timestamp 1731220534
transform 1 0 1520 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5993_6
timestamp 1731220534
transform 1 0 1616 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5992_6
timestamp 1731220534
transform 1 0 1568 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5991_6
timestamp 1731220534
transform 1 0 1512 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5990_6
timestamp 1731220534
transform 1 0 1456 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5989_6
timestamp 1731220534
transform 1 0 1464 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5988_6
timestamp 1731220534
transform 1 0 1408 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5987_6
timestamp 1731220534
transform 1 0 1416 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5986_6
timestamp 1731220534
transform 1 0 1488 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5985_6
timestamp 1731220534
transform 1 0 1560 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5984_6
timestamp 1731220534
transform 1 0 1544 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5983_6
timestamp 1731220534
transform 1 0 1496 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5982_6
timestamp 1731220534
transform 1 0 1448 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5981_6
timestamp 1731220534
transform 1 0 1408 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5980_6
timestamp 1731220534
transform 1 0 1368 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5979_6
timestamp 1731220534
transform 1 0 1328 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5978_6
timestamp 1731220534
transform 1 0 1288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5977_6
timestamp 1731220534
transform 1 0 1256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5976_6
timestamp 1731220534
transform 1 0 1216 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5975_6
timestamp 1731220534
transform 1 0 1176 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5974_6
timestamp 1731220534
transform 1 0 1200 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5973_6
timestamp 1731220534
transform 1 0 1272 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5972_6
timestamp 1731220534
transform 1 0 1344 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5971_6
timestamp 1731220534
transform 1 0 1344 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5970_6
timestamp 1731220534
transform 1 0 1280 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5969_6
timestamp 1731220534
transform 1 0 1304 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5968_6
timestamp 1731220534
transform 1 0 1360 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5967_6
timestamp 1731220534
transform 1 0 1408 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5966_6
timestamp 1731220534
transform 1 0 1384 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5965_6
timestamp 1731220534
transform 1 0 1320 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5964_6
timestamp 1731220534
transform 1 0 1440 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5963_6
timestamp 1731220534
transform 1 0 1488 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5962_6
timestamp 1731220534
transform 1 0 1536 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5961_6
timestamp 1731220534
transform 1 0 1584 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5960_6
timestamp 1731220534
transform 1 0 1616 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5959_6
timestamp 1731220534
transform 1 0 1616 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5958_6
timestamp 1731220534
transform 1 0 1616 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5957_6
timestamp 1731220534
transform 1 0 1584 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5956_6
timestamp 1731220534
transform 1 0 1536 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5955_6
timestamp 1731220534
transform 1 0 1488 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5954_6
timestamp 1731220534
transform 1 0 1576 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5953_6
timestamp 1731220534
transform 1 0 1512 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5952_6
timestamp 1731220534
transform 1 0 1456 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5951_6
timestamp 1731220534
transform 1 0 1400 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5950_6
timestamp 1731220534
transform 1 0 1336 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5949_6
timestamp 1731220534
transform 1 0 1440 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5948_6
timestamp 1731220534
transform 1 0 1392 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5947_6
timestamp 1731220534
transform 1 0 1344 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5946_6
timestamp 1731220534
transform 1 0 1296 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5945_6
timestamp 1731220534
transform 1 0 1248 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5944_6
timestamp 1731220534
transform 1 0 1200 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5943_6
timestamp 1731220534
transform 1 0 1160 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5942_6
timestamp 1731220534
transform 1 0 1200 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5941_6
timestamp 1731220534
transform 1 0 1240 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5940_6
timestamp 1731220534
transform 1 0 1280 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5939_6
timestamp 1731220534
transform 1 0 1376 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5938_6
timestamp 1731220534
transform 1 0 1328 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5937_6
timestamp 1731220534
transform 1 0 1312 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5936_6
timestamp 1731220534
transform 1 0 1256 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5935_6
timestamp 1731220534
transform 1 0 1368 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5934_6
timestamp 1731220534
transform 1 0 1424 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5933_6
timestamp 1731220534
transform 1 0 1488 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5932_6
timestamp 1731220534
transform 1 0 1472 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5931_6
timestamp 1731220534
transform 1 0 1424 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5930_6
timestamp 1731220534
transform 1 0 1528 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5929_6
timestamp 1731220534
transform 1 0 1616 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5928_6
timestamp 1731220534
transform 1 0 1584 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5927_6
timestamp 1731220534
transform 1 0 1568 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5926_6
timestamp 1731220534
transform 1 0 1616 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5925_6
timestamp 1731220534
transform 1 0 1616 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5924_6
timestamp 1731220534
transform 1 0 1616 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5923_6
timestamp 1731220534
transform 1 0 1616 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5922_6
timestamp 1731220534
transform 1 0 1616 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5921_6
timestamp 1731220534
transform 1 0 1576 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5920_6
timestamp 1731220534
transform 1 0 1616 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5919_6
timestamp 1731220534
transform 1 0 1576 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5918_6
timestamp 1731220534
transform 1 0 1520 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5917_6
timestamp 1731220534
transform 1 0 1464 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5916_6
timestamp 1731220534
transform 1 0 1464 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5915_6
timestamp 1731220534
transform 1 0 1552 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5914_6
timestamp 1731220534
transform 1 0 1568 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5913_6
timestamp 1731220534
transform 1 0 1496 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5912_6
timestamp 1731220534
transform 1 0 1424 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5911_6
timestamp 1731220534
transform 1 0 1352 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5910_6
timestamp 1731220534
transform 1 0 1568 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5909_6
timestamp 1731220534
transform 1 0 1504 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5908_6
timestamp 1731220534
transform 1 0 1440 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5907_6
timestamp 1731220534
transform 1 0 1376 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5906_6
timestamp 1731220534
transform 1 0 1320 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5905_6
timestamp 1731220534
transform 1 0 1504 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5904_6
timestamp 1731220534
transform 1 0 1440 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5903_6
timestamp 1731220534
transform 1 0 1384 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5902_6
timestamp 1731220534
transform 1 0 1328 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5901_6
timestamp 1731220534
transform 1 0 1272 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5900_6
timestamp 1731220534
transform 1 0 1224 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5899_6
timestamp 1731220534
transform 1 0 1376 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5898_6
timestamp 1731220534
transform 1 0 1328 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5897_6
timestamp 1731220534
transform 1 0 1280 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5896_6
timestamp 1731220534
transform 1 0 1232 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5895_6
timestamp 1731220534
transform 1 0 1184 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5894_6
timestamp 1731220534
transform 1 0 1136 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5893_6
timestamp 1731220534
transform 1 0 1088 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5892_6
timestamp 1731220534
transform 1 0 1032 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5891_6
timestamp 1731220534
transform 1 0 976 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5890_6
timestamp 1731220534
transform 1 0 912 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5889_6
timestamp 1731220534
transform 1 0 1064 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5888_6
timestamp 1731220534
transform 1 0 1120 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5887_6
timestamp 1731220534
transform 1 0 1176 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5886_6
timestamp 1731220534
transform 1 0 1152 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5885_6
timestamp 1731220534
transform 1 0 1208 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5884_6
timestamp 1731220534
transform 1 0 1264 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5883_6
timestamp 1731220534
transform 1 0 1280 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5882_6
timestamp 1731220534
transform 1 0 1200 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5881_6
timestamp 1731220534
transform 1 0 1208 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5880_6
timestamp 1731220534
transform 1 0 1288 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5879_6
timestamp 1731220534
transform 1 0 1376 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5878_6
timestamp 1731220534
transform 1 0 1408 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5877_6
timestamp 1731220534
transform 1 0 1344 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5876_6
timestamp 1731220534
transform 1 0 1280 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5875_6
timestamp 1731220534
transform 1 0 1216 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5874_6
timestamp 1731220534
transform 1 0 1152 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5873_6
timestamp 1731220534
transform 1 0 1232 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5872_6
timestamp 1731220534
transform 1 0 1288 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5871_6
timestamp 1731220534
transform 1 0 1344 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5870_6
timestamp 1731220534
transform 1 0 1400 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5869_6
timestamp 1731220534
transform 1 0 1456 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5868_6
timestamp 1731220534
transform 1 0 1512 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5867_6
timestamp 1731220534
transform 1 0 1464 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5866_6
timestamp 1731220534
transform 1 0 1408 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5865_6
timestamp 1731220534
transform 1 0 1352 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5864_6
timestamp 1731220534
transform 1 0 1520 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5863_6
timestamp 1731220534
transform 1 0 1584 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5862_6
timestamp 1731220534
transform 1 0 1584 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5861_6
timestamp 1731220534
transform 1 0 1528 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5860_6
timestamp 1731220534
transform 1 0 1472 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5859_6
timestamp 1731220534
transform 1 0 1416 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5858_6
timestamp 1731220534
transform 1 0 1360 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5857_6
timestamp 1731220534
transform 1 0 1304 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5856_6
timestamp 1731220534
transform 1 0 1456 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5855_6
timestamp 1731220534
transform 1 0 1392 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5854_6
timestamp 1731220534
transform 1 0 1336 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5853_6
timestamp 1731220534
transform 1 0 1280 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5852_6
timestamp 1731220534
transform 1 0 1224 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5851_6
timestamp 1731220534
transform 1 0 1160 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5850_6
timestamp 1731220534
transform 1 0 1376 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5849_6
timestamp 1731220534
transform 1 0 1312 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5848_6
timestamp 1731220534
transform 1 0 1248 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5847_6
timestamp 1731220534
transform 1 0 1192 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5846_6
timestamp 1731220534
transform 1 0 1136 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5845_6
timestamp 1731220534
transform 1 0 1224 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5844_6
timestamp 1731220534
transform 1 0 1280 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5843_6
timestamp 1731220534
transform 1 0 1336 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5842_6
timestamp 1731220534
transform 1 0 1280 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5841_6
timestamp 1731220534
transform 1 0 1336 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5840_6
timestamp 1731220534
transform 1 0 1392 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5839_6
timestamp 1731220534
transform 1 0 1376 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5838_6
timestamp 1731220534
transform 1 0 1328 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5837_6
timestamp 1731220534
transform 1 0 1424 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5836_6
timestamp 1731220534
transform 1 0 1472 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5835_6
timestamp 1731220534
transform 1 0 1528 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5834_6
timestamp 1731220534
transform 1 0 1536 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5833_6
timestamp 1731220534
transform 1 0 1488 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5832_6
timestamp 1731220534
transform 1 0 1440 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5831_6
timestamp 1731220534
transform 1 0 1424 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5830_6
timestamp 1731220534
transform 1 0 1384 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5829_6
timestamp 1731220534
transform 1 0 1464 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5828_6
timestamp 1731220534
transform 1 0 1504 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5827_6
timestamp 1731220534
transform 1 0 1544 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5826_6
timestamp 1731220534
transform 1 0 1616 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5825_6
timestamp 1731220534
transform 1 0 1584 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5824_6
timestamp 1731220534
transform 1 0 1584 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5823_6
timestamp 1731220534
transform 1 0 1616 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5822_6
timestamp 1731220534
transform 1 0 1616 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5821_6
timestamp 1731220534
transform 1 0 1584 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5820_6
timestamp 1731220534
transform 1 0 1616 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5819_6
timestamp 1731220534
transform 1 0 1616 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5818_6
timestamp 1731220534
transform 1 0 1584 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5817_6
timestamp 1731220534
transform 1 0 1536 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5816_6
timestamp 1731220534
transform 1 0 1584 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5815_6
timestamp 1731220534
transform 1 0 1544 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5814_6
timestamp 1731220534
transform 1 0 1496 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5813_6
timestamp 1731220534
transform 1 0 1456 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5812_6
timestamp 1731220534
transform 1 0 1408 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5811_6
timestamp 1731220534
transform 1 0 1352 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5810_6
timestamp 1731220534
transform 1 0 1488 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5809_6
timestamp 1731220534
transform 1 0 1440 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5808_6
timestamp 1731220534
transform 1 0 1384 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5807_6
timestamp 1731220534
transform 1 0 1328 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5806_6
timestamp 1731220534
transform 1 0 1552 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5805_6
timestamp 1731220534
transform 1 0 1472 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5804_6
timestamp 1731220534
transform 1 0 1400 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5803_6
timestamp 1731220534
transform 1 0 1336 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5802_6
timestamp 1731220534
transform 1 0 1272 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5801_6
timestamp 1731220534
transform 1 0 1208 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5800_6
timestamp 1731220534
transform 1 0 1536 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5799_6
timestamp 1731220534
transform 1 0 1440 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5798_6
timestamp 1731220534
transform 1 0 1352 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5797_6
timestamp 1731220534
transform 1 0 1272 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5796_6
timestamp 1731220534
transform 1 0 1200 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5795_6
timestamp 1731220534
transform 1 0 1136 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5794_6
timestamp 1731220534
transform 1 0 1528 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5793_6
timestamp 1731220534
transform 1 0 1416 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5792_6
timestamp 1731220534
transform 1 0 1312 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5791_6
timestamp 1731220534
transform 1 0 1224 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5790_6
timestamp 1731220534
transform 1 0 1152 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5789_6
timestamp 1731220534
transform 1 0 1088 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5788_6
timestamp 1731220534
transform 1 0 1136 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5787_6
timestamp 1731220534
transform 1 0 1200 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5786_6
timestamp 1731220534
transform 1 0 1272 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5785_6
timestamp 1731220534
transform 1 0 1536 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5784_6
timestamp 1731220534
transform 1 0 1440 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5783_6
timestamp 1731220534
transform 1 0 1352 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5782_6
timestamp 1731220534
transform 1 0 1336 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5781_6
timestamp 1731220534
transform 1 0 1272 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5780_6
timestamp 1731220534
transform 1 0 1208 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5779_6
timestamp 1731220534
transform 1 0 1400 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5778_6
timestamp 1731220534
transform 1 0 1552 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5777_6
timestamp 1731220534
transform 1 0 1472 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5776_6
timestamp 1731220534
transform 1 0 1424 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5775_6
timestamp 1731220534
transform 1 0 1360 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5774_6
timestamp 1731220534
transform 1 0 1296 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5773_6
timestamp 1731220534
transform 1 0 1560 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5772_6
timestamp 1731220534
transform 1 0 1488 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5771_6
timestamp 1731220534
transform 1 0 1456 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5770_6
timestamp 1731220534
transform 1 0 1408 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5769_6
timestamp 1731220534
transform 1 0 1352 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5768_6
timestamp 1731220534
transform 1 0 1496 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5767_6
timestamp 1731220534
transform 1 0 1552 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5766_6
timestamp 1731220534
transform 1 0 1544 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5765_6
timestamp 1731220534
transform 1 0 1584 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5764_6
timestamp 1731220534
transform 1 0 1616 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5763_6
timestamp 1731220534
transform 1 0 1616 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5762_6
timestamp 1731220534
transform 1 0 1616 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5761_6
timestamp 1731220534
transform 1 0 1616 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5760_6
timestamp 1731220534
transform 1 0 1616 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5759_6
timestamp 1731220534
transform 1 0 1616 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5758_6
timestamp 1731220534
transform 1 0 1616 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5757_6
timestamp 1731220534
transform 1 0 1616 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5756_6
timestamp 1731220534
transform 1 0 1616 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5755_6
timestamp 1731220534
transform 1 0 1616 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5754_6
timestamp 1731220534
transform 1 0 1616 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5753_6
timestamp 1731220534
transform 1 0 1616 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5752_6
timestamp 1731220534
transform 1 0 1616 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5751_6
timestamp 1731220534
transform 1 0 1576 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5750_6
timestamp 1731220534
transform 1 0 1520 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5749_6
timestamp 1731220534
transform 1 0 1576 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5748_6
timestamp 1731220534
transform 1 0 1576 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5747_6
timestamp 1731220534
transform 1 0 1520 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5746_6
timestamp 1731220534
transform 1 0 1464 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5745_6
timestamp 1731220534
transform 1 0 1400 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5744_6
timestamp 1731220534
transform 1 0 1328 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5743_6
timestamp 1731220534
transform 1 0 1344 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5742_6
timestamp 1731220534
transform 1 0 1464 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5741_6
timestamp 1731220534
transform 1 0 1408 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5740_6
timestamp 1731220534
transform 1 0 1392 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5739_6
timestamp 1731220534
transform 1 0 1472 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5738_6
timestamp 1731220534
transform 1 0 1552 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5737_6
timestamp 1731220534
transform 1 0 1512 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5736_6
timestamp 1731220534
transform 1 0 1448 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5735_6
timestamp 1731220534
transform 1 0 1384 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5734_6
timestamp 1731220534
transform 1 0 1512 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5733_6
timestamp 1731220534
transform 1 0 1464 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5732_6
timestamp 1731220534
transform 1 0 1416 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5731_6
timestamp 1731220534
transform 1 0 1368 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5730_6
timestamp 1731220534
transform 1 0 1328 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5729_6
timestamp 1731220534
transform 1 0 1280 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5728_6
timestamp 1731220534
transform 1 0 1224 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5727_6
timestamp 1731220534
transform 1 0 1240 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5726_6
timestamp 1731220534
transform 1 0 1312 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5725_6
timestamp 1731220534
transform 1 0 1312 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5724_6
timestamp 1731220534
transform 1 0 1240 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5723_6
timestamp 1731220534
transform 1 0 1272 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5722_6
timestamp 1731220534
transform 1 0 1256 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5721_6
timestamp 1731220534
transform 1 0 1560 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5720_6
timestamp 1731220534
transform 1 0 1480 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5719_6
timestamp 1731220534
transform 1 0 1408 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5718_6
timestamp 1731220534
transform 1 0 1344 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5717_6
timestamp 1731220534
transform 1 0 1288 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5716_6
timestamp 1731220534
transform 1 0 1248 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5715_6
timestamp 1731220534
transform 1 0 1472 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5714_6
timestamp 1731220534
transform 1 0 1392 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5713_6
timestamp 1731220534
transform 1 0 1320 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5712_6
timestamp 1731220534
transform 1 0 1256 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5711_6
timestamp 1731220534
transform 1 0 1200 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5710_6
timestamp 1731220534
transform 1 0 1152 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5709_6
timestamp 1731220534
transform 1 0 1208 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5708_6
timestamp 1731220534
transform 1 0 1176 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5707_6
timestamp 1731220534
transform 1 0 1144 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5706_6
timestamp 1731220534
transform 1 0 1104 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5705_6
timestamp 1731220534
transform 1 0 1056 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5704_6
timestamp 1731220534
transform 1 0 1000 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5703_6
timestamp 1731220534
transform 1 0 1008 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5702_6
timestamp 1731220534
transform 1 0 1064 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5701_6
timestamp 1731220534
transform 1 0 1112 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5700_6
timestamp 1731220534
transform 1 0 1288 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5699_6
timestamp 1731220534
transform 1 0 1224 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5698_6
timestamp 1731220534
transform 1 0 1160 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5697_6
timestamp 1731220534
transform 1 0 1096 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5696_6
timestamp 1731220534
transform 1 0 1024 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5695_6
timestamp 1731220534
transform 1 0 960 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5694_6
timestamp 1731220534
transform 1 0 1232 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5693_6
timestamp 1731220534
transform 1 0 1168 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5692_6
timestamp 1731220534
transform 1 0 1096 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5691_6
timestamp 1731220534
transform 1 0 1024 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5690_6
timestamp 1731220534
transform 1 0 952 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5689_6
timestamp 1731220534
transform 1 0 880 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5688_6
timestamp 1731220534
transform 1 0 1144 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5687_6
timestamp 1731220534
transform 1 0 1080 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5686_6
timestamp 1731220534
transform 1 0 1016 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5685_6
timestamp 1731220534
transform 1 0 952 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5684_6
timestamp 1731220534
transform 1 0 880 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5683_6
timestamp 1731220534
transform 1 0 816 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5682_6
timestamp 1731220534
transform 1 0 1072 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5681_6
timestamp 1731220534
transform 1 0 1016 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5680_6
timestamp 1731220534
transform 1 0 952 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5679_6
timestamp 1731220534
transform 1 0 888 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5678_6
timestamp 1731220534
transform 1 0 824 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5677_6
timestamp 1731220534
transform 1 0 768 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5676_6
timestamp 1731220534
transform 1 0 760 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5675_6
timestamp 1731220534
transform 1 0 712 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5674_6
timestamp 1731220534
transform 1 0 712 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5673_6
timestamp 1731220534
transform 1 0 656 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5672_6
timestamp 1731220534
transform 1 0 808 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5671_6
timestamp 1731220534
transform 1 0 864 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5670_6
timestamp 1731220534
transform 1 0 1032 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5669_6
timestamp 1731220534
transform 1 0 976 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5668_6
timestamp 1731220534
transform 1 0 920 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5667_6
timestamp 1731220534
transform 1 0 880 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5666_6
timestamp 1731220534
transform 1 0 816 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5665_6
timestamp 1731220534
transform 1 0 760 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5664_6
timestamp 1731220534
transform 1 0 944 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5663_6
timestamp 1731220534
transform 1 0 1072 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5662_6
timestamp 1731220534
transform 1 0 1008 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5661_6
timestamp 1731220534
transform 1 0 960 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5660_6
timestamp 1731220534
transform 1 0 896 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5659_6
timestamp 1731220534
transform 1 0 832 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5658_6
timestamp 1731220534
transform 1 0 1152 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5657_6
timestamp 1731220534
transform 1 0 1088 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5656_6
timestamp 1731220534
transform 1 0 1024 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5655_6
timestamp 1731220534
transform 1 0 1016 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5654_6
timestamp 1731220534
transform 1 0 960 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5653_6
timestamp 1731220534
transform 1 0 904 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5652_6
timestamp 1731220534
transform 1 0 1080 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5651_6
timestamp 1731220534
transform 1 0 1272 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5650_6
timestamp 1731220534
transform 1 0 1208 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5649_6
timestamp 1731220534
transform 1 0 1144 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5648_6
timestamp 1731220534
transform 1 0 1104 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5647_6
timestamp 1731220534
transform 1 0 1032 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5646_6
timestamp 1731220534
transform 1 0 960 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5645_6
timestamp 1731220534
transform 1 0 1168 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5644_6
timestamp 1731220534
transform 1 0 1232 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5643_6
timestamp 1731220534
transform 1 0 1296 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5642_6
timestamp 1731220534
transform 1 0 1272 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5641_6
timestamp 1731220534
transform 1 0 1216 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5640_6
timestamp 1731220534
transform 1 0 1152 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5639_6
timestamp 1731220534
transform 1 0 1088 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5638_6
timestamp 1731220534
transform 1 0 1024 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5637_6
timestamp 1731220534
transform 1 0 952 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5636_6
timestamp 1731220534
transform 1 0 1216 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5635_6
timestamp 1731220534
transform 1 0 1152 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5634_6
timestamp 1731220534
transform 1 0 1088 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5633_6
timestamp 1731220534
transform 1 0 1024 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5632_6
timestamp 1731220534
transform 1 0 960 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5631_6
timestamp 1731220534
transform 1 0 896 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5630_6
timestamp 1731220534
transform 1 0 1160 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5629_6
timestamp 1731220534
transform 1 0 1096 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5628_6
timestamp 1731220534
transform 1 0 1032 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5627_6
timestamp 1731220534
transform 1 0 968 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5626_6
timestamp 1731220534
transform 1 0 904 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5625_6
timestamp 1731220534
transform 1 0 840 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5624_6
timestamp 1731220534
transform 1 0 1080 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5623_6
timestamp 1731220534
transform 1 0 1016 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5622_6
timestamp 1731220534
transform 1 0 952 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5621_6
timestamp 1731220534
transform 1 0 896 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5620_6
timestamp 1731220534
transform 1 0 840 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5619_6
timestamp 1731220534
transform 1 0 792 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5618_6
timestamp 1731220534
transform 1 0 792 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5617_6
timestamp 1731220534
transform 1 0 840 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5616_6
timestamp 1731220534
transform 1 0 896 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5615_6
timestamp 1731220534
transform 1 0 960 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5614_6
timestamp 1731220534
transform 1 0 1096 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5613_6
timestamp 1731220534
transform 1 0 1032 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5612_6
timestamp 1731220534
transform 1 0 1032 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5611_6
timestamp 1731220534
transform 1 0 968 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5610_6
timestamp 1731220534
transform 1 0 904 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5609_6
timestamp 1731220534
transform 1 0 1104 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5608_6
timestamp 1731220534
transform 1 0 1176 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5607_6
timestamp 1731220534
transform 1 0 1240 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5606_6
timestamp 1731220534
transform 1 0 1288 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5605_6
timestamp 1731220534
transform 1 0 1224 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5604_6
timestamp 1731220534
transform 1 0 1160 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5603_6
timestamp 1731220534
transform 1 0 1088 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5602_6
timestamp 1731220534
transform 1 0 1016 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5601_6
timestamp 1731220534
transform 1 0 944 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5600_6
timestamp 1731220534
transform 1 0 1176 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5599_6
timestamp 1731220534
transform 1 0 1112 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5598_6
timestamp 1731220534
transform 1 0 1048 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5597_6
timestamp 1731220534
transform 1 0 984 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5596_6
timestamp 1731220534
transform 1 0 920 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5595_6
timestamp 1731220534
transform 1 0 952 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5594_6
timestamp 1731220534
transform 1 0 1080 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5593_6
timestamp 1731220534
transform 1 0 1016 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5592_6
timestamp 1731220534
transform 1 0 968 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5591_6
timestamp 1731220534
transform 1 0 1040 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5590_6
timestamp 1731220534
transform 1 0 1120 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5589_6
timestamp 1731220534
transform 1 0 1120 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5588_6
timestamp 1731220534
transform 1 0 1040 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5587_6
timestamp 1731220534
transform 1 0 1096 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5586_6
timestamp 1731220534
transform 1 0 1040 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5585_6
timestamp 1731220534
transform 1 0 984 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5584_6
timestamp 1731220534
transform 1 0 1000 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5583_6
timestamp 1731220534
transform 1 0 936 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5582_6
timestamp 1731220534
transform 1 0 872 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5581_6
timestamp 1731220534
transform 1 0 872 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5580_6
timestamp 1731220534
transform 1 0 816 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5579_6
timestamp 1731220534
transform 1 0 928 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5578_6
timestamp 1731220534
transform 1 0 960 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5577_6
timestamp 1731220534
transform 1 0 888 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5576_6
timestamp 1731220534
transform 1 0 824 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5575_6
timestamp 1731220534
transform 1 0 784 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5574_6
timestamp 1731220534
transform 1 0 840 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5573_6
timestamp 1731220534
transform 1 0 904 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5572_6
timestamp 1731220534
transform 1 0 880 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5571_6
timestamp 1731220534
transform 1 0 816 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5570_6
timestamp 1731220534
transform 1 0 752 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5569_6
timestamp 1731220534
transform 1 0 728 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5568_6
timestamp 1731220534
transform 1 0 792 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5567_6
timestamp 1731220534
transform 1 0 856 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5566_6
timestamp 1731220534
transform 1 0 864 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5565_6
timestamp 1731220534
transform 1 0 784 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5564_6
timestamp 1731220534
transform 1 0 696 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5563_6
timestamp 1731220534
transform 1 0 840 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5562_6
timestamp 1731220534
transform 1 0 784 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5561_6
timestamp 1731220534
transform 1 0 728 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5560_6
timestamp 1731220534
transform 1 0 664 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5559_6
timestamp 1731220534
transform 1 0 744 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5558_6
timestamp 1731220534
transform 1 0 696 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5557_6
timestamp 1731220534
transform 1 0 528 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5556_6
timestamp 1731220534
transform 1 0 464 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5555_6
timestamp 1731220534
transform 1 0 464 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5554_6
timestamp 1731220534
transform 1 0 528 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5553_6
timestamp 1731220534
transform 1 0 584 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5552_6
timestamp 1731220534
transform 1 0 656 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5551_6
timestamp 1731220534
transform 1 0 592 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5550_6
timestamp 1731220534
transform 1 0 528 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5549_6
timestamp 1731220534
transform 1 0 464 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5548_6
timestamp 1731220534
transform 1 0 680 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5547_6
timestamp 1731220534
transform 1 0 608 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5546_6
timestamp 1731220534
transform 1 0 536 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5545_6
timestamp 1731220534
transform 1 0 472 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5544_6
timestamp 1731220534
transform 1 0 704 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5543_6
timestamp 1731220534
transform 1 0 624 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5542_6
timestamp 1731220534
transform 1 0 552 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5541_6
timestamp 1731220534
transform 1 0 496 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5540_6
timestamp 1731220534
transform 1 0 648 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5539_6
timestamp 1731220534
transform 1 0 568 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5538_6
timestamp 1731220534
transform 1 0 496 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5537_6
timestamp 1731220534
transform 1 0 432 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5536_6
timestamp 1731220534
transform 1 0 384 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5535_6
timestamp 1731220534
transform 1 0 344 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5534_6
timestamp 1731220534
transform 1 0 304 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5533_6
timestamp 1731220534
transform 1 0 448 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5532_6
timestamp 1731220534
transform 1 0 416 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5531_6
timestamp 1731220534
transform 1 0 384 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5530_6
timestamp 1731220534
transform 1 0 352 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5529_6
timestamp 1731220534
transform 1 0 320 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5528_6
timestamp 1731220534
transform 1 0 288 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5527_6
timestamp 1731220534
transform 1 0 416 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5526_6
timestamp 1731220534
transform 1 0 376 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5525_6
timestamp 1731220534
transform 1 0 336 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5524_6
timestamp 1731220534
transform 1 0 304 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5523_6
timestamp 1731220534
transform 1 0 272 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5522_6
timestamp 1731220534
transform 1 0 240 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5521_6
timestamp 1731220534
transform 1 0 400 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5520_6
timestamp 1731220534
transform 1 0 336 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5519_6
timestamp 1731220534
transform 1 0 280 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5518_6
timestamp 1731220534
transform 1 0 232 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5517_6
timestamp 1731220534
transform 1 0 192 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5516_6
timestamp 1731220534
transform 1 0 160 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5515_6
timestamp 1731220534
transform 1 0 400 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5514_6
timestamp 1731220534
transform 1 0 328 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5513_6
timestamp 1731220534
transform 1 0 264 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5512_6
timestamp 1731220534
transform 1 0 200 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5511_6
timestamp 1731220534
transform 1 0 160 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5510_6
timestamp 1731220534
transform 1 0 128 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5509_6
timestamp 1731220534
transform 1 0 400 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5508_6
timestamp 1731220534
transform 1 0 328 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5507_6
timestamp 1731220534
transform 1 0 264 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5506_6
timestamp 1731220534
transform 1 0 200 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5505_6
timestamp 1731220534
transform 1 0 160 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5504_6
timestamp 1731220534
transform 1 0 128 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5503_6
timestamp 1731220534
transform 1 0 128 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5502_6
timestamp 1731220534
transform 1 0 160 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5501_6
timestamp 1731220534
transform 1 0 208 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5500_6
timestamp 1731220534
transform 1 0 408 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5499_6
timestamp 1731220534
transform 1 0 336 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5498_6
timestamp 1731220534
transform 1 0 272 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5497_6
timestamp 1731220534
transform 1 0 224 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5496_6
timestamp 1731220534
transform 1 0 168 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5495_6
timestamp 1731220534
transform 1 0 128 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5494_6
timestamp 1731220534
transform 1 0 440 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5493_6
timestamp 1731220534
transform 1 0 360 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5492_6
timestamp 1731220534
transform 1 0 288 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5491_6
timestamp 1731220534
transform 1 0 272 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5490_6
timestamp 1731220534
transform 1 0 240 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5489_6
timestamp 1731220534
transform 1 0 208 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5488_6
timestamp 1731220534
transform 1 0 312 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5487_6
timestamp 1731220534
transform 1 0 392 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5486_6
timestamp 1731220534
transform 1 0 352 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5485_6
timestamp 1731220534
transform 1 0 336 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5484_6
timestamp 1731220534
transform 1 0 304 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5483_6
timestamp 1731220534
transform 1 0 272 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5482_6
timestamp 1731220534
transform 1 0 368 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5481_6
timestamp 1731220534
transform 1 0 400 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5480_6
timestamp 1731220534
transform 1 0 432 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5479_6
timestamp 1731220534
transform 1 0 480 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5478_6
timestamp 1731220534
transform 1 0 448 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5477_6
timestamp 1731220534
transform 1 0 416 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5476_6
timestamp 1731220534
transform 1 0 384 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5475_6
timestamp 1731220534
transform 1 0 352 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5474_6
timestamp 1731220534
transform 1 0 320 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5473_6
timestamp 1731220534
transform 1 0 288 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5472_6
timestamp 1731220534
transform 1 0 464 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5471_6
timestamp 1731220534
transform 1 0 416 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5470_6
timestamp 1731220534
transform 1 0 360 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5469_6
timestamp 1731220534
transform 1 0 312 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5468_6
timestamp 1731220534
transform 1 0 272 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5467_6
timestamp 1731220534
transform 1 0 240 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5466_6
timestamp 1731220534
transform 1 0 480 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5465_6
timestamp 1731220534
transform 1 0 400 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5464_6
timestamp 1731220534
transform 1 0 328 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5463_6
timestamp 1731220534
transform 1 0 264 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5462_6
timestamp 1731220534
transform 1 0 208 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5461_6
timestamp 1731220534
transform 1 0 160 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5460_6
timestamp 1731220534
transform 1 0 320 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5459_6
timestamp 1731220534
transform 1 0 272 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5458_6
timestamp 1731220534
transform 1 0 224 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5457_6
timestamp 1731220534
transform 1 0 192 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5456_6
timestamp 1731220534
transform 1 0 160 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5455_6
timestamp 1731220534
transform 1 0 128 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5454_6
timestamp 1731220534
transform 1 0 232 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5453_6
timestamp 1731220534
transform 1 0 192 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5452_6
timestamp 1731220534
transform 1 0 160 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5451_6
timestamp 1731220534
transform 1 0 128 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5450_6
timestamp 1731220534
transform 1 0 280 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5449_6
timestamp 1731220534
transform 1 0 248 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5448_6
timestamp 1731220534
transform 1 0 200 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5447_6
timestamp 1731220534
transform 1 0 144 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5446_6
timestamp 1731220534
transform 1 0 168 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5445_6
timestamp 1731220534
transform 1 0 216 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5444_6
timestamp 1731220534
transform 1 0 192 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5443_6
timestamp 1731220534
transform 1 0 160 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5442_6
timestamp 1731220534
transform 1 0 128 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5441_6
timestamp 1731220534
transform 1 0 160 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5440_6
timestamp 1731220534
transform 1 0 128 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5439_6
timestamp 1731220534
transform 1 0 128 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5438_6
timestamp 1731220534
transform 1 0 160 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5437_6
timestamp 1731220534
transform 1 0 224 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5436_6
timestamp 1731220534
transform 1 0 168 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5435_6
timestamp 1731220534
transform 1 0 128 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5434_6
timestamp 1731220534
transform 1 0 128 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5433_6
timestamp 1731220534
transform 1 0 160 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5432_6
timestamp 1731220534
transform 1 0 200 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5431_6
timestamp 1731220534
transform 1 0 224 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5430_6
timestamp 1731220534
transform 1 0 168 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5429_6
timestamp 1731220534
transform 1 0 128 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5428_6
timestamp 1731220534
transform 1 0 128 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5427_6
timestamp 1731220534
transform 1 0 160 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5426_6
timestamp 1731220534
transform 1 0 192 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5425_6
timestamp 1731220534
transform 1 0 224 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5424_6
timestamp 1731220534
transform 1 0 256 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5423_6
timestamp 1731220534
transform 1 0 288 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5422_6
timestamp 1731220534
transform 1 0 320 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5421_6
timestamp 1731220534
transform 1 0 352 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5420_6
timestamp 1731220534
transform 1 0 384 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5419_6
timestamp 1731220534
transform 1 0 416 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5418_6
timestamp 1731220534
transform 1 0 392 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5417_6
timestamp 1731220534
transform 1 0 336 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5416_6
timestamp 1731220534
transform 1 0 280 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5415_6
timestamp 1731220534
transform 1 0 248 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5414_6
timestamp 1731220534
transform 1 0 296 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5413_6
timestamp 1731220534
transform 1 0 336 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5412_6
timestamp 1731220534
transform 1 0 440 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5411_6
timestamp 1731220534
transform 1 0 376 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5410_6
timestamp 1731220534
transform 1 0 312 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5409_6
timestamp 1731220534
transform 1 0 240 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5408_6
timestamp 1731220534
transform 1 0 288 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5407_6
timestamp 1731220534
transform 1 0 360 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5406_6
timestamp 1731220534
transform 1 0 432 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5405_6
timestamp 1731220534
transform 1 0 384 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5404_6
timestamp 1731220534
transform 1 0 320 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5403_6
timestamp 1731220534
transform 1 0 256 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5402_6
timestamp 1731220534
transform 1 0 200 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5401_6
timestamp 1731220534
transform 1 0 232 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5400_6
timestamp 1731220534
transform 1 0 288 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5399_6
timestamp 1731220534
transform 1 0 344 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5398_6
timestamp 1731220534
transform 1 0 400 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5397_6
timestamp 1731220534
transform 1 0 408 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5396_6
timestamp 1731220534
transform 1 0 360 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5395_6
timestamp 1731220534
transform 1 0 312 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5394_6
timestamp 1731220534
transform 1 0 264 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5393_6
timestamp 1731220534
transform 1 0 304 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5392_6
timestamp 1731220534
transform 1 0 432 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5391_6
timestamp 1731220534
transform 1 0 360 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5390_6
timestamp 1731220534
transform 1 0 320 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5389_6
timestamp 1731220534
transform 1 0 368 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5388_6
timestamp 1731220534
transform 1 0 416 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5387_6
timestamp 1731220534
transform 1 0 472 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5386_6
timestamp 1731220534
transform 1 0 424 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5385_6
timestamp 1731220534
transform 1 0 368 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5384_6
timestamp 1731220534
transform 1 0 488 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5383_6
timestamp 1731220534
transform 1 0 552 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5382_6
timestamp 1731220534
transform 1 0 616 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5381_6
timestamp 1731220534
transform 1 0 608 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5380_6
timestamp 1731220534
transform 1 0 536 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5379_6
timestamp 1731220534
transform 1 0 688 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5378_6
timestamp 1731220534
transform 1 0 672 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5377_6
timestamp 1731220534
transform 1 0 592 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5376_6
timestamp 1731220534
transform 1 0 512 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5375_6
timestamp 1731220534
transform 1 0 464 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5374_6
timestamp 1731220534
transform 1 0 520 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5373_6
timestamp 1731220534
transform 1 0 584 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5372_6
timestamp 1731220534
transform 1 0 656 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5371_6
timestamp 1731220534
transform 1 0 624 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5370_6
timestamp 1731220534
transform 1 0 568 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5369_6
timestamp 1731220534
transform 1 0 512 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5368_6
timestamp 1731220534
transform 1 0 456 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5367_6
timestamp 1731220534
transform 1 0 448 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5366_6
timestamp 1731220534
transform 1 0 512 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5365_6
timestamp 1731220534
transform 1 0 680 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5364_6
timestamp 1731220534
transform 1 0 744 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5363_6
timestamp 1731220534
transform 1 0 680 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5362_6
timestamp 1731220534
transform 1 0 624 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5361_6
timestamp 1731220534
transform 1 0 656 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5360_6
timestamp 1731220534
transform 1 0 736 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5359_6
timestamp 1731220534
transform 1 0 816 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5358_6
timestamp 1731220534
transform 1 0 888 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5357_6
timestamp 1731220534
transform 1 0 1024 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5356_6
timestamp 1731220534
transform 1 0 944 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5355_6
timestamp 1731220534
transform 1 0 872 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5354_6
timestamp 1731220534
transform 1 0 800 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5353_6
timestamp 1731220534
transform 1 0 736 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5352_6
timestamp 1731220534
transform 1 0 808 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5351_6
timestamp 1731220534
transform 1 0 872 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5350_6
timestamp 1731220534
transform 1 0 944 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5349_6
timestamp 1731220534
transform 1 0 1024 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5348_6
timestamp 1731220534
transform 1 0 1032 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5347_6
timestamp 1731220534
transform 1 0 976 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5346_6
timestamp 1731220534
transform 1 0 912 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5345_6
timestamp 1731220534
transform 1 0 848 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5344_6
timestamp 1731220534
transform 1 0 864 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5343_6
timestamp 1731220534
transform 1 0 984 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5342_6
timestamp 1731220534
transform 1 0 928 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5341_6
timestamp 1731220534
transform 1 0 904 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5340_6
timestamp 1731220534
transform 1 0 832 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5339_6
timestamp 1731220534
transform 1 0 976 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5338_6
timestamp 1731220534
transform 1 0 1048 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5337_6
timestamp 1731220534
transform 1 0 1120 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5336_6
timestamp 1731220534
transform 1 0 1192 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5335_6
timestamp 1731220534
transform 1 0 1120 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5334_6
timestamp 1731220534
transform 1 0 1080 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5333_6
timestamp 1731220534
transform 1 0 1032 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5332_6
timestamp 1731220534
transform 1 0 1088 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5331_6
timestamp 1731220534
transform 1 0 1144 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5330_6
timestamp 1731220534
transform 1 0 1104 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5329_6
timestamp 1731220534
transform 1 0 1184 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5328_6
timestamp 1731220534
transform 1 0 1264 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5327_6
timestamp 1731220534
transform 1 0 1256 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5326_6
timestamp 1731220534
transform 1 0 1184 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5325_6
timestamp 1731220534
transform 1 0 1104 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5324_6
timestamp 1731220534
transform 1 0 1248 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5323_6
timestamp 1731220534
transform 1 0 1192 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5322_6
timestamp 1731220534
transform 1 0 1136 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5321_6
timestamp 1731220534
transform 1 0 1080 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5320_6
timestamp 1731220534
transform 1 0 1024 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5319_6
timestamp 1731220534
transform 1 0 960 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5318_6
timestamp 1731220534
transform 1 0 1208 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5317_6
timestamp 1731220534
transform 1 0 1136 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5316_6
timestamp 1731220534
transform 1 0 1064 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5315_6
timestamp 1731220534
transform 1 0 992 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5314_6
timestamp 1731220534
transform 1 0 920 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5313_6
timestamp 1731220534
transform 1 0 848 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5312_6
timestamp 1731220534
transform 1 0 1136 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5311_6
timestamp 1731220534
transform 1 0 1072 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5310_6
timestamp 1731220534
transform 1 0 1008 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5309_6
timestamp 1731220534
transform 1 0 944 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5308_6
timestamp 1731220534
transform 1 0 888 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5307_6
timestamp 1731220534
transform 1 0 824 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5306_6
timestamp 1731220534
transform 1 0 1136 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5305_6
timestamp 1731220534
transform 1 0 1096 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5304_6
timestamp 1731220534
transform 1 0 1056 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5303_6
timestamp 1731220534
transform 1 0 1008 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5302_6
timestamp 1731220534
transform 1 0 968 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5301_6
timestamp 1731220534
transform 1 0 928 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5300_6
timestamp 1731220534
transform 1 0 888 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5299_6
timestamp 1731220534
transform 1 0 856 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5298_6
timestamp 1731220534
transform 1 0 824 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5297_6
timestamp 1731220534
transform 1 0 792 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5296_6
timestamp 1731220534
transform 1 0 760 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5295_6
timestamp 1731220534
transform 1 0 728 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5294_6
timestamp 1731220534
transform 1 0 696 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5293_6
timestamp 1731220534
transform 1 0 664 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5292_6
timestamp 1731220534
transform 1 0 632 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5291_6
timestamp 1731220534
transform 1 0 600 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5290_6
timestamp 1731220534
transform 1 0 568 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5289_6
timestamp 1731220534
transform 1 0 536 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5288_6
timestamp 1731220534
transform 1 0 496 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5287_6
timestamp 1731220534
transform 1 0 456 0 1 80
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5286_6
timestamp 1731220534
transform 1 0 760 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5285_6
timestamp 1731220534
transform 1 0 696 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5284_6
timestamp 1731220534
transform 1 0 632 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5283_6
timestamp 1731220534
transform 1 0 568 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5282_6
timestamp 1731220534
transform 1 0 504 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5281_6
timestamp 1731220534
transform 1 0 448 0 -1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5280_6
timestamp 1731220534
transform 1 0 768 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5279_6
timestamp 1731220534
transform 1 0 688 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5278_6
timestamp 1731220534
transform 1 0 608 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5277_6
timestamp 1731220534
transform 1 0 464 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5276_6
timestamp 1731220534
transform 1 0 408 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5275_6
timestamp 1731220534
transform 1 0 368 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5274_6
timestamp 1731220534
transform 1 0 528 0 1 176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5273_6
timestamp 1731220534
transform 1 0 584 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5272_6
timestamp 1731220534
transform 1 0 512 0 -1 256
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5271_6
timestamp 1731220534
transform 1 0 496 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5270_6
timestamp 1731220534
transform 1 0 560 0 1 260
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5269_6
timestamp 1731220534
transform 1 0 568 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5268_6
timestamp 1731220534
transform 1 0 624 0 -1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5267_6
timestamp 1731220534
transform 1 0 680 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5266_6
timestamp 1731220534
transform 1 0 792 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5265_6
timestamp 1731220534
transform 1 0 736 0 1 340
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5264_6
timestamp 1731220534
transform 1 0 728 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5263_6
timestamp 1731220534
transform 1 0 800 0 -1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5262_6
timestamp 1731220534
transform 1 0 752 0 1 424
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5261_6
timestamp 1731220534
transform 1 0 840 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5260_6
timestamp 1731220534
transform 1 0 768 0 -1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5259_6
timestamp 1731220534
transform 1 0 744 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5258_6
timestamp 1731220534
transform 1 0 680 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5257_6
timestamp 1731220534
transform 1 0 808 0 1 504
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5256_6
timestamp 1731220534
transform 1 0 760 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5255_6
timestamp 1731220534
transform 1 0 696 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5254_6
timestamp 1731220534
transform 1 0 624 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5253_6
timestamp 1731220534
transform 1 0 552 0 -1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5252_6
timestamp 1731220534
transform 1 0 768 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5251_6
timestamp 1731220534
transform 1 0 712 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5250_6
timestamp 1731220534
transform 1 0 656 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5249_6
timestamp 1731220534
transform 1 0 608 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5248_6
timestamp 1731220534
transform 1 0 560 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5247_6
timestamp 1731220534
transform 1 0 512 0 1 588
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5246_6
timestamp 1731220534
transform 1 0 728 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5245_6
timestamp 1731220534
transform 1 0 680 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5244_6
timestamp 1731220534
transform 1 0 632 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5243_6
timestamp 1731220534
transform 1 0 584 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5242_6
timestamp 1731220534
transform 1 0 544 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5241_6
timestamp 1731220534
transform 1 0 512 0 -1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5240_6
timestamp 1731220534
transform 1 0 696 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5239_6
timestamp 1731220534
transform 1 0 640 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5238_6
timestamp 1731220534
transform 1 0 584 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5237_6
timestamp 1731220534
transform 1 0 536 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5236_6
timestamp 1731220534
transform 1 0 496 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5235_6
timestamp 1731220534
transform 1 0 464 0 1 668
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5234_6
timestamp 1731220534
transform 1 0 432 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5233_6
timestamp 1731220534
transform 1 0 480 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5232_6
timestamp 1731220534
transform 1 0 536 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5231_6
timestamp 1731220534
transform 1 0 600 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5230_6
timestamp 1731220534
transform 1 0 664 0 -1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5229_6
timestamp 1731220534
transform 1 0 608 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5228_6
timestamp 1731220534
transform 1 0 520 0 1 752
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5227_6
timestamp 1731220534
transform 1 0 472 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5226_6
timestamp 1731220534
transform 1 0 536 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5225_6
timestamp 1731220534
transform 1 0 600 0 -1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5224_6
timestamp 1731220534
transform 1 0 592 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5223_6
timestamp 1731220534
transform 1 0 648 0 1 836
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5222_6
timestamp 1731220534
transform 1 0 640 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5221_6
timestamp 1731220534
transform 1 0 696 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5220_6
timestamp 1731220534
transform 1 0 744 0 -1 920
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5219_6
timestamp 1731220534
transform 1 0 720 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5218_6
timestamp 1731220534
transform 1 0 784 0 1 924
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5217_6
timestamp 1731220534
transform 1 0 752 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5216_6
timestamp 1731220534
transform 1 0 824 0 -1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5215_6
timestamp 1731220534
transform 1 0 872 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5214_6
timestamp 1731220534
transform 1 0 792 0 1 1004
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5213_6
timestamp 1731220534
transform 1 0 728 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5212_6
timestamp 1731220534
transform 1 0 808 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5211_6
timestamp 1731220534
transform 1 0 888 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5210_6
timestamp 1731220534
transform 1 0 848 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5209_6
timestamp 1731220534
transform 1 0 784 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5208_6
timestamp 1731220534
transform 1 0 720 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5207_6
timestamp 1731220534
transform 1 0 656 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5206_6
timestamp 1731220534
transform 1 0 592 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5205_6
timestamp 1731220534
transform 1 0 520 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5204_6
timestamp 1731220534
transform 1 0 776 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5203_6
timestamp 1731220534
transform 1 0 720 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5202_6
timestamp 1731220534
transform 1 0 656 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5201_6
timestamp 1731220534
transform 1 0 592 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5200_6
timestamp 1731220534
transform 1 0 528 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5199_6
timestamp 1731220534
transform 1 0 464 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5198_6
timestamp 1731220534
transform 1 0 704 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5197_6
timestamp 1731220534
transform 1 0 648 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5196_6
timestamp 1731220534
transform 1 0 592 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5195_6
timestamp 1731220534
transform 1 0 536 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5194_6
timestamp 1731220534
transform 1 0 480 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5193_6
timestamp 1731220534
transform 1 0 424 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5192_6
timestamp 1731220534
transform 1 0 600 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5191_6
timestamp 1731220534
transform 1 0 544 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5190_6
timestamp 1731220534
transform 1 0 488 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5189_6
timestamp 1731220534
transform 1 0 432 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5188_6
timestamp 1731220534
transform 1 0 424 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5187_6
timestamp 1731220534
transform 1 0 480 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5186_6
timestamp 1731220534
transform 1 0 536 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5185_6
timestamp 1731220534
transform 1 0 656 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5184_6
timestamp 1731220534
transform 1 0 600 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5183_6
timestamp 1731220534
transform 1 0 560 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5182_6
timestamp 1731220534
transform 1 0 504 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5181_6
timestamp 1731220534
transform 1 0 448 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5180_6
timestamp 1731220534
transform 1 0 624 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5179_6
timestamp 1731220534
transform 1 0 752 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5178_6
timestamp 1731220534
transform 1 0 688 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5177_6
timestamp 1731220534
transform 1 0 656 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5176_6
timestamp 1731220534
transform 1 0 576 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5175_6
timestamp 1731220534
transform 1 0 496 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5174_6
timestamp 1731220534
transform 1 0 808 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5173_6
timestamp 1731220534
transform 1 0 736 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5172_6
timestamp 1731220534
transform 1 0 672 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5171_6
timestamp 1731220534
transform 1 0 592 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5170_6
timestamp 1731220534
transform 1 0 512 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5169_6
timestamp 1731220534
transform 1 0 752 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5168_6
timestamp 1731220534
transform 1 0 824 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5167_6
timestamp 1731220534
transform 1 0 896 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5166_6
timestamp 1731220534
transform 1 0 840 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5165_6
timestamp 1731220534
transform 1 0 896 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5164_6
timestamp 1731220534
transform 1 0 952 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5163_6
timestamp 1731220534
transform 1 0 936 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5162_6
timestamp 1731220534
transform 1 0 912 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5161_6
timestamp 1731220534
transform 1 0 1000 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5160_6
timestamp 1731220534
transform 1 0 1088 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5159_6
timestamp 1731220534
transform 1 0 1176 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5158_6
timestamp 1731220534
transform 1 0 1192 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5157_6
timestamp 1731220534
transform 1 0 1112 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5156_6
timestamp 1731220534
transform 1 0 1032 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5155_6
timestamp 1731220534
transform 1 0 944 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5154_6
timestamp 1731220534
transform 1 0 1016 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5153_6
timestamp 1731220534
transform 1 0 1096 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5152_6
timestamp 1731220534
transform 1 0 1168 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5151_6
timestamp 1731220534
transform 1 0 1096 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5150_6
timestamp 1731220534
transform 1 0 1024 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5149_6
timestamp 1731220534
transform 1 0 1168 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5148_6
timestamp 1731220534
transform 1 0 1168 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5147_6
timestamp 1731220534
transform 1 0 1112 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5146_6
timestamp 1731220534
transform 1 0 1056 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5145_6
timestamp 1731220534
transform 1 0 1000 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5144_6
timestamp 1731220534
transform 1 0 944 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5143_6
timestamp 1731220534
transform 1 0 888 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5142_6
timestamp 1731220534
transform 1 0 832 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5141_6
timestamp 1731220534
transform 1 0 864 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5140_6
timestamp 1731220534
transform 1 0 944 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5139_6
timestamp 1731220534
transform 1 0 936 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5138_6
timestamp 1731220534
transform 1 0 864 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5137_6
timestamp 1731220534
transform 1 0 792 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5136_6
timestamp 1731220534
transform 1 0 792 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5135_6
timestamp 1731220534
transform 1 0 864 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5134_6
timestamp 1731220534
transform 1 0 824 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5133_6
timestamp 1731220534
transform 1 0 872 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5132_6
timestamp 1731220534
transform 1 0 808 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5131_6
timestamp 1731220534
transform 1 0 736 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5130_6
timestamp 1731220534
transform 1 0 776 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5129_6
timestamp 1731220534
transform 1 0 712 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5128_6
timestamp 1731220534
transform 1 0 656 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5127_6
timestamp 1731220534
transform 1 0 592 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5126_6
timestamp 1731220534
transform 1 0 520 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5125_6
timestamp 1731220534
transform 1 0 520 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5124_6
timestamp 1731220534
transform 1 0 592 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5123_6
timestamp 1731220534
transform 1 0 664 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5122_6
timestamp 1731220534
transform 1 0 752 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5121_6
timestamp 1731220534
transform 1 0 688 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5120_6
timestamp 1731220534
transform 1 0 624 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5119_6
timestamp 1731220534
transform 1 0 656 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5118_6
timestamp 1731220534
transform 1 0 720 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5117_6
timestamp 1731220534
transform 1 0 720 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5116_6
timestamp 1731220534
transform 1 0 656 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5115_6
timestamp 1731220534
transform 1 0 624 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5114_6
timestamp 1731220534
transform 1 0 704 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5113_6
timestamp 1731220534
transform 1 0 784 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5112_6
timestamp 1731220534
transform 1 0 776 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5111_6
timestamp 1731220534
transform 1 0 720 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5110_6
timestamp 1731220534
transform 1 0 656 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5109_6
timestamp 1731220534
transform 1 0 600 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5108_6
timestamp 1731220534
transform 1 0 544 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5107_6
timestamp 1731220534
transform 1 0 496 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5106_6
timestamp 1731220534
transform 1 0 480 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5105_6
timestamp 1731220534
transform 1 0 408 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5104_6
timestamp 1731220534
transform 1 0 552 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5103_6
timestamp 1731220534
transform 1 0 592 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5102_6
timestamp 1731220534
transform 1 0 528 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5101_6
timestamp 1731220534
transform 1 0 464 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_5100_6
timestamp 1731220534
transform 1 0 472 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_599_6
timestamp 1731220534
transform 1 0 528 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_598_6
timestamp 1731220534
transform 1 0 592 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_597_6
timestamp 1731220534
transform 1 0 560 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_596_6
timestamp 1731220534
transform 1 0 504 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_595_6
timestamp 1731220534
transform 1 0 448 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_594_6
timestamp 1731220534
transform 1 0 400 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_593_6
timestamp 1731220534
transform 1 0 352 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_592_6
timestamp 1731220534
transform 1 0 328 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_591_6
timestamp 1731220534
transform 1 0 376 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_590_6
timestamp 1731220534
transform 1 0 424 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_589_6
timestamp 1731220534
transform 1 0 408 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_588_6
timestamp 1731220534
transform 1 0 352 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_587_6
timestamp 1731220534
transform 1 0 296 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_586_6
timestamp 1731220534
transform 1 0 240 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_585_6
timestamp 1731220534
transform 1 0 176 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_584_6
timestamp 1731220534
transform 1 0 272 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_583_6
timestamp 1731220534
transform 1 0 216 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_582_6
timestamp 1731220534
transform 1 0 208 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_581_6
timestamp 1731220534
transform 1 0 256 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_580_6
timestamp 1731220534
transform 1 0 304 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_579_6
timestamp 1731220534
transform 1 0 448 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_578_6
timestamp 1731220534
transform 1 0 368 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_577_6
timestamp 1731220534
transform 1 0 288 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_576_6
timestamp 1731220534
transform 1 0 216 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_575_6
timestamp 1731220534
transform 1 0 160 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_574_6
timestamp 1731220534
transform 1 0 216 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_573_6
timestamp 1731220534
transform 1 0 288 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_572_6
timestamp 1731220534
transform 1 0 368 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_571_6
timestamp 1731220534
transform 1 0 448 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_570_6
timestamp 1731220534
transform 1 0 432 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_569_6
timestamp 1731220534
transform 1 0 352 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_568_6
timestamp 1731220534
transform 1 0 280 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_567_6
timestamp 1731220534
transform 1 0 216 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_566_6
timestamp 1731220534
transform 1 0 280 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_565_6
timestamp 1731220534
transform 1 0 352 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_564_6
timestamp 1731220534
transform 1 0 424 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_563_6
timestamp 1731220534
transform 1 0 392 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_562_6
timestamp 1731220534
transform 1 0 344 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_561_6
timestamp 1731220534
transform 1 0 288 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_560_6
timestamp 1731220534
transform 1 0 232 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_559_6
timestamp 1731220534
transform 1 0 368 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_558_6
timestamp 1731220534
transform 1 0 320 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_557_6
timestamp 1731220534
transform 1 0 272 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_556_6
timestamp 1731220534
transform 1 0 272 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_555_6
timestamp 1731220534
transform 1 0 320 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_554_6
timestamp 1731220534
transform 1 0 376 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_553_6
timestamp 1731220534
transform 1 0 376 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_552_6
timestamp 1731220534
transform 1 0 328 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_551_6
timestamp 1731220534
transform 1 0 272 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_550_6
timestamp 1731220534
transform 1 0 280 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_549_6
timestamp 1731220534
transform 1 0 344 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_548_6
timestamp 1731220534
transform 1 0 408 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_547_6
timestamp 1731220534
transform 1 0 456 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_546_6
timestamp 1731220534
transform 1 0 392 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_545_6
timestamp 1731220534
transform 1 0 328 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_544_6
timestamp 1731220534
transform 1 0 272 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_543_6
timestamp 1731220534
transform 1 0 240 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_542_6
timestamp 1731220534
transform 1 0 208 0 -1 1088
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_541_6
timestamp 1731220534
transform 1 0 264 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_540_6
timestamp 1731220534
transform 1 0 208 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_539_6
timestamp 1731220534
transform 1 0 168 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_538_6
timestamp 1731220534
transform 1 0 136 0 1 1092
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_537_6
timestamp 1731220534
transform 1 0 128 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_536_6
timestamp 1731220534
transform 1 0 160 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_535_6
timestamp 1731220534
transform 1 0 216 0 -1 1176
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_534_6
timestamp 1731220534
transform 1 0 216 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_533_6
timestamp 1731220534
transform 1 0 160 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_532_6
timestamp 1731220534
transform 1 0 128 0 1 1180
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_531_6
timestamp 1731220534
transform 1 0 128 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_530_6
timestamp 1731220534
transform 1 0 160 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_529_6
timestamp 1731220534
transform 1 0 216 0 -1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_528_6
timestamp 1731220534
transform 1 0 224 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_527_6
timestamp 1731220534
transform 1 0 176 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_526_6
timestamp 1731220534
transform 1 0 128 0 1 1264
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_525_6
timestamp 1731220534
transform 1 0 128 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_524_6
timestamp 1731220534
transform 1 0 176 0 -1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_523_6
timestamp 1731220534
transform 1 0 160 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_522_6
timestamp 1731220534
transform 1 0 128 0 1 1348
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_521_6
timestamp 1731220534
transform 1 0 208 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_520_6
timestamp 1731220534
transform 1 0 160 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_519_6
timestamp 1731220534
transform 1 0 128 0 -1 1428
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_518_6
timestamp 1731220534
transform 1 0 128 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_517_6
timestamp 1731220534
transform 1 0 160 0 1 1432
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_516_6
timestamp 1731220534
transform 1 0 128 0 -1 1512
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_515_6
timestamp 1731220534
transform 1 0 128 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_514_6
timestamp 1731220534
transform 1 0 160 0 1 1516
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_513_6
timestamp 1731220534
transform 1 0 160 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_512_6
timestamp 1731220534
transform 1 0 128 0 -1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_511_6
timestamp 1731220534
transform 1 0 128 0 1 1596
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_510_6
timestamp 1731220534
transform 1 0 128 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_59_6
timestamp 1731220534
transform 1 0 160 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_58_6
timestamp 1731220534
transform 1 0 208 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_57_6
timestamp 1731220534
transform 1 0 272 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_56_6
timestamp 1731220534
transform 1 0 336 0 -1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_55_6
timestamp 1731220534
transform 1 0 312 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_54_6
timestamp 1731220534
transform 1 0 280 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_53_6
timestamp 1731220534
transform 1 0 248 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_52_6
timestamp 1731220534
transform 1 0 352 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_51_6
timestamp 1731220534
transform 1 0 400 0 1 1676
box 8 7 28 34
use _0_0std_0_0cells_0_0INVX1  tst_50_6
timestamp 1731220534
transform 1 0 448 0 1 1676
box 8 7 28 34
<< end >>
