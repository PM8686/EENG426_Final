VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.600000 BY 0.300000 ;
END CoreSite

LAYER li
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.056250 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.225000 ;
   PITCH 0.600000 0.600000 ;
END li

LAYER mcon
    TYPE CUT ;
    SPACING 0.225000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END mcon

LAYER met1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.150000 ;
   AREA 0.084375 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met1

LAYER v1
    TYPE CUT ;
    SPACING 0.075000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.075000 ;
END v1

LAYER met2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.150000 ;
   AREA 0.073125 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met2

LAYER v2
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v2

LAYER met3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met3

LAYER v3
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.450000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v3

LAYER met4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met4

LAYER v4
    TYPE CUT ;
    SPACING 0.450000 ;
    WIDTH 1.200000 ;
    ENCLOSURE ABOVE 0.150000 0.150000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END v4

LAYER met5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.650000 ;
   AREA 4.005000 ;
   WIDTH 1.650000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 1.650000 ;
   PITCH 3.300000 3.300000 ;
END met5

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA mcon_C DEFAULT
   LAYER li ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER mcon ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END mcon_C

VIA v1_C DEFAULT
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER met2 ;
     RECT -0.225000 -0.150000 0.225000 0.150000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_C

VIA v3_Ch
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Ch

VIA v3_Cv
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER met4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER met5 ;
     RECT -0.750000 -0.750000 0.750000 0.750000 ;
END v4_C

MACRO _0_0cell_0_0gcelem2x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0gcelem2x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 6.600000 BY 4.800000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 4.350000 0.900000 4.425000 1.125000 ;
        RECT 4.425000 0.900000 4.650000 1.125000 ;
        RECT 4.650000 0.900000 4.725000 1.125000 ;
        RECT 4.500000 0.600000 4.725000 0.900000 ;
        RECT 4.500000 0.300000 4.800000 0.600000 ;
        END
        ANTENNAGATEAREA 0.247500 ;
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.750000 3.900000 3.825000 4.125000 ;
        RECT 3.825000 3.900000 4.050000 4.125000 ;
        RECT 4.050000 3.900000 4.425000 4.125000 ;
        RECT 4.200000 4.200000 4.500000 4.500000 ;
        RECT 4.200000 4.125000 4.425000 4.200000 ;
        END
        ANTENNAGATEAREA 0.247500 ;
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 3.675000 1.800000 3.900000 2.025000 ;
        RECT 3.675000 1.725000 3.900000 1.800000 ;
        RECT 3.675000 2.925000 3.900000 3.000000 ;
        RECT 3.675000 2.700000 3.900000 2.925000 ;
        RECT 3.675000 2.475000 3.900000 2.700000 ;
        RECT 3.675000 2.250000 3.900000 2.475000 ;
        RECT 3.675000 2.025000 3.900000 2.250000 ;
        RECT 6.000000 2.700000 6.300000 3.000000 ;
        RECT 6.000000 2.400000 6.225000 2.700000 ;
        RECT 6.000000 2.175000 6.225000 2.400000 ;
        RECT 6.000000 2.100000 6.225000 2.175000 ;
        LAYER mcon ;
        RECT 3.675000 2.250000 3.900000 2.475000 ;
        RECT 6.000000 2.175000 6.225000 2.400000 ;
        LAYER met1 ;
        RECT 5.925000 2.175000 6.000000 2.250000 ;
        RECT 5.925000 2.100000 6.300000 2.175000 ;
        RECT 6.000000 2.175000 6.225000 2.400000 ;
        RECT 6.225000 2.175000 6.300000 2.400000 ;
        RECT 3.600000 2.475000 3.975000 2.550000 ;
        RECT 3.600000 2.250000 3.675000 2.475000 ;
        RECT 3.600000 2.175000 3.975000 2.250000 ;
        RECT 3.675000 2.250000 3.900000 2.475000 ;
        RECT 3.900000 2.400000 3.975000 2.475000 ;
        RECT 3.900000 2.250000 6.000000 2.400000 ;
        RECT 5.925000 2.400000 6.300000 2.475000 ;
        END
        ANTENNAGATEAREA 0.360000 ;
        ANTENNADIFFAREA 0.697500 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.675000 3.000000 0.900000 3.075000 ;
        RECT 0.675000 2.775000 0.900000 3.000000 ;
        RECT 0.675000 2.700000 0.900000 2.775000 ;
        RECT 1.575000 1.425000 1.800000 2.775000 ;
        RECT 1.575000 1.200000 1.800000 1.425000 ;
        RECT 1.575000 1.125000 1.800000 1.200000 ;
        RECT 1.575000 3.000000 1.800000 3.075000 ;
        RECT 1.575000 2.775000 1.800000 3.000000 ;
        RECT 4.575000 3.000000 4.800000 3.075000 ;
        RECT 4.575000 2.775000 4.800000 3.000000 ;
        RECT 4.575000 2.700000 4.800000 2.775000 ;
        LAYER mcon ;
        RECT 0.675000 2.775000 0.900000 3.000000 ;
        RECT 1.575000 2.775000 1.800000 3.000000 ;
        RECT 4.575000 2.775000 4.800000 3.000000 ;
        LAYER met1 ;
        RECT 0.600000 3.000000 4.875000 3.075000 ;
        RECT 0.600000 2.775000 0.675000 3.000000 ;
        RECT 0.600000 2.700000 4.875000 2.775000 ;
        RECT 0.675000 2.775000 0.900000 3.000000 ;
        RECT 0.900000 2.775000 1.575000 3.000000 ;
        RECT 1.575000 2.775000 1.800000 3.000000 ;
        RECT 1.800000 2.775000 4.575000 3.000000 ;
        RECT 4.575000 2.775000 4.800000 3.000000 ;
        RECT 4.800000 2.775000 4.875000 3.000000 ;
        END
        ANTENNAGATEAREA 0.945000 ;
        ANTENNADIFFAREA 0.495000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.675000 1.950000 0.900000 2.025000 ;
        RECT 0.675000 1.725000 0.900000 1.950000 ;
        RECT 0.675000 1.650000 0.900000 1.725000 ;
        RECT 1.125000 3.600000 1.350000 3.675000 ;
        RECT 1.125000 3.375000 1.350000 3.600000 ;
        RECT 1.125000 1.950000 1.350000 3.375000 ;
        RECT 1.125000 1.725000 1.350000 1.950000 ;
        RECT 1.125000 1.650000 1.350000 1.725000 ;
        RECT 4.500000 1.725000 4.575000 1.950000 ;
        RECT 4.575000 1.725000 4.800000 1.950000 ;
        RECT 4.800000 1.725000 4.875000 1.950000 ;
        LAYER mcon ;
        RECT 0.675000 1.725000 0.900000 1.950000 ;
        RECT 1.125000 1.725000 1.350000 1.950000 ;
        RECT 4.575000 1.725000 4.800000 1.950000 ;
        LAYER met1 ;
        RECT 0.600000 1.950000 4.875000 2.025000 ;
        RECT 0.600000 1.725000 0.675000 1.950000 ;
        RECT 0.600000 1.650000 4.875000 1.725000 ;
        RECT 0.675000 1.725000 0.900000 1.950000 ;
        RECT 0.900000 1.725000 1.125000 1.950000 ;
        RECT 1.125000 1.725000 1.350000 1.950000 ;
        RECT 1.350000 1.725000 4.575000 1.950000 ;
        RECT 4.575000 1.725000 4.800000 1.950000 ;
        RECT 4.800000 1.725000 4.875000 1.950000 ;
        END
        ANTENNAGATEAREA 0.472500 ;
        ANTENNADIFFAREA 0.427500 ;
    END GND
    OBS
        LAYER li ;
        RECT 3.150000 3.600000 3.375000 3.675000 ;
        RECT 3.150000 3.375000 3.375000 3.600000 ;
        RECT 3.150000 3.300000 3.375000 3.375000 ;
        RECT 5.250000 3.600000 5.475000 3.675000 ;
        RECT 5.250000 3.375000 5.475000 3.600000 ;
        RECT 5.250000 2.925000 5.475000 3.375000 ;
        RECT 5.250000 2.700000 5.475000 2.925000 ;
        RECT 5.250000 2.025000 5.475000 2.700000 ;
        RECT 5.250000 1.800000 5.475000 2.025000 ;
        RECT 5.250000 1.725000 5.475000 1.800000 ;
        LAYER met1 ;
        RECT 3.075000 3.600000 5.550000 3.675000 ;
        RECT 3.075000 3.375000 3.150000 3.600000 ;
        RECT 3.075000 3.300000 5.550000 3.375000 ;
        RECT 3.150000 3.375000 3.375000 3.600000 ;
        RECT 3.375000 3.375000 5.250000 3.600000 ;
        RECT 5.250000 3.375000 5.475000 3.600000 ;
        RECT 5.475000 3.375000 5.550000 3.600000 ;
    END
END _0_0cell_0_0gcelem2x0

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 2.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.525000 1.725000 0.900000 1.800000 ;
        RECT 0.525000 1.500000 0.600000 1.725000 ;
        RECT 0.525000 1.425000 0.900000 1.500000 ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        RECT 0.825000 1.500000 0.900000 1.725000 ;
        LAYER mcon ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        LAYER met1 ;
        RECT 0.525000 1.725000 0.900000 1.800000 ;
        RECT 0.525000 1.500000 0.600000 1.725000 ;
        RECT 0.525000 1.425000 0.900000 1.500000 ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        RECT 0.825000 1.500000 0.900000 1.725000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.525000 0.525000 0.900000 0.600000 ;
        RECT 0.525000 0.300000 0.600000 0.525000 ;
        RECT 0.525000 0.225000 0.900000 0.300000 ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        RECT 0.825000 0.300000 0.900000 0.525000 ;
        LAYER mcon ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        LAYER met1 ;
        RECT 0.525000 0.525000 0.900000 0.600000 ;
        RECT 0.525000 0.300000 0.600000 0.525000 ;
        RECT 0.525000 0.225000 0.900000 0.300000 ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        RECT 0.825000 0.300000 0.900000 0.525000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 258.000000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 258.000000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

