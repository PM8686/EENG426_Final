magic
tech sky130l
timestamp 1731220652
<< m2 >>
rect 718 2557 724 2558
rect 110 2556 116 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 718 2553 719 2557
rect 723 2553 724 2557
rect 718 2552 724 2553
rect 774 2557 780 2558
rect 774 2553 775 2557
rect 779 2553 780 2557
rect 774 2552 780 2553
rect 830 2557 836 2558
rect 830 2553 831 2557
rect 835 2553 836 2557
rect 830 2552 836 2553
rect 886 2557 892 2558
rect 886 2553 887 2557
rect 891 2553 892 2557
rect 886 2552 892 2553
rect 942 2557 948 2558
rect 942 2553 943 2557
rect 947 2553 948 2557
rect 942 2552 948 2553
rect 1286 2556 1292 2557
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 110 2551 116 2552
rect 1286 2551 1292 2552
rect 110 2539 116 2540
rect 110 2535 111 2539
rect 115 2535 116 2539
rect 1286 2539 1292 2540
rect 110 2534 116 2535
rect 702 2536 708 2537
rect 702 2532 703 2536
rect 707 2532 708 2536
rect 702 2531 708 2532
rect 758 2536 764 2537
rect 758 2532 759 2536
rect 763 2532 764 2536
rect 758 2531 764 2532
rect 814 2536 820 2537
rect 814 2532 815 2536
rect 819 2532 820 2536
rect 814 2531 820 2532
rect 870 2536 876 2537
rect 870 2532 871 2536
rect 875 2532 876 2536
rect 870 2531 876 2532
rect 926 2536 932 2537
rect 926 2532 927 2536
rect 931 2532 932 2536
rect 1286 2535 1287 2539
rect 1291 2535 1292 2539
rect 1286 2534 1292 2535
rect 1398 2533 1404 2534
rect 926 2531 932 2532
rect 1326 2532 1332 2533
rect 1326 2528 1327 2532
rect 1331 2528 1332 2532
rect 1398 2529 1399 2533
rect 1403 2529 1404 2533
rect 1398 2528 1404 2529
rect 1454 2533 1460 2534
rect 1454 2529 1455 2533
rect 1459 2529 1460 2533
rect 1454 2528 1460 2529
rect 1510 2533 1516 2534
rect 1510 2529 1511 2533
rect 1515 2529 1516 2533
rect 1510 2528 1516 2529
rect 1566 2533 1572 2534
rect 1566 2529 1567 2533
rect 1571 2529 1572 2533
rect 1566 2528 1572 2529
rect 1622 2533 1628 2534
rect 1622 2529 1623 2533
rect 1627 2529 1628 2533
rect 1622 2528 1628 2529
rect 1678 2533 1684 2534
rect 1678 2529 1679 2533
rect 1683 2529 1684 2533
rect 1678 2528 1684 2529
rect 1734 2533 1740 2534
rect 1734 2529 1735 2533
rect 1739 2529 1740 2533
rect 1734 2528 1740 2529
rect 1790 2533 1796 2534
rect 1790 2529 1791 2533
rect 1795 2529 1796 2533
rect 1790 2528 1796 2529
rect 1846 2533 1852 2534
rect 1846 2529 1847 2533
rect 1851 2529 1852 2533
rect 1846 2528 1852 2529
rect 1902 2533 1908 2534
rect 1902 2529 1903 2533
rect 1907 2529 1908 2533
rect 1902 2528 1908 2529
rect 1958 2533 1964 2534
rect 1958 2529 1959 2533
rect 1963 2529 1964 2533
rect 1958 2528 1964 2529
rect 2014 2533 2020 2534
rect 2014 2529 2015 2533
rect 2019 2529 2020 2533
rect 2014 2528 2020 2529
rect 2070 2533 2076 2534
rect 2070 2529 2071 2533
rect 2075 2529 2076 2533
rect 2070 2528 2076 2529
rect 2126 2533 2132 2534
rect 2126 2529 2127 2533
rect 2131 2529 2132 2533
rect 2126 2528 2132 2529
rect 2182 2533 2188 2534
rect 2182 2529 2183 2533
rect 2187 2529 2188 2533
rect 2182 2528 2188 2529
rect 2502 2532 2508 2533
rect 2502 2528 2503 2532
rect 2507 2528 2508 2532
rect 1326 2527 1332 2528
rect 2502 2527 2508 2528
rect 166 2524 172 2525
rect 110 2521 116 2522
rect 110 2517 111 2521
rect 115 2517 116 2521
rect 166 2520 167 2524
rect 171 2520 172 2524
rect 166 2519 172 2520
rect 222 2524 228 2525
rect 222 2520 223 2524
rect 227 2520 228 2524
rect 222 2519 228 2520
rect 278 2524 284 2525
rect 278 2520 279 2524
rect 283 2520 284 2524
rect 278 2519 284 2520
rect 342 2524 348 2525
rect 342 2520 343 2524
rect 347 2520 348 2524
rect 342 2519 348 2520
rect 406 2524 412 2525
rect 406 2520 407 2524
rect 411 2520 412 2524
rect 406 2519 412 2520
rect 478 2524 484 2525
rect 478 2520 479 2524
rect 483 2520 484 2524
rect 478 2519 484 2520
rect 558 2524 564 2525
rect 558 2520 559 2524
rect 563 2520 564 2524
rect 558 2519 564 2520
rect 638 2524 644 2525
rect 638 2520 639 2524
rect 643 2520 644 2524
rect 638 2519 644 2520
rect 718 2524 724 2525
rect 718 2520 719 2524
rect 723 2520 724 2524
rect 718 2519 724 2520
rect 798 2524 804 2525
rect 798 2520 799 2524
rect 803 2520 804 2524
rect 798 2519 804 2520
rect 878 2524 884 2525
rect 878 2520 879 2524
rect 883 2520 884 2524
rect 878 2519 884 2520
rect 958 2524 964 2525
rect 958 2520 959 2524
rect 963 2520 964 2524
rect 958 2519 964 2520
rect 1038 2524 1044 2525
rect 1038 2520 1039 2524
rect 1043 2520 1044 2524
rect 1038 2519 1044 2520
rect 1286 2521 1292 2522
rect 110 2516 116 2517
rect 1286 2517 1287 2521
rect 1291 2517 1292 2521
rect 1286 2516 1292 2517
rect 1326 2515 1332 2516
rect 1326 2511 1327 2515
rect 1331 2511 1332 2515
rect 2502 2515 2508 2516
rect 1326 2510 1332 2511
rect 1382 2512 1388 2513
rect 1382 2508 1383 2512
rect 1387 2508 1388 2512
rect 1382 2507 1388 2508
rect 1438 2512 1444 2513
rect 1438 2508 1439 2512
rect 1443 2508 1444 2512
rect 1438 2507 1444 2508
rect 1494 2512 1500 2513
rect 1494 2508 1495 2512
rect 1499 2508 1500 2512
rect 1494 2507 1500 2508
rect 1550 2512 1556 2513
rect 1550 2508 1551 2512
rect 1555 2508 1556 2512
rect 1550 2507 1556 2508
rect 1606 2512 1612 2513
rect 1606 2508 1607 2512
rect 1611 2508 1612 2512
rect 1606 2507 1612 2508
rect 1662 2512 1668 2513
rect 1662 2508 1663 2512
rect 1667 2508 1668 2512
rect 1662 2507 1668 2508
rect 1718 2512 1724 2513
rect 1718 2508 1719 2512
rect 1723 2508 1724 2512
rect 1718 2507 1724 2508
rect 1774 2512 1780 2513
rect 1774 2508 1775 2512
rect 1779 2508 1780 2512
rect 1774 2507 1780 2508
rect 1830 2512 1836 2513
rect 1830 2508 1831 2512
rect 1835 2508 1836 2512
rect 1830 2507 1836 2508
rect 1886 2512 1892 2513
rect 1886 2508 1887 2512
rect 1891 2508 1892 2512
rect 1886 2507 1892 2508
rect 1942 2512 1948 2513
rect 1942 2508 1943 2512
rect 1947 2508 1948 2512
rect 1942 2507 1948 2508
rect 1998 2512 2004 2513
rect 1998 2508 1999 2512
rect 2003 2508 2004 2512
rect 1998 2507 2004 2508
rect 2054 2512 2060 2513
rect 2054 2508 2055 2512
rect 2059 2508 2060 2512
rect 2054 2507 2060 2508
rect 2110 2512 2116 2513
rect 2110 2508 2111 2512
rect 2115 2508 2116 2512
rect 2110 2507 2116 2508
rect 2166 2512 2172 2513
rect 2166 2508 2167 2512
rect 2171 2508 2172 2512
rect 2502 2511 2503 2515
rect 2507 2511 2508 2515
rect 2502 2510 2508 2511
rect 2166 2507 2172 2508
rect 110 2504 116 2505
rect 1286 2504 1292 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 110 2499 116 2500
rect 182 2503 188 2504
rect 182 2499 183 2503
rect 187 2499 188 2503
rect 182 2498 188 2499
rect 238 2503 244 2504
rect 238 2499 239 2503
rect 243 2499 244 2503
rect 238 2498 244 2499
rect 294 2503 300 2504
rect 294 2499 295 2503
rect 299 2499 300 2503
rect 294 2498 300 2499
rect 358 2503 364 2504
rect 358 2499 359 2503
rect 363 2499 364 2503
rect 358 2498 364 2499
rect 422 2503 428 2504
rect 422 2499 423 2503
rect 427 2499 428 2503
rect 422 2498 428 2499
rect 494 2503 500 2504
rect 494 2499 495 2503
rect 499 2499 500 2503
rect 494 2498 500 2499
rect 574 2503 580 2504
rect 574 2499 575 2503
rect 579 2499 580 2503
rect 574 2498 580 2499
rect 654 2503 660 2504
rect 654 2499 655 2503
rect 659 2499 660 2503
rect 654 2498 660 2499
rect 734 2503 740 2504
rect 734 2499 735 2503
rect 739 2499 740 2503
rect 734 2498 740 2499
rect 814 2503 820 2504
rect 814 2499 815 2503
rect 819 2499 820 2503
rect 814 2498 820 2499
rect 894 2503 900 2504
rect 894 2499 895 2503
rect 899 2499 900 2503
rect 894 2498 900 2499
rect 974 2503 980 2504
rect 974 2499 975 2503
rect 979 2499 980 2503
rect 974 2498 980 2499
rect 1054 2503 1060 2504
rect 1054 2499 1055 2503
rect 1059 2499 1060 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1054 2498 1060 2499
rect 1350 2492 1356 2493
rect 1326 2489 1332 2490
rect 1326 2485 1327 2489
rect 1331 2485 1332 2489
rect 1350 2488 1351 2492
rect 1355 2488 1356 2492
rect 1350 2487 1356 2488
rect 1422 2492 1428 2493
rect 1422 2488 1423 2492
rect 1427 2488 1428 2492
rect 1422 2487 1428 2488
rect 1510 2492 1516 2493
rect 1510 2488 1511 2492
rect 1515 2488 1516 2492
rect 1510 2487 1516 2488
rect 1598 2492 1604 2493
rect 1598 2488 1599 2492
rect 1603 2488 1604 2492
rect 1598 2487 1604 2488
rect 1686 2492 1692 2493
rect 1686 2488 1687 2492
rect 1691 2488 1692 2492
rect 1686 2487 1692 2488
rect 1774 2492 1780 2493
rect 1774 2488 1775 2492
rect 1779 2488 1780 2492
rect 1774 2487 1780 2488
rect 1862 2492 1868 2493
rect 1862 2488 1863 2492
rect 1867 2488 1868 2492
rect 1862 2487 1868 2488
rect 1950 2492 1956 2493
rect 1950 2488 1951 2492
rect 1955 2488 1956 2492
rect 1950 2487 1956 2488
rect 2038 2492 2044 2493
rect 2038 2488 2039 2492
rect 2043 2488 2044 2492
rect 2038 2487 2044 2488
rect 2126 2492 2132 2493
rect 2126 2488 2127 2492
rect 2131 2488 2132 2492
rect 2126 2487 2132 2488
rect 2502 2489 2508 2490
rect 1326 2484 1332 2485
rect 2502 2485 2503 2489
rect 2507 2485 2508 2489
rect 2502 2484 2508 2485
rect 1326 2472 1332 2473
rect 2502 2472 2508 2473
rect 1326 2468 1327 2472
rect 1331 2468 1332 2472
rect 1326 2467 1332 2468
rect 1366 2471 1372 2472
rect 1366 2467 1367 2471
rect 1371 2467 1372 2471
rect 1366 2466 1372 2467
rect 1438 2471 1444 2472
rect 1438 2467 1439 2471
rect 1443 2467 1444 2471
rect 1438 2466 1444 2467
rect 1526 2471 1532 2472
rect 1526 2467 1527 2471
rect 1531 2467 1532 2471
rect 1526 2466 1532 2467
rect 1614 2471 1620 2472
rect 1614 2467 1615 2471
rect 1619 2467 1620 2471
rect 1614 2466 1620 2467
rect 1702 2471 1708 2472
rect 1702 2467 1703 2471
rect 1707 2467 1708 2471
rect 1702 2466 1708 2467
rect 1790 2471 1796 2472
rect 1790 2467 1791 2471
rect 1795 2467 1796 2471
rect 1790 2466 1796 2467
rect 1878 2471 1884 2472
rect 1878 2467 1879 2471
rect 1883 2467 1884 2471
rect 1878 2466 1884 2467
rect 1966 2471 1972 2472
rect 1966 2467 1967 2471
rect 1971 2467 1972 2471
rect 1966 2466 1972 2467
rect 2054 2471 2060 2472
rect 2054 2467 2055 2471
rect 2059 2467 2060 2471
rect 2054 2466 2060 2467
rect 2142 2471 2148 2472
rect 2142 2467 2143 2471
rect 2147 2467 2148 2471
rect 2502 2468 2503 2472
rect 2507 2468 2508 2472
rect 2502 2467 2508 2468
rect 2142 2466 2148 2467
rect 182 2453 188 2454
rect 110 2452 116 2453
rect 110 2448 111 2452
rect 115 2448 116 2452
rect 182 2449 183 2453
rect 187 2449 188 2453
rect 182 2448 188 2449
rect 246 2453 252 2454
rect 246 2449 247 2453
rect 251 2449 252 2453
rect 246 2448 252 2449
rect 326 2453 332 2454
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 414 2453 420 2454
rect 414 2449 415 2453
rect 419 2449 420 2453
rect 414 2448 420 2449
rect 502 2453 508 2454
rect 502 2449 503 2453
rect 507 2449 508 2453
rect 502 2448 508 2449
rect 598 2453 604 2454
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 598 2448 604 2449
rect 694 2453 700 2454
rect 694 2449 695 2453
rect 699 2449 700 2453
rect 694 2448 700 2449
rect 790 2453 796 2454
rect 790 2449 791 2453
rect 795 2449 796 2453
rect 790 2448 796 2449
rect 878 2453 884 2454
rect 878 2449 879 2453
rect 883 2449 884 2453
rect 878 2448 884 2449
rect 966 2453 972 2454
rect 966 2449 967 2453
rect 971 2449 972 2453
rect 966 2448 972 2449
rect 1062 2453 1068 2454
rect 1062 2449 1063 2453
rect 1067 2449 1068 2453
rect 1062 2448 1068 2449
rect 1158 2453 1164 2454
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1158 2448 1164 2449
rect 1286 2452 1292 2453
rect 1286 2448 1287 2452
rect 1291 2448 1292 2452
rect 110 2447 116 2448
rect 1286 2447 1292 2448
rect 110 2435 116 2436
rect 110 2431 111 2435
rect 115 2431 116 2435
rect 1286 2435 1292 2436
rect 110 2430 116 2431
rect 166 2432 172 2433
rect 166 2428 167 2432
rect 171 2428 172 2432
rect 166 2427 172 2428
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 486 2432 492 2433
rect 486 2428 487 2432
rect 491 2428 492 2432
rect 486 2427 492 2428
rect 582 2432 588 2433
rect 582 2428 583 2432
rect 587 2428 588 2432
rect 582 2427 588 2428
rect 678 2432 684 2433
rect 678 2428 679 2432
rect 683 2428 684 2432
rect 678 2427 684 2428
rect 774 2432 780 2433
rect 774 2428 775 2432
rect 779 2428 780 2432
rect 774 2427 780 2428
rect 862 2432 868 2433
rect 862 2428 863 2432
rect 867 2428 868 2432
rect 862 2427 868 2428
rect 950 2432 956 2433
rect 950 2428 951 2432
rect 955 2428 956 2432
rect 950 2427 956 2428
rect 1046 2432 1052 2433
rect 1046 2428 1047 2432
rect 1051 2428 1052 2432
rect 1046 2427 1052 2428
rect 1142 2432 1148 2433
rect 1142 2428 1143 2432
rect 1147 2428 1148 2432
rect 1286 2431 1287 2435
rect 1291 2431 1292 2435
rect 1286 2430 1292 2431
rect 1142 2427 1148 2428
rect 150 2416 156 2417
rect 110 2413 116 2414
rect 110 2409 111 2413
rect 115 2409 116 2413
rect 150 2412 151 2416
rect 155 2412 156 2416
rect 150 2411 156 2412
rect 230 2416 236 2417
rect 230 2412 231 2416
rect 235 2412 236 2416
rect 230 2411 236 2412
rect 318 2416 324 2417
rect 318 2412 319 2416
rect 323 2412 324 2416
rect 318 2411 324 2412
rect 414 2416 420 2417
rect 414 2412 415 2416
rect 419 2412 420 2416
rect 414 2411 420 2412
rect 518 2416 524 2417
rect 518 2412 519 2416
rect 523 2412 524 2416
rect 518 2411 524 2412
rect 622 2416 628 2417
rect 622 2412 623 2416
rect 627 2412 628 2416
rect 622 2411 628 2412
rect 726 2416 732 2417
rect 726 2412 727 2416
rect 731 2412 732 2416
rect 726 2411 732 2412
rect 830 2416 836 2417
rect 830 2412 831 2416
rect 835 2412 836 2416
rect 830 2411 836 2412
rect 934 2416 940 2417
rect 934 2412 935 2416
rect 939 2412 940 2416
rect 934 2411 940 2412
rect 1038 2416 1044 2417
rect 1038 2412 1039 2416
rect 1043 2412 1044 2416
rect 1038 2411 1044 2412
rect 1150 2416 1156 2417
rect 1150 2412 1151 2416
rect 1155 2412 1156 2416
rect 1150 2411 1156 2412
rect 1286 2413 1292 2414
rect 1366 2413 1372 2414
rect 110 2408 116 2409
rect 1286 2409 1287 2413
rect 1291 2409 1292 2413
rect 1286 2408 1292 2409
rect 1326 2412 1332 2413
rect 1326 2408 1327 2412
rect 1331 2408 1332 2412
rect 1366 2409 1367 2413
rect 1371 2409 1372 2413
rect 1366 2408 1372 2409
rect 1438 2413 1444 2414
rect 1438 2409 1439 2413
rect 1443 2409 1444 2413
rect 1438 2408 1444 2409
rect 1542 2413 1548 2414
rect 1542 2409 1543 2413
rect 1547 2409 1548 2413
rect 1542 2408 1548 2409
rect 1638 2413 1644 2414
rect 1638 2409 1639 2413
rect 1643 2409 1644 2413
rect 1638 2408 1644 2409
rect 1734 2413 1740 2414
rect 1734 2409 1735 2413
rect 1739 2409 1740 2413
rect 1734 2408 1740 2409
rect 1822 2413 1828 2414
rect 1822 2409 1823 2413
rect 1827 2409 1828 2413
rect 1822 2408 1828 2409
rect 1910 2413 1916 2414
rect 1910 2409 1911 2413
rect 1915 2409 1916 2413
rect 1910 2408 1916 2409
rect 2006 2413 2012 2414
rect 2006 2409 2007 2413
rect 2011 2409 2012 2413
rect 2006 2408 2012 2409
rect 2102 2413 2108 2414
rect 2102 2409 2103 2413
rect 2107 2409 2108 2413
rect 2102 2408 2108 2409
rect 2502 2412 2508 2413
rect 2502 2408 2503 2412
rect 2507 2408 2508 2412
rect 1326 2407 1332 2408
rect 2502 2407 2508 2408
rect 110 2396 116 2397
rect 1286 2396 1292 2397
rect 110 2392 111 2396
rect 115 2392 116 2396
rect 110 2391 116 2392
rect 166 2395 172 2396
rect 166 2391 167 2395
rect 171 2391 172 2395
rect 166 2390 172 2391
rect 246 2395 252 2396
rect 246 2391 247 2395
rect 251 2391 252 2395
rect 246 2390 252 2391
rect 334 2395 340 2396
rect 334 2391 335 2395
rect 339 2391 340 2395
rect 334 2390 340 2391
rect 430 2395 436 2396
rect 430 2391 431 2395
rect 435 2391 436 2395
rect 430 2390 436 2391
rect 534 2395 540 2396
rect 534 2391 535 2395
rect 539 2391 540 2395
rect 534 2390 540 2391
rect 638 2395 644 2396
rect 638 2391 639 2395
rect 643 2391 644 2395
rect 638 2390 644 2391
rect 742 2395 748 2396
rect 742 2391 743 2395
rect 747 2391 748 2395
rect 742 2390 748 2391
rect 846 2395 852 2396
rect 846 2391 847 2395
rect 851 2391 852 2395
rect 846 2390 852 2391
rect 950 2395 956 2396
rect 950 2391 951 2395
rect 955 2391 956 2395
rect 950 2390 956 2391
rect 1054 2395 1060 2396
rect 1054 2391 1055 2395
rect 1059 2391 1060 2395
rect 1054 2390 1060 2391
rect 1166 2395 1172 2396
rect 1166 2391 1167 2395
rect 1171 2391 1172 2395
rect 1286 2392 1287 2396
rect 1291 2392 1292 2396
rect 1286 2391 1292 2392
rect 1326 2395 1332 2396
rect 1326 2391 1327 2395
rect 1331 2391 1332 2395
rect 2502 2395 2508 2396
rect 1166 2390 1172 2391
rect 1326 2390 1332 2391
rect 1350 2392 1356 2393
rect 1350 2388 1351 2392
rect 1355 2388 1356 2392
rect 1350 2387 1356 2388
rect 1422 2392 1428 2393
rect 1422 2388 1423 2392
rect 1427 2388 1428 2392
rect 1422 2387 1428 2388
rect 1526 2392 1532 2393
rect 1526 2388 1527 2392
rect 1531 2388 1532 2392
rect 1526 2387 1532 2388
rect 1622 2392 1628 2393
rect 1622 2388 1623 2392
rect 1627 2388 1628 2392
rect 1622 2387 1628 2388
rect 1718 2392 1724 2393
rect 1718 2388 1719 2392
rect 1723 2388 1724 2392
rect 1718 2387 1724 2388
rect 1806 2392 1812 2393
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1894 2392 1900 2393
rect 1894 2388 1895 2392
rect 1899 2388 1900 2392
rect 1894 2387 1900 2388
rect 1990 2392 1996 2393
rect 1990 2388 1991 2392
rect 1995 2388 1996 2392
rect 1990 2387 1996 2388
rect 2086 2392 2092 2393
rect 2086 2388 2087 2392
rect 2091 2388 2092 2392
rect 2502 2391 2503 2395
rect 2507 2391 2508 2395
rect 2502 2390 2508 2391
rect 2086 2387 2092 2388
rect 1350 2372 1356 2373
rect 1326 2369 1332 2370
rect 1326 2365 1327 2369
rect 1331 2365 1332 2369
rect 1350 2368 1351 2372
rect 1355 2368 1356 2372
rect 1350 2367 1356 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1494 2372 1500 2373
rect 1494 2368 1495 2372
rect 1499 2368 1500 2372
rect 1494 2367 1500 2368
rect 1582 2372 1588 2373
rect 1582 2368 1583 2372
rect 1587 2368 1588 2372
rect 1582 2367 1588 2368
rect 1670 2372 1676 2373
rect 1670 2368 1671 2372
rect 1675 2368 1676 2372
rect 1670 2367 1676 2368
rect 1750 2372 1756 2373
rect 1750 2368 1751 2372
rect 1755 2368 1756 2372
rect 1750 2367 1756 2368
rect 1830 2372 1836 2373
rect 1830 2368 1831 2372
rect 1835 2368 1836 2372
rect 1830 2367 1836 2368
rect 1918 2372 1924 2373
rect 1918 2368 1919 2372
rect 1923 2368 1924 2372
rect 1918 2367 1924 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2094 2372 2100 2373
rect 2094 2368 2095 2372
rect 2099 2368 2100 2372
rect 2094 2367 2100 2368
rect 2502 2369 2508 2370
rect 1326 2364 1332 2365
rect 2502 2365 2503 2369
rect 2507 2365 2508 2369
rect 2502 2364 2508 2365
rect 1326 2352 1332 2353
rect 2502 2352 2508 2353
rect 1326 2348 1327 2352
rect 1331 2348 1332 2352
rect 1326 2347 1332 2348
rect 1366 2351 1372 2352
rect 1366 2347 1367 2351
rect 1371 2347 1372 2351
rect 1366 2346 1372 2347
rect 1422 2351 1428 2352
rect 1422 2347 1423 2351
rect 1427 2347 1428 2351
rect 1422 2346 1428 2347
rect 1510 2351 1516 2352
rect 1510 2347 1511 2351
rect 1515 2347 1516 2351
rect 1510 2346 1516 2347
rect 1598 2351 1604 2352
rect 1598 2347 1599 2351
rect 1603 2347 1604 2351
rect 1598 2346 1604 2347
rect 1686 2351 1692 2352
rect 1686 2347 1687 2351
rect 1691 2347 1692 2351
rect 1686 2346 1692 2347
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2347 1772 2351
rect 1766 2346 1772 2347
rect 1846 2351 1852 2352
rect 1846 2347 1847 2351
rect 1851 2347 1852 2351
rect 1846 2346 1852 2347
rect 1934 2351 1940 2352
rect 1934 2347 1935 2351
rect 1939 2347 1940 2351
rect 1934 2346 1940 2347
rect 2022 2351 2028 2352
rect 2022 2347 2023 2351
rect 2027 2347 2028 2351
rect 2022 2346 2028 2347
rect 2110 2351 2116 2352
rect 2110 2347 2111 2351
rect 2115 2347 2116 2351
rect 2502 2348 2503 2352
rect 2507 2348 2508 2352
rect 2502 2347 2508 2348
rect 2110 2346 2116 2347
rect 174 2345 180 2346
rect 110 2344 116 2345
rect 110 2340 111 2344
rect 115 2340 116 2344
rect 174 2341 175 2345
rect 179 2341 180 2345
rect 174 2340 180 2341
rect 278 2345 284 2346
rect 278 2341 279 2345
rect 283 2341 284 2345
rect 278 2340 284 2341
rect 390 2345 396 2346
rect 390 2341 391 2345
rect 395 2341 396 2345
rect 390 2340 396 2341
rect 502 2345 508 2346
rect 502 2341 503 2345
rect 507 2341 508 2345
rect 502 2340 508 2341
rect 622 2345 628 2346
rect 622 2341 623 2345
rect 627 2341 628 2345
rect 622 2340 628 2341
rect 742 2345 748 2346
rect 742 2341 743 2345
rect 747 2341 748 2345
rect 742 2340 748 2341
rect 870 2345 876 2346
rect 870 2341 871 2345
rect 875 2341 876 2345
rect 870 2340 876 2341
rect 998 2345 1004 2346
rect 998 2341 999 2345
rect 1003 2341 1004 2345
rect 998 2340 1004 2341
rect 1126 2345 1132 2346
rect 1126 2341 1127 2345
rect 1131 2341 1132 2345
rect 1126 2340 1132 2341
rect 1286 2344 1292 2345
rect 1286 2340 1287 2344
rect 1291 2340 1292 2344
rect 110 2339 116 2340
rect 1286 2339 1292 2340
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 1286 2327 1292 2328
rect 110 2322 116 2323
rect 158 2324 164 2325
rect 158 2320 159 2324
rect 163 2320 164 2324
rect 158 2319 164 2320
rect 262 2324 268 2325
rect 262 2320 263 2324
rect 267 2320 268 2324
rect 262 2319 268 2320
rect 374 2324 380 2325
rect 374 2320 375 2324
rect 379 2320 380 2324
rect 374 2319 380 2320
rect 486 2324 492 2325
rect 486 2320 487 2324
rect 491 2320 492 2324
rect 486 2319 492 2320
rect 606 2324 612 2325
rect 606 2320 607 2324
rect 611 2320 612 2324
rect 606 2319 612 2320
rect 726 2324 732 2325
rect 726 2320 727 2324
rect 731 2320 732 2324
rect 726 2319 732 2320
rect 854 2324 860 2325
rect 854 2320 855 2324
rect 859 2320 860 2324
rect 854 2319 860 2320
rect 982 2324 988 2325
rect 982 2320 983 2324
rect 987 2320 988 2324
rect 982 2319 988 2320
rect 1110 2324 1116 2325
rect 1110 2320 1111 2324
rect 1115 2320 1116 2324
rect 1286 2323 1287 2327
rect 1291 2323 1292 2327
rect 1286 2322 1292 2323
rect 1110 2319 1116 2320
rect 206 2308 212 2309
rect 110 2305 116 2306
rect 110 2301 111 2305
rect 115 2301 116 2305
rect 206 2304 207 2308
rect 211 2304 212 2308
rect 206 2303 212 2304
rect 286 2308 292 2309
rect 286 2304 287 2308
rect 291 2304 292 2308
rect 286 2303 292 2304
rect 374 2308 380 2309
rect 374 2304 375 2308
rect 379 2304 380 2308
rect 374 2303 380 2304
rect 470 2308 476 2309
rect 470 2304 471 2308
rect 475 2304 476 2308
rect 470 2303 476 2304
rect 558 2308 564 2309
rect 558 2304 559 2308
rect 563 2304 564 2308
rect 558 2303 564 2304
rect 646 2308 652 2309
rect 646 2304 647 2308
rect 651 2304 652 2308
rect 646 2303 652 2304
rect 734 2308 740 2309
rect 734 2304 735 2308
rect 739 2304 740 2308
rect 734 2303 740 2304
rect 814 2308 820 2309
rect 814 2304 815 2308
rect 819 2304 820 2308
rect 814 2303 820 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 990 2308 996 2309
rect 990 2304 991 2308
rect 995 2304 996 2308
rect 990 2303 996 2304
rect 1078 2308 1084 2309
rect 1078 2304 1079 2308
rect 1083 2304 1084 2308
rect 1078 2303 1084 2304
rect 1286 2305 1292 2306
rect 110 2300 116 2301
rect 1286 2301 1287 2305
rect 1291 2301 1292 2305
rect 1286 2300 1292 2301
rect 1366 2297 1372 2298
rect 1326 2296 1332 2297
rect 1326 2292 1327 2296
rect 1331 2292 1332 2296
rect 1366 2293 1367 2297
rect 1371 2293 1372 2297
rect 1366 2292 1372 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1542 2297 1548 2298
rect 1542 2293 1543 2297
rect 1547 2293 1548 2297
rect 1542 2292 1548 2293
rect 1638 2297 1644 2298
rect 1638 2293 1639 2297
rect 1643 2293 1644 2297
rect 1638 2292 1644 2293
rect 1734 2297 1740 2298
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1830 2297 1836 2298
rect 1830 2293 1831 2297
rect 1835 2293 1836 2297
rect 1830 2292 1836 2293
rect 1926 2297 1932 2298
rect 1926 2293 1927 2297
rect 1931 2293 1932 2297
rect 1926 2292 1932 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2110 2297 2116 2298
rect 2110 2293 2111 2297
rect 2115 2293 2116 2297
rect 2110 2292 2116 2293
rect 2206 2297 2212 2298
rect 2206 2293 2207 2297
rect 2211 2293 2212 2297
rect 2206 2292 2212 2293
rect 2502 2296 2508 2297
rect 2502 2292 2503 2296
rect 2507 2292 2508 2296
rect 1326 2291 1332 2292
rect 2502 2291 2508 2292
rect 110 2288 116 2289
rect 1286 2288 1292 2289
rect 110 2284 111 2288
rect 115 2284 116 2288
rect 110 2283 116 2284
rect 222 2287 228 2288
rect 222 2283 223 2287
rect 227 2283 228 2287
rect 222 2282 228 2283
rect 302 2287 308 2288
rect 302 2283 303 2287
rect 307 2283 308 2287
rect 302 2282 308 2283
rect 390 2287 396 2288
rect 390 2283 391 2287
rect 395 2283 396 2287
rect 390 2282 396 2283
rect 486 2287 492 2288
rect 486 2283 487 2287
rect 491 2283 492 2287
rect 486 2282 492 2283
rect 574 2287 580 2288
rect 574 2283 575 2287
rect 579 2283 580 2287
rect 574 2282 580 2283
rect 662 2287 668 2288
rect 662 2283 663 2287
rect 667 2283 668 2287
rect 662 2282 668 2283
rect 750 2287 756 2288
rect 750 2283 751 2287
rect 755 2283 756 2287
rect 750 2282 756 2283
rect 830 2287 836 2288
rect 830 2283 831 2287
rect 835 2283 836 2287
rect 830 2282 836 2283
rect 918 2287 924 2288
rect 918 2283 919 2287
rect 923 2283 924 2287
rect 918 2282 924 2283
rect 1006 2287 1012 2288
rect 1006 2283 1007 2287
rect 1011 2283 1012 2287
rect 1006 2282 1012 2283
rect 1094 2287 1100 2288
rect 1094 2283 1095 2287
rect 1099 2283 1100 2287
rect 1286 2284 1287 2288
rect 1291 2284 1292 2288
rect 1286 2283 1292 2284
rect 1094 2282 1100 2283
rect 1326 2279 1332 2280
rect 1326 2275 1327 2279
rect 1331 2275 1332 2279
rect 2502 2279 2508 2280
rect 1326 2274 1332 2275
rect 1350 2276 1356 2277
rect 1350 2272 1351 2276
rect 1355 2272 1356 2276
rect 1350 2271 1356 2272
rect 1438 2276 1444 2277
rect 1438 2272 1439 2276
rect 1443 2272 1444 2276
rect 1438 2271 1444 2272
rect 1526 2276 1532 2277
rect 1526 2272 1527 2276
rect 1531 2272 1532 2276
rect 1526 2271 1532 2272
rect 1622 2276 1628 2277
rect 1622 2272 1623 2276
rect 1627 2272 1628 2276
rect 1622 2271 1628 2272
rect 1718 2276 1724 2277
rect 1718 2272 1719 2276
rect 1723 2272 1724 2276
rect 1718 2271 1724 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1814 2271 1820 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1998 2276 2004 2277
rect 1998 2272 1999 2276
rect 2003 2272 2004 2276
rect 1998 2271 2004 2272
rect 2094 2276 2100 2277
rect 2094 2272 2095 2276
rect 2099 2272 2100 2276
rect 2094 2271 2100 2272
rect 2190 2276 2196 2277
rect 2190 2272 2191 2276
rect 2195 2272 2196 2276
rect 2502 2275 2503 2279
rect 2507 2275 2508 2279
rect 2502 2274 2508 2275
rect 2190 2271 2196 2272
rect 1454 2264 1460 2265
rect 1326 2261 1332 2262
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1454 2260 1455 2264
rect 1459 2260 1460 2264
rect 1454 2259 1460 2260
rect 1542 2264 1548 2265
rect 1542 2260 1543 2264
rect 1547 2260 1548 2264
rect 1542 2259 1548 2260
rect 1638 2264 1644 2265
rect 1638 2260 1639 2264
rect 1643 2260 1644 2264
rect 1638 2259 1644 2260
rect 1734 2264 1740 2265
rect 1734 2260 1735 2264
rect 1739 2260 1740 2264
rect 1734 2259 1740 2260
rect 1838 2264 1844 2265
rect 1838 2260 1839 2264
rect 1843 2260 1844 2264
rect 1838 2259 1844 2260
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 1934 2259 1940 2260
rect 2030 2264 2036 2265
rect 2030 2260 2031 2264
rect 2035 2260 2036 2264
rect 2030 2259 2036 2260
rect 2118 2264 2124 2265
rect 2118 2260 2119 2264
rect 2123 2260 2124 2264
rect 2118 2259 2124 2260
rect 2214 2264 2220 2265
rect 2214 2260 2215 2264
rect 2219 2260 2220 2264
rect 2214 2259 2220 2260
rect 2310 2264 2316 2265
rect 2310 2260 2311 2264
rect 2315 2260 2316 2264
rect 2310 2259 2316 2260
rect 2502 2261 2508 2262
rect 1326 2256 1332 2257
rect 2502 2257 2503 2261
rect 2507 2257 2508 2261
rect 2502 2256 2508 2257
rect 1326 2244 1332 2245
rect 2502 2244 2508 2245
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1326 2239 1332 2240
rect 1470 2243 1476 2244
rect 1470 2239 1471 2243
rect 1475 2239 1476 2243
rect 1470 2238 1476 2239
rect 1558 2243 1564 2244
rect 1558 2239 1559 2243
rect 1563 2239 1564 2243
rect 1558 2238 1564 2239
rect 1654 2243 1660 2244
rect 1654 2239 1655 2243
rect 1659 2239 1660 2243
rect 1654 2238 1660 2239
rect 1750 2243 1756 2244
rect 1750 2239 1751 2243
rect 1755 2239 1756 2243
rect 1750 2238 1756 2239
rect 1854 2243 1860 2244
rect 1854 2239 1855 2243
rect 1859 2239 1860 2243
rect 1854 2238 1860 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 2046 2243 2052 2244
rect 2046 2239 2047 2243
rect 2051 2239 2052 2243
rect 2046 2238 2052 2239
rect 2134 2243 2140 2244
rect 2134 2239 2135 2243
rect 2139 2239 2140 2243
rect 2134 2238 2140 2239
rect 2230 2243 2236 2244
rect 2230 2239 2231 2243
rect 2235 2239 2236 2243
rect 2230 2238 2236 2239
rect 2326 2243 2332 2244
rect 2326 2239 2327 2243
rect 2331 2239 2332 2243
rect 2502 2240 2503 2244
rect 2507 2240 2508 2244
rect 2502 2239 2508 2240
rect 2326 2238 2332 2239
rect 262 2233 268 2234
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 262 2229 263 2233
rect 267 2229 268 2233
rect 262 2228 268 2229
rect 318 2233 324 2234
rect 318 2229 319 2233
rect 323 2229 324 2233
rect 318 2228 324 2229
rect 382 2233 388 2234
rect 382 2229 383 2233
rect 387 2229 388 2233
rect 382 2228 388 2229
rect 446 2233 452 2234
rect 446 2229 447 2233
rect 451 2229 452 2233
rect 446 2228 452 2229
rect 502 2233 508 2234
rect 502 2229 503 2233
rect 507 2229 508 2233
rect 502 2228 508 2229
rect 558 2233 564 2234
rect 558 2229 559 2233
rect 563 2229 564 2233
rect 558 2228 564 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 670 2233 676 2234
rect 670 2229 671 2233
rect 675 2229 676 2233
rect 670 2228 676 2229
rect 726 2233 732 2234
rect 726 2229 727 2233
rect 731 2229 732 2233
rect 726 2228 732 2229
rect 790 2233 796 2234
rect 790 2229 791 2233
rect 795 2229 796 2233
rect 790 2228 796 2229
rect 854 2233 860 2234
rect 854 2229 855 2233
rect 859 2229 860 2233
rect 854 2228 860 2229
rect 918 2233 924 2234
rect 918 2229 919 2233
rect 923 2229 924 2233
rect 918 2228 924 2229
rect 982 2233 988 2234
rect 982 2229 983 2233
rect 987 2229 988 2233
rect 982 2228 988 2229
rect 1046 2233 1052 2234
rect 1046 2229 1047 2233
rect 1051 2229 1052 2233
rect 1046 2228 1052 2229
rect 1110 2233 1116 2234
rect 1110 2229 1111 2233
rect 1115 2229 1116 2233
rect 1110 2228 1116 2229
rect 1286 2232 1292 2233
rect 1286 2228 1287 2232
rect 1291 2228 1292 2232
rect 110 2227 116 2228
rect 1286 2227 1292 2228
rect 110 2215 116 2216
rect 110 2211 111 2215
rect 115 2211 116 2215
rect 1286 2215 1292 2216
rect 110 2210 116 2211
rect 246 2212 252 2213
rect 246 2208 247 2212
rect 251 2208 252 2212
rect 246 2207 252 2208
rect 302 2212 308 2213
rect 302 2208 303 2212
rect 307 2208 308 2212
rect 302 2207 308 2208
rect 366 2212 372 2213
rect 366 2208 367 2212
rect 371 2208 372 2212
rect 366 2207 372 2208
rect 430 2212 436 2213
rect 430 2208 431 2212
rect 435 2208 436 2212
rect 430 2207 436 2208
rect 486 2212 492 2213
rect 486 2208 487 2212
rect 491 2208 492 2212
rect 486 2207 492 2208
rect 542 2212 548 2213
rect 542 2208 543 2212
rect 547 2208 548 2212
rect 542 2207 548 2208
rect 598 2212 604 2213
rect 598 2208 599 2212
rect 603 2208 604 2212
rect 598 2207 604 2208
rect 654 2212 660 2213
rect 654 2208 655 2212
rect 659 2208 660 2212
rect 654 2207 660 2208
rect 710 2212 716 2213
rect 710 2208 711 2212
rect 715 2208 716 2212
rect 710 2207 716 2208
rect 774 2212 780 2213
rect 774 2208 775 2212
rect 779 2208 780 2212
rect 774 2207 780 2208
rect 838 2212 844 2213
rect 838 2208 839 2212
rect 843 2208 844 2212
rect 838 2207 844 2208
rect 902 2212 908 2213
rect 902 2208 903 2212
rect 907 2208 908 2212
rect 902 2207 908 2208
rect 966 2212 972 2213
rect 966 2208 967 2212
rect 971 2208 972 2212
rect 966 2207 972 2208
rect 1030 2212 1036 2213
rect 1030 2208 1031 2212
rect 1035 2208 1036 2212
rect 1030 2207 1036 2208
rect 1094 2212 1100 2213
rect 1094 2208 1095 2212
rect 1099 2208 1100 2212
rect 1286 2211 1287 2215
rect 1291 2211 1292 2215
rect 1286 2210 1292 2211
rect 1094 2207 1100 2208
rect 334 2196 340 2197
rect 110 2193 116 2194
rect 110 2189 111 2193
rect 115 2189 116 2193
rect 334 2192 335 2196
rect 339 2192 340 2196
rect 334 2191 340 2192
rect 390 2196 396 2197
rect 390 2192 391 2196
rect 395 2192 396 2196
rect 390 2191 396 2192
rect 446 2196 452 2197
rect 446 2192 447 2196
rect 451 2192 452 2196
rect 446 2191 452 2192
rect 502 2196 508 2197
rect 502 2192 503 2196
rect 507 2192 508 2196
rect 502 2191 508 2192
rect 558 2196 564 2197
rect 558 2192 559 2196
rect 563 2192 564 2196
rect 558 2191 564 2192
rect 1286 2193 1292 2194
rect 110 2188 116 2189
rect 1286 2189 1287 2193
rect 1291 2189 1292 2193
rect 1566 2189 1572 2190
rect 1286 2188 1292 2189
rect 1326 2188 1332 2189
rect 1326 2184 1327 2188
rect 1331 2184 1332 2188
rect 1566 2185 1567 2189
rect 1571 2185 1572 2189
rect 1566 2184 1572 2185
rect 1622 2189 1628 2190
rect 1622 2185 1623 2189
rect 1627 2185 1628 2189
rect 1622 2184 1628 2185
rect 1678 2189 1684 2190
rect 1678 2185 1679 2189
rect 1683 2185 1684 2189
rect 1678 2184 1684 2185
rect 1742 2189 1748 2190
rect 1742 2185 1743 2189
rect 1747 2185 1748 2189
rect 1742 2184 1748 2185
rect 1806 2189 1812 2190
rect 1806 2185 1807 2189
rect 1811 2185 1812 2189
rect 1806 2184 1812 2185
rect 1870 2189 1876 2190
rect 1870 2185 1871 2189
rect 1875 2185 1876 2189
rect 1870 2184 1876 2185
rect 1926 2189 1932 2190
rect 1926 2185 1927 2189
rect 1931 2185 1932 2189
rect 1926 2184 1932 2185
rect 1982 2189 1988 2190
rect 1982 2185 1983 2189
rect 1987 2185 1988 2189
rect 1982 2184 1988 2185
rect 2038 2189 2044 2190
rect 2038 2185 2039 2189
rect 2043 2185 2044 2189
rect 2038 2184 2044 2185
rect 2094 2189 2100 2190
rect 2094 2185 2095 2189
rect 2099 2185 2100 2189
rect 2094 2184 2100 2185
rect 2158 2189 2164 2190
rect 2158 2185 2159 2189
rect 2163 2185 2164 2189
rect 2158 2184 2164 2185
rect 2222 2189 2228 2190
rect 2222 2185 2223 2189
rect 2227 2185 2228 2189
rect 2222 2184 2228 2185
rect 2286 2189 2292 2190
rect 2286 2185 2287 2189
rect 2291 2185 2292 2189
rect 2286 2184 2292 2185
rect 2342 2189 2348 2190
rect 2342 2185 2343 2189
rect 2347 2185 2348 2189
rect 2342 2184 2348 2185
rect 2398 2189 2404 2190
rect 2398 2185 2399 2189
rect 2403 2185 2404 2189
rect 2398 2184 2404 2185
rect 2454 2189 2460 2190
rect 2454 2185 2455 2189
rect 2459 2185 2460 2189
rect 2454 2184 2460 2185
rect 2502 2188 2508 2189
rect 2502 2184 2503 2188
rect 2507 2184 2508 2188
rect 1326 2183 1332 2184
rect 2502 2183 2508 2184
rect 110 2176 116 2177
rect 1286 2176 1292 2177
rect 110 2172 111 2176
rect 115 2172 116 2176
rect 110 2171 116 2172
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 350 2170 356 2171
rect 406 2175 412 2176
rect 406 2171 407 2175
rect 411 2171 412 2175
rect 406 2170 412 2171
rect 462 2175 468 2176
rect 462 2171 463 2175
rect 467 2171 468 2175
rect 462 2170 468 2171
rect 518 2175 524 2176
rect 518 2171 519 2175
rect 523 2171 524 2175
rect 518 2170 524 2171
rect 574 2175 580 2176
rect 574 2171 575 2175
rect 579 2171 580 2175
rect 1286 2172 1287 2176
rect 1291 2172 1292 2176
rect 1286 2171 1292 2172
rect 1326 2171 1332 2172
rect 574 2170 580 2171
rect 1326 2167 1327 2171
rect 1331 2167 1332 2171
rect 2502 2171 2508 2172
rect 1326 2166 1332 2167
rect 1550 2168 1556 2169
rect 1550 2164 1551 2168
rect 1555 2164 1556 2168
rect 1550 2163 1556 2164
rect 1606 2168 1612 2169
rect 1606 2164 1607 2168
rect 1611 2164 1612 2168
rect 1606 2163 1612 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1726 2168 1732 2169
rect 1726 2164 1727 2168
rect 1731 2164 1732 2168
rect 1726 2163 1732 2164
rect 1790 2168 1796 2169
rect 1790 2164 1791 2168
rect 1795 2164 1796 2168
rect 1790 2163 1796 2164
rect 1854 2168 1860 2169
rect 1854 2164 1855 2168
rect 1859 2164 1860 2168
rect 1854 2163 1860 2164
rect 1910 2168 1916 2169
rect 1910 2164 1911 2168
rect 1915 2164 1916 2168
rect 1910 2163 1916 2164
rect 1966 2168 1972 2169
rect 1966 2164 1967 2168
rect 1971 2164 1972 2168
rect 1966 2163 1972 2164
rect 2022 2168 2028 2169
rect 2022 2164 2023 2168
rect 2027 2164 2028 2168
rect 2022 2163 2028 2164
rect 2078 2168 2084 2169
rect 2078 2164 2079 2168
rect 2083 2164 2084 2168
rect 2078 2163 2084 2164
rect 2142 2168 2148 2169
rect 2142 2164 2143 2168
rect 2147 2164 2148 2168
rect 2142 2163 2148 2164
rect 2206 2168 2212 2169
rect 2206 2164 2207 2168
rect 2211 2164 2212 2168
rect 2206 2163 2212 2164
rect 2270 2168 2276 2169
rect 2270 2164 2271 2168
rect 2275 2164 2276 2168
rect 2270 2163 2276 2164
rect 2326 2168 2332 2169
rect 2326 2164 2327 2168
rect 2331 2164 2332 2168
rect 2326 2163 2332 2164
rect 2382 2168 2388 2169
rect 2382 2164 2383 2168
rect 2387 2164 2388 2168
rect 2382 2163 2388 2164
rect 2438 2168 2444 2169
rect 2438 2164 2439 2168
rect 2443 2164 2444 2168
rect 2502 2167 2503 2171
rect 2507 2167 2508 2171
rect 2502 2166 2508 2167
rect 2438 2163 2444 2164
rect 1662 2144 1668 2145
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1718 2144 1724 2145
rect 1718 2140 1719 2144
rect 1723 2140 1724 2144
rect 1718 2139 1724 2140
rect 1790 2144 1796 2145
rect 1790 2140 1791 2144
rect 1795 2140 1796 2144
rect 1790 2139 1796 2140
rect 1870 2144 1876 2145
rect 1870 2140 1871 2144
rect 1875 2140 1876 2144
rect 1870 2139 1876 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2078 2144 2084 2145
rect 2078 2140 2079 2144
rect 2083 2140 2084 2144
rect 2078 2139 2084 2140
rect 2198 2144 2204 2145
rect 2198 2140 2199 2144
rect 2203 2140 2204 2144
rect 2198 2139 2204 2140
rect 2326 2144 2332 2145
rect 2326 2140 2327 2144
rect 2331 2140 2332 2144
rect 2326 2139 2332 2140
rect 2438 2144 2444 2145
rect 2438 2140 2439 2144
rect 2443 2140 2444 2144
rect 2438 2139 2444 2140
rect 2502 2141 2508 2142
rect 1326 2136 1332 2137
rect 2502 2137 2503 2141
rect 2507 2137 2508 2141
rect 2502 2136 2508 2137
rect 414 2125 420 2126
rect 110 2124 116 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 414 2121 415 2125
rect 419 2121 420 2125
rect 414 2120 420 2121
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 606 2125 612 2126
rect 606 2121 607 2125
rect 611 2121 612 2125
rect 606 2120 612 2121
rect 710 2125 716 2126
rect 710 2121 711 2125
rect 715 2121 716 2125
rect 710 2120 716 2121
rect 814 2125 820 2126
rect 814 2121 815 2125
rect 819 2121 820 2125
rect 814 2120 820 2121
rect 926 2125 932 2126
rect 926 2121 927 2125
rect 931 2121 932 2125
rect 926 2120 932 2121
rect 1038 2125 1044 2126
rect 1038 2121 1039 2125
rect 1043 2121 1044 2125
rect 1038 2120 1044 2121
rect 1150 2125 1156 2126
rect 1150 2121 1151 2125
rect 1155 2121 1156 2125
rect 1150 2120 1156 2121
rect 1238 2125 1244 2126
rect 1238 2121 1239 2125
rect 1243 2121 1244 2125
rect 1238 2120 1244 2121
rect 1286 2124 1292 2125
rect 1286 2120 1287 2124
rect 1291 2120 1292 2124
rect 110 2119 116 2120
rect 1286 2119 1292 2120
rect 1326 2124 1332 2125
rect 2502 2124 2508 2125
rect 1326 2120 1327 2124
rect 1331 2120 1332 2124
rect 1326 2119 1332 2120
rect 1678 2123 1684 2124
rect 1678 2119 1679 2123
rect 1683 2119 1684 2123
rect 1678 2118 1684 2119
rect 1734 2123 1740 2124
rect 1734 2119 1735 2123
rect 1739 2119 1740 2123
rect 1734 2118 1740 2119
rect 1806 2123 1812 2124
rect 1806 2119 1807 2123
rect 1811 2119 1812 2123
rect 1806 2118 1812 2119
rect 1886 2123 1892 2124
rect 1886 2119 1887 2123
rect 1891 2119 1892 2123
rect 1886 2118 1892 2119
rect 1982 2123 1988 2124
rect 1982 2119 1983 2123
rect 1987 2119 1988 2123
rect 1982 2118 1988 2119
rect 2094 2123 2100 2124
rect 2094 2119 2095 2123
rect 2099 2119 2100 2123
rect 2094 2118 2100 2119
rect 2214 2123 2220 2124
rect 2214 2119 2215 2123
rect 2219 2119 2220 2123
rect 2214 2118 2220 2119
rect 2342 2123 2348 2124
rect 2342 2119 2343 2123
rect 2347 2119 2348 2123
rect 2342 2118 2348 2119
rect 2454 2123 2460 2124
rect 2454 2119 2455 2123
rect 2459 2119 2460 2123
rect 2502 2120 2503 2124
rect 2507 2120 2508 2124
rect 2502 2119 2508 2120
rect 2454 2118 2460 2119
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 1286 2107 1292 2108
rect 110 2102 116 2103
rect 398 2104 404 2105
rect 398 2100 399 2104
rect 403 2100 404 2104
rect 398 2099 404 2100
rect 494 2104 500 2105
rect 494 2100 495 2104
rect 499 2100 500 2104
rect 494 2099 500 2100
rect 590 2104 596 2105
rect 590 2100 591 2104
rect 595 2100 596 2104
rect 590 2099 596 2100
rect 694 2104 700 2105
rect 694 2100 695 2104
rect 699 2100 700 2104
rect 694 2099 700 2100
rect 798 2104 804 2105
rect 798 2100 799 2104
rect 803 2100 804 2104
rect 798 2099 804 2100
rect 910 2104 916 2105
rect 910 2100 911 2104
rect 915 2100 916 2104
rect 910 2099 916 2100
rect 1022 2104 1028 2105
rect 1022 2100 1023 2104
rect 1027 2100 1028 2104
rect 1022 2099 1028 2100
rect 1134 2104 1140 2105
rect 1134 2100 1135 2104
rect 1139 2100 1140 2104
rect 1134 2099 1140 2100
rect 1222 2104 1228 2105
rect 1222 2100 1223 2104
rect 1227 2100 1228 2104
rect 1286 2103 1287 2107
rect 1291 2103 1292 2107
rect 1286 2102 1292 2103
rect 1222 2099 1228 2100
rect 374 2092 380 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 446 2092 452 2093
rect 446 2088 447 2092
rect 451 2088 452 2092
rect 446 2087 452 2088
rect 518 2092 524 2093
rect 518 2088 519 2092
rect 523 2088 524 2092
rect 518 2087 524 2088
rect 598 2092 604 2093
rect 598 2088 599 2092
rect 603 2088 604 2092
rect 598 2087 604 2088
rect 678 2092 684 2093
rect 678 2088 679 2092
rect 683 2088 684 2092
rect 678 2087 684 2088
rect 758 2092 764 2093
rect 758 2088 759 2092
rect 763 2088 764 2092
rect 758 2087 764 2088
rect 830 2092 836 2093
rect 830 2088 831 2092
rect 835 2088 836 2092
rect 830 2087 836 2088
rect 902 2092 908 2093
rect 902 2088 903 2092
rect 907 2088 908 2092
rect 902 2087 908 2088
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 1030 2092 1036 2093
rect 1030 2088 1031 2092
rect 1035 2088 1036 2092
rect 1030 2087 1036 2088
rect 1102 2092 1108 2093
rect 1102 2088 1103 2092
rect 1107 2088 1108 2092
rect 1102 2087 1108 2088
rect 1166 2092 1172 2093
rect 1166 2088 1167 2092
rect 1171 2088 1172 2092
rect 1166 2087 1172 2088
rect 1222 2092 1228 2093
rect 1222 2088 1223 2092
rect 1227 2088 1228 2092
rect 1222 2087 1228 2088
rect 1286 2089 1292 2090
rect 110 2084 116 2085
rect 1286 2085 1287 2089
rect 1291 2085 1292 2089
rect 1286 2084 1292 2085
rect 110 2072 116 2073
rect 1286 2072 1292 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 390 2071 396 2072
rect 390 2067 391 2071
rect 395 2067 396 2071
rect 390 2066 396 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 534 2071 540 2072
rect 534 2067 535 2071
rect 539 2067 540 2071
rect 534 2066 540 2067
rect 614 2071 620 2072
rect 614 2067 615 2071
rect 619 2067 620 2071
rect 614 2066 620 2067
rect 694 2071 700 2072
rect 694 2067 695 2071
rect 699 2067 700 2071
rect 694 2066 700 2067
rect 774 2071 780 2072
rect 774 2067 775 2071
rect 779 2067 780 2071
rect 774 2066 780 2067
rect 846 2071 852 2072
rect 846 2067 847 2071
rect 851 2067 852 2071
rect 846 2066 852 2067
rect 918 2071 924 2072
rect 918 2067 919 2071
rect 923 2067 924 2071
rect 918 2066 924 2067
rect 982 2071 988 2072
rect 982 2067 983 2071
rect 987 2067 988 2071
rect 982 2066 988 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1118 2071 1124 2072
rect 1118 2067 1119 2071
rect 1123 2067 1124 2071
rect 1118 2066 1124 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 1238 2071 1244 2072
rect 1238 2067 1239 2071
rect 1243 2067 1244 2071
rect 1286 2068 1287 2072
rect 1291 2068 1292 2072
rect 1286 2067 1292 2068
rect 1238 2066 1244 2067
rect 1366 2061 1372 2062
rect 1326 2060 1332 2061
rect 1326 2056 1327 2060
rect 1331 2056 1332 2060
rect 1366 2057 1367 2061
rect 1371 2057 1372 2061
rect 1366 2056 1372 2057
rect 1422 2061 1428 2062
rect 1422 2057 1423 2061
rect 1427 2057 1428 2061
rect 1422 2056 1428 2057
rect 1502 2061 1508 2062
rect 1502 2057 1503 2061
rect 1507 2057 1508 2061
rect 1502 2056 1508 2057
rect 1590 2061 1596 2062
rect 1590 2057 1591 2061
rect 1595 2057 1596 2061
rect 1590 2056 1596 2057
rect 1678 2061 1684 2062
rect 1678 2057 1679 2061
rect 1683 2057 1684 2061
rect 1678 2056 1684 2057
rect 1782 2061 1788 2062
rect 1782 2057 1783 2061
rect 1787 2057 1788 2061
rect 1782 2056 1788 2057
rect 1894 2061 1900 2062
rect 1894 2057 1895 2061
rect 1899 2057 1900 2061
rect 1894 2056 1900 2057
rect 2022 2061 2028 2062
rect 2022 2057 2023 2061
rect 2027 2057 2028 2061
rect 2022 2056 2028 2057
rect 2166 2061 2172 2062
rect 2166 2057 2167 2061
rect 2171 2057 2172 2061
rect 2166 2056 2172 2057
rect 2318 2061 2324 2062
rect 2318 2057 2319 2061
rect 2323 2057 2324 2061
rect 2318 2056 2324 2057
rect 2454 2061 2460 2062
rect 2454 2057 2455 2061
rect 2459 2057 2460 2061
rect 2454 2056 2460 2057
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 1326 2055 1332 2056
rect 2502 2055 2508 2056
rect 1326 2043 1332 2044
rect 1326 2039 1327 2043
rect 1331 2039 1332 2043
rect 2502 2043 2508 2044
rect 1326 2038 1332 2039
rect 1350 2040 1356 2041
rect 1350 2036 1351 2040
rect 1355 2036 1356 2040
rect 1350 2035 1356 2036
rect 1406 2040 1412 2041
rect 1406 2036 1407 2040
rect 1411 2036 1412 2040
rect 1406 2035 1412 2036
rect 1486 2040 1492 2041
rect 1486 2036 1487 2040
rect 1491 2036 1492 2040
rect 1486 2035 1492 2036
rect 1574 2040 1580 2041
rect 1574 2036 1575 2040
rect 1579 2036 1580 2040
rect 1574 2035 1580 2036
rect 1662 2040 1668 2041
rect 1662 2036 1663 2040
rect 1667 2036 1668 2040
rect 1662 2035 1668 2036
rect 1766 2040 1772 2041
rect 1766 2036 1767 2040
rect 1771 2036 1772 2040
rect 1766 2035 1772 2036
rect 1878 2040 1884 2041
rect 1878 2036 1879 2040
rect 1883 2036 1884 2040
rect 1878 2035 1884 2036
rect 2006 2040 2012 2041
rect 2006 2036 2007 2040
rect 2011 2036 2012 2040
rect 2006 2035 2012 2036
rect 2150 2040 2156 2041
rect 2150 2036 2151 2040
rect 2155 2036 2156 2040
rect 2150 2035 2156 2036
rect 2302 2040 2308 2041
rect 2302 2036 2303 2040
rect 2307 2036 2308 2040
rect 2302 2035 2308 2036
rect 2438 2040 2444 2041
rect 2438 2036 2439 2040
rect 2443 2036 2444 2040
rect 2502 2039 2503 2043
rect 2507 2039 2508 2043
rect 2502 2038 2508 2039
rect 2438 2035 2444 2036
rect 1350 2028 1356 2029
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1350 2024 1351 2028
rect 1355 2024 1356 2028
rect 1350 2023 1356 2024
rect 1422 2028 1428 2029
rect 1422 2024 1423 2028
rect 1427 2024 1428 2028
rect 1422 2023 1428 2024
rect 1518 2028 1524 2029
rect 1518 2024 1519 2028
rect 1523 2024 1524 2028
rect 1518 2023 1524 2024
rect 1614 2028 1620 2029
rect 1614 2024 1615 2028
rect 1619 2024 1620 2028
rect 1614 2023 1620 2024
rect 1718 2028 1724 2029
rect 1718 2024 1719 2028
rect 1723 2024 1724 2028
rect 1718 2023 1724 2024
rect 1822 2028 1828 2029
rect 1822 2024 1823 2028
rect 1827 2024 1828 2028
rect 1822 2023 1828 2024
rect 1934 2028 1940 2029
rect 1934 2024 1935 2028
rect 1939 2024 1940 2028
rect 1934 2023 1940 2024
rect 2054 2028 2060 2029
rect 2054 2024 2055 2028
rect 2059 2024 2060 2028
rect 2054 2023 2060 2024
rect 2182 2028 2188 2029
rect 2182 2024 2183 2028
rect 2187 2024 2188 2028
rect 2182 2023 2188 2024
rect 2318 2028 2324 2029
rect 2318 2024 2319 2028
rect 2323 2024 2324 2028
rect 2318 2023 2324 2024
rect 2438 2028 2444 2029
rect 2438 2024 2439 2028
rect 2443 2024 2444 2028
rect 2438 2023 2444 2024
rect 2502 2025 2508 2026
rect 1326 2020 1332 2021
rect 2502 2021 2503 2025
rect 2507 2021 2508 2025
rect 2502 2020 2508 2021
rect 294 2017 300 2018
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 294 2013 295 2017
rect 299 2013 300 2017
rect 294 2012 300 2013
rect 374 2017 380 2018
rect 374 2013 375 2017
rect 379 2013 380 2017
rect 374 2012 380 2013
rect 462 2017 468 2018
rect 462 2013 463 2017
rect 467 2013 468 2017
rect 462 2012 468 2013
rect 550 2017 556 2018
rect 550 2013 551 2017
rect 555 2013 556 2017
rect 550 2012 556 2013
rect 638 2017 644 2018
rect 638 2013 639 2017
rect 643 2013 644 2017
rect 638 2012 644 2013
rect 718 2017 724 2018
rect 718 2013 719 2017
rect 723 2013 724 2017
rect 718 2012 724 2013
rect 798 2017 804 2018
rect 798 2013 799 2017
rect 803 2013 804 2017
rect 798 2012 804 2013
rect 886 2017 892 2018
rect 886 2013 887 2017
rect 891 2013 892 2017
rect 886 2012 892 2013
rect 974 2017 980 2018
rect 974 2013 975 2017
rect 979 2013 980 2017
rect 974 2012 980 2013
rect 1062 2017 1068 2018
rect 1062 2013 1063 2017
rect 1067 2013 1068 2017
rect 1062 2012 1068 2013
rect 1286 2016 1292 2017
rect 1286 2012 1287 2016
rect 1291 2012 1292 2016
rect 110 2011 116 2012
rect 1286 2011 1292 2012
rect 1326 2008 1332 2009
rect 2502 2008 2508 2009
rect 1326 2004 1327 2008
rect 1331 2004 1332 2008
rect 1326 2003 1332 2004
rect 1366 2007 1372 2008
rect 1366 2003 1367 2007
rect 1371 2003 1372 2007
rect 1366 2002 1372 2003
rect 1438 2007 1444 2008
rect 1438 2003 1439 2007
rect 1443 2003 1444 2007
rect 1438 2002 1444 2003
rect 1534 2007 1540 2008
rect 1534 2003 1535 2007
rect 1539 2003 1540 2007
rect 1534 2002 1540 2003
rect 1630 2007 1636 2008
rect 1630 2003 1631 2007
rect 1635 2003 1636 2007
rect 1630 2002 1636 2003
rect 1734 2007 1740 2008
rect 1734 2003 1735 2007
rect 1739 2003 1740 2007
rect 1734 2002 1740 2003
rect 1838 2007 1844 2008
rect 1838 2003 1839 2007
rect 1843 2003 1844 2007
rect 1838 2002 1844 2003
rect 1950 2007 1956 2008
rect 1950 2003 1951 2007
rect 1955 2003 1956 2007
rect 1950 2002 1956 2003
rect 2070 2007 2076 2008
rect 2070 2003 2071 2007
rect 2075 2003 2076 2007
rect 2070 2002 2076 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2334 2007 2340 2008
rect 2334 2003 2335 2007
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2454 2007 2460 2008
rect 2454 2003 2455 2007
rect 2459 2003 2460 2007
rect 2502 2004 2503 2008
rect 2507 2004 2508 2008
rect 2502 2003 2508 2004
rect 2454 2002 2460 2003
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1286 1999 1292 2000
rect 110 1994 116 1995
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 358 1996 364 1997
rect 358 1992 359 1996
rect 363 1992 364 1996
rect 358 1991 364 1992
rect 446 1996 452 1997
rect 446 1992 447 1996
rect 451 1992 452 1996
rect 446 1991 452 1992
rect 534 1996 540 1997
rect 534 1992 535 1996
rect 539 1992 540 1996
rect 534 1991 540 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 702 1996 708 1997
rect 702 1992 703 1996
rect 707 1992 708 1996
rect 702 1991 708 1992
rect 782 1996 788 1997
rect 782 1992 783 1996
rect 787 1992 788 1996
rect 782 1991 788 1992
rect 870 1996 876 1997
rect 870 1992 871 1996
rect 875 1992 876 1996
rect 870 1991 876 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1286 1995 1287 1999
rect 1291 1995 1292 1999
rect 1286 1994 1292 1995
rect 1046 1991 1052 1992
rect 134 1980 140 1981
rect 110 1977 116 1978
rect 110 1973 111 1977
rect 115 1973 116 1977
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 206 1980 212 1981
rect 206 1976 207 1980
rect 211 1976 212 1980
rect 206 1975 212 1976
rect 286 1980 292 1981
rect 286 1976 287 1980
rect 291 1976 292 1980
rect 286 1975 292 1976
rect 382 1980 388 1981
rect 382 1976 383 1980
rect 387 1976 388 1980
rect 382 1975 388 1976
rect 486 1980 492 1981
rect 486 1976 487 1980
rect 491 1976 492 1980
rect 486 1975 492 1976
rect 590 1980 596 1981
rect 590 1976 591 1980
rect 595 1976 596 1980
rect 590 1975 596 1976
rect 694 1980 700 1981
rect 694 1976 695 1980
rect 699 1976 700 1980
rect 694 1975 700 1976
rect 798 1980 804 1981
rect 798 1976 799 1980
rect 803 1976 804 1980
rect 798 1975 804 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1014 1980 1020 1981
rect 1014 1976 1015 1980
rect 1019 1976 1020 1980
rect 1014 1975 1020 1976
rect 1286 1977 1292 1978
rect 110 1972 116 1973
rect 1286 1973 1287 1977
rect 1291 1973 1292 1977
rect 1286 1972 1292 1973
rect 110 1960 116 1961
rect 1286 1960 1292 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 110 1955 116 1956
rect 150 1959 156 1960
rect 150 1955 151 1959
rect 155 1955 156 1959
rect 150 1954 156 1955
rect 222 1959 228 1960
rect 222 1955 223 1959
rect 227 1955 228 1959
rect 222 1954 228 1955
rect 302 1959 308 1960
rect 302 1955 303 1959
rect 307 1955 308 1959
rect 302 1954 308 1955
rect 398 1959 404 1960
rect 398 1955 399 1959
rect 403 1955 404 1959
rect 398 1954 404 1955
rect 502 1959 508 1960
rect 502 1955 503 1959
rect 507 1955 508 1959
rect 502 1954 508 1955
rect 606 1959 612 1960
rect 606 1955 607 1959
rect 611 1955 612 1959
rect 606 1954 612 1955
rect 710 1959 716 1960
rect 710 1955 711 1959
rect 715 1955 716 1959
rect 710 1954 716 1955
rect 814 1959 820 1960
rect 814 1955 815 1959
rect 819 1955 820 1959
rect 814 1954 820 1955
rect 918 1959 924 1960
rect 918 1955 919 1959
rect 923 1955 924 1959
rect 918 1954 924 1955
rect 1030 1959 1036 1960
rect 1030 1955 1031 1959
rect 1035 1955 1036 1959
rect 1286 1956 1287 1960
rect 1291 1956 1292 1960
rect 1286 1955 1292 1956
rect 1030 1954 1036 1955
rect 1454 1953 1460 1954
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1542 1953 1548 1954
rect 1542 1949 1543 1953
rect 1547 1949 1548 1953
rect 1542 1948 1548 1949
rect 1638 1953 1644 1954
rect 1638 1949 1639 1953
rect 1643 1949 1644 1953
rect 1638 1948 1644 1949
rect 1734 1953 1740 1954
rect 1734 1949 1735 1953
rect 1739 1949 1740 1953
rect 1734 1948 1740 1949
rect 1838 1953 1844 1954
rect 1838 1949 1839 1953
rect 1843 1949 1844 1953
rect 1838 1948 1844 1949
rect 1942 1953 1948 1954
rect 1942 1949 1943 1953
rect 1947 1949 1948 1953
rect 1942 1948 1948 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2046 1948 2052 1949
rect 2150 1953 2156 1954
rect 2150 1949 2151 1953
rect 2155 1949 2156 1953
rect 2150 1948 2156 1949
rect 2254 1953 2260 1954
rect 2254 1949 2255 1953
rect 2259 1949 2260 1953
rect 2254 1948 2260 1949
rect 2366 1953 2372 1954
rect 2366 1949 2367 1953
rect 2371 1949 2372 1953
rect 2366 1948 2372 1949
rect 2454 1953 2460 1954
rect 2454 1949 2455 1953
rect 2459 1949 2460 1953
rect 2454 1948 2460 1949
rect 2502 1952 2508 1953
rect 2502 1948 2503 1952
rect 2507 1948 2508 1952
rect 1326 1947 1332 1948
rect 2502 1947 2508 1948
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 2502 1935 2508 1936
rect 1326 1930 1332 1931
rect 1438 1932 1444 1933
rect 1438 1928 1439 1932
rect 1443 1928 1444 1932
rect 1438 1927 1444 1928
rect 1526 1932 1532 1933
rect 1526 1928 1527 1932
rect 1531 1928 1532 1932
rect 1526 1927 1532 1928
rect 1622 1932 1628 1933
rect 1622 1928 1623 1932
rect 1627 1928 1628 1932
rect 1622 1927 1628 1928
rect 1718 1932 1724 1933
rect 1718 1928 1719 1932
rect 1723 1928 1724 1932
rect 1718 1927 1724 1928
rect 1822 1932 1828 1933
rect 1822 1928 1823 1932
rect 1827 1928 1828 1932
rect 1822 1927 1828 1928
rect 1926 1932 1932 1933
rect 1926 1928 1927 1932
rect 1931 1928 1932 1932
rect 1926 1927 1932 1928
rect 2030 1932 2036 1933
rect 2030 1928 2031 1932
rect 2035 1928 2036 1932
rect 2030 1927 2036 1928
rect 2134 1932 2140 1933
rect 2134 1928 2135 1932
rect 2139 1928 2140 1932
rect 2134 1927 2140 1928
rect 2238 1932 2244 1933
rect 2238 1928 2239 1932
rect 2243 1928 2244 1932
rect 2238 1927 2244 1928
rect 2350 1932 2356 1933
rect 2350 1928 2351 1932
rect 2355 1928 2356 1932
rect 2350 1927 2356 1928
rect 2438 1932 2444 1933
rect 2438 1928 2439 1932
rect 2443 1928 2444 1932
rect 2502 1931 2503 1935
rect 2507 1931 2508 1935
rect 2502 1930 2508 1931
rect 2438 1927 2444 1928
rect 1526 1916 1532 1917
rect 1326 1913 1332 1914
rect 1326 1909 1327 1913
rect 1331 1909 1332 1913
rect 1526 1912 1527 1916
rect 1531 1912 1532 1916
rect 1526 1911 1532 1912
rect 1614 1916 1620 1917
rect 1614 1912 1615 1916
rect 1619 1912 1620 1916
rect 1614 1911 1620 1912
rect 1710 1916 1716 1917
rect 1710 1912 1711 1916
rect 1715 1912 1716 1916
rect 1710 1911 1716 1912
rect 1814 1916 1820 1917
rect 1814 1912 1815 1916
rect 1819 1912 1820 1916
rect 1814 1911 1820 1912
rect 1918 1916 1924 1917
rect 1918 1912 1919 1916
rect 1923 1912 1924 1916
rect 1918 1911 1924 1912
rect 2014 1916 2020 1917
rect 2014 1912 2015 1916
rect 2019 1912 2020 1916
rect 2014 1911 2020 1912
rect 2110 1916 2116 1917
rect 2110 1912 2111 1916
rect 2115 1912 2116 1916
rect 2110 1911 2116 1912
rect 2198 1916 2204 1917
rect 2198 1912 2199 1916
rect 2203 1912 2204 1916
rect 2198 1911 2204 1912
rect 2286 1916 2292 1917
rect 2286 1912 2287 1916
rect 2291 1912 2292 1916
rect 2286 1911 2292 1912
rect 2374 1916 2380 1917
rect 2374 1912 2375 1916
rect 2379 1912 2380 1916
rect 2374 1911 2380 1912
rect 2438 1916 2444 1917
rect 2438 1912 2439 1916
rect 2443 1912 2444 1916
rect 2438 1911 2444 1912
rect 2502 1913 2508 1914
rect 1326 1908 1332 1909
rect 2502 1909 2503 1913
rect 2507 1909 2508 1913
rect 2502 1908 2508 1909
rect 150 1901 156 1902
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 150 1897 151 1901
rect 155 1897 156 1901
rect 150 1896 156 1897
rect 238 1901 244 1902
rect 238 1897 239 1901
rect 243 1897 244 1901
rect 238 1896 244 1897
rect 374 1901 380 1902
rect 374 1897 375 1901
rect 379 1897 380 1901
rect 374 1896 380 1897
rect 526 1901 532 1902
rect 526 1897 527 1901
rect 531 1897 532 1901
rect 526 1896 532 1897
rect 686 1901 692 1902
rect 686 1897 687 1901
rect 691 1897 692 1901
rect 686 1896 692 1897
rect 862 1901 868 1902
rect 862 1897 863 1901
rect 867 1897 868 1901
rect 862 1896 868 1897
rect 1038 1901 1044 1902
rect 1038 1897 1039 1901
rect 1043 1897 1044 1901
rect 1038 1896 1044 1897
rect 1286 1900 1292 1901
rect 1286 1896 1287 1900
rect 1291 1896 1292 1900
rect 110 1895 116 1896
rect 1286 1895 1292 1896
rect 1326 1896 1332 1897
rect 2502 1896 2508 1897
rect 1326 1892 1327 1896
rect 1331 1892 1332 1896
rect 1326 1891 1332 1892
rect 1542 1895 1548 1896
rect 1542 1891 1543 1895
rect 1547 1891 1548 1895
rect 1542 1890 1548 1891
rect 1630 1895 1636 1896
rect 1630 1891 1631 1895
rect 1635 1891 1636 1895
rect 1630 1890 1636 1891
rect 1726 1895 1732 1896
rect 1726 1891 1727 1895
rect 1731 1891 1732 1895
rect 1726 1890 1732 1891
rect 1830 1895 1836 1896
rect 1830 1891 1831 1895
rect 1835 1891 1836 1895
rect 1830 1890 1836 1891
rect 1934 1895 1940 1896
rect 1934 1891 1935 1895
rect 1939 1891 1940 1895
rect 1934 1890 1940 1891
rect 2030 1895 2036 1896
rect 2030 1891 2031 1895
rect 2035 1891 2036 1895
rect 2030 1890 2036 1891
rect 2126 1895 2132 1896
rect 2126 1891 2127 1895
rect 2131 1891 2132 1895
rect 2126 1890 2132 1891
rect 2214 1895 2220 1896
rect 2214 1891 2215 1895
rect 2219 1891 2220 1895
rect 2214 1890 2220 1891
rect 2302 1895 2308 1896
rect 2302 1891 2303 1895
rect 2307 1891 2308 1895
rect 2302 1890 2308 1891
rect 2390 1895 2396 1896
rect 2390 1891 2391 1895
rect 2395 1891 2396 1895
rect 2390 1890 2396 1891
rect 2454 1895 2460 1896
rect 2454 1891 2455 1895
rect 2459 1891 2460 1895
rect 2502 1892 2503 1896
rect 2507 1892 2508 1896
rect 2502 1891 2508 1892
rect 2454 1890 2460 1891
rect 110 1883 116 1884
rect 110 1879 111 1883
rect 115 1879 116 1883
rect 1286 1883 1292 1884
rect 110 1878 116 1879
rect 134 1880 140 1881
rect 134 1876 135 1880
rect 139 1876 140 1880
rect 134 1875 140 1876
rect 222 1880 228 1881
rect 222 1876 223 1880
rect 227 1876 228 1880
rect 222 1875 228 1876
rect 358 1880 364 1881
rect 358 1876 359 1880
rect 363 1876 364 1880
rect 358 1875 364 1876
rect 510 1880 516 1881
rect 510 1876 511 1880
rect 515 1876 516 1880
rect 510 1875 516 1876
rect 670 1880 676 1881
rect 670 1876 671 1880
rect 675 1876 676 1880
rect 670 1875 676 1876
rect 846 1880 852 1881
rect 846 1876 847 1880
rect 851 1876 852 1880
rect 846 1875 852 1876
rect 1022 1880 1028 1881
rect 1022 1876 1023 1880
rect 1027 1876 1028 1880
rect 1286 1879 1287 1883
rect 1291 1879 1292 1883
rect 1286 1878 1292 1879
rect 1022 1875 1028 1876
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 190 1868 196 1869
rect 190 1864 191 1868
rect 195 1864 196 1868
rect 190 1863 196 1864
rect 262 1868 268 1869
rect 262 1864 263 1868
rect 267 1864 268 1868
rect 262 1863 268 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 406 1868 412 1869
rect 406 1864 407 1868
rect 411 1864 412 1868
rect 406 1863 412 1864
rect 478 1868 484 1869
rect 478 1864 479 1868
rect 483 1864 484 1868
rect 478 1863 484 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 614 1868 620 1869
rect 614 1864 615 1868
rect 619 1864 620 1868
rect 614 1863 620 1864
rect 678 1868 684 1869
rect 678 1864 679 1868
rect 683 1864 684 1868
rect 678 1863 684 1864
rect 742 1868 748 1869
rect 742 1864 743 1868
rect 747 1864 748 1868
rect 742 1863 748 1864
rect 814 1868 820 1869
rect 814 1864 815 1868
rect 819 1864 820 1868
rect 814 1863 820 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 958 1868 964 1869
rect 958 1864 959 1868
rect 963 1864 964 1868
rect 958 1863 964 1864
rect 1038 1868 1044 1869
rect 1038 1864 1039 1868
rect 1043 1864 1044 1868
rect 1038 1863 1044 1864
rect 1286 1865 1292 1866
rect 110 1860 116 1861
rect 1286 1861 1287 1865
rect 1291 1861 1292 1865
rect 1286 1860 1292 1861
rect 110 1848 116 1849
rect 1286 1848 1292 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 150 1847 156 1848
rect 150 1843 151 1847
rect 155 1843 156 1847
rect 150 1842 156 1843
rect 206 1847 212 1848
rect 206 1843 207 1847
rect 211 1843 212 1847
rect 206 1842 212 1843
rect 278 1847 284 1848
rect 278 1843 279 1847
rect 283 1843 284 1847
rect 278 1842 284 1843
rect 350 1847 356 1848
rect 350 1843 351 1847
rect 355 1843 356 1847
rect 350 1842 356 1843
rect 422 1847 428 1848
rect 422 1843 423 1847
rect 427 1843 428 1847
rect 422 1842 428 1843
rect 494 1847 500 1848
rect 494 1843 495 1847
rect 499 1843 500 1847
rect 494 1842 500 1843
rect 566 1847 572 1848
rect 566 1843 567 1847
rect 571 1843 572 1847
rect 566 1842 572 1843
rect 630 1847 636 1848
rect 630 1843 631 1847
rect 635 1843 636 1847
rect 630 1842 636 1843
rect 694 1847 700 1848
rect 694 1843 695 1847
rect 699 1843 700 1847
rect 694 1842 700 1843
rect 758 1847 764 1848
rect 758 1843 759 1847
rect 763 1843 764 1847
rect 758 1842 764 1843
rect 830 1847 836 1848
rect 830 1843 831 1847
rect 835 1843 836 1847
rect 830 1842 836 1843
rect 902 1847 908 1848
rect 902 1843 903 1847
rect 907 1843 908 1847
rect 902 1842 908 1843
rect 974 1847 980 1848
rect 974 1843 975 1847
rect 979 1843 980 1847
rect 974 1842 980 1843
rect 1054 1847 1060 1848
rect 1054 1843 1055 1847
rect 1059 1843 1060 1847
rect 1286 1844 1287 1848
rect 1291 1844 1292 1848
rect 1534 1845 1540 1846
rect 1286 1843 1292 1844
rect 1326 1844 1332 1845
rect 1054 1842 1060 1843
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1534 1841 1535 1845
rect 1539 1841 1540 1845
rect 1534 1840 1540 1841
rect 1606 1845 1612 1846
rect 1606 1841 1607 1845
rect 1611 1841 1612 1845
rect 1606 1840 1612 1841
rect 1686 1845 1692 1846
rect 1686 1841 1687 1845
rect 1691 1841 1692 1845
rect 1686 1840 1692 1841
rect 1782 1845 1788 1846
rect 1782 1841 1783 1845
rect 1787 1841 1788 1845
rect 1782 1840 1788 1841
rect 1878 1845 1884 1846
rect 1878 1841 1879 1845
rect 1883 1841 1884 1845
rect 1878 1840 1884 1841
rect 1982 1845 1988 1846
rect 1982 1841 1983 1845
rect 1987 1841 1988 1845
rect 1982 1840 1988 1841
rect 2078 1845 2084 1846
rect 2078 1841 2079 1845
rect 2083 1841 2084 1845
rect 2078 1840 2084 1841
rect 2174 1845 2180 1846
rect 2174 1841 2175 1845
rect 2179 1841 2180 1845
rect 2174 1840 2180 1841
rect 2270 1845 2276 1846
rect 2270 1841 2271 1845
rect 2275 1841 2276 1845
rect 2270 1840 2276 1841
rect 2366 1845 2372 1846
rect 2366 1841 2367 1845
rect 2371 1841 2372 1845
rect 2366 1840 2372 1841
rect 2454 1845 2460 1846
rect 2454 1841 2455 1845
rect 2459 1841 2460 1845
rect 2454 1840 2460 1841
rect 2502 1844 2508 1845
rect 2502 1840 2503 1844
rect 2507 1840 2508 1844
rect 1326 1839 1332 1840
rect 2502 1839 2508 1840
rect 1326 1827 1332 1828
rect 1326 1823 1327 1827
rect 1331 1823 1332 1827
rect 2502 1827 2508 1828
rect 1326 1822 1332 1823
rect 1518 1824 1524 1825
rect 1518 1820 1519 1824
rect 1523 1820 1524 1824
rect 1518 1819 1524 1820
rect 1590 1824 1596 1825
rect 1590 1820 1591 1824
rect 1595 1820 1596 1824
rect 1590 1819 1596 1820
rect 1670 1824 1676 1825
rect 1670 1820 1671 1824
rect 1675 1820 1676 1824
rect 1670 1819 1676 1820
rect 1766 1824 1772 1825
rect 1766 1820 1767 1824
rect 1771 1820 1772 1824
rect 1766 1819 1772 1820
rect 1862 1824 1868 1825
rect 1862 1820 1863 1824
rect 1867 1820 1868 1824
rect 1862 1819 1868 1820
rect 1966 1824 1972 1825
rect 1966 1820 1967 1824
rect 1971 1820 1972 1824
rect 1966 1819 1972 1820
rect 2062 1824 2068 1825
rect 2062 1820 2063 1824
rect 2067 1820 2068 1824
rect 2062 1819 2068 1820
rect 2158 1824 2164 1825
rect 2158 1820 2159 1824
rect 2163 1820 2164 1824
rect 2158 1819 2164 1820
rect 2254 1824 2260 1825
rect 2254 1820 2255 1824
rect 2259 1820 2260 1824
rect 2254 1819 2260 1820
rect 2350 1824 2356 1825
rect 2350 1820 2351 1824
rect 2355 1820 2356 1824
rect 2350 1819 2356 1820
rect 2438 1824 2444 1825
rect 2438 1820 2439 1824
rect 2443 1820 2444 1824
rect 2502 1823 2503 1827
rect 2507 1823 2508 1827
rect 2502 1822 2508 1823
rect 2438 1819 2444 1820
rect 1462 1808 1468 1809
rect 1326 1805 1332 1806
rect 1326 1801 1327 1805
rect 1331 1801 1332 1805
rect 1462 1804 1463 1808
rect 1467 1804 1468 1808
rect 1462 1803 1468 1804
rect 1558 1808 1564 1809
rect 1558 1804 1559 1808
rect 1563 1804 1564 1808
rect 1558 1803 1564 1804
rect 1662 1808 1668 1809
rect 1662 1804 1663 1808
rect 1667 1804 1668 1808
rect 1662 1803 1668 1804
rect 1766 1808 1772 1809
rect 1766 1804 1767 1808
rect 1771 1804 1772 1808
rect 1766 1803 1772 1804
rect 1878 1808 1884 1809
rect 1878 1804 1879 1808
rect 1883 1804 1884 1808
rect 1878 1803 1884 1804
rect 1982 1808 1988 1809
rect 1982 1804 1983 1808
rect 1987 1804 1988 1808
rect 1982 1803 1988 1804
rect 2086 1808 2092 1809
rect 2086 1804 2087 1808
rect 2091 1804 2092 1808
rect 2086 1803 2092 1804
rect 2182 1808 2188 1809
rect 2182 1804 2183 1808
rect 2187 1804 2188 1808
rect 2182 1803 2188 1804
rect 2270 1808 2276 1809
rect 2270 1804 2271 1808
rect 2275 1804 2276 1808
rect 2270 1803 2276 1804
rect 2366 1808 2372 1809
rect 2366 1804 2367 1808
rect 2371 1804 2372 1808
rect 2366 1803 2372 1804
rect 2438 1808 2444 1809
rect 2438 1804 2439 1808
rect 2443 1804 2444 1808
rect 2438 1803 2444 1804
rect 2502 1805 2508 1806
rect 1326 1800 1332 1801
rect 2502 1801 2503 1805
rect 2507 1801 2508 1805
rect 2502 1800 2508 1801
rect 150 1789 156 1790
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 150 1785 151 1789
rect 155 1785 156 1789
rect 150 1784 156 1785
rect 230 1789 236 1790
rect 230 1785 231 1789
rect 235 1785 236 1789
rect 230 1784 236 1785
rect 334 1789 340 1790
rect 334 1785 335 1789
rect 339 1785 340 1789
rect 334 1784 340 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 534 1789 540 1790
rect 534 1785 535 1789
rect 539 1785 540 1789
rect 534 1784 540 1785
rect 630 1789 636 1790
rect 630 1785 631 1789
rect 635 1785 636 1789
rect 630 1784 636 1785
rect 718 1789 724 1790
rect 718 1785 719 1789
rect 723 1785 724 1789
rect 718 1784 724 1785
rect 798 1789 804 1790
rect 798 1785 799 1789
rect 803 1785 804 1789
rect 798 1784 804 1785
rect 878 1789 884 1790
rect 878 1785 879 1789
rect 883 1785 884 1789
rect 878 1784 884 1785
rect 958 1789 964 1790
rect 958 1785 959 1789
rect 963 1785 964 1789
rect 958 1784 964 1785
rect 1038 1789 1044 1790
rect 1038 1785 1039 1789
rect 1043 1785 1044 1789
rect 1038 1784 1044 1785
rect 1118 1789 1124 1790
rect 1118 1785 1119 1789
rect 1123 1785 1124 1789
rect 1118 1784 1124 1785
rect 1286 1788 1292 1789
rect 1286 1784 1287 1788
rect 1291 1784 1292 1788
rect 110 1783 116 1784
rect 1286 1783 1292 1784
rect 1326 1788 1332 1789
rect 2502 1788 2508 1789
rect 1326 1784 1327 1788
rect 1331 1784 1332 1788
rect 1326 1783 1332 1784
rect 1478 1787 1484 1788
rect 1478 1783 1479 1787
rect 1483 1783 1484 1787
rect 1478 1782 1484 1783
rect 1574 1787 1580 1788
rect 1574 1783 1575 1787
rect 1579 1783 1580 1787
rect 1574 1782 1580 1783
rect 1678 1787 1684 1788
rect 1678 1783 1679 1787
rect 1683 1783 1684 1787
rect 1678 1782 1684 1783
rect 1782 1787 1788 1788
rect 1782 1783 1783 1787
rect 1787 1783 1788 1787
rect 1782 1782 1788 1783
rect 1894 1787 1900 1788
rect 1894 1783 1895 1787
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1998 1787 2004 1788
rect 1998 1783 1999 1787
rect 2003 1783 2004 1787
rect 1998 1782 2004 1783
rect 2102 1787 2108 1788
rect 2102 1783 2103 1787
rect 2107 1783 2108 1787
rect 2102 1782 2108 1783
rect 2198 1787 2204 1788
rect 2198 1783 2199 1787
rect 2203 1783 2204 1787
rect 2198 1782 2204 1783
rect 2286 1787 2292 1788
rect 2286 1783 2287 1787
rect 2291 1783 2292 1787
rect 2286 1782 2292 1783
rect 2382 1787 2388 1788
rect 2382 1783 2383 1787
rect 2387 1783 2388 1787
rect 2382 1782 2388 1783
rect 2454 1787 2460 1788
rect 2454 1783 2455 1787
rect 2459 1783 2460 1787
rect 2502 1784 2503 1788
rect 2507 1784 2508 1788
rect 2502 1783 2508 1784
rect 2454 1782 2460 1783
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1286 1771 1292 1772
rect 110 1766 116 1767
rect 134 1768 140 1769
rect 134 1764 135 1768
rect 139 1764 140 1768
rect 134 1763 140 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 318 1768 324 1769
rect 318 1764 319 1768
rect 323 1764 324 1768
rect 318 1763 324 1764
rect 422 1768 428 1769
rect 422 1764 423 1768
rect 427 1764 428 1768
rect 422 1763 428 1764
rect 518 1768 524 1769
rect 518 1764 519 1768
rect 523 1764 524 1768
rect 518 1763 524 1764
rect 614 1768 620 1769
rect 614 1764 615 1768
rect 619 1764 620 1768
rect 614 1763 620 1764
rect 702 1768 708 1769
rect 702 1764 703 1768
rect 707 1764 708 1768
rect 702 1763 708 1764
rect 782 1768 788 1769
rect 782 1764 783 1768
rect 787 1764 788 1768
rect 782 1763 788 1764
rect 862 1768 868 1769
rect 862 1764 863 1768
rect 867 1764 868 1768
rect 862 1763 868 1764
rect 942 1768 948 1769
rect 942 1764 943 1768
rect 947 1764 948 1768
rect 942 1763 948 1764
rect 1022 1768 1028 1769
rect 1022 1764 1023 1768
rect 1027 1764 1028 1768
rect 1022 1763 1028 1764
rect 1102 1768 1108 1769
rect 1102 1764 1103 1768
rect 1107 1764 1108 1768
rect 1286 1767 1287 1771
rect 1291 1767 1292 1771
rect 1286 1766 1292 1767
rect 1102 1763 1108 1764
rect 134 1752 140 1753
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 134 1748 135 1752
rect 139 1748 140 1752
rect 134 1747 140 1748
rect 238 1752 244 1753
rect 238 1748 239 1752
rect 243 1748 244 1752
rect 238 1747 244 1748
rect 350 1752 356 1753
rect 350 1748 351 1752
rect 355 1748 356 1752
rect 350 1747 356 1748
rect 462 1752 468 1753
rect 462 1748 463 1752
rect 467 1748 468 1752
rect 462 1747 468 1748
rect 574 1752 580 1753
rect 574 1748 575 1752
rect 579 1748 580 1752
rect 574 1747 580 1748
rect 678 1752 684 1753
rect 678 1748 679 1752
rect 683 1748 684 1752
rect 678 1747 684 1748
rect 782 1752 788 1753
rect 782 1748 783 1752
rect 787 1748 788 1752
rect 782 1747 788 1748
rect 886 1752 892 1753
rect 886 1748 887 1752
rect 891 1748 892 1752
rect 886 1747 892 1748
rect 990 1752 996 1753
rect 990 1748 991 1752
rect 995 1748 996 1752
rect 990 1747 996 1748
rect 1102 1752 1108 1753
rect 1102 1748 1103 1752
rect 1107 1748 1108 1752
rect 1102 1747 1108 1748
rect 1286 1749 1292 1750
rect 110 1744 116 1745
rect 1286 1745 1287 1749
rect 1291 1745 1292 1749
rect 1286 1744 1292 1745
rect 1374 1733 1380 1734
rect 110 1732 116 1733
rect 1286 1732 1292 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 150 1731 156 1732
rect 150 1727 151 1731
rect 155 1727 156 1731
rect 150 1726 156 1727
rect 254 1731 260 1732
rect 254 1727 255 1731
rect 259 1727 260 1731
rect 254 1726 260 1727
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 478 1731 484 1732
rect 478 1727 479 1731
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 590 1731 596 1732
rect 590 1727 591 1731
rect 595 1727 596 1731
rect 590 1726 596 1727
rect 694 1731 700 1732
rect 694 1727 695 1731
rect 699 1727 700 1731
rect 694 1726 700 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 902 1731 908 1732
rect 902 1727 903 1731
rect 907 1727 908 1731
rect 902 1726 908 1727
rect 1006 1731 1012 1732
rect 1006 1727 1007 1731
rect 1011 1727 1012 1731
rect 1006 1726 1012 1727
rect 1118 1731 1124 1732
rect 1118 1727 1119 1731
rect 1123 1727 1124 1731
rect 1286 1728 1287 1732
rect 1291 1728 1292 1732
rect 1286 1727 1292 1728
rect 1326 1732 1332 1733
rect 1326 1728 1327 1732
rect 1331 1728 1332 1732
rect 1374 1729 1375 1733
rect 1379 1729 1380 1733
rect 1374 1728 1380 1729
rect 1470 1733 1476 1734
rect 1470 1729 1471 1733
rect 1475 1729 1476 1733
rect 1470 1728 1476 1729
rect 1566 1733 1572 1734
rect 1566 1729 1567 1733
rect 1571 1729 1572 1733
rect 1566 1728 1572 1729
rect 1670 1733 1676 1734
rect 1670 1729 1671 1733
rect 1675 1729 1676 1733
rect 1670 1728 1676 1729
rect 1774 1733 1780 1734
rect 1774 1729 1775 1733
rect 1779 1729 1780 1733
rect 1774 1728 1780 1729
rect 1886 1733 1892 1734
rect 1886 1729 1887 1733
rect 1891 1729 1892 1733
rect 1886 1728 1892 1729
rect 1998 1733 2004 1734
rect 1998 1729 1999 1733
rect 2003 1729 2004 1733
rect 1998 1728 2004 1729
rect 2110 1733 2116 1734
rect 2110 1729 2111 1733
rect 2115 1729 2116 1733
rect 2110 1728 2116 1729
rect 2230 1733 2236 1734
rect 2230 1729 2231 1733
rect 2235 1729 2236 1733
rect 2230 1728 2236 1729
rect 2350 1733 2356 1734
rect 2350 1729 2351 1733
rect 2355 1729 2356 1733
rect 2350 1728 2356 1729
rect 2454 1733 2460 1734
rect 2454 1729 2455 1733
rect 2459 1729 2460 1733
rect 2454 1728 2460 1729
rect 2502 1732 2508 1733
rect 2502 1728 2503 1732
rect 2507 1728 2508 1732
rect 1326 1727 1332 1728
rect 2502 1727 2508 1728
rect 1118 1726 1124 1727
rect 1326 1715 1332 1716
rect 1326 1711 1327 1715
rect 1331 1711 1332 1715
rect 2502 1715 2508 1716
rect 1326 1710 1332 1711
rect 1358 1712 1364 1713
rect 1358 1708 1359 1712
rect 1363 1708 1364 1712
rect 1358 1707 1364 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1550 1712 1556 1713
rect 1550 1708 1551 1712
rect 1555 1708 1556 1712
rect 1550 1707 1556 1708
rect 1654 1712 1660 1713
rect 1654 1708 1655 1712
rect 1659 1708 1660 1712
rect 1654 1707 1660 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1870 1712 1876 1713
rect 1870 1708 1871 1712
rect 1875 1708 1876 1712
rect 1870 1707 1876 1708
rect 1982 1712 1988 1713
rect 1982 1708 1983 1712
rect 1987 1708 1988 1712
rect 1982 1707 1988 1708
rect 2094 1712 2100 1713
rect 2094 1708 2095 1712
rect 2099 1708 2100 1712
rect 2094 1707 2100 1708
rect 2214 1712 2220 1713
rect 2214 1708 2215 1712
rect 2219 1708 2220 1712
rect 2214 1707 2220 1708
rect 2334 1712 2340 1713
rect 2334 1708 2335 1712
rect 2339 1708 2340 1712
rect 2334 1707 2340 1708
rect 2438 1712 2444 1713
rect 2438 1708 2439 1712
rect 2443 1708 2444 1712
rect 2502 1711 2503 1715
rect 2507 1711 2508 1715
rect 2502 1710 2508 1711
rect 2438 1707 2444 1708
rect 1350 1700 1356 1701
rect 1326 1697 1332 1698
rect 1326 1693 1327 1697
rect 1331 1693 1332 1697
rect 1350 1696 1351 1700
rect 1355 1696 1356 1700
rect 1350 1695 1356 1696
rect 1430 1700 1436 1701
rect 1430 1696 1431 1700
rect 1435 1696 1436 1700
rect 1430 1695 1436 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1646 1700 1652 1701
rect 1646 1696 1647 1700
rect 1651 1696 1652 1700
rect 1646 1695 1652 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 2014 1700 2020 1701
rect 2014 1696 2015 1700
rect 2019 1696 2020 1700
rect 2014 1695 2020 1696
rect 2158 1700 2164 1701
rect 2158 1696 2159 1700
rect 2163 1696 2164 1700
rect 2158 1695 2164 1696
rect 2310 1700 2316 1701
rect 2310 1696 2311 1700
rect 2315 1696 2316 1700
rect 2310 1695 2316 1696
rect 2438 1700 2444 1701
rect 2438 1696 2439 1700
rect 2443 1696 2444 1700
rect 2438 1695 2444 1696
rect 2502 1697 2508 1698
rect 1326 1692 1332 1693
rect 2502 1693 2503 1697
rect 2507 1693 2508 1697
rect 2502 1692 2508 1693
rect 1326 1680 1332 1681
rect 2502 1680 2508 1681
rect 190 1677 196 1678
rect 110 1676 116 1677
rect 110 1672 111 1676
rect 115 1672 116 1676
rect 190 1673 191 1677
rect 195 1673 196 1677
rect 190 1672 196 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 350 1677 356 1678
rect 350 1673 351 1677
rect 355 1673 356 1677
rect 350 1672 356 1673
rect 438 1677 444 1678
rect 438 1673 439 1677
rect 443 1673 444 1677
rect 438 1672 444 1673
rect 534 1677 540 1678
rect 534 1673 535 1677
rect 539 1673 540 1677
rect 534 1672 540 1673
rect 638 1677 644 1678
rect 638 1673 639 1677
rect 643 1673 644 1677
rect 638 1672 644 1673
rect 742 1677 748 1678
rect 742 1673 743 1677
rect 747 1673 748 1677
rect 742 1672 748 1673
rect 846 1677 852 1678
rect 846 1673 847 1677
rect 851 1673 852 1677
rect 846 1672 852 1673
rect 950 1677 956 1678
rect 950 1673 951 1677
rect 955 1673 956 1677
rect 950 1672 956 1673
rect 1062 1677 1068 1678
rect 1062 1673 1063 1677
rect 1067 1673 1068 1677
rect 1062 1672 1068 1673
rect 1174 1677 1180 1678
rect 1174 1673 1175 1677
rect 1179 1673 1180 1677
rect 1174 1672 1180 1673
rect 1286 1676 1292 1677
rect 1286 1672 1287 1676
rect 1291 1672 1292 1676
rect 1326 1676 1327 1680
rect 1331 1676 1332 1680
rect 1326 1675 1332 1676
rect 1366 1679 1372 1680
rect 1366 1675 1367 1679
rect 1371 1675 1372 1679
rect 1366 1674 1372 1675
rect 1446 1679 1452 1680
rect 1446 1675 1447 1679
rect 1451 1675 1452 1679
rect 1446 1674 1452 1675
rect 1550 1679 1556 1680
rect 1550 1675 1551 1679
rect 1555 1675 1556 1679
rect 1550 1674 1556 1675
rect 1662 1679 1668 1680
rect 1662 1675 1663 1679
rect 1667 1675 1668 1679
rect 1662 1674 1668 1675
rect 1774 1679 1780 1680
rect 1774 1675 1775 1679
rect 1779 1675 1780 1679
rect 1774 1674 1780 1675
rect 1894 1679 1900 1680
rect 1894 1675 1895 1679
rect 1899 1675 1900 1679
rect 1894 1674 1900 1675
rect 2030 1679 2036 1680
rect 2030 1675 2031 1679
rect 2035 1675 2036 1679
rect 2030 1674 2036 1675
rect 2174 1679 2180 1680
rect 2174 1675 2175 1679
rect 2179 1675 2180 1679
rect 2174 1674 2180 1675
rect 2326 1679 2332 1680
rect 2326 1675 2327 1679
rect 2331 1675 2332 1679
rect 2326 1674 2332 1675
rect 2454 1679 2460 1680
rect 2454 1675 2455 1679
rect 2459 1675 2460 1679
rect 2502 1676 2503 1680
rect 2507 1676 2508 1680
rect 2502 1675 2508 1676
rect 2454 1674 2460 1675
rect 110 1671 116 1672
rect 1286 1671 1292 1672
rect 110 1659 116 1660
rect 110 1655 111 1659
rect 115 1655 116 1659
rect 1286 1659 1292 1660
rect 110 1654 116 1655
rect 174 1656 180 1657
rect 174 1652 175 1656
rect 179 1652 180 1656
rect 174 1651 180 1652
rect 254 1656 260 1657
rect 254 1652 255 1656
rect 259 1652 260 1656
rect 254 1651 260 1652
rect 334 1656 340 1657
rect 334 1652 335 1656
rect 339 1652 340 1656
rect 334 1651 340 1652
rect 422 1656 428 1657
rect 422 1652 423 1656
rect 427 1652 428 1656
rect 422 1651 428 1652
rect 518 1656 524 1657
rect 518 1652 519 1656
rect 523 1652 524 1656
rect 518 1651 524 1652
rect 622 1656 628 1657
rect 622 1652 623 1656
rect 627 1652 628 1656
rect 622 1651 628 1652
rect 726 1656 732 1657
rect 726 1652 727 1656
rect 731 1652 732 1656
rect 726 1651 732 1652
rect 830 1656 836 1657
rect 830 1652 831 1656
rect 835 1652 836 1656
rect 830 1651 836 1652
rect 934 1656 940 1657
rect 934 1652 935 1656
rect 939 1652 940 1656
rect 934 1651 940 1652
rect 1046 1656 1052 1657
rect 1046 1652 1047 1656
rect 1051 1652 1052 1656
rect 1046 1651 1052 1652
rect 1158 1656 1164 1657
rect 1158 1652 1159 1656
rect 1163 1652 1164 1656
rect 1286 1655 1287 1659
rect 1291 1655 1292 1659
rect 1286 1654 1292 1655
rect 1158 1651 1164 1652
rect 214 1644 220 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 270 1644 276 1645
rect 270 1640 271 1644
rect 275 1640 276 1644
rect 270 1639 276 1640
rect 334 1644 340 1645
rect 334 1640 335 1644
rect 339 1640 340 1644
rect 334 1639 340 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 478 1644 484 1645
rect 478 1640 479 1644
rect 483 1640 484 1644
rect 478 1639 484 1640
rect 558 1644 564 1645
rect 558 1640 559 1644
rect 563 1640 564 1644
rect 558 1639 564 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 742 1644 748 1645
rect 742 1640 743 1644
rect 747 1640 748 1644
rect 742 1639 748 1640
rect 838 1644 844 1645
rect 838 1640 839 1644
rect 843 1640 844 1644
rect 838 1639 844 1640
rect 942 1644 948 1645
rect 942 1640 943 1644
rect 947 1640 948 1644
rect 942 1639 948 1640
rect 1054 1644 1060 1645
rect 1054 1640 1055 1644
rect 1059 1640 1060 1644
rect 1054 1639 1060 1640
rect 1174 1644 1180 1645
rect 1174 1640 1175 1644
rect 1179 1640 1180 1644
rect 1174 1639 1180 1640
rect 1286 1641 1292 1642
rect 110 1636 116 1637
rect 1286 1637 1287 1641
rect 1291 1637 1292 1641
rect 1286 1636 1292 1637
rect 110 1624 116 1625
rect 1286 1624 1292 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 230 1623 236 1624
rect 230 1619 231 1623
rect 235 1619 236 1623
rect 230 1618 236 1619
rect 286 1623 292 1624
rect 286 1619 287 1623
rect 291 1619 292 1623
rect 286 1618 292 1619
rect 350 1623 356 1624
rect 350 1619 351 1623
rect 355 1619 356 1623
rect 350 1618 356 1619
rect 422 1623 428 1624
rect 422 1619 423 1623
rect 427 1619 428 1623
rect 422 1618 428 1619
rect 494 1623 500 1624
rect 494 1619 495 1623
rect 499 1619 500 1623
rect 494 1618 500 1619
rect 574 1623 580 1624
rect 574 1619 575 1623
rect 579 1619 580 1623
rect 574 1618 580 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 758 1623 764 1624
rect 758 1619 759 1623
rect 763 1619 764 1623
rect 758 1618 764 1619
rect 854 1623 860 1624
rect 854 1619 855 1623
rect 859 1619 860 1623
rect 854 1618 860 1619
rect 958 1623 964 1624
rect 958 1619 959 1623
rect 963 1619 964 1623
rect 958 1618 964 1619
rect 1070 1623 1076 1624
rect 1070 1619 1071 1623
rect 1075 1619 1076 1623
rect 1070 1618 1076 1619
rect 1190 1623 1196 1624
rect 1190 1619 1191 1623
rect 1195 1619 1196 1623
rect 1286 1620 1287 1624
rect 1291 1620 1292 1624
rect 1366 1621 1372 1622
rect 1286 1619 1292 1620
rect 1326 1620 1332 1621
rect 1190 1618 1196 1619
rect 1326 1616 1327 1620
rect 1331 1616 1332 1620
rect 1366 1617 1367 1621
rect 1371 1617 1372 1621
rect 1366 1616 1372 1617
rect 1430 1621 1436 1622
rect 1430 1617 1431 1621
rect 1435 1617 1436 1621
rect 1430 1616 1436 1617
rect 1518 1621 1524 1622
rect 1518 1617 1519 1621
rect 1523 1617 1524 1621
rect 1518 1616 1524 1617
rect 1598 1621 1604 1622
rect 1598 1617 1599 1621
rect 1603 1617 1604 1621
rect 1598 1616 1604 1617
rect 1678 1621 1684 1622
rect 1678 1617 1679 1621
rect 1683 1617 1684 1621
rect 1678 1616 1684 1617
rect 1750 1621 1756 1622
rect 1750 1617 1751 1621
rect 1755 1617 1756 1621
rect 1750 1616 1756 1617
rect 1838 1621 1844 1622
rect 1838 1617 1839 1621
rect 1843 1617 1844 1621
rect 1838 1616 1844 1617
rect 1934 1621 1940 1622
rect 1934 1617 1935 1621
rect 1939 1617 1940 1621
rect 1934 1616 1940 1617
rect 2054 1621 2060 1622
rect 2054 1617 2055 1621
rect 2059 1617 2060 1621
rect 2054 1616 2060 1617
rect 2182 1621 2188 1622
rect 2182 1617 2183 1621
rect 2187 1617 2188 1621
rect 2182 1616 2188 1617
rect 2326 1621 2332 1622
rect 2326 1617 2327 1621
rect 2331 1617 2332 1621
rect 2326 1616 2332 1617
rect 2454 1621 2460 1622
rect 2454 1617 2455 1621
rect 2459 1617 2460 1621
rect 2454 1616 2460 1617
rect 2502 1620 2508 1621
rect 2502 1616 2503 1620
rect 2507 1616 2508 1620
rect 1326 1615 1332 1616
rect 2502 1615 2508 1616
rect 1326 1603 1332 1604
rect 1326 1599 1327 1603
rect 1331 1599 1332 1603
rect 2502 1603 2508 1604
rect 1326 1598 1332 1599
rect 1350 1600 1356 1601
rect 1350 1596 1351 1600
rect 1355 1596 1356 1600
rect 1350 1595 1356 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1502 1600 1508 1601
rect 1502 1596 1503 1600
rect 1507 1596 1508 1600
rect 1502 1595 1508 1596
rect 1582 1600 1588 1601
rect 1582 1596 1583 1600
rect 1587 1596 1588 1600
rect 1582 1595 1588 1596
rect 1662 1600 1668 1601
rect 1662 1596 1663 1600
rect 1667 1596 1668 1600
rect 1662 1595 1668 1596
rect 1734 1600 1740 1601
rect 1734 1596 1735 1600
rect 1739 1596 1740 1600
rect 1734 1595 1740 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1918 1600 1924 1601
rect 1918 1596 1919 1600
rect 1923 1596 1924 1600
rect 1918 1595 1924 1596
rect 2038 1600 2044 1601
rect 2038 1596 2039 1600
rect 2043 1596 2044 1600
rect 2038 1595 2044 1596
rect 2166 1600 2172 1601
rect 2166 1596 2167 1600
rect 2171 1596 2172 1600
rect 2166 1595 2172 1596
rect 2310 1600 2316 1601
rect 2310 1596 2311 1600
rect 2315 1596 2316 1600
rect 2310 1595 2316 1596
rect 2438 1600 2444 1601
rect 2438 1596 2439 1600
rect 2443 1596 2444 1600
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2438 1595 2444 1596
rect 1350 1584 1356 1585
rect 1326 1581 1332 1582
rect 1326 1577 1327 1581
rect 1331 1577 1332 1581
rect 1350 1580 1351 1584
rect 1355 1580 1356 1584
rect 1350 1579 1356 1580
rect 1422 1584 1428 1585
rect 1422 1580 1423 1584
rect 1427 1580 1428 1584
rect 1422 1579 1428 1580
rect 1526 1584 1532 1585
rect 1526 1580 1527 1584
rect 1531 1580 1532 1584
rect 1526 1579 1532 1580
rect 1646 1584 1652 1585
rect 1646 1580 1647 1584
rect 1651 1580 1652 1584
rect 1646 1579 1652 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1934 1584 1940 1585
rect 1934 1580 1935 1584
rect 1939 1580 1940 1584
rect 1934 1579 1940 1580
rect 2102 1584 2108 1585
rect 2102 1580 2103 1584
rect 2107 1580 2108 1584
rect 2102 1579 2108 1580
rect 2278 1584 2284 1585
rect 2278 1580 2279 1584
rect 2283 1580 2284 1584
rect 2278 1579 2284 1580
rect 2438 1584 2444 1585
rect 2438 1580 2439 1584
rect 2443 1580 2444 1584
rect 2438 1579 2444 1580
rect 2502 1581 2508 1582
rect 1326 1576 1332 1577
rect 2502 1577 2503 1581
rect 2507 1577 2508 1581
rect 2502 1576 2508 1577
rect 286 1573 292 1574
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 286 1569 287 1573
rect 291 1569 292 1573
rect 286 1568 292 1569
rect 350 1573 356 1574
rect 350 1569 351 1573
rect 355 1569 356 1573
rect 350 1568 356 1569
rect 422 1573 428 1574
rect 422 1569 423 1573
rect 427 1569 428 1573
rect 422 1568 428 1569
rect 502 1573 508 1574
rect 502 1569 503 1573
rect 507 1569 508 1573
rect 502 1568 508 1569
rect 598 1573 604 1574
rect 598 1569 599 1573
rect 603 1569 604 1573
rect 598 1568 604 1569
rect 702 1573 708 1574
rect 702 1569 703 1573
rect 707 1569 708 1573
rect 702 1568 708 1569
rect 814 1573 820 1574
rect 814 1569 815 1573
rect 819 1569 820 1573
rect 814 1568 820 1569
rect 934 1573 940 1574
rect 934 1569 935 1573
rect 939 1569 940 1573
rect 934 1568 940 1569
rect 1062 1573 1068 1574
rect 1062 1569 1063 1573
rect 1067 1569 1068 1573
rect 1062 1568 1068 1569
rect 1190 1573 1196 1574
rect 1190 1569 1191 1573
rect 1195 1569 1196 1573
rect 1190 1568 1196 1569
rect 1286 1572 1292 1573
rect 1286 1568 1287 1572
rect 1291 1568 1292 1572
rect 110 1567 116 1568
rect 1286 1567 1292 1568
rect 1326 1564 1332 1565
rect 2502 1564 2508 1565
rect 1326 1560 1327 1564
rect 1331 1560 1332 1564
rect 1326 1559 1332 1560
rect 1366 1563 1372 1564
rect 1366 1559 1367 1563
rect 1371 1559 1372 1563
rect 1366 1558 1372 1559
rect 1438 1563 1444 1564
rect 1438 1559 1439 1563
rect 1443 1559 1444 1563
rect 1438 1558 1444 1559
rect 1542 1563 1548 1564
rect 1542 1559 1543 1563
rect 1547 1559 1548 1563
rect 1542 1558 1548 1559
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1559 1668 1563
rect 1662 1558 1668 1559
rect 1798 1563 1804 1564
rect 1798 1559 1799 1563
rect 1803 1559 1804 1563
rect 1798 1558 1804 1559
rect 1950 1563 1956 1564
rect 1950 1559 1951 1563
rect 1955 1559 1956 1563
rect 1950 1558 1956 1559
rect 2118 1563 2124 1564
rect 2118 1559 2119 1563
rect 2123 1559 2124 1563
rect 2118 1558 2124 1559
rect 2294 1563 2300 1564
rect 2294 1559 2295 1563
rect 2299 1559 2300 1563
rect 2294 1558 2300 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2502 1560 2503 1564
rect 2507 1560 2508 1564
rect 2502 1559 2508 1560
rect 2454 1558 2460 1559
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1286 1555 1292 1556
rect 110 1550 116 1551
rect 270 1552 276 1553
rect 270 1548 271 1552
rect 275 1548 276 1552
rect 270 1547 276 1548
rect 334 1552 340 1553
rect 334 1548 335 1552
rect 339 1548 340 1552
rect 334 1547 340 1548
rect 406 1552 412 1553
rect 406 1548 407 1552
rect 411 1548 412 1552
rect 406 1547 412 1548
rect 486 1552 492 1553
rect 486 1548 487 1552
rect 491 1548 492 1552
rect 486 1547 492 1548
rect 582 1552 588 1553
rect 582 1548 583 1552
rect 587 1548 588 1552
rect 582 1547 588 1548
rect 686 1552 692 1553
rect 686 1548 687 1552
rect 691 1548 692 1552
rect 686 1547 692 1548
rect 798 1552 804 1553
rect 798 1548 799 1552
rect 803 1548 804 1552
rect 798 1547 804 1548
rect 918 1552 924 1553
rect 918 1548 919 1552
rect 923 1548 924 1552
rect 918 1547 924 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1174 1552 1180 1553
rect 1174 1548 1175 1552
rect 1179 1548 1180 1552
rect 1286 1551 1287 1555
rect 1291 1551 1292 1555
rect 1286 1550 1292 1551
rect 1174 1547 1180 1548
rect 470 1532 476 1533
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 470 1528 471 1532
rect 475 1528 476 1532
rect 470 1527 476 1528
rect 550 1532 556 1533
rect 550 1528 551 1532
rect 555 1528 556 1532
rect 550 1527 556 1528
rect 638 1532 644 1533
rect 638 1528 639 1532
rect 643 1528 644 1532
rect 638 1527 644 1528
rect 734 1532 740 1533
rect 734 1528 735 1532
rect 739 1528 740 1532
rect 734 1527 740 1528
rect 838 1532 844 1533
rect 838 1528 839 1532
rect 843 1528 844 1532
rect 838 1527 844 1528
rect 950 1532 956 1533
rect 950 1528 951 1532
rect 955 1528 956 1532
rect 950 1527 956 1528
rect 1062 1532 1068 1533
rect 1062 1528 1063 1532
rect 1067 1528 1068 1532
rect 1062 1527 1068 1528
rect 1174 1532 1180 1533
rect 1174 1528 1175 1532
rect 1179 1528 1180 1532
rect 1174 1527 1180 1528
rect 1286 1529 1292 1530
rect 110 1524 116 1525
rect 1286 1525 1287 1529
rect 1291 1525 1292 1529
rect 1286 1524 1292 1525
rect 1366 1513 1372 1514
rect 110 1512 116 1513
rect 1286 1512 1292 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 486 1511 492 1512
rect 486 1507 487 1511
rect 491 1507 492 1511
rect 486 1506 492 1507
rect 566 1511 572 1512
rect 566 1507 567 1511
rect 571 1507 572 1511
rect 566 1506 572 1507
rect 654 1511 660 1512
rect 654 1507 655 1511
rect 659 1507 660 1511
rect 654 1506 660 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 854 1511 860 1512
rect 854 1507 855 1511
rect 859 1507 860 1511
rect 854 1506 860 1507
rect 966 1511 972 1512
rect 966 1507 967 1511
rect 971 1507 972 1511
rect 966 1506 972 1507
rect 1078 1511 1084 1512
rect 1078 1507 1079 1511
rect 1083 1507 1084 1511
rect 1078 1506 1084 1507
rect 1190 1511 1196 1512
rect 1190 1507 1191 1511
rect 1195 1507 1196 1511
rect 1286 1508 1287 1512
rect 1291 1508 1292 1512
rect 1286 1507 1292 1508
rect 1326 1512 1332 1513
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1366 1509 1367 1513
rect 1371 1509 1372 1513
rect 1366 1508 1372 1509
rect 1438 1513 1444 1514
rect 1438 1509 1439 1513
rect 1443 1509 1444 1513
rect 1438 1508 1444 1509
rect 1542 1513 1548 1514
rect 1542 1509 1543 1513
rect 1547 1509 1548 1513
rect 1542 1508 1548 1509
rect 1646 1513 1652 1514
rect 1646 1509 1647 1513
rect 1651 1509 1652 1513
rect 1646 1508 1652 1509
rect 1750 1513 1756 1514
rect 1750 1509 1751 1513
rect 1755 1509 1756 1513
rect 1750 1508 1756 1509
rect 1854 1513 1860 1514
rect 1854 1509 1855 1513
rect 1859 1509 1860 1513
rect 1854 1508 1860 1509
rect 1958 1513 1964 1514
rect 1958 1509 1959 1513
rect 1963 1509 1964 1513
rect 1958 1508 1964 1509
rect 2054 1513 2060 1514
rect 2054 1509 2055 1513
rect 2059 1509 2060 1513
rect 2054 1508 2060 1509
rect 2150 1513 2156 1514
rect 2150 1509 2151 1513
rect 2155 1509 2156 1513
rect 2150 1508 2156 1509
rect 2246 1513 2252 1514
rect 2246 1509 2247 1513
rect 2251 1509 2252 1513
rect 2246 1508 2252 1509
rect 2342 1513 2348 1514
rect 2342 1509 2343 1513
rect 2347 1509 2348 1513
rect 2342 1508 2348 1509
rect 2438 1513 2444 1514
rect 2438 1509 2439 1513
rect 2443 1509 2444 1513
rect 2438 1508 2444 1509
rect 2502 1512 2508 1513
rect 2502 1508 2503 1512
rect 2507 1508 2508 1512
rect 1326 1507 1332 1508
rect 2502 1507 2508 1508
rect 1190 1506 1196 1507
rect 1326 1495 1332 1496
rect 1326 1491 1327 1495
rect 1331 1491 1332 1495
rect 2502 1495 2508 1496
rect 1326 1490 1332 1491
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1422 1492 1428 1493
rect 1422 1488 1423 1492
rect 1427 1488 1428 1492
rect 1422 1487 1428 1488
rect 1526 1492 1532 1493
rect 1526 1488 1527 1492
rect 1531 1488 1532 1492
rect 1526 1487 1532 1488
rect 1630 1492 1636 1493
rect 1630 1488 1631 1492
rect 1635 1488 1636 1492
rect 1630 1487 1636 1488
rect 1734 1492 1740 1493
rect 1734 1488 1735 1492
rect 1739 1488 1740 1492
rect 1734 1487 1740 1488
rect 1838 1492 1844 1493
rect 1838 1488 1839 1492
rect 1843 1488 1844 1492
rect 1838 1487 1844 1488
rect 1942 1492 1948 1493
rect 1942 1488 1943 1492
rect 1947 1488 1948 1492
rect 1942 1487 1948 1488
rect 2038 1492 2044 1493
rect 2038 1488 2039 1492
rect 2043 1488 2044 1492
rect 2038 1487 2044 1488
rect 2134 1492 2140 1493
rect 2134 1488 2135 1492
rect 2139 1488 2140 1492
rect 2134 1487 2140 1488
rect 2230 1492 2236 1493
rect 2230 1488 2231 1492
rect 2235 1488 2236 1492
rect 2230 1487 2236 1488
rect 2326 1492 2332 1493
rect 2326 1488 2327 1492
rect 2331 1488 2332 1492
rect 2326 1487 2332 1488
rect 2422 1492 2428 1493
rect 2422 1488 2423 1492
rect 2427 1488 2428 1492
rect 2502 1491 2503 1495
rect 2507 1491 2508 1495
rect 2502 1490 2508 1491
rect 2422 1487 2428 1488
rect 1350 1476 1356 1477
rect 1326 1473 1332 1474
rect 1326 1469 1327 1473
rect 1331 1469 1332 1473
rect 1350 1472 1351 1476
rect 1355 1472 1356 1476
rect 1350 1471 1356 1472
rect 1422 1476 1428 1477
rect 1422 1472 1423 1476
rect 1427 1472 1428 1476
rect 1422 1471 1428 1472
rect 1518 1476 1524 1477
rect 1518 1472 1519 1476
rect 1523 1472 1524 1476
rect 1518 1471 1524 1472
rect 1614 1476 1620 1477
rect 1614 1472 1615 1476
rect 1619 1472 1620 1476
rect 1614 1471 1620 1472
rect 1710 1476 1716 1477
rect 1710 1472 1711 1476
rect 1715 1472 1716 1476
rect 1710 1471 1716 1472
rect 1814 1476 1820 1477
rect 1814 1472 1815 1476
rect 1819 1472 1820 1476
rect 1814 1471 1820 1472
rect 1926 1476 1932 1477
rect 1926 1472 1927 1476
rect 1931 1472 1932 1476
rect 1926 1471 1932 1472
rect 2046 1476 2052 1477
rect 2046 1472 2047 1476
rect 2051 1472 2052 1476
rect 2046 1471 2052 1472
rect 2174 1476 2180 1477
rect 2174 1472 2175 1476
rect 2179 1472 2180 1476
rect 2174 1471 2180 1472
rect 2302 1476 2308 1477
rect 2302 1472 2303 1476
rect 2307 1472 2308 1476
rect 2302 1471 2308 1472
rect 2438 1476 2444 1477
rect 2438 1472 2439 1476
rect 2443 1472 2444 1476
rect 2438 1471 2444 1472
rect 2502 1473 2508 1474
rect 1326 1468 1332 1469
rect 2502 1469 2503 1473
rect 2507 1469 2508 1473
rect 2502 1468 2508 1469
rect 374 1461 380 1462
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 374 1457 375 1461
rect 379 1457 380 1461
rect 374 1456 380 1457
rect 462 1461 468 1462
rect 462 1457 463 1461
rect 467 1457 468 1461
rect 462 1456 468 1457
rect 558 1461 564 1462
rect 558 1457 559 1461
rect 563 1457 564 1461
rect 558 1456 564 1457
rect 654 1461 660 1462
rect 654 1457 655 1461
rect 659 1457 660 1461
rect 654 1456 660 1457
rect 750 1461 756 1462
rect 750 1457 751 1461
rect 755 1457 756 1461
rect 750 1456 756 1457
rect 854 1461 860 1462
rect 854 1457 855 1461
rect 859 1457 860 1461
rect 854 1456 860 1457
rect 958 1461 964 1462
rect 958 1457 959 1461
rect 963 1457 964 1461
rect 958 1456 964 1457
rect 1062 1461 1068 1462
rect 1062 1457 1063 1461
rect 1067 1457 1068 1461
rect 1062 1456 1068 1457
rect 1166 1461 1172 1462
rect 1166 1457 1167 1461
rect 1171 1457 1172 1461
rect 1166 1456 1172 1457
rect 1286 1460 1292 1461
rect 1286 1456 1287 1460
rect 1291 1456 1292 1460
rect 110 1455 116 1456
rect 1286 1455 1292 1456
rect 1326 1456 1332 1457
rect 2502 1456 2508 1457
rect 1326 1452 1327 1456
rect 1331 1452 1332 1456
rect 1326 1451 1332 1452
rect 1366 1455 1372 1456
rect 1366 1451 1367 1455
rect 1371 1451 1372 1455
rect 1366 1450 1372 1451
rect 1438 1455 1444 1456
rect 1438 1451 1439 1455
rect 1443 1451 1444 1455
rect 1438 1450 1444 1451
rect 1534 1455 1540 1456
rect 1534 1451 1535 1455
rect 1539 1451 1540 1455
rect 1534 1450 1540 1451
rect 1630 1455 1636 1456
rect 1630 1451 1631 1455
rect 1635 1451 1636 1455
rect 1630 1450 1636 1451
rect 1726 1455 1732 1456
rect 1726 1451 1727 1455
rect 1731 1451 1732 1455
rect 1726 1450 1732 1451
rect 1830 1455 1836 1456
rect 1830 1451 1831 1455
rect 1835 1451 1836 1455
rect 1830 1450 1836 1451
rect 1942 1455 1948 1456
rect 1942 1451 1943 1455
rect 1947 1451 1948 1455
rect 1942 1450 1948 1451
rect 2062 1455 2068 1456
rect 2062 1451 2063 1455
rect 2067 1451 2068 1455
rect 2062 1450 2068 1451
rect 2190 1455 2196 1456
rect 2190 1451 2191 1455
rect 2195 1451 2196 1455
rect 2190 1450 2196 1451
rect 2318 1455 2324 1456
rect 2318 1451 2319 1455
rect 2323 1451 2324 1455
rect 2318 1450 2324 1451
rect 2454 1455 2460 1456
rect 2454 1451 2455 1455
rect 2459 1451 2460 1455
rect 2502 1452 2503 1456
rect 2507 1452 2508 1456
rect 2502 1451 2508 1452
rect 2454 1450 2460 1451
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 1286 1443 1292 1444
rect 110 1438 116 1439
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 446 1440 452 1441
rect 446 1436 447 1440
rect 451 1436 452 1440
rect 446 1435 452 1436
rect 542 1440 548 1441
rect 542 1436 543 1440
rect 547 1436 548 1440
rect 542 1435 548 1436
rect 638 1440 644 1441
rect 638 1436 639 1440
rect 643 1436 644 1440
rect 638 1435 644 1436
rect 734 1440 740 1441
rect 734 1436 735 1440
rect 739 1436 740 1440
rect 734 1435 740 1436
rect 838 1440 844 1441
rect 838 1436 839 1440
rect 843 1436 844 1440
rect 838 1435 844 1436
rect 942 1440 948 1441
rect 942 1436 943 1440
rect 947 1436 948 1440
rect 942 1435 948 1436
rect 1046 1440 1052 1441
rect 1046 1436 1047 1440
rect 1051 1436 1052 1440
rect 1046 1435 1052 1436
rect 1150 1440 1156 1441
rect 1150 1436 1151 1440
rect 1155 1436 1156 1440
rect 1286 1439 1287 1443
rect 1291 1439 1292 1443
rect 1286 1438 1292 1439
rect 1150 1435 1156 1436
rect 230 1428 236 1429
rect 110 1425 116 1426
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 230 1424 231 1428
rect 235 1424 236 1428
rect 230 1423 236 1424
rect 318 1428 324 1429
rect 318 1424 319 1428
rect 323 1424 324 1428
rect 318 1423 324 1424
rect 414 1428 420 1429
rect 414 1424 415 1428
rect 419 1424 420 1428
rect 414 1423 420 1424
rect 510 1428 516 1429
rect 510 1424 511 1428
rect 515 1424 516 1428
rect 510 1423 516 1424
rect 614 1428 620 1429
rect 614 1424 615 1428
rect 619 1424 620 1428
rect 614 1423 620 1424
rect 710 1428 716 1429
rect 710 1424 711 1428
rect 715 1424 716 1428
rect 710 1423 716 1424
rect 806 1428 812 1429
rect 806 1424 807 1428
rect 811 1424 812 1428
rect 806 1423 812 1424
rect 894 1428 900 1429
rect 894 1424 895 1428
rect 899 1424 900 1428
rect 894 1423 900 1424
rect 990 1428 996 1429
rect 990 1424 991 1428
rect 995 1424 996 1428
rect 990 1423 996 1424
rect 1086 1428 1092 1429
rect 1086 1424 1087 1428
rect 1091 1424 1092 1428
rect 1086 1423 1092 1424
rect 1286 1425 1292 1426
rect 110 1420 116 1421
rect 1286 1421 1287 1425
rect 1291 1421 1292 1425
rect 1286 1420 1292 1421
rect 110 1408 116 1409
rect 1286 1408 1292 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 246 1407 252 1408
rect 246 1403 247 1407
rect 251 1403 252 1407
rect 246 1402 252 1403
rect 334 1407 340 1408
rect 334 1403 335 1407
rect 339 1403 340 1407
rect 334 1402 340 1403
rect 430 1407 436 1408
rect 430 1403 431 1407
rect 435 1403 436 1407
rect 430 1402 436 1403
rect 526 1407 532 1408
rect 526 1403 527 1407
rect 531 1403 532 1407
rect 526 1402 532 1403
rect 630 1407 636 1408
rect 630 1403 631 1407
rect 635 1403 636 1407
rect 630 1402 636 1403
rect 726 1407 732 1408
rect 726 1403 727 1407
rect 731 1403 732 1407
rect 726 1402 732 1403
rect 822 1407 828 1408
rect 822 1403 823 1407
rect 827 1403 828 1407
rect 822 1402 828 1403
rect 910 1407 916 1408
rect 910 1403 911 1407
rect 915 1403 916 1407
rect 910 1402 916 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1102 1407 1108 1408
rect 1102 1403 1103 1407
rect 1107 1403 1108 1407
rect 1286 1404 1287 1408
rect 1291 1404 1292 1408
rect 1286 1403 1292 1404
rect 1102 1402 1108 1403
rect 1366 1401 1372 1402
rect 1326 1400 1332 1401
rect 1326 1396 1327 1400
rect 1331 1396 1332 1400
rect 1366 1397 1367 1401
rect 1371 1397 1372 1401
rect 1366 1396 1372 1397
rect 1422 1401 1428 1402
rect 1422 1397 1423 1401
rect 1427 1397 1428 1401
rect 1422 1396 1428 1397
rect 1502 1401 1508 1402
rect 1502 1397 1503 1401
rect 1507 1397 1508 1401
rect 1502 1396 1508 1397
rect 1590 1401 1596 1402
rect 1590 1397 1591 1401
rect 1595 1397 1596 1401
rect 1590 1396 1596 1397
rect 1678 1401 1684 1402
rect 1678 1397 1679 1401
rect 1683 1397 1684 1401
rect 1678 1396 1684 1397
rect 1774 1401 1780 1402
rect 1774 1397 1775 1401
rect 1779 1397 1780 1401
rect 1774 1396 1780 1397
rect 1878 1401 1884 1402
rect 1878 1397 1879 1401
rect 1883 1397 1884 1401
rect 1878 1396 1884 1397
rect 1990 1401 1996 1402
rect 1990 1397 1991 1401
rect 1995 1397 1996 1401
rect 1990 1396 1996 1397
rect 2110 1401 2116 1402
rect 2110 1397 2111 1401
rect 2115 1397 2116 1401
rect 2110 1396 2116 1397
rect 2230 1401 2236 1402
rect 2230 1397 2231 1401
rect 2235 1397 2236 1401
rect 2230 1396 2236 1397
rect 2350 1401 2356 1402
rect 2350 1397 2351 1401
rect 2355 1397 2356 1401
rect 2350 1396 2356 1397
rect 2454 1401 2460 1402
rect 2454 1397 2455 1401
rect 2459 1397 2460 1401
rect 2454 1396 2460 1397
rect 2502 1400 2508 1401
rect 2502 1396 2503 1400
rect 2507 1396 2508 1400
rect 1326 1395 1332 1396
rect 2502 1395 2508 1396
rect 1326 1383 1332 1384
rect 1326 1379 1327 1383
rect 1331 1379 1332 1383
rect 2502 1383 2508 1384
rect 1326 1378 1332 1379
rect 1350 1380 1356 1381
rect 1350 1376 1351 1380
rect 1355 1376 1356 1380
rect 1350 1375 1356 1376
rect 1406 1380 1412 1381
rect 1406 1376 1407 1380
rect 1411 1376 1412 1380
rect 1406 1375 1412 1376
rect 1486 1380 1492 1381
rect 1486 1376 1487 1380
rect 1491 1376 1492 1380
rect 1486 1375 1492 1376
rect 1574 1380 1580 1381
rect 1574 1376 1575 1380
rect 1579 1376 1580 1380
rect 1574 1375 1580 1376
rect 1662 1380 1668 1381
rect 1662 1376 1663 1380
rect 1667 1376 1668 1380
rect 1662 1375 1668 1376
rect 1758 1380 1764 1381
rect 1758 1376 1759 1380
rect 1763 1376 1764 1380
rect 1758 1375 1764 1376
rect 1862 1380 1868 1381
rect 1862 1376 1863 1380
rect 1867 1376 1868 1380
rect 1862 1375 1868 1376
rect 1974 1380 1980 1381
rect 1974 1376 1975 1380
rect 1979 1376 1980 1380
rect 1974 1375 1980 1376
rect 2094 1380 2100 1381
rect 2094 1376 2095 1380
rect 2099 1376 2100 1380
rect 2094 1375 2100 1376
rect 2214 1380 2220 1381
rect 2214 1376 2215 1380
rect 2219 1376 2220 1380
rect 2214 1375 2220 1376
rect 2334 1380 2340 1381
rect 2334 1376 2335 1380
rect 2339 1376 2340 1380
rect 2334 1375 2340 1376
rect 2438 1380 2444 1381
rect 2438 1376 2439 1380
rect 2443 1376 2444 1380
rect 2502 1379 2503 1383
rect 2507 1379 2508 1383
rect 2502 1378 2508 1379
rect 2438 1375 2444 1376
rect 1350 1364 1356 1365
rect 1326 1361 1332 1362
rect 150 1357 156 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 150 1353 151 1357
rect 155 1353 156 1357
rect 150 1352 156 1353
rect 214 1357 220 1358
rect 214 1353 215 1357
rect 219 1353 220 1357
rect 214 1352 220 1353
rect 310 1357 316 1358
rect 310 1353 311 1357
rect 315 1353 316 1357
rect 310 1352 316 1353
rect 406 1357 412 1358
rect 406 1353 407 1357
rect 411 1353 412 1357
rect 406 1352 412 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 606 1357 612 1358
rect 606 1353 607 1357
rect 611 1353 612 1357
rect 606 1352 612 1353
rect 702 1357 708 1358
rect 702 1353 703 1357
rect 707 1353 708 1357
rect 702 1352 708 1353
rect 798 1357 804 1358
rect 798 1353 799 1357
rect 803 1353 804 1357
rect 798 1352 804 1353
rect 894 1357 900 1358
rect 894 1353 895 1357
rect 899 1353 900 1357
rect 894 1352 900 1353
rect 998 1357 1004 1358
rect 1326 1357 1327 1361
rect 1331 1357 1332 1361
rect 1350 1360 1351 1364
rect 1355 1360 1356 1364
rect 1350 1359 1356 1360
rect 1406 1364 1412 1365
rect 1406 1360 1407 1364
rect 1411 1360 1412 1364
rect 1406 1359 1412 1360
rect 1478 1364 1484 1365
rect 1478 1360 1479 1364
rect 1483 1360 1484 1364
rect 1478 1359 1484 1360
rect 1566 1364 1572 1365
rect 1566 1360 1567 1364
rect 1571 1360 1572 1364
rect 1566 1359 1572 1360
rect 1654 1364 1660 1365
rect 1654 1360 1655 1364
rect 1659 1360 1660 1364
rect 1654 1359 1660 1360
rect 1750 1364 1756 1365
rect 1750 1360 1751 1364
rect 1755 1360 1756 1364
rect 1750 1359 1756 1360
rect 1854 1364 1860 1365
rect 1854 1360 1855 1364
rect 1859 1360 1860 1364
rect 1854 1359 1860 1360
rect 1966 1364 1972 1365
rect 1966 1360 1967 1364
rect 1971 1360 1972 1364
rect 1966 1359 1972 1360
rect 2078 1364 2084 1365
rect 2078 1360 2079 1364
rect 2083 1360 2084 1364
rect 2078 1359 2084 1360
rect 2198 1364 2204 1365
rect 2198 1360 2199 1364
rect 2203 1360 2204 1364
rect 2198 1359 2204 1360
rect 2326 1364 2332 1365
rect 2326 1360 2327 1364
rect 2331 1360 2332 1364
rect 2326 1359 2332 1360
rect 2438 1364 2444 1365
rect 2438 1360 2439 1364
rect 2443 1360 2444 1364
rect 2438 1359 2444 1360
rect 2502 1361 2508 1362
rect 998 1353 999 1357
rect 1003 1353 1004 1357
rect 998 1352 1004 1353
rect 1286 1356 1292 1357
rect 1326 1356 1332 1357
rect 2502 1357 2503 1361
rect 2507 1357 2508 1361
rect 2502 1356 2508 1357
rect 1286 1352 1287 1356
rect 1291 1352 1292 1356
rect 110 1351 116 1352
rect 1286 1351 1292 1352
rect 1326 1344 1332 1345
rect 2502 1344 2508 1345
rect 1326 1340 1327 1344
rect 1331 1340 1332 1344
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 1286 1339 1292 1340
rect 1326 1339 1332 1340
rect 1366 1343 1372 1344
rect 1366 1339 1367 1343
rect 1371 1339 1372 1343
rect 110 1334 116 1335
rect 134 1336 140 1337
rect 134 1332 135 1336
rect 139 1332 140 1336
rect 134 1331 140 1332
rect 198 1336 204 1337
rect 198 1332 199 1336
rect 203 1332 204 1336
rect 198 1331 204 1332
rect 294 1336 300 1337
rect 294 1332 295 1336
rect 299 1332 300 1336
rect 294 1331 300 1332
rect 390 1336 396 1337
rect 390 1332 391 1336
rect 395 1332 396 1336
rect 390 1331 396 1332
rect 494 1336 500 1337
rect 494 1332 495 1336
rect 499 1332 500 1336
rect 494 1331 500 1332
rect 590 1336 596 1337
rect 590 1332 591 1336
rect 595 1332 596 1336
rect 590 1331 596 1332
rect 686 1336 692 1337
rect 686 1332 687 1336
rect 691 1332 692 1336
rect 686 1331 692 1332
rect 782 1336 788 1337
rect 782 1332 783 1336
rect 787 1332 788 1336
rect 782 1331 788 1332
rect 878 1336 884 1337
rect 878 1332 879 1336
rect 883 1332 884 1336
rect 878 1331 884 1332
rect 982 1336 988 1337
rect 982 1332 983 1336
rect 987 1332 988 1336
rect 1286 1335 1287 1339
rect 1291 1335 1292 1339
rect 1366 1338 1372 1339
rect 1422 1343 1428 1344
rect 1422 1339 1423 1343
rect 1427 1339 1428 1343
rect 1422 1338 1428 1339
rect 1494 1343 1500 1344
rect 1494 1339 1495 1343
rect 1499 1339 1500 1343
rect 1494 1338 1500 1339
rect 1582 1343 1588 1344
rect 1582 1339 1583 1343
rect 1587 1339 1588 1343
rect 1582 1338 1588 1339
rect 1670 1343 1676 1344
rect 1670 1339 1671 1343
rect 1675 1339 1676 1343
rect 1670 1338 1676 1339
rect 1766 1343 1772 1344
rect 1766 1339 1767 1343
rect 1771 1339 1772 1343
rect 1766 1338 1772 1339
rect 1870 1343 1876 1344
rect 1870 1339 1871 1343
rect 1875 1339 1876 1343
rect 1870 1338 1876 1339
rect 1982 1343 1988 1344
rect 1982 1339 1983 1343
rect 1987 1339 1988 1343
rect 1982 1338 1988 1339
rect 2094 1343 2100 1344
rect 2094 1339 2095 1343
rect 2099 1339 2100 1343
rect 2094 1338 2100 1339
rect 2214 1343 2220 1344
rect 2214 1339 2215 1343
rect 2219 1339 2220 1343
rect 2214 1338 2220 1339
rect 2342 1343 2348 1344
rect 2342 1339 2343 1343
rect 2347 1339 2348 1343
rect 2342 1338 2348 1339
rect 2454 1343 2460 1344
rect 2454 1339 2455 1343
rect 2459 1339 2460 1343
rect 2502 1340 2503 1344
rect 2507 1340 2508 1344
rect 2502 1339 2508 1340
rect 2454 1338 2460 1339
rect 1286 1334 1292 1335
rect 982 1331 988 1332
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 414 1324 420 1325
rect 414 1320 415 1324
rect 419 1320 420 1324
rect 414 1319 420 1320
rect 510 1324 516 1325
rect 510 1320 511 1324
rect 515 1320 516 1324
rect 510 1319 516 1320
rect 598 1324 604 1325
rect 598 1320 599 1324
rect 603 1320 604 1324
rect 598 1319 604 1320
rect 686 1324 692 1325
rect 686 1320 687 1324
rect 691 1320 692 1324
rect 686 1319 692 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 878 1324 884 1325
rect 878 1320 879 1324
rect 883 1320 884 1324
rect 878 1319 884 1320
rect 1286 1321 1292 1322
rect 110 1316 116 1317
rect 1286 1317 1287 1321
rect 1291 1317 1292 1321
rect 1286 1316 1292 1317
rect 110 1304 116 1305
rect 1286 1304 1292 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 150 1303 156 1304
rect 150 1299 151 1303
rect 155 1299 156 1303
rect 150 1298 156 1299
rect 230 1303 236 1304
rect 230 1299 231 1303
rect 235 1299 236 1303
rect 230 1298 236 1299
rect 334 1303 340 1304
rect 334 1299 335 1303
rect 339 1299 340 1303
rect 334 1298 340 1299
rect 430 1303 436 1304
rect 430 1299 431 1303
rect 435 1299 436 1303
rect 430 1298 436 1299
rect 526 1303 532 1304
rect 526 1299 527 1303
rect 531 1299 532 1303
rect 526 1298 532 1299
rect 614 1303 620 1304
rect 614 1299 615 1303
rect 619 1299 620 1303
rect 614 1298 620 1299
rect 702 1303 708 1304
rect 702 1299 703 1303
rect 707 1299 708 1303
rect 702 1298 708 1299
rect 798 1303 804 1304
rect 798 1299 799 1303
rect 803 1299 804 1303
rect 798 1298 804 1299
rect 894 1303 900 1304
rect 894 1299 895 1303
rect 899 1299 900 1303
rect 1286 1300 1287 1304
rect 1291 1300 1292 1304
rect 1286 1299 1292 1300
rect 894 1298 900 1299
rect 1366 1285 1372 1286
rect 1326 1284 1332 1285
rect 1326 1280 1327 1284
rect 1331 1280 1332 1284
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 1422 1285 1428 1286
rect 1422 1281 1423 1285
rect 1427 1281 1428 1285
rect 1422 1280 1428 1281
rect 1518 1285 1524 1286
rect 1518 1281 1519 1285
rect 1523 1281 1524 1285
rect 1518 1280 1524 1281
rect 1614 1285 1620 1286
rect 1614 1281 1615 1285
rect 1619 1281 1620 1285
rect 1614 1280 1620 1281
rect 1718 1285 1724 1286
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1718 1280 1724 1281
rect 1822 1285 1828 1286
rect 1822 1281 1823 1285
rect 1827 1281 1828 1285
rect 1822 1280 1828 1281
rect 1918 1285 1924 1286
rect 1918 1281 1919 1285
rect 1923 1281 1924 1285
rect 1918 1280 1924 1281
rect 2014 1285 2020 1286
rect 2014 1281 2015 1285
rect 2019 1281 2020 1285
rect 2014 1280 2020 1281
rect 2102 1285 2108 1286
rect 2102 1281 2103 1285
rect 2107 1281 2108 1285
rect 2102 1280 2108 1281
rect 2182 1285 2188 1286
rect 2182 1281 2183 1285
rect 2187 1281 2188 1285
rect 2182 1280 2188 1281
rect 2254 1285 2260 1286
rect 2254 1281 2255 1285
rect 2259 1281 2260 1285
rect 2254 1280 2260 1281
rect 2326 1285 2332 1286
rect 2326 1281 2327 1285
rect 2331 1281 2332 1285
rect 2326 1280 2332 1281
rect 2398 1285 2404 1286
rect 2398 1281 2399 1285
rect 2403 1281 2404 1285
rect 2398 1280 2404 1281
rect 2454 1285 2460 1286
rect 2454 1281 2455 1285
rect 2459 1281 2460 1285
rect 2454 1280 2460 1281
rect 2502 1284 2508 1285
rect 2502 1280 2503 1284
rect 2507 1280 2508 1284
rect 1326 1279 1332 1280
rect 2502 1279 2508 1280
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1263 1332 1267
rect 2502 1267 2508 1268
rect 1326 1262 1332 1263
rect 1350 1264 1356 1265
rect 1350 1260 1351 1264
rect 1355 1260 1356 1264
rect 1350 1259 1356 1260
rect 1406 1264 1412 1265
rect 1406 1260 1407 1264
rect 1411 1260 1412 1264
rect 1406 1259 1412 1260
rect 1502 1264 1508 1265
rect 1502 1260 1503 1264
rect 1507 1260 1508 1264
rect 1502 1259 1508 1260
rect 1598 1264 1604 1265
rect 1598 1260 1599 1264
rect 1603 1260 1604 1264
rect 1598 1259 1604 1260
rect 1702 1264 1708 1265
rect 1702 1260 1703 1264
rect 1707 1260 1708 1264
rect 1702 1259 1708 1260
rect 1806 1264 1812 1265
rect 1806 1260 1807 1264
rect 1811 1260 1812 1264
rect 1806 1259 1812 1260
rect 1902 1264 1908 1265
rect 1902 1260 1903 1264
rect 1907 1260 1908 1264
rect 1902 1259 1908 1260
rect 1998 1264 2004 1265
rect 1998 1260 1999 1264
rect 2003 1260 2004 1264
rect 1998 1259 2004 1260
rect 2086 1264 2092 1265
rect 2086 1260 2087 1264
rect 2091 1260 2092 1264
rect 2086 1259 2092 1260
rect 2166 1264 2172 1265
rect 2166 1260 2167 1264
rect 2171 1260 2172 1264
rect 2166 1259 2172 1260
rect 2238 1264 2244 1265
rect 2238 1260 2239 1264
rect 2243 1260 2244 1264
rect 2238 1259 2244 1260
rect 2310 1264 2316 1265
rect 2310 1260 2311 1264
rect 2315 1260 2316 1264
rect 2310 1259 2316 1260
rect 2382 1264 2388 1265
rect 2382 1260 2383 1264
rect 2387 1260 2388 1264
rect 2382 1259 2388 1260
rect 2438 1264 2444 1265
rect 2438 1260 2439 1264
rect 2443 1260 2444 1264
rect 2502 1263 2503 1267
rect 2507 1263 2508 1267
rect 2502 1262 2508 1263
rect 2438 1259 2444 1260
rect 190 1253 196 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 190 1249 191 1253
rect 195 1249 196 1253
rect 190 1248 196 1249
rect 246 1253 252 1254
rect 246 1249 247 1253
rect 251 1249 252 1253
rect 246 1248 252 1249
rect 302 1253 308 1254
rect 302 1249 303 1253
rect 307 1249 308 1253
rect 302 1248 308 1249
rect 366 1253 372 1254
rect 366 1249 367 1253
rect 371 1249 372 1253
rect 366 1248 372 1249
rect 438 1253 444 1254
rect 438 1249 439 1253
rect 443 1249 444 1253
rect 438 1248 444 1249
rect 526 1253 532 1254
rect 526 1249 527 1253
rect 531 1249 532 1253
rect 526 1248 532 1249
rect 638 1253 644 1254
rect 638 1249 639 1253
rect 643 1249 644 1253
rect 638 1248 644 1249
rect 774 1253 780 1254
rect 774 1249 775 1253
rect 779 1249 780 1253
rect 774 1248 780 1249
rect 926 1253 932 1254
rect 926 1249 927 1253
rect 931 1249 932 1253
rect 926 1248 932 1249
rect 1094 1253 1100 1254
rect 1094 1249 1095 1253
rect 1099 1249 1100 1253
rect 1094 1248 1100 1249
rect 1238 1253 1244 1254
rect 1238 1249 1239 1253
rect 1243 1249 1244 1253
rect 1238 1248 1244 1249
rect 1286 1252 1292 1253
rect 1286 1248 1287 1252
rect 1291 1248 1292 1252
rect 110 1247 116 1248
rect 1286 1247 1292 1248
rect 1350 1236 1356 1237
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1286 1235 1292 1236
rect 110 1230 116 1231
rect 174 1232 180 1233
rect 174 1228 175 1232
rect 179 1228 180 1232
rect 174 1227 180 1228
rect 230 1232 236 1233
rect 230 1228 231 1232
rect 235 1228 236 1232
rect 230 1227 236 1228
rect 286 1232 292 1233
rect 286 1228 287 1232
rect 291 1228 292 1232
rect 286 1227 292 1228
rect 350 1232 356 1233
rect 350 1228 351 1232
rect 355 1228 356 1232
rect 350 1227 356 1228
rect 422 1232 428 1233
rect 422 1228 423 1232
rect 427 1228 428 1232
rect 422 1227 428 1228
rect 510 1232 516 1233
rect 510 1228 511 1232
rect 515 1228 516 1232
rect 510 1227 516 1228
rect 622 1232 628 1233
rect 622 1228 623 1232
rect 627 1228 628 1232
rect 622 1227 628 1228
rect 758 1232 764 1233
rect 758 1228 759 1232
rect 763 1228 764 1232
rect 758 1227 764 1228
rect 910 1232 916 1233
rect 910 1228 911 1232
rect 915 1228 916 1232
rect 910 1227 916 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1222 1232 1228 1233
rect 1222 1228 1223 1232
rect 1227 1228 1228 1232
rect 1286 1231 1287 1235
rect 1291 1231 1292 1235
rect 1286 1230 1292 1231
rect 1326 1233 1332 1234
rect 1326 1229 1327 1233
rect 1331 1229 1332 1233
rect 1350 1232 1351 1236
rect 1355 1232 1356 1236
rect 1350 1231 1356 1232
rect 1446 1236 1452 1237
rect 1446 1232 1447 1236
rect 1451 1232 1452 1236
rect 1446 1231 1452 1232
rect 1574 1236 1580 1237
rect 1574 1232 1575 1236
rect 1579 1232 1580 1236
rect 1574 1231 1580 1232
rect 1694 1236 1700 1237
rect 1694 1232 1695 1236
rect 1699 1232 1700 1236
rect 1694 1231 1700 1232
rect 1814 1236 1820 1237
rect 1814 1232 1815 1236
rect 1819 1232 1820 1236
rect 1814 1231 1820 1232
rect 1926 1236 1932 1237
rect 1926 1232 1927 1236
rect 1931 1232 1932 1236
rect 1926 1231 1932 1232
rect 2030 1236 2036 1237
rect 2030 1232 2031 1236
rect 2035 1232 2036 1236
rect 2030 1231 2036 1232
rect 2126 1236 2132 1237
rect 2126 1232 2127 1236
rect 2131 1232 2132 1236
rect 2126 1231 2132 1232
rect 2214 1236 2220 1237
rect 2214 1232 2215 1236
rect 2219 1232 2220 1236
rect 2214 1231 2220 1232
rect 2294 1236 2300 1237
rect 2294 1232 2295 1236
rect 2299 1232 2300 1236
rect 2294 1231 2300 1232
rect 2374 1236 2380 1237
rect 2374 1232 2375 1236
rect 2379 1232 2380 1236
rect 2374 1231 2380 1232
rect 2438 1236 2444 1237
rect 2438 1232 2439 1236
rect 2443 1232 2444 1236
rect 2438 1231 2444 1232
rect 2502 1233 2508 1234
rect 1326 1228 1332 1229
rect 2502 1229 2503 1233
rect 2507 1229 2508 1233
rect 2502 1228 2508 1229
rect 1222 1227 1228 1228
rect 350 1220 356 1221
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 350 1216 351 1220
rect 355 1216 356 1220
rect 350 1215 356 1216
rect 406 1220 412 1221
rect 406 1216 407 1220
rect 411 1216 412 1220
rect 406 1215 412 1216
rect 462 1220 468 1221
rect 462 1216 463 1220
rect 467 1216 468 1220
rect 462 1215 468 1216
rect 518 1220 524 1221
rect 518 1216 519 1220
rect 523 1216 524 1220
rect 518 1215 524 1216
rect 574 1220 580 1221
rect 574 1216 575 1220
rect 579 1216 580 1220
rect 574 1215 580 1216
rect 630 1220 636 1221
rect 630 1216 631 1220
rect 635 1216 636 1220
rect 630 1215 636 1216
rect 686 1220 692 1221
rect 686 1216 687 1220
rect 691 1216 692 1220
rect 686 1215 692 1216
rect 742 1220 748 1221
rect 742 1216 743 1220
rect 747 1216 748 1220
rect 742 1215 748 1216
rect 798 1220 804 1221
rect 798 1216 799 1220
rect 803 1216 804 1220
rect 798 1215 804 1216
rect 854 1220 860 1221
rect 854 1216 855 1220
rect 859 1216 860 1220
rect 854 1215 860 1216
rect 910 1220 916 1221
rect 910 1216 911 1220
rect 915 1216 916 1220
rect 910 1215 916 1216
rect 1286 1217 1292 1218
rect 110 1212 116 1213
rect 1286 1213 1287 1217
rect 1291 1213 1292 1217
rect 1286 1212 1292 1213
rect 1326 1216 1332 1217
rect 2502 1216 2508 1217
rect 1326 1212 1327 1216
rect 1331 1212 1332 1216
rect 1326 1211 1332 1212
rect 1366 1215 1372 1216
rect 1366 1211 1367 1215
rect 1371 1211 1372 1215
rect 1366 1210 1372 1211
rect 1462 1215 1468 1216
rect 1462 1211 1463 1215
rect 1467 1211 1468 1215
rect 1462 1210 1468 1211
rect 1590 1215 1596 1216
rect 1590 1211 1591 1215
rect 1595 1211 1596 1215
rect 1590 1210 1596 1211
rect 1710 1215 1716 1216
rect 1710 1211 1711 1215
rect 1715 1211 1716 1215
rect 1710 1210 1716 1211
rect 1830 1215 1836 1216
rect 1830 1211 1831 1215
rect 1835 1211 1836 1215
rect 1830 1210 1836 1211
rect 1942 1215 1948 1216
rect 1942 1211 1943 1215
rect 1947 1211 1948 1215
rect 1942 1210 1948 1211
rect 2046 1215 2052 1216
rect 2046 1211 2047 1215
rect 2051 1211 2052 1215
rect 2046 1210 2052 1211
rect 2142 1215 2148 1216
rect 2142 1211 2143 1215
rect 2147 1211 2148 1215
rect 2142 1210 2148 1211
rect 2230 1215 2236 1216
rect 2230 1211 2231 1215
rect 2235 1211 2236 1215
rect 2230 1210 2236 1211
rect 2310 1215 2316 1216
rect 2310 1211 2311 1215
rect 2315 1211 2316 1215
rect 2310 1210 2316 1211
rect 2390 1215 2396 1216
rect 2390 1211 2391 1215
rect 2395 1211 2396 1215
rect 2390 1210 2396 1211
rect 2454 1215 2460 1216
rect 2454 1211 2455 1215
rect 2459 1211 2460 1215
rect 2502 1212 2503 1216
rect 2507 1212 2508 1216
rect 2502 1211 2508 1212
rect 2454 1210 2460 1211
rect 110 1200 116 1201
rect 1286 1200 1292 1201
rect 110 1196 111 1200
rect 115 1196 116 1200
rect 110 1195 116 1196
rect 366 1199 372 1200
rect 366 1195 367 1199
rect 371 1195 372 1199
rect 366 1194 372 1195
rect 422 1199 428 1200
rect 422 1195 423 1199
rect 427 1195 428 1199
rect 422 1194 428 1195
rect 478 1199 484 1200
rect 478 1195 479 1199
rect 483 1195 484 1199
rect 478 1194 484 1195
rect 534 1199 540 1200
rect 534 1195 535 1199
rect 539 1195 540 1199
rect 534 1194 540 1195
rect 590 1199 596 1200
rect 590 1195 591 1199
rect 595 1195 596 1199
rect 590 1194 596 1195
rect 646 1199 652 1200
rect 646 1195 647 1199
rect 651 1195 652 1199
rect 646 1194 652 1195
rect 702 1199 708 1200
rect 702 1195 703 1199
rect 707 1195 708 1199
rect 702 1194 708 1195
rect 758 1199 764 1200
rect 758 1195 759 1199
rect 763 1195 764 1199
rect 758 1194 764 1195
rect 814 1199 820 1200
rect 814 1195 815 1199
rect 819 1195 820 1199
rect 814 1194 820 1195
rect 870 1199 876 1200
rect 870 1195 871 1199
rect 875 1195 876 1199
rect 870 1194 876 1195
rect 926 1199 932 1200
rect 926 1195 927 1199
rect 931 1195 932 1199
rect 1286 1196 1287 1200
rect 1291 1196 1292 1200
rect 1286 1195 1292 1196
rect 926 1194 932 1195
rect 1366 1165 1372 1166
rect 1326 1164 1332 1165
rect 1326 1160 1327 1164
rect 1331 1160 1332 1164
rect 1366 1161 1367 1165
rect 1371 1161 1372 1165
rect 1366 1160 1372 1161
rect 1470 1165 1476 1166
rect 1470 1161 1471 1165
rect 1475 1161 1476 1165
rect 1470 1160 1476 1161
rect 1598 1165 1604 1166
rect 1598 1161 1599 1165
rect 1603 1161 1604 1165
rect 1598 1160 1604 1161
rect 1734 1165 1740 1166
rect 1734 1161 1735 1165
rect 1739 1161 1740 1165
rect 1734 1160 1740 1161
rect 1862 1165 1868 1166
rect 1862 1161 1863 1165
rect 1867 1161 1868 1165
rect 1862 1160 1868 1161
rect 1982 1165 1988 1166
rect 1982 1161 1983 1165
rect 1987 1161 1988 1165
rect 1982 1160 1988 1161
rect 2086 1165 2092 1166
rect 2086 1161 2087 1165
rect 2091 1161 2092 1165
rect 2086 1160 2092 1161
rect 2190 1165 2196 1166
rect 2190 1161 2191 1165
rect 2195 1161 2196 1165
rect 2190 1160 2196 1161
rect 2286 1165 2292 1166
rect 2286 1161 2287 1165
rect 2291 1161 2292 1165
rect 2286 1160 2292 1161
rect 2382 1165 2388 1166
rect 2382 1161 2383 1165
rect 2387 1161 2388 1165
rect 2382 1160 2388 1161
rect 2454 1165 2460 1166
rect 2454 1161 2455 1165
rect 2459 1161 2460 1165
rect 2454 1160 2460 1161
rect 2502 1164 2508 1165
rect 2502 1160 2503 1164
rect 2507 1160 2508 1164
rect 1326 1159 1332 1160
rect 2502 1159 2508 1160
rect 1326 1147 1332 1148
rect 422 1145 428 1146
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 422 1141 423 1145
rect 427 1141 428 1145
rect 422 1140 428 1141
rect 478 1145 484 1146
rect 478 1141 479 1145
rect 483 1141 484 1145
rect 478 1140 484 1141
rect 534 1145 540 1146
rect 534 1141 535 1145
rect 539 1141 540 1145
rect 534 1140 540 1141
rect 590 1145 596 1146
rect 590 1141 591 1145
rect 595 1141 596 1145
rect 590 1140 596 1141
rect 646 1145 652 1146
rect 646 1141 647 1145
rect 651 1141 652 1145
rect 646 1140 652 1141
rect 702 1145 708 1146
rect 702 1141 703 1145
rect 707 1141 708 1145
rect 702 1140 708 1141
rect 758 1145 764 1146
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 814 1145 820 1146
rect 814 1141 815 1145
rect 819 1141 820 1145
rect 814 1140 820 1141
rect 870 1145 876 1146
rect 870 1141 871 1145
rect 875 1141 876 1145
rect 870 1140 876 1141
rect 926 1145 932 1146
rect 926 1141 927 1145
rect 931 1141 932 1145
rect 926 1140 932 1141
rect 982 1145 988 1146
rect 982 1141 983 1145
rect 987 1141 988 1145
rect 982 1140 988 1141
rect 1286 1144 1292 1145
rect 1286 1140 1287 1144
rect 1291 1140 1292 1144
rect 1326 1143 1327 1147
rect 1331 1143 1332 1147
rect 2502 1147 2508 1148
rect 1326 1142 1332 1143
rect 1350 1144 1356 1145
rect 110 1139 116 1140
rect 1286 1139 1292 1140
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1454 1144 1460 1145
rect 1454 1140 1455 1144
rect 1459 1140 1460 1144
rect 1454 1139 1460 1140
rect 1582 1144 1588 1145
rect 1582 1140 1583 1144
rect 1587 1140 1588 1144
rect 1582 1139 1588 1140
rect 1718 1144 1724 1145
rect 1718 1140 1719 1144
rect 1723 1140 1724 1144
rect 1718 1139 1724 1140
rect 1846 1144 1852 1145
rect 1846 1140 1847 1144
rect 1851 1140 1852 1144
rect 1846 1139 1852 1140
rect 1966 1144 1972 1145
rect 1966 1140 1967 1144
rect 1971 1140 1972 1144
rect 1966 1139 1972 1140
rect 2070 1144 2076 1145
rect 2070 1140 2071 1144
rect 2075 1140 2076 1144
rect 2070 1139 2076 1140
rect 2174 1144 2180 1145
rect 2174 1140 2175 1144
rect 2179 1140 2180 1144
rect 2174 1139 2180 1140
rect 2270 1144 2276 1145
rect 2270 1140 2271 1144
rect 2275 1140 2276 1144
rect 2270 1139 2276 1140
rect 2366 1144 2372 1145
rect 2366 1140 2367 1144
rect 2371 1140 2372 1144
rect 2366 1139 2372 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2502 1143 2503 1147
rect 2507 1143 2508 1147
rect 2502 1142 2508 1143
rect 2438 1139 2444 1140
rect 1366 1128 1372 1129
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 1286 1127 1292 1128
rect 110 1122 116 1123
rect 406 1124 412 1125
rect 406 1120 407 1124
rect 411 1120 412 1124
rect 406 1119 412 1120
rect 462 1124 468 1125
rect 462 1120 463 1124
rect 467 1120 468 1124
rect 462 1119 468 1120
rect 518 1124 524 1125
rect 518 1120 519 1124
rect 523 1120 524 1124
rect 518 1119 524 1120
rect 574 1124 580 1125
rect 574 1120 575 1124
rect 579 1120 580 1124
rect 574 1119 580 1120
rect 630 1124 636 1125
rect 630 1120 631 1124
rect 635 1120 636 1124
rect 630 1119 636 1120
rect 686 1124 692 1125
rect 686 1120 687 1124
rect 691 1120 692 1124
rect 686 1119 692 1120
rect 742 1124 748 1125
rect 742 1120 743 1124
rect 747 1120 748 1124
rect 742 1119 748 1120
rect 798 1124 804 1125
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 798 1119 804 1120
rect 854 1124 860 1125
rect 854 1120 855 1124
rect 859 1120 860 1124
rect 854 1119 860 1120
rect 910 1124 916 1125
rect 910 1120 911 1124
rect 915 1120 916 1124
rect 910 1119 916 1120
rect 966 1124 972 1125
rect 966 1120 967 1124
rect 971 1120 972 1124
rect 1286 1123 1287 1127
rect 1291 1123 1292 1127
rect 1286 1122 1292 1123
rect 1326 1125 1332 1126
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1366 1124 1367 1128
rect 1371 1124 1372 1128
rect 1366 1123 1372 1124
rect 1446 1128 1452 1129
rect 1446 1124 1447 1128
rect 1451 1124 1452 1128
rect 1446 1123 1452 1124
rect 1534 1128 1540 1129
rect 1534 1124 1535 1128
rect 1539 1124 1540 1128
rect 1534 1123 1540 1124
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1806 1128 1812 1129
rect 1806 1124 1807 1128
rect 1811 1124 1812 1128
rect 1806 1123 1812 1124
rect 1894 1128 1900 1129
rect 1894 1124 1895 1128
rect 1899 1124 1900 1128
rect 1894 1123 1900 1124
rect 1982 1128 1988 1129
rect 1982 1124 1983 1128
rect 1987 1124 1988 1128
rect 1982 1123 1988 1124
rect 2070 1128 2076 1129
rect 2070 1124 2071 1128
rect 2075 1124 2076 1128
rect 2070 1123 2076 1124
rect 2158 1128 2164 1129
rect 2158 1124 2159 1128
rect 2163 1124 2164 1128
rect 2158 1123 2164 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 2438 1128 2444 1129
rect 2438 1124 2439 1128
rect 2443 1124 2444 1128
rect 2438 1123 2444 1124
rect 2502 1125 2508 1126
rect 1326 1120 1332 1121
rect 2502 1121 2503 1125
rect 2507 1121 2508 1125
rect 2502 1120 2508 1121
rect 966 1119 972 1120
rect 222 1108 228 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 222 1104 223 1108
rect 227 1104 228 1108
rect 222 1103 228 1104
rect 310 1108 316 1109
rect 310 1104 311 1108
rect 315 1104 316 1108
rect 310 1103 316 1104
rect 398 1108 404 1109
rect 398 1104 399 1108
rect 403 1104 404 1108
rect 398 1103 404 1104
rect 494 1108 500 1109
rect 494 1104 495 1108
rect 499 1104 500 1108
rect 494 1103 500 1104
rect 590 1108 596 1109
rect 590 1104 591 1108
rect 595 1104 596 1108
rect 590 1103 596 1104
rect 678 1108 684 1109
rect 678 1104 679 1108
rect 683 1104 684 1108
rect 678 1103 684 1104
rect 766 1108 772 1109
rect 766 1104 767 1108
rect 771 1104 772 1108
rect 766 1103 772 1104
rect 846 1108 852 1109
rect 846 1104 847 1108
rect 851 1104 852 1108
rect 846 1103 852 1104
rect 926 1108 932 1109
rect 926 1104 927 1108
rect 931 1104 932 1108
rect 926 1103 932 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1102 1108 1108 1109
rect 1102 1104 1103 1108
rect 1107 1104 1108 1108
rect 1326 1108 1332 1109
rect 2502 1108 2508 1109
rect 1102 1103 1108 1104
rect 1286 1105 1292 1106
rect 110 1100 116 1101
rect 1286 1101 1287 1105
rect 1291 1101 1292 1105
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1326 1103 1332 1104
rect 1382 1107 1388 1108
rect 1382 1103 1383 1107
rect 1387 1103 1388 1107
rect 1382 1102 1388 1103
rect 1462 1107 1468 1108
rect 1462 1103 1463 1107
rect 1467 1103 1468 1107
rect 1462 1102 1468 1103
rect 1550 1107 1556 1108
rect 1550 1103 1551 1107
rect 1555 1103 1556 1107
rect 1550 1102 1556 1103
rect 1646 1107 1652 1108
rect 1646 1103 1647 1107
rect 1651 1103 1652 1107
rect 1646 1102 1652 1103
rect 1734 1107 1740 1108
rect 1734 1103 1735 1107
rect 1739 1103 1740 1107
rect 1734 1102 1740 1103
rect 1822 1107 1828 1108
rect 1822 1103 1823 1107
rect 1827 1103 1828 1107
rect 1822 1102 1828 1103
rect 1910 1107 1916 1108
rect 1910 1103 1911 1107
rect 1915 1103 1916 1107
rect 1910 1102 1916 1103
rect 1998 1107 2004 1108
rect 1998 1103 1999 1107
rect 2003 1103 2004 1107
rect 1998 1102 2004 1103
rect 2086 1107 2092 1108
rect 2086 1103 2087 1107
rect 2091 1103 2092 1107
rect 2086 1102 2092 1103
rect 2174 1107 2180 1108
rect 2174 1103 2175 1107
rect 2179 1103 2180 1107
rect 2174 1102 2180 1103
rect 2270 1107 2276 1108
rect 2270 1103 2271 1107
rect 2275 1103 2276 1107
rect 2270 1102 2276 1103
rect 2374 1107 2380 1108
rect 2374 1103 2375 1107
rect 2379 1103 2380 1107
rect 2374 1102 2380 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2502 1104 2503 1108
rect 2507 1104 2508 1108
rect 2502 1103 2508 1104
rect 2454 1102 2460 1103
rect 1286 1100 1292 1101
rect 110 1088 116 1089
rect 1286 1088 1292 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 238 1087 244 1088
rect 238 1083 239 1087
rect 243 1083 244 1087
rect 238 1082 244 1083
rect 326 1087 332 1088
rect 326 1083 327 1087
rect 331 1083 332 1087
rect 326 1082 332 1083
rect 414 1087 420 1088
rect 414 1083 415 1087
rect 419 1083 420 1087
rect 414 1082 420 1083
rect 510 1087 516 1088
rect 510 1083 511 1087
rect 515 1083 516 1087
rect 510 1082 516 1083
rect 606 1087 612 1088
rect 606 1083 607 1087
rect 611 1083 612 1087
rect 606 1082 612 1083
rect 694 1087 700 1088
rect 694 1083 695 1087
rect 699 1083 700 1087
rect 694 1082 700 1083
rect 782 1087 788 1088
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 862 1087 868 1088
rect 862 1083 863 1087
rect 867 1083 868 1087
rect 862 1082 868 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 942 1082 948 1083
rect 1030 1087 1036 1088
rect 1030 1083 1031 1087
rect 1035 1083 1036 1087
rect 1030 1082 1036 1083
rect 1118 1087 1124 1088
rect 1118 1083 1119 1087
rect 1123 1083 1124 1087
rect 1286 1084 1287 1088
rect 1291 1084 1292 1088
rect 1286 1083 1292 1084
rect 1118 1082 1124 1083
rect 1430 1049 1436 1050
rect 1326 1048 1332 1049
rect 1326 1044 1327 1048
rect 1331 1044 1332 1048
rect 1430 1045 1431 1049
rect 1435 1045 1436 1049
rect 1430 1044 1436 1045
rect 1494 1049 1500 1050
rect 1494 1045 1495 1049
rect 1499 1045 1500 1049
rect 1494 1044 1500 1045
rect 1566 1049 1572 1050
rect 1566 1045 1567 1049
rect 1571 1045 1572 1049
rect 1566 1044 1572 1045
rect 1638 1049 1644 1050
rect 1638 1045 1639 1049
rect 1643 1045 1644 1049
rect 1638 1044 1644 1045
rect 1702 1049 1708 1050
rect 1702 1045 1703 1049
rect 1707 1045 1708 1049
rect 1702 1044 1708 1045
rect 1766 1049 1772 1050
rect 1766 1045 1767 1049
rect 1771 1045 1772 1049
rect 1766 1044 1772 1045
rect 1838 1049 1844 1050
rect 1838 1045 1839 1049
rect 1843 1045 1844 1049
rect 1838 1044 1844 1045
rect 1918 1049 1924 1050
rect 1918 1045 1919 1049
rect 1923 1045 1924 1049
rect 1918 1044 1924 1045
rect 2006 1049 2012 1050
rect 2006 1045 2007 1049
rect 2011 1045 2012 1049
rect 2006 1044 2012 1045
rect 2110 1049 2116 1050
rect 2110 1045 2111 1049
rect 2115 1045 2116 1049
rect 2110 1044 2116 1045
rect 2230 1049 2236 1050
rect 2230 1045 2231 1049
rect 2235 1045 2236 1049
rect 2230 1044 2236 1045
rect 2350 1049 2356 1050
rect 2350 1045 2351 1049
rect 2355 1045 2356 1049
rect 2350 1044 2356 1045
rect 2454 1049 2460 1050
rect 2454 1045 2455 1049
rect 2459 1045 2460 1049
rect 2454 1044 2460 1045
rect 2502 1048 2508 1049
rect 2502 1044 2503 1048
rect 2507 1044 2508 1048
rect 1326 1043 1332 1044
rect 2502 1043 2508 1044
rect 150 1033 156 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 150 1029 151 1033
rect 155 1029 156 1033
rect 150 1028 156 1029
rect 206 1033 212 1034
rect 206 1029 207 1033
rect 211 1029 212 1033
rect 206 1028 212 1029
rect 302 1033 308 1034
rect 302 1029 303 1033
rect 307 1029 308 1033
rect 302 1028 308 1029
rect 414 1033 420 1034
rect 414 1029 415 1033
rect 419 1029 420 1033
rect 414 1028 420 1029
rect 534 1033 540 1034
rect 534 1029 535 1033
rect 539 1029 540 1033
rect 534 1028 540 1029
rect 654 1033 660 1034
rect 654 1029 655 1033
rect 659 1029 660 1033
rect 654 1028 660 1029
rect 766 1033 772 1034
rect 766 1029 767 1033
rect 771 1029 772 1033
rect 766 1028 772 1029
rect 878 1033 884 1034
rect 878 1029 879 1033
rect 883 1029 884 1033
rect 878 1028 884 1029
rect 982 1033 988 1034
rect 982 1029 983 1033
rect 987 1029 988 1033
rect 982 1028 988 1029
rect 1094 1033 1100 1034
rect 1094 1029 1095 1033
rect 1099 1029 1100 1033
rect 1094 1028 1100 1029
rect 1206 1033 1212 1034
rect 1206 1029 1207 1033
rect 1211 1029 1212 1033
rect 1206 1028 1212 1029
rect 1286 1032 1292 1033
rect 1286 1028 1287 1032
rect 1291 1028 1292 1032
rect 110 1027 116 1028
rect 1286 1027 1292 1028
rect 1326 1031 1332 1032
rect 1326 1027 1327 1031
rect 1331 1027 1332 1031
rect 2502 1031 2508 1032
rect 1326 1026 1332 1027
rect 1414 1028 1420 1029
rect 1414 1024 1415 1028
rect 1419 1024 1420 1028
rect 1414 1023 1420 1024
rect 1478 1028 1484 1029
rect 1478 1024 1479 1028
rect 1483 1024 1484 1028
rect 1478 1023 1484 1024
rect 1550 1028 1556 1029
rect 1550 1024 1551 1028
rect 1555 1024 1556 1028
rect 1550 1023 1556 1024
rect 1622 1028 1628 1029
rect 1622 1024 1623 1028
rect 1627 1024 1628 1028
rect 1622 1023 1628 1024
rect 1686 1028 1692 1029
rect 1686 1024 1687 1028
rect 1691 1024 1692 1028
rect 1686 1023 1692 1024
rect 1750 1028 1756 1029
rect 1750 1024 1751 1028
rect 1755 1024 1756 1028
rect 1750 1023 1756 1024
rect 1822 1028 1828 1029
rect 1822 1024 1823 1028
rect 1827 1024 1828 1028
rect 1822 1023 1828 1024
rect 1902 1028 1908 1029
rect 1902 1024 1903 1028
rect 1907 1024 1908 1028
rect 1902 1023 1908 1024
rect 1990 1028 1996 1029
rect 1990 1024 1991 1028
rect 1995 1024 1996 1028
rect 1990 1023 1996 1024
rect 2094 1028 2100 1029
rect 2094 1024 2095 1028
rect 2099 1024 2100 1028
rect 2094 1023 2100 1024
rect 2214 1028 2220 1029
rect 2214 1024 2215 1028
rect 2219 1024 2220 1028
rect 2214 1023 2220 1024
rect 2334 1028 2340 1029
rect 2334 1024 2335 1028
rect 2339 1024 2340 1028
rect 2334 1023 2340 1024
rect 2438 1028 2444 1029
rect 2438 1024 2439 1028
rect 2443 1024 2444 1028
rect 2502 1027 2503 1031
rect 2507 1027 2508 1031
rect 2502 1026 2508 1027
rect 2438 1023 2444 1024
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 1286 1015 1292 1016
rect 110 1010 116 1011
rect 134 1012 140 1013
rect 134 1008 135 1012
rect 139 1008 140 1012
rect 134 1007 140 1008
rect 190 1012 196 1013
rect 190 1008 191 1012
rect 195 1008 196 1012
rect 190 1007 196 1008
rect 286 1012 292 1013
rect 286 1008 287 1012
rect 291 1008 292 1012
rect 286 1007 292 1008
rect 398 1012 404 1013
rect 398 1008 399 1012
rect 403 1008 404 1012
rect 398 1007 404 1008
rect 518 1012 524 1013
rect 518 1008 519 1012
rect 523 1008 524 1012
rect 518 1007 524 1008
rect 638 1012 644 1013
rect 638 1008 639 1012
rect 643 1008 644 1012
rect 638 1007 644 1008
rect 750 1012 756 1013
rect 750 1008 751 1012
rect 755 1008 756 1012
rect 750 1007 756 1008
rect 862 1012 868 1013
rect 862 1008 863 1012
rect 867 1008 868 1012
rect 862 1007 868 1008
rect 966 1012 972 1013
rect 966 1008 967 1012
rect 971 1008 972 1012
rect 966 1007 972 1008
rect 1078 1012 1084 1013
rect 1078 1008 1079 1012
rect 1083 1008 1084 1012
rect 1078 1007 1084 1008
rect 1190 1012 1196 1013
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1286 1011 1287 1015
rect 1291 1011 1292 1015
rect 1286 1010 1292 1011
rect 1190 1007 1196 1008
rect 1510 1008 1516 1009
rect 1326 1005 1332 1006
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1566 1008 1572 1009
rect 1566 1004 1567 1008
rect 1571 1004 1572 1008
rect 1566 1003 1572 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1734 1008 1740 1009
rect 1734 1004 1735 1008
rect 1739 1004 1740 1008
rect 1734 1003 1740 1004
rect 1806 1008 1812 1009
rect 1806 1004 1807 1008
rect 1811 1004 1812 1008
rect 1806 1003 1812 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1982 1008 1988 1009
rect 1982 1004 1983 1008
rect 1987 1004 1988 1008
rect 1982 1003 1988 1004
rect 2094 1008 2100 1009
rect 2094 1004 2095 1008
rect 2099 1004 2100 1008
rect 2094 1003 2100 1004
rect 2214 1008 2220 1009
rect 2214 1004 2215 1008
rect 2219 1004 2220 1008
rect 2214 1003 2220 1004
rect 2334 1008 2340 1009
rect 2334 1004 2335 1008
rect 2339 1004 2340 1008
rect 2334 1003 2340 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 134 996 140 997
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 134 992 135 996
rect 139 992 140 996
rect 134 991 140 992
rect 214 996 220 997
rect 214 992 215 996
rect 219 992 220 996
rect 214 991 220 992
rect 326 996 332 997
rect 326 992 327 996
rect 331 992 332 996
rect 326 991 332 992
rect 438 996 444 997
rect 438 992 439 996
rect 443 992 444 996
rect 438 991 444 992
rect 550 996 556 997
rect 550 992 551 996
rect 555 992 556 996
rect 550 991 556 992
rect 662 996 668 997
rect 662 992 663 996
rect 667 992 668 996
rect 662 991 668 992
rect 758 996 764 997
rect 758 992 759 996
rect 763 992 764 996
rect 758 991 764 992
rect 846 996 852 997
rect 846 992 847 996
rect 851 992 852 996
rect 846 991 852 992
rect 934 996 940 997
rect 934 992 935 996
rect 939 992 940 996
rect 934 991 940 992
rect 1014 996 1020 997
rect 1014 992 1015 996
rect 1019 992 1020 996
rect 1014 991 1020 992
rect 1086 996 1092 997
rect 1086 992 1087 996
rect 1091 992 1092 996
rect 1086 991 1092 992
rect 1166 996 1172 997
rect 1166 992 1167 996
rect 1171 992 1172 996
rect 1166 991 1172 992
rect 1222 996 1228 997
rect 1222 992 1223 996
rect 1227 992 1228 996
rect 1222 991 1228 992
rect 1286 993 1292 994
rect 110 988 116 989
rect 1286 989 1287 993
rect 1291 989 1292 993
rect 1286 988 1292 989
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1582 987 1588 988
rect 1582 983 1583 987
rect 1587 983 1588 987
rect 1582 982 1588 983
rect 1638 987 1644 988
rect 1638 983 1639 987
rect 1643 983 1644 987
rect 1638 982 1644 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1750 987 1756 988
rect 1750 983 1751 987
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1822 987 1828 988
rect 1822 983 1823 987
rect 1827 983 1828 987
rect 1822 982 1828 983
rect 1902 987 1908 988
rect 1902 983 1903 987
rect 1907 983 1908 987
rect 1902 982 1908 983
rect 1998 987 2004 988
rect 1998 983 1999 987
rect 2003 983 2004 987
rect 1998 982 2004 983
rect 2110 987 2116 988
rect 2110 983 2111 987
rect 2115 983 2116 987
rect 2110 982 2116 983
rect 2230 987 2236 988
rect 2230 983 2231 987
rect 2235 983 2236 987
rect 2230 982 2236 983
rect 2350 987 2356 988
rect 2350 983 2351 987
rect 2355 983 2356 987
rect 2350 982 2356 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2454 982 2460 983
rect 110 976 116 977
rect 1286 976 1292 977
rect 110 972 111 976
rect 115 972 116 976
rect 110 971 116 972
rect 150 975 156 976
rect 150 971 151 975
rect 155 971 156 975
rect 150 970 156 971
rect 230 975 236 976
rect 230 971 231 975
rect 235 971 236 975
rect 230 970 236 971
rect 342 975 348 976
rect 342 971 343 975
rect 347 971 348 975
rect 342 970 348 971
rect 454 975 460 976
rect 454 971 455 975
rect 459 971 460 975
rect 454 970 460 971
rect 566 975 572 976
rect 566 971 567 975
rect 571 971 572 975
rect 566 970 572 971
rect 678 975 684 976
rect 678 971 679 975
rect 683 971 684 975
rect 678 970 684 971
rect 774 975 780 976
rect 774 971 775 975
rect 779 971 780 975
rect 774 970 780 971
rect 862 975 868 976
rect 862 971 863 975
rect 867 971 868 975
rect 862 970 868 971
rect 950 975 956 976
rect 950 971 951 975
rect 955 971 956 975
rect 950 970 956 971
rect 1030 975 1036 976
rect 1030 971 1031 975
rect 1035 971 1036 975
rect 1030 970 1036 971
rect 1102 975 1108 976
rect 1102 971 1103 975
rect 1107 971 1108 975
rect 1102 970 1108 971
rect 1182 975 1188 976
rect 1182 971 1183 975
rect 1187 971 1188 975
rect 1182 970 1188 971
rect 1238 975 1244 976
rect 1238 971 1239 975
rect 1243 971 1244 975
rect 1286 972 1287 976
rect 1291 972 1292 976
rect 1286 971 1292 972
rect 1238 970 1244 971
rect 150 925 156 926
rect 110 924 116 925
rect 110 920 111 924
rect 115 920 116 924
rect 150 921 151 925
rect 155 921 156 925
rect 150 920 156 921
rect 206 925 212 926
rect 206 921 207 925
rect 211 921 212 925
rect 206 920 212 921
rect 294 925 300 926
rect 294 921 295 925
rect 299 921 300 925
rect 294 920 300 921
rect 398 925 404 926
rect 398 921 399 925
rect 403 921 404 925
rect 398 920 404 921
rect 510 925 516 926
rect 510 921 511 925
rect 515 921 516 925
rect 510 920 516 921
rect 622 925 628 926
rect 622 921 623 925
rect 627 921 628 925
rect 622 920 628 921
rect 734 925 740 926
rect 734 921 735 925
rect 739 921 740 925
rect 734 920 740 921
rect 830 925 836 926
rect 830 921 831 925
rect 835 921 836 925
rect 830 920 836 921
rect 926 925 932 926
rect 926 921 927 925
rect 931 921 932 925
rect 926 920 932 921
rect 1014 925 1020 926
rect 1014 921 1015 925
rect 1019 921 1020 925
rect 1014 920 1020 921
rect 1094 925 1100 926
rect 1094 921 1095 925
rect 1099 921 1100 925
rect 1094 920 1100 921
rect 1174 925 1180 926
rect 1174 921 1175 925
rect 1179 921 1180 925
rect 1174 920 1180 921
rect 1238 925 1244 926
rect 1238 921 1239 925
rect 1243 921 1244 925
rect 1238 920 1244 921
rect 1286 924 1292 925
rect 1286 920 1287 924
rect 1291 920 1292 924
rect 1366 921 1372 922
rect 110 919 116 920
rect 1286 919 1292 920
rect 1326 920 1332 921
rect 1326 916 1327 920
rect 1331 916 1332 920
rect 1366 917 1367 921
rect 1371 917 1372 921
rect 1366 916 1372 917
rect 1438 921 1444 922
rect 1438 917 1439 921
rect 1443 917 1444 921
rect 1438 916 1444 917
rect 1526 921 1532 922
rect 1526 917 1527 921
rect 1531 917 1532 921
rect 1526 916 1532 917
rect 1614 921 1620 922
rect 1614 917 1615 921
rect 1619 917 1620 921
rect 1614 916 1620 917
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1790 921 1796 922
rect 1790 917 1791 921
rect 1795 917 1796 921
rect 1790 916 1796 917
rect 1894 921 1900 922
rect 1894 917 1895 921
rect 1899 917 1900 921
rect 1894 916 1900 917
rect 2014 921 2020 922
rect 2014 917 2015 921
rect 2019 917 2020 921
rect 2014 916 2020 917
rect 2150 921 2156 922
rect 2150 917 2151 921
rect 2155 917 2156 921
rect 2150 916 2156 917
rect 2294 921 2300 922
rect 2294 917 2295 921
rect 2299 917 2300 921
rect 2294 916 2300 917
rect 2438 921 2444 922
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2438 916 2444 917
rect 2502 920 2508 921
rect 2502 916 2503 920
rect 2507 916 2508 920
rect 1326 915 1332 916
rect 2502 915 2508 916
rect 110 907 116 908
rect 110 903 111 907
rect 115 903 116 907
rect 1286 907 1292 908
rect 110 902 116 903
rect 134 904 140 905
rect 134 900 135 904
rect 139 900 140 904
rect 134 899 140 900
rect 190 904 196 905
rect 190 900 191 904
rect 195 900 196 904
rect 190 899 196 900
rect 278 904 284 905
rect 278 900 279 904
rect 283 900 284 904
rect 278 899 284 900
rect 382 904 388 905
rect 382 900 383 904
rect 387 900 388 904
rect 382 899 388 900
rect 494 904 500 905
rect 494 900 495 904
rect 499 900 500 904
rect 494 899 500 900
rect 606 904 612 905
rect 606 900 607 904
rect 611 900 612 904
rect 606 899 612 900
rect 718 904 724 905
rect 718 900 719 904
rect 723 900 724 904
rect 718 899 724 900
rect 814 904 820 905
rect 814 900 815 904
rect 819 900 820 904
rect 814 899 820 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 998 904 1004 905
rect 998 900 999 904
rect 1003 900 1004 904
rect 998 899 1004 900
rect 1078 904 1084 905
rect 1078 900 1079 904
rect 1083 900 1084 904
rect 1078 899 1084 900
rect 1158 904 1164 905
rect 1158 900 1159 904
rect 1163 900 1164 904
rect 1158 899 1164 900
rect 1222 904 1228 905
rect 1222 900 1223 904
rect 1227 900 1228 904
rect 1286 903 1287 907
rect 1291 903 1292 907
rect 1286 902 1292 903
rect 1326 903 1332 904
rect 1222 899 1228 900
rect 1326 899 1327 903
rect 1331 899 1332 903
rect 2502 903 2508 904
rect 1326 898 1332 899
rect 1350 900 1356 901
rect 1350 896 1351 900
rect 1355 896 1356 900
rect 1350 895 1356 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1510 900 1516 901
rect 1510 896 1511 900
rect 1515 896 1516 900
rect 1510 895 1516 896
rect 1598 900 1604 901
rect 1598 896 1599 900
rect 1603 896 1604 900
rect 1598 895 1604 896
rect 1678 900 1684 901
rect 1678 896 1679 900
rect 1683 896 1684 900
rect 1678 895 1684 896
rect 1774 900 1780 901
rect 1774 896 1775 900
rect 1779 896 1780 900
rect 1774 895 1780 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1998 900 2004 901
rect 1998 896 1999 900
rect 2003 896 2004 900
rect 1998 895 2004 896
rect 2134 900 2140 901
rect 2134 896 2135 900
rect 2139 896 2140 900
rect 2134 895 2140 896
rect 2278 900 2284 901
rect 2278 896 2279 900
rect 2283 896 2284 900
rect 2278 895 2284 896
rect 2422 900 2428 901
rect 2422 896 2423 900
rect 2427 896 2428 900
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2422 895 2428 896
rect 246 888 252 889
rect 110 885 116 886
rect 110 881 111 885
rect 115 881 116 885
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 342 888 348 889
rect 342 884 343 888
rect 347 884 348 888
rect 342 883 348 884
rect 438 888 444 889
rect 438 884 439 888
rect 443 884 444 888
rect 438 883 444 884
rect 542 888 548 889
rect 542 884 543 888
rect 547 884 548 888
rect 542 883 548 884
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 742 888 748 889
rect 742 884 743 888
rect 747 884 748 888
rect 742 883 748 884
rect 838 888 844 889
rect 838 884 839 888
rect 843 884 844 888
rect 838 883 844 884
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 1006 888 1012 889
rect 1006 884 1007 888
rect 1011 884 1012 888
rect 1006 883 1012 884
rect 1086 888 1092 889
rect 1086 884 1087 888
rect 1091 884 1092 888
rect 1086 883 1092 884
rect 1166 888 1172 889
rect 1166 884 1167 888
rect 1171 884 1172 888
rect 1166 883 1172 884
rect 1222 888 1228 889
rect 1222 884 1223 888
rect 1227 884 1228 888
rect 1222 883 1228 884
rect 1286 885 1292 886
rect 110 880 116 881
rect 1286 881 1287 885
rect 1291 881 1292 885
rect 1286 880 1292 881
rect 1486 880 1492 881
rect 1326 877 1332 878
rect 1326 873 1327 877
rect 1331 873 1332 877
rect 1486 876 1487 880
rect 1491 876 1492 880
rect 1486 875 1492 876
rect 1558 880 1564 881
rect 1558 876 1559 880
rect 1563 876 1564 880
rect 1558 875 1564 876
rect 1622 880 1628 881
rect 1622 876 1623 880
rect 1627 876 1628 880
rect 1622 875 1628 876
rect 1686 880 1692 881
rect 1686 876 1687 880
rect 1691 876 1692 880
rect 1686 875 1692 876
rect 1750 880 1756 881
rect 1750 876 1751 880
rect 1755 876 1756 880
rect 1750 875 1756 876
rect 1814 880 1820 881
rect 1814 876 1815 880
rect 1819 876 1820 880
rect 1814 875 1820 876
rect 1886 880 1892 881
rect 1886 876 1887 880
rect 1891 876 1892 880
rect 1886 875 1892 876
rect 1974 880 1980 881
rect 1974 876 1975 880
rect 1979 876 1980 880
rect 1974 875 1980 876
rect 2078 880 2084 881
rect 2078 876 2079 880
rect 2083 876 2084 880
rect 2078 875 2084 876
rect 2198 880 2204 881
rect 2198 876 2199 880
rect 2203 876 2204 880
rect 2198 875 2204 876
rect 2318 880 2324 881
rect 2318 876 2319 880
rect 2323 876 2324 880
rect 2318 875 2324 876
rect 2438 880 2444 881
rect 2438 876 2439 880
rect 2443 876 2444 880
rect 2438 875 2444 876
rect 2502 877 2508 878
rect 1326 872 1332 873
rect 2502 873 2503 877
rect 2507 873 2508 877
rect 2502 872 2508 873
rect 110 868 116 869
rect 1286 868 1292 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 262 867 268 868
rect 262 863 263 867
rect 267 863 268 867
rect 262 862 268 863
rect 358 867 364 868
rect 358 863 359 867
rect 363 863 364 867
rect 358 862 364 863
rect 454 867 460 868
rect 454 863 455 867
rect 459 863 460 867
rect 454 862 460 863
rect 558 867 564 868
rect 558 863 559 867
rect 563 863 564 867
rect 558 862 564 863
rect 662 867 668 868
rect 662 863 663 867
rect 667 863 668 867
rect 662 862 668 863
rect 758 867 764 868
rect 758 863 759 867
rect 763 863 764 867
rect 758 862 764 863
rect 854 867 860 868
rect 854 863 855 867
rect 859 863 860 867
rect 854 862 860 863
rect 942 867 948 868
rect 942 863 943 867
rect 947 863 948 867
rect 942 862 948 863
rect 1022 867 1028 868
rect 1022 863 1023 867
rect 1027 863 1028 867
rect 1022 862 1028 863
rect 1102 867 1108 868
rect 1102 863 1103 867
rect 1107 863 1108 867
rect 1102 862 1108 863
rect 1182 867 1188 868
rect 1182 863 1183 867
rect 1187 863 1188 867
rect 1182 862 1188 863
rect 1238 867 1244 868
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 1286 864 1287 868
rect 1291 864 1292 868
rect 1286 863 1292 864
rect 1238 862 1244 863
rect 1326 860 1332 861
rect 2502 860 2508 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1502 859 1508 860
rect 1502 855 1503 859
rect 1507 855 1508 859
rect 1502 854 1508 855
rect 1574 859 1580 860
rect 1574 855 1575 859
rect 1579 855 1580 859
rect 1574 854 1580 855
rect 1638 859 1644 860
rect 1638 855 1639 859
rect 1643 855 1644 859
rect 1638 854 1644 855
rect 1702 859 1708 860
rect 1702 855 1703 859
rect 1707 855 1708 859
rect 1702 854 1708 855
rect 1766 859 1772 860
rect 1766 855 1767 859
rect 1771 855 1772 859
rect 1766 854 1772 855
rect 1830 859 1836 860
rect 1830 855 1831 859
rect 1835 855 1836 859
rect 1830 854 1836 855
rect 1902 859 1908 860
rect 1902 855 1903 859
rect 1907 855 1908 859
rect 1902 854 1908 855
rect 1990 859 1996 860
rect 1990 855 1991 859
rect 1995 855 1996 859
rect 1990 854 1996 855
rect 2094 859 2100 860
rect 2094 855 2095 859
rect 2099 855 2100 859
rect 2094 854 2100 855
rect 2214 859 2220 860
rect 2214 855 2215 859
rect 2219 855 2220 859
rect 2214 854 2220 855
rect 2334 859 2340 860
rect 2334 855 2335 859
rect 2339 855 2340 859
rect 2334 854 2340 855
rect 2454 859 2460 860
rect 2454 855 2455 859
rect 2459 855 2460 859
rect 2502 856 2503 860
rect 2507 856 2508 860
rect 2502 855 2508 856
rect 2454 854 2460 855
rect 238 813 244 814
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 238 809 239 813
rect 243 809 244 813
rect 238 808 244 809
rect 302 813 308 814
rect 302 809 303 813
rect 307 809 308 813
rect 302 808 308 809
rect 382 813 388 814
rect 382 809 383 813
rect 387 809 388 813
rect 382 808 388 809
rect 462 813 468 814
rect 462 809 463 813
rect 467 809 468 813
rect 462 808 468 809
rect 550 813 556 814
rect 550 809 551 813
rect 555 809 556 813
rect 550 808 556 809
rect 638 813 644 814
rect 638 809 639 813
rect 643 809 644 813
rect 638 808 644 809
rect 726 813 732 814
rect 726 809 727 813
rect 731 809 732 813
rect 726 808 732 809
rect 806 813 812 814
rect 806 809 807 813
rect 811 809 812 813
rect 806 808 812 809
rect 894 813 900 814
rect 894 809 895 813
rect 899 809 900 813
rect 894 808 900 809
rect 982 813 988 814
rect 982 809 983 813
rect 987 809 988 813
rect 982 808 988 809
rect 1070 813 1076 814
rect 1070 809 1071 813
rect 1075 809 1076 813
rect 1070 808 1076 809
rect 1286 812 1292 813
rect 1286 808 1287 812
rect 1291 808 1292 812
rect 110 807 116 808
rect 1286 807 1292 808
rect 1438 801 1444 802
rect 1326 800 1332 801
rect 1326 796 1327 800
rect 1331 796 1332 800
rect 1438 797 1439 801
rect 1443 797 1444 801
rect 1438 796 1444 797
rect 1510 801 1516 802
rect 1510 797 1511 801
rect 1515 797 1516 801
rect 1510 796 1516 797
rect 1590 801 1596 802
rect 1590 797 1591 801
rect 1595 797 1596 801
rect 1590 796 1596 797
rect 1670 801 1676 802
rect 1670 797 1671 801
rect 1675 797 1676 801
rect 1670 796 1676 797
rect 1758 801 1764 802
rect 1758 797 1759 801
rect 1763 797 1764 801
rect 1758 796 1764 797
rect 1846 801 1852 802
rect 1846 797 1847 801
rect 1851 797 1852 801
rect 1846 796 1852 797
rect 1934 801 1940 802
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 2022 801 2028 802
rect 2022 797 2023 801
rect 2027 797 2028 801
rect 2022 796 2028 797
rect 2110 801 2116 802
rect 2110 797 2111 801
rect 2115 797 2116 801
rect 2110 796 2116 797
rect 2198 801 2204 802
rect 2198 797 2199 801
rect 2203 797 2204 801
rect 2198 796 2204 797
rect 2286 801 2292 802
rect 2286 797 2287 801
rect 2291 797 2292 801
rect 2286 796 2292 797
rect 2382 801 2388 802
rect 2382 797 2383 801
rect 2387 797 2388 801
rect 2382 796 2388 797
rect 2454 801 2460 802
rect 2454 797 2455 801
rect 2459 797 2460 801
rect 2454 796 2460 797
rect 2502 800 2508 801
rect 2502 796 2503 800
rect 2507 796 2508 800
rect 110 795 116 796
rect 110 791 111 795
rect 115 791 116 795
rect 1286 795 1292 796
rect 1326 795 1332 796
rect 2502 795 2508 796
rect 110 790 116 791
rect 222 792 228 793
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 286 792 292 793
rect 286 788 287 792
rect 291 788 292 792
rect 286 787 292 788
rect 366 792 372 793
rect 366 788 367 792
rect 371 788 372 792
rect 366 787 372 788
rect 446 792 452 793
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 534 792 540 793
rect 534 788 535 792
rect 539 788 540 792
rect 534 787 540 788
rect 622 792 628 793
rect 622 788 623 792
rect 627 788 628 792
rect 622 787 628 788
rect 710 792 716 793
rect 710 788 711 792
rect 715 788 716 792
rect 710 787 716 788
rect 790 792 796 793
rect 790 788 791 792
rect 795 788 796 792
rect 790 787 796 788
rect 878 792 884 793
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 966 792 972 793
rect 966 788 967 792
rect 971 788 972 792
rect 966 787 972 788
rect 1054 792 1060 793
rect 1054 788 1055 792
rect 1059 788 1060 792
rect 1286 791 1287 795
rect 1291 791 1292 795
rect 1286 790 1292 791
rect 1054 787 1060 788
rect 1326 783 1332 784
rect 1326 779 1327 783
rect 1331 779 1332 783
rect 2502 783 2508 784
rect 1326 778 1332 779
rect 1422 780 1428 781
rect 150 776 156 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 150 772 151 776
rect 155 772 156 776
rect 150 771 156 772
rect 246 776 252 777
rect 246 772 247 776
rect 251 772 252 776
rect 246 771 252 772
rect 342 776 348 777
rect 342 772 343 776
rect 347 772 348 776
rect 342 771 348 772
rect 438 776 444 777
rect 438 772 439 776
rect 443 772 444 776
rect 438 771 444 772
rect 526 776 532 777
rect 526 772 527 776
rect 531 772 532 776
rect 526 771 532 772
rect 606 776 612 777
rect 606 772 607 776
rect 611 772 612 776
rect 606 771 612 772
rect 678 776 684 777
rect 678 772 679 776
rect 683 772 684 776
rect 678 771 684 772
rect 750 776 756 777
rect 750 772 751 776
rect 755 772 756 776
rect 750 771 756 772
rect 822 776 828 777
rect 822 772 823 776
rect 827 772 828 776
rect 822 771 828 772
rect 894 776 900 777
rect 894 772 895 776
rect 899 772 900 776
rect 894 771 900 772
rect 974 776 980 777
rect 974 772 975 776
rect 979 772 980 776
rect 1422 776 1423 780
rect 1427 776 1428 780
rect 1422 775 1428 776
rect 1494 780 1500 781
rect 1494 776 1495 780
rect 1499 776 1500 780
rect 1494 775 1500 776
rect 1574 780 1580 781
rect 1574 776 1575 780
rect 1579 776 1580 780
rect 1574 775 1580 776
rect 1654 780 1660 781
rect 1654 776 1655 780
rect 1659 776 1660 780
rect 1654 775 1660 776
rect 1742 780 1748 781
rect 1742 776 1743 780
rect 1747 776 1748 780
rect 1742 775 1748 776
rect 1830 780 1836 781
rect 1830 776 1831 780
rect 1835 776 1836 780
rect 1830 775 1836 776
rect 1918 780 1924 781
rect 1918 776 1919 780
rect 1923 776 1924 780
rect 1918 775 1924 776
rect 2006 780 2012 781
rect 2006 776 2007 780
rect 2011 776 2012 780
rect 2006 775 2012 776
rect 2094 780 2100 781
rect 2094 776 2095 780
rect 2099 776 2100 780
rect 2094 775 2100 776
rect 2182 780 2188 781
rect 2182 776 2183 780
rect 2187 776 2188 780
rect 2182 775 2188 776
rect 2270 780 2276 781
rect 2270 776 2271 780
rect 2275 776 2276 780
rect 2270 775 2276 776
rect 2366 780 2372 781
rect 2366 776 2367 780
rect 2371 776 2372 780
rect 2366 775 2372 776
rect 2438 780 2444 781
rect 2438 776 2439 780
rect 2443 776 2444 780
rect 2502 779 2503 783
rect 2507 779 2508 783
rect 2502 778 2508 779
rect 2438 775 2444 776
rect 974 771 980 772
rect 1286 773 1292 774
rect 110 768 116 769
rect 1286 769 1287 773
rect 1291 769 1292 773
rect 1286 768 1292 769
rect 1350 764 1356 765
rect 1326 761 1332 762
rect 1326 757 1327 761
rect 1331 757 1332 761
rect 1350 760 1351 764
rect 1355 760 1356 764
rect 1350 759 1356 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1566 764 1572 765
rect 1566 760 1567 764
rect 1571 760 1572 764
rect 1566 759 1572 760
rect 1686 764 1692 765
rect 1686 760 1687 764
rect 1691 760 1692 764
rect 1686 759 1692 760
rect 1806 764 1812 765
rect 1806 760 1807 764
rect 1811 760 1812 764
rect 1806 759 1812 760
rect 1926 764 1932 765
rect 1926 760 1927 764
rect 1931 760 1932 764
rect 1926 759 1932 760
rect 2038 764 2044 765
rect 2038 760 2039 764
rect 2043 760 2044 764
rect 2038 759 2044 760
rect 2142 764 2148 765
rect 2142 760 2143 764
rect 2147 760 2148 764
rect 2142 759 2148 760
rect 2246 764 2252 765
rect 2246 760 2247 764
rect 2251 760 2252 764
rect 2246 759 2252 760
rect 2350 764 2356 765
rect 2350 760 2351 764
rect 2355 760 2356 764
rect 2350 759 2356 760
rect 2438 764 2444 765
rect 2438 760 2439 764
rect 2443 760 2444 764
rect 2438 759 2444 760
rect 2502 761 2508 762
rect 110 756 116 757
rect 1286 756 1292 757
rect 1326 756 1332 757
rect 2502 757 2503 761
rect 2507 757 2508 761
rect 2502 756 2508 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 166 750 172 751
rect 262 755 268 756
rect 262 751 263 755
rect 267 751 268 755
rect 262 750 268 751
rect 358 755 364 756
rect 358 751 359 755
rect 363 751 364 755
rect 358 750 364 751
rect 454 755 460 756
rect 454 751 455 755
rect 459 751 460 755
rect 454 750 460 751
rect 542 755 548 756
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 694 755 700 756
rect 694 751 695 755
rect 699 751 700 755
rect 694 750 700 751
rect 766 755 772 756
rect 766 751 767 755
rect 771 751 772 755
rect 766 750 772 751
rect 838 755 844 756
rect 838 751 839 755
rect 843 751 844 755
rect 838 750 844 751
rect 910 755 916 756
rect 910 751 911 755
rect 915 751 916 755
rect 910 750 916 751
rect 990 755 996 756
rect 990 751 991 755
rect 995 751 996 755
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 990 750 996 751
rect 1326 744 1332 745
rect 2502 744 2508 745
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 1326 739 1332 740
rect 1366 743 1372 744
rect 1366 739 1367 743
rect 1371 739 1372 743
rect 1366 738 1372 739
rect 1462 743 1468 744
rect 1462 739 1463 743
rect 1467 739 1468 743
rect 1462 738 1468 739
rect 1582 743 1588 744
rect 1582 739 1583 743
rect 1587 739 1588 743
rect 1582 738 1588 739
rect 1702 743 1708 744
rect 1702 739 1703 743
rect 1707 739 1708 743
rect 1702 738 1708 739
rect 1822 743 1828 744
rect 1822 739 1823 743
rect 1827 739 1828 743
rect 1822 738 1828 739
rect 1942 743 1948 744
rect 1942 739 1943 743
rect 1947 739 1948 743
rect 1942 738 1948 739
rect 2054 743 2060 744
rect 2054 739 2055 743
rect 2059 739 2060 743
rect 2054 738 2060 739
rect 2158 743 2164 744
rect 2158 739 2159 743
rect 2163 739 2164 743
rect 2158 738 2164 739
rect 2262 743 2268 744
rect 2262 739 2263 743
rect 2267 739 2268 743
rect 2262 738 2268 739
rect 2366 743 2372 744
rect 2366 739 2367 743
rect 2371 739 2372 743
rect 2366 738 2372 739
rect 2454 743 2460 744
rect 2454 739 2455 743
rect 2459 739 2460 743
rect 2502 740 2503 744
rect 2507 740 2508 744
rect 2502 739 2508 740
rect 2454 738 2460 739
rect 174 701 180 702
rect 110 700 116 701
rect 110 696 111 700
rect 115 696 116 700
rect 174 697 175 701
rect 179 697 180 701
rect 174 696 180 697
rect 262 701 268 702
rect 262 697 263 701
rect 267 697 268 701
rect 262 696 268 697
rect 342 701 348 702
rect 342 697 343 701
rect 347 697 348 701
rect 342 696 348 697
rect 422 701 428 702
rect 422 697 423 701
rect 427 697 428 701
rect 422 696 428 697
rect 502 701 508 702
rect 502 697 503 701
rect 507 697 508 701
rect 502 696 508 697
rect 574 701 580 702
rect 574 697 575 701
rect 579 697 580 701
rect 574 696 580 697
rect 638 701 644 702
rect 638 697 639 701
rect 643 697 644 701
rect 638 696 644 697
rect 702 701 708 702
rect 702 697 703 701
rect 707 697 708 701
rect 702 696 708 697
rect 766 701 772 702
rect 766 697 767 701
rect 771 697 772 701
rect 766 696 772 697
rect 838 701 844 702
rect 838 697 839 701
rect 843 697 844 701
rect 838 696 844 697
rect 910 701 916 702
rect 910 697 911 701
rect 915 697 916 701
rect 910 696 916 697
rect 1286 700 1292 701
rect 1286 696 1287 700
rect 1291 696 1292 700
rect 110 695 116 696
rect 1286 695 1292 696
rect 1366 689 1372 690
rect 1326 688 1332 689
rect 1326 684 1327 688
rect 1331 684 1332 688
rect 1366 685 1367 689
rect 1371 685 1372 689
rect 1366 684 1372 685
rect 1430 689 1436 690
rect 1430 685 1431 689
rect 1435 685 1436 689
rect 1430 684 1436 685
rect 1534 689 1540 690
rect 1534 685 1535 689
rect 1539 685 1540 689
rect 1534 684 1540 685
rect 1638 689 1644 690
rect 1638 685 1639 689
rect 1643 685 1644 689
rect 1638 684 1644 685
rect 1750 689 1756 690
rect 1750 685 1751 689
rect 1755 685 1756 689
rect 1750 684 1756 685
rect 1862 689 1868 690
rect 1862 685 1863 689
rect 1867 685 1868 689
rect 1862 684 1868 685
rect 1966 689 1972 690
rect 1966 685 1967 689
rect 1971 685 1972 689
rect 1966 684 1972 685
rect 2062 689 2068 690
rect 2062 685 2063 689
rect 2067 685 2068 689
rect 2062 684 2068 685
rect 2150 689 2156 690
rect 2150 685 2151 689
rect 2155 685 2156 689
rect 2150 684 2156 685
rect 2230 689 2236 690
rect 2230 685 2231 689
rect 2235 685 2236 689
rect 2230 684 2236 685
rect 2310 689 2316 690
rect 2310 685 2311 689
rect 2315 685 2316 689
rect 2310 684 2316 685
rect 2390 689 2396 690
rect 2390 685 2391 689
rect 2395 685 2396 689
rect 2390 684 2396 685
rect 2454 689 2460 690
rect 2454 685 2455 689
rect 2459 685 2460 689
rect 2454 684 2460 685
rect 2502 688 2508 689
rect 2502 684 2503 688
rect 2507 684 2508 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1286 683 1292 684
rect 1326 683 1332 684
rect 2502 683 2508 684
rect 110 678 116 679
rect 158 680 164 681
rect 158 676 159 680
rect 163 676 164 680
rect 158 675 164 676
rect 246 680 252 681
rect 246 676 247 680
rect 251 676 252 680
rect 246 675 252 676
rect 326 680 332 681
rect 326 676 327 680
rect 331 676 332 680
rect 326 675 332 676
rect 406 680 412 681
rect 406 676 407 680
rect 411 676 412 680
rect 406 675 412 676
rect 486 680 492 681
rect 486 676 487 680
rect 491 676 492 680
rect 486 675 492 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 686 680 692 681
rect 686 676 687 680
rect 691 676 692 680
rect 686 675 692 676
rect 750 680 756 681
rect 750 676 751 680
rect 755 676 756 680
rect 750 675 756 676
rect 822 680 828 681
rect 822 676 823 680
rect 827 676 828 680
rect 822 675 828 676
rect 894 680 900 681
rect 894 676 895 680
rect 899 676 900 680
rect 1286 679 1287 683
rect 1291 679 1292 683
rect 1286 678 1292 679
rect 894 675 900 676
rect 1326 671 1332 672
rect 214 668 220 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 214 664 215 668
rect 219 664 220 668
rect 214 663 220 664
rect 294 668 300 669
rect 294 664 295 668
rect 299 664 300 668
rect 294 663 300 664
rect 374 668 380 669
rect 374 664 375 668
rect 379 664 380 668
rect 374 663 380 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 526 668 532 669
rect 526 664 527 668
rect 531 664 532 668
rect 526 663 532 664
rect 590 668 596 669
rect 590 664 591 668
rect 595 664 596 668
rect 590 663 596 664
rect 654 668 660 669
rect 654 664 655 668
rect 659 664 660 668
rect 654 663 660 664
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 782 668 788 669
rect 782 664 783 668
rect 787 664 788 668
rect 782 663 788 664
rect 846 668 852 669
rect 846 664 847 668
rect 851 664 852 668
rect 846 663 852 664
rect 918 668 924 669
rect 918 664 919 668
rect 923 664 924 668
rect 1326 667 1327 671
rect 1331 667 1332 671
rect 2502 671 2508 672
rect 1326 666 1332 667
rect 1350 668 1356 669
rect 918 663 924 664
rect 1286 665 1292 666
rect 110 660 116 661
rect 1286 661 1287 665
rect 1291 661 1292 665
rect 1350 664 1351 668
rect 1355 664 1356 668
rect 1350 663 1356 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1414 663 1420 664
rect 1518 668 1524 669
rect 1518 664 1519 668
rect 1523 664 1524 668
rect 1518 663 1524 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1734 668 1740 669
rect 1734 664 1735 668
rect 1739 664 1740 668
rect 1734 663 1740 664
rect 1846 668 1852 669
rect 1846 664 1847 668
rect 1851 664 1852 668
rect 1846 663 1852 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2134 668 2140 669
rect 2134 664 2135 668
rect 2139 664 2140 668
rect 2134 663 2140 664
rect 2214 668 2220 669
rect 2214 664 2215 668
rect 2219 664 2220 668
rect 2214 663 2220 664
rect 2294 668 2300 669
rect 2294 664 2295 668
rect 2299 664 2300 668
rect 2294 663 2300 664
rect 2374 668 2380 669
rect 2374 664 2375 668
rect 2379 664 2380 668
rect 2374 663 2380 664
rect 2438 668 2444 669
rect 2438 664 2439 668
rect 2443 664 2444 668
rect 2502 667 2503 671
rect 2507 667 2508 671
rect 2502 666 2508 667
rect 2438 663 2444 664
rect 1286 660 1292 661
rect 110 648 116 649
rect 1286 648 1292 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 230 647 236 648
rect 230 643 231 647
rect 235 643 236 647
rect 230 642 236 643
rect 310 647 316 648
rect 310 643 311 647
rect 315 643 316 647
rect 310 642 316 643
rect 390 647 396 648
rect 390 643 391 647
rect 395 643 396 647
rect 390 642 396 643
rect 470 647 476 648
rect 470 643 471 647
rect 475 643 476 647
rect 470 642 476 643
rect 542 647 548 648
rect 542 643 543 647
rect 547 643 548 647
rect 542 642 548 643
rect 606 647 612 648
rect 606 643 607 647
rect 611 643 612 647
rect 606 642 612 643
rect 670 647 676 648
rect 670 643 671 647
rect 675 643 676 647
rect 670 642 676 643
rect 734 647 740 648
rect 734 643 735 647
rect 739 643 740 647
rect 734 642 740 643
rect 798 647 804 648
rect 798 643 799 647
rect 803 643 804 647
rect 798 642 804 643
rect 862 647 868 648
rect 862 643 863 647
rect 867 643 868 647
rect 862 642 868 643
rect 934 647 940 648
rect 934 643 935 647
rect 939 643 940 647
rect 1286 644 1287 648
rect 1291 644 1292 648
rect 1478 648 1484 649
rect 1286 643 1292 644
rect 1326 645 1332 646
rect 934 642 940 643
rect 1326 641 1327 645
rect 1331 641 1332 645
rect 1478 644 1479 648
rect 1483 644 1484 648
rect 1478 643 1484 644
rect 1558 648 1564 649
rect 1558 644 1559 648
rect 1563 644 1564 648
rect 1558 643 1564 644
rect 1646 648 1652 649
rect 1646 644 1647 648
rect 1651 644 1652 648
rect 1646 643 1652 644
rect 1734 648 1740 649
rect 1734 644 1735 648
rect 1739 644 1740 648
rect 1734 643 1740 644
rect 1830 648 1836 649
rect 1830 644 1831 648
rect 1835 644 1836 648
rect 1830 643 1836 644
rect 1918 648 1924 649
rect 1918 644 1919 648
rect 1923 644 1924 648
rect 1918 643 1924 644
rect 2006 648 2012 649
rect 2006 644 2007 648
rect 2011 644 2012 648
rect 2006 643 2012 644
rect 2086 648 2092 649
rect 2086 644 2087 648
rect 2091 644 2092 648
rect 2086 643 2092 644
rect 2166 648 2172 649
rect 2166 644 2167 648
rect 2171 644 2172 648
rect 2166 643 2172 644
rect 2238 648 2244 649
rect 2238 644 2239 648
rect 2243 644 2244 648
rect 2238 643 2244 644
rect 2310 648 2316 649
rect 2310 644 2311 648
rect 2315 644 2316 648
rect 2310 643 2316 644
rect 2382 648 2388 649
rect 2382 644 2383 648
rect 2387 644 2388 648
rect 2382 643 2388 644
rect 2438 648 2444 649
rect 2438 644 2439 648
rect 2443 644 2444 648
rect 2438 643 2444 644
rect 2502 645 2508 646
rect 1326 640 1332 641
rect 2502 641 2503 645
rect 2507 641 2508 645
rect 2502 640 2508 641
rect 1326 628 1332 629
rect 2502 628 2508 629
rect 1326 624 1327 628
rect 1331 624 1332 628
rect 1326 623 1332 624
rect 1494 627 1500 628
rect 1494 623 1495 627
rect 1499 623 1500 627
rect 1494 622 1500 623
rect 1574 627 1580 628
rect 1574 623 1575 627
rect 1579 623 1580 627
rect 1574 622 1580 623
rect 1662 627 1668 628
rect 1662 623 1663 627
rect 1667 623 1668 627
rect 1662 622 1668 623
rect 1750 627 1756 628
rect 1750 623 1751 627
rect 1755 623 1756 627
rect 1750 622 1756 623
rect 1846 627 1852 628
rect 1846 623 1847 627
rect 1851 623 1852 627
rect 1846 622 1852 623
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 1934 622 1940 623
rect 2022 627 2028 628
rect 2022 623 2023 627
rect 2027 623 2028 627
rect 2022 622 2028 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2182 627 2188 628
rect 2182 623 2183 627
rect 2187 623 2188 627
rect 2182 622 2188 623
rect 2254 627 2260 628
rect 2254 623 2255 627
rect 2259 623 2260 627
rect 2254 622 2260 623
rect 2326 627 2332 628
rect 2326 623 2327 627
rect 2331 623 2332 627
rect 2326 622 2332 623
rect 2398 627 2404 628
rect 2398 623 2399 627
rect 2403 623 2404 627
rect 2398 622 2404 623
rect 2454 627 2460 628
rect 2454 623 2455 627
rect 2459 623 2460 627
rect 2502 624 2503 628
rect 2507 624 2508 628
rect 2502 623 2508 624
rect 2454 622 2460 623
rect 206 593 212 594
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 206 589 207 593
rect 211 589 212 593
rect 206 588 212 589
rect 302 593 308 594
rect 302 589 303 593
rect 307 589 308 593
rect 302 588 308 589
rect 406 593 412 594
rect 406 589 407 593
rect 411 589 412 593
rect 406 588 412 589
rect 502 593 508 594
rect 502 589 503 593
rect 507 589 508 593
rect 502 588 508 589
rect 598 593 604 594
rect 598 589 599 593
rect 603 589 604 593
rect 598 588 604 589
rect 686 593 692 594
rect 686 589 687 593
rect 691 589 692 593
rect 686 588 692 589
rect 766 593 772 594
rect 766 589 767 593
rect 771 589 772 593
rect 766 588 772 589
rect 846 593 852 594
rect 846 589 847 593
rect 851 589 852 593
rect 846 588 852 589
rect 926 593 932 594
rect 926 589 927 593
rect 931 589 932 593
rect 926 588 932 589
rect 1006 593 1012 594
rect 1006 589 1007 593
rect 1011 589 1012 593
rect 1006 588 1012 589
rect 1086 593 1092 594
rect 1086 589 1087 593
rect 1091 589 1092 593
rect 1086 588 1092 589
rect 1286 592 1292 593
rect 1286 588 1287 592
rect 1291 588 1292 592
rect 110 587 116 588
rect 1286 587 1292 588
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1286 575 1292 576
rect 110 570 116 571
rect 190 572 196 573
rect 190 568 191 572
rect 195 568 196 572
rect 190 567 196 568
rect 286 572 292 573
rect 286 568 287 572
rect 291 568 292 572
rect 286 567 292 568
rect 390 572 396 573
rect 390 568 391 572
rect 395 568 396 572
rect 390 567 396 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 670 572 676 573
rect 670 568 671 572
rect 675 568 676 572
rect 670 567 676 568
rect 750 572 756 573
rect 750 568 751 572
rect 755 568 756 572
rect 750 567 756 568
rect 830 572 836 573
rect 830 568 831 572
rect 835 568 836 572
rect 830 567 836 568
rect 910 572 916 573
rect 910 568 911 572
rect 915 568 916 572
rect 910 567 916 568
rect 990 572 996 573
rect 990 568 991 572
rect 995 568 996 572
rect 990 567 996 568
rect 1070 572 1076 573
rect 1070 568 1071 572
rect 1075 568 1076 572
rect 1286 571 1287 575
rect 1291 571 1292 575
rect 1454 573 1460 574
rect 1286 570 1292 571
rect 1326 572 1332 573
rect 1070 567 1076 568
rect 1326 568 1327 572
rect 1331 568 1332 572
rect 1454 569 1455 573
rect 1459 569 1460 573
rect 1454 568 1460 569
rect 1558 573 1564 574
rect 1558 569 1559 573
rect 1563 569 1564 573
rect 1558 568 1564 569
rect 1670 573 1676 574
rect 1670 569 1671 573
rect 1675 569 1676 573
rect 1670 568 1676 569
rect 1774 573 1780 574
rect 1774 569 1775 573
rect 1779 569 1780 573
rect 1774 568 1780 569
rect 1878 573 1884 574
rect 1878 569 1879 573
rect 1883 569 1884 573
rect 1878 568 1884 569
rect 1982 573 1988 574
rect 1982 569 1983 573
rect 1987 569 1988 573
rect 1982 568 1988 569
rect 2086 573 2092 574
rect 2086 569 2087 573
rect 2091 569 2092 573
rect 2086 568 2092 569
rect 2182 573 2188 574
rect 2182 569 2183 573
rect 2187 569 2188 573
rect 2182 568 2188 569
rect 2278 573 2284 574
rect 2278 569 2279 573
rect 2283 569 2284 573
rect 2278 568 2284 569
rect 2374 573 2380 574
rect 2374 569 2375 573
rect 2379 569 2380 573
rect 2374 568 2380 569
rect 2454 573 2460 574
rect 2454 569 2455 573
rect 2459 569 2460 573
rect 2454 568 2460 569
rect 2502 572 2508 573
rect 2502 568 2503 572
rect 2507 568 2508 572
rect 1326 567 1332 568
rect 2502 567 2508 568
rect 174 556 180 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 270 556 276 557
rect 270 552 271 556
rect 275 552 276 556
rect 270 551 276 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 486 556 492 557
rect 486 552 487 556
rect 491 552 492 556
rect 486 551 492 552
rect 590 556 596 557
rect 590 552 591 556
rect 595 552 596 556
rect 590 551 596 552
rect 694 556 700 557
rect 694 552 695 556
rect 699 552 700 556
rect 694 551 700 552
rect 790 556 796 557
rect 790 552 791 556
rect 795 552 796 556
rect 790 551 796 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 966 556 972 557
rect 966 552 967 556
rect 971 552 972 556
rect 966 551 972 552
rect 1054 556 1060 557
rect 1054 552 1055 556
rect 1059 552 1060 556
rect 1054 551 1060 552
rect 1150 556 1156 557
rect 1150 552 1151 556
rect 1155 552 1156 556
rect 1326 555 1332 556
rect 1150 551 1156 552
rect 1286 553 1292 554
rect 110 548 116 549
rect 1286 549 1287 553
rect 1291 549 1292 553
rect 1326 551 1327 555
rect 1331 551 1332 555
rect 2502 555 2508 556
rect 1326 550 1332 551
rect 1438 552 1444 553
rect 1286 548 1292 549
rect 1438 548 1439 552
rect 1443 548 1444 552
rect 1438 547 1444 548
rect 1542 552 1548 553
rect 1542 548 1543 552
rect 1547 548 1548 552
rect 1542 547 1548 548
rect 1654 552 1660 553
rect 1654 548 1655 552
rect 1659 548 1660 552
rect 1654 547 1660 548
rect 1758 552 1764 553
rect 1758 548 1759 552
rect 1763 548 1764 552
rect 1758 547 1764 548
rect 1862 552 1868 553
rect 1862 548 1863 552
rect 1867 548 1868 552
rect 1862 547 1868 548
rect 1966 552 1972 553
rect 1966 548 1967 552
rect 1971 548 1972 552
rect 1966 547 1972 548
rect 2070 552 2076 553
rect 2070 548 2071 552
rect 2075 548 2076 552
rect 2070 547 2076 548
rect 2166 552 2172 553
rect 2166 548 2167 552
rect 2171 548 2172 552
rect 2166 547 2172 548
rect 2262 552 2268 553
rect 2262 548 2263 552
rect 2267 548 2268 552
rect 2262 547 2268 548
rect 2358 552 2364 553
rect 2358 548 2359 552
rect 2363 548 2364 552
rect 2358 547 2364 548
rect 2438 552 2444 553
rect 2438 548 2439 552
rect 2443 548 2444 552
rect 2502 551 2503 555
rect 2507 551 2508 555
rect 2502 550 2508 551
rect 2438 547 2444 548
rect 110 536 116 537
rect 1286 536 1292 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 190 535 196 536
rect 190 531 191 535
rect 195 531 196 535
rect 190 530 196 531
rect 286 535 292 536
rect 286 531 287 535
rect 291 531 292 535
rect 286 530 292 531
rect 390 535 396 536
rect 390 531 391 535
rect 395 531 396 535
rect 390 530 396 531
rect 502 535 508 536
rect 502 531 503 535
rect 507 531 508 535
rect 502 530 508 531
rect 606 535 612 536
rect 606 531 607 535
rect 611 531 612 535
rect 606 530 612 531
rect 710 535 716 536
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 806 535 812 536
rect 806 531 807 535
rect 811 531 812 535
rect 806 530 812 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 982 535 988 536
rect 982 531 983 535
rect 987 531 988 535
rect 982 530 988 531
rect 1070 535 1076 536
rect 1070 531 1071 535
rect 1075 531 1076 535
rect 1070 530 1076 531
rect 1166 535 1172 536
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1286 532 1287 536
rect 1291 532 1292 536
rect 1366 536 1372 537
rect 1286 531 1292 532
rect 1326 533 1332 534
rect 1166 530 1172 531
rect 1326 529 1327 533
rect 1331 529 1332 533
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1446 536 1452 537
rect 1446 532 1447 536
rect 1451 532 1452 536
rect 1446 531 1452 532
rect 1526 536 1532 537
rect 1526 532 1527 536
rect 1531 532 1532 536
rect 1526 531 1532 532
rect 1614 536 1620 537
rect 1614 532 1615 536
rect 1619 532 1620 536
rect 1614 531 1620 532
rect 1710 536 1716 537
rect 1710 532 1711 536
rect 1715 532 1716 536
rect 1710 531 1716 532
rect 1798 536 1804 537
rect 1798 532 1799 536
rect 1803 532 1804 536
rect 1798 531 1804 532
rect 1886 536 1892 537
rect 1886 532 1887 536
rect 1891 532 1892 536
rect 1886 531 1892 532
rect 1974 536 1980 537
rect 1974 532 1975 536
rect 1979 532 1980 536
rect 1974 531 1980 532
rect 2062 536 2068 537
rect 2062 532 2063 536
rect 2067 532 2068 536
rect 2062 531 2068 532
rect 2150 536 2156 537
rect 2150 532 2151 536
rect 2155 532 2156 536
rect 2150 531 2156 532
rect 2246 536 2252 537
rect 2246 532 2247 536
rect 2251 532 2252 536
rect 2246 531 2252 532
rect 2342 536 2348 537
rect 2342 532 2343 536
rect 2347 532 2348 536
rect 2342 531 2348 532
rect 2438 536 2444 537
rect 2438 532 2439 536
rect 2443 532 2444 536
rect 2438 531 2444 532
rect 2502 533 2508 534
rect 1326 528 1332 529
rect 2502 529 2503 533
rect 2507 529 2508 533
rect 2502 528 2508 529
rect 1326 516 1332 517
rect 2502 516 2508 517
rect 1326 512 1327 516
rect 1331 512 1332 516
rect 1326 511 1332 512
rect 1382 515 1388 516
rect 1382 511 1383 515
rect 1387 511 1388 515
rect 1382 510 1388 511
rect 1462 515 1468 516
rect 1462 511 1463 515
rect 1467 511 1468 515
rect 1462 510 1468 511
rect 1542 515 1548 516
rect 1542 511 1543 515
rect 1547 511 1548 515
rect 1542 510 1548 511
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 1726 515 1732 516
rect 1726 511 1727 515
rect 1731 511 1732 515
rect 1726 510 1732 511
rect 1814 515 1820 516
rect 1814 511 1815 515
rect 1819 511 1820 515
rect 1814 510 1820 511
rect 1902 515 1908 516
rect 1902 511 1903 515
rect 1907 511 1908 515
rect 1902 510 1908 511
rect 1990 515 1996 516
rect 1990 511 1991 515
rect 1995 511 1996 515
rect 1990 510 1996 511
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2166 515 2172 516
rect 2166 511 2167 515
rect 2171 511 2172 515
rect 2166 510 2172 511
rect 2262 515 2268 516
rect 2262 511 2263 515
rect 2267 511 2268 515
rect 2262 510 2268 511
rect 2358 515 2364 516
rect 2358 511 2359 515
rect 2363 511 2364 515
rect 2358 510 2364 511
rect 2454 515 2460 516
rect 2454 511 2455 515
rect 2459 511 2460 515
rect 2502 512 2503 516
rect 2507 512 2508 516
rect 2502 511 2508 512
rect 2454 510 2460 511
rect 150 481 156 482
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 150 477 151 481
rect 155 477 156 481
rect 150 476 156 477
rect 246 481 252 482
rect 246 477 247 481
rect 251 477 252 481
rect 246 476 252 477
rect 366 481 372 482
rect 366 477 367 481
rect 371 477 372 481
rect 366 476 372 477
rect 486 481 492 482
rect 486 477 487 481
rect 491 477 492 481
rect 486 476 492 477
rect 614 481 620 482
rect 614 477 615 481
rect 619 477 620 481
rect 614 476 620 477
rect 734 481 740 482
rect 734 477 735 481
rect 739 477 740 481
rect 734 476 740 477
rect 846 481 852 482
rect 846 477 847 481
rect 851 477 852 481
rect 846 476 852 477
rect 950 481 956 482
rect 950 477 951 481
rect 955 477 956 481
rect 950 476 956 477
rect 1054 481 1060 482
rect 1054 477 1055 481
rect 1059 477 1060 481
rect 1054 476 1060 477
rect 1158 481 1164 482
rect 1158 477 1159 481
rect 1163 477 1164 481
rect 1158 476 1164 477
rect 1238 481 1244 482
rect 1238 477 1239 481
rect 1243 477 1244 481
rect 1238 476 1244 477
rect 1286 480 1292 481
rect 1286 476 1287 480
rect 1291 476 1292 480
rect 110 475 116 476
rect 1286 475 1292 476
rect 110 463 116 464
rect 110 459 111 463
rect 115 459 116 463
rect 1286 463 1292 464
rect 110 458 116 459
rect 134 460 140 461
rect 134 456 135 460
rect 139 456 140 460
rect 134 455 140 456
rect 230 460 236 461
rect 230 456 231 460
rect 235 456 236 460
rect 230 455 236 456
rect 350 460 356 461
rect 350 456 351 460
rect 355 456 356 460
rect 350 455 356 456
rect 470 460 476 461
rect 470 456 471 460
rect 475 456 476 460
rect 470 455 476 456
rect 598 460 604 461
rect 598 456 599 460
rect 603 456 604 460
rect 598 455 604 456
rect 718 460 724 461
rect 718 456 719 460
rect 723 456 724 460
rect 718 455 724 456
rect 830 460 836 461
rect 830 456 831 460
rect 835 456 836 460
rect 830 455 836 456
rect 934 460 940 461
rect 934 456 935 460
rect 939 456 940 460
rect 934 455 940 456
rect 1038 460 1044 461
rect 1038 456 1039 460
rect 1043 456 1044 460
rect 1038 455 1044 456
rect 1142 460 1148 461
rect 1142 456 1143 460
rect 1147 456 1148 460
rect 1142 455 1148 456
rect 1222 460 1228 461
rect 1222 456 1223 460
rect 1227 456 1228 460
rect 1286 459 1287 463
rect 1291 459 1292 463
rect 1366 461 1372 462
rect 1286 458 1292 459
rect 1326 460 1332 461
rect 1222 455 1228 456
rect 1326 456 1327 460
rect 1331 456 1332 460
rect 1366 457 1367 461
rect 1371 457 1372 461
rect 1366 456 1372 457
rect 1430 461 1436 462
rect 1430 457 1431 461
rect 1435 457 1436 461
rect 1430 456 1436 457
rect 1518 461 1524 462
rect 1518 457 1519 461
rect 1523 457 1524 461
rect 1518 456 1524 457
rect 1614 461 1620 462
rect 1614 457 1615 461
rect 1619 457 1620 461
rect 1614 456 1620 457
rect 1710 461 1716 462
rect 1710 457 1711 461
rect 1715 457 1716 461
rect 1710 456 1716 457
rect 1814 461 1820 462
rect 1814 457 1815 461
rect 1819 457 1820 461
rect 1814 456 1820 457
rect 1926 461 1932 462
rect 1926 457 1927 461
rect 1931 457 1932 461
rect 1926 456 1932 457
rect 2054 461 2060 462
rect 2054 457 2055 461
rect 2059 457 2060 461
rect 2054 456 2060 457
rect 2190 461 2196 462
rect 2190 457 2191 461
rect 2195 457 2196 461
rect 2190 456 2196 457
rect 2334 461 2340 462
rect 2334 457 2335 461
rect 2339 457 2340 461
rect 2334 456 2340 457
rect 2454 461 2460 462
rect 2454 457 2455 461
rect 2459 457 2460 461
rect 2454 456 2460 457
rect 2502 460 2508 461
rect 2502 456 2503 460
rect 2507 456 2508 460
rect 1326 455 1332 456
rect 2502 455 2508 456
rect 134 444 140 445
rect 110 441 116 442
rect 110 437 111 441
rect 115 437 116 441
rect 134 440 135 444
rect 139 440 140 444
rect 134 439 140 440
rect 190 444 196 445
rect 190 440 191 444
rect 195 440 196 444
rect 190 439 196 440
rect 246 444 252 445
rect 246 440 247 444
rect 251 440 252 444
rect 246 439 252 440
rect 302 444 308 445
rect 302 440 303 444
rect 307 440 308 444
rect 302 439 308 440
rect 382 444 388 445
rect 382 440 383 444
rect 387 440 388 444
rect 382 439 388 440
rect 470 444 476 445
rect 470 440 471 444
rect 475 440 476 444
rect 470 439 476 440
rect 566 444 572 445
rect 566 440 567 444
rect 571 440 572 444
rect 566 439 572 440
rect 670 444 676 445
rect 670 440 671 444
rect 675 440 676 444
rect 670 439 676 440
rect 782 444 788 445
rect 782 440 783 444
rect 787 440 788 444
rect 782 439 788 440
rect 894 444 900 445
rect 894 440 895 444
rect 899 440 900 444
rect 894 439 900 440
rect 1006 444 1012 445
rect 1006 440 1007 444
rect 1011 440 1012 444
rect 1006 439 1012 440
rect 1126 444 1132 445
rect 1126 440 1127 444
rect 1131 440 1132 444
rect 1126 439 1132 440
rect 1222 444 1228 445
rect 1222 440 1223 444
rect 1227 440 1228 444
rect 1326 443 1332 444
rect 1222 439 1228 440
rect 1286 441 1292 442
rect 110 436 116 437
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1326 439 1327 443
rect 1331 439 1332 443
rect 2502 443 2508 444
rect 1326 438 1332 439
rect 1350 440 1356 441
rect 1286 436 1292 437
rect 1350 436 1351 440
rect 1355 436 1356 440
rect 1350 435 1356 436
rect 1414 440 1420 441
rect 1414 436 1415 440
rect 1419 436 1420 440
rect 1414 435 1420 436
rect 1502 440 1508 441
rect 1502 436 1503 440
rect 1507 436 1508 440
rect 1502 435 1508 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1694 440 1700 441
rect 1694 436 1695 440
rect 1699 436 1700 440
rect 1694 435 1700 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1910 440 1916 441
rect 1910 436 1911 440
rect 1915 436 1916 440
rect 1910 435 1916 436
rect 2038 440 2044 441
rect 2038 436 2039 440
rect 2043 436 2044 440
rect 2038 435 2044 436
rect 2174 440 2180 441
rect 2174 436 2175 440
rect 2179 436 2180 440
rect 2174 435 2180 436
rect 2318 440 2324 441
rect 2318 436 2319 440
rect 2323 436 2324 440
rect 2318 435 2324 436
rect 2438 440 2444 441
rect 2438 436 2439 440
rect 2443 436 2444 440
rect 2502 439 2503 443
rect 2507 439 2508 443
rect 2502 438 2508 439
rect 2438 435 2444 436
rect 110 424 116 425
rect 1286 424 1292 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 150 423 156 424
rect 150 419 151 423
rect 155 419 156 423
rect 150 418 156 419
rect 206 423 212 424
rect 206 419 207 423
rect 211 419 212 423
rect 206 418 212 419
rect 262 423 268 424
rect 262 419 263 423
rect 267 419 268 423
rect 262 418 268 419
rect 318 423 324 424
rect 318 419 319 423
rect 323 419 324 423
rect 318 418 324 419
rect 398 423 404 424
rect 398 419 399 423
rect 403 419 404 423
rect 398 418 404 419
rect 486 423 492 424
rect 486 419 487 423
rect 491 419 492 423
rect 486 418 492 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 686 423 692 424
rect 686 419 687 423
rect 691 419 692 423
rect 686 418 692 419
rect 798 423 804 424
rect 798 419 799 423
rect 803 419 804 423
rect 798 418 804 419
rect 910 423 916 424
rect 910 419 911 423
rect 915 419 916 423
rect 910 418 916 419
rect 1022 423 1028 424
rect 1022 419 1023 423
rect 1027 419 1028 423
rect 1022 418 1028 419
rect 1142 423 1148 424
rect 1142 419 1143 423
rect 1147 419 1148 423
rect 1142 418 1148 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1286 420 1287 424
rect 1291 420 1292 424
rect 1350 424 1356 425
rect 1286 419 1292 420
rect 1326 421 1332 422
rect 1238 418 1244 419
rect 1326 417 1327 421
rect 1331 417 1332 421
rect 1350 420 1351 424
rect 1355 420 1356 424
rect 1350 419 1356 420
rect 1422 424 1428 425
rect 1422 420 1423 424
rect 1427 420 1428 424
rect 1422 419 1428 420
rect 1510 424 1516 425
rect 1510 420 1511 424
rect 1515 420 1516 424
rect 1510 419 1516 420
rect 1598 424 1604 425
rect 1598 420 1599 424
rect 1603 420 1604 424
rect 1598 419 1604 420
rect 1678 424 1684 425
rect 1678 420 1679 424
rect 1683 420 1684 424
rect 1678 419 1684 420
rect 1774 424 1780 425
rect 1774 420 1775 424
rect 1779 420 1780 424
rect 1774 419 1780 420
rect 1886 424 1892 425
rect 1886 420 1887 424
rect 1891 420 1892 424
rect 1886 419 1892 420
rect 2014 424 2020 425
rect 2014 420 2015 424
rect 2019 420 2020 424
rect 2014 419 2020 420
rect 2158 424 2164 425
rect 2158 420 2159 424
rect 2163 420 2164 424
rect 2158 419 2164 420
rect 2310 424 2316 425
rect 2310 420 2311 424
rect 2315 420 2316 424
rect 2310 419 2316 420
rect 2438 424 2444 425
rect 2438 420 2439 424
rect 2443 420 2444 424
rect 2438 419 2444 420
rect 2502 421 2508 422
rect 1326 416 1332 417
rect 2502 417 2503 421
rect 2507 417 2508 421
rect 2502 416 2508 417
rect 1326 404 1332 405
rect 2502 404 2508 405
rect 1326 400 1327 404
rect 1331 400 1332 404
rect 1326 399 1332 400
rect 1366 403 1372 404
rect 1366 399 1367 403
rect 1371 399 1372 403
rect 1366 398 1372 399
rect 1438 403 1444 404
rect 1438 399 1439 403
rect 1443 399 1444 403
rect 1438 398 1444 399
rect 1526 403 1532 404
rect 1526 399 1527 403
rect 1531 399 1532 403
rect 1526 398 1532 399
rect 1614 403 1620 404
rect 1614 399 1615 403
rect 1619 399 1620 403
rect 1614 398 1620 399
rect 1694 403 1700 404
rect 1694 399 1695 403
rect 1699 399 1700 403
rect 1694 398 1700 399
rect 1790 403 1796 404
rect 1790 399 1791 403
rect 1795 399 1796 403
rect 1790 398 1796 399
rect 1902 403 1908 404
rect 1902 399 1903 403
rect 1907 399 1908 403
rect 1902 398 1908 399
rect 2030 403 2036 404
rect 2030 399 2031 403
rect 2035 399 2036 403
rect 2030 398 2036 399
rect 2174 403 2180 404
rect 2174 399 2175 403
rect 2179 399 2180 403
rect 2174 398 2180 399
rect 2326 403 2332 404
rect 2326 399 2327 403
rect 2331 399 2332 403
rect 2326 398 2332 399
rect 2454 403 2460 404
rect 2454 399 2455 403
rect 2459 399 2460 403
rect 2502 400 2503 404
rect 2507 400 2508 404
rect 2502 399 2508 400
rect 2454 398 2460 399
rect 150 365 156 366
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 150 361 151 365
rect 155 361 156 365
rect 150 360 156 361
rect 206 365 212 366
rect 206 361 207 365
rect 211 361 212 365
rect 206 360 212 361
rect 278 365 284 366
rect 278 361 279 365
rect 283 361 284 365
rect 278 360 284 361
rect 358 365 364 366
rect 358 361 359 365
rect 363 361 364 365
rect 358 360 364 361
rect 430 365 436 366
rect 430 361 431 365
rect 435 361 436 365
rect 430 360 436 361
rect 510 365 516 366
rect 510 361 511 365
rect 515 361 516 365
rect 510 360 516 361
rect 590 365 596 366
rect 590 361 591 365
rect 595 361 596 365
rect 590 360 596 361
rect 670 365 676 366
rect 670 361 671 365
rect 675 361 676 365
rect 670 360 676 361
rect 750 365 756 366
rect 750 361 751 365
rect 755 361 756 365
rect 750 360 756 361
rect 822 365 828 366
rect 822 361 823 365
rect 827 361 828 365
rect 822 360 828 361
rect 894 365 900 366
rect 894 361 895 365
rect 899 361 900 365
rect 894 360 900 361
rect 966 365 972 366
rect 966 361 967 365
rect 971 361 972 365
rect 966 360 972 361
rect 1038 365 1044 366
rect 1038 361 1039 365
rect 1043 361 1044 365
rect 1038 360 1044 361
rect 1110 365 1116 366
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 1182 365 1188 366
rect 1182 361 1183 365
rect 1187 361 1188 365
rect 1182 360 1188 361
rect 1238 365 1244 366
rect 1238 361 1239 365
rect 1243 361 1244 365
rect 1238 360 1244 361
rect 1286 364 1292 365
rect 1286 360 1287 364
rect 1291 360 1292 364
rect 110 359 116 360
rect 1286 359 1292 360
rect 1678 349 1684 350
rect 1326 348 1332 349
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 1286 347 1292 348
rect 110 342 116 343
rect 134 344 140 345
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 190 344 196 345
rect 190 340 191 344
rect 195 340 196 344
rect 190 339 196 340
rect 262 344 268 345
rect 262 340 263 344
rect 267 340 268 344
rect 262 339 268 340
rect 342 344 348 345
rect 342 340 343 344
rect 347 340 348 344
rect 342 339 348 340
rect 414 344 420 345
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 806 344 812 345
rect 806 340 807 344
rect 811 340 812 344
rect 806 339 812 340
rect 878 344 884 345
rect 878 340 879 344
rect 883 340 884 344
rect 878 339 884 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1022 344 1028 345
rect 1022 340 1023 344
rect 1027 340 1028 344
rect 1022 339 1028 340
rect 1094 344 1100 345
rect 1094 340 1095 344
rect 1099 340 1100 344
rect 1094 339 1100 340
rect 1166 344 1172 345
rect 1166 340 1167 344
rect 1171 340 1172 344
rect 1166 339 1172 340
rect 1222 344 1228 345
rect 1222 340 1223 344
rect 1227 340 1228 344
rect 1286 343 1287 347
rect 1291 343 1292 347
rect 1326 344 1327 348
rect 1331 344 1332 348
rect 1678 345 1679 349
rect 1683 345 1684 349
rect 1678 344 1684 345
rect 1734 349 1740 350
rect 1734 345 1735 349
rect 1739 345 1740 349
rect 1734 344 1740 345
rect 1806 349 1812 350
rect 1806 345 1807 349
rect 1811 345 1812 349
rect 1806 344 1812 345
rect 1902 349 1908 350
rect 1902 345 1903 349
rect 1907 345 1908 349
rect 1902 344 1908 345
rect 2022 349 2028 350
rect 2022 345 2023 349
rect 2027 345 2028 349
rect 2022 344 2028 345
rect 2158 349 2164 350
rect 2158 345 2159 349
rect 2163 345 2164 349
rect 2158 344 2164 345
rect 2302 349 2308 350
rect 2302 345 2303 349
rect 2307 345 2308 349
rect 2302 344 2308 345
rect 2454 349 2460 350
rect 2454 345 2455 349
rect 2459 345 2460 349
rect 2454 344 2460 345
rect 2502 348 2508 349
rect 2502 344 2503 348
rect 2507 344 2508 348
rect 1326 343 1332 344
rect 2502 343 2508 344
rect 1286 342 1292 343
rect 1222 339 1228 340
rect 1326 331 1332 332
rect 1326 327 1327 331
rect 1331 327 1332 331
rect 2502 331 2508 332
rect 1326 326 1332 327
rect 1662 328 1668 329
rect 134 324 140 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 134 320 135 324
rect 139 320 140 324
rect 134 319 140 320
rect 198 324 204 325
rect 198 320 199 324
rect 203 320 204 324
rect 198 319 204 320
rect 286 324 292 325
rect 286 320 287 324
rect 291 320 292 324
rect 286 319 292 320
rect 374 324 380 325
rect 374 320 375 324
rect 379 320 380 324
rect 374 319 380 320
rect 454 324 460 325
rect 454 320 455 324
rect 459 320 460 324
rect 454 319 460 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 630 324 636 325
rect 630 320 631 324
rect 635 320 636 324
rect 630 319 636 320
rect 726 324 732 325
rect 726 320 727 324
rect 731 320 732 324
rect 726 319 732 320
rect 822 324 828 325
rect 822 320 823 324
rect 827 320 828 324
rect 822 319 828 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 1030 324 1036 325
rect 1030 320 1031 324
rect 1035 320 1036 324
rect 1030 319 1036 320
rect 1134 324 1140 325
rect 1134 320 1135 324
rect 1139 320 1140 324
rect 1134 319 1140 320
rect 1222 324 1228 325
rect 1222 320 1223 324
rect 1227 320 1228 324
rect 1662 324 1663 328
rect 1667 324 1668 328
rect 1662 323 1668 324
rect 1718 328 1724 329
rect 1718 324 1719 328
rect 1723 324 1724 328
rect 1718 323 1724 324
rect 1790 328 1796 329
rect 1790 324 1791 328
rect 1795 324 1796 328
rect 1790 323 1796 324
rect 1886 328 1892 329
rect 1886 324 1887 328
rect 1891 324 1892 328
rect 1886 323 1892 324
rect 2006 328 2012 329
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 2142 328 2148 329
rect 2142 324 2143 328
rect 2147 324 2148 328
rect 2142 323 2148 324
rect 2286 328 2292 329
rect 2286 324 2287 328
rect 2291 324 2292 328
rect 2286 323 2292 324
rect 2438 328 2444 329
rect 2438 324 2439 328
rect 2443 324 2444 328
rect 2502 327 2503 331
rect 2507 327 2508 331
rect 2502 326 2508 327
rect 2438 323 2444 324
rect 1222 319 1228 320
rect 1286 321 1292 322
rect 110 316 116 317
rect 1286 317 1287 321
rect 1291 317 1292 321
rect 1286 316 1292 317
rect 1350 316 1356 317
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1350 312 1351 316
rect 1355 312 1356 316
rect 1350 311 1356 312
rect 1430 316 1436 317
rect 1430 312 1431 316
rect 1435 312 1436 316
rect 1430 311 1436 312
rect 1526 316 1532 317
rect 1526 312 1527 316
rect 1531 312 1532 316
rect 1526 311 1532 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1710 316 1716 317
rect 1710 312 1711 316
rect 1715 312 1716 316
rect 1710 311 1716 312
rect 1806 316 1812 317
rect 1806 312 1807 316
rect 1811 312 1812 316
rect 1806 311 1812 312
rect 1910 316 1916 317
rect 1910 312 1911 316
rect 1915 312 1916 316
rect 1910 311 1916 312
rect 2022 316 2028 317
rect 2022 312 2023 316
rect 2027 312 2028 316
rect 2022 311 2028 312
rect 2150 316 2156 317
rect 2150 312 2151 316
rect 2155 312 2156 316
rect 2150 311 2156 312
rect 2286 316 2292 317
rect 2286 312 2287 316
rect 2291 312 2292 316
rect 2286 311 2292 312
rect 2422 316 2428 317
rect 2422 312 2423 316
rect 2427 312 2428 316
rect 2422 311 2428 312
rect 2502 313 2508 314
rect 1326 308 1332 309
rect 2502 309 2503 313
rect 2507 309 2508 313
rect 2502 308 2508 309
rect 110 304 116 305
rect 1286 304 1292 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 150 303 156 304
rect 150 299 151 303
rect 155 299 156 303
rect 150 298 156 299
rect 214 303 220 304
rect 214 299 215 303
rect 219 299 220 303
rect 214 298 220 299
rect 302 303 308 304
rect 302 299 303 303
rect 307 299 308 303
rect 302 298 308 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 470 303 476 304
rect 470 299 471 303
rect 475 299 476 303
rect 470 298 476 299
rect 558 303 564 304
rect 558 299 559 303
rect 563 299 564 303
rect 558 298 564 299
rect 646 303 652 304
rect 646 299 647 303
rect 651 299 652 303
rect 646 298 652 299
rect 742 303 748 304
rect 742 299 743 303
rect 747 299 748 303
rect 742 298 748 299
rect 838 303 844 304
rect 838 299 839 303
rect 843 299 844 303
rect 838 298 844 299
rect 942 303 948 304
rect 942 299 943 303
rect 947 299 948 303
rect 942 298 948 299
rect 1046 303 1052 304
rect 1046 299 1047 303
rect 1051 299 1052 303
rect 1046 298 1052 299
rect 1150 303 1156 304
rect 1150 299 1151 303
rect 1155 299 1156 303
rect 1150 298 1156 299
rect 1238 303 1244 304
rect 1238 299 1239 303
rect 1243 299 1244 303
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1238 298 1244 299
rect 1326 296 1332 297
rect 2502 296 2508 297
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1326 291 1332 292
rect 1366 295 1372 296
rect 1366 291 1367 295
rect 1371 291 1372 295
rect 1366 290 1372 291
rect 1446 295 1452 296
rect 1446 291 1447 295
rect 1451 291 1452 295
rect 1446 290 1452 291
rect 1542 295 1548 296
rect 1542 291 1543 295
rect 1547 291 1548 295
rect 1542 290 1548 291
rect 1638 295 1644 296
rect 1638 291 1639 295
rect 1643 291 1644 295
rect 1638 290 1644 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1822 295 1828 296
rect 1822 291 1823 295
rect 1827 291 1828 295
rect 1822 290 1828 291
rect 1926 295 1932 296
rect 1926 291 1927 295
rect 1931 291 1932 295
rect 1926 290 1932 291
rect 2038 295 2044 296
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2166 295 2172 296
rect 2166 291 2167 295
rect 2171 291 2172 295
rect 2166 290 2172 291
rect 2302 295 2308 296
rect 2302 291 2303 295
rect 2307 291 2308 295
rect 2302 290 2308 291
rect 2438 295 2444 296
rect 2438 291 2439 295
rect 2443 291 2444 295
rect 2502 292 2503 296
rect 2507 292 2508 296
rect 2502 291 2508 292
rect 2438 290 2444 291
rect 150 245 156 246
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 150 241 151 245
rect 155 241 156 245
rect 150 240 156 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 326 245 332 246
rect 326 241 327 245
rect 331 241 332 245
rect 326 240 332 241
rect 422 245 428 246
rect 422 241 423 245
rect 427 241 428 245
rect 422 240 428 241
rect 518 245 524 246
rect 518 241 519 245
rect 523 241 524 245
rect 518 240 524 241
rect 614 245 620 246
rect 614 241 615 245
rect 619 241 620 245
rect 614 240 620 241
rect 710 245 716 246
rect 710 241 711 245
rect 715 241 716 245
rect 710 240 716 241
rect 806 245 812 246
rect 806 241 807 245
rect 811 241 812 245
rect 806 240 812 241
rect 902 245 908 246
rect 902 241 903 245
rect 907 241 908 245
rect 902 240 908 241
rect 1006 245 1012 246
rect 1006 241 1007 245
rect 1011 241 1012 245
rect 1006 240 1012 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1214 245 1220 246
rect 1214 241 1215 245
rect 1219 241 1220 245
rect 1214 240 1220 241
rect 1286 244 1292 245
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1366 241 1372 242
rect 110 239 116 240
rect 1286 239 1292 240
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1438 241 1444 242
rect 1438 237 1439 241
rect 1443 237 1444 241
rect 1438 236 1444 237
rect 1534 241 1540 242
rect 1534 237 1535 241
rect 1539 237 1540 241
rect 1534 236 1540 237
rect 1630 241 1636 242
rect 1630 237 1631 241
rect 1635 237 1636 241
rect 1630 236 1636 237
rect 1726 241 1732 242
rect 1726 237 1727 241
rect 1731 237 1732 241
rect 1726 236 1732 237
rect 1814 241 1820 242
rect 1814 237 1815 241
rect 1819 237 1820 241
rect 1814 236 1820 237
rect 1902 241 1908 242
rect 1902 237 1903 241
rect 1907 237 1908 241
rect 1902 236 1908 237
rect 1998 241 2004 242
rect 1998 237 1999 241
rect 2003 237 2004 241
rect 1998 236 2004 237
rect 2102 241 2108 242
rect 2102 237 2103 241
rect 2107 237 2108 241
rect 2102 236 2108 237
rect 2214 241 2220 242
rect 2214 237 2215 241
rect 2219 237 2220 241
rect 2214 236 2220 237
rect 2334 241 2340 242
rect 2334 237 2335 241
rect 2339 237 2340 241
rect 2334 236 2340 237
rect 2454 241 2460 242
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2454 236 2460 237
rect 2502 240 2508 241
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 1326 235 1332 236
rect 2502 235 2508 236
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1286 227 1292 228
rect 110 222 116 223
rect 134 224 140 225
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 214 224 220 225
rect 214 220 215 224
rect 219 220 220 224
rect 214 219 220 220
rect 310 224 316 225
rect 310 220 311 224
rect 315 220 316 224
rect 310 219 316 220
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 502 224 508 225
rect 502 220 503 224
rect 507 220 508 224
rect 502 219 508 220
rect 598 224 604 225
rect 598 220 599 224
rect 603 220 604 224
rect 598 219 604 220
rect 694 224 700 225
rect 694 220 695 224
rect 699 220 700 224
rect 694 219 700 220
rect 790 224 796 225
rect 790 220 791 224
rect 795 220 796 224
rect 790 219 796 220
rect 886 224 892 225
rect 886 220 887 224
rect 891 220 892 224
rect 886 219 892 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1094 224 1100 225
rect 1094 220 1095 224
rect 1099 220 1100 224
rect 1094 219 1100 220
rect 1198 224 1204 225
rect 1198 220 1199 224
rect 1203 220 1204 224
rect 1286 223 1287 227
rect 1291 223 1292 227
rect 1286 222 1292 223
rect 1326 223 1332 224
rect 1198 219 1204 220
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1422 220 1428 221
rect 1422 216 1423 220
rect 1427 216 1428 220
rect 1422 215 1428 216
rect 1518 220 1524 221
rect 1518 216 1519 220
rect 1523 216 1524 220
rect 1518 215 1524 216
rect 1614 220 1620 221
rect 1614 216 1615 220
rect 1619 216 1620 220
rect 1614 215 1620 216
rect 1710 220 1716 221
rect 1710 216 1711 220
rect 1715 216 1716 220
rect 1710 215 1716 216
rect 1798 220 1804 221
rect 1798 216 1799 220
rect 1803 216 1804 220
rect 1798 215 1804 216
rect 1886 220 1892 221
rect 1886 216 1887 220
rect 1891 216 1892 220
rect 1886 215 1892 216
rect 1982 220 1988 221
rect 1982 216 1983 220
rect 1987 216 1988 220
rect 1982 215 1988 216
rect 2086 220 2092 221
rect 2086 216 2087 220
rect 2091 216 2092 220
rect 2086 215 2092 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2318 220 2324 221
rect 2318 216 2319 220
rect 2323 216 2324 220
rect 2318 215 2324 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 158 204 164 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 158 200 159 204
rect 163 200 164 204
rect 158 199 164 200
rect 238 204 244 205
rect 238 200 239 204
rect 243 200 244 204
rect 238 199 244 200
rect 326 204 332 205
rect 326 200 327 204
rect 331 200 332 204
rect 326 199 332 200
rect 414 204 420 205
rect 414 200 415 204
rect 419 200 420 204
rect 414 199 420 200
rect 510 204 516 205
rect 510 200 511 204
rect 515 200 516 204
rect 510 199 516 200
rect 606 204 612 205
rect 606 200 607 204
rect 611 200 612 204
rect 606 199 612 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 782 204 788 205
rect 782 200 783 204
rect 787 200 788 204
rect 782 199 788 200
rect 870 204 876 205
rect 870 200 871 204
rect 875 200 876 204
rect 870 199 876 200
rect 958 204 964 205
rect 958 200 959 204
rect 963 200 964 204
rect 958 199 964 200
rect 1046 204 1052 205
rect 1046 200 1047 204
rect 1051 200 1052 204
rect 1046 199 1052 200
rect 1134 204 1140 205
rect 1134 200 1135 204
rect 1139 200 1140 204
rect 1390 204 1396 205
rect 1134 199 1140 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1390 200 1391 204
rect 1395 200 1396 204
rect 1390 199 1396 200
rect 1494 204 1500 205
rect 1494 200 1495 204
rect 1499 200 1500 204
rect 1494 199 1500 200
rect 1598 204 1604 205
rect 1598 200 1599 204
rect 1603 200 1604 204
rect 1598 199 1604 200
rect 1710 204 1716 205
rect 1710 200 1711 204
rect 1715 200 1716 204
rect 1710 199 1716 200
rect 1814 204 1820 205
rect 1814 200 1815 204
rect 1819 200 1820 204
rect 1814 199 1820 200
rect 1918 204 1924 205
rect 1918 200 1919 204
rect 1923 200 1924 204
rect 1918 199 1924 200
rect 2014 204 2020 205
rect 2014 200 2015 204
rect 2019 200 2020 204
rect 2014 199 2020 200
rect 2110 204 2116 205
rect 2110 200 2111 204
rect 2115 200 2116 204
rect 2110 199 2116 200
rect 2198 204 2204 205
rect 2198 200 2199 204
rect 2203 200 2204 204
rect 2198 199 2204 200
rect 2286 204 2292 205
rect 2286 200 2287 204
rect 2291 200 2292 204
rect 2286 199 2292 200
rect 2374 204 2380 205
rect 2374 200 2375 204
rect 2379 200 2380 204
rect 2374 199 2380 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 174 183 180 184
rect 174 179 175 183
rect 179 179 180 183
rect 174 178 180 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 179 260 183
rect 254 178 260 179
rect 342 183 348 184
rect 342 179 343 183
rect 347 179 348 183
rect 342 178 348 179
rect 430 183 436 184
rect 430 179 431 183
rect 435 179 436 183
rect 430 178 436 179
rect 526 183 532 184
rect 526 179 527 183
rect 531 179 532 183
rect 526 178 532 179
rect 622 183 628 184
rect 622 179 623 183
rect 627 179 628 183
rect 622 178 628 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 798 183 804 184
rect 798 179 799 183
rect 803 179 804 183
rect 798 178 804 179
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 974 183 980 184
rect 974 179 975 183
rect 979 179 980 183
rect 974 178 980 179
rect 1062 183 1068 184
rect 1062 179 1063 183
rect 1067 179 1068 183
rect 1062 178 1068 179
rect 1150 183 1156 184
rect 1150 179 1151 183
rect 1155 179 1156 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1406 183 1412 184
rect 1406 179 1407 183
rect 1411 179 1412 183
rect 1150 178 1156 179
rect 1406 178 1412 179
rect 1510 183 1516 184
rect 1510 179 1511 183
rect 1515 179 1516 183
rect 1510 178 1516 179
rect 1614 183 1620 184
rect 1614 179 1615 183
rect 1619 179 1620 183
rect 1614 178 1620 179
rect 1726 183 1732 184
rect 1726 179 1727 183
rect 1731 179 1732 183
rect 1726 178 1732 179
rect 1830 183 1836 184
rect 1830 179 1831 183
rect 1835 179 1836 183
rect 1830 178 1836 179
rect 1934 183 1940 184
rect 1934 179 1935 183
rect 1939 179 1940 183
rect 1934 178 1940 179
rect 2030 183 2036 184
rect 2030 179 2031 183
rect 2035 179 2036 183
rect 2030 178 2036 179
rect 2126 183 2132 184
rect 2126 179 2127 183
rect 2131 179 2132 183
rect 2126 178 2132 179
rect 2214 183 2220 184
rect 2214 179 2215 183
rect 2219 179 2220 183
rect 2214 178 2220 179
rect 2302 183 2308 184
rect 2302 179 2303 183
rect 2307 179 2308 183
rect 2302 178 2308 179
rect 2390 183 2396 184
rect 2390 179 2391 183
rect 2395 179 2396 183
rect 2390 178 2396 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2454 178 2460 179
rect 150 113 156 114
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 150 109 151 113
rect 155 109 156 113
rect 150 108 156 109
rect 206 113 212 114
rect 206 109 207 113
rect 211 109 212 113
rect 206 108 212 109
rect 262 113 268 114
rect 262 109 263 113
rect 267 109 268 113
rect 262 108 268 109
rect 318 113 324 114
rect 318 109 319 113
rect 323 109 324 113
rect 318 108 324 109
rect 374 113 380 114
rect 374 109 375 113
rect 379 109 380 113
rect 374 108 380 109
rect 430 113 436 114
rect 430 109 431 113
rect 435 109 436 113
rect 430 108 436 109
rect 486 113 492 114
rect 486 109 487 113
rect 491 109 492 113
rect 486 108 492 109
rect 550 113 556 114
rect 550 109 551 113
rect 555 109 556 113
rect 550 108 556 109
rect 622 113 628 114
rect 622 109 623 113
rect 627 109 628 113
rect 622 108 628 109
rect 686 113 692 114
rect 686 109 687 113
rect 691 109 692 113
rect 686 108 692 109
rect 750 113 756 114
rect 750 109 751 113
rect 755 109 756 113
rect 750 108 756 109
rect 814 113 820 114
rect 814 109 815 113
rect 819 109 820 113
rect 814 108 820 109
rect 878 113 884 114
rect 878 109 879 113
rect 883 109 884 113
rect 878 108 884 109
rect 942 113 948 114
rect 942 109 943 113
rect 947 109 948 113
rect 942 108 948 109
rect 1006 113 1012 114
rect 1006 109 1007 113
rect 1011 109 1012 113
rect 1006 108 1012 109
rect 1070 113 1076 114
rect 1070 109 1071 113
rect 1075 109 1076 113
rect 1070 108 1076 109
rect 1134 113 1140 114
rect 1134 109 1135 113
rect 1139 109 1140 113
rect 1134 108 1140 109
rect 1198 113 1204 114
rect 1366 113 1372 114
rect 1198 109 1199 113
rect 1203 109 1204 113
rect 1198 108 1204 109
rect 1286 112 1292 113
rect 1286 108 1287 112
rect 1291 108 1292 112
rect 110 107 116 108
rect 1286 107 1292 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1814 113 1820 114
rect 1814 109 1815 113
rect 1819 109 1820 113
rect 1814 108 1820 109
rect 1870 113 1876 114
rect 1870 109 1871 113
rect 1875 109 1876 113
rect 1870 108 1876 109
rect 1926 113 1932 114
rect 1926 109 1927 113
rect 1931 109 1932 113
rect 1926 108 1932 109
rect 1982 113 1988 114
rect 1982 109 1983 113
rect 1987 109 1988 113
rect 1982 108 1988 109
rect 2038 113 2044 114
rect 2038 109 2039 113
rect 2043 109 2044 113
rect 2038 108 2044 109
rect 2094 113 2100 114
rect 2094 109 2095 113
rect 2099 109 2100 113
rect 2094 108 2100 109
rect 2158 113 2164 114
rect 2158 109 2159 113
rect 2163 109 2164 113
rect 2158 108 2164 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2286 113 2292 114
rect 2286 109 2287 113
rect 2291 109 2292 113
rect 2286 108 2292 109
rect 2342 113 2348 114
rect 2342 109 2343 113
rect 2347 109 2348 113
rect 2342 108 2348 109
rect 2398 113 2404 114
rect 2398 109 2399 113
rect 2403 109 2404 113
rect 2398 108 2404 109
rect 2454 113 2460 114
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 1326 107 1332 108
rect 2502 107 2508 108
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1286 95 1292 96
rect 110 90 116 91
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 246 92 252 93
rect 246 88 247 92
rect 251 88 252 92
rect 246 87 252 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 358 92 364 93
rect 358 88 359 92
rect 363 88 364 92
rect 358 87 364 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 606 92 612 93
rect 606 88 607 92
rect 611 88 612 92
rect 606 87 612 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 798 92 804 93
rect 798 88 799 92
rect 803 88 804 92
rect 798 87 804 88
rect 862 92 868 93
rect 862 88 863 92
rect 867 88 868 92
rect 862 87 868 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1054 92 1060 93
rect 1054 88 1055 92
rect 1059 88 1060 92
rect 1054 87 1060 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1182 92 1188 93
rect 1182 88 1183 92
rect 1187 88 1188 92
rect 1286 91 1287 95
rect 1291 91 1292 95
rect 1286 90 1292 91
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1182 87 1188 88
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1798 92 1804 93
rect 1798 88 1799 92
rect 1803 88 1804 92
rect 1798 87 1804 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1910 92 1916 93
rect 1910 88 1911 92
rect 1915 88 1916 92
rect 1910 87 1916 88
rect 1966 92 1972 93
rect 1966 88 1967 92
rect 1971 88 1972 92
rect 1966 87 1972 88
rect 2022 92 2028 93
rect 2022 88 2023 92
rect 2027 88 2028 92
rect 2022 87 2028 88
rect 2078 92 2084 93
rect 2078 88 2079 92
rect 2083 88 2084 92
rect 2078 87 2084 88
rect 2142 92 2148 93
rect 2142 88 2143 92
rect 2147 88 2148 92
rect 2142 87 2148 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2270 92 2276 93
rect 2270 88 2271 92
rect 2275 88 2276 92
rect 2270 87 2276 88
rect 2326 92 2332 93
rect 2326 88 2327 92
rect 2331 88 2332 92
rect 2326 87 2332 88
rect 2382 92 2388 93
rect 2382 88 2383 92
rect 2387 88 2388 92
rect 2382 87 2388 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
<< m3c >>
rect 111 2552 115 2556
rect 719 2553 723 2557
rect 775 2553 779 2557
rect 831 2553 835 2557
rect 887 2553 891 2557
rect 943 2553 947 2557
rect 1287 2552 1291 2556
rect 111 2535 115 2539
rect 703 2532 707 2536
rect 759 2532 763 2536
rect 815 2532 819 2536
rect 871 2532 875 2536
rect 927 2532 931 2536
rect 1287 2535 1291 2539
rect 1327 2528 1331 2532
rect 1399 2529 1403 2533
rect 1455 2529 1459 2533
rect 1511 2529 1515 2533
rect 1567 2529 1571 2533
rect 1623 2529 1627 2533
rect 1679 2529 1683 2533
rect 1735 2529 1739 2533
rect 1791 2529 1795 2533
rect 1847 2529 1851 2533
rect 1903 2529 1907 2533
rect 1959 2529 1963 2533
rect 2015 2529 2019 2533
rect 2071 2529 2075 2533
rect 2127 2529 2131 2533
rect 2183 2529 2187 2533
rect 2503 2528 2507 2532
rect 111 2517 115 2521
rect 167 2520 171 2524
rect 223 2520 227 2524
rect 279 2520 283 2524
rect 343 2520 347 2524
rect 407 2520 411 2524
rect 479 2520 483 2524
rect 559 2520 563 2524
rect 639 2520 643 2524
rect 719 2520 723 2524
rect 799 2520 803 2524
rect 879 2520 883 2524
rect 959 2520 963 2524
rect 1039 2520 1043 2524
rect 1287 2517 1291 2521
rect 1327 2511 1331 2515
rect 1383 2508 1387 2512
rect 1439 2508 1443 2512
rect 1495 2508 1499 2512
rect 1551 2508 1555 2512
rect 1607 2508 1611 2512
rect 1663 2508 1667 2512
rect 1719 2508 1723 2512
rect 1775 2508 1779 2512
rect 1831 2508 1835 2512
rect 1887 2508 1891 2512
rect 1943 2508 1947 2512
rect 1999 2508 2003 2512
rect 2055 2508 2059 2512
rect 2111 2508 2115 2512
rect 2167 2508 2171 2512
rect 2503 2511 2507 2515
rect 111 2500 115 2504
rect 183 2499 187 2503
rect 239 2499 243 2503
rect 295 2499 299 2503
rect 359 2499 363 2503
rect 423 2499 427 2503
rect 495 2499 499 2503
rect 575 2499 579 2503
rect 655 2499 659 2503
rect 735 2499 739 2503
rect 815 2499 819 2503
rect 895 2499 899 2503
rect 975 2499 979 2503
rect 1055 2499 1059 2503
rect 1287 2500 1291 2504
rect 1327 2485 1331 2489
rect 1351 2488 1355 2492
rect 1423 2488 1427 2492
rect 1511 2488 1515 2492
rect 1599 2488 1603 2492
rect 1687 2488 1691 2492
rect 1775 2488 1779 2492
rect 1863 2488 1867 2492
rect 1951 2488 1955 2492
rect 2039 2488 2043 2492
rect 2127 2488 2131 2492
rect 2503 2485 2507 2489
rect 1327 2468 1331 2472
rect 1367 2467 1371 2471
rect 1439 2467 1443 2471
rect 1527 2467 1531 2471
rect 1615 2467 1619 2471
rect 1703 2467 1707 2471
rect 1791 2467 1795 2471
rect 1879 2467 1883 2471
rect 1967 2467 1971 2471
rect 2055 2467 2059 2471
rect 2143 2467 2147 2471
rect 2503 2468 2507 2472
rect 111 2448 115 2452
rect 183 2449 187 2453
rect 247 2449 251 2453
rect 327 2449 331 2453
rect 415 2449 419 2453
rect 503 2449 507 2453
rect 599 2449 603 2453
rect 695 2449 699 2453
rect 791 2449 795 2453
rect 879 2449 883 2453
rect 967 2449 971 2453
rect 1063 2449 1067 2453
rect 1159 2449 1163 2453
rect 1287 2448 1291 2452
rect 111 2431 115 2435
rect 167 2428 171 2432
rect 231 2428 235 2432
rect 311 2428 315 2432
rect 399 2428 403 2432
rect 487 2428 491 2432
rect 583 2428 587 2432
rect 679 2428 683 2432
rect 775 2428 779 2432
rect 863 2428 867 2432
rect 951 2428 955 2432
rect 1047 2428 1051 2432
rect 1143 2428 1147 2432
rect 1287 2431 1291 2435
rect 111 2409 115 2413
rect 151 2412 155 2416
rect 231 2412 235 2416
rect 319 2412 323 2416
rect 415 2412 419 2416
rect 519 2412 523 2416
rect 623 2412 627 2416
rect 727 2412 731 2416
rect 831 2412 835 2416
rect 935 2412 939 2416
rect 1039 2412 1043 2416
rect 1151 2412 1155 2416
rect 1287 2409 1291 2413
rect 1327 2408 1331 2412
rect 1367 2409 1371 2413
rect 1439 2409 1443 2413
rect 1543 2409 1547 2413
rect 1639 2409 1643 2413
rect 1735 2409 1739 2413
rect 1823 2409 1827 2413
rect 1911 2409 1915 2413
rect 2007 2409 2011 2413
rect 2103 2409 2107 2413
rect 2503 2408 2507 2412
rect 111 2392 115 2396
rect 167 2391 171 2395
rect 247 2391 251 2395
rect 335 2391 339 2395
rect 431 2391 435 2395
rect 535 2391 539 2395
rect 639 2391 643 2395
rect 743 2391 747 2395
rect 847 2391 851 2395
rect 951 2391 955 2395
rect 1055 2391 1059 2395
rect 1167 2391 1171 2395
rect 1287 2392 1291 2396
rect 1327 2391 1331 2395
rect 1351 2388 1355 2392
rect 1423 2388 1427 2392
rect 1527 2388 1531 2392
rect 1623 2388 1627 2392
rect 1719 2388 1723 2392
rect 1807 2388 1811 2392
rect 1895 2388 1899 2392
rect 1991 2388 1995 2392
rect 2087 2388 2091 2392
rect 2503 2391 2507 2395
rect 1327 2365 1331 2369
rect 1351 2368 1355 2372
rect 1407 2368 1411 2372
rect 1495 2368 1499 2372
rect 1583 2368 1587 2372
rect 1671 2368 1675 2372
rect 1751 2368 1755 2372
rect 1831 2368 1835 2372
rect 1919 2368 1923 2372
rect 2007 2368 2011 2372
rect 2095 2368 2099 2372
rect 2503 2365 2507 2369
rect 1327 2348 1331 2352
rect 1367 2347 1371 2351
rect 1423 2347 1427 2351
rect 1511 2347 1515 2351
rect 1599 2347 1603 2351
rect 1687 2347 1691 2351
rect 1767 2347 1771 2351
rect 1847 2347 1851 2351
rect 1935 2347 1939 2351
rect 2023 2347 2027 2351
rect 2111 2347 2115 2351
rect 2503 2348 2507 2352
rect 111 2340 115 2344
rect 175 2341 179 2345
rect 279 2341 283 2345
rect 391 2341 395 2345
rect 503 2341 507 2345
rect 623 2341 627 2345
rect 743 2341 747 2345
rect 871 2341 875 2345
rect 999 2341 1003 2345
rect 1127 2341 1131 2345
rect 1287 2340 1291 2344
rect 111 2323 115 2327
rect 159 2320 163 2324
rect 263 2320 267 2324
rect 375 2320 379 2324
rect 487 2320 491 2324
rect 607 2320 611 2324
rect 727 2320 731 2324
rect 855 2320 859 2324
rect 983 2320 987 2324
rect 1111 2320 1115 2324
rect 1287 2323 1291 2327
rect 111 2301 115 2305
rect 207 2304 211 2308
rect 287 2304 291 2308
rect 375 2304 379 2308
rect 471 2304 475 2308
rect 559 2304 563 2308
rect 647 2304 651 2308
rect 735 2304 739 2308
rect 815 2304 819 2308
rect 903 2304 907 2308
rect 991 2304 995 2308
rect 1079 2304 1083 2308
rect 1287 2301 1291 2305
rect 1327 2292 1331 2296
rect 1367 2293 1371 2297
rect 1455 2293 1459 2297
rect 1543 2293 1547 2297
rect 1639 2293 1643 2297
rect 1735 2293 1739 2297
rect 1831 2293 1835 2297
rect 1927 2293 1931 2297
rect 2015 2293 2019 2297
rect 2111 2293 2115 2297
rect 2207 2293 2211 2297
rect 2503 2292 2507 2296
rect 111 2284 115 2288
rect 223 2283 227 2287
rect 303 2283 307 2287
rect 391 2283 395 2287
rect 487 2283 491 2287
rect 575 2283 579 2287
rect 663 2283 667 2287
rect 751 2283 755 2287
rect 831 2283 835 2287
rect 919 2283 923 2287
rect 1007 2283 1011 2287
rect 1095 2283 1099 2287
rect 1287 2284 1291 2288
rect 1327 2275 1331 2279
rect 1351 2272 1355 2276
rect 1439 2272 1443 2276
rect 1527 2272 1531 2276
rect 1623 2272 1627 2276
rect 1719 2272 1723 2276
rect 1815 2272 1819 2276
rect 1911 2272 1915 2276
rect 1999 2272 2003 2276
rect 2095 2272 2099 2276
rect 2191 2272 2195 2276
rect 2503 2275 2507 2279
rect 1327 2257 1331 2261
rect 1455 2260 1459 2264
rect 1543 2260 1547 2264
rect 1639 2260 1643 2264
rect 1735 2260 1739 2264
rect 1839 2260 1843 2264
rect 1935 2260 1939 2264
rect 2031 2260 2035 2264
rect 2119 2260 2123 2264
rect 2215 2260 2219 2264
rect 2311 2260 2315 2264
rect 2503 2257 2507 2261
rect 1327 2240 1331 2244
rect 1471 2239 1475 2243
rect 1559 2239 1563 2243
rect 1655 2239 1659 2243
rect 1751 2239 1755 2243
rect 1855 2239 1859 2243
rect 1951 2239 1955 2243
rect 2047 2239 2051 2243
rect 2135 2239 2139 2243
rect 2231 2239 2235 2243
rect 2327 2239 2331 2243
rect 2503 2240 2507 2244
rect 111 2228 115 2232
rect 263 2229 267 2233
rect 319 2229 323 2233
rect 383 2229 387 2233
rect 447 2229 451 2233
rect 503 2229 507 2233
rect 559 2229 563 2233
rect 615 2229 619 2233
rect 671 2229 675 2233
rect 727 2229 731 2233
rect 791 2229 795 2233
rect 855 2229 859 2233
rect 919 2229 923 2233
rect 983 2229 987 2233
rect 1047 2229 1051 2233
rect 1111 2229 1115 2233
rect 1287 2228 1291 2232
rect 111 2211 115 2215
rect 247 2208 251 2212
rect 303 2208 307 2212
rect 367 2208 371 2212
rect 431 2208 435 2212
rect 487 2208 491 2212
rect 543 2208 547 2212
rect 599 2208 603 2212
rect 655 2208 659 2212
rect 711 2208 715 2212
rect 775 2208 779 2212
rect 839 2208 843 2212
rect 903 2208 907 2212
rect 967 2208 971 2212
rect 1031 2208 1035 2212
rect 1095 2208 1099 2212
rect 1287 2211 1291 2215
rect 111 2189 115 2193
rect 335 2192 339 2196
rect 391 2192 395 2196
rect 447 2192 451 2196
rect 503 2192 507 2196
rect 559 2192 563 2196
rect 1287 2189 1291 2193
rect 1327 2184 1331 2188
rect 1567 2185 1571 2189
rect 1623 2185 1627 2189
rect 1679 2185 1683 2189
rect 1743 2185 1747 2189
rect 1807 2185 1811 2189
rect 1871 2185 1875 2189
rect 1927 2185 1931 2189
rect 1983 2185 1987 2189
rect 2039 2185 2043 2189
rect 2095 2185 2099 2189
rect 2159 2185 2163 2189
rect 2223 2185 2227 2189
rect 2287 2185 2291 2189
rect 2343 2185 2347 2189
rect 2399 2185 2403 2189
rect 2455 2185 2459 2189
rect 2503 2184 2507 2188
rect 111 2172 115 2176
rect 351 2171 355 2175
rect 407 2171 411 2175
rect 463 2171 467 2175
rect 519 2171 523 2175
rect 575 2171 579 2175
rect 1287 2172 1291 2176
rect 1327 2167 1331 2171
rect 1551 2164 1555 2168
rect 1607 2164 1611 2168
rect 1663 2164 1667 2168
rect 1727 2164 1731 2168
rect 1791 2164 1795 2168
rect 1855 2164 1859 2168
rect 1911 2164 1915 2168
rect 1967 2164 1971 2168
rect 2023 2164 2027 2168
rect 2079 2164 2083 2168
rect 2143 2164 2147 2168
rect 2207 2164 2211 2168
rect 2271 2164 2275 2168
rect 2327 2164 2331 2168
rect 2383 2164 2387 2168
rect 2439 2164 2443 2168
rect 2503 2167 2507 2171
rect 1327 2137 1331 2141
rect 1663 2140 1667 2144
rect 1719 2140 1723 2144
rect 1791 2140 1795 2144
rect 1871 2140 1875 2144
rect 1967 2140 1971 2144
rect 2079 2140 2083 2144
rect 2199 2140 2203 2144
rect 2327 2140 2331 2144
rect 2439 2140 2443 2144
rect 2503 2137 2507 2141
rect 111 2120 115 2124
rect 415 2121 419 2125
rect 511 2121 515 2125
rect 607 2121 611 2125
rect 711 2121 715 2125
rect 815 2121 819 2125
rect 927 2121 931 2125
rect 1039 2121 1043 2125
rect 1151 2121 1155 2125
rect 1239 2121 1243 2125
rect 1287 2120 1291 2124
rect 1327 2120 1331 2124
rect 1679 2119 1683 2123
rect 1735 2119 1739 2123
rect 1807 2119 1811 2123
rect 1887 2119 1891 2123
rect 1983 2119 1987 2123
rect 2095 2119 2099 2123
rect 2215 2119 2219 2123
rect 2343 2119 2347 2123
rect 2455 2119 2459 2123
rect 2503 2120 2507 2124
rect 111 2103 115 2107
rect 399 2100 403 2104
rect 495 2100 499 2104
rect 591 2100 595 2104
rect 695 2100 699 2104
rect 799 2100 803 2104
rect 911 2100 915 2104
rect 1023 2100 1027 2104
rect 1135 2100 1139 2104
rect 1223 2100 1227 2104
rect 1287 2103 1291 2107
rect 111 2085 115 2089
rect 375 2088 379 2092
rect 447 2088 451 2092
rect 519 2088 523 2092
rect 599 2088 603 2092
rect 679 2088 683 2092
rect 759 2088 763 2092
rect 831 2088 835 2092
rect 903 2088 907 2092
rect 967 2088 971 2092
rect 1031 2088 1035 2092
rect 1103 2088 1107 2092
rect 1167 2088 1171 2092
rect 1223 2088 1227 2092
rect 1287 2085 1291 2089
rect 111 2068 115 2072
rect 391 2067 395 2071
rect 463 2067 467 2071
rect 535 2067 539 2071
rect 615 2067 619 2071
rect 695 2067 699 2071
rect 775 2067 779 2071
rect 847 2067 851 2071
rect 919 2067 923 2071
rect 983 2067 987 2071
rect 1047 2067 1051 2071
rect 1119 2067 1123 2071
rect 1183 2067 1187 2071
rect 1239 2067 1243 2071
rect 1287 2068 1291 2072
rect 1327 2056 1331 2060
rect 1367 2057 1371 2061
rect 1423 2057 1427 2061
rect 1503 2057 1507 2061
rect 1591 2057 1595 2061
rect 1679 2057 1683 2061
rect 1783 2057 1787 2061
rect 1895 2057 1899 2061
rect 2023 2057 2027 2061
rect 2167 2057 2171 2061
rect 2319 2057 2323 2061
rect 2455 2057 2459 2061
rect 2503 2056 2507 2060
rect 1327 2039 1331 2043
rect 1351 2036 1355 2040
rect 1407 2036 1411 2040
rect 1487 2036 1491 2040
rect 1575 2036 1579 2040
rect 1663 2036 1667 2040
rect 1767 2036 1771 2040
rect 1879 2036 1883 2040
rect 2007 2036 2011 2040
rect 2151 2036 2155 2040
rect 2303 2036 2307 2040
rect 2439 2036 2443 2040
rect 2503 2039 2507 2043
rect 1327 2021 1331 2025
rect 1351 2024 1355 2028
rect 1423 2024 1427 2028
rect 1519 2024 1523 2028
rect 1615 2024 1619 2028
rect 1719 2024 1723 2028
rect 1823 2024 1827 2028
rect 1935 2024 1939 2028
rect 2055 2024 2059 2028
rect 2183 2024 2187 2028
rect 2319 2024 2323 2028
rect 2439 2024 2443 2028
rect 2503 2021 2507 2025
rect 111 2012 115 2016
rect 295 2013 299 2017
rect 375 2013 379 2017
rect 463 2013 467 2017
rect 551 2013 555 2017
rect 639 2013 643 2017
rect 719 2013 723 2017
rect 799 2013 803 2017
rect 887 2013 891 2017
rect 975 2013 979 2017
rect 1063 2013 1067 2017
rect 1287 2012 1291 2016
rect 1327 2004 1331 2008
rect 1367 2003 1371 2007
rect 1439 2003 1443 2007
rect 1535 2003 1539 2007
rect 1631 2003 1635 2007
rect 1735 2003 1739 2007
rect 1839 2003 1843 2007
rect 1951 2003 1955 2007
rect 2071 2003 2075 2007
rect 2199 2003 2203 2007
rect 2335 2003 2339 2007
rect 2455 2003 2459 2007
rect 2503 2004 2507 2008
rect 111 1995 115 1999
rect 279 1992 283 1996
rect 359 1992 363 1996
rect 447 1992 451 1996
rect 535 1992 539 1996
rect 623 1992 627 1996
rect 703 1992 707 1996
rect 783 1992 787 1996
rect 871 1992 875 1996
rect 959 1992 963 1996
rect 1047 1992 1051 1996
rect 1287 1995 1291 1999
rect 111 1973 115 1977
rect 135 1976 139 1980
rect 207 1976 211 1980
rect 287 1976 291 1980
rect 383 1976 387 1980
rect 487 1976 491 1980
rect 591 1976 595 1980
rect 695 1976 699 1980
rect 799 1976 803 1980
rect 903 1976 907 1980
rect 1015 1976 1019 1980
rect 1287 1973 1291 1977
rect 111 1956 115 1960
rect 151 1955 155 1959
rect 223 1955 227 1959
rect 303 1955 307 1959
rect 399 1955 403 1959
rect 503 1955 507 1959
rect 607 1955 611 1959
rect 711 1955 715 1959
rect 815 1955 819 1959
rect 919 1955 923 1959
rect 1031 1955 1035 1959
rect 1287 1956 1291 1960
rect 1327 1948 1331 1952
rect 1455 1949 1459 1953
rect 1543 1949 1547 1953
rect 1639 1949 1643 1953
rect 1735 1949 1739 1953
rect 1839 1949 1843 1953
rect 1943 1949 1947 1953
rect 2047 1949 2051 1953
rect 2151 1949 2155 1953
rect 2255 1949 2259 1953
rect 2367 1949 2371 1953
rect 2455 1949 2459 1953
rect 2503 1948 2507 1952
rect 1327 1931 1331 1935
rect 1439 1928 1443 1932
rect 1527 1928 1531 1932
rect 1623 1928 1627 1932
rect 1719 1928 1723 1932
rect 1823 1928 1827 1932
rect 1927 1928 1931 1932
rect 2031 1928 2035 1932
rect 2135 1928 2139 1932
rect 2239 1928 2243 1932
rect 2351 1928 2355 1932
rect 2439 1928 2443 1932
rect 2503 1931 2507 1935
rect 1327 1909 1331 1913
rect 1527 1912 1531 1916
rect 1615 1912 1619 1916
rect 1711 1912 1715 1916
rect 1815 1912 1819 1916
rect 1919 1912 1923 1916
rect 2015 1912 2019 1916
rect 2111 1912 2115 1916
rect 2199 1912 2203 1916
rect 2287 1912 2291 1916
rect 2375 1912 2379 1916
rect 2439 1912 2443 1916
rect 2503 1909 2507 1913
rect 111 1896 115 1900
rect 151 1897 155 1901
rect 239 1897 243 1901
rect 375 1897 379 1901
rect 527 1897 531 1901
rect 687 1897 691 1901
rect 863 1897 867 1901
rect 1039 1897 1043 1901
rect 1287 1896 1291 1900
rect 1327 1892 1331 1896
rect 1543 1891 1547 1895
rect 1631 1891 1635 1895
rect 1727 1891 1731 1895
rect 1831 1891 1835 1895
rect 1935 1891 1939 1895
rect 2031 1891 2035 1895
rect 2127 1891 2131 1895
rect 2215 1891 2219 1895
rect 2303 1891 2307 1895
rect 2391 1891 2395 1895
rect 2455 1891 2459 1895
rect 2503 1892 2507 1896
rect 111 1879 115 1883
rect 135 1876 139 1880
rect 223 1876 227 1880
rect 359 1876 363 1880
rect 511 1876 515 1880
rect 671 1876 675 1880
rect 847 1876 851 1880
rect 1023 1876 1027 1880
rect 1287 1879 1291 1883
rect 111 1861 115 1865
rect 135 1864 139 1868
rect 191 1864 195 1868
rect 263 1864 267 1868
rect 335 1864 339 1868
rect 407 1864 411 1868
rect 479 1864 483 1868
rect 551 1864 555 1868
rect 615 1864 619 1868
rect 679 1864 683 1868
rect 743 1864 747 1868
rect 815 1864 819 1868
rect 887 1864 891 1868
rect 959 1864 963 1868
rect 1039 1864 1043 1868
rect 1287 1861 1291 1865
rect 111 1844 115 1848
rect 151 1843 155 1847
rect 207 1843 211 1847
rect 279 1843 283 1847
rect 351 1843 355 1847
rect 423 1843 427 1847
rect 495 1843 499 1847
rect 567 1843 571 1847
rect 631 1843 635 1847
rect 695 1843 699 1847
rect 759 1843 763 1847
rect 831 1843 835 1847
rect 903 1843 907 1847
rect 975 1843 979 1847
rect 1055 1843 1059 1847
rect 1287 1844 1291 1848
rect 1327 1840 1331 1844
rect 1535 1841 1539 1845
rect 1607 1841 1611 1845
rect 1687 1841 1691 1845
rect 1783 1841 1787 1845
rect 1879 1841 1883 1845
rect 1983 1841 1987 1845
rect 2079 1841 2083 1845
rect 2175 1841 2179 1845
rect 2271 1841 2275 1845
rect 2367 1841 2371 1845
rect 2455 1841 2459 1845
rect 2503 1840 2507 1844
rect 1327 1823 1331 1827
rect 1519 1820 1523 1824
rect 1591 1820 1595 1824
rect 1671 1820 1675 1824
rect 1767 1820 1771 1824
rect 1863 1820 1867 1824
rect 1967 1820 1971 1824
rect 2063 1820 2067 1824
rect 2159 1820 2163 1824
rect 2255 1820 2259 1824
rect 2351 1820 2355 1824
rect 2439 1820 2443 1824
rect 2503 1823 2507 1827
rect 1327 1801 1331 1805
rect 1463 1804 1467 1808
rect 1559 1804 1563 1808
rect 1663 1804 1667 1808
rect 1767 1804 1771 1808
rect 1879 1804 1883 1808
rect 1983 1804 1987 1808
rect 2087 1804 2091 1808
rect 2183 1804 2187 1808
rect 2271 1804 2275 1808
rect 2367 1804 2371 1808
rect 2439 1804 2443 1808
rect 2503 1801 2507 1805
rect 111 1784 115 1788
rect 151 1785 155 1789
rect 231 1785 235 1789
rect 335 1785 339 1789
rect 439 1785 443 1789
rect 535 1785 539 1789
rect 631 1785 635 1789
rect 719 1785 723 1789
rect 799 1785 803 1789
rect 879 1785 883 1789
rect 959 1785 963 1789
rect 1039 1785 1043 1789
rect 1119 1785 1123 1789
rect 1287 1784 1291 1788
rect 1327 1784 1331 1788
rect 1479 1783 1483 1787
rect 1575 1783 1579 1787
rect 1679 1783 1683 1787
rect 1783 1783 1787 1787
rect 1895 1783 1899 1787
rect 1999 1783 2003 1787
rect 2103 1783 2107 1787
rect 2199 1783 2203 1787
rect 2287 1783 2291 1787
rect 2383 1783 2387 1787
rect 2455 1783 2459 1787
rect 2503 1784 2507 1788
rect 111 1767 115 1771
rect 135 1764 139 1768
rect 215 1764 219 1768
rect 319 1764 323 1768
rect 423 1764 427 1768
rect 519 1764 523 1768
rect 615 1764 619 1768
rect 703 1764 707 1768
rect 783 1764 787 1768
rect 863 1764 867 1768
rect 943 1764 947 1768
rect 1023 1764 1027 1768
rect 1103 1764 1107 1768
rect 1287 1767 1291 1771
rect 111 1745 115 1749
rect 135 1748 139 1752
rect 239 1748 243 1752
rect 351 1748 355 1752
rect 463 1748 467 1752
rect 575 1748 579 1752
rect 679 1748 683 1752
rect 783 1748 787 1752
rect 887 1748 891 1752
rect 991 1748 995 1752
rect 1103 1748 1107 1752
rect 1287 1745 1291 1749
rect 111 1728 115 1732
rect 151 1727 155 1731
rect 255 1727 259 1731
rect 367 1727 371 1731
rect 479 1727 483 1731
rect 591 1727 595 1731
rect 695 1727 699 1731
rect 799 1727 803 1731
rect 903 1727 907 1731
rect 1007 1727 1011 1731
rect 1119 1727 1123 1731
rect 1287 1728 1291 1732
rect 1327 1728 1331 1732
rect 1375 1729 1379 1733
rect 1471 1729 1475 1733
rect 1567 1729 1571 1733
rect 1671 1729 1675 1733
rect 1775 1729 1779 1733
rect 1887 1729 1891 1733
rect 1999 1729 2003 1733
rect 2111 1729 2115 1733
rect 2231 1729 2235 1733
rect 2351 1729 2355 1733
rect 2455 1729 2459 1733
rect 2503 1728 2507 1732
rect 1327 1711 1331 1715
rect 1359 1708 1363 1712
rect 1455 1708 1459 1712
rect 1551 1708 1555 1712
rect 1655 1708 1659 1712
rect 1759 1708 1763 1712
rect 1871 1708 1875 1712
rect 1983 1708 1987 1712
rect 2095 1708 2099 1712
rect 2215 1708 2219 1712
rect 2335 1708 2339 1712
rect 2439 1708 2443 1712
rect 2503 1711 2507 1715
rect 1327 1693 1331 1697
rect 1351 1696 1355 1700
rect 1431 1696 1435 1700
rect 1535 1696 1539 1700
rect 1647 1696 1651 1700
rect 1759 1696 1763 1700
rect 1879 1696 1883 1700
rect 2015 1696 2019 1700
rect 2159 1696 2163 1700
rect 2311 1696 2315 1700
rect 2439 1696 2443 1700
rect 2503 1693 2507 1697
rect 111 1672 115 1676
rect 191 1673 195 1677
rect 271 1673 275 1677
rect 351 1673 355 1677
rect 439 1673 443 1677
rect 535 1673 539 1677
rect 639 1673 643 1677
rect 743 1673 747 1677
rect 847 1673 851 1677
rect 951 1673 955 1677
rect 1063 1673 1067 1677
rect 1175 1673 1179 1677
rect 1287 1672 1291 1676
rect 1327 1676 1331 1680
rect 1367 1675 1371 1679
rect 1447 1675 1451 1679
rect 1551 1675 1555 1679
rect 1663 1675 1667 1679
rect 1775 1675 1779 1679
rect 1895 1675 1899 1679
rect 2031 1675 2035 1679
rect 2175 1675 2179 1679
rect 2327 1675 2331 1679
rect 2455 1675 2459 1679
rect 2503 1676 2507 1680
rect 111 1655 115 1659
rect 175 1652 179 1656
rect 255 1652 259 1656
rect 335 1652 339 1656
rect 423 1652 427 1656
rect 519 1652 523 1656
rect 623 1652 627 1656
rect 727 1652 731 1656
rect 831 1652 835 1656
rect 935 1652 939 1656
rect 1047 1652 1051 1656
rect 1159 1652 1163 1656
rect 1287 1655 1291 1659
rect 111 1637 115 1641
rect 215 1640 219 1644
rect 271 1640 275 1644
rect 335 1640 339 1644
rect 407 1640 411 1644
rect 479 1640 483 1644
rect 559 1640 563 1644
rect 647 1640 651 1644
rect 743 1640 747 1644
rect 839 1640 843 1644
rect 943 1640 947 1644
rect 1055 1640 1059 1644
rect 1175 1640 1179 1644
rect 1287 1637 1291 1641
rect 111 1620 115 1624
rect 231 1619 235 1623
rect 287 1619 291 1623
rect 351 1619 355 1623
rect 423 1619 427 1623
rect 495 1619 499 1623
rect 575 1619 579 1623
rect 663 1619 667 1623
rect 759 1619 763 1623
rect 855 1619 859 1623
rect 959 1619 963 1623
rect 1071 1619 1075 1623
rect 1191 1619 1195 1623
rect 1287 1620 1291 1624
rect 1327 1616 1331 1620
rect 1367 1617 1371 1621
rect 1431 1617 1435 1621
rect 1519 1617 1523 1621
rect 1599 1617 1603 1621
rect 1679 1617 1683 1621
rect 1751 1617 1755 1621
rect 1839 1617 1843 1621
rect 1935 1617 1939 1621
rect 2055 1617 2059 1621
rect 2183 1617 2187 1621
rect 2327 1617 2331 1621
rect 2455 1617 2459 1621
rect 2503 1616 2507 1620
rect 1327 1599 1331 1603
rect 1351 1596 1355 1600
rect 1415 1596 1419 1600
rect 1503 1596 1507 1600
rect 1583 1596 1587 1600
rect 1663 1596 1667 1600
rect 1735 1596 1739 1600
rect 1823 1596 1827 1600
rect 1919 1596 1923 1600
rect 2039 1596 2043 1600
rect 2167 1596 2171 1600
rect 2311 1596 2315 1600
rect 2439 1596 2443 1600
rect 2503 1599 2507 1603
rect 1327 1577 1331 1581
rect 1351 1580 1355 1584
rect 1423 1580 1427 1584
rect 1527 1580 1531 1584
rect 1647 1580 1651 1584
rect 1783 1580 1787 1584
rect 1935 1580 1939 1584
rect 2103 1580 2107 1584
rect 2279 1580 2283 1584
rect 2439 1580 2443 1584
rect 2503 1577 2507 1581
rect 111 1568 115 1572
rect 287 1569 291 1573
rect 351 1569 355 1573
rect 423 1569 427 1573
rect 503 1569 507 1573
rect 599 1569 603 1573
rect 703 1569 707 1573
rect 815 1569 819 1573
rect 935 1569 939 1573
rect 1063 1569 1067 1573
rect 1191 1569 1195 1573
rect 1287 1568 1291 1572
rect 1327 1560 1331 1564
rect 1367 1559 1371 1563
rect 1439 1559 1443 1563
rect 1543 1559 1547 1563
rect 1663 1559 1667 1563
rect 1799 1559 1803 1563
rect 1951 1559 1955 1563
rect 2119 1559 2123 1563
rect 2295 1559 2299 1563
rect 2455 1559 2459 1563
rect 2503 1560 2507 1564
rect 111 1551 115 1555
rect 271 1548 275 1552
rect 335 1548 339 1552
rect 407 1548 411 1552
rect 487 1548 491 1552
rect 583 1548 587 1552
rect 687 1548 691 1552
rect 799 1548 803 1552
rect 919 1548 923 1552
rect 1047 1548 1051 1552
rect 1175 1548 1179 1552
rect 1287 1551 1291 1555
rect 111 1525 115 1529
rect 471 1528 475 1532
rect 551 1528 555 1532
rect 639 1528 643 1532
rect 735 1528 739 1532
rect 839 1528 843 1532
rect 951 1528 955 1532
rect 1063 1528 1067 1532
rect 1175 1528 1179 1532
rect 1287 1525 1291 1529
rect 111 1508 115 1512
rect 487 1507 491 1511
rect 567 1507 571 1511
rect 655 1507 659 1511
rect 751 1507 755 1511
rect 855 1507 859 1511
rect 967 1507 971 1511
rect 1079 1507 1083 1511
rect 1191 1507 1195 1511
rect 1287 1508 1291 1512
rect 1327 1508 1331 1512
rect 1367 1509 1371 1513
rect 1439 1509 1443 1513
rect 1543 1509 1547 1513
rect 1647 1509 1651 1513
rect 1751 1509 1755 1513
rect 1855 1509 1859 1513
rect 1959 1509 1963 1513
rect 2055 1509 2059 1513
rect 2151 1509 2155 1513
rect 2247 1509 2251 1513
rect 2343 1509 2347 1513
rect 2439 1509 2443 1513
rect 2503 1508 2507 1512
rect 1327 1491 1331 1495
rect 1351 1488 1355 1492
rect 1423 1488 1427 1492
rect 1527 1488 1531 1492
rect 1631 1488 1635 1492
rect 1735 1488 1739 1492
rect 1839 1488 1843 1492
rect 1943 1488 1947 1492
rect 2039 1488 2043 1492
rect 2135 1488 2139 1492
rect 2231 1488 2235 1492
rect 2327 1488 2331 1492
rect 2423 1488 2427 1492
rect 2503 1491 2507 1495
rect 1327 1469 1331 1473
rect 1351 1472 1355 1476
rect 1423 1472 1427 1476
rect 1519 1472 1523 1476
rect 1615 1472 1619 1476
rect 1711 1472 1715 1476
rect 1815 1472 1819 1476
rect 1927 1472 1931 1476
rect 2047 1472 2051 1476
rect 2175 1472 2179 1476
rect 2303 1472 2307 1476
rect 2439 1472 2443 1476
rect 2503 1469 2507 1473
rect 111 1456 115 1460
rect 375 1457 379 1461
rect 463 1457 467 1461
rect 559 1457 563 1461
rect 655 1457 659 1461
rect 751 1457 755 1461
rect 855 1457 859 1461
rect 959 1457 963 1461
rect 1063 1457 1067 1461
rect 1167 1457 1171 1461
rect 1287 1456 1291 1460
rect 1327 1452 1331 1456
rect 1367 1451 1371 1455
rect 1439 1451 1443 1455
rect 1535 1451 1539 1455
rect 1631 1451 1635 1455
rect 1727 1451 1731 1455
rect 1831 1451 1835 1455
rect 1943 1451 1947 1455
rect 2063 1451 2067 1455
rect 2191 1451 2195 1455
rect 2319 1451 2323 1455
rect 2455 1451 2459 1455
rect 2503 1452 2507 1456
rect 111 1439 115 1443
rect 359 1436 363 1440
rect 447 1436 451 1440
rect 543 1436 547 1440
rect 639 1436 643 1440
rect 735 1436 739 1440
rect 839 1436 843 1440
rect 943 1436 947 1440
rect 1047 1436 1051 1440
rect 1151 1436 1155 1440
rect 1287 1439 1291 1443
rect 111 1421 115 1425
rect 231 1424 235 1428
rect 319 1424 323 1428
rect 415 1424 419 1428
rect 511 1424 515 1428
rect 615 1424 619 1428
rect 711 1424 715 1428
rect 807 1424 811 1428
rect 895 1424 899 1428
rect 991 1424 995 1428
rect 1087 1424 1091 1428
rect 1287 1421 1291 1425
rect 111 1404 115 1408
rect 247 1403 251 1407
rect 335 1403 339 1407
rect 431 1403 435 1407
rect 527 1403 531 1407
rect 631 1403 635 1407
rect 727 1403 731 1407
rect 823 1403 827 1407
rect 911 1403 915 1407
rect 1007 1403 1011 1407
rect 1103 1403 1107 1407
rect 1287 1404 1291 1408
rect 1327 1396 1331 1400
rect 1367 1397 1371 1401
rect 1423 1397 1427 1401
rect 1503 1397 1507 1401
rect 1591 1397 1595 1401
rect 1679 1397 1683 1401
rect 1775 1397 1779 1401
rect 1879 1397 1883 1401
rect 1991 1397 1995 1401
rect 2111 1397 2115 1401
rect 2231 1397 2235 1401
rect 2351 1397 2355 1401
rect 2455 1397 2459 1401
rect 2503 1396 2507 1400
rect 1327 1379 1331 1383
rect 1351 1376 1355 1380
rect 1407 1376 1411 1380
rect 1487 1376 1491 1380
rect 1575 1376 1579 1380
rect 1663 1376 1667 1380
rect 1759 1376 1763 1380
rect 1863 1376 1867 1380
rect 1975 1376 1979 1380
rect 2095 1376 2099 1380
rect 2215 1376 2219 1380
rect 2335 1376 2339 1380
rect 2439 1376 2443 1380
rect 2503 1379 2507 1383
rect 111 1352 115 1356
rect 151 1353 155 1357
rect 215 1353 219 1357
rect 311 1353 315 1357
rect 407 1353 411 1357
rect 511 1353 515 1357
rect 607 1353 611 1357
rect 703 1353 707 1357
rect 799 1353 803 1357
rect 895 1353 899 1357
rect 1327 1357 1331 1361
rect 1351 1360 1355 1364
rect 1407 1360 1411 1364
rect 1479 1360 1483 1364
rect 1567 1360 1571 1364
rect 1655 1360 1659 1364
rect 1751 1360 1755 1364
rect 1855 1360 1859 1364
rect 1967 1360 1971 1364
rect 2079 1360 2083 1364
rect 2199 1360 2203 1364
rect 2327 1360 2331 1364
rect 2439 1360 2443 1364
rect 999 1353 1003 1357
rect 2503 1357 2507 1361
rect 1287 1352 1291 1356
rect 1327 1340 1331 1344
rect 111 1335 115 1339
rect 1367 1339 1371 1343
rect 135 1332 139 1336
rect 199 1332 203 1336
rect 295 1332 299 1336
rect 391 1332 395 1336
rect 495 1332 499 1336
rect 591 1332 595 1336
rect 687 1332 691 1336
rect 783 1332 787 1336
rect 879 1332 883 1336
rect 983 1332 987 1336
rect 1287 1335 1291 1339
rect 1423 1339 1427 1343
rect 1495 1339 1499 1343
rect 1583 1339 1587 1343
rect 1671 1339 1675 1343
rect 1767 1339 1771 1343
rect 1871 1339 1875 1343
rect 1983 1339 1987 1343
rect 2095 1339 2099 1343
rect 2215 1339 2219 1343
rect 2343 1339 2347 1343
rect 2455 1339 2459 1343
rect 2503 1340 2507 1344
rect 111 1317 115 1321
rect 135 1320 139 1324
rect 215 1320 219 1324
rect 319 1320 323 1324
rect 415 1320 419 1324
rect 511 1320 515 1324
rect 599 1320 603 1324
rect 687 1320 691 1324
rect 783 1320 787 1324
rect 879 1320 883 1324
rect 1287 1317 1291 1321
rect 111 1300 115 1304
rect 151 1299 155 1303
rect 231 1299 235 1303
rect 335 1299 339 1303
rect 431 1299 435 1303
rect 527 1299 531 1303
rect 615 1299 619 1303
rect 703 1299 707 1303
rect 799 1299 803 1303
rect 895 1299 899 1303
rect 1287 1300 1291 1304
rect 1327 1280 1331 1284
rect 1367 1281 1371 1285
rect 1423 1281 1427 1285
rect 1519 1281 1523 1285
rect 1615 1281 1619 1285
rect 1719 1281 1723 1285
rect 1823 1281 1827 1285
rect 1919 1281 1923 1285
rect 2015 1281 2019 1285
rect 2103 1281 2107 1285
rect 2183 1281 2187 1285
rect 2255 1281 2259 1285
rect 2327 1281 2331 1285
rect 2399 1281 2403 1285
rect 2455 1281 2459 1285
rect 2503 1280 2507 1284
rect 1327 1263 1331 1267
rect 1351 1260 1355 1264
rect 1407 1260 1411 1264
rect 1503 1260 1507 1264
rect 1599 1260 1603 1264
rect 1703 1260 1707 1264
rect 1807 1260 1811 1264
rect 1903 1260 1907 1264
rect 1999 1260 2003 1264
rect 2087 1260 2091 1264
rect 2167 1260 2171 1264
rect 2239 1260 2243 1264
rect 2311 1260 2315 1264
rect 2383 1260 2387 1264
rect 2439 1260 2443 1264
rect 2503 1263 2507 1267
rect 111 1248 115 1252
rect 191 1249 195 1253
rect 247 1249 251 1253
rect 303 1249 307 1253
rect 367 1249 371 1253
rect 439 1249 443 1253
rect 527 1249 531 1253
rect 639 1249 643 1253
rect 775 1249 779 1253
rect 927 1249 931 1253
rect 1095 1249 1099 1253
rect 1239 1249 1243 1253
rect 1287 1248 1291 1252
rect 111 1231 115 1235
rect 175 1228 179 1232
rect 231 1228 235 1232
rect 287 1228 291 1232
rect 351 1228 355 1232
rect 423 1228 427 1232
rect 511 1228 515 1232
rect 623 1228 627 1232
rect 759 1228 763 1232
rect 911 1228 915 1232
rect 1079 1228 1083 1232
rect 1223 1228 1227 1232
rect 1287 1231 1291 1235
rect 1327 1229 1331 1233
rect 1351 1232 1355 1236
rect 1447 1232 1451 1236
rect 1575 1232 1579 1236
rect 1695 1232 1699 1236
rect 1815 1232 1819 1236
rect 1927 1232 1931 1236
rect 2031 1232 2035 1236
rect 2127 1232 2131 1236
rect 2215 1232 2219 1236
rect 2295 1232 2299 1236
rect 2375 1232 2379 1236
rect 2439 1232 2443 1236
rect 2503 1229 2507 1233
rect 111 1213 115 1217
rect 351 1216 355 1220
rect 407 1216 411 1220
rect 463 1216 467 1220
rect 519 1216 523 1220
rect 575 1216 579 1220
rect 631 1216 635 1220
rect 687 1216 691 1220
rect 743 1216 747 1220
rect 799 1216 803 1220
rect 855 1216 859 1220
rect 911 1216 915 1220
rect 1287 1213 1291 1217
rect 1327 1212 1331 1216
rect 1367 1211 1371 1215
rect 1463 1211 1467 1215
rect 1591 1211 1595 1215
rect 1711 1211 1715 1215
rect 1831 1211 1835 1215
rect 1943 1211 1947 1215
rect 2047 1211 2051 1215
rect 2143 1211 2147 1215
rect 2231 1211 2235 1215
rect 2311 1211 2315 1215
rect 2391 1211 2395 1215
rect 2455 1211 2459 1215
rect 2503 1212 2507 1216
rect 111 1196 115 1200
rect 367 1195 371 1199
rect 423 1195 427 1199
rect 479 1195 483 1199
rect 535 1195 539 1199
rect 591 1195 595 1199
rect 647 1195 651 1199
rect 703 1195 707 1199
rect 759 1195 763 1199
rect 815 1195 819 1199
rect 871 1195 875 1199
rect 927 1195 931 1199
rect 1287 1196 1291 1200
rect 1327 1160 1331 1164
rect 1367 1161 1371 1165
rect 1471 1161 1475 1165
rect 1599 1161 1603 1165
rect 1735 1161 1739 1165
rect 1863 1161 1867 1165
rect 1983 1161 1987 1165
rect 2087 1161 2091 1165
rect 2191 1161 2195 1165
rect 2287 1161 2291 1165
rect 2383 1161 2387 1165
rect 2455 1161 2459 1165
rect 2503 1160 2507 1164
rect 111 1140 115 1144
rect 423 1141 427 1145
rect 479 1141 483 1145
rect 535 1141 539 1145
rect 591 1141 595 1145
rect 647 1141 651 1145
rect 703 1141 707 1145
rect 759 1141 763 1145
rect 815 1141 819 1145
rect 871 1141 875 1145
rect 927 1141 931 1145
rect 983 1141 987 1145
rect 1287 1140 1291 1144
rect 1327 1143 1331 1147
rect 1351 1140 1355 1144
rect 1455 1140 1459 1144
rect 1583 1140 1587 1144
rect 1719 1140 1723 1144
rect 1847 1140 1851 1144
rect 1967 1140 1971 1144
rect 2071 1140 2075 1144
rect 2175 1140 2179 1144
rect 2271 1140 2275 1144
rect 2367 1140 2371 1144
rect 2439 1140 2443 1144
rect 2503 1143 2507 1147
rect 111 1123 115 1127
rect 407 1120 411 1124
rect 463 1120 467 1124
rect 519 1120 523 1124
rect 575 1120 579 1124
rect 631 1120 635 1124
rect 687 1120 691 1124
rect 743 1120 747 1124
rect 799 1120 803 1124
rect 855 1120 859 1124
rect 911 1120 915 1124
rect 967 1120 971 1124
rect 1287 1123 1291 1127
rect 1327 1121 1331 1125
rect 1367 1124 1371 1128
rect 1447 1124 1451 1128
rect 1535 1124 1539 1128
rect 1631 1124 1635 1128
rect 1719 1124 1723 1128
rect 1807 1124 1811 1128
rect 1895 1124 1899 1128
rect 1983 1124 1987 1128
rect 2071 1124 2075 1128
rect 2159 1124 2163 1128
rect 2255 1124 2259 1128
rect 2359 1124 2363 1128
rect 2439 1124 2443 1128
rect 2503 1121 2507 1125
rect 111 1101 115 1105
rect 223 1104 227 1108
rect 311 1104 315 1108
rect 399 1104 403 1108
rect 495 1104 499 1108
rect 591 1104 595 1108
rect 679 1104 683 1108
rect 767 1104 771 1108
rect 847 1104 851 1108
rect 927 1104 931 1108
rect 1015 1104 1019 1108
rect 1103 1104 1107 1108
rect 1287 1101 1291 1105
rect 1327 1104 1331 1108
rect 1383 1103 1387 1107
rect 1463 1103 1467 1107
rect 1551 1103 1555 1107
rect 1647 1103 1651 1107
rect 1735 1103 1739 1107
rect 1823 1103 1827 1107
rect 1911 1103 1915 1107
rect 1999 1103 2003 1107
rect 2087 1103 2091 1107
rect 2175 1103 2179 1107
rect 2271 1103 2275 1107
rect 2375 1103 2379 1107
rect 2455 1103 2459 1107
rect 2503 1104 2507 1108
rect 111 1084 115 1088
rect 239 1083 243 1087
rect 327 1083 331 1087
rect 415 1083 419 1087
rect 511 1083 515 1087
rect 607 1083 611 1087
rect 695 1083 699 1087
rect 783 1083 787 1087
rect 863 1083 867 1087
rect 943 1083 947 1087
rect 1031 1083 1035 1087
rect 1119 1083 1123 1087
rect 1287 1084 1291 1088
rect 1327 1044 1331 1048
rect 1431 1045 1435 1049
rect 1495 1045 1499 1049
rect 1567 1045 1571 1049
rect 1639 1045 1643 1049
rect 1703 1045 1707 1049
rect 1767 1045 1771 1049
rect 1839 1045 1843 1049
rect 1919 1045 1923 1049
rect 2007 1045 2011 1049
rect 2111 1045 2115 1049
rect 2231 1045 2235 1049
rect 2351 1045 2355 1049
rect 2455 1045 2459 1049
rect 2503 1044 2507 1048
rect 111 1028 115 1032
rect 151 1029 155 1033
rect 207 1029 211 1033
rect 303 1029 307 1033
rect 415 1029 419 1033
rect 535 1029 539 1033
rect 655 1029 659 1033
rect 767 1029 771 1033
rect 879 1029 883 1033
rect 983 1029 987 1033
rect 1095 1029 1099 1033
rect 1207 1029 1211 1033
rect 1287 1028 1291 1032
rect 1327 1027 1331 1031
rect 1415 1024 1419 1028
rect 1479 1024 1483 1028
rect 1551 1024 1555 1028
rect 1623 1024 1627 1028
rect 1687 1024 1691 1028
rect 1751 1024 1755 1028
rect 1823 1024 1827 1028
rect 1903 1024 1907 1028
rect 1991 1024 1995 1028
rect 2095 1024 2099 1028
rect 2215 1024 2219 1028
rect 2335 1024 2339 1028
rect 2439 1024 2443 1028
rect 2503 1027 2507 1031
rect 111 1011 115 1015
rect 135 1008 139 1012
rect 191 1008 195 1012
rect 287 1008 291 1012
rect 399 1008 403 1012
rect 519 1008 523 1012
rect 639 1008 643 1012
rect 751 1008 755 1012
rect 863 1008 867 1012
rect 967 1008 971 1012
rect 1079 1008 1083 1012
rect 1191 1008 1195 1012
rect 1287 1011 1291 1015
rect 1327 1001 1331 1005
rect 1511 1004 1515 1008
rect 1567 1004 1571 1008
rect 1623 1004 1627 1008
rect 1679 1004 1683 1008
rect 1735 1004 1739 1008
rect 1807 1004 1811 1008
rect 1887 1004 1891 1008
rect 1983 1004 1987 1008
rect 2095 1004 2099 1008
rect 2215 1004 2219 1008
rect 2335 1004 2339 1008
rect 2439 1004 2443 1008
rect 2503 1001 2507 1005
rect 111 989 115 993
rect 135 992 139 996
rect 215 992 219 996
rect 327 992 331 996
rect 439 992 443 996
rect 551 992 555 996
rect 663 992 667 996
rect 759 992 763 996
rect 847 992 851 996
rect 935 992 939 996
rect 1015 992 1019 996
rect 1087 992 1091 996
rect 1167 992 1171 996
rect 1223 992 1227 996
rect 1287 989 1291 993
rect 1327 984 1331 988
rect 1527 983 1531 987
rect 1583 983 1587 987
rect 1639 983 1643 987
rect 1695 983 1699 987
rect 1751 983 1755 987
rect 1823 983 1827 987
rect 1903 983 1907 987
rect 1999 983 2003 987
rect 2111 983 2115 987
rect 2231 983 2235 987
rect 2351 983 2355 987
rect 2455 983 2459 987
rect 2503 984 2507 988
rect 111 972 115 976
rect 151 971 155 975
rect 231 971 235 975
rect 343 971 347 975
rect 455 971 459 975
rect 567 971 571 975
rect 679 971 683 975
rect 775 971 779 975
rect 863 971 867 975
rect 951 971 955 975
rect 1031 971 1035 975
rect 1103 971 1107 975
rect 1183 971 1187 975
rect 1239 971 1243 975
rect 1287 972 1291 976
rect 111 920 115 924
rect 151 921 155 925
rect 207 921 211 925
rect 295 921 299 925
rect 399 921 403 925
rect 511 921 515 925
rect 623 921 627 925
rect 735 921 739 925
rect 831 921 835 925
rect 927 921 931 925
rect 1015 921 1019 925
rect 1095 921 1099 925
rect 1175 921 1179 925
rect 1239 921 1243 925
rect 1287 920 1291 924
rect 1327 916 1331 920
rect 1367 917 1371 921
rect 1439 917 1443 921
rect 1527 917 1531 921
rect 1615 917 1619 921
rect 1695 917 1699 921
rect 1791 917 1795 921
rect 1895 917 1899 921
rect 2015 917 2019 921
rect 2151 917 2155 921
rect 2295 917 2299 921
rect 2439 917 2443 921
rect 2503 916 2507 920
rect 111 903 115 907
rect 135 900 139 904
rect 191 900 195 904
rect 279 900 283 904
rect 383 900 387 904
rect 495 900 499 904
rect 607 900 611 904
rect 719 900 723 904
rect 815 900 819 904
rect 911 900 915 904
rect 999 900 1003 904
rect 1079 900 1083 904
rect 1159 900 1163 904
rect 1223 900 1227 904
rect 1287 903 1291 907
rect 1327 899 1331 903
rect 1351 896 1355 900
rect 1423 896 1427 900
rect 1511 896 1515 900
rect 1599 896 1603 900
rect 1679 896 1683 900
rect 1775 896 1779 900
rect 1879 896 1883 900
rect 1999 896 2003 900
rect 2135 896 2139 900
rect 2279 896 2283 900
rect 2423 896 2427 900
rect 2503 899 2507 903
rect 111 881 115 885
rect 247 884 251 888
rect 343 884 347 888
rect 439 884 443 888
rect 543 884 547 888
rect 647 884 651 888
rect 743 884 747 888
rect 839 884 843 888
rect 927 884 931 888
rect 1007 884 1011 888
rect 1087 884 1091 888
rect 1167 884 1171 888
rect 1223 884 1227 888
rect 1287 881 1291 885
rect 1327 873 1331 877
rect 1487 876 1491 880
rect 1559 876 1563 880
rect 1623 876 1627 880
rect 1687 876 1691 880
rect 1751 876 1755 880
rect 1815 876 1819 880
rect 1887 876 1891 880
rect 1975 876 1979 880
rect 2079 876 2083 880
rect 2199 876 2203 880
rect 2319 876 2323 880
rect 2439 876 2443 880
rect 2503 873 2507 877
rect 111 864 115 868
rect 263 863 267 867
rect 359 863 363 867
rect 455 863 459 867
rect 559 863 563 867
rect 663 863 667 867
rect 759 863 763 867
rect 855 863 859 867
rect 943 863 947 867
rect 1023 863 1027 867
rect 1103 863 1107 867
rect 1183 863 1187 867
rect 1239 863 1243 867
rect 1287 864 1291 868
rect 1327 856 1331 860
rect 1503 855 1507 859
rect 1575 855 1579 859
rect 1639 855 1643 859
rect 1703 855 1707 859
rect 1767 855 1771 859
rect 1831 855 1835 859
rect 1903 855 1907 859
rect 1991 855 1995 859
rect 2095 855 2099 859
rect 2215 855 2219 859
rect 2335 855 2339 859
rect 2455 855 2459 859
rect 2503 856 2507 860
rect 111 808 115 812
rect 239 809 243 813
rect 303 809 307 813
rect 383 809 387 813
rect 463 809 467 813
rect 551 809 555 813
rect 639 809 643 813
rect 727 809 731 813
rect 807 809 811 813
rect 895 809 899 813
rect 983 809 987 813
rect 1071 809 1075 813
rect 1287 808 1291 812
rect 1327 796 1331 800
rect 1439 797 1443 801
rect 1511 797 1515 801
rect 1591 797 1595 801
rect 1671 797 1675 801
rect 1759 797 1763 801
rect 1847 797 1851 801
rect 1935 797 1939 801
rect 2023 797 2027 801
rect 2111 797 2115 801
rect 2199 797 2203 801
rect 2287 797 2291 801
rect 2383 797 2387 801
rect 2455 797 2459 801
rect 2503 796 2507 800
rect 111 791 115 795
rect 223 788 227 792
rect 287 788 291 792
rect 367 788 371 792
rect 447 788 451 792
rect 535 788 539 792
rect 623 788 627 792
rect 711 788 715 792
rect 791 788 795 792
rect 879 788 883 792
rect 967 788 971 792
rect 1055 788 1059 792
rect 1287 791 1291 795
rect 1327 779 1331 783
rect 111 769 115 773
rect 151 772 155 776
rect 247 772 251 776
rect 343 772 347 776
rect 439 772 443 776
rect 527 772 531 776
rect 607 772 611 776
rect 679 772 683 776
rect 751 772 755 776
rect 823 772 827 776
rect 895 772 899 776
rect 975 772 979 776
rect 1423 776 1427 780
rect 1495 776 1499 780
rect 1575 776 1579 780
rect 1655 776 1659 780
rect 1743 776 1747 780
rect 1831 776 1835 780
rect 1919 776 1923 780
rect 2007 776 2011 780
rect 2095 776 2099 780
rect 2183 776 2187 780
rect 2271 776 2275 780
rect 2367 776 2371 780
rect 2439 776 2443 780
rect 2503 779 2507 783
rect 1287 769 1291 773
rect 1327 757 1331 761
rect 1351 760 1355 764
rect 1447 760 1451 764
rect 1567 760 1571 764
rect 1687 760 1691 764
rect 1807 760 1811 764
rect 1927 760 1931 764
rect 2039 760 2043 764
rect 2143 760 2147 764
rect 2247 760 2251 764
rect 2351 760 2355 764
rect 2439 760 2443 764
rect 2503 757 2507 761
rect 111 752 115 756
rect 167 751 171 755
rect 263 751 267 755
rect 359 751 363 755
rect 455 751 459 755
rect 543 751 547 755
rect 623 751 627 755
rect 695 751 699 755
rect 767 751 771 755
rect 839 751 843 755
rect 911 751 915 755
rect 991 751 995 755
rect 1287 752 1291 756
rect 1327 740 1331 744
rect 1367 739 1371 743
rect 1463 739 1467 743
rect 1583 739 1587 743
rect 1703 739 1707 743
rect 1823 739 1827 743
rect 1943 739 1947 743
rect 2055 739 2059 743
rect 2159 739 2163 743
rect 2263 739 2267 743
rect 2367 739 2371 743
rect 2455 739 2459 743
rect 2503 740 2507 744
rect 111 696 115 700
rect 175 697 179 701
rect 263 697 267 701
rect 343 697 347 701
rect 423 697 427 701
rect 503 697 507 701
rect 575 697 579 701
rect 639 697 643 701
rect 703 697 707 701
rect 767 697 771 701
rect 839 697 843 701
rect 911 697 915 701
rect 1287 696 1291 700
rect 1327 684 1331 688
rect 1367 685 1371 689
rect 1431 685 1435 689
rect 1535 685 1539 689
rect 1639 685 1643 689
rect 1751 685 1755 689
rect 1863 685 1867 689
rect 1967 685 1971 689
rect 2063 685 2067 689
rect 2151 685 2155 689
rect 2231 685 2235 689
rect 2311 685 2315 689
rect 2391 685 2395 689
rect 2455 685 2459 689
rect 2503 684 2507 688
rect 111 679 115 683
rect 159 676 163 680
rect 247 676 251 680
rect 327 676 331 680
rect 407 676 411 680
rect 487 676 491 680
rect 559 676 563 680
rect 623 676 627 680
rect 687 676 691 680
rect 751 676 755 680
rect 823 676 827 680
rect 895 676 899 680
rect 1287 679 1291 683
rect 111 661 115 665
rect 215 664 219 668
rect 295 664 299 668
rect 375 664 379 668
rect 455 664 459 668
rect 527 664 531 668
rect 591 664 595 668
rect 655 664 659 668
rect 719 664 723 668
rect 783 664 787 668
rect 847 664 851 668
rect 919 664 923 668
rect 1327 667 1331 671
rect 1287 661 1291 665
rect 1351 664 1355 668
rect 1415 664 1419 668
rect 1519 664 1523 668
rect 1623 664 1627 668
rect 1735 664 1739 668
rect 1847 664 1851 668
rect 1951 664 1955 668
rect 2047 664 2051 668
rect 2135 664 2139 668
rect 2215 664 2219 668
rect 2295 664 2299 668
rect 2375 664 2379 668
rect 2439 664 2443 668
rect 2503 667 2507 671
rect 111 644 115 648
rect 231 643 235 647
rect 311 643 315 647
rect 391 643 395 647
rect 471 643 475 647
rect 543 643 547 647
rect 607 643 611 647
rect 671 643 675 647
rect 735 643 739 647
rect 799 643 803 647
rect 863 643 867 647
rect 935 643 939 647
rect 1287 644 1291 648
rect 1327 641 1331 645
rect 1479 644 1483 648
rect 1559 644 1563 648
rect 1647 644 1651 648
rect 1735 644 1739 648
rect 1831 644 1835 648
rect 1919 644 1923 648
rect 2007 644 2011 648
rect 2087 644 2091 648
rect 2167 644 2171 648
rect 2239 644 2243 648
rect 2311 644 2315 648
rect 2383 644 2387 648
rect 2439 644 2443 648
rect 2503 641 2507 645
rect 1327 624 1331 628
rect 1495 623 1499 627
rect 1575 623 1579 627
rect 1663 623 1667 627
rect 1751 623 1755 627
rect 1847 623 1851 627
rect 1935 623 1939 627
rect 2023 623 2027 627
rect 2103 623 2107 627
rect 2183 623 2187 627
rect 2255 623 2259 627
rect 2327 623 2331 627
rect 2399 623 2403 627
rect 2455 623 2459 627
rect 2503 624 2507 628
rect 111 588 115 592
rect 207 589 211 593
rect 303 589 307 593
rect 407 589 411 593
rect 503 589 507 593
rect 599 589 603 593
rect 687 589 691 593
rect 767 589 771 593
rect 847 589 851 593
rect 927 589 931 593
rect 1007 589 1011 593
rect 1087 589 1091 593
rect 1287 588 1291 592
rect 111 571 115 575
rect 191 568 195 572
rect 287 568 291 572
rect 391 568 395 572
rect 487 568 491 572
rect 583 568 587 572
rect 671 568 675 572
rect 751 568 755 572
rect 831 568 835 572
rect 911 568 915 572
rect 991 568 995 572
rect 1071 568 1075 572
rect 1287 571 1291 575
rect 1327 568 1331 572
rect 1455 569 1459 573
rect 1559 569 1563 573
rect 1671 569 1675 573
rect 1775 569 1779 573
rect 1879 569 1883 573
rect 1983 569 1987 573
rect 2087 569 2091 573
rect 2183 569 2187 573
rect 2279 569 2283 573
rect 2375 569 2379 573
rect 2455 569 2459 573
rect 2503 568 2507 572
rect 111 549 115 553
rect 175 552 179 556
rect 271 552 275 556
rect 375 552 379 556
rect 487 552 491 556
rect 591 552 595 556
rect 695 552 699 556
rect 791 552 795 556
rect 879 552 883 556
rect 967 552 971 556
rect 1055 552 1059 556
rect 1151 552 1155 556
rect 1287 549 1291 553
rect 1327 551 1331 555
rect 1439 548 1443 552
rect 1543 548 1547 552
rect 1655 548 1659 552
rect 1759 548 1763 552
rect 1863 548 1867 552
rect 1967 548 1971 552
rect 2071 548 2075 552
rect 2167 548 2171 552
rect 2263 548 2267 552
rect 2359 548 2363 552
rect 2439 548 2443 552
rect 2503 551 2507 555
rect 111 532 115 536
rect 191 531 195 535
rect 287 531 291 535
rect 391 531 395 535
rect 503 531 507 535
rect 607 531 611 535
rect 711 531 715 535
rect 807 531 811 535
rect 895 531 899 535
rect 983 531 987 535
rect 1071 531 1075 535
rect 1167 531 1171 535
rect 1287 532 1291 536
rect 1327 529 1331 533
rect 1367 532 1371 536
rect 1447 532 1451 536
rect 1527 532 1531 536
rect 1615 532 1619 536
rect 1711 532 1715 536
rect 1799 532 1803 536
rect 1887 532 1891 536
rect 1975 532 1979 536
rect 2063 532 2067 536
rect 2151 532 2155 536
rect 2247 532 2251 536
rect 2343 532 2347 536
rect 2439 532 2443 536
rect 2503 529 2507 533
rect 1327 512 1331 516
rect 1383 511 1387 515
rect 1463 511 1467 515
rect 1543 511 1547 515
rect 1631 511 1635 515
rect 1727 511 1731 515
rect 1815 511 1819 515
rect 1903 511 1907 515
rect 1991 511 1995 515
rect 2079 511 2083 515
rect 2167 511 2171 515
rect 2263 511 2267 515
rect 2359 511 2363 515
rect 2455 511 2459 515
rect 2503 512 2507 516
rect 111 476 115 480
rect 151 477 155 481
rect 247 477 251 481
rect 367 477 371 481
rect 487 477 491 481
rect 615 477 619 481
rect 735 477 739 481
rect 847 477 851 481
rect 951 477 955 481
rect 1055 477 1059 481
rect 1159 477 1163 481
rect 1239 477 1243 481
rect 1287 476 1291 480
rect 111 459 115 463
rect 135 456 139 460
rect 231 456 235 460
rect 351 456 355 460
rect 471 456 475 460
rect 599 456 603 460
rect 719 456 723 460
rect 831 456 835 460
rect 935 456 939 460
rect 1039 456 1043 460
rect 1143 456 1147 460
rect 1223 456 1227 460
rect 1287 459 1291 463
rect 1327 456 1331 460
rect 1367 457 1371 461
rect 1431 457 1435 461
rect 1519 457 1523 461
rect 1615 457 1619 461
rect 1711 457 1715 461
rect 1815 457 1819 461
rect 1927 457 1931 461
rect 2055 457 2059 461
rect 2191 457 2195 461
rect 2335 457 2339 461
rect 2455 457 2459 461
rect 2503 456 2507 460
rect 111 437 115 441
rect 135 440 139 444
rect 191 440 195 444
rect 247 440 251 444
rect 303 440 307 444
rect 383 440 387 444
rect 471 440 475 444
rect 567 440 571 444
rect 671 440 675 444
rect 783 440 787 444
rect 895 440 899 444
rect 1007 440 1011 444
rect 1127 440 1131 444
rect 1223 440 1227 444
rect 1287 437 1291 441
rect 1327 439 1331 443
rect 1351 436 1355 440
rect 1415 436 1419 440
rect 1503 436 1507 440
rect 1599 436 1603 440
rect 1695 436 1699 440
rect 1799 436 1803 440
rect 1911 436 1915 440
rect 2039 436 2043 440
rect 2175 436 2179 440
rect 2319 436 2323 440
rect 2439 436 2443 440
rect 2503 439 2507 443
rect 111 420 115 424
rect 151 419 155 423
rect 207 419 211 423
rect 263 419 267 423
rect 319 419 323 423
rect 399 419 403 423
rect 487 419 491 423
rect 583 419 587 423
rect 687 419 691 423
rect 799 419 803 423
rect 911 419 915 423
rect 1023 419 1027 423
rect 1143 419 1147 423
rect 1239 419 1243 423
rect 1287 420 1291 424
rect 1327 417 1331 421
rect 1351 420 1355 424
rect 1423 420 1427 424
rect 1511 420 1515 424
rect 1599 420 1603 424
rect 1679 420 1683 424
rect 1775 420 1779 424
rect 1887 420 1891 424
rect 2015 420 2019 424
rect 2159 420 2163 424
rect 2311 420 2315 424
rect 2439 420 2443 424
rect 2503 417 2507 421
rect 1327 400 1331 404
rect 1367 399 1371 403
rect 1439 399 1443 403
rect 1527 399 1531 403
rect 1615 399 1619 403
rect 1695 399 1699 403
rect 1791 399 1795 403
rect 1903 399 1907 403
rect 2031 399 2035 403
rect 2175 399 2179 403
rect 2327 399 2331 403
rect 2455 399 2459 403
rect 2503 400 2507 404
rect 111 360 115 364
rect 151 361 155 365
rect 207 361 211 365
rect 279 361 283 365
rect 359 361 363 365
rect 431 361 435 365
rect 511 361 515 365
rect 591 361 595 365
rect 671 361 675 365
rect 751 361 755 365
rect 823 361 827 365
rect 895 361 899 365
rect 967 361 971 365
rect 1039 361 1043 365
rect 1111 361 1115 365
rect 1183 361 1187 365
rect 1239 361 1243 365
rect 1287 360 1291 364
rect 111 343 115 347
rect 135 340 139 344
rect 191 340 195 344
rect 263 340 267 344
rect 343 340 347 344
rect 415 340 419 344
rect 495 340 499 344
rect 575 340 579 344
rect 655 340 659 344
rect 735 340 739 344
rect 807 340 811 344
rect 879 340 883 344
rect 951 340 955 344
rect 1023 340 1027 344
rect 1095 340 1099 344
rect 1167 340 1171 344
rect 1223 340 1227 344
rect 1287 343 1291 347
rect 1327 344 1331 348
rect 1679 345 1683 349
rect 1735 345 1739 349
rect 1807 345 1811 349
rect 1903 345 1907 349
rect 2023 345 2027 349
rect 2159 345 2163 349
rect 2303 345 2307 349
rect 2455 345 2459 349
rect 2503 344 2507 348
rect 1327 327 1331 331
rect 111 317 115 321
rect 135 320 139 324
rect 199 320 203 324
rect 287 320 291 324
rect 375 320 379 324
rect 455 320 459 324
rect 543 320 547 324
rect 631 320 635 324
rect 727 320 731 324
rect 823 320 827 324
rect 927 320 931 324
rect 1031 320 1035 324
rect 1135 320 1139 324
rect 1223 320 1227 324
rect 1663 324 1667 328
rect 1719 324 1723 328
rect 1791 324 1795 328
rect 1887 324 1891 328
rect 2007 324 2011 328
rect 2143 324 2147 328
rect 2287 324 2291 328
rect 2439 324 2443 328
rect 2503 327 2507 331
rect 1287 317 1291 321
rect 1327 309 1331 313
rect 1351 312 1355 316
rect 1431 312 1435 316
rect 1527 312 1531 316
rect 1623 312 1627 316
rect 1711 312 1715 316
rect 1807 312 1811 316
rect 1911 312 1915 316
rect 2023 312 2027 316
rect 2151 312 2155 316
rect 2287 312 2291 316
rect 2423 312 2427 316
rect 2503 309 2507 313
rect 111 300 115 304
rect 151 299 155 303
rect 215 299 219 303
rect 303 299 307 303
rect 391 299 395 303
rect 471 299 475 303
rect 559 299 563 303
rect 647 299 651 303
rect 743 299 747 303
rect 839 299 843 303
rect 943 299 947 303
rect 1047 299 1051 303
rect 1151 299 1155 303
rect 1239 299 1243 303
rect 1287 300 1291 304
rect 1327 292 1331 296
rect 1367 291 1371 295
rect 1447 291 1451 295
rect 1543 291 1547 295
rect 1639 291 1643 295
rect 1727 291 1731 295
rect 1823 291 1827 295
rect 1927 291 1931 295
rect 2039 291 2043 295
rect 2167 291 2171 295
rect 2303 291 2307 295
rect 2439 291 2443 295
rect 2503 292 2507 296
rect 111 240 115 244
rect 151 241 155 245
rect 231 241 235 245
rect 327 241 331 245
rect 423 241 427 245
rect 519 241 523 245
rect 615 241 619 245
rect 711 241 715 245
rect 807 241 811 245
rect 903 241 907 245
rect 1007 241 1011 245
rect 1111 241 1115 245
rect 1215 241 1219 245
rect 1287 240 1291 244
rect 1327 236 1331 240
rect 1367 237 1371 241
rect 1439 237 1443 241
rect 1535 237 1539 241
rect 1631 237 1635 241
rect 1727 237 1731 241
rect 1815 237 1819 241
rect 1903 237 1907 241
rect 1999 237 2003 241
rect 2103 237 2107 241
rect 2215 237 2219 241
rect 2335 237 2339 241
rect 2455 237 2459 241
rect 2503 236 2507 240
rect 111 223 115 227
rect 135 220 139 224
rect 215 220 219 224
rect 311 220 315 224
rect 407 220 411 224
rect 503 220 507 224
rect 599 220 603 224
rect 695 220 699 224
rect 791 220 795 224
rect 887 220 891 224
rect 991 220 995 224
rect 1095 220 1099 224
rect 1199 220 1203 224
rect 1287 223 1291 227
rect 1327 219 1331 223
rect 1351 216 1355 220
rect 1423 216 1427 220
rect 1519 216 1523 220
rect 1615 216 1619 220
rect 1711 216 1715 220
rect 1799 216 1803 220
rect 1887 216 1891 220
rect 1983 216 1987 220
rect 2087 216 2091 220
rect 2199 216 2203 220
rect 2319 216 2323 220
rect 2439 216 2443 220
rect 2503 219 2507 223
rect 111 197 115 201
rect 159 200 163 204
rect 239 200 243 204
rect 327 200 331 204
rect 415 200 419 204
rect 511 200 515 204
rect 607 200 611 204
rect 695 200 699 204
rect 783 200 787 204
rect 871 200 875 204
rect 959 200 963 204
rect 1047 200 1051 204
rect 1135 200 1139 204
rect 1287 197 1291 201
rect 1327 197 1331 201
rect 1391 200 1395 204
rect 1495 200 1499 204
rect 1599 200 1603 204
rect 1711 200 1715 204
rect 1815 200 1819 204
rect 1919 200 1923 204
rect 2015 200 2019 204
rect 2111 200 2115 204
rect 2199 200 2203 204
rect 2287 200 2291 204
rect 2375 200 2379 204
rect 2439 200 2443 204
rect 2503 197 2507 201
rect 111 180 115 184
rect 175 179 179 183
rect 255 179 259 183
rect 343 179 347 183
rect 431 179 435 183
rect 527 179 531 183
rect 623 179 627 183
rect 711 179 715 183
rect 799 179 803 183
rect 887 179 891 183
rect 975 179 979 183
rect 1063 179 1067 183
rect 1151 179 1155 183
rect 1287 180 1291 184
rect 1327 180 1331 184
rect 1407 179 1411 183
rect 1511 179 1515 183
rect 1615 179 1619 183
rect 1727 179 1731 183
rect 1831 179 1835 183
rect 1935 179 1939 183
rect 2031 179 2035 183
rect 2127 179 2131 183
rect 2215 179 2219 183
rect 2303 179 2307 183
rect 2391 179 2395 183
rect 2455 179 2459 183
rect 2503 180 2507 184
rect 111 108 115 112
rect 151 109 155 113
rect 207 109 211 113
rect 263 109 267 113
rect 319 109 323 113
rect 375 109 379 113
rect 431 109 435 113
rect 487 109 491 113
rect 551 109 555 113
rect 623 109 627 113
rect 687 109 691 113
rect 751 109 755 113
rect 815 109 819 113
rect 879 109 883 113
rect 943 109 947 113
rect 1007 109 1011 113
rect 1071 109 1075 113
rect 1135 109 1139 113
rect 1199 109 1203 113
rect 1287 108 1291 112
rect 1327 108 1331 112
rect 1367 109 1371 113
rect 1423 109 1427 113
rect 1479 109 1483 113
rect 1535 109 1539 113
rect 1591 109 1595 113
rect 1647 109 1651 113
rect 1703 109 1707 113
rect 1759 109 1763 113
rect 1815 109 1819 113
rect 1871 109 1875 113
rect 1927 109 1931 113
rect 1983 109 1987 113
rect 2039 109 2043 113
rect 2095 109 2099 113
rect 2159 109 2163 113
rect 2223 109 2227 113
rect 2287 109 2291 113
rect 2343 109 2347 113
rect 2399 109 2403 113
rect 2455 109 2459 113
rect 2503 108 2507 112
rect 111 91 115 95
rect 135 88 139 92
rect 191 88 195 92
rect 247 88 251 92
rect 303 88 307 92
rect 359 88 363 92
rect 415 88 419 92
rect 471 88 475 92
rect 535 88 539 92
rect 607 88 611 92
rect 671 88 675 92
rect 735 88 739 92
rect 799 88 803 92
rect 863 88 867 92
rect 927 88 931 92
rect 991 88 995 92
rect 1055 88 1059 92
rect 1119 88 1123 92
rect 1183 88 1187 92
rect 1287 91 1291 95
rect 1327 91 1331 95
rect 1351 88 1355 92
rect 1407 88 1411 92
rect 1463 88 1467 92
rect 1519 88 1523 92
rect 1575 88 1579 92
rect 1631 88 1635 92
rect 1687 88 1691 92
rect 1743 88 1747 92
rect 1799 88 1803 92
rect 1855 88 1859 92
rect 1911 88 1915 92
rect 1967 88 1971 92
rect 2023 88 2027 92
rect 2079 88 2083 92
rect 2143 88 2147 92
rect 2207 88 2211 92
rect 2271 88 2275 92
rect 2327 88 2331 92
rect 2383 88 2387 92
rect 2439 88 2443 92
rect 2503 91 2507 95
<< m3 >>
rect 111 2582 115 2583
rect 111 2577 115 2578
rect 719 2582 723 2583
rect 719 2577 723 2578
rect 775 2582 779 2583
rect 775 2577 779 2578
rect 831 2582 835 2583
rect 831 2577 835 2578
rect 887 2582 891 2583
rect 887 2577 891 2578
rect 943 2582 947 2583
rect 943 2577 947 2578
rect 1287 2582 1291 2583
rect 1287 2577 1291 2578
rect 112 2557 114 2577
rect 720 2558 722 2577
rect 776 2558 778 2577
rect 832 2558 834 2577
rect 888 2558 890 2577
rect 944 2558 946 2577
rect 718 2557 724 2558
rect 110 2556 116 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 718 2553 719 2557
rect 723 2553 724 2557
rect 718 2552 724 2553
rect 774 2557 780 2558
rect 774 2553 775 2557
rect 779 2553 780 2557
rect 774 2552 780 2553
rect 830 2557 836 2558
rect 830 2553 831 2557
rect 835 2553 836 2557
rect 830 2552 836 2553
rect 886 2557 892 2558
rect 886 2553 887 2557
rect 891 2553 892 2557
rect 886 2552 892 2553
rect 942 2557 948 2558
rect 1288 2557 1290 2577
rect 1327 2558 1331 2559
rect 942 2553 943 2557
rect 947 2553 948 2557
rect 942 2552 948 2553
rect 1286 2556 1292 2557
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1327 2553 1331 2554
rect 1399 2558 1403 2559
rect 1399 2553 1403 2554
rect 1455 2558 1459 2559
rect 1455 2553 1459 2554
rect 1511 2558 1515 2559
rect 1511 2553 1515 2554
rect 1567 2558 1571 2559
rect 1567 2553 1571 2554
rect 1623 2558 1627 2559
rect 1623 2553 1627 2554
rect 1679 2558 1683 2559
rect 1679 2553 1683 2554
rect 1735 2558 1739 2559
rect 1735 2553 1739 2554
rect 1791 2558 1795 2559
rect 1791 2553 1795 2554
rect 1847 2558 1851 2559
rect 1847 2553 1851 2554
rect 1903 2558 1907 2559
rect 1903 2553 1907 2554
rect 1959 2558 1963 2559
rect 1959 2553 1963 2554
rect 2015 2558 2019 2559
rect 2015 2553 2019 2554
rect 2071 2558 2075 2559
rect 2071 2553 2075 2554
rect 2127 2558 2131 2559
rect 2127 2553 2131 2554
rect 2183 2558 2187 2559
rect 2183 2553 2187 2554
rect 2503 2558 2507 2559
rect 2503 2553 2507 2554
rect 110 2551 116 2552
rect 1286 2551 1292 2552
rect 110 2539 116 2540
rect 110 2535 111 2539
rect 115 2535 116 2539
rect 1286 2539 1292 2540
rect 110 2534 116 2535
rect 702 2536 708 2537
rect 112 2531 114 2534
rect 702 2532 703 2536
rect 707 2532 708 2536
rect 702 2531 708 2532
rect 758 2536 764 2537
rect 758 2532 759 2536
rect 763 2532 764 2536
rect 758 2531 764 2532
rect 814 2536 820 2537
rect 814 2532 815 2536
rect 819 2532 820 2536
rect 814 2531 820 2532
rect 870 2536 876 2537
rect 870 2532 871 2536
rect 875 2532 876 2536
rect 870 2531 876 2532
rect 926 2536 932 2537
rect 926 2532 927 2536
rect 931 2532 932 2536
rect 1286 2535 1287 2539
rect 1291 2535 1292 2539
rect 1286 2534 1292 2535
rect 926 2531 932 2532
rect 1288 2531 1290 2534
rect 1328 2533 1330 2553
rect 1400 2534 1402 2553
rect 1456 2534 1458 2553
rect 1512 2534 1514 2553
rect 1568 2534 1570 2553
rect 1624 2534 1626 2553
rect 1680 2534 1682 2553
rect 1736 2534 1738 2553
rect 1792 2534 1794 2553
rect 1848 2534 1850 2553
rect 1904 2534 1906 2553
rect 1960 2534 1962 2553
rect 2016 2534 2018 2553
rect 2072 2534 2074 2553
rect 2128 2534 2130 2553
rect 2184 2534 2186 2553
rect 1398 2533 1404 2534
rect 1326 2532 1332 2533
rect 111 2530 115 2531
rect 111 2525 115 2526
rect 167 2530 171 2531
rect 167 2525 171 2526
rect 223 2530 227 2531
rect 223 2525 227 2526
rect 279 2530 283 2531
rect 279 2525 283 2526
rect 343 2530 347 2531
rect 343 2525 347 2526
rect 407 2530 411 2531
rect 407 2525 411 2526
rect 479 2530 483 2531
rect 479 2525 483 2526
rect 559 2530 563 2531
rect 559 2525 563 2526
rect 639 2530 643 2531
rect 639 2525 643 2526
rect 703 2530 707 2531
rect 703 2525 707 2526
rect 719 2530 723 2531
rect 719 2525 723 2526
rect 759 2530 763 2531
rect 759 2525 763 2526
rect 799 2530 803 2531
rect 799 2525 803 2526
rect 815 2530 819 2531
rect 815 2525 819 2526
rect 871 2530 875 2531
rect 871 2525 875 2526
rect 879 2530 883 2531
rect 879 2525 883 2526
rect 927 2530 931 2531
rect 927 2525 931 2526
rect 959 2530 963 2531
rect 959 2525 963 2526
rect 1039 2530 1043 2531
rect 1039 2525 1043 2526
rect 1287 2530 1291 2531
rect 1326 2528 1327 2532
rect 1331 2528 1332 2532
rect 1398 2529 1399 2533
rect 1403 2529 1404 2533
rect 1398 2528 1404 2529
rect 1454 2533 1460 2534
rect 1454 2529 1455 2533
rect 1459 2529 1460 2533
rect 1454 2528 1460 2529
rect 1510 2533 1516 2534
rect 1510 2529 1511 2533
rect 1515 2529 1516 2533
rect 1510 2528 1516 2529
rect 1566 2533 1572 2534
rect 1566 2529 1567 2533
rect 1571 2529 1572 2533
rect 1566 2528 1572 2529
rect 1622 2533 1628 2534
rect 1622 2529 1623 2533
rect 1627 2529 1628 2533
rect 1622 2528 1628 2529
rect 1678 2533 1684 2534
rect 1678 2529 1679 2533
rect 1683 2529 1684 2533
rect 1678 2528 1684 2529
rect 1734 2533 1740 2534
rect 1734 2529 1735 2533
rect 1739 2529 1740 2533
rect 1734 2528 1740 2529
rect 1790 2533 1796 2534
rect 1790 2529 1791 2533
rect 1795 2529 1796 2533
rect 1790 2528 1796 2529
rect 1846 2533 1852 2534
rect 1846 2529 1847 2533
rect 1851 2529 1852 2533
rect 1846 2528 1852 2529
rect 1902 2533 1908 2534
rect 1902 2529 1903 2533
rect 1907 2529 1908 2533
rect 1902 2528 1908 2529
rect 1958 2533 1964 2534
rect 1958 2529 1959 2533
rect 1963 2529 1964 2533
rect 1958 2528 1964 2529
rect 2014 2533 2020 2534
rect 2014 2529 2015 2533
rect 2019 2529 2020 2533
rect 2014 2528 2020 2529
rect 2070 2533 2076 2534
rect 2070 2529 2071 2533
rect 2075 2529 2076 2533
rect 2070 2528 2076 2529
rect 2126 2533 2132 2534
rect 2126 2529 2127 2533
rect 2131 2529 2132 2533
rect 2126 2528 2132 2529
rect 2182 2533 2188 2534
rect 2504 2533 2506 2553
rect 2182 2529 2183 2533
rect 2187 2529 2188 2533
rect 2182 2528 2188 2529
rect 2502 2532 2508 2533
rect 2502 2528 2503 2532
rect 2507 2528 2508 2532
rect 1326 2527 1332 2528
rect 2502 2527 2508 2528
rect 1287 2525 1291 2526
rect 112 2522 114 2525
rect 166 2524 172 2525
rect 110 2521 116 2522
rect 110 2517 111 2521
rect 115 2517 116 2521
rect 166 2520 167 2524
rect 171 2520 172 2524
rect 166 2519 172 2520
rect 222 2524 228 2525
rect 222 2520 223 2524
rect 227 2520 228 2524
rect 222 2519 228 2520
rect 278 2524 284 2525
rect 278 2520 279 2524
rect 283 2520 284 2524
rect 278 2519 284 2520
rect 342 2524 348 2525
rect 342 2520 343 2524
rect 347 2520 348 2524
rect 342 2519 348 2520
rect 406 2524 412 2525
rect 406 2520 407 2524
rect 411 2520 412 2524
rect 406 2519 412 2520
rect 478 2524 484 2525
rect 478 2520 479 2524
rect 483 2520 484 2524
rect 478 2519 484 2520
rect 558 2524 564 2525
rect 558 2520 559 2524
rect 563 2520 564 2524
rect 558 2519 564 2520
rect 638 2524 644 2525
rect 638 2520 639 2524
rect 643 2520 644 2524
rect 638 2519 644 2520
rect 718 2524 724 2525
rect 718 2520 719 2524
rect 723 2520 724 2524
rect 718 2519 724 2520
rect 798 2524 804 2525
rect 798 2520 799 2524
rect 803 2520 804 2524
rect 798 2519 804 2520
rect 878 2524 884 2525
rect 878 2520 879 2524
rect 883 2520 884 2524
rect 878 2519 884 2520
rect 958 2524 964 2525
rect 958 2520 959 2524
rect 963 2520 964 2524
rect 958 2519 964 2520
rect 1038 2524 1044 2525
rect 1038 2520 1039 2524
rect 1043 2520 1044 2524
rect 1288 2522 1290 2525
rect 1038 2519 1044 2520
rect 1286 2521 1292 2522
rect 110 2516 116 2517
rect 1286 2517 1287 2521
rect 1291 2517 1292 2521
rect 1286 2516 1292 2517
rect 1326 2515 1332 2516
rect 1326 2511 1327 2515
rect 1331 2511 1332 2515
rect 2502 2515 2508 2516
rect 1326 2510 1332 2511
rect 1382 2512 1388 2513
rect 110 2504 116 2505
rect 1286 2504 1292 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 110 2499 116 2500
rect 182 2503 188 2504
rect 182 2499 183 2503
rect 187 2499 188 2503
rect 112 2479 114 2499
rect 182 2498 188 2499
rect 238 2503 244 2504
rect 238 2499 239 2503
rect 243 2499 244 2503
rect 238 2498 244 2499
rect 294 2503 300 2504
rect 294 2499 295 2503
rect 299 2499 300 2503
rect 294 2498 300 2499
rect 358 2503 364 2504
rect 358 2499 359 2503
rect 363 2499 364 2503
rect 358 2498 364 2499
rect 422 2503 428 2504
rect 422 2499 423 2503
rect 427 2499 428 2503
rect 422 2498 428 2499
rect 494 2503 500 2504
rect 494 2499 495 2503
rect 499 2499 500 2503
rect 494 2498 500 2499
rect 574 2503 580 2504
rect 574 2499 575 2503
rect 579 2499 580 2503
rect 574 2498 580 2499
rect 654 2503 660 2504
rect 654 2499 655 2503
rect 659 2499 660 2503
rect 654 2498 660 2499
rect 734 2503 740 2504
rect 734 2499 735 2503
rect 739 2499 740 2503
rect 734 2498 740 2499
rect 814 2503 820 2504
rect 814 2499 815 2503
rect 819 2499 820 2503
rect 814 2498 820 2499
rect 894 2503 900 2504
rect 894 2499 895 2503
rect 899 2499 900 2503
rect 894 2498 900 2499
rect 974 2503 980 2504
rect 974 2499 975 2503
rect 979 2499 980 2503
rect 974 2498 980 2499
rect 1054 2503 1060 2504
rect 1054 2499 1055 2503
rect 1059 2499 1060 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1328 2499 1330 2510
rect 1382 2508 1383 2512
rect 1387 2508 1388 2512
rect 1382 2507 1388 2508
rect 1438 2512 1444 2513
rect 1438 2508 1439 2512
rect 1443 2508 1444 2512
rect 1438 2507 1444 2508
rect 1494 2512 1500 2513
rect 1494 2508 1495 2512
rect 1499 2508 1500 2512
rect 1494 2507 1500 2508
rect 1550 2512 1556 2513
rect 1550 2508 1551 2512
rect 1555 2508 1556 2512
rect 1550 2507 1556 2508
rect 1606 2512 1612 2513
rect 1606 2508 1607 2512
rect 1611 2508 1612 2512
rect 1606 2507 1612 2508
rect 1662 2512 1668 2513
rect 1662 2508 1663 2512
rect 1667 2508 1668 2512
rect 1662 2507 1668 2508
rect 1718 2512 1724 2513
rect 1718 2508 1719 2512
rect 1723 2508 1724 2512
rect 1718 2507 1724 2508
rect 1774 2512 1780 2513
rect 1774 2508 1775 2512
rect 1779 2508 1780 2512
rect 1774 2507 1780 2508
rect 1830 2512 1836 2513
rect 1830 2508 1831 2512
rect 1835 2508 1836 2512
rect 1830 2507 1836 2508
rect 1886 2512 1892 2513
rect 1886 2508 1887 2512
rect 1891 2508 1892 2512
rect 1886 2507 1892 2508
rect 1942 2512 1948 2513
rect 1942 2508 1943 2512
rect 1947 2508 1948 2512
rect 1942 2507 1948 2508
rect 1998 2512 2004 2513
rect 1998 2508 1999 2512
rect 2003 2508 2004 2512
rect 1998 2507 2004 2508
rect 2054 2512 2060 2513
rect 2054 2508 2055 2512
rect 2059 2508 2060 2512
rect 2054 2507 2060 2508
rect 2110 2512 2116 2513
rect 2110 2508 2111 2512
rect 2115 2508 2116 2512
rect 2110 2507 2116 2508
rect 2166 2512 2172 2513
rect 2166 2508 2167 2512
rect 2171 2508 2172 2512
rect 2502 2511 2503 2515
rect 2507 2511 2508 2515
rect 2502 2510 2508 2511
rect 2166 2507 2172 2508
rect 1384 2499 1386 2507
rect 1440 2499 1442 2507
rect 1496 2499 1498 2507
rect 1552 2499 1554 2507
rect 1608 2499 1610 2507
rect 1664 2499 1666 2507
rect 1720 2499 1722 2507
rect 1776 2499 1778 2507
rect 1832 2499 1834 2507
rect 1888 2499 1890 2507
rect 1944 2499 1946 2507
rect 2000 2499 2002 2507
rect 2056 2499 2058 2507
rect 2112 2499 2114 2507
rect 2168 2499 2170 2507
rect 2504 2499 2506 2510
rect 1054 2498 1060 2499
rect 184 2479 186 2498
rect 240 2479 242 2498
rect 296 2479 298 2498
rect 360 2479 362 2498
rect 424 2479 426 2498
rect 496 2479 498 2498
rect 576 2479 578 2498
rect 656 2479 658 2498
rect 736 2479 738 2498
rect 816 2479 818 2498
rect 896 2479 898 2498
rect 976 2479 978 2498
rect 1056 2479 1058 2498
rect 1288 2479 1290 2499
rect 1327 2498 1331 2499
rect 1327 2493 1331 2494
rect 1351 2498 1355 2499
rect 1351 2493 1355 2494
rect 1383 2498 1387 2499
rect 1383 2493 1387 2494
rect 1423 2498 1427 2499
rect 1423 2493 1427 2494
rect 1439 2498 1443 2499
rect 1439 2493 1443 2494
rect 1495 2498 1499 2499
rect 1495 2493 1499 2494
rect 1511 2498 1515 2499
rect 1511 2493 1515 2494
rect 1551 2498 1555 2499
rect 1551 2493 1555 2494
rect 1599 2498 1603 2499
rect 1599 2493 1603 2494
rect 1607 2498 1611 2499
rect 1607 2493 1611 2494
rect 1663 2498 1667 2499
rect 1663 2493 1667 2494
rect 1687 2498 1691 2499
rect 1687 2493 1691 2494
rect 1719 2498 1723 2499
rect 1719 2493 1723 2494
rect 1775 2498 1779 2499
rect 1775 2493 1779 2494
rect 1831 2498 1835 2499
rect 1831 2493 1835 2494
rect 1863 2498 1867 2499
rect 1863 2493 1867 2494
rect 1887 2498 1891 2499
rect 1887 2493 1891 2494
rect 1943 2498 1947 2499
rect 1943 2493 1947 2494
rect 1951 2498 1955 2499
rect 1951 2493 1955 2494
rect 1999 2498 2003 2499
rect 1999 2493 2003 2494
rect 2039 2498 2043 2499
rect 2039 2493 2043 2494
rect 2055 2498 2059 2499
rect 2055 2493 2059 2494
rect 2111 2498 2115 2499
rect 2111 2493 2115 2494
rect 2127 2498 2131 2499
rect 2127 2493 2131 2494
rect 2167 2498 2171 2499
rect 2167 2493 2171 2494
rect 2503 2498 2507 2499
rect 2503 2493 2507 2494
rect 1328 2490 1330 2493
rect 1350 2492 1356 2493
rect 1326 2489 1332 2490
rect 1326 2485 1327 2489
rect 1331 2485 1332 2489
rect 1350 2488 1351 2492
rect 1355 2488 1356 2492
rect 1350 2487 1356 2488
rect 1422 2492 1428 2493
rect 1422 2488 1423 2492
rect 1427 2488 1428 2492
rect 1422 2487 1428 2488
rect 1510 2492 1516 2493
rect 1510 2488 1511 2492
rect 1515 2488 1516 2492
rect 1510 2487 1516 2488
rect 1598 2492 1604 2493
rect 1598 2488 1599 2492
rect 1603 2488 1604 2492
rect 1598 2487 1604 2488
rect 1686 2492 1692 2493
rect 1686 2488 1687 2492
rect 1691 2488 1692 2492
rect 1686 2487 1692 2488
rect 1774 2492 1780 2493
rect 1774 2488 1775 2492
rect 1779 2488 1780 2492
rect 1774 2487 1780 2488
rect 1862 2492 1868 2493
rect 1862 2488 1863 2492
rect 1867 2488 1868 2492
rect 1862 2487 1868 2488
rect 1950 2492 1956 2493
rect 1950 2488 1951 2492
rect 1955 2488 1956 2492
rect 1950 2487 1956 2488
rect 2038 2492 2044 2493
rect 2038 2488 2039 2492
rect 2043 2488 2044 2492
rect 2038 2487 2044 2488
rect 2126 2492 2132 2493
rect 2126 2488 2127 2492
rect 2131 2488 2132 2492
rect 2504 2490 2506 2493
rect 2126 2487 2132 2488
rect 2502 2489 2508 2490
rect 1326 2484 1332 2485
rect 2502 2485 2503 2489
rect 2507 2485 2508 2489
rect 2502 2484 2508 2485
rect 111 2478 115 2479
rect 111 2473 115 2474
rect 183 2478 187 2479
rect 183 2473 187 2474
rect 239 2478 243 2479
rect 239 2473 243 2474
rect 247 2478 251 2479
rect 247 2473 251 2474
rect 295 2478 299 2479
rect 295 2473 299 2474
rect 327 2478 331 2479
rect 327 2473 331 2474
rect 359 2478 363 2479
rect 359 2473 363 2474
rect 415 2478 419 2479
rect 415 2473 419 2474
rect 423 2478 427 2479
rect 423 2473 427 2474
rect 495 2478 499 2479
rect 495 2473 499 2474
rect 503 2478 507 2479
rect 503 2473 507 2474
rect 575 2478 579 2479
rect 575 2473 579 2474
rect 599 2478 603 2479
rect 599 2473 603 2474
rect 655 2478 659 2479
rect 655 2473 659 2474
rect 695 2478 699 2479
rect 695 2473 699 2474
rect 735 2478 739 2479
rect 735 2473 739 2474
rect 791 2478 795 2479
rect 791 2473 795 2474
rect 815 2478 819 2479
rect 815 2473 819 2474
rect 879 2478 883 2479
rect 879 2473 883 2474
rect 895 2478 899 2479
rect 895 2473 899 2474
rect 967 2478 971 2479
rect 967 2473 971 2474
rect 975 2478 979 2479
rect 975 2473 979 2474
rect 1055 2478 1059 2479
rect 1055 2473 1059 2474
rect 1063 2478 1067 2479
rect 1063 2473 1067 2474
rect 1159 2478 1163 2479
rect 1159 2473 1163 2474
rect 1287 2478 1291 2479
rect 1287 2473 1291 2474
rect 112 2453 114 2473
rect 184 2454 186 2473
rect 248 2454 250 2473
rect 328 2454 330 2473
rect 416 2454 418 2473
rect 504 2454 506 2473
rect 600 2454 602 2473
rect 696 2454 698 2473
rect 792 2454 794 2473
rect 880 2454 882 2473
rect 968 2454 970 2473
rect 1064 2454 1066 2473
rect 1160 2454 1162 2473
rect 182 2453 188 2454
rect 110 2452 116 2453
rect 110 2448 111 2452
rect 115 2448 116 2452
rect 182 2449 183 2453
rect 187 2449 188 2453
rect 182 2448 188 2449
rect 246 2453 252 2454
rect 246 2449 247 2453
rect 251 2449 252 2453
rect 246 2448 252 2449
rect 326 2453 332 2454
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 414 2453 420 2454
rect 414 2449 415 2453
rect 419 2449 420 2453
rect 414 2448 420 2449
rect 502 2453 508 2454
rect 502 2449 503 2453
rect 507 2449 508 2453
rect 502 2448 508 2449
rect 598 2453 604 2454
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 598 2448 604 2449
rect 694 2453 700 2454
rect 694 2449 695 2453
rect 699 2449 700 2453
rect 694 2448 700 2449
rect 790 2453 796 2454
rect 790 2449 791 2453
rect 795 2449 796 2453
rect 790 2448 796 2449
rect 878 2453 884 2454
rect 878 2449 879 2453
rect 883 2449 884 2453
rect 878 2448 884 2449
rect 966 2453 972 2454
rect 966 2449 967 2453
rect 971 2449 972 2453
rect 966 2448 972 2449
rect 1062 2453 1068 2454
rect 1062 2449 1063 2453
rect 1067 2449 1068 2453
rect 1062 2448 1068 2449
rect 1158 2453 1164 2454
rect 1288 2453 1290 2473
rect 1326 2472 1332 2473
rect 2502 2472 2508 2473
rect 1326 2468 1327 2472
rect 1331 2468 1332 2472
rect 1326 2467 1332 2468
rect 1366 2471 1372 2472
rect 1366 2467 1367 2471
rect 1371 2467 1372 2471
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1158 2448 1164 2449
rect 1286 2452 1292 2453
rect 1286 2448 1287 2452
rect 1291 2448 1292 2452
rect 110 2447 116 2448
rect 1286 2447 1292 2448
rect 1328 2439 1330 2467
rect 1366 2466 1372 2467
rect 1438 2471 1444 2472
rect 1438 2467 1439 2471
rect 1443 2467 1444 2471
rect 1438 2466 1444 2467
rect 1526 2471 1532 2472
rect 1526 2467 1527 2471
rect 1531 2467 1532 2471
rect 1526 2466 1532 2467
rect 1614 2471 1620 2472
rect 1614 2467 1615 2471
rect 1619 2467 1620 2471
rect 1614 2466 1620 2467
rect 1702 2471 1708 2472
rect 1702 2467 1703 2471
rect 1707 2467 1708 2471
rect 1702 2466 1708 2467
rect 1790 2471 1796 2472
rect 1790 2467 1791 2471
rect 1795 2467 1796 2471
rect 1790 2466 1796 2467
rect 1878 2471 1884 2472
rect 1878 2467 1879 2471
rect 1883 2467 1884 2471
rect 1878 2466 1884 2467
rect 1966 2471 1972 2472
rect 1966 2467 1967 2471
rect 1971 2467 1972 2471
rect 1966 2466 1972 2467
rect 2054 2471 2060 2472
rect 2054 2467 2055 2471
rect 2059 2467 2060 2471
rect 2054 2466 2060 2467
rect 2142 2471 2148 2472
rect 2142 2467 2143 2471
rect 2147 2467 2148 2471
rect 2502 2468 2503 2472
rect 2507 2468 2508 2472
rect 2502 2467 2508 2468
rect 2142 2466 2148 2467
rect 1368 2439 1370 2466
rect 1440 2439 1442 2466
rect 1528 2439 1530 2466
rect 1616 2439 1618 2466
rect 1704 2439 1706 2466
rect 1792 2439 1794 2466
rect 1880 2439 1882 2466
rect 1968 2439 1970 2466
rect 2056 2439 2058 2466
rect 2144 2439 2146 2466
rect 2504 2439 2506 2467
rect 1327 2438 1331 2439
rect 110 2435 116 2436
rect 110 2431 111 2435
rect 115 2431 116 2435
rect 1286 2435 1292 2436
rect 110 2430 116 2431
rect 166 2432 172 2433
rect 112 2423 114 2430
rect 166 2428 167 2432
rect 171 2428 172 2432
rect 166 2427 172 2428
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 486 2432 492 2433
rect 486 2428 487 2432
rect 491 2428 492 2432
rect 486 2427 492 2428
rect 582 2432 588 2433
rect 582 2428 583 2432
rect 587 2428 588 2432
rect 582 2427 588 2428
rect 678 2432 684 2433
rect 678 2428 679 2432
rect 683 2428 684 2432
rect 678 2427 684 2428
rect 774 2432 780 2433
rect 774 2428 775 2432
rect 779 2428 780 2432
rect 774 2427 780 2428
rect 862 2432 868 2433
rect 862 2428 863 2432
rect 867 2428 868 2432
rect 862 2427 868 2428
rect 950 2432 956 2433
rect 950 2428 951 2432
rect 955 2428 956 2432
rect 950 2427 956 2428
rect 1046 2432 1052 2433
rect 1046 2428 1047 2432
rect 1051 2428 1052 2432
rect 1046 2427 1052 2428
rect 1142 2432 1148 2433
rect 1142 2428 1143 2432
rect 1147 2428 1148 2432
rect 1286 2431 1287 2435
rect 1291 2431 1292 2435
rect 1327 2433 1331 2434
rect 1367 2438 1371 2439
rect 1367 2433 1371 2434
rect 1439 2438 1443 2439
rect 1439 2433 1443 2434
rect 1527 2438 1531 2439
rect 1527 2433 1531 2434
rect 1543 2438 1547 2439
rect 1543 2433 1547 2434
rect 1615 2438 1619 2439
rect 1615 2433 1619 2434
rect 1639 2438 1643 2439
rect 1639 2433 1643 2434
rect 1703 2438 1707 2439
rect 1703 2433 1707 2434
rect 1735 2438 1739 2439
rect 1735 2433 1739 2434
rect 1791 2438 1795 2439
rect 1791 2433 1795 2434
rect 1823 2438 1827 2439
rect 1823 2433 1827 2434
rect 1879 2438 1883 2439
rect 1879 2433 1883 2434
rect 1911 2438 1915 2439
rect 1911 2433 1915 2434
rect 1967 2438 1971 2439
rect 1967 2433 1971 2434
rect 2007 2438 2011 2439
rect 2007 2433 2011 2434
rect 2055 2438 2059 2439
rect 2055 2433 2059 2434
rect 2103 2438 2107 2439
rect 2103 2433 2107 2434
rect 2143 2438 2147 2439
rect 2143 2433 2147 2434
rect 2503 2438 2507 2439
rect 2503 2433 2507 2434
rect 1286 2430 1292 2431
rect 1142 2427 1148 2428
rect 168 2423 170 2427
rect 232 2423 234 2427
rect 312 2423 314 2427
rect 400 2423 402 2427
rect 488 2423 490 2427
rect 584 2423 586 2427
rect 680 2423 682 2427
rect 776 2423 778 2427
rect 864 2423 866 2427
rect 952 2423 954 2427
rect 1048 2423 1050 2427
rect 1144 2423 1146 2427
rect 1288 2423 1290 2430
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 151 2422 155 2423
rect 151 2417 155 2418
rect 167 2422 171 2423
rect 167 2417 171 2418
rect 231 2422 235 2423
rect 231 2417 235 2418
rect 311 2422 315 2423
rect 311 2417 315 2418
rect 319 2422 323 2423
rect 319 2417 323 2418
rect 399 2422 403 2423
rect 399 2417 403 2418
rect 415 2422 419 2423
rect 415 2417 419 2418
rect 487 2422 491 2423
rect 487 2417 491 2418
rect 519 2422 523 2423
rect 519 2417 523 2418
rect 583 2422 587 2423
rect 583 2417 587 2418
rect 623 2422 627 2423
rect 623 2417 627 2418
rect 679 2422 683 2423
rect 679 2417 683 2418
rect 727 2422 731 2423
rect 727 2417 731 2418
rect 775 2422 779 2423
rect 775 2417 779 2418
rect 831 2422 835 2423
rect 831 2417 835 2418
rect 863 2422 867 2423
rect 863 2417 867 2418
rect 935 2422 939 2423
rect 935 2417 939 2418
rect 951 2422 955 2423
rect 951 2417 955 2418
rect 1039 2422 1043 2423
rect 1039 2417 1043 2418
rect 1047 2422 1051 2423
rect 1047 2417 1051 2418
rect 1143 2422 1147 2423
rect 1143 2417 1147 2418
rect 1151 2422 1155 2423
rect 1151 2417 1155 2418
rect 1287 2422 1291 2423
rect 1287 2417 1291 2418
rect 112 2414 114 2417
rect 150 2416 156 2417
rect 110 2413 116 2414
rect 110 2409 111 2413
rect 115 2409 116 2413
rect 150 2412 151 2416
rect 155 2412 156 2416
rect 150 2411 156 2412
rect 230 2416 236 2417
rect 230 2412 231 2416
rect 235 2412 236 2416
rect 230 2411 236 2412
rect 318 2416 324 2417
rect 318 2412 319 2416
rect 323 2412 324 2416
rect 318 2411 324 2412
rect 414 2416 420 2417
rect 414 2412 415 2416
rect 419 2412 420 2416
rect 414 2411 420 2412
rect 518 2416 524 2417
rect 518 2412 519 2416
rect 523 2412 524 2416
rect 518 2411 524 2412
rect 622 2416 628 2417
rect 622 2412 623 2416
rect 627 2412 628 2416
rect 622 2411 628 2412
rect 726 2416 732 2417
rect 726 2412 727 2416
rect 731 2412 732 2416
rect 726 2411 732 2412
rect 830 2416 836 2417
rect 830 2412 831 2416
rect 835 2412 836 2416
rect 830 2411 836 2412
rect 934 2416 940 2417
rect 934 2412 935 2416
rect 939 2412 940 2416
rect 934 2411 940 2412
rect 1038 2416 1044 2417
rect 1038 2412 1039 2416
rect 1043 2412 1044 2416
rect 1038 2411 1044 2412
rect 1150 2416 1156 2417
rect 1150 2412 1151 2416
rect 1155 2412 1156 2416
rect 1288 2414 1290 2417
rect 1150 2411 1156 2412
rect 1286 2413 1292 2414
rect 1328 2413 1330 2433
rect 1368 2414 1370 2433
rect 1440 2414 1442 2433
rect 1544 2414 1546 2433
rect 1640 2414 1642 2433
rect 1736 2414 1738 2433
rect 1824 2414 1826 2433
rect 1912 2414 1914 2433
rect 2008 2414 2010 2433
rect 2104 2414 2106 2433
rect 1366 2413 1372 2414
rect 110 2408 116 2409
rect 1286 2409 1287 2413
rect 1291 2409 1292 2413
rect 1286 2408 1292 2409
rect 1326 2412 1332 2413
rect 1326 2408 1327 2412
rect 1331 2408 1332 2412
rect 1366 2409 1367 2413
rect 1371 2409 1372 2413
rect 1366 2408 1372 2409
rect 1438 2413 1444 2414
rect 1438 2409 1439 2413
rect 1443 2409 1444 2413
rect 1438 2408 1444 2409
rect 1542 2413 1548 2414
rect 1542 2409 1543 2413
rect 1547 2409 1548 2413
rect 1542 2408 1548 2409
rect 1638 2413 1644 2414
rect 1638 2409 1639 2413
rect 1643 2409 1644 2413
rect 1638 2408 1644 2409
rect 1734 2413 1740 2414
rect 1734 2409 1735 2413
rect 1739 2409 1740 2413
rect 1734 2408 1740 2409
rect 1822 2413 1828 2414
rect 1822 2409 1823 2413
rect 1827 2409 1828 2413
rect 1822 2408 1828 2409
rect 1910 2413 1916 2414
rect 1910 2409 1911 2413
rect 1915 2409 1916 2413
rect 1910 2408 1916 2409
rect 2006 2413 2012 2414
rect 2006 2409 2007 2413
rect 2011 2409 2012 2413
rect 2006 2408 2012 2409
rect 2102 2413 2108 2414
rect 2504 2413 2506 2433
rect 2102 2409 2103 2413
rect 2107 2409 2108 2413
rect 2102 2408 2108 2409
rect 2502 2412 2508 2413
rect 2502 2408 2503 2412
rect 2507 2408 2508 2412
rect 1326 2407 1332 2408
rect 2502 2407 2508 2408
rect 110 2396 116 2397
rect 1286 2396 1292 2397
rect 110 2392 111 2396
rect 115 2392 116 2396
rect 110 2391 116 2392
rect 166 2395 172 2396
rect 166 2391 167 2395
rect 171 2391 172 2395
rect 112 2371 114 2391
rect 166 2390 172 2391
rect 246 2395 252 2396
rect 246 2391 247 2395
rect 251 2391 252 2395
rect 246 2390 252 2391
rect 334 2395 340 2396
rect 334 2391 335 2395
rect 339 2391 340 2395
rect 334 2390 340 2391
rect 430 2395 436 2396
rect 430 2391 431 2395
rect 435 2391 436 2395
rect 430 2390 436 2391
rect 534 2395 540 2396
rect 534 2391 535 2395
rect 539 2391 540 2395
rect 534 2390 540 2391
rect 638 2395 644 2396
rect 638 2391 639 2395
rect 643 2391 644 2395
rect 638 2390 644 2391
rect 742 2395 748 2396
rect 742 2391 743 2395
rect 747 2391 748 2395
rect 742 2390 748 2391
rect 846 2395 852 2396
rect 846 2391 847 2395
rect 851 2391 852 2395
rect 846 2390 852 2391
rect 950 2395 956 2396
rect 950 2391 951 2395
rect 955 2391 956 2395
rect 950 2390 956 2391
rect 1054 2395 1060 2396
rect 1054 2391 1055 2395
rect 1059 2391 1060 2395
rect 1054 2390 1060 2391
rect 1166 2395 1172 2396
rect 1166 2391 1167 2395
rect 1171 2391 1172 2395
rect 1286 2392 1287 2396
rect 1291 2392 1292 2396
rect 1286 2391 1292 2392
rect 1326 2395 1332 2396
rect 1326 2391 1327 2395
rect 1331 2391 1332 2395
rect 2502 2395 2508 2396
rect 1166 2390 1172 2391
rect 168 2371 170 2390
rect 248 2371 250 2390
rect 336 2371 338 2390
rect 432 2371 434 2390
rect 536 2371 538 2390
rect 640 2371 642 2390
rect 744 2371 746 2390
rect 848 2371 850 2390
rect 952 2371 954 2390
rect 1056 2371 1058 2390
rect 1168 2371 1170 2390
rect 1288 2371 1290 2391
rect 1326 2390 1332 2391
rect 1350 2392 1356 2393
rect 1328 2379 1330 2390
rect 1350 2388 1351 2392
rect 1355 2388 1356 2392
rect 1350 2387 1356 2388
rect 1422 2392 1428 2393
rect 1422 2388 1423 2392
rect 1427 2388 1428 2392
rect 1422 2387 1428 2388
rect 1526 2392 1532 2393
rect 1526 2388 1527 2392
rect 1531 2388 1532 2392
rect 1526 2387 1532 2388
rect 1622 2392 1628 2393
rect 1622 2388 1623 2392
rect 1627 2388 1628 2392
rect 1622 2387 1628 2388
rect 1718 2392 1724 2393
rect 1718 2388 1719 2392
rect 1723 2388 1724 2392
rect 1718 2387 1724 2388
rect 1806 2392 1812 2393
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1894 2392 1900 2393
rect 1894 2388 1895 2392
rect 1899 2388 1900 2392
rect 1894 2387 1900 2388
rect 1990 2392 1996 2393
rect 1990 2388 1991 2392
rect 1995 2388 1996 2392
rect 1990 2387 1996 2388
rect 2086 2392 2092 2393
rect 2086 2388 2087 2392
rect 2091 2388 2092 2392
rect 2502 2391 2503 2395
rect 2507 2391 2508 2395
rect 2502 2390 2508 2391
rect 2086 2387 2092 2388
rect 1352 2379 1354 2387
rect 1424 2379 1426 2387
rect 1528 2379 1530 2387
rect 1624 2379 1626 2387
rect 1720 2379 1722 2387
rect 1808 2379 1810 2387
rect 1896 2379 1898 2387
rect 1992 2379 1994 2387
rect 2088 2379 2090 2387
rect 2504 2379 2506 2390
rect 1327 2378 1331 2379
rect 1327 2373 1331 2374
rect 1351 2378 1355 2379
rect 1351 2373 1355 2374
rect 1407 2378 1411 2379
rect 1407 2373 1411 2374
rect 1423 2378 1427 2379
rect 1423 2373 1427 2374
rect 1495 2378 1499 2379
rect 1495 2373 1499 2374
rect 1527 2378 1531 2379
rect 1527 2373 1531 2374
rect 1583 2378 1587 2379
rect 1583 2373 1587 2374
rect 1623 2378 1627 2379
rect 1623 2373 1627 2374
rect 1671 2378 1675 2379
rect 1671 2373 1675 2374
rect 1719 2378 1723 2379
rect 1719 2373 1723 2374
rect 1751 2378 1755 2379
rect 1751 2373 1755 2374
rect 1807 2378 1811 2379
rect 1807 2373 1811 2374
rect 1831 2378 1835 2379
rect 1831 2373 1835 2374
rect 1895 2378 1899 2379
rect 1895 2373 1899 2374
rect 1919 2378 1923 2379
rect 1919 2373 1923 2374
rect 1991 2378 1995 2379
rect 1991 2373 1995 2374
rect 2007 2378 2011 2379
rect 2007 2373 2011 2374
rect 2087 2378 2091 2379
rect 2087 2373 2091 2374
rect 2095 2378 2099 2379
rect 2095 2373 2099 2374
rect 2503 2378 2507 2379
rect 2503 2373 2507 2374
rect 111 2370 115 2371
rect 111 2365 115 2366
rect 167 2370 171 2371
rect 167 2365 171 2366
rect 175 2370 179 2371
rect 175 2365 179 2366
rect 247 2370 251 2371
rect 247 2365 251 2366
rect 279 2370 283 2371
rect 279 2365 283 2366
rect 335 2370 339 2371
rect 335 2365 339 2366
rect 391 2370 395 2371
rect 391 2365 395 2366
rect 431 2370 435 2371
rect 431 2365 435 2366
rect 503 2370 507 2371
rect 503 2365 507 2366
rect 535 2370 539 2371
rect 535 2365 539 2366
rect 623 2370 627 2371
rect 623 2365 627 2366
rect 639 2370 643 2371
rect 639 2365 643 2366
rect 743 2370 747 2371
rect 743 2365 747 2366
rect 847 2370 851 2371
rect 847 2365 851 2366
rect 871 2370 875 2371
rect 871 2365 875 2366
rect 951 2370 955 2371
rect 951 2365 955 2366
rect 999 2370 1003 2371
rect 999 2365 1003 2366
rect 1055 2370 1059 2371
rect 1055 2365 1059 2366
rect 1127 2370 1131 2371
rect 1127 2365 1131 2366
rect 1167 2370 1171 2371
rect 1167 2365 1171 2366
rect 1287 2370 1291 2371
rect 1328 2370 1330 2373
rect 1350 2372 1356 2373
rect 1287 2365 1291 2366
rect 1326 2369 1332 2370
rect 1326 2365 1327 2369
rect 1331 2365 1332 2369
rect 1350 2368 1351 2372
rect 1355 2368 1356 2372
rect 1350 2367 1356 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1494 2372 1500 2373
rect 1494 2368 1495 2372
rect 1499 2368 1500 2372
rect 1494 2367 1500 2368
rect 1582 2372 1588 2373
rect 1582 2368 1583 2372
rect 1587 2368 1588 2372
rect 1582 2367 1588 2368
rect 1670 2372 1676 2373
rect 1670 2368 1671 2372
rect 1675 2368 1676 2372
rect 1670 2367 1676 2368
rect 1750 2372 1756 2373
rect 1750 2368 1751 2372
rect 1755 2368 1756 2372
rect 1750 2367 1756 2368
rect 1830 2372 1836 2373
rect 1830 2368 1831 2372
rect 1835 2368 1836 2372
rect 1830 2367 1836 2368
rect 1918 2372 1924 2373
rect 1918 2368 1919 2372
rect 1923 2368 1924 2372
rect 1918 2367 1924 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2094 2372 2100 2373
rect 2094 2368 2095 2372
rect 2099 2368 2100 2372
rect 2504 2370 2506 2373
rect 2094 2367 2100 2368
rect 2502 2369 2508 2370
rect 112 2345 114 2365
rect 176 2346 178 2365
rect 280 2346 282 2365
rect 392 2346 394 2365
rect 504 2346 506 2365
rect 624 2346 626 2365
rect 744 2346 746 2365
rect 872 2346 874 2365
rect 1000 2346 1002 2365
rect 1128 2346 1130 2365
rect 174 2345 180 2346
rect 110 2344 116 2345
rect 110 2340 111 2344
rect 115 2340 116 2344
rect 174 2341 175 2345
rect 179 2341 180 2345
rect 174 2340 180 2341
rect 278 2345 284 2346
rect 278 2341 279 2345
rect 283 2341 284 2345
rect 278 2340 284 2341
rect 390 2345 396 2346
rect 390 2341 391 2345
rect 395 2341 396 2345
rect 390 2340 396 2341
rect 502 2345 508 2346
rect 502 2341 503 2345
rect 507 2341 508 2345
rect 502 2340 508 2341
rect 622 2345 628 2346
rect 622 2341 623 2345
rect 627 2341 628 2345
rect 622 2340 628 2341
rect 742 2345 748 2346
rect 742 2341 743 2345
rect 747 2341 748 2345
rect 742 2340 748 2341
rect 870 2345 876 2346
rect 870 2341 871 2345
rect 875 2341 876 2345
rect 870 2340 876 2341
rect 998 2345 1004 2346
rect 998 2341 999 2345
rect 1003 2341 1004 2345
rect 998 2340 1004 2341
rect 1126 2345 1132 2346
rect 1288 2345 1290 2365
rect 1326 2364 1332 2365
rect 2502 2365 2503 2369
rect 2507 2365 2508 2369
rect 2502 2364 2508 2365
rect 1326 2352 1332 2353
rect 2502 2352 2508 2353
rect 1326 2348 1327 2352
rect 1331 2348 1332 2352
rect 1326 2347 1332 2348
rect 1366 2351 1372 2352
rect 1366 2347 1367 2351
rect 1371 2347 1372 2351
rect 1126 2341 1127 2345
rect 1131 2341 1132 2345
rect 1126 2340 1132 2341
rect 1286 2344 1292 2345
rect 1286 2340 1287 2344
rect 1291 2340 1292 2344
rect 110 2339 116 2340
rect 1286 2339 1292 2340
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 1286 2327 1292 2328
rect 110 2322 116 2323
rect 158 2324 164 2325
rect 112 2315 114 2322
rect 158 2320 159 2324
rect 163 2320 164 2324
rect 158 2319 164 2320
rect 262 2324 268 2325
rect 262 2320 263 2324
rect 267 2320 268 2324
rect 262 2319 268 2320
rect 374 2324 380 2325
rect 374 2320 375 2324
rect 379 2320 380 2324
rect 374 2319 380 2320
rect 486 2324 492 2325
rect 486 2320 487 2324
rect 491 2320 492 2324
rect 486 2319 492 2320
rect 606 2324 612 2325
rect 606 2320 607 2324
rect 611 2320 612 2324
rect 606 2319 612 2320
rect 726 2324 732 2325
rect 726 2320 727 2324
rect 731 2320 732 2324
rect 726 2319 732 2320
rect 854 2324 860 2325
rect 854 2320 855 2324
rect 859 2320 860 2324
rect 854 2319 860 2320
rect 982 2324 988 2325
rect 982 2320 983 2324
rect 987 2320 988 2324
rect 982 2319 988 2320
rect 1110 2324 1116 2325
rect 1110 2320 1111 2324
rect 1115 2320 1116 2324
rect 1286 2323 1287 2327
rect 1291 2323 1292 2327
rect 1328 2323 1330 2347
rect 1366 2346 1372 2347
rect 1422 2351 1428 2352
rect 1422 2347 1423 2351
rect 1427 2347 1428 2351
rect 1422 2346 1428 2347
rect 1510 2351 1516 2352
rect 1510 2347 1511 2351
rect 1515 2347 1516 2351
rect 1510 2346 1516 2347
rect 1598 2351 1604 2352
rect 1598 2347 1599 2351
rect 1603 2347 1604 2351
rect 1598 2346 1604 2347
rect 1686 2351 1692 2352
rect 1686 2347 1687 2351
rect 1691 2347 1692 2351
rect 1686 2346 1692 2347
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2347 1772 2351
rect 1766 2346 1772 2347
rect 1846 2351 1852 2352
rect 1846 2347 1847 2351
rect 1851 2347 1852 2351
rect 1846 2346 1852 2347
rect 1934 2351 1940 2352
rect 1934 2347 1935 2351
rect 1939 2347 1940 2351
rect 1934 2346 1940 2347
rect 2022 2351 2028 2352
rect 2022 2347 2023 2351
rect 2027 2347 2028 2351
rect 2022 2346 2028 2347
rect 2110 2351 2116 2352
rect 2110 2347 2111 2351
rect 2115 2347 2116 2351
rect 2502 2348 2503 2352
rect 2507 2348 2508 2352
rect 2502 2347 2508 2348
rect 2110 2346 2116 2347
rect 1368 2323 1370 2346
rect 1424 2323 1426 2346
rect 1512 2323 1514 2346
rect 1600 2323 1602 2346
rect 1688 2323 1690 2346
rect 1768 2323 1770 2346
rect 1848 2323 1850 2346
rect 1936 2323 1938 2346
rect 2024 2323 2026 2346
rect 2112 2323 2114 2346
rect 2504 2323 2506 2347
rect 1286 2322 1292 2323
rect 1327 2322 1331 2323
rect 1110 2319 1116 2320
rect 160 2315 162 2319
rect 264 2315 266 2319
rect 376 2315 378 2319
rect 488 2315 490 2319
rect 608 2315 610 2319
rect 728 2315 730 2319
rect 856 2315 858 2319
rect 984 2315 986 2319
rect 1112 2315 1114 2319
rect 1288 2315 1290 2322
rect 1327 2317 1331 2318
rect 1367 2322 1371 2323
rect 1367 2317 1371 2318
rect 1423 2322 1427 2323
rect 1423 2317 1427 2318
rect 1455 2322 1459 2323
rect 1455 2317 1459 2318
rect 1511 2322 1515 2323
rect 1511 2317 1515 2318
rect 1543 2322 1547 2323
rect 1543 2317 1547 2318
rect 1599 2322 1603 2323
rect 1599 2317 1603 2318
rect 1639 2322 1643 2323
rect 1639 2317 1643 2318
rect 1687 2322 1691 2323
rect 1687 2317 1691 2318
rect 1735 2322 1739 2323
rect 1735 2317 1739 2318
rect 1767 2322 1771 2323
rect 1767 2317 1771 2318
rect 1831 2322 1835 2323
rect 1831 2317 1835 2318
rect 1847 2322 1851 2323
rect 1847 2317 1851 2318
rect 1927 2322 1931 2323
rect 1927 2317 1931 2318
rect 1935 2322 1939 2323
rect 1935 2317 1939 2318
rect 2015 2322 2019 2323
rect 2015 2317 2019 2318
rect 2023 2322 2027 2323
rect 2023 2317 2027 2318
rect 2111 2322 2115 2323
rect 2111 2317 2115 2318
rect 2207 2322 2211 2323
rect 2207 2317 2211 2318
rect 2503 2322 2507 2323
rect 2503 2317 2507 2318
rect 111 2314 115 2315
rect 111 2309 115 2310
rect 159 2314 163 2315
rect 159 2309 163 2310
rect 207 2314 211 2315
rect 207 2309 211 2310
rect 263 2314 267 2315
rect 263 2309 267 2310
rect 287 2314 291 2315
rect 287 2309 291 2310
rect 375 2314 379 2315
rect 375 2309 379 2310
rect 471 2314 475 2315
rect 471 2309 475 2310
rect 487 2314 491 2315
rect 487 2309 491 2310
rect 559 2314 563 2315
rect 559 2309 563 2310
rect 607 2314 611 2315
rect 607 2309 611 2310
rect 647 2314 651 2315
rect 647 2309 651 2310
rect 727 2314 731 2315
rect 727 2309 731 2310
rect 735 2314 739 2315
rect 735 2309 739 2310
rect 815 2314 819 2315
rect 815 2309 819 2310
rect 855 2314 859 2315
rect 855 2309 859 2310
rect 903 2314 907 2315
rect 903 2309 907 2310
rect 983 2314 987 2315
rect 983 2309 987 2310
rect 991 2314 995 2315
rect 991 2309 995 2310
rect 1079 2314 1083 2315
rect 1079 2309 1083 2310
rect 1111 2314 1115 2315
rect 1111 2309 1115 2310
rect 1287 2314 1291 2315
rect 1287 2309 1291 2310
rect 112 2306 114 2309
rect 206 2308 212 2309
rect 110 2305 116 2306
rect 110 2301 111 2305
rect 115 2301 116 2305
rect 206 2304 207 2308
rect 211 2304 212 2308
rect 206 2303 212 2304
rect 286 2308 292 2309
rect 286 2304 287 2308
rect 291 2304 292 2308
rect 286 2303 292 2304
rect 374 2308 380 2309
rect 374 2304 375 2308
rect 379 2304 380 2308
rect 374 2303 380 2304
rect 470 2308 476 2309
rect 470 2304 471 2308
rect 475 2304 476 2308
rect 470 2303 476 2304
rect 558 2308 564 2309
rect 558 2304 559 2308
rect 563 2304 564 2308
rect 558 2303 564 2304
rect 646 2308 652 2309
rect 646 2304 647 2308
rect 651 2304 652 2308
rect 646 2303 652 2304
rect 734 2308 740 2309
rect 734 2304 735 2308
rect 739 2304 740 2308
rect 734 2303 740 2304
rect 814 2308 820 2309
rect 814 2304 815 2308
rect 819 2304 820 2308
rect 814 2303 820 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 990 2308 996 2309
rect 990 2304 991 2308
rect 995 2304 996 2308
rect 990 2303 996 2304
rect 1078 2308 1084 2309
rect 1078 2304 1079 2308
rect 1083 2304 1084 2308
rect 1288 2306 1290 2309
rect 1078 2303 1084 2304
rect 1286 2305 1292 2306
rect 110 2300 116 2301
rect 1286 2301 1287 2305
rect 1291 2301 1292 2305
rect 1286 2300 1292 2301
rect 1328 2297 1330 2317
rect 1368 2298 1370 2317
rect 1456 2298 1458 2317
rect 1544 2298 1546 2317
rect 1640 2298 1642 2317
rect 1736 2298 1738 2317
rect 1832 2298 1834 2317
rect 1928 2298 1930 2317
rect 2016 2298 2018 2317
rect 2112 2298 2114 2317
rect 2208 2298 2210 2317
rect 1366 2297 1372 2298
rect 1326 2296 1332 2297
rect 1326 2292 1327 2296
rect 1331 2292 1332 2296
rect 1366 2293 1367 2297
rect 1371 2293 1372 2297
rect 1366 2292 1372 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1542 2297 1548 2298
rect 1542 2293 1543 2297
rect 1547 2293 1548 2297
rect 1542 2292 1548 2293
rect 1638 2297 1644 2298
rect 1638 2293 1639 2297
rect 1643 2293 1644 2297
rect 1638 2292 1644 2293
rect 1734 2297 1740 2298
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1830 2297 1836 2298
rect 1830 2293 1831 2297
rect 1835 2293 1836 2297
rect 1830 2292 1836 2293
rect 1926 2297 1932 2298
rect 1926 2293 1927 2297
rect 1931 2293 1932 2297
rect 1926 2292 1932 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2110 2297 2116 2298
rect 2110 2293 2111 2297
rect 2115 2293 2116 2297
rect 2110 2292 2116 2293
rect 2206 2297 2212 2298
rect 2504 2297 2506 2317
rect 2206 2293 2207 2297
rect 2211 2293 2212 2297
rect 2206 2292 2212 2293
rect 2502 2296 2508 2297
rect 2502 2292 2503 2296
rect 2507 2292 2508 2296
rect 1326 2291 1332 2292
rect 2502 2291 2508 2292
rect 110 2288 116 2289
rect 1286 2288 1292 2289
rect 110 2284 111 2288
rect 115 2284 116 2288
rect 110 2283 116 2284
rect 222 2287 228 2288
rect 222 2283 223 2287
rect 227 2283 228 2287
rect 112 2259 114 2283
rect 222 2282 228 2283
rect 302 2287 308 2288
rect 302 2283 303 2287
rect 307 2283 308 2287
rect 302 2282 308 2283
rect 390 2287 396 2288
rect 390 2283 391 2287
rect 395 2283 396 2287
rect 390 2282 396 2283
rect 486 2287 492 2288
rect 486 2283 487 2287
rect 491 2283 492 2287
rect 486 2282 492 2283
rect 574 2287 580 2288
rect 574 2283 575 2287
rect 579 2283 580 2287
rect 574 2282 580 2283
rect 662 2287 668 2288
rect 662 2283 663 2287
rect 667 2283 668 2287
rect 662 2282 668 2283
rect 750 2287 756 2288
rect 750 2283 751 2287
rect 755 2283 756 2287
rect 750 2282 756 2283
rect 830 2287 836 2288
rect 830 2283 831 2287
rect 835 2283 836 2287
rect 830 2282 836 2283
rect 918 2287 924 2288
rect 918 2283 919 2287
rect 923 2283 924 2287
rect 918 2282 924 2283
rect 1006 2287 1012 2288
rect 1006 2283 1007 2287
rect 1011 2283 1012 2287
rect 1006 2282 1012 2283
rect 1094 2287 1100 2288
rect 1094 2283 1095 2287
rect 1099 2283 1100 2287
rect 1286 2284 1287 2288
rect 1291 2284 1292 2288
rect 1286 2283 1292 2284
rect 1094 2282 1100 2283
rect 224 2259 226 2282
rect 304 2259 306 2282
rect 392 2259 394 2282
rect 488 2259 490 2282
rect 576 2259 578 2282
rect 664 2259 666 2282
rect 752 2259 754 2282
rect 832 2259 834 2282
rect 920 2259 922 2282
rect 1008 2259 1010 2282
rect 1096 2259 1098 2282
rect 1288 2259 1290 2283
rect 1326 2279 1332 2280
rect 1326 2275 1327 2279
rect 1331 2275 1332 2279
rect 2502 2279 2508 2280
rect 1326 2274 1332 2275
rect 1350 2276 1356 2277
rect 1328 2271 1330 2274
rect 1350 2272 1351 2276
rect 1355 2272 1356 2276
rect 1350 2271 1356 2272
rect 1438 2276 1444 2277
rect 1438 2272 1439 2276
rect 1443 2272 1444 2276
rect 1438 2271 1444 2272
rect 1526 2276 1532 2277
rect 1526 2272 1527 2276
rect 1531 2272 1532 2276
rect 1526 2271 1532 2272
rect 1622 2276 1628 2277
rect 1622 2272 1623 2276
rect 1627 2272 1628 2276
rect 1622 2271 1628 2272
rect 1718 2276 1724 2277
rect 1718 2272 1719 2276
rect 1723 2272 1724 2276
rect 1718 2271 1724 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1814 2271 1820 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1998 2276 2004 2277
rect 1998 2272 1999 2276
rect 2003 2272 2004 2276
rect 1998 2271 2004 2272
rect 2094 2276 2100 2277
rect 2094 2272 2095 2276
rect 2099 2272 2100 2276
rect 2094 2271 2100 2272
rect 2190 2276 2196 2277
rect 2190 2272 2191 2276
rect 2195 2272 2196 2276
rect 2502 2275 2503 2279
rect 2507 2275 2508 2279
rect 2502 2274 2508 2275
rect 2190 2271 2196 2272
rect 2504 2271 2506 2274
rect 1327 2270 1331 2271
rect 1327 2265 1331 2266
rect 1351 2270 1355 2271
rect 1351 2265 1355 2266
rect 1439 2270 1443 2271
rect 1439 2265 1443 2266
rect 1455 2270 1459 2271
rect 1455 2265 1459 2266
rect 1527 2270 1531 2271
rect 1527 2265 1531 2266
rect 1543 2270 1547 2271
rect 1543 2265 1547 2266
rect 1623 2270 1627 2271
rect 1623 2265 1627 2266
rect 1639 2270 1643 2271
rect 1639 2265 1643 2266
rect 1719 2270 1723 2271
rect 1719 2265 1723 2266
rect 1735 2270 1739 2271
rect 1735 2265 1739 2266
rect 1815 2270 1819 2271
rect 1815 2265 1819 2266
rect 1839 2270 1843 2271
rect 1839 2265 1843 2266
rect 1911 2270 1915 2271
rect 1911 2265 1915 2266
rect 1935 2270 1939 2271
rect 1935 2265 1939 2266
rect 1999 2270 2003 2271
rect 1999 2265 2003 2266
rect 2031 2270 2035 2271
rect 2031 2265 2035 2266
rect 2095 2270 2099 2271
rect 2095 2265 2099 2266
rect 2119 2270 2123 2271
rect 2119 2265 2123 2266
rect 2191 2270 2195 2271
rect 2191 2265 2195 2266
rect 2215 2270 2219 2271
rect 2215 2265 2219 2266
rect 2311 2270 2315 2271
rect 2311 2265 2315 2266
rect 2503 2270 2507 2271
rect 2503 2265 2507 2266
rect 1328 2262 1330 2265
rect 1454 2264 1460 2265
rect 1326 2261 1332 2262
rect 111 2258 115 2259
rect 111 2253 115 2254
rect 223 2258 227 2259
rect 223 2253 227 2254
rect 263 2258 267 2259
rect 263 2253 267 2254
rect 303 2258 307 2259
rect 303 2253 307 2254
rect 319 2258 323 2259
rect 319 2253 323 2254
rect 383 2258 387 2259
rect 383 2253 387 2254
rect 391 2258 395 2259
rect 391 2253 395 2254
rect 447 2258 451 2259
rect 447 2253 451 2254
rect 487 2258 491 2259
rect 487 2253 491 2254
rect 503 2258 507 2259
rect 503 2253 507 2254
rect 559 2258 563 2259
rect 559 2253 563 2254
rect 575 2258 579 2259
rect 575 2253 579 2254
rect 615 2258 619 2259
rect 615 2253 619 2254
rect 663 2258 667 2259
rect 663 2253 667 2254
rect 671 2258 675 2259
rect 671 2253 675 2254
rect 727 2258 731 2259
rect 727 2253 731 2254
rect 751 2258 755 2259
rect 751 2253 755 2254
rect 791 2258 795 2259
rect 791 2253 795 2254
rect 831 2258 835 2259
rect 831 2253 835 2254
rect 855 2258 859 2259
rect 855 2253 859 2254
rect 919 2258 923 2259
rect 919 2253 923 2254
rect 983 2258 987 2259
rect 983 2253 987 2254
rect 1007 2258 1011 2259
rect 1007 2253 1011 2254
rect 1047 2258 1051 2259
rect 1047 2253 1051 2254
rect 1095 2258 1099 2259
rect 1095 2253 1099 2254
rect 1111 2258 1115 2259
rect 1111 2253 1115 2254
rect 1287 2258 1291 2259
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1454 2260 1455 2264
rect 1459 2260 1460 2264
rect 1454 2259 1460 2260
rect 1542 2264 1548 2265
rect 1542 2260 1543 2264
rect 1547 2260 1548 2264
rect 1542 2259 1548 2260
rect 1638 2264 1644 2265
rect 1638 2260 1639 2264
rect 1643 2260 1644 2264
rect 1638 2259 1644 2260
rect 1734 2264 1740 2265
rect 1734 2260 1735 2264
rect 1739 2260 1740 2264
rect 1734 2259 1740 2260
rect 1838 2264 1844 2265
rect 1838 2260 1839 2264
rect 1843 2260 1844 2264
rect 1838 2259 1844 2260
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 1934 2259 1940 2260
rect 2030 2264 2036 2265
rect 2030 2260 2031 2264
rect 2035 2260 2036 2264
rect 2030 2259 2036 2260
rect 2118 2264 2124 2265
rect 2118 2260 2119 2264
rect 2123 2260 2124 2264
rect 2118 2259 2124 2260
rect 2214 2264 2220 2265
rect 2214 2260 2215 2264
rect 2219 2260 2220 2264
rect 2214 2259 2220 2260
rect 2310 2264 2316 2265
rect 2310 2260 2311 2264
rect 2315 2260 2316 2264
rect 2504 2262 2506 2265
rect 2310 2259 2316 2260
rect 2502 2261 2508 2262
rect 1326 2256 1332 2257
rect 2502 2257 2503 2261
rect 2507 2257 2508 2261
rect 2502 2256 2508 2257
rect 1287 2253 1291 2254
rect 112 2233 114 2253
rect 264 2234 266 2253
rect 320 2234 322 2253
rect 384 2234 386 2253
rect 448 2234 450 2253
rect 504 2234 506 2253
rect 560 2234 562 2253
rect 616 2234 618 2253
rect 672 2234 674 2253
rect 728 2234 730 2253
rect 792 2234 794 2253
rect 856 2234 858 2253
rect 920 2234 922 2253
rect 984 2234 986 2253
rect 1048 2234 1050 2253
rect 1112 2234 1114 2253
rect 262 2233 268 2234
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 262 2229 263 2233
rect 267 2229 268 2233
rect 262 2228 268 2229
rect 318 2233 324 2234
rect 318 2229 319 2233
rect 323 2229 324 2233
rect 318 2228 324 2229
rect 382 2233 388 2234
rect 382 2229 383 2233
rect 387 2229 388 2233
rect 382 2228 388 2229
rect 446 2233 452 2234
rect 446 2229 447 2233
rect 451 2229 452 2233
rect 446 2228 452 2229
rect 502 2233 508 2234
rect 502 2229 503 2233
rect 507 2229 508 2233
rect 502 2228 508 2229
rect 558 2233 564 2234
rect 558 2229 559 2233
rect 563 2229 564 2233
rect 558 2228 564 2229
rect 614 2233 620 2234
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 670 2233 676 2234
rect 670 2229 671 2233
rect 675 2229 676 2233
rect 670 2228 676 2229
rect 726 2233 732 2234
rect 726 2229 727 2233
rect 731 2229 732 2233
rect 726 2228 732 2229
rect 790 2233 796 2234
rect 790 2229 791 2233
rect 795 2229 796 2233
rect 790 2228 796 2229
rect 854 2233 860 2234
rect 854 2229 855 2233
rect 859 2229 860 2233
rect 854 2228 860 2229
rect 918 2233 924 2234
rect 918 2229 919 2233
rect 923 2229 924 2233
rect 918 2228 924 2229
rect 982 2233 988 2234
rect 982 2229 983 2233
rect 987 2229 988 2233
rect 982 2228 988 2229
rect 1046 2233 1052 2234
rect 1046 2229 1047 2233
rect 1051 2229 1052 2233
rect 1046 2228 1052 2229
rect 1110 2233 1116 2234
rect 1288 2233 1290 2253
rect 1326 2244 1332 2245
rect 2502 2244 2508 2245
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1326 2239 1332 2240
rect 1470 2243 1476 2244
rect 1470 2239 1471 2243
rect 1475 2239 1476 2243
rect 1110 2229 1111 2233
rect 1115 2229 1116 2233
rect 1110 2228 1116 2229
rect 1286 2232 1292 2233
rect 1286 2228 1287 2232
rect 1291 2228 1292 2232
rect 110 2227 116 2228
rect 1286 2227 1292 2228
rect 110 2215 116 2216
rect 110 2211 111 2215
rect 115 2211 116 2215
rect 1286 2215 1292 2216
rect 1328 2215 1330 2239
rect 1470 2238 1476 2239
rect 1558 2243 1564 2244
rect 1558 2239 1559 2243
rect 1563 2239 1564 2243
rect 1558 2238 1564 2239
rect 1654 2243 1660 2244
rect 1654 2239 1655 2243
rect 1659 2239 1660 2243
rect 1654 2238 1660 2239
rect 1750 2243 1756 2244
rect 1750 2239 1751 2243
rect 1755 2239 1756 2243
rect 1750 2238 1756 2239
rect 1854 2243 1860 2244
rect 1854 2239 1855 2243
rect 1859 2239 1860 2243
rect 1854 2238 1860 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 2046 2243 2052 2244
rect 2046 2239 2047 2243
rect 2051 2239 2052 2243
rect 2046 2238 2052 2239
rect 2134 2243 2140 2244
rect 2134 2239 2135 2243
rect 2139 2239 2140 2243
rect 2134 2238 2140 2239
rect 2230 2243 2236 2244
rect 2230 2239 2231 2243
rect 2235 2239 2236 2243
rect 2230 2238 2236 2239
rect 2326 2243 2332 2244
rect 2326 2239 2327 2243
rect 2331 2239 2332 2243
rect 2502 2240 2503 2244
rect 2507 2240 2508 2244
rect 2502 2239 2508 2240
rect 2326 2238 2332 2239
rect 1472 2215 1474 2238
rect 1560 2215 1562 2238
rect 1656 2215 1658 2238
rect 1752 2215 1754 2238
rect 1856 2215 1858 2238
rect 1952 2215 1954 2238
rect 2048 2215 2050 2238
rect 2136 2215 2138 2238
rect 2232 2215 2234 2238
rect 2328 2215 2330 2238
rect 2504 2215 2506 2239
rect 110 2210 116 2211
rect 246 2212 252 2213
rect 112 2203 114 2210
rect 246 2208 247 2212
rect 251 2208 252 2212
rect 246 2207 252 2208
rect 302 2212 308 2213
rect 302 2208 303 2212
rect 307 2208 308 2212
rect 302 2207 308 2208
rect 366 2212 372 2213
rect 366 2208 367 2212
rect 371 2208 372 2212
rect 366 2207 372 2208
rect 430 2212 436 2213
rect 430 2208 431 2212
rect 435 2208 436 2212
rect 430 2207 436 2208
rect 486 2212 492 2213
rect 486 2208 487 2212
rect 491 2208 492 2212
rect 486 2207 492 2208
rect 542 2212 548 2213
rect 542 2208 543 2212
rect 547 2208 548 2212
rect 542 2207 548 2208
rect 598 2212 604 2213
rect 598 2208 599 2212
rect 603 2208 604 2212
rect 598 2207 604 2208
rect 654 2212 660 2213
rect 654 2208 655 2212
rect 659 2208 660 2212
rect 654 2207 660 2208
rect 710 2212 716 2213
rect 710 2208 711 2212
rect 715 2208 716 2212
rect 710 2207 716 2208
rect 774 2212 780 2213
rect 774 2208 775 2212
rect 779 2208 780 2212
rect 774 2207 780 2208
rect 838 2212 844 2213
rect 838 2208 839 2212
rect 843 2208 844 2212
rect 838 2207 844 2208
rect 902 2212 908 2213
rect 902 2208 903 2212
rect 907 2208 908 2212
rect 902 2207 908 2208
rect 966 2212 972 2213
rect 966 2208 967 2212
rect 971 2208 972 2212
rect 966 2207 972 2208
rect 1030 2212 1036 2213
rect 1030 2208 1031 2212
rect 1035 2208 1036 2212
rect 1030 2207 1036 2208
rect 1094 2212 1100 2213
rect 1094 2208 1095 2212
rect 1099 2208 1100 2212
rect 1286 2211 1287 2215
rect 1291 2211 1292 2215
rect 1286 2210 1292 2211
rect 1327 2214 1331 2215
rect 1094 2207 1100 2208
rect 248 2203 250 2207
rect 304 2203 306 2207
rect 368 2203 370 2207
rect 432 2203 434 2207
rect 488 2203 490 2207
rect 544 2203 546 2207
rect 600 2203 602 2207
rect 656 2203 658 2207
rect 712 2203 714 2207
rect 776 2203 778 2207
rect 840 2203 842 2207
rect 904 2203 906 2207
rect 968 2203 970 2207
rect 1032 2203 1034 2207
rect 1096 2203 1098 2207
rect 1288 2203 1290 2210
rect 1327 2209 1331 2210
rect 1471 2214 1475 2215
rect 1471 2209 1475 2210
rect 1559 2214 1563 2215
rect 1559 2209 1563 2210
rect 1567 2214 1571 2215
rect 1567 2209 1571 2210
rect 1623 2214 1627 2215
rect 1623 2209 1627 2210
rect 1655 2214 1659 2215
rect 1655 2209 1659 2210
rect 1679 2214 1683 2215
rect 1679 2209 1683 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1751 2214 1755 2215
rect 1751 2209 1755 2210
rect 1807 2214 1811 2215
rect 1807 2209 1811 2210
rect 1855 2214 1859 2215
rect 1855 2209 1859 2210
rect 1871 2214 1875 2215
rect 1871 2209 1875 2210
rect 1927 2214 1931 2215
rect 1927 2209 1931 2210
rect 1951 2214 1955 2215
rect 1951 2209 1955 2210
rect 1983 2214 1987 2215
rect 1983 2209 1987 2210
rect 2039 2214 2043 2215
rect 2039 2209 2043 2210
rect 2047 2214 2051 2215
rect 2047 2209 2051 2210
rect 2095 2214 2099 2215
rect 2095 2209 2099 2210
rect 2135 2214 2139 2215
rect 2135 2209 2139 2210
rect 2159 2214 2163 2215
rect 2159 2209 2163 2210
rect 2223 2214 2227 2215
rect 2223 2209 2227 2210
rect 2231 2214 2235 2215
rect 2231 2209 2235 2210
rect 2287 2214 2291 2215
rect 2287 2209 2291 2210
rect 2327 2214 2331 2215
rect 2327 2209 2331 2210
rect 2343 2214 2347 2215
rect 2343 2209 2347 2210
rect 2399 2214 2403 2215
rect 2399 2209 2403 2210
rect 2455 2214 2459 2215
rect 2455 2209 2459 2210
rect 2503 2214 2507 2215
rect 2503 2209 2507 2210
rect 111 2202 115 2203
rect 111 2197 115 2198
rect 247 2202 251 2203
rect 247 2197 251 2198
rect 303 2202 307 2203
rect 303 2197 307 2198
rect 335 2202 339 2203
rect 335 2197 339 2198
rect 367 2202 371 2203
rect 367 2197 371 2198
rect 391 2202 395 2203
rect 391 2197 395 2198
rect 431 2202 435 2203
rect 431 2197 435 2198
rect 447 2202 451 2203
rect 447 2197 451 2198
rect 487 2202 491 2203
rect 487 2197 491 2198
rect 503 2202 507 2203
rect 503 2197 507 2198
rect 543 2202 547 2203
rect 543 2197 547 2198
rect 559 2202 563 2203
rect 559 2197 563 2198
rect 599 2202 603 2203
rect 599 2197 603 2198
rect 655 2202 659 2203
rect 655 2197 659 2198
rect 711 2202 715 2203
rect 711 2197 715 2198
rect 775 2202 779 2203
rect 775 2197 779 2198
rect 839 2202 843 2203
rect 839 2197 843 2198
rect 903 2202 907 2203
rect 903 2197 907 2198
rect 967 2202 971 2203
rect 967 2197 971 2198
rect 1031 2202 1035 2203
rect 1031 2197 1035 2198
rect 1095 2202 1099 2203
rect 1095 2197 1099 2198
rect 1287 2202 1291 2203
rect 1287 2197 1291 2198
rect 112 2194 114 2197
rect 334 2196 340 2197
rect 110 2193 116 2194
rect 110 2189 111 2193
rect 115 2189 116 2193
rect 334 2192 335 2196
rect 339 2192 340 2196
rect 334 2191 340 2192
rect 390 2196 396 2197
rect 390 2192 391 2196
rect 395 2192 396 2196
rect 390 2191 396 2192
rect 446 2196 452 2197
rect 446 2192 447 2196
rect 451 2192 452 2196
rect 446 2191 452 2192
rect 502 2196 508 2197
rect 502 2192 503 2196
rect 507 2192 508 2196
rect 502 2191 508 2192
rect 558 2196 564 2197
rect 558 2192 559 2196
rect 563 2192 564 2196
rect 1288 2194 1290 2197
rect 558 2191 564 2192
rect 1286 2193 1292 2194
rect 110 2188 116 2189
rect 1286 2189 1287 2193
rect 1291 2189 1292 2193
rect 1328 2189 1330 2209
rect 1568 2190 1570 2209
rect 1624 2190 1626 2209
rect 1680 2190 1682 2209
rect 1744 2190 1746 2209
rect 1808 2190 1810 2209
rect 1872 2190 1874 2209
rect 1928 2190 1930 2209
rect 1984 2190 1986 2209
rect 2040 2190 2042 2209
rect 2096 2190 2098 2209
rect 2160 2190 2162 2209
rect 2224 2190 2226 2209
rect 2288 2190 2290 2209
rect 2344 2190 2346 2209
rect 2400 2190 2402 2209
rect 2456 2190 2458 2209
rect 1566 2189 1572 2190
rect 1286 2188 1292 2189
rect 1326 2188 1332 2189
rect 1326 2184 1327 2188
rect 1331 2184 1332 2188
rect 1566 2185 1567 2189
rect 1571 2185 1572 2189
rect 1566 2184 1572 2185
rect 1622 2189 1628 2190
rect 1622 2185 1623 2189
rect 1627 2185 1628 2189
rect 1622 2184 1628 2185
rect 1678 2189 1684 2190
rect 1678 2185 1679 2189
rect 1683 2185 1684 2189
rect 1678 2184 1684 2185
rect 1742 2189 1748 2190
rect 1742 2185 1743 2189
rect 1747 2185 1748 2189
rect 1742 2184 1748 2185
rect 1806 2189 1812 2190
rect 1806 2185 1807 2189
rect 1811 2185 1812 2189
rect 1806 2184 1812 2185
rect 1870 2189 1876 2190
rect 1870 2185 1871 2189
rect 1875 2185 1876 2189
rect 1870 2184 1876 2185
rect 1926 2189 1932 2190
rect 1926 2185 1927 2189
rect 1931 2185 1932 2189
rect 1926 2184 1932 2185
rect 1982 2189 1988 2190
rect 1982 2185 1983 2189
rect 1987 2185 1988 2189
rect 1982 2184 1988 2185
rect 2038 2189 2044 2190
rect 2038 2185 2039 2189
rect 2043 2185 2044 2189
rect 2038 2184 2044 2185
rect 2094 2189 2100 2190
rect 2094 2185 2095 2189
rect 2099 2185 2100 2189
rect 2094 2184 2100 2185
rect 2158 2189 2164 2190
rect 2158 2185 2159 2189
rect 2163 2185 2164 2189
rect 2158 2184 2164 2185
rect 2222 2189 2228 2190
rect 2222 2185 2223 2189
rect 2227 2185 2228 2189
rect 2222 2184 2228 2185
rect 2286 2189 2292 2190
rect 2286 2185 2287 2189
rect 2291 2185 2292 2189
rect 2286 2184 2292 2185
rect 2342 2189 2348 2190
rect 2342 2185 2343 2189
rect 2347 2185 2348 2189
rect 2342 2184 2348 2185
rect 2398 2189 2404 2190
rect 2398 2185 2399 2189
rect 2403 2185 2404 2189
rect 2398 2184 2404 2185
rect 2454 2189 2460 2190
rect 2504 2189 2506 2209
rect 2454 2185 2455 2189
rect 2459 2185 2460 2189
rect 2454 2184 2460 2185
rect 2502 2188 2508 2189
rect 2502 2184 2503 2188
rect 2507 2184 2508 2188
rect 1326 2183 1332 2184
rect 2502 2183 2508 2184
rect 110 2176 116 2177
rect 1286 2176 1292 2177
rect 110 2172 111 2176
rect 115 2172 116 2176
rect 110 2171 116 2172
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 112 2151 114 2171
rect 350 2170 356 2171
rect 406 2175 412 2176
rect 406 2171 407 2175
rect 411 2171 412 2175
rect 406 2170 412 2171
rect 462 2175 468 2176
rect 462 2171 463 2175
rect 467 2171 468 2175
rect 462 2170 468 2171
rect 518 2175 524 2176
rect 518 2171 519 2175
rect 523 2171 524 2175
rect 518 2170 524 2171
rect 574 2175 580 2176
rect 574 2171 575 2175
rect 579 2171 580 2175
rect 1286 2172 1287 2176
rect 1291 2172 1292 2176
rect 1286 2171 1292 2172
rect 1326 2171 1332 2172
rect 574 2170 580 2171
rect 352 2151 354 2170
rect 408 2151 410 2170
rect 464 2151 466 2170
rect 520 2151 522 2170
rect 576 2151 578 2170
rect 1288 2151 1290 2171
rect 1326 2167 1327 2171
rect 1331 2167 1332 2171
rect 2502 2171 2508 2172
rect 1326 2166 1332 2167
rect 1550 2168 1556 2169
rect 1328 2151 1330 2166
rect 1550 2164 1551 2168
rect 1555 2164 1556 2168
rect 1550 2163 1556 2164
rect 1606 2168 1612 2169
rect 1606 2164 1607 2168
rect 1611 2164 1612 2168
rect 1606 2163 1612 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1726 2168 1732 2169
rect 1726 2164 1727 2168
rect 1731 2164 1732 2168
rect 1726 2163 1732 2164
rect 1790 2168 1796 2169
rect 1790 2164 1791 2168
rect 1795 2164 1796 2168
rect 1790 2163 1796 2164
rect 1854 2168 1860 2169
rect 1854 2164 1855 2168
rect 1859 2164 1860 2168
rect 1854 2163 1860 2164
rect 1910 2168 1916 2169
rect 1910 2164 1911 2168
rect 1915 2164 1916 2168
rect 1910 2163 1916 2164
rect 1966 2168 1972 2169
rect 1966 2164 1967 2168
rect 1971 2164 1972 2168
rect 1966 2163 1972 2164
rect 2022 2168 2028 2169
rect 2022 2164 2023 2168
rect 2027 2164 2028 2168
rect 2022 2163 2028 2164
rect 2078 2168 2084 2169
rect 2078 2164 2079 2168
rect 2083 2164 2084 2168
rect 2078 2163 2084 2164
rect 2142 2168 2148 2169
rect 2142 2164 2143 2168
rect 2147 2164 2148 2168
rect 2142 2163 2148 2164
rect 2206 2168 2212 2169
rect 2206 2164 2207 2168
rect 2211 2164 2212 2168
rect 2206 2163 2212 2164
rect 2270 2168 2276 2169
rect 2270 2164 2271 2168
rect 2275 2164 2276 2168
rect 2270 2163 2276 2164
rect 2326 2168 2332 2169
rect 2326 2164 2327 2168
rect 2331 2164 2332 2168
rect 2326 2163 2332 2164
rect 2382 2168 2388 2169
rect 2382 2164 2383 2168
rect 2387 2164 2388 2168
rect 2382 2163 2388 2164
rect 2438 2168 2444 2169
rect 2438 2164 2439 2168
rect 2443 2164 2444 2168
rect 2502 2167 2503 2171
rect 2507 2167 2508 2171
rect 2502 2166 2508 2167
rect 2438 2163 2444 2164
rect 1552 2151 1554 2163
rect 1608 2151 1610 2163
rect 1664 2151 1666 2163
rect 1728 2151 1730 2163
rect 1792 2151 1794 2163
rect 1856 2151 1858 2163
rect 1912 2151 1914 2163
rect 1968 2151 1970 2163
rect 2024 2151 2026 2163
rect 2080 2151 2082 2163
rect 2144 2151 2146 2163
rect 2208 2151 2210 2163
rect 2272 2151 2274 2163
rect 2328 2151 2330 2163
rect 2384 2151 2386 2163
rect 2440 2151 2442 2163
rect 2504 2151 2506 2166
rect 111 2150 115 2151
rect 111 2145 115 2146
rect 351 2150 355 2151
rect 351 2145 355 2146
rect 407 2150 411 2151
rect 407 2145 411 2146
rect 415 2150 419 2151
rect 415 2145 419 2146
rect 463 2150 467 2151
rect 463 2145 467 2146
rect 511 2150 515 2151
rect 511 2145 515 2146
rect 519 2150 523 2151
rect 519 2145 523 2146
rect 575 2150 579 2151
rect 575 2145 579 2146
rect 607 2150 611 2151
rect 607 2145 611 2146
rect 711 2150 715 2151
rect 711 2145 715 2146
rect 815 2150 819 2151
rect 815 2145 819 2146
rect 927 2150 931 2151
rect 927 2145 931 2146
rect 1039 2150 1043 2151
rect 1039 2145 1043 2146
rect 1151 2150 1155 2151
rect 1151 2145 1155 2146
rect 1239 2150 1243 2151
rect 1239 2145 1243 2146
rect 1287 2150 1291 2151
rect 1287 2145 1291 2146
rect 1327 2150 1331 2151
rect 1327 2145 1331 2146
rect 1551 2150 1555 2151
rect 1551 2145 1555 2146
rect 1607 2150 1611 2151
rect 1607 2145 1611 2146
rect 1663 2150 1667 2151
rect 1663 2145 1667 2146
rect 1719 2150 1723 2151
rect 1719 2145 1723 2146
rect 1727 2150 1731 2151
rect 1727 2145 1731 2146
rect 1791 2150 1795 2151
rect 1791 2145 1795 2146
rect 1855 2150 1859 2151
rect 1855 2145 1859 2146
rect 1871 2150 1875 2151
rect 1871 2145 1875 2146
rect 1911 2150 1915 2151
rect 1911 2145 1915 2146
rect 1967 2150 1971 2151
rect 1967 2145 1971 2146
rect 2023 2150 2027 2151
rect 2023 2145 2027 2146
rect 2079 2150 2083 2151
rect 2079 2145 2083 2146
rect 2143 2150 2147 2151
rect 2143 2145 2147 2146
rect 2199 2150 2203 2151
rect 2199 2145 2203 2146
rect 2207 2150 2211 2151
rect 2207 2145 2211 2146
rect 2271 2150 2275 2151
rect 2271 2145 2275 2146
rect 2327 2150 2331 2151
rect 2327 2145 2331 2146
rect 2383 2150 2387 2151
rect 2383 2145 2387 2146
rect 2439 2150 2443 2151
rect 2439 2145 2443 2146
rect 2503 2150 2507 2151
rect 2503 2145 2507 2146
rect 112 2125 114 2145
rect 416 2126 418 2145
rect 512 2126 514 2145
rect 608 2126 610 2145
rect 712 2126 714 2145
rect 816 2126 818 2145
rect 928 2126 930 2145
rect 1040 2126 1042 2145
rect 1152 2126 1154 2145
rect 1240 2126 1242 2145
rect 414 2125 420 2126
rect 110 2124 116 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 414 2121 415 2125
rect 419 2121 420 2125
rect 414 2120 420 2121
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 606 2125 612 2126
rect 606 2121 607 2125
rect 611 2121 612 2125
rect 606 2120 612 2121
rect 710 2125 716 2126
rect 710 2121 711 2125
rect 715 2121 716 2125
rect 710 2120 716 2121
rect 814 2125 820 2126
rect 814 2121 815 2125
rect 819 2121 820 2125
rect 814 2120 820 2121
rect 926 2125 932 2126
rect 926 2121 927 2125
rect 931 2121 932 2125
rect 926 2120 932 2121
rect 1038 2125 1044 2126
rect 1038 2121 1039 2125
rect 1043 2121 1044 2125
rect 1038 2120 1044 2121
rect 1150 2125 1156 2126
rect 1150 2121 1151 2125
rect 1155 2121 1156 2125
rect 1150 2120 1156 2121
rect 1238 2125 1244 2126
rect 1288 2125 1290 2145
rect 1328 2142 1330 2145
rect 1662 2144 1668 2145
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1718 2144 1724 2145
rect 1718 2140 1719 2144
rect 1723 2140 1724 2144
rect 1718 2139 1724 2140
rect 1790 2144 1796 2145
rect 1790 2140 1791 2144
rect 1795 2140 1796 2144
rect 1790 2139 1796 2140
rect 1870 2144 1876 2145
rect 1870 2140 1871 2144
rect 1875 2140 1876 2144
rect 1870 2139 1876 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2078 2144 2084 2145
rect 2078 2140 2079 2144
rect 2083 2140 2084 2144
rect 2078 2139 2084 2140
rect 2198 2144 2204 2145
rect 2198 2140 2199 2144
rect 2203 2140 2204 2144
rect 2198 2139 2204 2140
rect 2326 2144 2332 2145
rect 2326 2140 2327 2144
rect 2331 2140 2332 2144
rect 2326 2139 2332 2140
rect 2438 2144 2444 2145
rect 2438 2140 2439 2144
rect 2443 2140 2444 2144
rect 2504 2142 2506 2145
rect 2438 2139 2444 2140
rect 2502 2141 2508 2142
rect 1326 2136 1332 2137
rect 2502 2137 2503 2141
rect 2507 2137 2508 2141
rect 2502 2136 2508 2137
rect 1238 2121 1239 2125
rect 1243 2121 1244 2125
rect 1238 2120 1244 2121
rect 1286 2124 1292 2125
rect 1286 2120 1287 2124
rect 1291 2120 1292 2124
rect 110 2119 116 2120
rect 1286 2119 1292 2120
rect 1326 2124 1332 2125
rect 2502 2124 2508 2125
rect 1326 2120 1327 2124
rect 1331 2120 1332 2124
rect 1326 2119 1332 2120
rect 1678 2123 1684 2124
rect 1678 2119 1679 2123
rect 1683 2119 1684 2123
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 1286 2107 1292 2108
rect 110 2102 116 2103
rect 398 2104 404 2105
rect 112 2099 114 2102
rect 398 2100 399 2104
rect 403 2100 404 2104
rect 398 2099 404 2100
rect 494 2104 500 2105
rect 494 2100 495 2104
rect 499 2100 500 2104
rect 494 2099 500 2100
rect 590 2104 596 2105
rect 590 2100 591 2104
rect 595 2100 596 2104
rect 590 2099 596 2100
rect 694 2104 700 2105
rect 694 2100 695 2104
rect 699 2100 700 2104
rect 694 2099 700 2100
rect 798 2104 804 2105
rect 798 2100 799 2104
rect 803 2100 804 2104
rect 798 2099 804 2100
rect 910 2104 916 2105
rect 910 2100 911 2104
rect 915 2100 916 2104
rect 910 2099 916 2100
rect 1022 2104 1028 2105
rect 1022 2100 1023 2104
rect 1027 2100 1028 2104
rect 1022 2099 1028 2100
rect 1134 2104 1140 2105
rect 1134 2100 1135 2104
rect 1139 2100 1140 2104
rect 1134 2099 1140 2100
rect 1222 2104 1228 2105
rect 1222 2100 1223 2104
rect 1227 2100 1228 2104
rect 1286 2103 1287 2107
rect 1291 2103 1292 2107
rect 1286 2102 1292 2103
rect 1222 2099 1228 2100
rect 1288 2099 1290 2102
rect 111 2098 115 2099
rect 111 2093 115 2094
rect 375 2098 379 2099
rect 375 2093 379 2094
rect 399 2098 403 2099
rect 399 2093 403 2094
rect 447 2098 451 2099
rect 447 2093 451 2094
rect 495 2098 499 2099
rect 495 2093 499 2094
rect 519 2098 523 2099
rect 519 2093 523 2094
rect 591 2098 595 2099
rect 591 2093 595 2094
rect 599 2098 603 2099
rect 599 2093 603 2094
rect 679 2098 683 2099
rect 679 2093 683 2094
rect 695 2098 699 2099
rect 695 2093 699 2094
rect 759 2098 763 2099
rect 759 2093 763 2094
rect 799 2098 803 2099
rect 799 2093 803 2094
rect 831 2098 835 2099
rect 831 2093 835 2094
rect 903 2098 907 2099
rect 903 2093 907 2094
rect 911 2098 915 2099
rect 911 2093 915 2094
rect 967 2098 971 2099
rect 967 2093 971 2094
rect 1023 2098 1027 2099
rect 1023 2093 1027 2094
rect 1031 2098 1035 2099
rect 1031 2093 1035 2094
rect 1103 2098 1107 2099
rect 1103 2093 1107 2094
rect 1135 2098 1139 2099
rect 1135 2093 1139 2094
rect 1167 2098 1171 2099
rect 1167 2093 1171 2094
rect 1223 2098 1227 2099
rect 1223 2093 1227 2094
rect 1287 2098 1291 2099
rect 1287 2093 1291 2094
rect 112 2090 114 2093
rect 374 2092 380 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 446 2092 452 2093
rect 446 2088 447 2092
rect 451 2088 452 2092
rect 446 2087 452 2088
rect 518 2092 524 2093
rect 518 2088 519 2092
rect 523 2088 524 2092
rect 518 2087 524 2088
rect 598 2092 604 2093
rect 598 2088 599 2092
rect 603 2088 604 2092
rect 598 2087 604 2088
rect 678 2092 684 2093
rect 678 2088 679 2092
rect 683 2088 684 2092
rect 678 2087 684 2088
rect 758 2092 764 2093
rect 758 2088 759 2092
rect 763 2088 764 2092
rect 758 2087 764 2088
rect 830 2092 836 2093
rect 830 2088 831 2092
rect 835 2088 836 2092
rect 830 2087 836 2088
rect 902 2092 908 2093
rect 902 2088 903 2092
rect 907 2088 908 2092
rect 902 2087 908 2088
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 1030 2092 1036 2093
rect 1030 2088 1031 2092
rect 1035 2088 1036 2092
rect 1030 2087 1036 2088
rect 1102 2092 1108 2093
rect 1102 2088 1103 2092
rect 1107 2088 1108 2092
rect 1102 2087 1108 2088
rect 1166 2092 1172 2093
rect 1166 2088 1167 2092
rect 1171 2088 1172 2092
rect 1166 2087 1172 2088
rect 1222 2092 1228 2093
rect 1222 2088 1223 2092
rect 1227 2088 1228 2092
rect 1288 2090 1290 2093
rect 1222 2087 1228 2088
rect 1286 2089 1292 2090
rect 110 2084 116 2085
rect 1286 2085 1287 2089
rect 1291 2085 1292 2089
rect 1328 2087 1330 2119
rect 1678 2118 1684 2119
rect 1734 2123 1740 2124
rect 1734 2119 1735 2123
rect 1739 2119 1740 2123
rect 1734 2118 1740 2119
rect 1806 2123 1812 2124
rect 1806 2119 1807 2123
rect 1811 2119 1812 2123
rect 1806 2118 1812 2119
rect 1886 2123 1892 2124
rect 1886 2119 1887 2123
rect 1891 2119 1892 2123
rect 1886 2118 1892 2119
rect 1982 2123 1988 2124
rect 1982 2119 1983 2123
rect 1987 2119 1988 2123
rect 1982 2118 1988 2119
rect 2094 2123 2100 2124
rect 2094 2119 2095 2123
rect 2099 2119 2100 2123
rect 2094 2118 2100 2119
rect 2214 2123 2220 2124
rect 2214 2119 2215 2123
rect 2219 2119 2220 2123
rect 2214 2118 2220 2119
rect 2342 2123 2348 2124
rect 2342 2119 2343 2123
rect 2347 2119 2348 2123
rect 2342 2118 2348 2119
rect 2454 2123 2460 2124
rect 2454 2119 2455 2123
rect 2459 2119 2460 2123
rect 2502 2120 2503 2124
rect 2507 2120 2508 2124
rect 2502 2119 2508 2120
rect 2454 2118 2460 2119
rect 1680 2087 1682 2118
rect 1736 2087 1738 2118
rect 1808 2087 1810 2118
rect 1888 2087 1890 2118
rect 1984 2087 1986 2118
rect 2096 2087 2098 2118
rect 2216 2087 2218 2118
rect 2344 2087 2346 2118
rect 2456 2087 2458 2118
rect 2504 2087 2506 2119
rect 1286 2084 1292 2085
rect 1327 2086 1331 2087
rect 1327 2081 1331 2082
rect 1367 2086 1371 2087
rect 1367 2081 1371 2082
rect 1423 2086 1427 2087
rect 1423 2081 1427 2082
rect 1503 2086 1507 2087
rect 1503 2081 1507 2082
rect 1591 2086 1595 2087
rect 1591 2081 1595 2082
rect 1679 2086 1683 2087
rect 1679 2081 1683 2082
rect 1735 2086 1739 2087
rect 1735 2081 1739 2082
rect 1783 2086 1787 2087
rect 1783 2081 1787 2082
rect 1807 2086 1811 2087
rect 1807 2081 1811 2082
rect 1887 2086 1891 2087
rect 1887 2081 1891 2082
rect 1895 2086 1899 2087
rect 1895 2081 1899 2082
rect 1983 2086 1987 2087
rect 1983 2081 1987 2082
rect 2023 2086 2027 2087
rect 2023 2081 2027 2082
rect 2095 2086 2099 2087
rect 2095 2081 2099 2082
rect 2167 2086 2171 2087
rect 2167 2081 2171 2082
rect 2215 2086 2219 2087
rect 2215 2081 2219 2082
rect 2319 2086 2323 2087
rect 2319 2081 2323 2082
rect 2343 2086 2347 2087
rect 2343 2081 2347 2082
rect 2455 2086 2459 2087
rect 2455 2081 2459 2082
rect 2503 2086 2507 2087
rect 2503 2081 2507 2082
rect 110 2072 116 2073
rect 1286 2072 1292 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 390 2071 396 2072
rect 390 2067 391 2071
rect 395 2067 396 2071
rect 112 2043 114 2067
rect 390 2066 396 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 534 2071 540 2072
rect 534 2067 535 2071
rect 539 2067 540 2071
rect 534 2066 540 2067
rect 614 2071 620 2072
rect 614 2067 615 2071
rect 619 2067 620 2071
rect 614 2066 620 2067
rect 694 2071 700 2072
rect 694 2067 695 2071
rect 699 2067 700 2071
rect 694 2066 700 2067
rect 774 2071 780 2072
rect 774 2067 775 2071
rect 779 2067 780 2071
rect 774 2066 780 2067
rect 846 2071 852 2072
rect 846 2067 847 2071
rect 851 2067 852 2071
rect 846 2066 852 2067
rect 918 2071 924 2072
rect 918 2067 919 2071
rect 923 2067 924 2071
rect 918 2066 924 2067
rect 982 2071 988 2072
rect 982 2067 983 2071
rect 987 2067 988 2071
rect 982 2066 988 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1118 2071 1124 2072
rect 1118 2067 1119 2071
rect 1123 2067 1124 2071
rect 1118 2066 1124 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 1238 2071 1244 2072
rect 1238 2067 1239 2071
rect 1243 2067 1244 2071
rect 1286 2068 1287 2072
rect 1291 2068 1292 2072
rect 1286 2067 1292 2068
rect 1238 2066 1244 2067
rect 392 2043 394 2066
rect 464 2043 466 2066
rect 536 2043 538 2066
rect 616 2043 618 2066
rect 696 2043 698 2066
rect 776 2043 778 2066
rect 848 2043 850 2066
rect 920 2043 922 2066
rect 984 2043 986 2066
rect 1048 2043 1050 2066
rect 1120 2043 1122 2066
rect 1184 2043 1186 2066
rect 1240 2043 1242 2066
rect 1288 2043 1290 2067
rect 1328 2061 1330 2081
rect 1368 2062 1370 2081
rect 1424 2062 1426 2081
rect 1504 2062 1506 2081
rect 1592 2062 1594 2081
rect 1680 2062 1682 2081
rect 1784 2062 1786 2081
rect 1896 2062 1898 2081
rect 2024 2062 2026 2081
rect 2168 2062 2170 2081
rect 2320 2062 2322 2081
rect 2456 2062 2458 2081
rect 1366 2061 1372 2062
rect 1326 2060 1332 2061
rect 1326 2056 1327 2060
rect 1331 2056 1332 2060
rect 1366 2057 1367 2061
rect 1371 2057 1372 2061
rect 1366 2056 1372 2057
rect 1422 2061 1428 2062
rect 1422 2057 1423 2061
rect 1427 2057 1428 2061
rect 1422 2056 1428 2057
rect 1502 2061 1508 2062
rect 1502 2057 1503 2061
rect 1507 2057 1508 2061
rect 1502 2056 1508 2057
rect 1590 2061 1596 2062
rect 1590 2057 1591 2061
rect 1595 2057 1596 2061
rect 1590 2056 1596 2057
rect 1678 2061 1684 2062
rect 1678 2057 1679 2061
rect 1683 2057 1684 2061
rect 1678 2056 1684 2057
rect 1782 2061 1788 2062
rect 1782 2057 1783 2061
rect 1787 2057 1788 2061
rect 1782 2056 1788 2057
rect 1894 2061 1900 2062
rect 1894 2057 1895 2061
rect 1899 2057 1900 2061
rect 1894 2056 1900 2057
rect 2022 2061 2028 2062
rect 2022 2057 2023 2061
rect 2027 2057 2028 2061
rect 2022 2056 2028 2057
rect 2166 2061 2172 2062
rect 2166 2057 2167 2061
rect 2171 2057 2172 2061
rect 2166 2056 2172 2057
rect 2318 2061 2324 2062
rect 2318 2057 2319 2061
rect 2323 2057 2324 2061
rect 2318 2056 2324 2057
rect 2454 2061 2460 2062
rect 2504 2061 2506 2081
rect 2454 2057 2455 2061
rect 2459 2057 2460 2061
rect 2454 2056 2460 2057
rect 2502 2060 2508 2061
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 1326 2055 1332 2056
rect 2502 2055 2508 2056
rect 1326 2043 1332 2044
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 295 2042 299 2043
rect 295 2037 299 2038
rect 375 2042 379 2043
rect 375 2037 379 2038
rect 391 2042 395 2043
rect 391 2037 395 2038
rect 463 2042 467 2043
rect 463 2037 467 2038
rect 535 2042 539 2043
rect 535 2037 539 2038
rect 551 2042 555 2043
rect 551 2037 555 2038
rect 615 2042 619 2043
rect 615 2037 619 2038
rect 639 2042 643 2043
rect 639 2037 643 2038
rect 695 2042 699 2043
rect 695 2037 699 2038
rect 719 2042 723 2043
rect 719 2037 723 2038
rect 775 2042 779 2043
rect 775 2037 779 2038
rect 799 2042 803 2043
rect 799 2037 803 2038
rect 847 2042 851 2043
rect 847 2037 851 2038
rect 887 2042 891 2043
rect 887 2037 891 2038
rect 919 2042 923 2043
rect 919 2037 923 2038
rect 975 2042 979 2043
rect 975 2037 979 2038
rect 983 2042 987 2043
rect 983 2037 987 2038
rect 1047 2042 1051 2043
rect 1047 2037 1051 2038
rect 1063 2042 1067 2043
rect 1063 2037 1067 2038
rect 1119 2042 1123 2043
rect 1119 2037 1123 2038
rect 1183 2042 1187 2043
rect 1183 2037 1187 2038
rect 1239 2042 1243 2043
rect 1239 2037 1243 2038
rect 1287 2042 1291 2043
rect 1326 2039 1327 2043
rect 1331 2039 1332 2043
rect 2502 2043 2508 2044
rect 1326 2038 1332 2039
rect 1350 2040 1356 2041
rect 1287 2037 1291 2038
rect 112 2017 114 2037
rect 296 2018 298 2037
rect 376 2018 378 2037
rect 464 2018 466 2037
rect 552 2018 554 2037
rect 640 2018 642 2037
rect 720 2018 722 2037
rect 800 2018 802 2037
rect 888 2018 890 2037
rect 976 2018 978 2037
rect 1064 2018 1066 2037
rect 294 2017 300 2018
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 294 2013 295 2017
rect 299 2013 300 2017
rect 294 2012 300 2013
rect 374 2017 380 2018
rect 374 2013 375 2017
rect 379 2013 380 2017
rect 374 2012 380 2013
rect 462 2017 468 2018
rect 462 2013 463 2017
rect 467 2013 468 2017
rect 462 2012 468 2013
rect 550 2017 556 2018
rect 550 2013 551 2017
rect 555 2013 556 2017
rect 550 2012 556 2013
rect 638 2017 644 2018
rect 638 2013 639 2017
rect 643 2013 644 2017
rect 638 2012 644 2013
rect 718 2017 724 2018
rect 718 2013 719 2017
rect 723 2013 724 2017
rect 718 2012 724 2013
rect 798 2017 804 2018
rect 798 2013 799 2017
rect 803 2013 804 2017
rect 798 2012 804 2013
rect 886 2017 892 2018
rect 886 2013 887 2017
rect 891 2013 892 2017
rect 886 2012 892 2013
rect 974 2017 980 2018
rect 974 2013 975 2017
rect 979 2013 980 2017
rect 974 2012 980 2013
rect 1062 2017 1068 2018
rect 1288 2017 1290 2037
rect 1328 2035 1330 2038
rect 1350 2036 1351 2040
rect 1355 2036 1356 2040
rect 1350 2035 1356 2036
rect 1406 2040 1412 2041
rect 1406 2036 1407 2040
rect 1411 2036 1412 2040
rect 1406 2035 1412 2036
rect 1486 2040 1492 2041
rect 1486 2036 1487 2040
rect 1491 2036 1492 2040
rect 1486 2035 1492 2036
rect 1574 2040 1580 2041
rect 1574 2036 1575 2040
rect 1579 2036 1580 2040
rect 1574 2035 1580 2036
rect 1662 2040 1668 2041
rect 1662 2036 1663 2040
rect 1667 2036 1668 2040
rect 1662 2035 1668 2036
rect 1766 2040 1772 2041
rect 1766 2036 1767 2040
rect 1771 2036 1772 2040
rect 1766 2035 1772 2036
rect 1878 2040 1884 2041
rect 1878 2036 1879 2040
rect 1883 2036 1884 2040
rect 1878 2035 1884 2036
rect 2006 2040 2012 2041
rect 2006 2036 2007 2040
rect 2011 2036 2012 2040
rect 2006 2035 2012 2036
rect 2150 2040 2156 2041
rect 2150 2036 2151 2040
rect 2155 2036 2156 2040
rect 2150 2035 2156 2036
rect 2302 2040 2308 2041
rect 2302 2036 2303 2040
rect 2307 2036 2308 2040
rect 2302 2035 2308 2036
rect 2438 2040 2444 2041
rect 2438 2036 2439 2040
rect 2443 2036 2444 2040
rect 2502 2039 2503 2043
rect 2507 2039 2508 2043
rect 2502 2038 2508 2039
rect 2438 2035 2444 2036
rect 2504 2035 2506 2038
rect 1327 2034 1331 2035
rect 1327 2029 1331 2030
rect 1351 2034 1355 2035
rect 1351 2029 1355 2030
rect 1407 2034 1411 2035
rect 1407 2029 1411 2030
rect 1423 2034 1427 2035
rect 1423 2029 1427 2030
rect 1487 2034 1491 2035
rect 1487 2029 1491 2030
rect 1519 2034 1523 2035
rect 1519 2029 1523 2030
rect 1575 2034 1579 2035
rect 1575 2029 1579 2030
rect 1615 2034 1619 2035
rect 1615 2029 1619 2030
rect 1663 2034 1667 2035
rect 1663 2029 1667 2030
rect 1719 2034 1723 2035
rect 1719 2029 1723 2030
rect 1767 2034 1771 2035
rect 1767 2029 1771 2030
rect 1823 2034 1827 2035
rect 1823 2029 1827 2030
rect 1879 2034 1883 2035
rect 1879 2029 1883 2030
rect 1935 2034 1939 2035
rect 1935 2029 1939 2030
rect 2007 2034 2011 2035
rect 2007 2029 2011 2030
rect 2055 2034 2059 2035
rect 2055 2029 2059 2030
rect 2151 2034 2155 2035
rect 2151 2029 2155 2030
rect 2183 2034 2187 2035
rect 2183 2029 2187 2030
rect 2303 2034 2307 2035
rect 2303 2029 2307 2030
rect 2319 2034 2323 2035
rect 2319 2029 2323 2030
rect 2439 2034 2443 2035
rect 2439 2029 2443 2030
rect 2503 2034 2507 2035
rect 2503 2029 2507 2030
rect 1328 2026 1330 2029
rect 1350 2028 1356 2029
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1350 2024 1351 2028
rect 1355 2024 1356 2028
rect 1350 2023 1356 2024
rect 1422 2028 1428 2029
rect 1422 2024 1423 2028
rect 1427 2024 1428 2028
rect 1422 2023 1428 2024
rect 1518 2028 1524 2029
rect 1518 2024 1519 2028
rect 1523 2024 1524 2028
rect 1518 2023 1524 2024
rect 1614 2028 1620 2029
rect 1614 2024 1615 2028
rect 1619 2024 1620 2028
rect 1614 2023 1620 2024
rect 1718 2028 1724 2029
rect 1718 2024 1719 2028
rect 1723 2024 1724 2028
rect 1718 2023 1724 2024
rect 1822 2028 1828 2029
rect 1822 2024 1823 2028
rect 1827 2024 1828 2028
rect 1822 2023 1828 2024
rect 1934 2028 1940 2029
rect 1934 2024 1935 2028
rect 1939 2024 1940 2028
rect 1934 2023 1940 2024
rect 2054 2028 2060 2029
rect 2054 2024 2055 2028
rect 2059 2024 2060 2028
rect 2054 2023 2060 2024
rect 2182 2028 2188 2029
rect 2182 2024 2183 2028
rect 2187 2024 2188 2028
rect 2182 2023 2188 2024
rect 2318 2028 2324 2029
rect 2318 2024 2319 2028
rect 2323 2024 2324 2028
rect 2318 2023 2324 2024
rect 2438 2028 2444 2029
rect 2438 2024 2439 2028
rect 2443 2024 2444 2028
rect 2504 2026 2506 2029
rect 2438 2023 2444 2024
rect 2502 2025 2508 2026
rect 1326 2020 1332 2021
rect 2502 2021 2503 2025
rect 2507 2021 2508 2025
rect 2502 2020 2508 2021
rect 1062 2013 1063 2017
rect 1067 2013 1068 2017
rect 1062 2012 1068 2013
rect 1286 2016 1292 2017
rect 1286 2012 1287 2016
rect 1291 2012 1292 2016
rect 110 2011 116 2012
rect 1286 2011 1292 2012
rect 1326 2008 1332 2009
rect 2502 2008 2508 2009
rect 1326 2004 1327 2008
rect 1331 2004 1332 2008
rect 1326 2003 1332 2004
rect 1366 2007 1372 2008
rect 1366 2003 1367 2007
rect 1371 2003 1372 2007
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1286 1999 1292 2000
rect 110 1994 116 1995
rect 278 1996 284 1997
rect 112 1987 114 1994
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 358 1996 364 1997
rect 358 1992 359 1996
rect 363 1992 364 1996
rect 358 1991 364 1992
rect 446 1996 452 1997
rect 446 1992 447 1996
rect 451 1992 452 1996
rect 446 1991 452 1992
rect 534 1996 540 1997
rect 534 1992 535 1996
rect 539 1992 540 1996
rect 534 1991 540 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 702 1996 708 1997
rect 702 1992 703 1996
rect 707 1992 708 1996
rect 702 1991 708 1992
rect 782 1996 788 1997
rect 782 1992 783 1996
rect 787 1992 788 1996
rect 782 1991 788 1992
rect 870 1996 876 1997
rect 870 1992 871 1996
rect 875 1992 876 1996
rect 870 1991 876 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1286 1995 1287 1999
rect 1291 1995 1292 1999
rect 1286 1994 1292 1995
rect 1046 1991 1052 1992
rect 280 1987 282 1991
rect 360 1987 362 1991
rect 448 1987 450 1991
rect 536 1987 538 1991
rect 624 1987 626 1991
rect 704 1987 706 1991
rect 784 1987 786 1991
rect 872 1987 874 1991
rect 960 1987 962 1991
rect 1048 1987 1050 1991
rect 1288 1987 1290 1994
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 135 1986 139 1987
rect 135 1981 139 1982
rect 207 1986 211 1987
rect 207 1981 211 1982
rect 279 1986 283 1987
rect 279 1981 283 1982
rect 287 1986 291 1987
rect 287 1981 291 1982
rect 359 1986 363 1987
rect 359 1981 363 1982
rect 383 1986 387 1987
rect 383 1981 387 1982
rect 447 1986 451 1987
rect 447 1981 451 1982
rect 487 1986 491 1987
rect 487 1981 491 1982
rect 535 1986 539 1987
rect 535 1981 539 1982
rect 591 1986 595 1987
rect 591 1981 595 1982
rect 623 1986 627 1987
rect 623 1981 627 1982
rect 695 1986 699 1987
rect 695 1981 699 1982
rect 703 1986 707 1987
rect 703 1981 707 1982
rect 783 1986 787 1987
rect 783 1981 787 1982
rect 799 1986 803 1987
rect 799 1981 803 1982
rect 871 1986 875 1987
rect 871 1981 875 1982
rect 903 1986 907 1987
rect 903 1981 907 1982
rect 959 1986 963 1987
rect 959 1981 963 1982
rect 1015 1986 1019 1987
rect 1015 1981 1019 1982
rect 1047 1986 1051 1987
rect 1047 1981 1051 1982
rect 1287 1986 1291 1987
rect 1287 1981 1291 1982
rect 112 1978 114 1981
rect 134 1980 140 1981
rect 110 1977 116 1978
rect 110 1973 111 1977
rect 115 1973 116 1977
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 206 1980 212 1981
rect 206 1976 207 1980
rect 211 1976 212 1980
rect 206 1975 212 1976
rect 286 1980 292 1981
rect 286 1976 287 1980
rect 291 1976 292 1980
rect 286 1975 292 1976
rect 382 1980 388 1981
rect 382 1976 383 1980
rect 387 1976 388 1980
rect 382 1975 388 1976
rect 486 1980 492 1981
rect 486 1976 487 1980
rect 491 1976 492 1980
rect 486 1975 492 1976
rect 590 1980 596 1981
rect 590 1976 591 1980
rect 595 1976 596 1980
rect 590 1975 596 1976
rect 694 1980 700 1981
rect 694 1976 695 1980
rect 699 1976 700 1980
rect 694 1975 700 1976
rect 798 1980 804 1981
rect 798 1976 799 1980
rect 803 1976 804 1980
rect 798 1975 804 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1014 1980 1020 1981
rect 1014 1976 1015 1980
rect 1019 1976 1020 1980
rect 1288 1978 1290 1981
rect 1328 1979 1330 2003
rect 1366 2002 1372 2003
rect 1438 2007 1444 2008
rect 1438 2003 1439 2007
rect 1443 2003 1444 2007
rect 1438 2002 1444 2003
rect 1534 2007 1540 2008
rect 1534 2003 1535 2007
rect 1539 2003 1540 2007
rect 1534 2002 1540 2003
rect 1630 2007 1636 2008
rect 1630 2003 1631 2007
rect 1635 2003 1636 2007
rect 1630 2002 1636 2003
rect 1734 2007 1740 2008
rect 1734 2003 1735 2007
rect 1739 2003 1740 2007
rect 1734 2002 1740 2003
rect 1838 2007 1844 2008
rect 1838 2003 1839 2007
rect 1843 2003 1844 2007
rect 1838 2002 1844 2003
rect 1950 2007 1956 2008
rect 1950 2003 1951 2007
rect 1955 2003 1956 2007
rect 1950 2002 1956 2003
rect 2070 2007 2076 2008
rect 2070 2003 2071 2007
rect 2075 2003 2076 2007
rect 2070 2002 2076 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2334 2007 2340 2008
rect 2334 2003 2335 2007
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2454 2007 2460 2008
rect 2454 2003 2455 2007
rect 2459 2003 2460 2007
rect 2502 2004 2503 2008
rect 2507 2004 2508 2008
rect 2502 2003 2508 2004
rect 2454 2002 2460 2003
rect 1368 1979 1370 2002
rect 1440 1979 1442 2002
rect 1536 1979 1538 2002
rect 1632 1979 1634 2002
rect 1736 1979 1738 2002
rect 1840 1979 1842 2002
rect 1952 1979 1954 2002
rect 2072 1979 2074 2002
rect 2200 1979 2202 2002
rect 2336 1979 2338 2002
rect 2456 1979 2458 2002
rect 2504 1979 2506 2003
rect 1327 1978 1331 1979
rect 1014 1975 1020 1976
rect 1286 1977 1292 1978
rect 110 1972 116 1973
rect 1286 1973 1287 1977
rect 1291 1973 1292 1977
rect 1327 1973 1331 1974
rect 1367 1978 1371 1979
rect 1367 1973 1371 1974
rect 1439 1978 1443 1979
rect 1439 1973 1443 1974
rect 1455 1978 1459 1979
rect 1455 1973 1459 1974
rect 1535 1978 1539 1979
rect 1535 1973 1539 1974
rect 1543 1978 1547 1979
rect 1543 1973 1547 1974
rect 1631 1978 1635 1979
rect 1631 1973 1635 1974
rect 1639 1978 1643 1979
rect 1639 1973 1643 1974
rect 1735 1978 1739 1979
rect 1735 1973 1739 1974
rect 1839 1978 1843 1979
rect 1839 1973 1843 1974
rect 1943 1978 1947 1979
rect 1943 1973 1947 1974
rect 1951 1978 1955 1979
rect 1951 1973 1955 1974
rect 2047 1978 2051 1979
rect 2047 1973 2051 1974
rect 2071 1978 2075 1979
rect 2071 1973 2075 1974
rect 2151 1978 2155 1979
rect 2151 1973 2155 1974
rect 2199 1978 2203 1979
rect 2199 1973 2203 1974
rect 2255 1978 2259 1979
rect 2255 1973 2259 1974
rect 2335 1978 2339 1979
rect 2335 1973 2339 1974
rect 2367 1978 2371 1979
rect 2367 1973 2371 1974
rect 2455 1978 2459 1979
rect 2455 1973 2459 1974
rect 2503 1978 2507 1979
rect 2503 1973 2507 1974
rect 1286 1972 1292 1973
rect 110 1960 116 1961
rect 1286 1960 1292 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 110 1955 116 1956
rect 150 1959 156 1960
rect 150 1955 151 1959
rect 155 1955 156 1959
rect 112 1927 114 1955
rect 150 1954 156 1955
rect 222 1959 228 1960
rect 222 1955 223 1959
rect 227 1955 228 1959
rect 222 1954 228 1955
rect 302 1959 308 1960
rect 302 1955 303 1959
rect 307 1955 308 1959
rect 302 1954 308 1955
rect 398 1959 404 1960
rect 398 1955 399 1959
rect 403 1955 404 1959
rect 398 1954 404 1955
rect 502 1959 508 1960
rect 502 1955 503 1959
rect 507 1955 508 1959
rect 502 1954 508 1955
rect 606 1959 612 1960
rect 606 1955 607 1959
rect 611 1955 612 1959
rect 606 1954 612 1955
rect 710 1959 716 1960
rect 710 1955 711 1959
rect 715 1955 716 1959
rect 710 1954 716 1955
rect 814 1959 820 1960
rect 814 1955 815 1959
rect 819 1955 820 1959
rect 814 1954 820 1955
rect 918 1959 924 1960
rect 918 1955 919 1959
rect 923 1955 924 1959
rect 918 1954 924 1955
rect 1030 1959 1036 1960
rect 1030 1955 1031 1959
rect 1035 1955 1036 1959
rect 1286 1956 1287 1960
rect 1291 1956 1292 1960
rect 1286 1955 1292 1956
rect 1030 1954 1036 1955
rect 152 1927 154 1954
rect 224 1927 226 1954
rect 304 1927 306 1954
rect 400 1927 402 1954
rect 504 1927 506 1954
rect 608 1927 610 1954
rect 712 1927 714 1954
rect 816 1927 818 1954
rect 920 1927 922 1954
rect 1032 1927 1034 1954
rect 1288 1927 1290 1955
rect 1328 1953 1330 1973
rect 1456 1954 1458 1973
rect 1544 1954 1546 1973
rect 1640 1954 1642 1973
rect 1736 1954 1738 1973
rect 1840 1954 1842 1973
rect 1944 1954 1946 1973
rect 2048 1954 2050 1973
rect 2152 1954 2154 1973
rect 2256 1954 2258 1973
rect 2368 1954 2370 1973
rect 2456 1954 2458 1973
rect 1454 1953 1460 1954
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1542 1953 1548 1954
rect 1542 1949 1543 1953
rect 1547 1949 1548 1953
rect 1542 1948 1548 1949
rect 1638 1953 1644 1954
rect 1638 1949 1639 1953
rect 1643 1949 1644 1953
rect 1638 1948 1644 1949
rect 1734 1953 1740 1954
rect 1734 1949 1735 1953
rect 1739 1949 1740 1953
rect 1734 1948 1740 1949
rect 1838 1953 1844 1954
rect 1838 1949 1839 1953
rect 1843 1949 1844 1953
rect 1838 1948 1844 1949
rect 1942 1953 1948 1954
rect 1942 1949 1943 1953
rect 1947 1949 1948 1953
rect 1942 1948 1948 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2046 1948 2052 1949
rect 2150 1953 2156 1954
rect 2150 1949 2151 1953
rect 2155 1949 2156 1953
rect 2150 1948 2156 1949
rect 2254 1953 2260 1954
rect 2254 1949 2255 1953
rect 2259 1949 2260 1953
rect 2254 1948 2260 1949
rect 2366 1953 2372 1954
rect 2366 1949 2367 1953
rect 2371 1949 2372 1953
rect 2366 1948 2372 1949
rect 2454 1953 2460 1954
rect 2504 1953 2506 1973
rect 2454 1949 2455 1953
rect 2459 1949 2460 1953
rect 2454 1948 2460 1949
rect 2502 1952 2508 1953
rect 2502 1948 2503 1952
rect 2507 1948 2508 1952
rect 1326 1947 1332 1948
rect 2502 1947 2508 1948
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 2502 1935 2508 1936
rect 1326 1930 1332 1931
rect 1438 1932 1444 1933
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 151 1926 155 1927
rect 151 1921 155 1922
rect 223 1926 227 1927
rect 223 1921 227 1922
rect 239 1926 243 1927
rect 239 1921 243 1922
rect 303 1926 307 1927
rect 303 1921 307 1922
rect 375 1926 379 1927
rect 375 1921 379 1922
rect 399 1926 403 1927
rect 399 1921 403 1922
rect 503 1926 507 1927
rect 503 1921 507 1922
rect 527 1926 531 1927
rect 527 1921 531 1922
rect 607 1926 611 1927
rect 607 1921 611 1922
rect 687 1926 691 1927
rect 687 1921 691 1922
rect 711 1926 715 1927
rect 711 1921 715 1922
rect 815 1926 819 1927
rect 815 1921 819 1922
rect 863 1926 867 1927
rect 863 1921 867 1922
rect 919 1926 923 1927
rect 919 1921 923 1922
rect 1031 1926 1035 1927
rect 1031 1921 1035 1922
rect 1039 1926 1043 1927
rect 1039 1921 1043 1922
rect 1287 1926 1291 1927
rect 1328 1923 1330 1930
rect 1438 1928 1439 1932
rect 1443 1928 1444 1932
rect 1438 1927 1444 1928
rect 1526 1932 1532 1933
rect 1526 1928 1527 1932
rect 1531 1928 1532 1932
rect 1526 1927 1532 1928
rect 1622 1932 1628 1933
rect 1622 1928 1623 1932
rect 1627 1928 1628 1932
rect 1622 1927 1628 1928
rect 1718 1932 1724 1933
rect 1718 1928 1719 1932
rect 1723 1928 1724 1932
rect 1718 1927 1724 1928
rect 1822 1932 1828 1933
rect 1822 1928 1823 1932
rect 1827 1928 1828 1932
rect 1822 1927 1828 1928
rect 1926 1932 1932 1933
rect 1926 1928 1927 1932
rect 1931 1928 1932 1932
rect 1926 1927 1932 1928
rect 2030 1932 2036 1933
rect 2030 1928 2031 1932
rect 2035 1928 2036 1932
rect 2030 1927 2036 1928
rect 2134 1932 2140 1933
rect 2134 1928 2135 1932
rect 2139 1928 2140 1932
rect 2134 1927 2140 1928
rect 2238 1932 2244 1933
rect 2238 1928 2239 1932
rect 2243 1928 2244 1932
rect 2238 1927 2244 1928
rect 2350 1932 2356 1933
rect 2350 1928 2351 1932
rect 2355 1928 2356 1932
rect 2350 1927 2356 1928
rect 2438 1932 2444 1933
rect 2438 1928 2439 1932
rect 2443 1928 2444 1932
rect 2502 1931 2503 1935
rect 2507 1931 2508 1935
rect 2502 1930 2508 1931
rect 2438 1927 2444 1928
rect 1440 1923 1442 1927
rect 1528 1923 1530 1927
rect 1624 1923 1626 1927
rect 1720 1923 1722 1927
rect 1824 1923 1826 1927
rect 1928 1923 1930 1927
rect 2032 1923 2034 1927
rect 2136 1923 2138 1927
rect 2240 1923 2242 1927
rect 2352 1923 2354 1927
rect 2440 1923 2442 1927
rect 2504 1923 2506 1930
rect 1287 1921 1291 1922
rect 1327 1922 1331 1923
rect 112 1901 114 1921
rect 152 1902 154 1921
rect 240 1902 242 1921
rect 376 1902 378 1921
rect 528 1902 530 1921
rect 688 1902 690 1921
rect 864 1902 866 1921
rect 1040 1902 1042 1921
rect 150 1901 156 1902
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 150 1897 151 1901
rect 155 1897 156 1901
rect 150 1896 156 1897
rect 238 1901 244 1902
rect 238 1897 239 1901
rect 243 1897 244 1901
rect 238 1896 244 1897
rect 374 1901 380 1902
rect 374 1897 375 1901
rect 379 1897 380 1901
rect 374 1896 380 1897
rect 526 1901 532 1902
rect 526 1897 527 1901
rect 531 1897 532 1901
rect 526 1896 532 1897
rect 686 1901 692 1902
rect 686 1897 687 1901
rect 691 1897 692 1901
rect 686 1896 692 1897
rect 862 1901 868 1902
rect 862 1897 863 1901
rect 867 1897 868 1901
rect 862 1896 868 1897
rect 1038 1901 1044 1902
rect 1288 1901 1290 1921
rect 1327 1917 1331 1918
rect 1439 1922 1443 1923
rect 1439 1917 1443 1918
rect 1527 1922 1531 1923
rect 1527 1917 1531 1918
rect 1615 1922 1619 1923
rect 1615 1917 1619 1918
rect 1623 1922 1627 1923
rect 1623 1917 1627 1918
rect 1711 1922 1715 1923
rect 1711 1917 1715 1918
rect 1719 1922 1723 1923
rect 1719 1917 1723 1918
rect 1815 1922 1819 1923
rect 1815 1917 1819 1918
rect 1823 1922 1827 1923
rect 1823 1917 1827 1918
rect 1919 1922 1923 1923
rect 1919 1917 1923 1918
rect 1927 1922 1931 1923
rect 1927 1917 1931 1918
rect 2015 1922 2019 1923
rect 2015 1917 2019 1918
rect 2031 1922 2035 1923
rect 2031 1917 2035 1918
rect 2111 1922 2115 1923
rect 2111 1917 2115 1918
rect 2135 1922 2139 1923
rect 2135 1917 2139 1918
rect 2199 1922 2203 1923
rect 2199 1917 2203 1918
rect 2239 1922 2243 1923
rect 2239 1917 2243 1918
rect 2287 1922 2291 1923
rect 2287 1917 2291 1918
rect 2351 1922 2355 1923
rect 2351 1917 2355 1918
rect 2375 1922 2379 1923
rect 2375 1917 2379 1918
rect 2439 1922 2443 1923
rect 2439 1917 2443 1918
rect 2503 1922 2507 1923
rect 2503 1917 2507 1918
rect 1328 1914 1330 1917
rect 1526 1916 1532 1917
rect 1326 1913 1332 1914
rect 1326 1909 1327 1913
rect 1331 1909 1332 1913
rect 1526 1912 1527 1916
rect 1531 1912 1532 1916
rect 1526 1911 1532 1912
rect 1614 1916 1620 1917
rect 1614 1912 1615 1916
rect 1619 1912 1620 1916
rect 1614 1911 1620 1912
rect 1710 1916 1716 1917
rect 1710 1912 1711 1916
rect 1715 1912 1716 1916
rect 1710 1911 1716 1912
rect 1814 1916 1820 1917
rect 1814 1912 1815 1916
rect 1819 1912 1820 1916
rect 1814 1911 1820 1912
rect 1918 1916 1924 1917
rect 1918 1912 1919 1916
rect 1923 1912 1924 1916
rect 1918 1911 1924 1912
rect 2014 1916 2020 1917
rect 2014 1912 2015 1916
rect 2019 1912 2020 1916
rect 2014 1911 2020 1912
rect 2110 1916 2116 1917
rect 2110 1912 2111 1916
rect 2115 1912 2116 1916
rect 2110 1911 2116 1912
rect 2198 1916 2204 1917
rect 2198 1912 2199 1916
rect 2203 1912 2204 1916
rect 2198 1911 2204 1912
rect 2286 1916 2292 1917
rect 2286 1912 2287 1916
rect 2291 1912 2292 1916
rect 2286 1911 2292 1912
rect 2374 1916 2380 1917
rect 2374 1912 2375 1916
rect 2379 1912 2380 1916
rect 2374 1911 2380 1912
rect 2438 1916 2444 1917
rect 2438 1912 2439 1916
rect 2443 1912 2444 1916
rect 2504 1914 2506 1917
rect 2438 1911 2444 1912
rect 2502 1913 2508 1914
rect 1326 1908 1332 1909
rect 2502 1909 2503 1913
rect 2507 1909 2508 1913
rect 2502 1908 2508 1909
rect 1038 1897 1039 1901
rect 1043 1897 1044 1901
rect 1038 1896 1044 1897
rect 1286 1900 1292 1901
rect 1286 1896 1287 1900
rect 1291 1896 1292 1900
rect 110 1895 116 1896
rect 1286 1895 1292 1896
rect 1326 1896 1332 1897
rect 2502 1896 2508 1897
rect 1326 1892 1327 1896
rect 1331 1892 1332 1896
rect 1326 1891 1332 1892
rect 1542 1895 1548 1896
rect 1542 1891 1543 1895
rect 1547 1891 1548 1895
rect 110 1883 116 1884
rect 110 1879 111 1883
rect 115 1879 116 1883
rect 1286 1883 1292 1884
rect 110 1878 116 1879
rect 134 1880 140 1881
rect 112 1875 114 1878
rect 134 1876 135 1880
rect 139 1876 140 1880
rect 134 1875 140 1876
rect 222 1880 228 1881
rect 222 1876 223 1880
rect 227 1876 228 1880
rect 222 1875 228 1876
rect 358 1880 364 1881
rect 358 1876 359 1880
rect 363 1876 364 1880
rect 358 1875 364 1876
rect 510 1880 516 1881
rect 510 1876 511 1880
rect 515 1876 516 1880
rect 510 1875 516 1876
rect 670 1880 676 1881
rect 670 1876 671 1880
rect 675 1876 676 1880
rect 670 1875 676 1876
rect 846 1880 852 1881
rect 846 1876 847 1880
rect 851 1876 852 1880
rect 846 1875 852 1876
rect 1022 1880 1028 1881
rect 1022 1876 1023 1880
rect 1027 1876 1028 1880
rect 1286 1879 1287 1883
rect 1291 1879 1292 1883
rect 1286 1878 1292 1879
rect 1022 1875 1028 1876
rect 1288 1875 1290 1878
rect 111 1874 115 1875
rect 111 1869 115 1870
rect 135 1874 139 1875
rect 135 1869 139 1870
rect 191 1874 195 1875
rect 191 1869 195 1870
rect 223 1874 227 1875
rect 223 1869 227 1870
rect 263 1874 267 1875
rect 263 1869 267 1870
rect 335 1874 339 1875
rect 335 1869 339 1870
rect 359 1874 363 1875
rect 359 1869 363 1870
rect 407 1874 411 1875
rect 407 1869 411 1870
rect 479 1874 483 1875
rect 479 1869 483 1870
rect 511 1874 515 1875
rect 511 1869 515 1870
rect 551 1874 555 1875
rect 551 1869 555 1870
rect 615 1874 619 1875
rect 615 1869 619 1870
rect 671 1874 675 1875
rect 671 1869 675 1870
rect 679 1874 683 1875
rect 679 1869 683 1870
rect 743 1874 747 1875
rect 743 1869 747 1870
rect 815 1874 819 1875
rect 815 1869 819 1870
rect 847 1874 851 1875
rect 847 1869 851 1870
rect 887 1874 891 1875
rect 887 1869 891 1870
rect 959 1874 963 1875
rect 959 1869 963 1870
rect 1023 1874 1027 1875
rect 1023 1869 1027 1870
rect 1039 1874 1043 1875
rect 1039 1869 1043 1870
rect 1287 1874 1291 1875
rect 1328 1871 1330 1891
rect 1542 1890 1548 1891
rect 1630 1895 1636 1896
rect 1630 1891 1631 1895
rect 1635 1891 1636 1895
rect 1630 1890 1636 1891
rect 1726 1895 1732 1896
rect 1726 1891 1727 1895
rect 1731 1891 1732 1895
rect 1726 1890 1732 1891
rect 1830 1895 1836 1896
rect 1830 1891 1831 1895
rect 1835 1891 1836 1895
rect 1830 1890 1836 1891
rect 1934 1895 1940 1896
rect 1934 1891 1935 1895
rect 1939 1891 1940 1895
rect 1934 1890 1940 1891
rect 2030 1895 2036 1896
rect 2030 1891 2031 1895
rect 2035 1891 2036 1895
rect 2030 1890 2036 1891
rect 2126 1895 2132 1896
rect 2126 1891 2127 1895
rect 2131 1891 2132 1895
rect 2126 1890 2132 1891
rect 2214 1895 2220 1896
rect 2214 1891 2215 1895
rect 2219 1891 2220 1895
rect 2214 1890 2220 1891
rect 2302 1895 2308 1896
rect 2302 1891 2303 1895
rect 2307 1891 2308 1895
rect 2302 1890 2308 1891
rect 2390 1895 2396 1896
rect 2390 1891 2391 1895
rect 2395 1891 2396 1895
rect 2390 1890 2396 1891
rect 2454 1895 2460 1896
rect 2454 1891 2455 1895
rect 2459 1891 2460 1895
rect 2502 1892 2503 1896
rect 2507 1892 2508 1896
rect 2502 1891 2508 1892
rect 2454 1890 2460 1891
rect 1544 1871 1546 1890
rect 1632 1871 1634 1890
rect 1728 1871 1730 1890
rect 1832 1871 1834 1890
rect 1936 1871 1938 1890
rect 2032 1871 2034 1890
rect 2128 1871 2130 1890
rect 2216 1871 2218 1890
rect 2304 1871 2306 1890
rect 2392 1871 2394 1890
rect 2456 1871 2458 1890
rect 2504 1871 2506 1891
rect 1287 1869 1291 1870
rect 1327 1870 1331 1871
rect 112 1866 114 1869
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 190 1868 196 1869
rect 190 1864 191 1868
rect 195 1864 196 1868
rect 190 1863 196 1864
rect 262 1868 268 1869
rect 262 1864 263 1868
rect 267 1864 268 1868
rect 262 1863 268 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 406 1868 412 1869
rect 406 1864 407 1868
rect 411 1864 412 1868
rect 406 1863 412 1864
rect 478 1868 484 1869
rect 478 1864 479 1868
rect 483 1864 484 1868
rect 478 1863 484 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 614 1868 620 1869
rect 614 1864 615 1868
rect 619 1864 620 1868
rect 614 1863 620 1864
rect 678 1868 684 1869
rect 678 1864 679 1868
rect 683 1864 684 1868
rect 678 1863 684 1864
rect 742 1868 748 1869
rect 742 1864 743 1868
rect 747 1864 748 1868
rect 742 1863 748 1864
rect 814 1868 820 1869
rect 814 1864 815 1868
rect 819 1864 820 1868
rect 814 1863 820 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 958 1868 964 1869
rect 958 1864 959 1868
rect 963 1864 964 1868
rect 958 1863 964 1864
rect 1038 1868 1044 1869
rect 1038 1864 1039 1868
rect 1043 1864 1044 1868
rect 1288 1866 1290 1869
rect 1038 1863 1044 1864
rect 1286 1865 1292 1866
rect 1327 1865 1331 1866
rect 1535 1870 1539 1871
rect 1535 1865 1539 1866
rect 1543 1870 1547 1871
rect 1543 1865 1547 1866
rect 1607 1870 1611 1871
rect 1607 1865 1611 1866
rect 1631 1870 1635 1871
rect 1631 1865 1635 1866
rect 1687 1870 1691 1871
rect 1687 1865 1691 1866
rect 1727 1870 1731 1871
rect 1727 1865 1731 1866
rect 1783 1870 1787 1871
rect 1783 1865 1787 1866
rect 1831 1870 1835 1871
rect 1831 1865 1835 1866
rect 1879 1870 1883 1871
rect 1879 1865 1883 1866
rect 1935 1870 1939 1871
rect 1935 1865 1939 1866
rect 1983 1870 1987 1871
rect 1983 1865 1987 1866
rect 2031 1870 2035 1871
rect 2031 1865 2035 1866
rect 2079 1870 2083 1871
rect 2079 1865 2083 1866
rect 2127 1870 2131 1871
rect 2127 1865 2131 1866
rect 2175 1870 2179 1871
rect 2175 1865 2179 1866
rect 2215 1870 2219 1871
rect 2215 1865 2219 1866
rect 2271 1870 2275 1871
rect 2271 1865 2275 1866
rect 2303 1870 2307 1871
rect 2303 1865 2307 1866
rect 2367 1870 2371 1871
rect 2367 1865 2371 1866
rect 2391 1870 2395 1871
rect 2391 1865 2395 1866
rect 2455 1870 2459 1871
rect 2455 1865 2459 1866
rect 2503 1870 2507 1871
rect 2503 1865 2507 1866
rect 110 1860 116 1861
rect 1286 1861 1287 1865
rect 1291 1861 1292 1865
rect 1286 1860 1292 1861
rect 110 1848 116 1849
rect 1286 1848 1292 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 150 1847 156 1848
rect 150 1843 151 1847
rect 155 1843 156 1847
rect 112 1815 114 1843
rect 150 1842 156 1843
rect 206 1847 212 1848
rect 206 1843 207 1847
rect 211 1843 212 1847
rect 206 1842 212 1843
rect 278 1847 284 1848
rect 278 1843 279 1847
rect 283 1843 284 1847
rect 278 1842 284 1843
rect 350 1847 356 1848
rect 350 1843 351 1847
rect 355 1843 356 1847
rect 350 1842 356 1843
rect 422 1847 428 1848
rect 422 1843 423 1847
rect 427 1843 428 1847
rect 422 1842 428 1843
rect 494 1847 500 1848
rect 494 1843 495 1847
rect 499 1843 500 1847
rect 494 1842 500 1843
rect 566 1847 572 1848
rect 566 1843 567 1847
rect 571 1843 572 1847
rect 566 1842 572 1843
rect 630 1847 636 1848
rect 630 1843 631 1847
rect 635 1843 636 1847
rect 630 1842 636 1843
rect 694 1847 700 1848
rect 694 1843 695 1847
rect 699 1843 700 1847
rect 694 1842 700 1843
rect 758 1847 764 1848
rect 758 1843 759 1847
rect 763 1843 764 1847
rect 758 1842 764 1843
rect 830 1847 836 1848
rect 830 1843 831 1847
rect 835 1843 836 1847
rect 830 1842 836 1843
rect 902 1847 908 1848
rect 902 1843 903 1847
rect 907 1843 908 1847
rect 902 1842 908 1843
rect 974 1847 980 1848
rect 974 1843 975 1847
rect 979 1843 980 1847
rect 974 1842 980 1843
rect 1054 1847 1060 1848
rect 1054 1843 1055 1847
rect 1059 1843 1060 1847
rect 1286 1844 1287 1848
rect 1291 1844 1292 1848
rect 1328 1845 1330 1865
rect 1536 1846 1538 1865
rect 1608 1846 1610 1865
rect 1688 1846 1690 1865
rect 1784 1846 1786 1865
rect 1880 1846 1882 1865
rect 1984 1846 1986 1865
rect 2080 1846 2082 1865
rect 2176 1846 2178 1865
rect 2272 1846 2274 1865
rect 2368 1846 2370 1865
rect 2456 1846 2458 1865
rect 1534 1845 1540 1846
rect 1286 1843 1292 1844
rect 1326 1844 1332 1845
rect 1054 1842 1060 1843
rect 152 1815 154 1842
rect 208 1815 210 1842
rect 280 1815 282 1842
rect 352 1815 354 1842
rect 424 1815 426 1842
rect 496 1815 498 1842
rect 568 1815 570 1842
rect 632 1815 634 1842
rect 696 1815 698 1842
rect 760 1815 762 1842
rect 832 1815 834 1842
rect 904 1815 906 1842
rect 976 1815 978 1842
rect 1056 1815 1058 1842
rect 1288 1815 1290 1843
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1534 1841 1535 1845
rect 1539 1841 1540 1845
rect 1534 1840 1540 1841
rect 1606 1845 1612 1846
rect 1606 1841 1607 1845
rect 1611 1841 1612 1845
rect 1606 1840 1612 1841
rect 1686 1845 1692 1846
rect 1686 1841 1687 1845
rect 1691 1841 1692 1845
rect 1686 1840 1692 1841
rect 1782 1845 1788 1846
rect 1782 1841 1783 1845
rect 1787 1841 1788 1845
rect 1782 1840 1788 1841
rect 1878 1845 1884 1846
rect 1878 1841 1879 1845
rect 1883 1841 1884 1845
rect 1878 1840 1884 1841
rect 1982 1845 1988 1846
rect 1982 1841 1983 1845
rect 1987 1841 1988 1845
rect 1982 1840 1988 1841
rect 2078 1845 2084 1846
rect 2078 1841 2079 1845
rect 2083 1841 2084 1845
rect 2078 1840 2084 1841
rect 2174 1845 2180 1846
rect 2174 1841 2175 1845
rect 2179 1841 2180 1845
rect 2174 1840 2180 1841
rect 2270 1845 2276 1846
rect 2270 1841 2271 1845
rect 2275 1841 2276 1845
rect 2270 1840 2276 1841
rect 2366 1845 2372 1846
rect 2366 1841 2367 1845
rect 2371 1841 2372 1845
rect 2366 1840 2372 1841
rect 2454 1845 2460 1846
rect 2504 1845 2506 1865
rect 2454 1841 2455 1845
rect 2459 1841 2460 1845
rect 2454 1840 2460 1841
rect 2502 1844 2508 1845
rect 2502 1840 2503 1844
rect 2507 1840 2508 1844
rect 1326 1839 1332 1840
rect 2502 1839 2508 1840
rect 1326 1827 1332 1828
rect 1326 1823 1327 1827
rect 1331 1823 1332 1827
rect 2502 1827 2508 1828
rect 1326 1822 1332 1823
rect 1518 1824 1524 1825
rect 1328 1815 1330 1822
rect 1518 1820 1519 1824
rect 1523 1820 1524 1824
rect 1518 1819 1524 1820
rect 1590 1824 1596 1825
rect 1590 1820 1591 1824
rect 1595 1820 1596 1824
rect 1590 1819 1596 1820
rect 1670 1824 1676 1825
rect 1670 1820 1671 1824
rect 1675 1820 1676 1824
rect 1670 1819 1676 1820
rect 1766 1824 1772 1825
rect 1766 1820 1767 1824
rect 1771 1820 1772 1824
rect 1766 1819 1772 1820
rect 1862 1824 1868 1825
rect 1862 1820 1863 1824
rect 1867 1820 1868 1824
rect 1862 1819 1868 1820
rect 1966 1824 1972 1825
rect 1966 1820 1967 1824
rect 1971 1820 1972 1824
rect 1966 1819 1972 1820
rect 2062 1824 2068 1825
rect 2062 1820 2063 1824
rect 2067 1820 2068 1824
rect 2062 1819 2068 1820
rect 2158 1824 2164 1825
rect 2158 1820 2159 1824
rect 2163 1820 2164 1824
rect 2158 1819 2164 1820
rect 2254 1824 2260 1825
rect 2254 1820 2255 1824
rect 2259 1820 2260 1824
rect 2254 1819 2260 1820
rect 2350 1824 2356 1825
rect 2350 1820 2351 1824
rect 2355 1820 2356 1824
rect 2350 1819 2356 1820
rect 2438 1824 2444 1825
rect 2438 1820 2439 1824
rect 2443 1820 2444 1824
rect 2502 1823 2503 1827
rect 2507 1823 2508 1827
rect 2502 1822 2508 1823
rect 2438 1819 2444 1820
rect 1520 1815 1522 1819
rect 1592 1815 1594 1819
rect 1672 1815 1674 1819
rect 1768 1815 1770 1819
rect 1864 1815 1866 1819
rect 1968 1815 1970 1819
rect 2064 1815 2066 1819
rect 2160 1815 2162 1819
rect 2256 1815 2258 1819
rect 2352 1815 2354 1819
rect 2440 1815 2442 1819
rect 2504 1815 2506 1822
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 151 1814 155 1815
rect 151 1809 155 1810
rect 207 1814 211 1815
rect 207 1809 211 1810
rect 231 1814 235 1815
rect 231 1809 235 1810
rect 279 1814 283 1815
rect 279 1809 283 1810
rect 335 1814 339 1815
rect 335 1809 339 1810
rect 351 1814 355 1815
rect 351 1809 355 1810
rect 423 1814 427 1815
rect 423 1809 427 1810
rect 439 1814 443 1815
rect 439 1809 443 1810
rect 495 1814 499 1815
rect 495 1809 499 1810
rect 535 1814 539 1815
rect 535 1809 539 1810
rect 567 1814 571 1815
rect 567 1809 571 1810
rect 631 1814 635 1815
rect 631 1809 635 1810
rect 695 1814 699 1815
rect 695 1809 699 1810
rect 719 1814 723 1815
rect 719 1809 723 1810
rect 759 1814 763 1815
rect 759 1809 763 1810
rect 799 1814 803 1815
rect 799 1809 803 1810
rect 831 1814 835 1815
rect 831 1809 835 1810
rect 879 1814 883 1815
rect 879 1809 883 1810
rect 903 1814 907 1815
rect 903 1809 907 1810
rect 959 1814 963 1815
rect 959 1809 963 1810
rect 975 1814 979 1815
rect 975 1809 979 1810
rect 1039 1814 1043 1815
rect 1039 1809 1043 1810
rect 1055 1814 1059 1815
rect 1055 1809 1059 1810
rect 1119 1814 1123 1815
rect 1119 1809 1123 1810
rect 1287 1814 1291 1815
rect 1287 1809 1291 1810
rect 1327 1814 1331 1815
rect 1327 1809 1331 1810
rect 1463 1814 1467 1815
rect 1463 1809 1467 1810
rect 1519 1814 1523 1815
rect 1519 1809 1523 1810
rect 1559 1814 1563 1815
rect 1559 1809 1563 1810
rect 1591 1814 1595 1815
rect 1591 1809 1595 1810
rect 1663 1814 1667 1815
rect 1663 1809 1667 1810
rect 1671 1814 1675 1815
rect 1671 1809 1675 1810
rect 1767 1814 1771 1815
rect 1767 1809 1771 1810
rect 1863 1814 1867 1815
rect 1863 1809 1867 1810
rect 1879 1814 1883 1815
rect 1879 1809 1883 1810
rect 1967 1814 1971 1815
rect 1967 1809 1971 1810
rect 1983 1814 1987 1815
rect 1983 1809 1987 1810
rect 2063 1814 2067 1815
rect 2063 1809 2067 1810
rect 2087 1814 2091 1815
rect 2087 1809 2091 1810
rect 2159 1814 2163 1815
rect 2159 1809 2163 1810
rect 2183 1814 2187 1815
rect 2183 1809 2187 1810
rect 2255 1814 2259 1815
rect 2255 1809 2259 1810
rect 2271 1814 2275 1815
rect 2271 1809 2275 1810
rect 2351 1814 2355 1815
rect 2351 1809 2355 1810
rect 2367 1814 2371 1815
rect 2367 1809 2371 1810
rect 2439 1814 2443 1815
rect 2439 1809 2443 1810
rect 2503 1814 2507 1815
rect 2503 1809 2507 1810
rect 112 1789 114 1809
rect 152 1790 154 1809
rect 232 1790 234 1809
rect 336 1790 338 1809
rect 440 1790 442 1809
rect 536 1790 538 1809
rect 632 1790 634 1809
rect 720 1790 722 1809
rect 800 1790 802 1809
rect 880 1790 882 1809
rect 960 1790 962 1809
rect 1040 1790 1042 1809
rect 1120 1790 1122 1809
rect 150 1789 156 1790
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 150 1785 151 1789
rect 155 1785 156 1789
rect 150 1784 156 1785
rect 230 1789 236 1790
rect 230 1785 231 1789
rect 235 1785 236 1789
rect 230 1784 236 1785
rect 334 1789 340 1790
rect 334 1785 335 1789
rect 339 1785 340 1789
rect 334 1784 340 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 534 1789 540 1790
rect 534 1785 535 1789
rect 539 1785 540 1789
rect 534 1784 540 1785
rect 630 1789 636 1790
rect 630 1785 631 1789
rect 635 1785 636 1789
rect 630 1784 636 1785
rect 718 1789 724 1790
rect 718 1785 719 1789
rect 723 1785 724 1789
rect 718 1784 724 1785
rect 798 1789 804 1790
rect 798 1785 799 1789
rect 803 1785 804 1789
rect 798 1784 804 1785
rect 878 1789 884 1790
rect 878 1785 879 1789
rect 883 1785 884 1789
rect 878 1784 884 1785
rect 958 1789 964 1790
rect 958 1785 959 1789
rect 963 1785 964 1789
rect 958 1784 964 1785
rect 1038 1789 1044 1790
rect 1038 1785 1039 1789
rect 1043 1785 1044 1789
rect 1038 1784 1044 1785
rect 1118 1789 1124 1790
rect 1288 1789 1290 1809
rect 1328 1806 1330 1809
rect 1462 1808 1468 1809
rect 1326 1805 1332 1806
rect 1326 1801 1327 1805
rect 1331 1801 1332 1805
rect 1462 1804 1463 1808
rect 1467 1804 1468 1808
rect 1462 1803 1468 1804
rect 1558 1808 1564 1809
rect 1558 1804 1559 1808
rect 1563 1804 1564 1808
rect 1558 1803 1564 1804
rect 1662 1808 1668 1809
rect 1662 1804 1663 1808
rect 1667 1804 1668 1808
rect 1662 1803 1668 1804
rect 1766 1808 1772 1809
rect 1766 1804 1767 1808
rect 1771 1804 1772 1808
rect 1766 1803 1772 1804
rect 1878 1808 1884 1809
rect 1878 1804 1879 1808
rect 1883 1804 1884 1808
rect 1878 1803 1884 1804
rect 1982 1808 1988 1809
rect 1982 1804 1983 1808
rect 1987 1804 1988 1808
rect 1982 1803 1988 1804
rect 2086 1808 2092 1809
rect 2086 1804 2087 1808
rect 2091 1804 2092 1808
rect 2086 1803 2092 1804
rect 2182 1808 2188 1809
rect 2182 1804 2183 1808
rect 2187 1804 2188 1808
rect 2182 1803 2188 1804
rect 2270 1808 2276 1809
rect 2270 1804 2271 1808
rect 2275 1804 2276 1808
rect 2270 1803 2276 1804
rect 2366 1808 2372 1809
rect 2366 1804 2367 1808
rect 2371 1804 2372 1808
rect 2366 1803 2372 1804
rect 2438 1808 2444 1809
rect 2438 1804 2439 1808
rect 2443 1804 2444 1808
rect 2504 1806 2506 1809
rect 2438 1803 2444 1804
rect 2502 1805 2508 1806
rect 1326 1800 1332 1801
rect 2502 1801 2503 1805
rect 2507 1801 2508 1805
rect 2502 1800 2508 1801
rect 1118 1785 1119 1789
rect 1123 1785 1124 1789
rect 1118 1784 1124 1785
rect 1286 1788 1292 1789
rect 1286 1784 1287 1788
rect 1291 1784 1292 1788
rect 110 1783 116 1784
rect 1286 1783 1292 1784
rect 1326 1788 1332 1789
rect 2502 1788 2508 1789
rect 1326 1784 1327 1788
rect 1331 1784 1332 1788
rect 1326 1783 1332 1784
rect 1478 1787 1484 1788
rect 1478 1783 1479 1787
rect 1483 1783 1484 1787
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1286 1771 1292 1772
rect 110 1766 116 1767
rect 134 1768 140 1769
rect 112 1759 114 1766
rect 134 1764 135 1768
rect 139 1764 140 1768
rect 134 1763 140 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 318 1768 324 1769
rect 318 1764 319 1768
rect 323 1764 324 1768
rect 318 1763 324 1764
rect 422 1768 428 1769
rect 422 1764 423 1768
rect 427 1764 428 1768
rect 422 1763 428 1764
rect 518 1768 524 1769
rect 518 1764 519 1768
rect 523 1764 524 1768
rect 518 1763 524 1764
rect 614 1768 620 1769
rect 614 1764 615 1768
rect 619 1764 620 1768
rect 614 1763 620 1764
rect 702 1768 708 1769
rect 702 1764 703 1768
rect 707 1764 708 1768
rect 702 1763 708 1764
rect 782 1768 788 1769
rect 782 1764 783 1768
rect 787 1764 788 1768
rect 782 1763 788 1764
rect 862 1768 868 1769
rect 862 1764 863 1768
rect 867 1764 868 1768
rect 862 1763 868 1764
rect 942 1768 948 1769
rect 942 1764 943 1768
rect 947 1764 948 1768
rect 942 1763 948 1764
rect 1022 1768 1028 1769
rect 1022 1764 1023 1768
rect 1027 1764 1028 1768
rect 1022 1763 1028 1764
rect 1102 1768 1108 1769
rect 1102 1764 1103 1768
rect 1107 1764 1108 1768
rect 1286 1767 1287 1771
rect 1291 1767 1292 1771
rect 1286 1766 1292 1767
rect 1102 1763 1108 1764
rect 136 1759 138 1763
rect 216 1759 218 1763
rect 320 1759 322 1763
rect 424 1759 426 1763
rect 520 1759 522 1763
rect 616 1759 618 1763
rect 704 1759 706 1763
rect 784 1759 786 1763
rect 864 1759 866 1763
rect 944 1759 946 1763
rect 1024 1759 1026 1763
rect 1104 1759 1106 1763
rect 1288 1759 1290 1766
rect 1328 1759 1330 1783
rect 1478 1782 1484 1783
rect 1574 1787 1580 1788
rect 1574 1783 1575 1787
rect 1579 1783 1580 1787
rect 1574 1782 1580 1783
rect 1678 1787 1684 1788
rect 1678 1783 1679 1787
rect 1683 1783 1684 1787
rect 1678 1782 1684 1783
rect 1782 1787 1788 1788
rect 1782 1783 1783 1787
rect 1787 1783 1788 1787
rect 1782 1782 1788 1783
rect 1894 1787 1900 1788
rect 1894 1783 1895 1787
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1998 1787 2004 1788
rect 1998 1783 1999 1787
rect 2003 1783 2004 1787
rect 1998 1782 2004 1783
rect 2102 1787 2108 1788
rect 2102 1783 2103 1787
rect 2107 1783 2108 1787
rect 2102 1782 2108 1783
rect 2198 1787 2204 1788
rect 2198 1783 2199 1787
rect 2203 1783 2204 1787
rect 2198 1782 2204 1783
rect 2286 1787 2292 1788
rect 2286 1783 2287 1787
rect 2291 1783 2292 1787
rect 2286 1782 2292 1783
rect 2382 1787 2388 1788
rect 2382 1783 2383 1787
rect 2387 1783 2388 1787
rect 2382 1782 2388 1783
rect 2454 1787 2460 1788
rect 2454 1783 2455 1787
rect 2459 1783 2460 1787
rect 2502 1784 2503 1788
rect 2507 1784 2508 1788
rect 2502 1783 2508 1784
rect 2454 1782 2460 1783
rect 1480 1759 1482 1782
rect 1576 1759 1578 1782
rect 1680 1759 1682 1782
rect 1784 1759 1786 1782
rect 1896 1759 1898 1782
rect 2000 1759 2002 1782
rect 2104 1759 2106 1782
rect 2200 1759 2202 1782
rect 2288 1759 2290 1782
rect 2384 1759 2386 1782
rect 2456 1759 2458 1782
rect 2504 1759 2506 1783
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 135 1758 139 1759
rect 135 1753 139 1754
rect 215 1758 219 1759
rect 215 1753 219 1754
rect 239 1758 243 1759
rect 239 1753 243 1754
rect 319 1758 323 1759
rect 319 1753 323 1754
rect 351 1758 355 1759
rect 351 1753 355 1754
rect 423 1758 427 1759
rect 423 1753 427 1754
rect 463 1758 467 1759
rect 463 1753 467 1754
rect 519 1758 523 1759
rect 519 1753 523 1754
rect 575 1758 579 1759
rect 575 1753 579 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 679 1758 683 1759
rect 679 1753 683 1754
rect 703 1758 707 1759
rect 703 1753 707 1754
rect 783 1758 787 1759
rect 783 1753 787 1754
rect 863 1758 867 1759
rect 863 1753 867 1754
rect 887 1758 891 1759
rect 887 1753 891 1754
rect 943 1758 947 1759
rect 943 1753 947 1754
rect 991 1758 995 1759
rect 991 1753 995 1754
rect 1023 1758 1027 1759
rect 1023 1753 1027 1754
rect 1103 1758 1107 1759
rect 1103 1753 1107 1754
rect 1287 1758 1291 1759
rect 1287 1753 1291 1754
rect 1327 1758 1331 1759
rect 1327 1753 1331 1754
rect 1375 1758 1379 1759
rect 1375 1753 1379 1754
rect 1471 1758 1475 1759
rect 1471 1753 1475 1754
rect 1479 1758 1483 1759
rect 1479 1753 1483 1754
rect 1567 1758 1571 1759
rect 1567 1753 1571 1754
rect 1575 1758 1579 1759
rect 1575 1753 1579 1754
rect 1671 1758 1675 1759
rect 1671 1753 1675 1754
rect 1679 1758 1683 1759
rect 1679 1753 1683 1754
rect 1775 1758 1779 1759
rect 1775 1753 1779 1754
rect 1783 1758 1787 1759
rect 1783 1753 1787 1754
rect 1887 1758 1891 1759
rect 1887 1753 1891 1754
rect 1895 1758 1899 1759
rect 1895 1753 1899 1754
rect 1999 1758 2003 1759
rect 1999 1753 2003 1754
rect 2103 1758 2107 1759
rect 2103 1753 2107 1754
rect 2111 1758 2115 1759
rect 2111 1753 2115 1754
rect 2199 1758 2203 1759
rect 2199 1753 2203 1754
rect 2231 1758 2235 1759
rect 2231 1753 2235 1754
rect 2287 1758 2291 1759
rect 2287 1753 2291 1754
rect 2351 1758 2355 1759
rect 2351 1753 2355 1754
rect 2383 1758 2387 1759
rect 2383 1753 2387 1754
rect 2455 1758 2459 1759
rect 2455 1753 2459 1754
rect 2503 1758 2507 1759
rect 2503 1753 2507 1754
rect 112 1750 114 1753
rect 134 1752 140 1753
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 134 1748 135 1752
rect 139 1748 140 1752
rect 134 1747 140 1748
rect 238 1752 244 1753
rect 238 1748 239 1752
rect 243 1748 244 1752
rect 238 1747 244 1748
rect 350 1752 356 1753
rect 350 1748 351 1752
rect 355 1748 356 1752
rect 350 1747 356 1748
rect 462 1752 468 1753
rect 462 1748 463 1752
rect 467 1748 468 1752
rect 462 1747 468 1748
rect 574 1752 580 1753
rect 574 1748 575 1752
rect 579 1748 580 1752
rect 574 1747 580 1748
rect 678 1752 684 1753
rect 678 1748 679 1752
rect 683 1748 684 1752
rect 678 1747 684 1748
rect 782 1752 788 1753
rect 782 1748 783 1752
rect 787 1748 788 1752
rect 782 1747 788 1748
rect 886 1752 892 1753
rect 886 1748 887 1752
rect 891 1748 892 1752
rect 886 1747 892 1748
rect 990 1752 996 1753
rect 990 1748 991 1752
rect 995 1748 996 1752
rect 990 1747 996 1748
rect 1102 1752 1108 1753
rect 1102 1748 1103 1752
rect 1107 1748 1108 1752
rect 1288 1750 1290 1753
rect 1102 1747 1108 1748
rect 1286 1749 1292 1750
rect 110 1744 116 1745
rect 1286 1745 1287 1749
rect 1291 1745 1292 1749
rect 1286 1744 1292 1745
rect 1328 1733 1330 1753
rect 1376 1734 1378 1753
rect 1472 1734 1474 1753
rect 1568 1734 1570 1753
rect 1672 1734 1674 1753
rect 1776 1734 1778 1753
rect 1888 1734 1890 1753
rect 2000 1734 2002 1753
rect 2112 1734 2114 1753
rect 2232 1734 2234 1753
rect 2352 1734 2354 1753
rect 2456 1734 2458 1753
rect 1374 1733 1380 1734
rect 110 1732 116 1733
rect 1286 1732 1292 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 150 1731 156 1732
rect 150 1727 151 1731
rect 155 1727 156 1731
rect 112 1703 114 1727
rect 150 1726 156 1727
rect 254 1731 260 1732
rect 254 1727 255 1731
rect 259 1727 260 1731
rect 254 1726 260 1727
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 478 1731 484 1732
rect 478 1727 479 1731
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 590 1731 596 1732
rect 590 1727 591 1731
rect 595 1727 596 1731
rect 590 1726 596 1727
rect 694 1731 700 1732
rect 694 1727 695 1731
rect 699 1727 700 1731
rect 694 1726 700 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 902 1731 908 1732
rect 902 1727 903 1731
rect 907 1727 908 1731
rect 902 1726 908 1727
rect 1006 1731 1012 1732
rect 1006 1727 1007 1731
rect 1011 1727 1012 1731
rect 1006 1726 1012 1727
rect 1118 1731 1124 1732
rect 1118 1727 1119 1731
rect 1123 1727 1124 1731
rect 1286 1728 1287 1732
rect 1291 1728 1292 1732
rect 1286 1727 1292 1728
rect 1326 1732 1332 1733
rect 1326 1728 1327 1732
rect 1331 1728 1332 1732
rect 1374 1729 1375 1733
rect 1379 1729 1380 1733
rect 1374 1728 1380 1729
rect 1470 1733 1476 1734
rect 1470 1729 1471 1733
rect 1475 1729 1476 1733
rect 1470 1728 1476 1729
rect 1566 1733 1572 1734
rect 1566 1729 1567 1733
rect 1571 1729 1572 1733
rect 1566 1728 1572 1729
rect 1670 1733 1676 1734
rect 1670 1729 1671 1733
rect 1675 1729 1676 1733
rect 1670 1728 1676 1729
rect 1774 1733 1780 1734
rect 1774 1729 1775 1733
rect 1779 1729 1780 1733
rect 1774 1728 1780 1729
rect 1886 1733 1892 1734
rect 1886 1729 1887 1733
rect 1891 1729 1892 1733
rect 1886 1728 1892 1729
rect 1998 1733 2004 1734
rect 1998 1729 1999 1733
rect 2003 1729 2004 1733
rect 1998 1728 2004 1729
rect 2110 1733 2116 1734
rect 2110 1729 2111 1733
rect 2115 1729 2116 1733
rect 2110 1728 2116 1729
rect 2230 1733 2236 1734
rect 2230 1729 2231 1733
rect 2235 1729 2236 1733
rect 2230 1728 2236 1729
rect 2350 1733 2356 1734
rect 2350 1729 2351 1733
rect 2355 1729 2356 1733
rect 2350 1728 2356 1729
rect 2454 1733 2460 1734
rect 2504 1733 2506 1753
rect 2454 1729 2455 1733
rect 2459 1729 2460 1733
rect 2454 1728 2460 1729
rect 2502 1732 2508 1733
rect 2502 1728 2503 1732
rect 2507 1728 2508 1732
rect 1326 1727 1332 1728
rect 2502 1727 2508 1728
rect 1118 1726 1124 1727
rect 152 1703 154 1726
rect 256 1703 258 1726
rect 368 1703 370 1726
rect 480 1703 482 1726
rect 592 1703 594 1726
rect 696 1703 698 1726
rect 800 1703 802 1726
rect 904 1703 906 1726
rect 1008 1703 1010 1726
rect 1120 1703 1122 1726
rect 1288 1703 1290 1727
rect 1326 1715 1332 1716
rect 1326 1711 1327 1715
rect 1331 1711 1332 1715
rect 2502 1715 2508 1716
rect 1326 1710 1332 1711
rect 1358 1712 1364 1713
rect 1328 1707 1330 1710
rect 1358 1708 1359 1712
rect 1363 1708 1364 1712
rect 1358 1707 1364 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1550 1712 1556 1713
rect 1550 1708 1551 1712
rect 1555 1708 1556 1712
rect 1550 1707 1556 1708
rect 1654 1712 1660 1713
rect 1654 1708 1655 1712
rect 1659 1708 1660 1712
rect 1654 1707 1660 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1870 1712 1876 1713
rect 1870 1708 1871 1712
rect 1875 1708 1876 1712
rect 1870 1707 1876 1708
rect 1982 1712 1988 1713
rect 1982 1708 1983 1712
rect 1987 1708 1988 1712
rect 1982 1707 1988 1708
rect 2094 1712 2100 1713
rect 2094 1708 2095 1712
rect 2099 1708 2100 1712
rect 2094 1707 2100 1708
rect 2214 1712 2220 1713
rect 2214 1708 2215 1712
rect 2219 1708 2220 1712
rect 2214 1707 2220 1708
rect 2334 1712 2340 1713
rect 2334 1708 2335 1712
rect 2339 1708 2340 1712
rect 2334 1707 2340 1708
rect 2438 1712 2444 1713
rect 2438 1708 2439 1712
rect 2443 1708 2444 1712
rect 2502 1711 2503 1715
rect 2507 1711 2508 1715
rect 2502 1710 2508 1711
rect 2438 1707 2444 1708
rect 2504 1707 2506 1710
rect 1327 1706 1331 1707
rect 111 1702 115 1703
rect 111 1697 115 1698
rect 151 1702 155 1703
rect 151 1697 155 1698
rect 191 1702 195 1703
rect 191 1697 195 1698
rect 255 1702 259 1703
rect 255 1697 259 1698
rect 271 1702 275 1703
rect 271 1697 275 1698
rect 351 1702 355 1703
rect 351 1697 355 1698
rect 367 1702 371 1703
rect 367 1697 371 1698
rect 439 1702 443 1703
rect 439 1697 443 1698
rect 479 1702 483 1703
rect 479 1697 483 1698
rect 535 1702 539 1703
rect 535 1697 539 1698
rect 591 1702 595 1703
rect 591 1697 595 1698
rect 639 1702 643 1703
rect 639 1697 643 1698
rect 695 1702 699 1703
rect 695 1697 699 1698
rect 743 1702 747 1703
rect 743 1697 747 1698
rect 799 1702 803 1703
rect 799 1697 803 1698
rect 847 1702 851 1703
rect 847 1697 851 1698
rect 903 1702 907 1703
rect 903 1697 907 1698
rect 951 1702 955 1703
rect 951 1697 955 1698
rect 1007 1702 1011 1703
rect 1007 1697 1011 1698
rect 1063 1702 1067 1703
rect 1063 1697 1067 1698
rect 1119 1702 1123 1703
rect 1119 1697 1123 1698
rect 1175 1702 1179 1703
rect 1175 1697 1179 1698
rect 1287 1702 1291 1703
rect 1327 1701 1331 1702
rect 1351 1706 1355 1707
rect 1351 1701 1355 1702
rect 1359 1706 1363 1707
rect 1359 1701 1363 1702
rect 1431 1706 1435 1707
rect 1431 1701 1435 1702
rect 1455 1706 1459 1707
rect 1455 1701 1459 1702
rect 1535 1706 1539 1707
rect 1535 1701 1539 1702
rect 1551 1706 1555 1707
rect 1551 1701 1555 1702
rect 1647 1706 1651 1707
rect 1647 1701 1651 1702
rect 1655 1706 1659 1707
rect 1655 1701 1659 1702
rect 1759 1706 1763 1707
rect 1759 1701 1763 1702
rect 1871 1706 1875 1707
rect 1871 1701 1875 1702
rect 1879 1706 1883 1707
rect 1879 1701 1883 1702
rect 1983 1706 1987 1707
rect 1983 1701 1987 1702
rect 2015 1706 2019 1707
rect 2015 1701 2019 1702
rect 2095 1706 2099 1707
rect 2095 1701 2099 1702
rect 2159 1706 2163 1707
rect 2159 1701 2163 1702
rect 2215 1706 2219 1707
rect 2215 1701 2219 1702
rect 2311 1706 2315 1707
rect 2311 1701 2315 1702
rect 2335 1706 2339 1707
rect 2335 1701 2339 1702
rect 2439 1706 2443 1707
rect 2439 1701 2443 1702
rect 2503 1706 2507 1707
rect 2503 1701 2507 1702
rect 1328 1698 1330 1701
rect 1350 1700 1356 1701
rect 1287 1697 1291 1698
rect 1326 1697 1332 1698
rect 112 1677 114 1697
rect 192 1678 194 1697
rect 272 1678 274 1697
rect 352 1678 354 1697
rect 440 1678 442 1697
rect 536 1678 538 1697
rect 640 1678 642 1697
rect 744 1678 746 1697
rect 848 1678 850 1697
rect 952 1678 954 1697
rect 1064 1678 1066 1697
rect 1176 1678 1178 1697
rect 190 1677 196 1678
rect 110 1676 116 1677
rect 110 1672 111 1676
rect 115 1672 116 1676
rect 190 1673 191 1677
rect 195 1673 196 1677
rect 190 1672 196 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 350 1677 356 1678
rect 350 1673 351 1677
rect 355 1673 356 1677
rect 350 1672 356 1673
rect 438 1677 444 1678
rect 438 1673 439 1677
rect 443 1673 444 1677
rect 438 1672 444 1673
rect 534 1677 540 1678
rect 534 1673 535 1677
rect 539 1673 540 1677
rect 534 1672 540 1673
rect 638 1677 644 1678
rect 638 1673 639 1677
rect 643 1673 644 1677
rect 638 1672 644 1673
rect 742 1677 748 1678
rect 742 1673 743 1677
rect 747 1673 748 1677
rect 742 1672 748 1673
rect 846 1677 852 1678
rect 846 1673 847 1677
rect 851 1673 852 1677
rect 846 1672 852 1673
rect 950 1677 956 1678
rect 950 1673 951 1677
rect 955 1673 956 1677
rect 950 1672 956 1673
rect 1062 1677 1068 1678
rect 1062 1673 1063 1677
rect 1067 1673 1068 1677
rect 1062 1672 1068 1673
rect 1174 1677 1180 1678
rect 1288 1677 1290 1697
rect 1326 1693 1327 1697
rect 1331 1693 1332 1697
rect 1350 1696 1351 1700
rect 1355 1696 1356 1700
rect 1350 1695 1356 1696
rect 1430 1700 1436 1701
rect 1430 1696 1431 1700
rect 1435 1696 1436 1700
rect 1430 1695 1436 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1646 1700 1652 1701
rect 1646 1696 1647 1700
rect 1651 1696 1652 1700
rect 1646 1695 1652 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 2014 1700 2020 1701
rect 2014 1696 2015 1700
rect 2019 1696 2020 1700
rect 2014 1695 2020 1696
rect 2158 1700 2164 1701
rect 2158 1696 2159 1700
rect 2163 1696 2164 1700
rect 2158 1695 2164 1696
rect 2310 1700 2316 1701
rect 2310 1696 2311 1700
rect 2315 1696 2316 1700
rect 2310 1695 2316 1696
rect 2438 1700 2444 1701
rect 2438 1696 2439 1700
rect 2443 1696 2444 1700
rect 2504 1698 2506 1701
rect 2438 1695 2444 1696
rect 2502 1697 2508 1698
rect 1326 1692 1332 1693
rect 2502 1693 2503 1697
rect 2507 1693 2508 1697
rect 2502 1692 2508 1693
rect 1326 1680 1332 1681
rect 2502 1680 2508 1681
rect 1174 1673 1175 1677
rect 1179 1673 1180 1677
rect 1174 1672 1180 1673
rect 1286 1676 1292 1677
rect 1286 1672 1287 1676
rect 1291 1672 1292 1676
rect 1326 1676 1327 1680
rect 1331 1676 1332 1680
rect 1326 1675 1332 1676
rect 1366 1679 1372 1680
rect 1366 1675 1367 1679
rect 1371 1675 1372 1679
rect 110 1671 116 1672
rect 1286 1671 1292 1672
rect 110 1659 116 1660
rect 110 1655 111 1659
rect 115 1655 116 1659
rect 1286 1659 1292 1660
rect 110 1654 116 1655
rect 174 1656 180 1657
rect 112 1651 114 1654
rect 174 1652 175 1656
rect 179 1652 180 1656
rect 174 1651 180 1652
rect 254 1656 260 1657
rect 254 1652 255 1656
rect 259 1652 260 1656
rect 254 1651 260 1652
rect 334 1656 340 1657
rect 334 1652 335 1656
rect 339 1652 340 1656
rect 334 1651 340 1652
rect 422 1656 428 1657
rect 422 1652 423 1656
rect 427 1652 428 1656
rect 422 1651 428 1652
rect 518 1656 524 1657
rect 518 1652 519 1656
rect 523 1652 524 1656
rect 518 1651 524 1652
rect 622 1656 628 1657
rect 622 1652 623 1656
rect 627 1652 628 1656
rect 622 1651 628 1652
rect 726 1656 732 1657
rect 726 1652 727 1656
rect 731 1652 732 1656
rect 726 1651 732 1652
rect 830 1656 836 1657
rect 830 1652 831 1656
rect 835 1652 836 1656
rect 830 1651 836 1652
rect 934 1656 940 1657
rect 934 1652 935 1656
rect 939 1652 940 1656
rect 934 1651 940 1652
rect 1046 1656 1052 1657
rect 1046 1652 1047 1656
rect 1051 1652 1052 1656
rect 1046 1651 1052 1652
rect 1158 1656 1164 1657
rect 1158 1652 1159 1656
rect 1163 1652 1164 1656
rect 1286 1655 1287 1659
rect 1291 1655 1292 1659
rect 1286 1654 1292 1655
rect 1158 1651 1164 1652
rect 1288 1651 1290 1654
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 175 1650 179 1651
rect 175 1645 179 1646
rect 215 1650 219 1651
rect 215 1645 219 1646
rect 255 1650 259 1651
rect 255 1645 259 1646
rect 271 1650 275 1651
rect 271 1645 275 1646
rect 335 1650 339 1651
rect 335 1645 339 1646
rect 407 1650 411 1651
rect 407 1645 411 1646
rect 423 1650 427 1651
rect 423 1645 427 1646
rect 479 1650 483 1651
rect 479 1645 483 1646
rect 519 1650 523 1651
rect 519 1645 523 1646
rect 559 1650 563 1651
rect 559 1645 563 1646
rect 623 1650 627 1651
rect 623 1645 627 1646
rect 647 1650 651 1651
rect 647 1645 651 1646
rect 727 1650 731 1651
rect 727 1645 731 1646
rect 743 1650 747 1651
rect 743 1645 747 1646
rect 831 1650 835 1651
rect 831 1645 835 1646
rect 839 1650 843 1651
rect 839 1645 843 1646
rect 935 1650 939 1651
rect 935 1645 939 1646
rect 943 1650 947 1651
rect 943 1645 947 1646
rect 1047 1650 1051 1651
rect 1047 1645 1051 1646
rect 1055 1650 1059 1651
rect 1055 1645 1059 1646
rect 1159 1650 1163 1651
rect 1159 1645 1163 1646
rect 1175 1650 1179 1651
rect 1175 1645 1179 1646
rect 1287 1650 1291 1651
rect 1328 1647 1330 1675
rect 1366 1674 1372 1675
rect 1446 1679 1452 1680
rect 1446 1675 1447 1679
rect 1451 1675 1452 1679
rect 1446 1674 1452 1675
rect 1550 1679 1556 1680
rect 1550 1675 1551 1679
rect 1555 1675 1556 1679
rect 1550 1674 1556 1675
rect 1662 1679 1668 1680
rect 1662 1675 1663 1679
rect 1667 1675 1668 1679
rect 1662 1674 1668 1675
rect 1774 1679 1780 1680
rect 1774 1675 1775 1679
rect 1779 1675 1780 1679
rect 1774 1674 1780 1675
rect 1894 1679 1900 1680
rect 1894 1675 1895 1679
rect 1899 1675 1900 1679
rect 1894 1674 1900 1675
rect 2030 1679 2036 1680
rect 2030 1675 2031 1679
rect 2035 1675 2036 1679
rect 2030 1674 2036 1675
rect 2174 1679 2180 1680
rect 2174 1675 2175 1679
rect 2179 1675 2180 1679
rect 2174 1674 2180 1675
rect 2326 1679 2332 1680
rect 2326 1675 2327 1679
rect 2331 1675 2332 1679
rect 2326 1674 2332 1675
rect 2454 1679 2460 1680
rect 2454 1675 2455 1679
rect 2459 1675 2460 1679
rect 2502 1676 2503 1680
rect 2507 1676 2508 1680
rect 2502 1675 2508 1676
rect 2454 1674 2460 1675
rect 1368 1647 1370 1674
rect 1448 1647 1450 1674
rect 1552 1647 1554 1674
rect 1664 1647 1666 1674
rect 1776 1647 1778 1674
rect 1896 1647 1898 1674
rect 2032 1647 2034 1674
rect 2176 1647 2178 1674
rect 2328 1647 2330 1674
rect 2456 1647 2458 1674
rect 2504 1647 2506 1675
rect 1287 1645 1291 1646
rect 1327 1646 1331 1647
rect 112 1642 114 1645
rect 214 1644 220 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 270 1644 276 1645
rect 270 1640 271 1644
rect 275 1640 276 1644
rect 270 1639 276 1640
rect 334 1644 340 1645
rect 334 1640 335 1644
rect 339 1640 340 1644
rect 334 1639 340 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 478 1644 484 1645
rect 478 1640 479 1644
rect 483 1640 484 1644
rect 478 1639 484 1640
rect 558 1644 564 1645
rect 558 1640 559 1644
rect 563 1640 564 1644
rect 558 1639 564 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 742 1644 748 1645
rect 742 1640 743 1644
rect 747 1640 748 1644
rect 742 1639 748 1640
rect 838 1644 844 1645
rect 838 1640 839 1644
rect 843 1640 844 1644
rect 838 1639 844 1640
rect 942 1644 948 1645
rect 942 1640 943 1644
rect 947 1640 948 1644
rect 942 1639 948 1640
rect 1054 1644 1060 1645
rect 1054 1640 1055 1644
rect 1059 1640 1060 1644
rect 1054 1639 1060 1640
rect 1174 1644 1180 1645
rect 1174 1640 1175 1644
rect 1179 1640 1180 1644
rect 1288 1642 1290 1645
rect 1174 1639 1180 1640
rect 1286 1641 1292 1642
rect 1327 1641 1331 1642
rect 1367 1646 1371 1647
rect 1367 1641 1371 1642
rect 1431 1646 1435 1647
rect 1431 1641 1435 1642
rect 1447 1646 1451 1647
rect 1447 1641 1451 1642
rect 1519 1646 1523 1647
rect 1519 1641 1523 1642
rect 1551 1646 1555 1647
rect 1551 1641 1555 1642
rect 1599 1646 1603 1647
rect 1599 1641 1603 1642
rect 1663 1646 1667 1647
rect 1663 1641 1667 1642
rect 1679 1646 1683 1647
rect 1679 1641 1683 1642
rect 1751 1646 1755 1647
rect 1751 1641 1755 1642
rect 1775 1646 1779 1647
rect 1775 1641 1779 1642
rect 1839 1646 1843 1647
rect 1839 1641 1843 1642
rect 1895 1646 1899 1647
rect 1895 1641 1899 1642
rect 1935 1646 1939 1647
rect 1935 1641 1939 1642
rect 2031 1646 2035 1647
rect 2031 1641 2035 1642
rect 2055 1646 2059 1647
rect 2055 1641 2059 1642
rect 2175 1646 2179 1647
rect 2175 1641 2179 1642
rect 2183 1646 2187 1647
rect 2183 1641 2187 1642
rect 2327 1646 2331 1647
rect 2327 1641 2331 1642
rect 2455 1646 2459 1647
rect 2455 1641 2459 1642
rect 2503 1646 2507 1647
rect 2503 1641 2507 1642
rect 110 1636 116 1637
rect 1286 1637 1287 1641
rect 1291 1637 1292 1641
rect 1286 1636 1292 1637
rect 110 1624 116 1625
rect 1286 1624 1292 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 230 1623 236 1624
rect 230 1619 231 1623
rect 235 1619 236 1623
rect 112 1599 114 1619
rect 230 1618 236 1619
rect 286 1623 292 1624
rect 286 1619 287 1623
rect 291 1619 292 1623
rect 286 1618 292 1619
rect 350 1623 356 1624
rect 350 1619 351 1623
rect 355 1619 356 1623
rect 350 1618 356 1619
rect 422 1623 428 1624
rect 422 1619 423 1623
rect 427 1619 428 1623
rect 422 1618 428 1619
rect 494 1623 500 1624
rect 494 1619 495 1623
rect 499 1619 500 1623
rect 494 1618 500 1619
rect 574 1623 580 1624
rect 574 1619 575 1623
rect 579 1619 580 1623
rect 574 1618 580 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 758 1623 764 1624
rect 758 1619 759 1623
rect 763 1619 764 1623
rect 758 1618 764 1619
rect 854 1623 860 1624
rect 854 1619 855 1623
rect 859 1619 860 1623
rect 854 1618 860 1619
rect 958 1623 964 1624
rect 958 1619 959 1623
rect 963 1619 964 1623
rect 958 1618 964 1619
rect 1070 1623 1076 1624
rect 1070 1619 1071 1623
rect 1075 1619 1076 1623
rect 1070 1618 1076 1619
rect 1190 1623 1196 1624
rect 1190 1619 1191 1623
rect 1195 1619 1196 1623
rect 1286 1620 1287 1624
rect 1291 1620 1292 1624
rect 1328 1621 1330 1641
rect 1368 1622 1370 1641
rect 1432 1622 1434 1641
rect 1520 1622 1522 1641
rect 1600 1622 1602 1641
rect 1680 1622 1682 1641
rect 1752 1622 1754 1641
rect 1840 1622 1842 1641
rect 1936 1622 1938 1641
rect 2056 1622 2058 1641
rect 2184 1622 2186 1641
rect 2328 1622 2330 1641
rect 2456 1622 2458 1641
rect 1366 1621 1372 1622
rect 1286 1619 1292 1620
rect 1326 1620 1332 1621
rect 1190 1618 1196 1619
rect 232 1599 234 1618
rect 288 1599 290 1618
rect 352 1599 354 1618
rect 424 1599 426 1618
rect 496 1599 498 1618
rect 576 1599 578 1618
rect 664 1599 666 1618
rect 760 1599 762 1618
rect 856 1599 858 1618
rect 960 1599 962 1618
rect 1072 1599 1074 1618
rect 1192 1599 1194 1618
rect 1288 1599 1290 1619
rect 1326 1616 1327 1620
rect 1331 1616 1332 1620
rect 1366 1617 1367 1621
rect 1371 1617 1372 1621
rect 1366 1616 1372 1617
rect 1430 1621 1436 1622
rect 1430 1617 1431 1621
rect 1435 1617 1436 1621
rect 1430 1616 1436 1617
rect 1518 1621 1524 1622
rect 1518 1617 1519 1621
rect 1523 1617 1524 1621
rect 1518 1616 1524 1617
rect 1598 1621 1604 1622
rect 1598 1617 1599 1621
rect 1603 1617 1604 1621
rect 1598 1616 1604 1617
rect 1678 1621 1684 1622
rect 1678 1617 1679 1621
rect 1683 1617 1684 1621
rect 1678 1616 1684 1617
rect 1750 1621 1756 1622
rect 1750 1617 1751 1621
rect 1755 1617 1756 1621
rect 1750 1616 1756 1617
rect 1838 1621 1844 1622
rect 1838 1617 1839 1621
rect 1843 1617 1844 1621
rect 1838 1616 1844 1617
rect 1934 1621 1940 1622
rect 1934 1617 1935 1621
rect 1939 1617 1940 1621
rect 1934 1616 1940 1617
rect 2054 1621 2060 1622
rect 2054 1617 2055 1621
rect 2059 1617 2060 1621
rect 2054 1616 2060 1617
rect 2182 1621 2188 1622
rect 2182 1617 2183 1621
rect 2187 1617 2188 1621
rect 2182 1616 2188 1617
rect 2326 1621 2332 1622
rect 2326 1617 2327 1621
rect 2331 1617 2332 1621
rect 2326 1616 2332 1617
rect 2454 1621 2460 1622
rect 2504 1621 2506 1641
rect 2454 1617 2455 1621
rect 2459 1617 2460 1621
rect 2454 1616 2460 1617
rect 2502 1620 2508 1621
rect 2502 1616 2503 1620
rect 2507 1616 2508 1620
rect 1326 1615 1332 1616
rect 2502 1615 2508 1616
rect 1326 1603 1332 1604
rect 1326 1599 1327 1603
rect 1331 1599 1332 1603
rect 2502 1603 2508 1604
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 231 1598 235 1599
rect 231 1593 235 1594
rect 287 1598 291 1599
rect 287 1593 291 1594
rect 351 1598 355 1599
rect 351 1593 355 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 495 1598 499 1599
rect 495 1593 499 1594
rect 503 1598 507 1599
rect 503 1593 507 1594
rect 575 1598 579 1599
rect 575 1593 579 1594
rect 599 1598 603 1599
rect 599 1593 603 1594
rect 663 1598 667 1599
rect 663 1593 667 1594
rect 703 1598 707 1599
rect 703 1593 707 1594
rect 759 1598 763 1599
rect 759 1593 763 1594
rect 815 1598 819 1599
rect 815 1593 819 1594
rect 855 1598 859 1599
rect 855 1593 859 1594
rect 935 1598 939 1599
rect 935 1593 939 1594
rect 959 1598 963 1599
rect 959 1593 963 1594
rect 1063 1598 1067 1599
rect 1063 1593 1067 1594
rect 1071 1598 1075 1599
rect 1071 1593 1075 1594
rect 1191 1598 1195 1599
rect 1191 1593 1195 1594
rect 1287 1598 1291 1599
rect 1326 1598 1332 1599
rect 1350 1600 1356 1601
rect 1287 1593 1291 1594
rect 112 1573 114 1593
rect 288 1574 290 1593
rect 352 1574 354 1593
rect 424 1574 426 1593
rect 504 1574 506 1593
rect 600 1574 602 1593
rect 704 1574 706 1593
rect 816 1574 818 1593
rect 936 1574 938 1593
rect 1064 1574 1066 1593
rect 1192 1574 1194 1593
rect 286 1573 292 1574
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 286 1569 287 1573
rect 291 1569 292 1573
rect 286 1568 292 1569
rect 350 1573 356 1574
rect 350 1569 351 1573
rect 355 1569 356 1573
rect 350 1568 356 1569
rect 422 1573 428 1574
rect 422 1569 423 1573
rect 427 1569 428 1573
rect 422 1568 428 1569
rect 502 1573 508 1574
rect 502 1569 503 1573
rect 507 1569 508 1573
rect 502 1568 508 1569
rect 598 1573 604 1574
rect 598 1569 599 1573
rect 603 1569 604 1573
rect 598 1568 604 1569
rect 702 1573 708 1574
rect 702 1569 703 1573
rect 707 1569 708 1573
rect 702 1568 708 1569
rect 814 1573 820 1574
rect 814 1569 815 1573
rect 819 1569 820 1573
rect 814 1568 820 1569
rect 934 1573 940 1574
rect 934 1569 935 1573
rect 939 1569 940 1573
rect 934 1568 940 1569
rect 1062 1573 1068 1574
rect 1062 1569 1063 1573
rect 1067 1569 1068 1573
rect 1062 1568 1068 1569
rect 1190 1573 1196 1574
rect 1288 1573 1290 1593
rect 1328 1591 1330 1598
rect 1350 1596 1351 1600
rect 1355 1596 1356 1600
rect 1350 1595 1356 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1502 1600 1508 1601
rect 1502 1596 1503 1600
rect 1507 1596 1508 1600
rect 1502 1595 1508 1596
rect 1582 1600 1588 1601
rect 1582 1596 1583 1600
rect 1587 1596 1588 1600
rect 1582 1595 1588 1596
rect 1662 1600 1668 1601
rect 1662 1596 1663 1600
rect 1667 1596 1668 1600
rect 1662 1595 1668 1596
rect 1734 1600 1740 1601
rect 1734 1596 1735 1600
rect 1739 1596 1740 1600
rect 1734 1595 1740 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1918 1600 1924 1601
rect 1918 1596 1919 1600
rect 1923 1596 1924 1600
rect 1918 1595 1924 1596
rect 2038 1600 2044 1601
rect 2038 1596 2039 1600
rect 2043 1596 2044 1600
rect 2038 1595 2044 1596
rect 2166 1600 2172 1601
rect 2166 1596 2167 1600
rect 2171 1596 2172 1600
rect 2166 1595 2172 1596
rect 2310 1600 2316 1601
rect 2310 1596 2311 1600
rect 2315 1596 2316 1600
rect 2310 1595 2316 1596
rect 2438 1600 2444 1601
rect 2438 1596 2439 1600
rect 2443 1596 2444 1600
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2438 1595 2444 1596
rect 1352 1591 1354 1595
rect 1416 1591 1418 1595
rect 1504 1591 1506 1595
rect 1584 1591 1586 1595
rect 1664 1591 1666 1595
rect 1736 1591 1738 1595
rect 1824 1591 1826 1595
rect 1920 1591 1922 1595
rect 2040 1591 2042 1595
rect 2168 1591 2170 1595
rect 2312 1591 2314 1595
rect 2440 1591 2442 1595
rect 2504 1591 2506 1598
rect 1327 1590 1331 1591
rect 1327 1585 1331 1586
rect 1351 1590 1355 1591
rect 1351 1585 1355 1586
rect 1415 1590 1419 1591
rect 1415 1585 1419 1586
rect 1423 1590 1427 1591
rect 1423 1585 1427 1586
rect 1503 1590 1507 1591
rect 1503 1585 1507 1586
rect 1527 1590 1531 1591
rect 1527 1585 1531 1586
rect 1583 1590 1587 1591
rect 1583 1585 1587 1586
rect 1647 1590 1651 1591
rect 1647 1585 1651 1586
rect 1663 1590 1667 1591
rect 1663 1585 1667 1586
rect 1735 1590 1739 1591
rect 1735 1585 1739 1586
rect 1783 1590 1787 1591
rect 1783 1585 1787 1586
rect 1823 1590 1827 1591
rect 1823 1585 1827 1586
rect 1919 1590 1923 1591
rect 1919 1585 1923 1586
rect 1935 1590 1939 1591
rect 1935 1585 1939 1586
rect 2039 1590 2043 1591
rect 2039 1585 2043 1586
rect 2103 1590 2107 1591
rect 2103 1585 2107 1586
rect 2167 1590 2171 1591
rect 2167 1585 2171 1586
rect 2279 1590 2283 1591
rect 2279 1585 2283 1586
rect 2311 1590 2315 1591
rect 2311 1585 2315 1586
rect 2439 1590 2443 1591
rect 2439 1585 2443 1586
rect 2503 1590 2507 1591
rect 2503 1585 2507 1586
rect 1328 1582 1330 1585
rect 1350 1584 1356 1585
rect 1326 1581 1332 1582
rect 1326 1577 1327 1581
rect 1331 1577 1332 1581
rect 1350 1580 1351 1584
rect 1355 1580 1356 1584
rect 1350 1579 1356 1580
rect 1422 1584 1428 1585
rect 1422 1580 1423 1584
rect 1427 1580 1428 1584
rect 1422 1579 1428 1580
rect 1526 1584 1532 1585
rect 1526 1580 1527 1584
rect 1531 1580 1532 1584
rect 1526 1579 1532 1580
rect 1646 1584 1652 1585
rect 1646 1580 1647 1584
rect 1651 1580 1652 1584
rect 1646 1579 1652 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1934 1584 1940 1585
rect 1934 1580 1935 1584
rect 1939 1580 1940 1584
rect 1934 1579 1940 1580
rect 2102 1584 2108 1585
rect 2102 1580 2103 1584
rect 2107 1580 2108 1584
rect 2102 1579 2108 1580
rect 2278 1584 2284 1585
rect 2278 1580 2279 1584
rect 2283 1580 2284 1584
rect 2278 1579 2284 1580
rect 2438 1584 2444 1585
rect 2438 1580 2439 1584
rect 2443 1580 2444 1584
rect 2504 1582 2506 1585
rect 2438 1579 2444 1580
rect 2502 1581 2508 1582
rect 1326 1576 1332 1577
rect 2502 1577 2503 1581
rect 2507 1577 2508 1581
rect 2502 1576 2508 1577
rect 1190 1569 1191 1573
rect 1195 1569 1196 1573
rect 1190 1568 1196 1569
rect 1286 1572 1292 1573
rect 1286 1568 1287 1572
rect 1291 1568 1292 1572
rect 110 1567 116 1568
rect 1286 1567 1292 1568
rect 1326 1564 1332 1565
rect 2502 1564 2508 1565
rect 1326 1560 1327 1564
rect 1331 1560 1332 1564
rect 1326 1559 1332 1560
rect 1366 1563 1372 1564
rect 1366 1559 1367 1563
rect 1371 1559 1372 1563
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1286 1555 1292 1556
rect 110 1550 116 1551
rect 270 1552 276 1553
rect 112 1539 114 1550
rect 270 1548 271 1552
rect 275 1548 276 1552
rect 270 1547 276 1548
rect 334 1552 340 1553
rect 334 1548 335 1552
rect 339 1548 340 1552
rect 334 1547 340 1548
rect 406 1552 412 1553
rect 406 1548 407 1552
rect 411 1548 412 1552
rect 406 1547 412 1548
rect 486 1552 492 1553
rect 486 1548 487 1552
rect 491 1548 492 1552
rect 486 1547 492 1548
rect 582 1552 588 1553
rect 582 1548 583 1552
rect 587 1548 588 1552
rect 582 1547 588 1548
rect 686 1552 692 1553
rect 686 1548 687 1552
rect 691 1548 692 1552
rect 686 1547 692 1548
rect 798 1552 804 1553
rect 798 1548 799 1552
rect 803 1548 804 1552
rect 798 1547 804 1548
rect 918 1552 924 1553
rect 918 1548 919 1552
rect 923 1548 924 1552
rect 918 1547 924 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1174 1552 1180 1553
rect 1174 1548 1175 1552
rect 1179 1548 1180 1552
rect 1286 1551 1287 1555
rect 1291 1551 1292 1555
rect 1286 1550 1292 1551
rect 1174 1547 1180 1548
rect 272 1539 274 1547
rect 336 1539 338 1547
rect 408 1539 410 1547
rect 488 1539 490 1547
rect 584 1539 586 1547
rect 688 1539 690 1547
rect 800 1539 802 1547
rect 920 1539 922 1547
rect 1048 1539 1050 1547
rect 1176 1539 1178 1547
rect 1288 1539 1290 1550
rect 1328 1539 1330 1559
rect 1366 1558 1372 1559
rect 1438 1563 1444 1564
rect 1438 1559 1439 1563
rect 1443 1559 1444 1563
rect 1438 1558 1444 1559
rect 1542 1563 1548 1564
rect 1542 1559 1543 1563
rect 1547 1559 1548 1563
rect 1542 1558 1548 1559
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1559 1668 1563
rect 1662 1558 1668 1559
rect 1798 1563 1804 1564
rect 1798 1559 1799 1563
rect 1803 1559 1804 1563
rect 1798 1558 1804 1559
rect 1950 1563 1956 1564
rect 1950 1559 1951 1563
rect 1955 1559 1956 1563
rect 1950 1558 1956 1559
rect 2118 1563 2124 1564
rect 2118 1559 2119 1563
rect 2123 1559 2124 1563
rect 2118 1558 2124 1559
rect 2294 1563 2300 1564
rect 2294 1559 2295 1563
rect 2299 1559 2300 1563
rect 2294 1558 2300 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2502 1560 2503 1564
rect 2507 1560 2508 1564
rect 2502 1559 2508 1560
rect 2454 1558 2460 1559
rect 1368 1539 1370 1558
rect 1440 1539 1442 1558
rect 1544 1539 1546 1558
rect 1664 1539 1666 1558
rect 1800 1539 1802 1558
rect 1952 1539 1954 1558
rect 2120 1539 2122 1558
rect 2296 1539 2298 1558
rect 2456 1539 2458 1558
rect 2504 1539 2506 1559
rect 111 1538 115 1539
rect 111 1533 115 1534
rect 271 1538 275 1539
rect 271 1533 275 1534
rect 335 1538 339 1539
rect 335 1533 339 1534
rect 407 1538 411 1539
rect 407 1533 411 1534
rect 471 1538 475 1539
rect 471 1533 475 1534
rect 487 1538 491 1539
rect 487 1533 491 1534
rect 551 1538 555 1539
rect 551 1533 555 1534
rect 583 1538 587 1539
rect 583 1533 587 1534
rect 639 1538 643 1539
rect 639 1533 643 1534
rect 687 1538 691 1539
rect 687 1533 691 1534
rect 735 1538 739 1539
rect 735 1533 739 1534
rect 799 1538 803 1539
rect 799 1533 803 1534
rect 839 1538 843 1539
rect 839 1533 843 1534
rect 919 1538 923 1539
rect 919 1533 923 1534
rect 951 1538 955 1539
rect 951 1533 955 1534
rect 1047 1538 1051 1539
rect 1047 1533 1051 1534
rect 1063 1538 1067 1539
rect 1063 1533 1067 1534
rect 1175 1538 1179 1539
rect 1175 1533 1179 1534
rect 1287 1538 1291 1539
rect 1287 1533 1291 1534
rect 1327 1538 1331 1539
rect 1327 1533 1331 1534
rect 1367 1538 1371 1539
rect 1367 1533 1371 1534
rect 1439 1538 1443 1539
rect 1439 1533 1443 1534
rect 1543 1538 1547 1539
rect 1543 1533 1547 1534
rect 1647 1538 1651 1539
rect 1647 1533 1651 1534
rect 1663 1538 1667 1539
rect 1663 1533 1667 1534
rect 1751 1538 1755 1539
rect 1751 1533 1755 1534
rect 1799 1538 1803 1539
rect 1799 1533 1803 1534
rect 1855 1538 1859 1539
rect 1855 1533 1859 1534
rect 1951 1538 1955 1539
rect 1951 1533 1955 1534
rect 1959 1538 1963 1539
rect 1959 1533 1963 1534
rect 2055 1538 2059 1539
rect 2055 1533 2059 1534
rect 2119 1538 2123 1539
rect 2119 1533 2123 1534
rect 2151 1538 2155 1539
rect 2151 1533 2155 1534
rect 2247 1538 2251 1539
rect 2247 1533 2251 1534
rect 2295 1538 2299 1539
rect 2295 1533 2299 1534
rect 2343 1538 2347 1539
rect 2343 1533 2347 1534
rect 2439 1538 2443 1539
rect 2439 1533 2443 1534
rect 2455 1538 2459 1539
rect 2455 1533 2459 1534
rect 2503 1538 2507 1539
rect 2503 1533 2507 1534
rect 112 1530 114 1533
rect 470 1532 476 1533
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 470 1528 471 1532
rect 475 1528 476 1532
rect 470 1527 476 1528
rect 550 1532 556 1533
rect 550 1528 551 1532
rect 555 1528 556 1532
rect 550 1527 556 1528
rect 638 1532 644 1533
rect 638 1528 639 1532
rect 643 1528 644 1532
rect 638 1527 644 1528
rect 734 1532 740 1533
rect 734 1528 735 1532
rect 739 1528 740 1532
rect 734 1527 740 1528
rect 838 1532 844 1533
rect 838 1528 839 1532
rect 843 1528 844 1532
rect 838 1527 844 1528
rect 950 1532 956 1533
rect 950 1528 951 1532
rect 955 1528 956 1532
rect 950 1527 956 1528
rect 1062 1532 1068 1533
rect 1062 1528 1063 1532
rect 1067 1528 1068 1532
rect 1062 1527 1068 1528
rect 1174 1532 1180 1533
rect 1174 1528 1175 1532
rect 1179 1528 1180 1532
rect 1288 1530 1290 1533
rect 1174 1527 1180 1528
rect 1286 1529 1292 1530
rect 110 1524 116 1525
rect 1286 1525 1287 1529
rect 1291 1525 1292 1529
rect 1286 1524 1292 1525
rect 1328 1513 1330 1533
rect 1368 1514 1370 1533
rect 1440 1514 1442 1533
rect 1544 1514 1546 1533
rect 1648 1514 1650 1533
rect 1752 1514 1754 1533
rect 1856 1514 1858 1533
rect 1960 1514 1962 1533
rect 2056 1514 2058 1533
rect 2152 1514 2154 1533
rect 2248 1514 2250 1533
rect 2344 1514 2346 1533
rect 2440 1514 2442 1533
rect 1366 1513 1372 1514
rect 110 1512 116 1513
rect 1286 1512 1292 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 486 1511 492 1512
rect 486 1507 487 1511
rect 491 1507 492 1511
rect 112 1487 114 1507
rect 486 1506 492 1507
rect 566 1511 572 1512
rect 566 1507 567 1511
rect 571 1507 572 1511
rect 566 1506 572 1507
rect 654 1511 660 1512
rect 654 1507 655 1511
rect 659 1507 660 1511
rect 654 1506 660 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 854 1511 860 1512
rect 854 1507 855 1511
rect 859 1507 860 1511
rect 854 1506 860 1507
rect 966 1511 972 1512
rect 966 1507 967 1511
rect 971 1507 972 1511
rect 966 1506 972 1507
rect 1078 1511 1084 1512
rect 1078 1507 1079 1511
rect 1083 1507 1084 1511
rect 1078 1506 1084 1507
rect 1190 1511 1196 1512
rect 1190 1507 1191 1511
rect 1195 1507 1196 1511
rect 1286 1508 1287 1512
rect 1291 1508 1292 1512
rect 1286 1507 1292 1508
rect 1326 1512 1332 1513
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1366 1509 1367 1513
rect 1371 1509 1372 1513
rect 1366 1508 1372 1509
rect 1438 1513 1444 1514
rect 1438 1509 1439 1513
rect 1443 1509 1444 1513
rect 1438 1508 1444 1509
rect 1542 1513 1548 1514
rect 1542 1509 1543 1513
rect 1547 1509 1548 1513
rect 1542 1508 1548 1509
rect 1646 1513 1652 1514
rect 1646 1509 1647 1513
rect 1651 1509 1652 1513
rect 1646 1508 1652 1509
rect 1750 1513 1756 1514
rect 1750 1509 1751 1513
rect 1755 1509 1756 1513
rect 1750 1508 1756 1509
rect 1854 1513 1860 1514
rect 1854 1509 1855 1513
rect 1859 1509 1860 1513
rect 1854 1508 1860 1509
rect 1958 1513 1964 1514
rect 1958 1509 1959 1513
rect 1963 1509 1964 1513
rect 1958 1508 1964 1509
rect 2054 1513 2060 1514
rect 2054 1509 2055 1513
rect 2059 1509 2060 1513
rect 2054 1508 2060 1509
rect 2150 1513 2156 1514
rect 2150 1509 2151 1513
rect 2155 1509 2156 1513
rect 2150 1508 2156 1509
rect 2246 1513 2252 1514
rect 2246 1509 2247 1513
rect 2251 1509 2252 1513
rect 2246 1508 2252 1509
rect 2342 1513 2348 1514
rect 2342 1509 2343 1513
rect 2347 1509 2348 1513
rect 2342 1508 2348 1509
rect 2438 1513 2444 1514
rect 2504 1513 2506 1533
rect 2438 1509 2439 1513
rect 2443 1509 2444 1513
rect 2438 1508 2444 1509
rect 2502 1512 2508 1513
rect 2502 1508 2503 1512
rect 2507 1508 2508 1512
rect 1326 1507 1332 1508
rect 2502 1507 2508 1508
rect 1190 1506 1196 1507
rect 488 1487 490 1506
rect 568 1487 570 1506
rect 656 1487 658 1506
rect 752 1487 754 1506
rect 856 1487 858 1506
rect 968 1487 970 1506
rect 1080 1487 1082 1506
rect 1192 1487 1194 1506
rect 1288 1487 1290 1507
rect 1326 1495 1332 1496
rect 1326 1491 1327 1495
rect 1331 1491 1332 1495
rect 2502 1495 2508 1496
rect 1326 1490 1332 1491
rect 1350 1492 1356 1493
rect 111 1486 115 1487
rect 111 1481 115 1482
rect 375 1486 379 1487
rect 375 1481 379 1482
rect 463 1486 467 1487
rect 463 1481 467 1482
rect 487 1486 491 1487
rect 487 1481 491 1482
rect 559 1486 563 1487
rect 559 1481 563 1482
rect 567 1486 571 1487
rect 567 1481 571 1482
rect 655 1486 659 1487
rect 655 1481 659 1482
rect 751 1486 755 1487
rect 751 1481 755 1482
rect 855 1486 859 1487
rect 855 1481 859 1482
rect 959 1486 963 1487
rect 959 1481 963 1482
rect 967 1486 971 1487
rect 967 1481 971 1482
rect 1063 1486 1067 1487
rect 1063 1481 1067 1482
rect 1079 1486 1083 1487
rect 1079 1481 1083 1482
rect 1167 1486 1171 1487
rect 1167 1481 1171 1482
rect 1191 1486 1195 1487
rect 1191 1481 1195 1482
rect 1287 1486 1291 1487
rect 1328 1483 1330 1490
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1422 1492 1428 1493
rect 1422 1488 1423 1492
rect 1427 1488 1428 1492
rect 1422 1487 1428 1488
rect 1526 1492 1532 1493
rect 1526 1488 1527 1492
rect 1531 1488 1532 1492
rect 1526 1487 1532 1488
rect 1630 1492 1636 1493
rect 1630 1488 1631 1492
rect 1635 1488 1636 1492
rect 1630 1487 1636 1488
rect 1734 1492 1740 1493
rect 1734 1488 1735 1492
rect 1739 1488 1740 1492
rect 1734 1487 1740 1488
rect 1838 1492 1844 1493
rect 1838 1488 1839 1492
rect 1843 1488 1844 1492
rect 1838 1487 1844 1488
rect 1942 1492 1948 1493
rect 1942 1488 1943 1492
rect 1947 1488 1948 1492
rect 1942 1487 1948 1488
rect 2038 1492 2044 1493
rect 2038 1488 2039 1492
rect 2043 1488 2044 1492
rect 2038 1487 2044 1488
rect 2134 1492 2140 1493
rect 2134 1488 2135 1492
rect 2139 1488 2140 1492
rect 2134 1487 2140 1488
rect 2230 1492 2236 1493
rect 2230 1488 2231 1492
rect 2235 1488 2236 1492
rect 2230 1487 2236 1488
rect 2326 1492 2332 1493
rect 2326 1488 2327 1492
rect 2331 1488 2332 1492
rect 2326 1487 2332 1488
rect 2422 1492 2428 1493
rect 2422 1488 2423 1492
rect 2427 1488 2428 1492
rect 2502 1491 2503 1495
rect 2507 1491 2508 1495
rect 2502 1490 2508 1491
rect 2422 1487 2428 1488
rect 1352 1483 1354 1487
rect 1424 1483 1426 1487
rect 1528 1483 1530 1487
rect 1632 1483 1634 1487
rect 1736 1483 1738 1487
rect 1840 1483 1842 1487
rect 1944 1483 1946 1487
rect 2040 1483 2042 1487
rect 2136 1483 2138 1487
rect 2232 1483 2234 1487
rect 2328 1483 2330 1487
rect 2424 1483 2426 1487
rect 2504 1483 2506 1490
rect 1287 1481 1291 1482
rect 1327 1482 1331 1483
rect 112 1461 114 1481
rect 376 1462 378 1481
rect 464 1462 466 1481
rect 560 1462 562 1481
rect 656 1462 658 1481
rect 752 1462 754 1481
rect 856 1462 858 1481
rect 960 1462 962 1481
rect 1064 1462 1066 1481
rect 1168 1462 1170 1481
rect 374 1461 380 1462
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 374 1457 375 1461
rect 379 1457 380 1461
rect 374 1456 380 1457
rect 462 1461 468 1462
rect 462 1457 463 1461
rect 467 1457 468 1461
rect 462 1456 468 1457
rect 558 1461 564 1462
rect 558 1457 559 1461
rect 563 1457 564 1461
rect 558 1456 564 1457
rect 654 1461 660 1462
rect 654 1457 655 1461
rect 659 1457 660 1461
rect 654 1456 660 1457
rect 750 1461 756 1462
rect 750 1457 751 1461
rect 755 1457 756 1461
rect 750 1456 756 1457
rect 854 1461 860 1462
rect 854 1457 855 1461
rect 859 1457 860 1461
rect 854 1456 860 1457
rect 958 1461 964 1462
rect 958 1457 959 1461
rect 963 1457 964 1461
rect 958 1456 964 1457
rect 1062 1461 1068 1462
rect 1062 1457 1063 1461
rect 1067 1457 1068 1461
rect 1062 1456 1068 1457
rect 1166 1461 1172 1462
rect 1288 1461 1290 1481
rect 1327 1477 1331 1478
rect 1351 1482 1355 1483
rect 1351 1477 1355 1478
rect 1423 1482 1427 1483
rect 1423 1477 1427 1478
rect 1519 1482 1523 1483
rect 1519 1477 1523 1478
rect 1527 1482 1531 1483
rect 1527 1477 1531 1478
rect 1615 1482 1619 1483
rect 1615 1477 1619 1478
rect 1631 1482 1635 1483
rect 1631 1477 1635 1478
rect 1711 1482 1715 1483
rect 1711 1477 1715 1478
rect 1735 1482 1739 1483
rect 1735 1477 1739 1478
rect 1815 1482 1819 1483
rect 1815 1477 1819 1478
rect 1839 1482 1843 1483
rect 1839 1477 1843 1478
rect 1927 1482 1931 1483
rect 1927 1477 1931 1478
rect 1943 1482 1947 1483
rect 1943 1477 1947 1478
rect 2039 1482 2043 1483
rect 2039 1477 2043 1478
rect 2047 1482 2051 1483
rect 2047 1477 2051 1478
rect 2135 1482 2139 1483
rect 2135 1477 2139 1478
rect 2175 1482 2179 1483
rect 2175 1477 2179 1478
rect 2231 1482 2235 1483
rect 2231 1477 2235 1478
rect 2303 1482 2307 1483
rect 2303 1477 2307 1478
rect 2327 1482 2331 1483
rect 2327 1477 2331 1478
rect 2423 1482 2427 1483
rect 2423 1477 2427 1478
rect 2439 1482 2443 1483
rect 2439 1477 2443 1478
rect 2503 1482 2507 1483
rect 2503 1477 2507 1478
rect 1328 1474 1330 1477
rect 1350 1476 1356 1477
rect 1326 1473 1332 1474
rect 1326 1469 1327 1473
rect 1331 1469 1332 1473
rect 1350 1472 1351 1476
rect 1355 1472 1356 1476
rect 1350 1471 1356 1472
rect 1422 1476 1428 1477
rect 1422 1472 1423 1476
rect 1427 1472 1428 1476
rect 1422 1471 1428 1472
rect 1518 1476 1524 1477
rect 1518 1472 1519 1476
rect 1523 1472 1524 1476
rect 1518 1471 1524 1472
rect 1614 1476 1620 1477
rect 1614 1472 1615 1476
rect 1619 1472 1620 1476
rect 1614 1471 1620 1472
rect 1710 1476 1716 1477
rect 1710 1472 1711 1476
rect 1715 1472 1716 1476
rect 1710 1471 1716 1472
rect 1814 1476 1820 1477
rect 1814 1472 1815 1476
rect 1819 1472 1820 1476
rect 1814 1471 1820 1472
rect 1926 1476 1932 1477
rect 1926 1472 1927 1476
rect 1931 1472 1932 1476
rect 1926 1471 1932 1472
rect 2046 1476 2052 1477
rect 2046 1472 2047 1476
rect 2051 1472 2052 1476
rect 2046 1471 2052 1472
rect 2174 1476 2180 1477
rect 2174 1472 2175 1476
rect 2179 1472 2180 1476
rect 2174 1471 2180 1472
rect 2302 1476 2308 1477
rect 2302 1472 2303 1476
rect 2307 1472 2308 1476
rect 2302 1471 2308 1472
rect 2438 1476 2444 1477
rect 2438 1472 2439 1476
rect 2443 1472 2444 1476
rect 2504 1474 2506 1477
rect 2438 1471 2444 1472
rect 2502 1473 2508 1474
rect 1326 1468 1332 1469
rect 2502 1469 2503 1473
rect 2507 1469 2508 1473
rect 2502 1468 2508 1469
rect 1166 1457 1167 1461
rect 1171 1457 1172 1461
rect 1166 1456 1172 1457
rect 1286 1460 1292 1461
rect 1286 1456 1287 1460
rect 1291 1456 1292 1460
rect 110 1455 116 1456
rect 1286 1455 1292 1456
rect 1326 1456 1332 1457
rect 2502 1456 2508 1457
rect 1326 1452 1327 1456
rect 1331 1452 1332 1456
rect 1326 1451 1332 1452
rect 1366 1455 1372 1456
rect 1366 1451 1367 1455
rect 1371 1451 1372 1455
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 1286 1443 1292 1444
rect 110 1438 116 1439
rect 358 1440 364 1441
rect 112 1435 114 1438
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 446 1440 452 1441
rect 446 1436 447 1440
rect 451 1436 452 1440
rect 446 1435 452 1436
rect 542 1440 548 1441
rect 542 1436 543 1440
rect 547 1436 548 1440
rect 542 1435 548 1436
rect 638 1440 644 1441
rect 638 1436 639 1440
rect 643 1436 644 1440
rect 638 1435 644 1436
rect 734 1440 740 1441
rect 734 1436 735 1440
rect 739 1436 740 1440
rect 734 1435 740 1436
rect 838 1440 844 1441
rect 838 1436 839 1440
rect 843 1436 844 1440
rect 838 1435 844 1436
rect 942 1440 948 1441
rect 942 1436 943 1440
rect 947 1436 948 1440
rect 942 1435 948 1436
rect 1046 1440 1052 1441
rect 1046 1436 1047 1440
rect 1051 1436 1052 1440
rect 1046 1435 1052 1436
rect 1150 1440 1156 1441
rect 1150 1436 1151 1440
rect 1155 1436 1156 1440
rect 1286 1439 1287 1443
rect 1291 1439 1292 1443
rect 1286 1438 1292 1439
rect 1150 1435 1156 1436
rect 1288 1435 1290 1438
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 231 1434 235 1435
rect 231 1429 235 1430
rect 319 1434 323 1435
rect 319 1429 323 1430
rect 359 1434 363 1435
rect 359 1429 363 1430
rect 415 1434 419 1435
rect 415 1429 419 1430
rect 447 1434 451 1435
rect 447 1429 451 1430
rect 511 1434 515 1435
rect 511 1429 515 1430
rect 543 1434 547 1435
rect 543 1429 547 1430
rect 615 1434 619 1435
rect 615 1429 619 1430
rect 639 1434 643 1435
rect 639 1429 643 1430
rect 711 1434 715 1435
rect 711 1429 715 1430
rect 735 1434 739 1435
rect 735 1429 739 1430
rect 807 1434 811 1435
rect 807 1429 811 1430
rect 839 1434 843 1435
rect 839 1429 843 1430
rect 895 1434 899 1435
rect 895 1429 899 1430
rect 943 1434 947 1435
rect 943 1429 947 1430
rect 991 1434 995 1435
rect 991 1429 995 1430
rect 1047 1434 1051 1435
rect 1047 1429 1051 1430
rect 1087 1434 1091 1435
rect 1087 1429 1091 1430
rect 1151 1434 1155 1435
rect 1151 1429 1155 1430
rect 1287 1434 1291 1435
rect 1287 1429 1291 1430
rect 112 1426 114 1429
rect 230 1428 236 1429
rect 110 1425 116 1426
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 230 1424 231 1428
rect 235 1424 236 1428
rect 230 1423 236 1424
rect 318 1428 324 1429
rect 318 1424 319 1428
rect 323 1424 324 1428
rect 318 1423 324 1424
rect 414 1428 420 1429
rect 414 1424 415 1428
rect 419 1424 420 1428
rect 414 1423 420 1424
rect 510 1428 516 1429
rect 510 1424 511 1428
rect 515 1424 516 1428
rect 510 1423 516 1424
rect 614 1428 620 1429
rect 614 1424 615 1428
rect 619 1424 620 1428
rect 614 1423 620 1424
rect 710 1428 716 1429
rect 710 1424 711 1428
rect 715 1424 716 1428
rect 710 1423 716 1424
rect 806 1428 812 1429
rect 806 1424 807 1428
rect 811 1424 812 1428
rect 806 1423 812 1424
rect 894 1428 900 1429
rect 894 1424 895 1428
rect 899 1424 900 1428
rect 894 1423 900 1424
rect 990 1428 996 1429
rect 990 1424 991 1428
rect 995 1424 996 1428
rect 990 1423 996 1424
rect 1086 1428 1092 1429
rect 1086 1424 1087 1428
rect 1091 1424 1092 1428
rect 1288 1426 1290 1429
rect 1328 1427 1330 1451
rect 1366 1450 1372 1451
rect 1438 1455 1444 1456
rect 1438 1451 1439 1455
rect 1443 1451 1444 1455
rect 1438 1450 1444 1451
rect 1534 1455 1540 1456
rect 1534 1451 1535 1455
rect 1539 1451 1540 1455
rect 1534 1450 1540 1451
rect 1630 1455 1636 1456
rect 1630 1451 1631 1455
rect 1635 1451 1636 1455
rect 1630 1450 1636 1451
rect 1726 1455 1732 1456
rect 1726 1451 1727 1455
rect 1731 1451 1732 1455
rect 1726 1450 1732 1451
rect 1830 1455 1836 1456
rect 1830 1451 1831 1455
rect 1835 1451 1836 1455
rect 1830 1450 1836 1451
rect 1942 1455 1948 1456
rect 1942 1451 1943 1455
rect 1947 1451 1948 1455
rect 1942 1450 1948 1451
rect 2062 1455 2068 1456
rect 2062 1451 2063 1455
rect 2067 1451 2068 1455
rect 2062 1450 2068 1451
rect 2190 1455 2196 1456
rect 2190 1451 2191 1455
rect 2195 1451 2196 1455
rect 2190 1450 2196 1451
rect 2318 1455 2324 1456
rect 2318 1451 2319 1455
rect 2323 1451 2324 1455
rect 2318 1450 2324 1451
rect 2454 1455 2460 1456
rect 2454 1451 2455 1455
rect 2459 1451 2460 1455
rect 2502 1452 2503 1456
rect 2507 1452 2508 1456
rect 2502 1451 2508 1452
rect 2454 1450 2460 1451
rect 1368 1427 1370 1450
rect 1440 1427 1442 1450
rect 1536 1427 1538 1450
rect 1632 1427 1634 1450
rect 1728 1427 1730 1450
rect 1832 1427 1834 1450
rect 1944 1427 1946 1450
rect 2064 1427 2066 1450
rect 2192 1427 2194 1450
rect 2320 1427 2322 1450
rect 2456 1427 2458 1450
rect 2504 1427 2506 1451
rect 1327 1426 1331 1427
rect 1086 1423 1092 1424
rect 1286 1425 1292 1426
rect 110 1420 116 1421
rect 1286 1421 1287 1425
rect 1291 1421 1292 1425
rect 1327 1421 1331 1422
rect 1367 1426 1371 1427
rect 1367 1421 1371 1422
rect 1423 1426 1427 1427
rect 1423 1421 1427 1422
rect 1439 1426 1443 1427
rect 1439 1421 1443 1422
rect 1503 1426 1507 1427
rect 1503 1421 1507 1422
rect 1535 1426 1539 1427
rect 1535 1421 1539 1422
rect 1591 1426 1595 1427
rect 1591 1421 1595 1422
rect 1631 1426 1635 1427
rect 1631 1421 1635 1422
rect 1679 1426 1683 1427
rect 1679 1421 1683 1422
rect 1727 1426 1731 1427
rect 1727 1421 1731 1422
rect 1775 1426 1779 1427
rect 1775 1421 1779 1422
rect 1831 1426 1835 1427
rect 1831 1421 1835 1422
rect 1879 1426 1883 1427
rect 1879 1421 1883 1422
rect 1943 1426 1947 1427
rect 1943 1421 1947 1422
rect 1991 1426 1995 1427
rect 1991 1421 1995 1422
rect 2063 1426 2067 1427
rect 2063 1421 2067 1422
rect 2111 1426 2115 1427
rect 2111 1421 2115 1422
rect 2191 1426 2195 1427
rect 2191 1421 2195 1422
rect 2231 1426 2235 1427
rect 2231 1421 2235 1422
rect 2319 1426 2323 1427
rect 2319 1421 2323 1422
rect 2351 1426 2355 1427
rect 2351 1421 2355 1422
rect 2455 1426 2459 1427
rect 2455 1421 2459 1422
rect 2503 1426 2507 1427
rect 2503 1421 2507 1422
rect 1286 1420 1292 1421
rect 110 1408 116 1409
rect 1286 1408 1292 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 246 1407 252 1408
rect 246 1403 247 1407
rect 251 1403 252 1407
rect 112 1383 114 1403
rect 246 1402 252 1403
rect 334 1407 340 1408
rect 334 1403 335 1407
rect 339 1403 340 1407
rect 334 1402 340 1403
rect 430 1407 436 1408
rect 430 1403 431 1407
rect 435 1403 436 1407
rect 430 1402 436 1403
rect 526 1407 532 1408
rect 526 1403 527 1407
rect 531 1403 532 1407
rect 526 1402 532 1403
rect 630 1407 636 1408
rect 630 1403 631 1407
rect 635 1403 636 1407
rect 630 1402 636 1403
rect 726 1407 732 1408
rect 726 1403 727 1407
rect 731 1403 732 1407
rect 726 1402 732 1403
rect 822 1407 828 1408
rect 822 1403 823 1407
rect 827 1403 828 1407
rect 822 1402 828 1403
rect 910 1407 916 1408
rect 910 1403 911 1407
rect 915 1403 916 1407
rect 910 1402 916 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1102 1407 1108 1408
rect 1102 1403 1103 1407
rect 1107 1403 1108 1407
rect 1286 1404 1287 1408
rect 1291 1404 1292 1408
rect 1286 1403 1292 1404
rect 1102 1402 1108 1403
rect 248 1383 250 1402
rect 336 1383 338 1402
rect 432 1383 434 1402
rect 528 1383 530 1402
rect 632 1383 634 1402
rect 728 1383 730 1402
rect 824 1383 826 1402
rect 912 1383 914 1402
rect 1008 1383 1010 1402
rect 1104 1383 1106 1402
rect 1288 1383 1290 1403
rect 1328 1401 1330 1421
rect 1368 1402 1370 1421
rect 1424 1402 1426 1421
rect 1504 1402 1506 1421
rect 1592 1402 1594 1421
rect 1680 1402 1682 1421
rect 1776 1402 1778 1421
rect 1880 1402 1882 1421
rect 1992 1402 1994 1421
rect 2112 1402 2114 1421
rect 2232 1402 2234 1421
rect 2352 1402 2354 1421
rect 2456 1402 2458 1421
rect 1366 1401 1372 1402
rect 1326 1400 1332 1401
rect 1326 1396 1327 1400
rect 1331 1396 1332 1400
rect 1366 1397 1367 1401
rect 1371 1397 1372 1401
rect 1366 1396 1372 1397
rect 1422 1401 1428 1402
rect 1422 1397 1423 1401
rect 1427 1397 1428 1401
rect 1422 1396 1428 1397
rect 1502 1401 1508 1402
rect 1502 1397 1503 1401
rect 1507 1397 1508 1401
rect 1502 1396 1508 1397
rect 1590 1401 1596 1402
rect 1590 1397 1591 1401
rect 1595 1397 1596 1401
rect 1590 1396 1596 1397
rect 1678 1401 1684 1402
rect 1678 1397 1679 1401
rect 1683 1397 1684 1401
rect 1678 1396 1684 1397
rect 1774 1401 1780 1402
rect 1774 1397 1775 1401
rect 1779 1397 1780 1401
rect 1774 1396 1780 1397
rect 1878 1401 1884 1402
rect 1878 1397 1879 1401
rect 1883 1397 1884 1401
rect 1878 1396 1884 1397
rect 1990 1401 1996 1402
rect 1990 1397 1991 1401
rect 1995 1397 1996 1401
rect 1990 1396 1996 1397
rect 2110 1401 2116 1402
rect 2110 1397 2111 1401
rect 2115 1397 2116 1401
rect 2110 1396 2116 1397
rect 2230 1401 2236 1402
rect 2230 1397 2231 1401
rect 2235 1397 2236 1401
rect 2230 1396 2236 1397
rect 2350 1401 2356 1402
rect 2350 1397 2351 1401
rect 2355 1397 2356 1401
rect 2350 1396 2356 1397
rect 2454 1401 2460 1402
rect 2504 1401 2506 1421
rect 2454 1397 2455 1401
rect 2459 1397 2460 1401
rect 2454 1396 2460 1397
rect 2502 1400 2508 1401
rect 2502 1396 2503 1400
rect 2507 1396 2508 1400
rect 1326 1395 1332 1396
rect 2502 1395 2508 1396
rect 1326 1383 1332 1384
rect 111 1382 115 1383
rect 111 1377 115 1378
rect 151 1382 155 1383
rect 151 1377 155 1378
rect 215 1382 219 1383
rect 215 1377 219 1378
rect 247 1382 251 1383
rect 247 1377 251 1378
rect 311 1382 315 1383
rect 311 1377 315 1378
rect 335 1382 339 1383
rect 335 1377 339 1378
rect 407 1382 411 1383
rect 407 1377 411 1378
rect 431 1382 435 1383
rect 431 1377 435 1378
rect 511 1382 515 1383
rect 511 1377 515 1378
rect 527 1382 531 1383
rect 527 1377 531 1378
rect 607 1382 611 1383
rect 607 1377 611 1378
rect 631 1382 635 1383
rect 631 1377 635 1378
rect 703 1382 707 1383
rect 703 1377 707 1378
rect 727 1382 731 1383
rect 727 1377 731 1378
rect 799 1382 803 1383
rect 799 1377 803 1378
rect 823 1382 827 1383
rect 823 1377 827 1378
rect 895 1382 899 1383
rect 895 1377 899 1378
rect 911 1382 915 1383
rect 911 1377 915 1378
rect 999 1382 1003 1383
rect 999 1377 1003 1378
rect 1007 1382 1011 1383
rect 1007 1377 1011 1378
rect 1103 1382 1107 1383
rect 1103 1377 1107 1378
rect 1287 1382 1291 1383
rect 1326 1379 1327 1383
rect 1331 1379 1332 1383
rect 2502 1383 2508 1384
rect 1326 1378 1332 1379
rect 1350 1380 1356 1381
rect 1287 1377 1291 1378
rect 112 1357 114 1377
rect 152 1358 154 1377
rect 216 1358 218 1377
rect 312 1358 314 1377
rect 408 1358 410 1377
rect 512 1358 514 1377
rect 608 1358 610 1377
rect 704 1358 706 1377
rect 800 1358 802 1377
rect 896 1358 898 1377
rect 1000 1358 1002 1377
rect 150 1357 156 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 150 1353 151 1357
rect 155 1353 156 1357
rect 150 1352 156 1353
rect 214 1357 220 1358
rect 214 1353 215 1357
rect 219 1353 220 1357
rect 214 1352 220 1353
rect 310 1357 316 1358
rect 310 1353 311 1357
rect 315 1353 316 1357
rect 310 1352 316 1353
rect 406 1357 412 1358
rect 406 1353 407 1357
rect 411 1353 412 1357
rect 406 1352 412 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 606 1357 612 1358
rect 606 1353 607 1357
rect 611 1353 612 1357
rect 606 1352 612 1353
rect 702 1357 708 1358
rect 702 1353 703 1357
rect 707 1353 708 1357
rect 702 1352 708 1353
rect 798 1357 804 1358
rect 798 1353 799 1357
rect 803 1353 804 1357
rect 798 1352 804 1353
rect 894 1357 900 1358
rect 894 1353 895 1357
rect 899 1353 900 1357
rect 894 1352 900 1353
rect 998 1357 1004 1358
rect 1288 1357 1290 1377
rect 1328 1371 1330 1378
rect 1350 1376 1351 1380
rect 1355 1376 1356 1380
rect 1350 1375 1356 1376
rect 1406 1380 1412 1381
rect 1406 1376 1407 1380
rect 1411 1376 1412 1380
rect 1406 1375 1412 1376
rect 1486 1380 1492 1381
rect 1486 1376 1487 1380
rect 1491 1376 1492 1380
rect 1486 1375 1492 1376
rect 1574 1380 1580 1381
rect 1574 1376 1575 1380
rect 1579 1376 1580 1380
rect 1574 1375 1580 1376
rect 1662 1380 1668 1381
rect 1662 1376 1663 1380
rect 1667 1376 1668 1380
rect 1662 1375 1668 1376
rect 1758 1380 1764 1381
rect 1758 1376 1759 1380
rect 1763 1376 1764 1380
rect 1758 1375 1764 1376
rect 1862 1380 1868 1381
rect 1862 1376 1863 1380
rect 1867 1376 1868 1380
rect 1862 1375 1868 1376
rect 1974 1380 1980 1381
rect 1974 1376 1975 1380
rect 1979 1376 1980 1380
rect 1974 1375 1980 1376
rect 2094 1380 2100 1381
rect 2094 1376 2095 1380
rect 2099 1376 2100 1380
rect 2094 1375 2100 1376
rect 2214 1380 2220 1381
rect 2214 1376 2215 1380
rect 2219 1376 2220 1380
rect 2214 1375 2220 1376
rect 2334 1380 2340 1381
rect 2334 1376 2335 1380
rect 2339 1376 2340 1380
rect 2334 1375 2340 1376
rect 2438 1380 2444 1381
rect 2438 1376 2439 1380
rect 2443 1376 2444 1380
rect 2502 1379 2503 1383
rect 2507 1379 2508 1383
rect 2502 1378 2508 1379
rect 2438 1375 2444 1376
rect 1352 1371 1354 1375
rect 1408 1371 1410 1375
rect 1488 1371 1490 1375
rect 1576 1371 1578 1375
rect 1664 1371 1666 1375
rect 1760 1371 1762 1375
rect 1864 1371 1866 1375
rect 1976 1371 1978 1375
rect 2096 1371 2098 1375
rect 2216 1371 2218 1375
rect 2336 1371 2338 1375
rect 2440 1371 2442 1375
rect 2504 1371 2506 1378
rect 1327 1370 1331 1371
rect 1327 1365 1331 1366
rect 1351 1370 1355 1371
rect 1351 1365 1355 1366
rect 1407 1370 1411 1371
rect 1407 1365 1411 1366
rect 1479 1370 1483 1371
rect 1479 1365 1483 1366
rect 1487 1370 1491 1371
rect 1487 1365 1491 1366
rect 1567 1370 1571 1371
rect 1567 1365 1571 1366
rect 1575 1370 1579 1371
rect 1575 1365 1579 1366
rect 1655 1370 1659 1371
rect 1655 1365 1659 1366
rect 1663 1370 1667 1371
rect 1663 1365 1667 1366
rect 1751 1370 1755 1371
rect 1751 1365 1755 1366
rect 1759 1370 1763 1371
rect 1759 1365 1763 1366
rect 1855 1370 1859 1371
rect 1855 1365 1859 1366
rect 1863 1370 1867 1371
rect 1863 1365 1867 1366
rect 1967 1370 1971 1371
rect 1967 1365 1971 1366
rect 1975 1370 1979 1371
rect 1975 1365 1979 1366
rect 2079 1370 2083 1371
rect 2079 1365 2083 1366
rect 2095 1370 2099 1371
rect 2095 1365 2099 1366
rect 2199 1370 2203 1371
rect 2199 1365 2203 1366
rect 2215 1370 2219 1371
rect 2215 1365 2219 1366
rect 2327 1370 2331 1371
rect 2327 1365 2331 1366
rect 2335 1370 2339 1371
rect 2335 1365 2339 1366
rect 2439 1370 2443 1371
rect 2439 1365 2443 1366
rect 2503 1370 2507 1371
rect 2503 1365 2507 1366
rect 1328 1362 1330 1365
rect 1350 1364 1356 1365
rect 1326 1361 1332 1362
rect 1326 1357 1327 1361
rect 1331 1357 1332 1361
rect 1350 1360 1351 1364
rect 1355 1360 1356 1364
rect 1350 1359 1356 1360
rect 1406 1364 1412 1365
rect 1406 1360 1407 1364
rect 1411 1360 1412 1364
rect 1406 1359 1412 1360
rect 1478 1364 1484 1365
rect 1478 1360 1479 1364
rect 1483 1360 1484 1364
rect 1478 1359 1484 1360
rect 1566 1364 1572 1365
rect 1566 1360 1567 1364
rect 1571 1360 1572 1364
rect 1566 1359 1572 1360
rect 1654 1364 1660 1365
rect 1654 1360 1655 1364
rect 1659 1360 1660 1364
rect 1654 1359 1660 1360
rect 1750 1364 1756 1365
rect 1750 1360 1751 1364
rect 1755 1360 1756 1364
rect 1750 1359 1756 1360
rect 1854 1364 1860 1365
rect 1854 1360 1855 1364
rect 1859 1360 1860 1364
rect 1854 1359 1860 1360
rect 1966 1364 1972 1365
rect 1966 1360 1967 1364
rect 1971 1360 1972 1364
rect 1966 1359 1972 1360
rect 2078 1364 2084 1365
rect 2078 1360 2079 1364
rect 2083 1360 2084 1364
rect 2078 1359 2084 1360
rect 2198 1364 2204 1365
rect 2198 1360 2199 1364
rect 2203 1360 2204 1364
rect 2198 1359 2204 1360
rect 2326 1364 2332 1365
rect 2326 1360 2327 1364
rect 2331 1360 2332 1364
rect 2326 1359 2332 1360
rect 2438 1364 2444 1365
rect 2438 1360 2439 1364
rect 2443 1360 2444 1364
rect 2504 1362 2506 1365
rect 2438 1359 2444 1360
rect 2502 1361 2508 1362
rect 998 1353 999 1357
rect 1003 1353 1004 1357
rect 998 1352 1004 1353
rect 1286 1356 1292 1357
rect 1326 1356 1332 1357
rect 2502 1357 2503 1361
rect 2507 1357 2508 1361
rect 2502 1356 2508 1357
rect 1286 1352 1287 1356
rect 1291 1352 1292 1356
rect 110 1351 116 1352
rect 1286 1351 1292 1352
rect 1326 1344 1332 1345
rect 2502 1344 2508 1345
rect 1326 1340 1327 1344
rect 1331 1340 1332 1344
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 1286 1339 1292 1340
rect 1326 1339 1332 1340
rect 1366 1343 1372 1344
rect 1366 1339 1367 1343
rect 1371 1339 1372 1343
rect 110 1334 116 1335
rect 134 1336 140 1337
rect 112 1331 114 1334
rect 134 1332 135 1336
rect 139 1332 140 1336
rect 134 1331 140 1332
rect 198 1336 204 1337
rect 198 1332 199 1336
rect 203 1332 204 1336
rect 198 1331 204 1332
rect 294 1336 300 1337
rect 294 1332 295 1336
rect 299 1332 300 1336
rect 294 1331 300 1332
rect 390 1336 396 1337
rect 390 1332 391 1336
rect 395 1332 396 1336
rect 390 1331 396 1332
rect 494 1336 500 1337
rect 494 1332 495 1336
rect 499 1332 500 1336
rect 494 1331 500 1332
rect 590 1336 596 1337
rect 590 1332 591 1336
rect 595 1332 596 1336
rect 590 1331 596 1332
rect 686 1336 692 1337
rect 686 1332 687 1336
rect 691 1332 692 1336
rect 686 1331 692 1332
rect 782 1336 788 1337
rect 782 1332 783 1336
rect 787 1332 788 1336
rect 782 1331 788 1332
rect 878 1336 884 1337
rect 878 1332 879 1336
rect 883 1332 884 1336
rect 878 1331 884 1332
rect 982 1336 988 1337
rect 982 1332 983 1336
rect 987 1332 988 1336
rect 1286 1335 1287 1339
rect 1291 1335 1292 1339
rect 1286 1334 1292 1335
rect 982 1331 988 1332
rect 1288 1331 1290 1334
rect 111 1330 115 1331
rect 111 1325 115 1326
rect 135 1330 139 1331
rect 135 1325 139 1326
rect 199 1330 203 1331
rect 199 1325 203 1326
rect 215 1330 219 1331
rect 215 1325 219 1326
rect 295 1330 299 1331
rect 295 1325 299 1326
rect 319 1330 323 1331
rect 319 1325 323 1326
rect 391 1330 395 1331
rect 391 1325 395 1326
rect 415 1330 419 1331
rect 415 1325 419 1326
rect 495 1330 499 1331
rect 495 1325 499 1326
rect 511 1330 515 1331
rect 511 1325 515 1326
rect 591 1330 595 1331
rect 591 1325 595 1326
rect 599 1330 603 1331
rect 599 1325 603 1326
rect 687 1330 691 1331
rect 687 1325 691 1326
rect 783 1330 787 1331
rect 783 1325 787 1326
rect 879 1330 883 1331
rect 879 1325 883 1326
rect 983 1330 987 1331
rect 983 1325 987 1326
rect 1287 1330 1291 1331
rect 1287 1325 1291 1326
rect 112 1322 114 1325
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 414 1324 420 1325
rect 414 1320 415 1324
rect 419 1320 420 1324
rect 414 1319 420 1320
rect 510 1324 516 1325
rect 510 1320 511 1324
rect 515 1320 516 1324
rect 510 1319 516 1320
rect 598 1324 604 1325
rect 598 1320 599 1324
rect 603 1320 604 1324
rect 598 1319 604 1320
rect 686 1324 692 1325
rect 686 1320 687 1324
rect 691 1320 692 1324
rect 686 1319 692 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 878 1324 884 1325
rect 878 1320 879 1324
rect 883 1320 884 1324
rect 1288 1322 1290 1325
rect 878 1319 884 1320
rect 1286 1321 1292 1322
rect 110 1316 116 1317
rect 1286 1317 1287 1321
rect 1291 1317 1292 1321
rect 1286 1316 1292 1317
rect 1328 1311 1330 1339
rect 1366 1338 1372 1339
rect 1422 1343 1428 1344
rect 1422 1339 1423 1343
rect 1427 1339 1428 1343
rect 1422 1338 1428 1339
rect 1494 1343 1500 1344
rect 1494 1339 1495 1343
rect 1499 1339 1500 1343
rect 1494 1338 1500 1339
rect 1582 1343 1588 1344
rect 1582 1339 1583 1343
rect 1587 1339 1588 1343
rect 1582 1338 1588 1339
rect 1670 1343 1676 1344
rect 1670 1339 1671 1343
rect 1675 1339 1676 1343
rect 1670 1338 1676 1339
rect 1766 1343 1772 1344
rect 1766 1339 1767 1343
rect 1771 1339 1772 1343
rect 1766 1338 1772 1339
rect 1870 1343 1876 1344
rect 1870 1339 1871 1343
rect 1875 1339 1876 1343
rect 1870 1338 1876 1339
rect 1982 1343 1988 1344
rect 1982 1339 1983 1343
rect 1987 1339 1988 1343
rect 1982 1338 1988 1339
rect 2094 1343 2100 1344
rect 2094 1339 2095 1343
rect 2099 1339 2100 1343
rect 2094 1338 2100 1339
rect 2214 1343 2220 1344
rect 2214 1339 2215 1343
rect 2219 1339 2220 1343
rect 2214 1338 2220 1339
rect 2342 1343 2348 1344
rect 2342 1339 2343 1343
rect 2347 1339 2348 1343
rect 2342 1338 2348 1339
rect 2454 1343 2460 1344
rect 2454 1339 2455 1343
rect 2459 1339 2460 1343
rect 2502 1340 2503 1344
rect 2507 1340 2508 1344
rect 2502 1339 2508 1340
rect 2454 1338 2460 1339
rect 1368 1311 1370 1338
rect 1424 1311 1426 1338
rect 1496 1311 1498 1338
rect 1584 1311 1586 1338
rect 1672 1311 1674 1338
rect 1768 1311 1770 1338
rect 1872 1311 1874 1338
rect 1984 1311 1986 1338
rect 2096 1311 2098 1338
rect 2216 1311 2218 1338
rect 2344 1311 2346 1338
rect 2456 1311 2458 1338
rect 2504 1311 2506 1339
rect 1327 1310 1331 1311
rect 1327 1305 1331 1306
rect 1367 1310 1371 1311
rect 1367 1305 1371 1306
rect 1423 1310 1427 1311
rect 1423 1305 1427 1306
rect 1495 1310 1499 1311
rect 1495 1305 1499 1306
rect 1519 1310 1523 1311
rect 1519 1305 1523 1306
rect 1583 1310 1587 1311
rect 1583 1305 1587 1306
rect 1615 1310 1619 1311
rect 1615 1305 1619 1306
rect 1671 1310 1675 1311
rect 1671 1305 1675 1306
rect 1719 1310 1723 1311
rect 1719 1305 1723 1306
rect 1767 1310 1771 1311
rect 1767 1305 1771 1306
rect 1823 1310 1827 1311
rect 1823 1305 1827 1306
rect 1871 1310 1875 1311
rect 1871 1305 1875 1306
rect 1919 1310 1923 1311
rect 1919 1305 1923 1306
rect 1983 1310 1987 1311
rect 1983 1305 1987 1306
rect 2015 1310 2019 1311
rect 2015 1305 2019 1306
rect 2095 1310 2099 1311
rect 2095 1305 2099 1306
rect 2103 1310 2107 1311
rect 2103 1305 2107 1306
rect 2183 1310 2187 1311
rect 2183 1305 2187 1306
rect 2215 1310 2219 1311
rect 2215 1305 2219 1306
rect 2255 1310 2259 1311
rect 2255 1305 2259 1306
rect 2327 1310 2331 1311
rect 2327 1305 2331 1306
rect 2343 1310 2347 1311
rect 2343 1305 2347 1306
rect 2399 1310 2403 1311
rect 2399 1305 2403 1306
rect 2455 1310 2459 1311
rect 2455 1305 2459 1306
rect 2503 1310 2507 1311
rect 2503 1305 2507 1306
rect 110 1304 116 1305
rect 1286 1304 1292 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 150 1303 156 1304
rect 150 1299 151 1303
rect 155 1299 156 1303
rect 112 1279 114 1299
rect 150 1298 156 1299
rect 230 1303 236 1304
rect 230 1299 231 1303
rect 235 1299 236 1303
rect 230 1298 236 1299
rect 334 1303 340 1304
rect 334 1299 335 1303
rect 339 1299 340 1303
rect 334 1298 340 1299
rect 430 1303 436 1304
rect 430 1299 431 1303
rect 435 1299 436 1303
rect 430 1298 436 1299
rect 526 1303 532 1304
rect 526 1299 527 1303
rect 531 1299 532 1303
rect 526 1298 532 1299
rect 614 1303 620 1304
rect 614 1299 615 1303
rect 619 1299 620 1303
rect 614 1298 620 1299
rect 702 1303 708 1304
rect 702 1299 703 1303
rect 707 1299 708 1303
rect 702 1298 708 1299
rect 798 1303 804 1304
rect 798 1299 799 1303
rect 803 1299 804 1303
rect 798 1298 804 1299
rect 894 1303 900 1304
rect 894 1299 895 1303
rect 899 1299 900 1303
rect 1286 1300 1287 1304
rect 1291 1300 1292 1304
rect 1286 1299 1292 1300
rect 894 1298 900 1299
rect 152 1279 154 1298
rect 232 1279 234 1298
rect 336 1279 338 1298
rect 432 1279 434 1298
rect 528 1279 530 1298
rect 616 1279 618 1298
rect 704 1279 706 1298
rect 800 1279 802 1298
rect 896 1279 898 1298
rect 1288 1279 1290 1299
rect 1328 1285 1330 1305
rect 1368 1286 1370 1305
rect 1424 1286 1426 1305
rect 1520 1286 1522 1305
rect 1616 1286 1618 1305
rect 1720 1286 1722 1305
rect 1824 1286 1826 1305
rect 1920 1286 1922 1305
rect 2016 1286 2018 1305
rect 2104 1286 2106 1305
rect 2184 1286 2186 1305
rect 2256 1286 2258 1305
rect 2328 1286 2330 1305
rect 2400 1286 2402 1305
rect 2456 1286 2458 1305
rect 1366 1285 1372 1286
rect 1326 1284 1332 1285
rect 1326 1280 1327 1284
rect 1331 1280 1332 1284
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 1422 1285 1428 1286
rect 1422 1281 1423 1285
rect 1427 1281 1428 1285
rect 1422 1280 1428 1281
rect 1518 1285 1524 1286
rect 1518 1281 1519 1285
rect 1523 1281 1524 1285
rect 1518 1280 1524 1281
rect 1614 1285 1620 1286
rect 1614 1281 1615 1285
rect 1619 1281 1620 1285
rect 1614 1280 1620 1281
rect 1718 1285 1724 1286
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1718 1280 1724 1281
rect 1822 1285 1828 1286
rect 1822 1281 1823 1285
rect 1827 1281 1828 1285
rect 1822 1280 1828 1281
rect 1918 1285 1924 1286
rect 1918 1281 1919 1285
rect 1923 1281 1924 1285
rect 1918 1280 1924 1281
rect 2014 1285 2020 1286
rect 2014 1281 2015 1285
rect 2019 1281 2020 1285
rect 2014 1280 2020 1281
rect 2102 1285 2108 1286
rect 2102 1281 2103 1285
rect 2107 1281 2108 1285
rect 2102 1280 2108 1281
rect 2182 1285 2188 1286
rect 2182 1281 2183 1285
rect 2187 1281 2188 1285
rect 2182 1280 2188 1281
rect 2254 1285 2260 1286
rect 2254 1281 2255 1285
rect 2259 1281 2260 1285
rect 2254 1280 2260 1281
rect 2326 1285 2332 1286
rect 2326 1281 2327 1285
rect 2331 1281 2332 1285
rect 2326 1280 2332 1281
rect 2398 1285 2404 1286
rect 2398 1281 2399 1285
rect 2403 1281 2404 1285
rect 2398 1280 2404 1281
rect 2454 1285 2460 1286
rect 2504 1285 2506 1305
rect 2454 1281 2455 1285
rect 2459 1281 2460 1285
rect 2454 1280 2460 1281
rect 2502 1284 2508 1285
rect 2502 1280 2503 1284
rect 2507 1280 2508 1284
rect 1326 1279 1332 1280
rect 2502 1279 2508 1280
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 151 1278 155 1279
rect 151 1273 155 1274
rect 191 1278 195 1279
rect 191 1273 195 1274
rect 231 1278 235 1279
rect 231 1273 235 1274
rect 247 1278 251 1279
rect 247 1273 251 1274
rect 303 1278 307 1279
rect 303 1273 307 1274
rect 335 1278 339 1279
rect 335 1273 339 1274
rect 367 1278 371 1279
rect 367 1273 371 1274
rect 431 1278 435 1279
rect 431 1273 435 1274
rect 439 1278 443 1279
rect 439 1273 443 1274
rect 527 1278 531 1279
rect 527 1273 531 1274
rect 615 1278 619 1279
rect 615 1273 619 1274
rect 639 1278 643 1279
rect 639 1273 643 1274
rect 703 1278 707 1279
rect 703 1273 707 1274
rect 775 1278 779 1279
rect 775 1273 779 1274
rect 799 1278 803 1279
rect 799 1273 803 1274
rect 895 1278 899 1279
rect 895 1273 899 1274
rect 927 1278 931 1279
rect 927 1273 931 1274
rect 1095 1278 1099 1279
rect 1095 1273 1099 1274
rect 1239 1278 1243 1279
rect 1239 1273 1243 1274
rect 1287 1278 1291 1279
rect 1287 1273 1291 1274
rect 112 1253 114 1273
rect 192 1254 194 1273
rect 248 1254 250 1273
rect 304 1254 306 1273
rect 368 1254 370 1273
rect 440 1254 442 1273
rect 528 1254 530 1273
rect 640 1254 642 1273
rect 776 1254 778 1273
rect 928 1254 930 1273
rect 1096 1254 1098 1273
rect 1240 1254 1242 1273
rect 190 1253 196 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 190 1249 191 1253
rect 195 1249 196 1253
rect 190 1248 196 1249
rect 246 1253 252 1254
rect 246 1249 247 1253
rect 251 1249 252 1253
rect 246 1248 252 1249
rect 302 1253 308 1254
rect 302 1249 303 1253
rect 307 1249 308 1253
rect 302 1248 308 1249
rect 366 1253 372 1254
rect 366 1249 367 1253
rect 371 1249 372 1253
rect 366 1248 372 1249
rect 438 1253 444 1254
rect 438 1249 439 1253
rect 443 1249 444 1253
rect 438 1248 444 1249
rect 526 1253 532 1254
rect 526 1249 527 1253
rect 531 1249 532 1253
rect 526 1248 532 1249
rect 638 1253 644 1254
rect 638 1249 639 1253
rect 643 1249 644 1253
rect 638 1248 644 1249
rect 774 1253 780 1254
rect 774 1249 775 1253
rect 779 1249 780 1253
rect 774 1248 780 1249
rect 926 1253 932 1254
rect 926 1249 927 1253
rect 931 1249 932 1253
rect 926 1248 932 1249
rect 1094 1253 1100 1254
rect 1094 1249 1095 1253
rect 1099 1249 1100 1253
rect 1094 1248 1100 1249
rect 1238 1253 1244 1254
rect 1288 1253 1290 1273
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1263 1332 1267
rect 2502 1267 2508 1268
rect 1326 1262 1332 1263
rect 1350 1264 1356 1265
rect 1238 1249 1239 1253
rect 1243 1249 1244 1253
rect 1238 1248 1244 1249
rect 1286 1252 1292 1253
rect 1286 1248 1287 1252
rect 1291 1248 1292 1252
rect 110 1247 116 1248
rect 1286 1247 1292 1248
rect 1328 1243 1330 1262
rect 1350 1260 1351 1264
rect 1355 1260 1356 1264
rect 1350 1259 1356 1260
rect 1406 1264 1412 1265
rect 1406 1260 1407 1264
rect 1411 1260 1412 1264
rect 1406 1259 1412 1260
rect 1502 1264 1508 1265
rect 1502 1260 1503 1264
rect 1507 1260 1508 1264
rect 1502 1259 1508 1260
rect 1598 1264 1604 1265
rect 1598 1260 1599 1264
rect 1603 1260 1604 1264
rect 1598 1259 1604 1260
rect 1702 1264 1708 1265
rect 1702 1260 1703 1264
rect 1707 1260 1708 1264
rect 1702 1259 1708 1260
rect 1806 1264 1812 1265
rect 1806 1260 1807 1264
rect 1811 1260 1812 1264
rect 1806 1259 1812 1260
rect 1902 1264 1908 1265
rect 1902 1260 1903 1264
rect 1907 1260 1908 1264
rect 1902 1259 1908 1260
rect 1998 1264 2004 1265
rect 1998 1260 1999 1264
rect 2003 1260 2004 1264
rect 1998 1259 2004 1260
rect 2086 1264 2092 1265
rect 2086 1260 2087 1264
rect 2091 1260 2092 1264
rect 2086 1259 2092 1260
rect 2166 1264 2172 1265
rect 2166 1260 2167 1264
rect 2171 1260 2172 1264
rect 2166 1259 2172 1260
rect 2238 1264 2244 1265
rect 2238 1260 2239 1264
rect 2243 1260 2244 1264
rect 2238 1259 2244 1260
rect 2310 1264 2316 1265
rect 2310 1260 2311 1264
rect 2315 1260 2316 1264
rect 2310 1259 2316 1260
rect 2382 1264 2388 1265
rect 2382 1260 2383 1264
rect 2387 1260 2388 1264
rect 2382 1259 2388 1260
rect 2438 1264 2444 1265
rect 2438 1260 2439 1264
rect 2443 1260 2444 1264
rect 2502 1263 2503 1267
rect 2507 1263 2508 1267
rect 2502 1262 2508 1263
rect 2438 1259 2444 1260
rect 1352 1243 1354 1259
rect 1408 1243 1410 1259
rect 1504 1243 1506 1259
rect 1600 1243 1602 1259
rect 1704 1243 1706 1259
rect 1808 1243 1810 1259
rect 1904 1243 1906 1259
rect 2000 1243 2002 1259
rect 2088 1243 2090 1259
rect 2168 1243 2170 1259
rect 2240 1243 2242 1259
rect 2312 1243 2314 1259
rect 2384 1243 2386 1259
rect 2440 1243 2442 1259
rect 2504 1243 2506 1262
rect 1327 1242 1331 1243
rect 1327 1237 1331 1238
rect 1351 1242 1355 1243
rect 1351 1237 1355 1238
rect 1407 1242 1411 1243
rect 1407 1237 1411 1238
rect 1447 1242 1451 1243
rect 1447 1237 1451 1238
rect 1503 1242 1507 1243
rect 1503 1237 1507 1238
rect 1575 1242 1579 1243
rect 1575 1237 1579 1238
rect 1599 1242 1603 1243
rect 1599 1237 1603 1238
rect 1695 1242 1699 1243
rect 1695 1237 1699 1238
rect 1703 1242 1707 1243
rect 1703 1237 1707 1238
rect 1807 1242 1811 1243
rect 1807 1237 1811 1238
rect 1815 1242 1819 1243
rect 1815 1237 1819 1238
rect 1903 1242 1907 1243
rect 1903 1237 1907 1238
rect 1927 1242 1931 1243
rect 1927 1237 1931 1238
rect 1999 1242 2003 1243
rect 1999 1237 2003 1238
rect 2031 1242 2035 1243
rect 2031 1237 2035 1238
rect 2087 1242 2091 1243
rect 2087 1237 2091 1238
rect 2127 1242 2131 1243
rect 2127 1237 2131 1238
rect 2167 1242 2171 1243
rect 2167 1237 2171 1238
rect 2215 1242 2219 1243
rect 2215 1237 2219 1238
rect 2239 1242 2243 1243
rect 2239 1237 2243 1238
rect 2295 1242 2299 1243
rect 2295 1237 2299 1238
rect 2311 1242 2315 1243
rect 2311 1237 2315 1238
rect 2375 1242 2379 1243
rect 2375 1237 2379 1238
rect 2383 1242 2387 1243
rect 2383 1237 2387 1238
rect 2439 1242 2443 1243
rect 2439 1237 2443 1238
rect 2503 1242 2507 1243
rect 2503 1237 2507 1238
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1286 1235 1292 1236
rect 110 1230 116 1231
rect 174 1232 180 1233
rect 112 1227 114 1230
rect 174 1228 175 1232
rect 179 1228 180 1232
rect 174 1227 180 1228
rect 230 1232 236 1233
rect 230 1228 231 1232
rect 235 1228 236 1232
rect 230 1227 236 1228
rect 286 1232 292 1233
rect 286 1228 287 1232
rect 291 1228 292 1232
rect 286 1227 292 1228
rect 350 1232 356 1233
rect 350 1228 351 1232
rect 355 1228 356 1232
rect 350 1227 356 1228
rect 422 1232 428 1233
rect 422 1228 423 1232
rect 427 1228 428 1232
rect 422 1227 428 1228
rect 510 1232 516 1233
rect 510 1228 511 1232
rect 515 1228 516 1232
rect 510 1227 516 1228
rect 622 1232 628 1233
rect 622 1228 623 1232
rect 627 1228 628 1232
rect 622 1227 628 1228
rect 758 1232 764 1233
rect 758 1228 759 1232
rect 763 1228 764 1232
rect 758 1227 764 1228
rect 910 1232 916 1233
rect 910 1228 911 1232
rect 915 1228 916 1232
rect 910 1227 916 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1222 1232 1228 1233
rect 1222 1228 1223 1232
rect 1227 1228 1228 1232
rect 1286 1231 1287 1235
rect 1291 1231 1292 1235
rect 1328 1234 1330 1237
rect 1350 1236 1356 1237
rect 1286 1230 1292 1231
rect 1326 1233 1332 1234
rect 1222 1227 1228 1228
rect 1288 1227 1290 1230
rect 1326 1229 1327 1233
rect 1331 1229 1332 1233
rect 1350 1232 1351 1236
rect 1355 1232 1356 1236
rect 1350 1231 1356 1232
rect 1446 1236 1452 1237
rect 1446 1232 1447 1236
rect 1451 1232 1452 1236
rect 1446 1231 1452 1232
rect 1574 1236 1580 1237
rect 1574 1232 1575 1236
rect 1579 1232 1580 1236
rect 1574 1231 1580 1232
rect 1694 1236 1700 1237
rect 1694 1232 1695 1236
rect 1699 1232 1700 1236
rect 1694 1231 1700 1232
rect 1814 1236 1820 1237
rect 1814 1232 1815 1236
rect 1819 1232 1820 1236
rect 1814 1231 1820 1232
rect 1926 1236 1932 1237
rect 1926 1232 1927 1236
rect 1931 1232 1932 1236
rect 1926 1231 1932 1232
rect 2030 1236 2036 1237
rect 2030 1232 2031 1236
rect 2035 1232 2036 1236
rect 2030 1231 2036 1232
rect 2126 1236 2132 1237
rect 2126 1232 2127 1236
rect 2131 1232 2132 1236
rect 2126 1231 2132 1232
rect 2214 1236 2220 1237
rect 2214 1232 2215 1236
rect 2219 1232 2220 1236
rect 2214 1231 2220 1232
rect 2294 1236 2300 1237
rect 2294 1232 2295 1236
rect 2299 1232 2300 1236
rect 2294 1231 2300 1232
rect 2374 1236 2380 1237
rect 2374 1232 2375 1236
rect 2379 1232 2380 1236
rect 2374 1231 2380 1232
rect 2438 1236 2444 1237
rect 2438 1232 2439 1236
rect 2443 1232 2444 1236
rect 2504 1234 2506 1237
rect 2438 1231 2444 1232
rect 2502 1233 2508 1234
rect 1326 1228 1332 1229
rect 2502 1229 2503 1233
rect 2507 1229 2508 1233
rect 2502 1228 2508 1229
rect 111 1226 115 1227
rect 111 1221 115 1222
rect 175 1226 179 1227
rect 175 1221 179 1222
rect 231 1226 235 1227
rect 231 1221 235 1222
rect 287 1226 291 1227
rect 287 1221 291 1222
rect 351 1226 355 1227
rect 351 1221 355 1222
rect 407 1226 411 1227
rect 407 1221 411 1222
rect 423 1226 427 1227
rect 423 1221 427 1222
rect 463 1226 467 1227
rect 463 1221 467 1222
rect 511 1226 515 1227
rect 511 1221 515 1222
rect 519 1226 523 1227
rect 519 1221 523 1222
rect 575 1226 579 1227
rect 575 1221 579 1222
rect 623 1226 627 1227
rect 623 1221 627 1222
rect 631 1226 635 1227
rect 631 1221 635 1222
rect 687 1226 691 1227
rect 687 1221 691 1222
rect 743 1226 747 1227
rect 743 1221 747 1222
rect 759 1226 763 1227
rect 759 1221 763 1222
rect 799 1226 803 1227
rect 799 1221 803 1222
rect 855 1226 859 1227
rect 855 1221 859 1222
rect 911 1226 915 1227
rect 911 1221 915 1222
rect 1079 1226 1083 1227
rect 1079 1221 1083 1222
rect 1223 1226 1227 1227
rect 1223 1221 1227 1222
rect 1287 1226 1291 1227
rect 1287 1221 1291 1222
rect 112 1218 114 1221
rect 350 1220 356 1221
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 350 1216 351 1220
rect 355 1216 356 1220
rect 350 1215 356 1216
rect 406 1220 412 1221
rect 406 1216 407 1220
rect 411 1216 412 1220
rect 406 1215 412 1216
rect 462 1220 468 1221
rect 462 1216 463 1220
rect 467 1216 468 1220
rect 462 1215 468 1216
rect 518 1220 524 1221
rect 518 1216 519 1220
rect 523 1216 524 1220
rect 518 1215 524 1216
rect 574 1220 580 1221
rect 574 1216 575 1220
rect 579 1216 580 1220
rect 574 1215 580 1216
rect 630 1220 636 1221
rect 630 1216 631 1220
rect 635 1216 636 1220
rect 630 1215 636 1216
rect 686 1220 692 1221
rect 686 1216 687 1220
rect 691 1216 692 1220
rect 686 1215 692 1216
rect 742 1220 748 1221
rect 742 1216 743 1220
rect 747 1216 748 1220
rect 742 1215 748 1216
rect 798 1220 804 1221
rect 798 1216 799 1220
rect 803 1216 804 1220
rect 798 1215 804 1216
rect 854 1220 860 1221
rect 854 1216 855 1220
rect 859 1216 860 1220
rect 854 1215 860 1216
rect 910 1220 916 1221
rect 910 1216 911 1220
rect 915 1216 916 1220
rect 1288 1218 1290 1221
rect 910 1215 916 1216
rect 1286 1217 1292 1218
rect 110 1212 116 1213
rect 1286 1213 1287 1217
rect 1291 1213 1292 1217
rect 1286 1212 1292 1213
rect 1326 1216 1332 1217
rect 2502 1216 2508 1217
rect 1326 1212 1327 1216
rect 1331 1212 1332 1216
rect 1326 1211 1332 1212
rect 1366 1215 1372 1216
rect 1366 1211 1367 1215
rect 1371 1211 1372 1215
rect 110 1200 116 1201
rect 1286 1200 1292 1201
rect 110 1196 111 1200
rect 115 1196 116 1200
rect 110 1195 116 1196
rect 366 1199 372 1200
rect 366 1195 367 1199
rect 371 1195 372 1199
rect 112 1171 114 1195
rect 366 1194 372 1195
rect 422 1199 428 1200
rect 422 1195 423 1199
rect 427 1195 428 1199
rect 422 1194 428 1195
rect 478 1199 484 1200
rect 478 1195 479 1199
rect 483 1195 484 1199
rect 478 1194 484 1195
rect 534 1199 540 1200
rect 534 1195 535 1199
rect 539 1195 540 1199
rect 534 1194 540 1195
rect 590 1199 596 1200
rect 590 1195 591 1199
rect 595 1195 596 1199
rect 590 1194 596 1195
rect 646 1199 652 1200
rect 646 1195 647 1199
rect 651 1195 652 1199
rect 646 1194 652 1195
rect 702 1199 708 1200
rect 702 1195 703 1199
rect 707 1195 708 1199
rect 702 1194 708 1195
rect 758 1199 764 1200
rect 758 1195 759 1199
rect 763 1195 764 1199
rect 758 1194 764 1195
rect 814 1199 820 1200
rect 814 1195 815 1199
rect 819 1195 820 1199
rect 814 1194 820 1195
rect 870 1199 876 1200
rect 870 1195 871 1199
rect 875 1195 876 1199
rect 870 1194 876 1195
rect 926 1199 932 1200
rect 926 1195 927 1199
rect 931 1195 932 1199
rect 1286 1196 1287 1200
rect 1291 1196 1292 1200
rect 1286 1195 1292 1196
rect 926 1194 932 1195
rect 368 1171 370 1194
rect 424 1171 426 1194
rect 480 1171 482 1194
rect 536 1171 538 1194
rect 592 1171 594 1194
rect 648 1171 650 1194
rect 704 1171 706 1194
rect 760 1171 762 1194
rect 816 1171 818 1194
rect 872 1171 874 1194
rect 928 1171 930 1194
rect 1288 1171 1290 1195
rect 1328 1191 1330 1211
rect 1366 1210 1372 1211
rect 1462 1215 1468 1216
rect 1462 1211 1463 1215
rect 1467 1211 1468 1215
rect 1462 1210 1468 1211
rect 1590 1215 1596 1216
rect 1590 1211 1591 1215
rect 1595 1211 1596 1215
rect 1590 1210 1596 1211
rect 1710 1215 1716 1216
rect 1710 1211 1711 1215
rect 1715 1211 1716 1215
rect 1710 1210 1716 1211
rect 1830 1215 1836 1216
rect 1830 1211 1831 1215
rect 1835 1211 1836 1215
rect 1830 1210 1836 1211
rect 1942 1215 1948 1216
rect 1942 1211 1943 1215
rect 1947 1211 1948 1215
rect 1942 1210 1948 1211
rect 2046 1215 2052 1216
rect 2046 1211 2047 1215
rect 2051 1211 2052 1215
rect 2046 1210 2052 1211
rect 2142 1215 2148 1216
rect 2142 1211 2143 1215
rect 2147 1211 2148 1215
rect 2142 1210 2148 1211
rect 2230 1215 2236 1216
rect 2230 1211 2231 1215
rect 2235 1211 2236 1215
rect 2230 1210 2236 1211
rect 2310 1215 2316 1216
rect 2310 1211 2311 1215
rect 2315 1211 2316 1215
rect 2310 1210 2316 1211
rect 2390 1215 2396 1216
rect 2390 1211 2391 1215
rect 2395 1211 2396 1215
rect 2390 1210 2396 1211
rect 2454 1215 2460 1216
rect 2454 1211 2455 1215
rect 2459 1211 2460 1215
rect 2502 1212 2503 1216
rect 2507 1212 2508 1216
rect 2502 1211 2508 1212
rect 2454 1210 2460 1211
rect 1368 1191 1370 1210
rect 1464 1191 1466 1210
rect 1592 1191 1594 1210
rect 1712 1191 1714 1210
rect 1832 1191 1834 1210
rect 1944 1191 1946 1210
rect 2048 1191 2050 1210
rect 2144 1191 2146 1210
rect 2232 1191 2234 1210
rect 2312 1191 2314 1210
rect 2392 1191 2394 1210
rect 2456 1191 2458 1210
rect 2504 1191 2506 1211
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1463 1190 1467 1191
rect 1463 1185 1467 1186
rect 1471 1190 1475 1191
rect 1471 1185 1475 1186
rect 1591 1190 1595 1191
rect 1591 1185 1595 1186
rect 1599 1190 1603 1191
rect 1599 1185 1603 1186
rect 1711 1190 1715 1191
rect 1711 1185 1715 1186
rect 1735 1190 1739 1191
rect 1735 1185 1739 1186
rect 1831 1190 1835 1191
rect 1831 1185 1835 1186
rect 1863 1190 1867 1191
rect 1863 1185 1867 1186
rect 1943 1190 1947 1191
rect 1943 1185 1947 1186
rect 1983 1190 1987 1191
rect 1983 1185 1987 1186
rect 2047 1190 2051 1191
rect 2047 1185 2051 1186
rect 2087 1190 2091 1191
rect 2087 1185 2091 1186
rect 2143 1190 2147 1191
rect 2143 1185 2147 1186
rect 2191 1190 2195 1191
rect 2191 1185 2195 1186
rect 2231 1190 2235 1191
rect 2231 1185 2235 1186
rect 2287 1190 2291 1191
rect 2287 1185 2291 1186
rect 2311 1190 2315 1191
rect 2311 1185 2315 1186
rect 2383 1190 2387 1191
rect 2383 1185 2387 1186
rect 2391 1190 2395 1191
rect 2391 1185 2395 1186
rect 2455 1190 2459 1191
rect 2455 1185 2459 1186
rect 2503 1190 2507 1191
rect 2503 1185 2507 1186
rect 111 1170 115 1171
rect 111 1165 115 1166
rect 367 1170 371 1171
rect 367 1165 371 1166
rect 423 1170 427 1171
rect 423 1165 427 1166
rect 479 1170 483 1171
rect 479 1165 483 1166
rect 535 1170 539 1171
rect 535 1165 539 1166
rect 591 1170 595 1171
rect 591 1165 595 1166
rect 647 1170 651 1171
rect 647 1165 651 1166
rect 703 1170 707 1171
rect 703 1165 707 1166
rect 759 1170 763 1171
rect 759 1165 763 1166
rect 815 1170 819 1171
rect 815 1165 819 1166
rect 871 1170 875 1171
rect 871 1165 875 1166
rect 927 1170 931 1171
rect 927 1165 931 1166
rect 983 1170 987 1171
rect 983 1165 987 1166
rect 1287 1170 1291 1171
rect 1287 1165 1291 1166
rect 1328 1165 1330 1185
rect 1368 1166 1370 1185
rect 1472 1166 1474 1185
rect 1600 1166 1602 1185
rect 1736 1166 1738 1185
rect 1864 1166 1866 1185
rect 1984 1166 1986 1185
rect 2088 1166 2090 1185
rect 2192 1166 2194 1185
rect 2288 1166 2290 1185
rect 2384 1166 2386 1185
rect 2456 1166 2458 1185
rect 1366 1165 1372 1166
rect 112 1145 114 1165
rect 424 1146 426 1165
rect 480 1146 482 1165
rect 536 1146 538 1165
rect 592 1146 594 1165
rect 648 1146 650 1165
rect 704 1146 706 1165
rect 760 1146 762 1165
rect 816 1146 818 1165
rect 872 1146 874 1165
rect 928 1146 930 1165
rect 984 1146 986 1165
rect 422 1145 428 1146
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 422 1141 423 1145
rect 427 1141 428 1145
rect 422 1140 428 1141
rect 478 1145 484 1146
rect 478 1141 479 1145
rect 483 1141 484 1145
rect 478 1140 484 1141
rect 534 1145 540 1146
rect 534 1141 535 1145
rect 539 1141 540 1145
rect 534 1140 540 1141
rect 590 1145 596 1146
rect 590 1141 591 1145
rect 595 1141 596 1145
rect 590 1140 596 1141
rect 646 1145 652 1146
rect 646 1141 647 1145
rect 651 1141 652 1145
rect 646 1140 652 1141
rect 702 1145 708 1146
rect 702 1141 703 1145
rect 707 1141 708 1145
rect 702 1140 708 1141
rect 758 1145 764 1146
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 814 1145 820 1146
rect 814 1141 815 1145
rect 819 1141 820 1145
rect 814 1140 820 1141
rect 870 1145 876 1146
rect 870 1141 871 1145
rect 875 1141 876 1145
rect 870 1140 876 1141
rect 926 1145 932 1146
rect 926 1141 927 1145
rect 931 1141 932 1145
rect 926 1140 932 1141
rect 982 1145 988 1146
rect 1288 1145 1290 1165
rect 1326 1164 1332 1165
rect 1326 1160 1327 1164
rect 1331 1160 1332 1164
rect 1366 1161 1367 1165
rect 1371 1161 1372 1165
rect 1366 1160 1372 1161
rect 1470 1165 1476 1166
rect 1470 1161 1471 1165
rect 1475 1161 1476 1165
rect 1470 1160 1476 1161
rect 1598 1165 1604 1166
rect 1598 1161 1599 1165
rect 1603 1161 1604 1165
rect 1598 1160 1604 1161
rect 1734 1165 1740 1166
rect 1734 1161 1735 1165
rect 1739 1161 1740 1165
rect 1734 1160 1740 1161
rect 1862 1165 1868 1166
rect 1862 1161 1863 1165
rect 1867 1161 1868 1165
rect 1862 1160 1868 1161
rect 1982 1165 1988 1166
rect 1982 1161 1983 1165
rect 1987 1161 1988 1165
rect 1982 1160 1988 1161
rect 2086 1165 2092 1166
rect 2086 1161 2087 1165
rect 2091 1161 2092 1165
rect 2086 1160 2092 1161
rect 2190 1165 2196 1166
rect 2190 1161 2191 1165
rect 2195 1161 2196 1165
rect 2190 1160 2196 1161
rect 2286 1165 2292 1166
rect 2286 1161 2287 1165
rect 2291 1161 2292 1165
rect 2286 1160 2292 1161
rect 2382 1165 2388 1166
rect 2382 1161 2383 1165
rect 2387 1161 2388 1165
rect 2382 1160 2388 1161
rect 2454 1165 2460 1166
rect 2504 1165 2506 1185
rect 2454 1161 2455 1165
rect 2459 1161 2460 1165
rect 2454 1160 2460 1161
rect 2502 1164 2508 1165
rect 2502 1160 2503 1164
rect 2507 1160 2508 1164
rect 1326 1159 1332 1160
rect 2502 1159 2508 1160
rect 1326 1147 1332 1148
rect 982 1141 983 1145
rect 987 1141 988 1145
rect 982 1140 988 1141
rect 1286 1144 1292 1145
rect 1286 1140 1287 1144
rect 1291 1140 1292 1144
rect 1326 1143 1327 1147
rect 1331 1143 1332 1147
rect 2502 1147 2508 1148
rect 1326 1142 1332 1143
rect 1350 1144 1356 1145
rect 110 1139 116 1140
rect 1286 1139 1292 1140
rect 1328 1135 1330 1142
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1454 1144 1460 1145
rect 1454 1140 1455 1144
rect 1459 1140 1460 1144
rect 1454 1139 1460 1140
rect 1582 1144 1588 1145
rect 1582 1140 1583 1144
rect 1587 1140 1588 1144
rect 1582 1139 1588 1140
rect 1718 1144 1724 1145
rect 1718 1140 1719 1144
rect 1723 1140 1724 1144
rect 1718 1139 1724 1140
rect 1846 1144 1852 1145
rect 1846 1140 1847 1144
rect 1851 1140 1852 1144
rect 1846 1139 1852 1140
rect 1966 1144 1972 1145
rect 1966 1140 1967 1144
rect 1971 1140 1972 1144
rect 1966 1139 1972 1140
rect 2070 1144 2076 1145
rect 2070 1140 2071 1144
rect 2075 1140 2076 1144
rect 2070 1139 2076 1140
rect 2174 1144 2180 1145
rect 2174 1140 2175 1144
rect 2179 1140 2180 1144
rect 2174 1139 2180 1140
rect 2270 1144 2276 1145
rect 2270 1140 2271 1144
rect 2275 1140 2276 1144
rect 2270 1139 2276 1140
rect 2366 1144 2372 1145
rect 2366 1140 2367 1144
rect 2371 1140 2372 1144
rect 2366 1139 2372 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2502 1143 2503 1147
rect 2507 1143 2508 1147
rect 2502 1142 2508 1143
rect 2438 1139 2444 1140
rect 1352 1135 1354 1139
rect 1456 1135 1458 1139
rect 1584 1135 1586 1139
rect 1720 1135 1722 1139
rect 1848 1135 1850 1139
rect 1968 1135 1970 1139
rect 2072 1135 2074 1139
rect 2176 1135 2178 1139
rect 2272 1135 2274 1139
rect 2368 1135 2370 1139
rect 2440 1135 2442 1139
rect 2504 1135 2506 1142
rect 1327 1134 1331 1135
rect 1327 1129 1331 1130
rect 1351 1134 1355 1135
rect 1351 1129 1355 1130
rect 1367 1134 1371 1135
rect 1367 1129 1371 1130
rect 1447 1134 1451 1135
rect 1447 1129 1451 1130
rect 1455 1134 1459 1135
rect 1455 1129 1459 1130
rect 1535 1134 1539 1135
rect 1535 1129 1539 1130
rect 1583 1134 1587 1135
rect 1583 1129 1587 1130
rect 1631 1134 1635 1135
rect 1631 1129 1635 1130
rect 1719 1134 1723 1135
rect 1719 1129 1723 1130
rect 1807 1134 1811 1135
rect 1807 1129 1811 1130
rect 1847 1134 1851 1135
rect 1847 1129 1851 1130
rect 1895 1134 1899 1135
rect 1895 1129 1899 1130
rect 1967 1134 1971 1135
rect 1967 1129 1971 1130
rect 1983 1134 1987 1135
rect 1983 1129 1987 1130
rect 2071 1134 2075 1135
rect 2071 1129 2075 1130
rect 2159 1134 2163 1135
rect 2159 1129 2163 1130
rect 2175 1134 2179 1135
rect 2175 1129 2179 1130
rect 2255 1134 2259 1135
rect 2255 1129 2259 1130
rect 2271 1134 2275 1135
rect 2271 1129 2275 1130
rect 2359 1134 2363 1135
rect 2359 1129 2363 1130
rect 2367 1134 2371 1135
rect 2367 1129 2371 1130
rect 2439 1134 2443 1135
rect 2439 1129 2443 1130
rect 2503 1134 2507 1135
rect 2503 1129 2507 1130
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 1286 1127 1292 1128
rect 110 1122 116 1123
rect 406 1124 412 1125
rect 112 1115 114 1122
rect 406 1120 407 1124
rect 411 1120 412 1124
rect 406 1119 412 1120
rect 462 1124 468 1125
rect 462 1120 463 1124
rect 467 1120 468 1124
rect 462 1119 468 1120
rect 518 1124 524 1125
rect 518 1120 519 1124
rect 523 1120 524 1124
rect 518 1119 524 1120
rect 574 1124 580 1125
rect 574 1120 575 1124
rect 579 1120 580 1124
rect 574 1119 580 1120
rect 630 1124 636 1125
rect 630 1120 631 1124
rect 635 1120 636 1124
rect 630 1119 636 1120
rect 686 1124 692 1125
rect 686 1120 687 1124
rect 691 1120 692 1124
rect 686 1119 692 1120
rect 742 1124 748 1125
rect 742 1120 743 1124
rect 747 1120 748 1124
rect 742 1119 748 1120
rect 798 1124 804 1125
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 798 1119 804 1120
rect 854 1124 860 1125
rect 854 1120 855 1124
rect 859 1120 860 1124
rect 854 1119 860 1120
rect 910 1124 916 1125
rect 910 1120 911 1124
rect 915 1120 916 1124
rect 910 1119 916 1120
rect 966 1124 972 1125
rect 966 1120 967 1124
rect 971 1120 972 1124
rect 1286 1123 1287 1127
rect 1291 1123 1292 1127
rect 1328 1126 1330 1129
rect 1366 1128 1372 1129
rect 1286 1122 1292 1123
rect 1326 1125 1332 1126
rect 966 1119 972 1120
rect 408 1115 410 1119
rect 464 1115 466 1119
rect 520 1115 522 1119
rect 576 1115 578 1119
rect 632 1115 634 1119
rect 688 1115 690 1119
rect 744 1115 746 1119
rect 800 1115 802 1119
rect 856 1115 858 1119
rect 912 1115 914 1119
rect 968 1115 970 1119
rect 1288 1115 1290 1122
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1366 1124 1367 1128
rect 1371 1124 1372 1128
rect 1366 1123 1372 1124
rect 1446 1128 1452 1129
rect 1446 1124 1447 1128
rect 1451 1124 1452 1128
rect 1446 1123 1452 1124
rect 1534 1128 1540 1129
rect 1534 1124 1535 1128
rect 1539 1124 1540 1128
rect 1534 1123 1540 1124
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1806 1128 1812 1129
rect 1806 1124 1807 1128
rect 1811 1124 1812 1128
rect 1806 1123 1812 1124
rect 1894 1128 1900 1129
rect 1894 1124 1895 1128
rect 1899 1124 1900 1128
rect 1894 1123 1900 1124
rect 1982 1128 1988 1129
rect 1982 1124 1983 1128
rect 1987 1124 1988 1128
rect 1982 1123 1988 1124
rect 2070 1128 2076 1129
rect 2070 1124 2071 1128
rect 2075 1124 2076 1128
rect 2070 1123 2076 1124
rect 2158 1128 2164 1129
rect 2158 1124 2159 1128
rect 2163 1124 2164 1128
rect 2158 1123 2164 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 2438 1128 2444 1129
rect 2438 1124 2439 1128
rect 2443 1124 2444 1128
rect 2504 1126 2506 1129
rect 2438 1123 2444 1124
rect 2502 1125 2508 1126
rect 1326 1120 1332 1121
rect 2502 1121 2503 1125
rect 2507 1121 2508 1125
rect 2502 1120 2508 1121
rect 111 1114 115 1115
rect 111 1109 115 1110
rect 223 1114 227 1115
rect 223 1109 227 1110
rect 311 1114 315 1115
rect 311 1109 315 1110
rect 399 1114 403 1115
rect 399 1109 403 1110
rect 407 1114 411 1115
rect 407 1109 411 1110
rect 463 1114 467 1115
rect 463 1109 467 1110
rect 495 1114 499 1115
rect 495 1109 499 1110
rect 519 1114 523 1115
rect 519 1109 523 1110
rect 575 1114 579 1115
rect 575 1109 579 1110
rect 591 1114 595 1115
rect 591 1109 595 1110
rect 631 1114 635 1115
rect 631 1109 635 1110
rect 679 1114 683 1115
rect 679 1109 683 1110
rect 687 1114 691 1115
rect 687 1109 691 1110
rect 743 1114 747 1115
rect 743 1109 747 1110
rect 767 1114 771 1115
rect 767 1109 771 1110
rect 799 1114 803 1115
rect 799 1109 803 1110
rect 847 1114 851 1115
rect 847 1109 851 1110
rect 855 1114 859 1115
rect 855 1109 859 1110
rect 911 1114 915 1115
rect 911 1109 915 1110
rect 927 1114 931 1115
rect 927 1109 931 1110
rect 967 1114 971 1115
rect 967 1109 971 1110
rect 1015 1114 1019 1115
rect 1015 1109 1019 1110
rect 1103 1114 1107 1115
rect 1103 1109 1107 1110
rect 1287 1114 1291 1115
rect 1287 1109 1291 1110
rect 112 1106 114 1109
rect 222 1108 228 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 222 1104 223 1108
rect 227 1104 228 1108
rect 222 1103 228 1104
rect 310 1108 316 1109
rect 310 1104 311 1108
rect 315 1104 316 1108
rect 310 1103 316 1104
rect 398 1108 404 1109
rect 398 1104 399 1108
rect 403 1104 404 1108
rect 398 1103 404 1104
rect 494 1108 500 1109
rect 494 1104 495 1108
rect 499 1104 500 1108
rect 494 1103 500 1104
rect 590 1108 596 1109
rect 590 1104 591 1108
rect 595 1104 596 1108
rect 590 1103 596 1104
rect 678 1108 684 1109
rect 678 1104 679 1108
rect 683 1104 684 1108
rect 678 1103 684 1104
rect 766 1108 772 1109
rect 766 1104 767 1108
rect 771 1104 772 1108
rect 766 1103 772 1104
rect 846 1108 852 1109
rect 846 1104 847 1108
rect 851 1104 852 1108
rect 846 1103 852 1104
rect 926 1108 932 1109
rect 926 1104 927 1108
rect 931 1104 932 1108
rect 926 1103 932 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1102 1108 1108 1109
rect 1102 1104 1103 1108
rect 1107 1104 1108 1108
rect 1288 1106 1290 1109
rect 1326 1108 1332 1109
rect 2502 1108 2508 1109
rect 1102 1103 1108 1104
rect 1286 1105 1292 1106
rect 110 1100 116 1101
rect 1286 1101 1287 1105
rect 1291 1101 1292 1105
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1326 1103 1332 1104
rect 1382 1107 1388 1108
rect 1382 1103 1383 1107
rect 1387 1103 1388 1107
rect 1286 1100 1292 1101
rect 110 1088 116 1089
rect 1286 1088 1292 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 238 1087 244 1088
rect 238 1083 239 1087
rect 243 1083 244 1087
rect 112 1059 114 1083
rect 238 1082 244 1083
rect 326 1087 332 1088
rect 326 1083 327 1087
rect 331 1083 332 1087
rect 326 1082 332 1083
rect 414 1087 420 1088
rect 414 1083 415 1087
rect 419 1083 420 1087
rect 414 1082 420 1083
rect 510 1087 516 1088
rect 510 1083 511 1087
rect 515 1083 516 1087
rect 510 1082 516 1083
rect 606 1087 612 1088
rect 606 1083 607 1087
rect 611 1083 612 1087
rect 606 1082 612 1083
rect 694 1087 700 1088
rect 694 1083 695 1087
rect 699 1083 700 1087
rect 694 1082 700 1083
rect 782 1087 788 1088
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 862 1087 868 1088
rect 862 1083 863 1087
rect 867 1083 868 1087
rect 862 1082 868 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 942 1082 948 1083
rect 1030 1087 1036 1088
rect 1030 1083 1031 1087
rect 1035 1083 1036 1087
rect 1030 1082 1036 1083
rect 1118 1087 1124 1088
rect 1118 1083 1119 1087
rect 1123 1083 1124 1087
rect 1286 1084 1287 1088
rect 1291 1084 1292 1088
rect 1286 1083 1292 1084
rect 1118 1082 1124 1083
rect 240 1059 242 1082
rect 328 1059 330 1082
rect 416 1059 418 1082
rect 512 1059 514 1082
rect 608 1059 610 1082
rect 696 1059 698 1082
rect 784 1059 786 1082
rect 864 1059 866 1082
rect 944 1059 946 1082
rect 1032 1059 1034 1082
rect 1120 1059 1122 1082
rect 1288 1059 1290 1083
rect 1328 1075 1330 1103
rect 1382 1102 1388 1103
rect 1462 1107 1468 1108
rect 1462 1103 1463 1107
rect 1467 1103 1468 1107
rect 1462 1102 1468 1103
rect 1550 1107 1556 1108
rect 1550 1103 1551 1107
rect 1555 1103 1556 1107
rect 1550 1102 1556 1103
rect 1646 1107 1652 1108
rect 1646 1103 1647 1107
rect 1651 1103 1652 1107
rect 1646 1102 1652 1103
rect 1734 1107 1740 1108
rect 1734 1103 1735 1107
rect 1739 1103 1740 1107
rect 1734 1102 1740 1103
rect 1822 1107 1828 1108
rect 1822 1103 1823 1107
rect 1827 1103 1828 1107
rect 1822 1102 1828 1103
rect 1910 1107 1916 1108
rect 1910 1103 1911 1107
rect 1915 1103 1916 1107
rect 1910 1102 1916 1103
rect 1998 1107 2004 1108
rect 1998 1103 1999 1107
rect 2003 1103 2004 1107
rect 1998 1102 2004 1103
rect 2086 1107 2092 1108
rect 2086 1103 2087 1107
rect 2091 1103 2092 1107
rect 2086 1102 2092 1103
rect 2174 1107 2180 1108
rect 2174 1103 2175 1107
rect 2179 1103 2180 1107
rect 2174 1102 2180 1103
rect 2270 1107 2276 1108
rect 2270 1103 2271 1107
rect 2275 1103 2276 1107
rect 2270 1102 2276 1103
rect 2374 1107 2380 1108
rect 2374 1103 2375 1107
rect 2379 1103 2380 1107
rect 2374 1102 2380 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2502 1104 2503 1108
rect 2507 1104 2508 1108
rect 2502 1103 2508 1104
rect 2454 1102 2460 1103
rect 1384 1075 1386 1102
rect 1464 1075 1466 1102
rect 1552 1075 1554 1102
rect 1648 1075 1650 1102
rect 1736 1075 1738 1102
rect 1824 1075 1826 1102
rect 1912 1075 1914 1102
rect 2000 1075 2002 1102
rect 2088 1075 2090 1102
rect 2176 1075 2178 1102
rect 2272 1075 2274 1102
rect 2376 1075 2378 1102
rect 2456 1075 2458 1102
rect 2504 1075 2506 1103
rect 1327 1074 1331 1075
rect 1327 1069 1331 1070
rect 1383 1074 1387 1075
rect 1383 1069 1387 1070
rect 1431 1074 1435 1075
rect 1431 1069 1435 1070
rect 1463 1074 1467 1075
rect 1463 1069 1467 1070
rect 1495 1074 1499 1075
rect 1495 1069 1499 1070
rect 1551 1074 1555 1075
rect 1551 1069 1555 1070
rect 1567 1074 1571 1075
rect 1567 1069 1571 1070
rect 1639 1074 1643 1075
rect 1639 1069 1643 1070
rect 1647 1074 1651 1075
rect 1647 1069 1651 1070
rect 1703 1074 1707 1075
rect 1703 1069 1707 1070
rect 1735 1074 1739 1075
rect 1735 1069 1739 1070
rect 1767 1074 1771 1075
rect 1767 1069 1771 1070
rect 1823 1074 1827 1075
rect 1823 1069 1827 1070
rect 1839 1074 1843 1075
rect 1839 1069 1843 1070
rect 1911 1074 1915 1075
rect 1911 1069 1915 1070
rect 1919 1074 1923 1075
rect 1919 1069 1923 1070
rect 1999 1074 2003 1075
rect 1999 1069 2003 1070
rect 2007 1074 2011 1075
rect 2007 1069 2011 1070
rect 2087 1074 2091 1075
rect 2087 1069 2091 1070
rect 2111 1074 2115 1075
rect 2111 1069 2115 1070
rect 2175 1074 2179 1075
rect 2175 1069 2179 1070
rect 2231 1074 2235 1075
rect 2231 1069 2235 1070
rect 2271 1074 2275 1075
rect 2271 1069 2275 1070
rect 2351 1074 2355 1075
rect 2351 1069 2355 1070
rect 2375 1074 2379 1075
rect 2375 1069 2379 1070
rect 2455 1074 2459 1075
rect 2455 1069 2459 1070
rect 2503 1074 2507 1075
rect 2503 1069 2507 1070
rect 111 1058 115 1059
rect 111 1053 115 1054
rect 151 1058 155 1059
rect 151 1053 155 1054
rect 207 1058 211 1059
rect 207 1053 211 1054
rect 239 1058 243 1059
rect 239 1053 243 1054
rect 303 1058 307 1059
rect 303 1053 307 1054
rect 327 1058 331 1059
rect 327 1053 331 1054
rect 415 1058 419 1059
rect 415 1053 419 1054
rect 511 1058 515 1059
rect 511 1053 515 1054
rect 535 1058 539 1059
rect 535 1053 539 1054
rect 607 1058 611 1059
rect 607 1053 611 1054
rect 655 1058 659 1059
rect 655 1053 659 1054
rect 695 1058 699 1059
rect 695 1053 699 1054
rect 767 1058 771 1059
rect 767 1053 771 1054
rect 783 1058 787 1059
rect 783 1053 787 1054
rect 863 1058 867 1059
rect 863 1053 867 1054
rect 879 1058 883 1059
rect 879 1053 883 1054
rect 943 1058 947 1059
rect 943 1053 947 1054
rect 983 1058 987 1059
rect 983 1053 987 1054
rect 1031 1058 1035 1059
rect 1031 1053 1035 1054
rect 1095 1058 1099 1059
rect 1095 1053 1099 1054
rect 1119 1058 1123 1059
rect 1119 1053 1123 1054
rect 1207 1058 1211 1059
rect 1207 1053 1211 1054
rect 1287 1058 1291 1059
rect 1287 1053 1291 1054
rect 112 1033 114 1053
rect 152 1034 154 1053
rect 208 1034 210 1053
rect 304 1034 306 1053
rect 416 1034 418 1053
rect 536 1034 538 1053
rect 656 1034 658 1053
rect 768 1034 770 1053
rect 880 1034 882 1053
rect 984 1034 986 1053
rect 1096 1034 1098 1053
rect 1208 1034 1210 1053
rect 150 1033 156 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 150 1029 151 1033
rect 155 1029 156 1033
rect 150 1028 156 1029
rect 206 1033 212 1034
rect 206 1029 207 1033
rect 211 1029 212 1033
rect 206 1028 212 1029
rect 302 1033 308 1034
rect 302 1029 303 1033
rect 307 1029 308 1033
rect 302 1028 308 1029
rect 414 1033 420 1034
rect 414 1029 415 1033
rect 419 1029 420 1033
rect 414 1028 420 1029
rect 534 1033 540 1034
rect 534 1029 535 1033
rect 539 1029 540 1033
rect 534 1028 540 1029
rect 654 1033 660 1034
rect 654 1029 655 1033
rect 659 1029 660 1033
rect 654 1028 660 1029
rect 766 1033 772 1034
rect 766 1029 767 1033
rect 771 1029 772 1033
rect 766 1028 772 1029
rect 878 1033 884 1034
rect 878 1029 879 1033
rect 883 1029 884 1033
rect 878 1028 884 1029
rect 982 1033 988 1034
rect 982 1029 983 1033
rect 987 1029 988 1033
rect 982 1028 988 1029
rect 1094 1033 1100 1034
rect 1094 1029 1095 1033
rect 1099 1029 1100 1033
rect 1094 1028 1100 1029
rect 1206 1033 1212 1034
rect 1288 1033 1290 1053
rect 1328 1049 1330 1069
rect 1432 1050 1434 1069
rect 1496 1050 1498 1069
rect 1568 1050 1570 1069
rect 1640 1050 1642 1069
rect 1704 1050 1706 1069
rect 1768 1050 1770 1069
rect 1840 1050 1842 1069
rect 1920 1050 1922 1069
rect 2008 1050 2010 1069
rect 2112 1050 2114 1069
rect 2232 1050 2234 1069
rect 2352 1050 2354 1069
rect 2456 1050 2458 1069
rect 1430 1049 1436 1050
rect 1326 1048 1332 1049
rect 1326 1044 1327 1048
rect 1331 1044 1332 1048
rect 1430 1045 1431 1049
rect 1435 1045 1436 1049
rect 1430 1044 1436 1045
rect 1494 1049 1500 1050
rect 1494 1045 1495 1049
rect 1499 1045 1500 1049
rect 1494 1044 1500 1045
rect 1566 1049 1572 1050
rect 1566 1045 1567 1049
rect 1571 1045 1572 1049
rect 1566 1044 1572 1045
rect 1638 1049 1644 1050
rect 1638 1045 1639 1049
rect 1643 1045 1644 1049
rect 1638 1044 1644 1045
rect 1702 1049 1708 1050
rect 1702 1045 1703 1049
rect 1707 1045 1708 1049
rect 1702 1044 1708 1045
rect 1766 1049 1772 1050
rect 1766 1045 1767 1049
rect 1771 1045 1772 1049
rect 1766 1044 1772 1045
rect 1838 1049 1844 1050
rect 1838 1045 1839 1049
rect 1843 1045 1844 1049
rect 1838 1044 1844 1045
rect 1918 1049 1924 1050
rect 1918 1045 1919 1049
rect 1923 1045 1924 1049
rect 1918 1044 1924 1045
rect 2006 1049 2012 1050
rect 2006 1045 2007 1049
rect 2011 1045 2012 1049
rect 2006 1044 2012 1045
rect 2110 1049 2116 1050
rect 2110 1045 2111 1049
rect 2115 1045 2116 1049
rect 2110 1044 2116 1045
rect 2230 1049 2236 1050
rect 2230 1045 2231 1049
rect 2235 1045 2236 1049
rect 2230 1044 2236 1045
rect 2350 1049 2356 1050
rect 2350 1045 2351 1049
rect 2355 1045 2356 1049
rect 2350 1044 2356 1045
rect 2454 1049 2460 1050
rect 2504 1049 2506 1069
rect 2454 1045 2455 1049
rect 2459 1045 2460 1049
rect 2454 1044 2460 1045
rect 2502 1048 2508 1049
rect 2502 1044 2503 1048
rect 2507 1044 2508 1048
rect 1326 1043 1332 1044
rect 2502 1043 2508 1044
rect 1206 1029 1207 1033
rect 1211 1029 1212 1033
rect 1206 1028 1212 1029
rect 1286 1032 1292 1033
rect 1286 1028 1287 1032
rect 1291 1028 1292 1032
rect 110 1027 116 1028
rect 1286 1027 1292 1028
rect 1326 1031 1332 1032
rect 1326 1027 1327 1031
rect 1331 1027 1332 1031
rect 2502 1031 2508 1032
rect 1326 1026 1332 1027
rect 1414 1028 1420 1029
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 1286 1015 1292 1016
rect 1328 1015 1330 1026
rect 1414 1024 1415 1028
rect 1419 1024 1420 1028
rect 1414 1023 1420 1024
rect 1478 1028 1484 1029
rect 1478 1024 1479 1028
rect 1483 1024 1484 1028
rect 1478 1023 1484 1024
rect 1550 1028 1556 1029
rect 1550 1024 1551 1028
rect 1555 1024 1556 1028
rect 1550 1023 1556 1024
rect 1622 1028 1628 1029
rect 1622 1024 1623 1028
rect 1627 1024 1628 1028
rect 1622 1023 1628 1024
rect 1686 1028 1692 1029
rect 1686 1024 1687 1028
rect 1691 1024 1692 1028
rect 1686 1023 1692 1024
rect 1750 1028 1756 1029
rect 1750 1024 1751 1028
rect 1755 1024 1756 1028
rect 1750 1023 1756 1024
rect 1822 1028 1828 1029
rect 1822 1024 1823 1028
rect 1827 1024 1828 1028
rect 1822 1023 1828 1024
rect 1902 1028 1908 1029
rect 1902 1024 1903 1028
rect 1907 1024 1908 1028
rect 1902 1023 1908 1024
rect 1990 1028 1996 1029
rect 1990 1024 1991 1028
rect 1995 1024 1996 1028
rect 1990 1023 1996 1024
rect 2094 1028 2100 1029
rect 2094 1024 2095 1028
rect 2099 1024 2100 1028
rect 2094 1023 2100 1024
rect 2214 1028 2220 1029
rect 2214 1024 2215 1028
rect 2219 1024 2220 1028
rect 2214 1023 2220 1024
rect 2334 1028 2340 1029
rect 2334 1024 2335 1028
rect 2339 1024 2340 1028
rect 2334 1023 2340 1024
rect 2438 1028 2444 1029
rect 2438 1024 2439 1028
rect 2443 1024 2444 1028
rect 2502 1027 2503 1031
rect 2507 1027 2508 1031
rect 2502 1026 2508 1027
rect 2438 1023 2444 1024
rect 1416 1015 1418 1023
rect 1480 1015 1482 1023
rect 1552 1015 1554 1023
rect 1624 1015 1626 1023
rect 1688 1015 1690 1023
rect 1752 1015 1754 1023
rect 1824 1015 1826 1023
rect 1904 1015 1906 1023
rect 1992 1015 1994 1023
rect 2096 1015 2098 1023
rect 2216 1015 2218 1023
rect 2336 1015 2338 1023
rect 2440 1015 2442 1023
rect 2504 1015 2506 1026
rect 110 1010 116 1011
rect 134 1012 140 1013
rect 112 1003 114 1010
rect 134 1008 135 1012
rect 139 1008 140 1012
rect 134 1007 140 1008
rect 190 1012 196 1013
rect 190 1008 191 1012
rect 195 1008 196 1012
rect 190 1007 196 1008
rect 286 1012 292 1013
rect 286 1008 287 1012
rect 291 1008 292 1012
rect 286 1007 292 1008
rect 398 1012 404 1013
rect 398 1008 399 1012
rect 403 1008 404 1012
rect 398 1007 404 1008
rect 518 1012 524 1013
rect 518 1008 519 1012
rect 523 1008 524 1012
rect 518 1007 524 1008
rect 638 1012 644 1013
rect 638 1008 639 1012
rect 643 1008 644 1012
rect 638 1007 644 1008
rect 750 1012 756 1013
rect 750 1008 751 1012
rect 755 1008 756 1012
rect 750 1007 756 1008
rect 862 1012 868 1013
rect 862 1008 863 1012
rect 867 1008 868 1012
rect 862 1007 868 1008
rect 966 1012 972 1013
rect 966 1008 967 1012
rect 971 1008 972 1012
rect 966 1007 972 1008
rect 1078 1012 1084 1013
rect 1078 1008 1079 1012
rect 1083 1008 1084 1012
rect 1078 1007 1084 1008
rect 1190 1012 1196 1013
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1286 1011 1287 1015
rect 1291 1011 1292 1015
rect 1286 1010 1292 1011
rect 1327 1014 1331 1015
rect 1190 1007 1196 1008
rect 136 1003 138 1007
rect 192 1003 194 1007
rect 288 1003 290 1007
rect 400 1003 402 1007
rect 520 1003 522 1007
rect 640 1003 642 1007
rect 752 1003 754 1007
rect 864 1003 866 1007
rect 968 1003 970 1007
rect 1080 1003 1082 1007
rect 1192 1003 1194 1007
rect 1288 1003 1290 1010
rect 1327 1009 1331 1010
rect 1415 1014 1419 1015
rect 1415 1009 1419 1010
rect 1479 1014 1483 1015
rect 1479 1009 1483 1010
rect 1511 1014 1515 1015
rect 1511 1009 1515 1010
rect 1551 1014 1555 1015
rect 1551 1009 1555 1010
rect 1567 1014 1571 1015
rect 1567 1009 1571 1010
rect 1623 1014 1627 1015
rect 1623 1009 1627 1010
rect 1679 1014 1683 1015
rect 1679 1009 1683 1010
rect 1687 1014 1691 1015
rect 1687 1009 1691 1010
rect 1735 1014 1739 1015
rect 1735 1009 1739 1010
rect 1751 1014 1755 1015
rect 1751 1009 1755 1010
rect 1807 1014 1811 1015
rect 1807 1009 1811 1010
rect 1823 1014 1827 1015
rect 1823 1009 1827 1010
rect 1887 1014 1891 1015
rect 1887 1009 1891 1010
rect 1903 1014 1907 1015
rect 1903 1009 1907 1010
rect 1983 1014 1987 1015
rect 1983 1009 1987 1010
rect 1991 1014 1995 1015
rect 1991 1009 1995 1010
rect 2095 1014 2099 1015
rect 2095 1009 2099 1010
rect 2215 1014 2219 1015
rect 2215 1009 2219 1010
rect 2335 1014 2339 1015
rect 2335 1009 2339 1010
rect 2439 1014 2443 1015
rect 2439 1009 2443 1010
rect 2503 1014 2507 1015
rect 2503 1009 2507 1010
rect 1328 1006 1330 1009
rect 1510 1008 1516 1009
rect 1326 1005 1332 1006
rect 111 1002 115 1003
rect 111 997 115 998
rect 135 1002 139 1003
rect 135 997 139 998
rect 191 1002 195 1003
rect 191 997 195 998
rect 215 1002 219 1003
rect 215 997 219 998
rect 287 1002 291 1003
rect 287 997 291 998
rect 327 1002 331 1003
rect 327 997 331 998
rect 399 1002 403 1003
rect 399 997 403 998
rect 439 1002 443 1003
rect 439 997 443 998
rect 519 1002 523 1003
rect 519 997 523 998
rect 551 1002 555 1003
rect 551 997 555 998
rect 639 1002 643 1003
rect 639 997 643 998
rect 663 1002 667 1003
rect 663 997 667 998
rect 751 1002 755 1003
rect 751 997 755 998
rect 759 1002 763 1003
rect 759 997 763 998
rect 847 1002 851 1003
rect 847 997 851 998
rect 863 1002 867 1003
rect 863 997 867 998
rect 935 1002 939 1003
rect 935 997 939 998
rect 967 1002 971 1003
rect 967 997 971 998
rect 1015 1002 1019 1003
rect 1015 997 1019 998
rect 1079 1002 1083 1003
rect 1079 997 1083 998
rect 1087 1002 1091 1003
rect 1087 997 1091 998
rect 1167 1002 1171 1003
rect 1167 997 1171 998
rect 1191 1002 1195 1003
rect 1191 997 1195 998
rect 1223 1002 1227 1003
rect 1223 997 1227 998
rect 1287 1002 1291 1003
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1566 1008 1572 1009
rect 1566 1004 1567 1008
rect 1571 1004 1572 1008
rect 1566 1003 1572 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1734 1008 1740 1009
rect 1734 1004 1735 1008
rect 1739 1004 1740 1008
rect 1734 1003 1740 1004
rect 1806 1008 1812 1009
rect 1806 1004 1807 1008
rect 1811 1004 1812 1008
rect 1806 1003 1812 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1982 1008 1988 1009
rect 1982 1004 1983 1008
rect 1987 1004 1988 1008
rect 1982 1003 1988 1004
rect 2094 1008 2100 1009
rect 2094 1004 2095 1008
rect 2099 1004 2100 1008
rect 2094 1003 2100 1004
rect 2214 1008 2220 1009
rect 2214 1004 2215 1008
rect 2219 1004 2220 1008
rect 2214 1003 2220 1004
rect 2334 1008 2340 1009
rect 2334 1004 2335 1008
rect 2339 1004 2340 1008
rect 2334 1003 2340 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2504 1006 2506 1009
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 1287 997 1291 998
rect 112 994 114 997
rect 134 996 140 997
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 134 992 135 996
rect 139 992 140 996
rect 134 991 140 992
rect 214 996 220 997
rect 214 992 215 996
rect 219 992 220 996
rect 214 991 220 992
rect 326 996 332 997
rect 326 992 327 996
rect 331 992 332 996
rect 326 991 332 992
rect 438 996 444 997
rect 438 992 439 996
rect 443 992 444 996
rect 438 991 444 992
rect 550 996 556 997
rect 550 992 551 996
rect 555 992 556 996
rect 550 991 556 992
rect 662 996 668 997
rect 662 992 663 996
rect 667 992 668 996
rect 662 991 668 992
rect 758 996 764 997
rect 758 992 759 996
rect 763 992 764 996
rect 758 991 764 992
rect 846 996 852 997
rect 846 992 847 996
rect 851 992 852 996
rect 846 991 852 992
rect 934 996 940 997
rect 934 992 935 996
rect 939 992 940 996
rect 934 991 940 992
rect 1014 996 1020 997
rect 1014 992 1015 996
rect 1019 992 1020 996
rect 1014 991 1020 992
rect 1086 996 1092 997
rect 1086 992 1087 996
rect 1091 992 1092 996
rect 1086 991 1092 992
rect 1166 996 1172 997
rect 1166 992 1167 996
rect 1171 992 1172 996
rect 1166 991 1172 992
rect 1222 996 1228 997
rect 1222 992 1223 996
rect 1227 992 1228 996
rect 1288 994 1290 997
rect 1222 991 1228 992
rect 1286 993 1292 994
rect 110 988 116 989
rect 1286 989 1287 993
rect 1291 989 1292 993
rect 1286 988 1292 989
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 110 976 116 977
rect 1286 976 1292 977
rect 110 972 111 976
rect 115 972 116 976
rect 110 971 116 972
rect 150 975 156 976
rect 150 971 151 975
rect 155 971 156 975
rect 112 951 114 971
rect 150 970 156 971
rect 230 975 236 976
rect 230 971 231 975
rect 235 971 236 975
rect 230 970 236 971
rect 342 975 348 976
rect 342 971 343 975
rect 347 971 348 975
rect 342 970 348 971
rect 454 975 460 976
rect 454 971 455 975
rect 459 971 460 975
rect 454 970 460 971
rect 566 975 572 976
rect 566 971 567 975
rect 571 971 572 975
rect 566 970 572 971
rect 678 975 684 976
rect 678 971 679 975
rect 683 971 684 975
rect 678 970 684 971
rect 774 975 780 976
rect 774 971 775 975
rect 779 971 780 975
rect 774 970 780 971
rect 862 975 868 976
rect 862 971 863 975
rect 867 971 868 975
rect 862 970 868 971
rect 950 975 956 976
rect 950 971 951 975
rect 955 971 956 975
rect 950 970 956 971
rect 1030 975 1036 976
rect 1030 971 1031 975
rect 1035 971 1036 975
rect 1030 970 1036 971
rect 1102 975 1108 976
rect 1102 971 1103 975
rect 1107 971 1108 975
rect 1102 970 1108 971
rect 1182 975 1188 976
rect 1182 971 1183 975
rect 1187 971 1188 975
rect 1182 970 1188 971
rect 1238 975 1244 976
rect 1238 971 1239 975
rect 1243 971 1244 975
rect 1286 972 1287 976
rect 1291 972 1292 976
rect 1286 971 1292 972
rect 1238 970 1244 971
rect 152 951 154 970
rect 232 951 234 970
rect 344 951 346 970
rect 456 951 458 970
rect 568 951 570 970
rect 680 951 682 970
rect 776 951 778 970
rect 864 951 866 970
rect 952 951 954 970
rect 1032 951 1034 970
rect 1104 951 1106 970
rect 1184 951 1186 970
rect 1240 951 1242 970
rect 1288 951 1290 971
rect 111 950 115 951
rect 111 945 115 946
rect 151 950 155 951
rect 151 945 155 946
rect 207 950 211 951
rect 207 945 211 946
rect 231 950 235 951
rect 231 945 235 946
rect 295 950 299 951
rect 295 945 299 946
rect 343 950 347 951
rect 343 945 347 946
rect 399 950 403 951
rect 399 945 403 946
rect 455 950 459 951
rect 455 945 459 946
rect 511 950 515 951
rect 511 945 515 946
rect 567 950 571 951
rect 567 945 571 946
rect 623 950 627 951
rect 623 945 627 946
rect 679 950 683 951
rect 679 945 683 946
rect 735 950 739 951
rect 735 945 739 946
rect 775 950 779 951
rect 775 945 779 946
rect 831 950 835 951
rect 831 945 835 946
rect 863 950 867 951
rect 863 945 867 946
rect 927 950 931 951
rect 927 945 931 946
rect 951 950 955 951
rect 951 945 955 946
rect 1015 950 1019 951
rect 1015 945 1019 946
rect 1031 950 1035 951
rect 1031 945 1035 946
rect 1095 950 1099 951
rect 1095 945 1099 946
rect 1103 950 1107 951
rect 1103 945 1107 946
rect 1175 950 1179 951
rect 1175 945 1179 946
rect 1183 950 1187 951
rect 1183 945 1187 946
rect 1239 950 1243 951
rect 1239 945 1243 946
rect 1287 950 1291 951
rect 1328 947 1330 983
rect 1526 982 1532 983
rect 1582 987 1588 988
rect 1582 983 1583 987
rect 1587 983 1588 987
rect 1582 982 1588 983
rect 1638 987 1644 988
rect 1638 983 1639 987
rect 1643 983 1644 987
rect 1638 982 1644 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1750 987 1756 988
rect 1750 983 1751 987
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1822 987 1828 988
rect 1822 983 1823 987
rect 1827 983 1828 987
rect 1822 982 1828 983
rect 1902 987 1908 988
rect 1902 983 1903 987
rect 1907 983 1908 987
rect 1902 982 1908 983
rect 1998 987 2004 988
rect 1998 983 1999 987
rect 2003 983 2004 987
rect 1998 982 2004 983
rect 2110 987 2116 988
rect 2110 983 2111 987
rect 2115 983 2116 987
rect 2110 982 2116 983
rect 2230 987 2236 988
rect 2230 983 2231 987
rect 2235 983 2236 987
rect 2230 982 2236 983
rect 2350 987 2356 988
rect 2350 983 2351 987
rect 2355 983 2356 987
rect 2350 982 2356 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2454 982 2460 983
rect 1528 947 1530 982
rect 1584 947 1586 982
rect 1640 947 1642 982
rect 1696 947 1698 982
rect 1752 947 1754 982
rect 1824 947 1826 982
rect 1904 947 1906 982
rect 2000 947 2002 982
rect 2112 947 2114 982
rect 2232 947 2234 982
rect 2352 947 2354 982
rect 2456 947 2458 982
rect 2504 947 2506 983
rect 1287 945 1291 946
rect 1327 946 1331 947
rect 112 925 114 945
rect 152 926 154 945
rect 208 926 210 945
rect 296 926 298 945
rect 400 926 402 945
rect 512 926 514 945
rect 624 926 626 945
rect 736 926 738 945
rect 832 926 834 945
rect 928 926 930 945
rect 1016 926 1018 945
rect 1096 926 1098 945
rect 1176 926 1178 945
rect 1240 926 1242 945
rect 150 925 156 926
rect 110 924 116 925
rect 110 920 111 924
rect 115 920 116 924
rect 150 921 151 925
rect 155 921 156 925
rect 150 920 156 921
rect 206 925 212 926
rect 206 921 207 925
rect 211 921 212 925
rect 206 920 212 921
rect 294 925 300 926
rect 294 921 295 925
rect 299 921 300 925
rect 294 920 300 921
rect 398 925 404 926
rect 398 921 399 925
rect 403 921 404 925
rect 398 920 404 921
rect 510 925 516 926
rect 510 921 511 925
rect 515 921 516 925
rect 510 920 516 921
rect 622 925 628 926
rect 622 921 623 925
rect 627 921 628 925
rect 622 920 628 921
rect 734 925 740 926
rect 734 921 735 925
rect 739 921 740 925
rect 734 920 740 921
rect 830 925 836 926
rect 830 921 831 925
rect 835 921 836 925
rect 830 920 836 921
rect 926 925 932 926
rect 926 921 927 925
rect 931 921 932 925
rect 926 920 932 921
rect 1014 925 1020 926
rect 1014 921 1015 925
rect 1019 921 1020 925
rect 1014 920 1020 921
rect 1094 925 1100 926
rect 1094 921 1095 925
rect 1099 921 1100 925
rect 1094 920 1100 921
rect 1174 925 1180 926
rect 1174 921 1175 925
rect 1179 921 1180 925
rect 1174 920 1180 921
rect 1238 925 1244 926
rect 1288 925 1290 945
rect 1327 941 1331 942
rect 1367 946 1371 947
rect 1367 941 1371 942
rect 1439 946 1443 947
rect 1439 941 1443 942
rect 1527 946 1531 947
rect 1527 941 1531 942
rect 1583 946 1587 947
rect 1583 941 1587 942
rect 1615 946 1619 947
rect 1615 941 1619 942
rect 1639 946 1643 947
rect 1639 941 1643 942
rect 1695 946 1699 947
rect 1695 941 1699 942
rect 1751 946 1755 947
rect 1751 941 1755 942
rect 1791 946 1795 947
rect 1791 941 1795 942
rect 1823 946 1827 947
rect 1823 941 1827 942
rect 1895 946 1899 947
rect 1895 941 1899 942
rect 1903 946 1907 947
rect 1903 941 1907 942
rect 1999 946 2003 947
rect 1999 941 2003 942
rect 2015 946 2019 947
rect 2015 941 2019 942
rect 2111 946 2115 947
rect 2111 941 2115 942
rect 2151 946 2155 947
rect 2151 941 2155 942
rect 2231 946 2235 947
rect 2231 941 2235 942
rect 2295 946 2299 947
rect 2295 941 2299 942
rect 2351 946 2355 947
rect 2351 941 2355 942
rect 2439 946 2443 947
rect 2439 941 2443 942
rect 2455 946 2459 947
rect 2455 941 2459 942
rect 2503 946 2507 947
rect 2503 941 2507 942
rect 1238 921 1239 925
rect 1243 921 1244 925
rect 1238 920 1244 921
rect 1286 924 1292 925
rect 1286 920 1287 924
rect 1291 920 1292 924
rect 1328 921 1330 941
rect 1368 922 1370 941
rect 1440 922 1442 941
rect 1528 922 1530 941
rect 1616 922 1618 941
rect 1696 922 1698 941
rect 1792 922 1794 941
rect 1896 922 1898 941
rect 2016 922 2018 941
rect 2152 922 2154 941
rect 2296 922 2298 941
rect 2440 922 2442 941
rect 1366 921 1372 922
rect 110 919 116 920
rect 1286 919 1292 920
rect 1326 920 1332 921
rect 1326 916 1327 920
rect 1331 916 1332 920
rect 1366 917 1367 921
rect 1371 917 1372 921
rect 1366 916 1372 917
rect 1438 921 1444 922
rect 1438 917 1439 921
rect 1443 917 1444 921
rect 1438 916 1444 917
rect 1526 921 1532 922
rect 1526 917 1527 921
rect 1531 917 1532 921
rect 1526 916 1532 917
rect 1614 921 1620 922
rect 1614 917 1615 921
rect 1619 917 1620 921
rect 1614 916 1620 917
rect 1694 921 1700 922
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1790 921 1796 922
rect 1790 917 1791 921
rect 1795 917 1796 921
rect 1790 916 1796 917
rect 1894 921 1900 922
rect 1894 917 1895 921
rect 1899 917 1900 921
rect 1894 916 1900 917
rect 2014 921 2020 922
rect 2014 917 2015 921
rect 2019 917 2020 921
rect 2014 916 2020 917
rect 2150 921 2156 922
rect 2150 917 2151 921
rect 2155 917 2156 921
rect 2150 916 2156 917
rect 2294 921 2300 922
rect 2294 917 2295 921
rect 2299 917 2300 921
rect 2294 916 2300 917
rect 2438 921 2444 922
rect 2504 921 2506 941
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2438 916 2444 917
rect 2502 920 2508 921
rect 2502 916 2503 920
rect 2507 916 2508 920
rect 1326 915 1332 916
rect 2502 915 2508 916
rect 110 907 116 908
rect 110 903 111 907
rect 115 903 116 907
rect 1286 907 1292 908
rect 110 902 116 903
rect 134 904 140 905
rect 112 895 114 902
rect 134 900 135 904
rect 139 900 140 904
rect 134 899 140 900
rect 190 904 196 905
rect 190 900 191 904
rect 195 900 196 904
rect 190 899 196 900
rect 278 904 284 905
rect 278 900 279 904
rect 283 900 284 904
rect 278 899 284 900
rect 382 904 388 905
rect 382 900 383 904
rect 387 900 388 904
rect 382 899 388 900
rect 494 904 500 905
rect 494 900 495 904
rect 499 900 500 904
rect 494 899 500 900
rect 606 904 612 905
rect 606 900 607 904
rect 611 900 612 904
rect 606 899 612 900
rect 718 904 724 905
rect 718 900 719 904
rect 723 900 724 904
rect 718 899 724 900
rect 814 904 820 905
rect 814 900 815 904
rect 819 900 820 904
rect 814 899 820 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 998 904 1004 905
rect 998 900 999 904
rect 1003 900 1004 904
rect 998 899 1004 900
rect 1078 904 1084 905
rect 1078 900 1079 904
rect 1083 900 1084 904
rect 1078 899 1084 900
rect 1158 904 1164 905
rect 1158 900 1159 904
rect 1163 900 1164 904
rect 1158 899 1164 900
rect 1222 904 1228 905
rect 1222 900 1223 904
rect 1227 900 1228 904
rect 1286 903 1287 907
rect 1291 903 1292 907
rect 1286 902 1292 903
rect 1326 903 1332 904
rect 1222 899 1228 900
rect 136 895 138 899
rect 192 895 194 899
rect 280 895 282 899
rect 384 895 386 899
rect 496 895 498 899
rect 608 895 610 899
rect 720 895 722 899
rect 816 895 818 899
rect 912 895 914 899
rect 1000 895 1002 899
rect 1080 895 1082 899
rect 1160 895 1162 899
rect 1224 895 1226 899
rect 1288 895 1290 902
rect 1326 899 1327 903
rect 1331 899 1332 903
rect 2502 903 2508 904
rect 1326 898 1332 899
rect 1350 900 1356 901
rect 111 894 115 895
rect 111 889 115 890
rect 135 894 139 895
rect 135 889 139 890
rect 191 894 195 895
rect 191 889 195 890
rect 247 894 251 895
rect 247 889 251 890
rect 279 894 283 895
rect 279 889 283 890
rect 343 894 347 895
rect 343 889 347 890
rect 383 894 387 895
rect 383 889 387 890
rect 439 894 443 895
rect 439 889 443 890
rect 495 894 499 895
rect 495 889 499 890
rect 543 894 547 895
rect 543 889 547 890
rect 607 894 611 895
rect 607 889 611 890
rect 647 894 651 895
rect 647 889 651 890
rect 719 894 723 895
rect 719 889 723 890
rect 743 894 747 895
rect 743 889 747 890
rect 815 894 819 895
rect 815 889 819 890
rect 839 894 843 895
rect 839 889 843 890
rect 911 894 915 895
rect 911 889 915 890
rect 927 894 931 895
rect 927 889 931 890
rect 999 894 1003 895
rect 999 889 1003 890
rect 1007 894 1011 895
rect 1007 889 1011 890
rect 1079 894 1083 895
rect 1079 889 1083 890
rect 1087 894 1091 895
rect 1087 889 1091 890
rect 1159 894 1163 895
rect 1159 889 1163 890
rect 1167 894 1171 895
rect 1167 889 1171 890
rect 1223 894 1227 895
rect 1223 889 1227 890
rect 1287 894 1291 895
rect 1287 889 1291 890
rect 112 886 114 889
rect 246 888 252 889
rect 110 885 116 886
rect 110 881 111 885
rect 115 881 116 885
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 342 888 348 889
rect 342 884 343 888
rect 347 884 348 888
rect 342 883 348 884
rect 438 888 444 889
rect 438 884 439 888
rect 443 884 444 888
rect 438 883 444 884
rect 542 888 548 889
rect 542 884 543 888
rect 547 884 548 888
rect 542 883 548 884
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 742 888 748 889
rect 742 884 743 888
rect 747 884 748 888
rect 742 883 748 884
rect 838 888 844 889
rect 838 884 839 888
rect 843 884 844 888
rect 838 883 844 884
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 1006 888 1012 889
rect 1006 884 1007 888
rect 1011 884 1012 888
rect 1006 883 1012 884
rect 1086 888 1092 889
rect 1086 884 1087 888
rect 1091 884 1092 888
rect 1086 883 1092 884
rect 1166 888 1172 889
rect 1166 884 1167 888
rect 1171 884 1172 888
rect 1166 883 1172 884
rect 1222 888 1228 889
rect 1222 884 1223 888
rect 1227 884 1228 888
rect 1288 886 1290 889
rect 1328 887 1330 898
rect 1350 896 1351 900
rect 1355 896 1356 900
rect 1350 895 1356 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1510 900 1516 901
rect 1510 896 1511 900
rect 1515 896 1516 900
rect 1510 895 1516 896
rect 1598 900 1604 901
rect 1598 896 1599 900
rect 1603 896 1604 900
rect 1598 895 1604 896
rect 1678 900 1684 901
rect 1678 896 1679 900
rect 1683 896 1684 900
rect 1678 895 1684 896
rect 1774 900 1780 901
rect 1774 896 1775 900
rect 1779 896 1780 900
rect 1774 895 1780 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1998 900 2004 901
rect 1998 896 1999 900
rect 2003 896 2004 900
rect 1998 895 2004 896
rect 2134 900 2140 901
rect 2134 896 2135 900
rect 2139 896 2140 900
rect 2134 895 2140 896
rect 2278 900 2284 901
rect 2278 896 2279 900
rect 2283 896 2284 900
rect 2278 895 2284 896
rect 2422 900 2428 901
rect 2422 896 2423 900
rect 2427 896 2428 900
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2422 895 2428 896
rect 1352 887 1354 895
rect 1424 887 1426 895
rect 1512 887 1514 895
rect 1600 887 1602 895
rect 1680 887 1682 895
rect 1776 887 1778 895
rect 1880 887 1882 895
rect 2000 887 2002 895
rect 2136 887 2138 895
rect 2280 887 2282 895
rect 2424 887 2426 895
rect 2504 887 2506 898
rect 1327 886 1331 887
rect 1222 883 1228 884
rect 1286 885 1292 886
rect 110 880 116 881
rect 1286 881 1287 885
rect 1291 881 1292 885
rect 1327 881 1331 882
rect 1351 886 1355 887
rect 1351 881 1355 882
rect 1423 886 1427 887
rect 1423 881 1427 882
rect 1487 886 1491 887
rect 1487 881 1491 882
rect 1511 886 1515 887
rect 1511 881 1515 882
rect 1559 886 1563 887
rect 1559 881 1563 882
rect 1599 886 1603 887
rect 1599 881 1603 882
rect 1623 886 1627 887
rect 1623 881 1627 882
rect 1679 886 1683 887
rect 1679 881 1683 882
rect 1687 886 1691 887
rect 1687 881 1691 882
rect 1751 886 1755 887
rect 1751 881 1755 882
rect 1775 886 1779 887
rect 1775 881 1779 882
rect 1815 886 1819 887
rect 1815 881 1819 882
rect 1879 886 1883 887
rect 1879 881 1883 882
rect 1887 886 1891 887
rect 1887 881 1891 882
rect 1975 886 1979 887
rect 1975 881 1979 882
rect 1999 886 2003 887
rect 1999 881 2003 882
rect 2079 886 2083 887
rect 2079 881 2083 882
rect 2135 886 2139 887
rect 2135 881 2139 882
rect 2199 886 2203 887
rect 2199 881 2203 882
rect 2279 886 2283 887
rect 2279 881 2283 882
rect 2319 886 2323 887
rect 2319 881 2323 882
rect 2423 886 2427 887
rect 2423 881 2427 882
rect 2439 886 2443 887
rect 2439 881 2443 882
rect 2503 886 2507 887
rect 2503 881 2507 882
rect 1286 880 1292 881
rect 1328 878 1330 881
rect 1486 880 1492 881
rect 1326 877 1332 878
rect 1326 873 1327 877
rect 1331 873 1332 877
rect 1486 876 1487 880
rect 1491 876 1492 880
rect 1486 875 1492 876
rect 1558 880 1564 881
rect 1558 876 1559 880
rect 1563 876 1564 880
rect 1558 875 1564 876
rect 1622 880 1628 881
rect 1622 876 1623 880
rect 1627 876 1628 880
rect 1622 875 1628 876
rect 1686 880 1692 881
rect 1686 876 1687 880
rect 1691 876 1692 880
rect 1686 875 1692 876
rect 1750 880 1756 881
rect 1750 876 1751 880
rect 1755 876 1756 880
rect 1750 875 1756 876
rect 1814 880 1820 881
rect 1814 876 1815 880
rect 1819 876 1820 880
rect 1814 875 1820 876
rect 1886 880 1892 881
rect 1886 876 1887 880
rect 1891 876 1892 880
rect 1886 875 1892 876
rect 1974 880 1980 881
rect 1974 876 1975 880
rect 1979 876 1980 880
rect 1974 875 1980 876
rect 2078 880 2084 881
rect 2078 876 2079 880
rect 2083 876 2084 880
rect 2078 875 2084 876
rect 2198 880 2204 881
rect 2198 876 2199 880
rect 2203 876 2204 880
rect 2198 875 2204 876
rect 2318 880 2324 881
rect 2318 876 2319 880
rect 2323 876 2324 880
rect 2318 875 2324 876
rect 2438 880 2444 881
rect 2438 876 2439 880
rect 2443 876 2444 880
rect 2504 878 2506 881
rect 2438 875 2444 876
rect 2502 877 2508 878
rect 1326 872 1332 873
rect 2502 873 2503 877
rect 2507 873 2508 877
rect 2502 872 2508 873
rect 110 868 116 869
rect 1286 868 1292 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 262 867 268 868
rect 262 863 263 867
rect 267 863 268 867
rect 112 839 114 863
rect 262 862 268 863
rect 358 867 364 868
rect 358 863 359 867
rect 363 863 364 867
rect 358 862 364 863
rect 454 867 460 868
rect 454 863 455 867
rect 459 863 460 867
rect 454 862 460 863
rect 558 867 564 868
rect 558 863 559 867
rect 563 863 564 867
rect 558 862 564 863
rect 662 867 668 868
rect 662 863 663 867
rect 667 863 668 867
rect 662 862 668 863
rect 758 867 764 868
rect 758 863 759 867
rect 763 863 764 867
rect 758 862 764 863
rect 854 867 860 868
rect 854 863 855 867
rect 859 863 860 867
rect 854 862 860 863
rect 942 867 948 868
rect 942 863 943 867
rect 947 863 948 867
rect 942 862 948 863
rect 1022 867 1028 868
rect 1022 863 1023 867
rect 1027 863 1028 867
rect 1022 862 1028 863
rect 1102 867 1108 868
rect 1102 863 1103 867
rect 1107 863 1108 867
rect 1102 862 1108 863
rect 1182 867 1188 868
rect 1182 863 1183 867
rect 1187 863 1188 867
rect 1182 862 1188 863
rect 1238 867 1244 868
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 1286 864 1287 868
rect 1291 864 1292 868
rect 1286 863 1292 864
rect 1238 862 1244 863
rect 264 839 266 862
rect 360 839 362 862
rect 456 839 458 862
rect 560 839 562 862
rect 664 839 666 862
rect 760 839 762 862
rect 856 839 858 862
rect 944 839 946 862
rect 1024 839 1026 862
rect 1104 839 1106 862
rect 1184 839 1186 862
rect 1240 839 1242 862
rect 1288 839 1290 863
rect 1326 860 1332 861
rect 2502 860 2508 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1502 859 1508 860
rect 1502 855 1503 859
rect 1507 855 1508 859
rect 111 838 115 839
rect 111 833 115 834
rect 239 838 243 839
rect 239 833 243 834
rect 263 838 267 839
rect 263 833 267 834
rect 303 838 307 839
rect 303 833 307 834
rect 359 838 363 839
rect 359 833 363 834
rect 383 838 387 839
rect 383 833 387 834
rect 455 838 459 839
rect 455 833 459 834
rect 463 838 467 839
rect 463 833 467 834
rect 551 838 555 839
rect 551 833 555 834
rect 559 838 563 839
rect 559 833 563 834
rect 639 838 643 839
rect 639 833 643 834
rect 663 838 667 839
rect 663 833 667 834
rect 727 838 731 839
rect 727 833 731 834
rect 759 838 763 839
rect 759 833 763 834
rect 807 838 811 839
rect 807 833 811 834
rect 855 838 859 839
rect 855 833 859 834
rect 895 838 899 839
rect 895 833 899 834
rect 943 838 947 839
rect 943 833 947 834
rect 983 838 987 839
rect 983 833 987 834
rect 1023 838 1027 839
rect 1023 833 1027 834
rect 1071 838 1075 839
rect 1071 833 1075 834
rect 1103 838 1107 839
rect 1103 833 1107 834
rect 1183 838 1187 839
rect 1183 833 1187 834
rect 1239 838 1243 839
rect 1239 833 1243 834
rect 1287 838 1291 839
rect 1287 833 1291 834
rect 112 813 114 833
rect 240 814 242 833
rect 304 814 306 833
rect 384 814 386 833
rect 464 814 466 833
rect 552 814 554 833
rect 640 814 642 833
rect 728 814 730 833
rect 808 814 810 833
rect 896 814 898 833
rect 984 814 986 833
rect 1072 814 1074 833
rect 238 813 244 814
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 238 809 239 813
rect 243 809 244 813
rect 238 808 244 809
rect 302 813 308 814
rect 302 809 303 813
rect 307 809 308 813
rect 302 808 308 809
rect 382 813 388 814
rect 382 809 383 813
rect 387 809 388 813
rect 382 808 388 809
rect 462 813 468 814
rect 462 809 463 813
rect 467 809 468 813
rect 462 808 468 809
rect 550 813 556 814
rect 550 809 551 813
rect 555 809 556 813
rect 550 808 556 809
rect 638 813 644 814
rect 638 809 639 813
rect 643 809 644 813
rect 638 808 644 809
rect 726 813 732 814
rect 726 809 727 813
rect 731 809 732 813
rect 726 808 732 809
rect 806 813 812 814
rect 806 809 807 813
rect 811 809 812 813
rect 806 808 812 809
rect 894 813 900 814
rect 894 809 895 813
rect 899 809 900 813
rect 894 808 900 809
rect 982 813 988 814
rect 982 809 983 813
rect 987 809 988 813
rect 982 808 988 809
rect 1070 813 1076 814
rect 1288 813 1290 833
rect 1328 827 1330 855
rect 1502 854 1508 855
rect 1574 859 1580 860
rect 1574 855 1575 859
rect 1579 855 1580 859
rect 1574 854 1580 855
rect 1638 859 1644 860
rect 1638 855 1639 859
rect 1643 855 1644 859
rect 1638 854 1644 855
rect 1702 859 1708 860
rect 1702 855 1703 859
rect 1707 855 1708 859
rect 1702 854 1708 855
rect 1766 859 1772 860
rect 1766 855 1767 859
rect 1771 855 1772 859
rect 1766 854 1772 855
rect 1830 859 1836 860
rect 1830 855 1831 859
rect 1835 855 1836 859
rect 1830 854 1836 855
rect 1902 859 1908 860
rect 1902 855 1903 859
rect 1907 855 1908 859
rect 1902 854 1908 855
rect 1990 859 1996 860
rect 1990 855 1991 859
rect 1995 855 1996 859
rect 1990 854 1996 855
rect 2094 859 2100 860
rect 2094 855 2095 859
rect 2099 855 2100 859
rect 2094 854 2100 855
rect 2214 859 2220 860
rect 2214 855 2215 859
rect 2219 855 2220 859
rect 2214 854 2220 855
rect 2334 859 2340 860
rect 2334 855 2335 859
rect 2339 855 2340 859
rect 2334 854 2340 855
rect 2454 859 2460 860
rect 2454 855 2455 859
rect 2459 855 2460 859
rect 2502 856 2503 860
rect 2507 856 2508 860
rect 2502 855 2508 856
rect 2454 854 2460 855
rect 1504 827 1506 854
rect 1576 827 1578 854
rect 1640 827 1642 854
rect 1704 827 1706 854
rect 1768 827 1770 854
rect 1832 827 1834 854
rect 1904 827 1906 854
rect 1992 827 1994 854
rect 2096 827 2098 854
rect 2216 827 2218 854
rect 2336 827 2338 854
rect 2456 827 2458 854
rect 2504 827 2506 855
rect 1327 826 1331 827
rect 1327 821 1331 822
rect 1439 826 1443 827
rect 1439 821 1443 822
rect 1503 826 1507 827
rect 1503 821 1507 822
rect 1511 826 1515 827
rect 1511 821 1515 822
rect 1575 826 1579 827
rect 1575 821 1579 822
rect 1591 826 1595 827
rect 1591 821 1595 822
rect 1639 826 1643 827
rect 1639 821 1643 822
rect 1671 826 1675 827
rect 1671 821 1675 822
rect 1703 826 1707 827
rect 1703 821 1707 822
rect 1759 826 1763 827
rect 1759 821 1763 822
rect 1767 826 1771 827
rect 1767 821 1771 822
rect 1831 826 1835 827
rect 1831 821 1835 822
rect 1847 826 1851 827
rect 1847 821 1851 822
rect 1903 826 1907 827
rect 1903 821 1907 822
rect 1935 826 1939 827
rect 1935 821 1939 822
rect 1991 826 1995 827
rect 1991 821 1995 822
rect 2023 826 2027 827
rect 2023 821 2027 822
rect 2095 826 2099 827
rect 2095 821 2099 822
rect 2111 826 2115 827
rect 2111 821 2115 822
rect 2199 826 2203 827
rect 2199 821 2203 822
rect 2215 826 2219 827
rect 2215 821 2219 822
rect 2287 826 2291 827
rect 2287 821 2291 822
rect 2335 826 2339 827
rect 2335 821 2339 822
rect 2383 826 2387 827
rect 2383 821 2387 822
rect 2455 826 2459 827
rect 2455 821 2459 822
rect 2503 826 2507 827
rect 2503 821 2507 822
rect 1070 809 1071 813
rect 1075 809 1076 813
rect 1070 808 1076 809
rect 1286 812 1292 813
rect 1286 808 1287 812
rect 1291 808 1292 812
rect 110 807 116 808
rect 1286 807 1292 808
rect 1328 801 1330 821
rect 1440 802 1442 821
rect 1512 802 1514 821
rect 1592 802 1594 821
rect 1672 802 1674 821
rect 1760 802 1762 821
rect 1848 802 1850 821
rect 1936 802 1938 821
rect 2024 802 2026 821
rect 2112 802 2114 821
rect 2200 802 2202 821
rect 2288 802 2290 821
rect 2384 802 2386 821
rect 2456 802 2458 821
rect 1438 801 1444 802
rect 1326 800 1332 801
rect 1326 796 1327 800
rect 1331 796 1332 800
rect 1438 797 1439 801
rect 1443 797 1444 801
rect 1438 796 1444 797
rect 1510 801 1516 802
rect 1510 797 1511 801
rect 1515 797 1516 801
rect 1510 796 1516 797
rect 1590 801 1596 802
rect 1590 797 1591 801
rect 1595 797 1596 801
rect 1590 796 1596 797
rect 1670 801 1676 802
rect 1670 797 1671 801
rect 1675 797 1676 801
rect 1670 796 1676 797
rect 1758 801 1764 802
rect 1758 797 1759 801
rect 1763 797 1764 801
rect 1758 796 1764 797
rect 1846 801 1852 802
rect 1846 797 1847 801
rect 1851 797 1852 801
rect 1846 796 1852 797
rect 1934 801 1940 802
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 2022 801 2028 802
rect 2022 797 2023 801
rect 2027 797 2028 801
rect 2022 796 2028 797
rect 2110 801 2116 802
rect 2110 797 2111 801
rect 2115 797 2116 801
rect 2110 796 2116 797
rect 2198 801 2204 802
rect 2198 797 2199 801
rect 2203 797 2204 801
rect 2198 796 2204 797
rect 2286 801 2292 802
rect 2286 797 2287 801
rect 2291 797 2292 801
rect 2286 796 2292 797
rect 2382 801 2388 802
rect 2382 797 2383 801
rect 2387 797 2388 801
rect 2382 796 2388 797
rect 2454 801 2460 802
rect 2504 801 2506 821
rect 2454 797 2455 801
rect 2459 797 2460 801
rect 2454 796 2460 797
rect 2502 800 2508 801
rect 2502 796 2503 800
rect 2507 796 2508 800
rect 110 795 116 796
rect 110 791 111 795
rect 115 791 116 795
rect 1286 795 1292 796
rect 1326 795 1332 796
rect 2502 795 2508 796
rect 110 790 116 791
rect 222 792 228 793
rect 112 783 114 790
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 286 792 292 793
rect 286 788 287 792
rect 291 788 292 792
rect 286 787 292 788
rect 366 792 372 793
rect 366 788 367 792
rect 371 788 372 792
rect 366 787 372 788
rect 446 792 452 793
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 534 792 540 793
rect 534 788 535 792
rect 539 788 540 792
rect 534 787 540 788
rect 622 792 628 793
rect 622 788 623 792
rect 627 788 628 792
rect 622 787 628 788
rect 710 792 716 793
rect 710 788 711 792
rect 715 788 716 792
rect 710 787 716 788
rect 790 792 796 793
rect 790 788 791 792
rect 795 788 796 792
rect 790 787 796 788
rect 878 792 884 793
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 966 792 972 793
rect 966 788 967 792
rect 971 788 972 792
rect 966 787 972 788
rect 1054 792 1060 793
rect 1054 788 1055 792
rect 1059 788 1060 792
rect 1286 791 1287 795
rect 1291 791 1292 795
rect 1286 790 1292 791
rect 1054 787 1060 788
rect 224 783 226 787
rect 288 783 290 787
rect 368 783 370 787
rect 448 783 450 787
rect 536 783 538 787
rect 624 783 626 787
rect 712 783 714 787
rect 792 783 794 787
rect 880 783 882 787
rect 968 783 970 787
rect 1056 783 1058 787
rect 1288 783 1290 790
rect 1326 783 1332 784
rect 111 782 115 783
rect 111 777 115 778
rect 151 782 155 783
rect 151 777 155 778
rect 223 782 227 783
rect 223 777 227 778
rect 247 782 251 783
rect 247 777 251 778
rect 287 782 291 783
rect 287 777 291 778
rect 343 782 347 783
rect 343 777 347 778
rect 367 782 371 783
rect 367 777 371 778
rect 439 782 443 783
rect 439 777 443 778
rect 447 782 451 783
rect 447 777 451 778
rect 527 782 531 783
rect 527 777 531 778
rect 535 782 539 783
rect 535 777 539 778
rect 607 782 611 783
rect 607 777 611 778
rect 623 782 627 783
rect 623 777 627 778
rect 679 782 683 783
rect 679 777 683 778
rect 711 782 715 783
rect 711 777 715 778
rect 751 782 755 783
rect 751 777 755 778
rect 791 782 795 783
rect 791 777 795 778
rect 823 782 827 783
rect 823 777 827 778
rect 879 782 883 783
rect 879 777 883 778
rect 895 782 899 783
rect 895 777 899 778
rect 967 782 971 783
rect 967 777 971 778
rect 975 782 979 783
rect 975 777 979 778
rect 1055 782 1059 783
rect 1055 777 1059 778
rect 1287 782 1291 783
rect 1326 779 1327 783
rect 1331 779 1332 783
rect 2502 783 2508 784
rect 1326 778 1332 779
rect 1422 780 1428 781
rect 1287 777 1291 778
rect 112 774 114 777
rect 150 776 156 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 150 772 151 776
rect 155 772 156 776
rect 150 771 156 772
rect 246 776 252 777
rect 246 772 247 776
rect 251 772 252 776
rect 246 771 252 772
rect 342 776 348 777
rect 342 772 343 776
rect 347 772 348 776
rect 342 771 348 772
rect 438 776 444 777
rect 438 772 439 776
rect 443 772 444 776
rect 438 771 444 772
rect 526 776 532 777
rect 526 772 527 776
rect 531 772 532 776
rect 526 771 532 772
rect 606 776 612 777
rect 606 772 607 776
rect 611 772 612 776
rect 606 771 612 772
rect 678 776 684 777
rect 678 772 679 776
rect 683 772 684 776
rect 678 771 684 772
rect 750 776 756 777
rect 750 772 751 776
rect 755 772 756 776
rect 750 771 756 772
rect 822 776 828 777
rect 822 772 823 776
rect 827 772 828 776
rect 822 771 828 772
rect 894 776 900 777
rect 894 772 895 776
rect 899 772 900 776
rect 894 771 900 772
rect 974 776 980 777
rect 974 772 975 776
rect 979 772 980 776
rect 1288 774 1290 777
rect 974 771 980 772
rect 1286 773 1292 774
rect 110 768 116 769
rect 1286 769 1287 773
rect 1291 769 1292 773
rect 1328 771 1330 778
rect 1422 776 1423 780
rect 1427 776 1428 780
rect 1422 775 1428 776
rect 1494 780 1500 781
rect 1494 776 1495 780
rect 1499 776 1500 780
rect 1494 775 1500 776
rect 1574 780 1580 781
rect 1574 776 1575 780
rect 1579 776 1580 780
rect 1574 775 1580 776
rect 1654 780 1660 781
rect 1654 776 1655 780
rect 1659 776 1660 780
rect 1654 775 1660 776
rect 1742 780 1748 781
rect 1742 776 1743 780
rect 1747 776 1748 780
rect 1742 775 1748 776
rect 1830 780 1836 781
rect 1830 776 1831 780
rect 1835 776 1836 780
rect 1830 775 1836 776
rect 1918 780 1924 781
rect 1918 776 1919 780
rect 1923 776 1924 780
rect 1918 775 1924 776
rect 2006 780 2012 781
rect 2006 776 2007 780
rect 2011 776 2012 780
rect 2006 775 2012 776
rect 2094 780 2100 781
rect 2094 776 2095 780
rect 2099 776 2100 780
rect 2094 775 2100 776
rect 2182 780 2188 781
rect 2182 776 2183 780
rect 2187 776 2188 780
rect 2182 775 2188 776
rect 2270 780 2276 781
rect 2270 776 2271 780
rect 2275 776 2276 780
rect 2270 775 2276 776
rect 2366 780 2372 781
rect 2366 776 2367 780
rect 2371 776 2372 780
rect 2366 775 2372 776
rect 2438 780 2444 781
rect 2438 776 2439 780
rect 2443 776 2444 780
rect 2502 779 2503 783
rect 2507 779 2508 783
rect 2502 778 2508 779
rect 2438 775 2444 776
rect 1424 771 1426 775
rect 1496 771 1498 775
rect 1576 771 1578 775
rect 1656 771 1658 775
rect 1744 771 1746 775
rect 1832 771 1834 775
rect 1920 771 1922 775
rect 2008 771 2010 775
rect 2096 771 2098 775
rect 2184 771 2186 775
rect 2272 771 2274 775
rect 2368 771 2370 775
rect 2440 771 2442 775
rect 2504 771 2506 778
rect 1286 768 1292 769
rect 1327 770 1331 771
rect 1327 765 1331 766
rect 1351 770 1355 771
rect 1351 765 1355 766
rect 1423 770 1427 771
rect 1423 765 1427 766
rect 1447 770 1451 771
rect 1447 765 1451 766
rect 1495 770 1499 771
rect 1495 765 1499 766
rect 1567 770 1571 771
rect 1567 765 1571 766
rect 1575 770 1579 771
rect 1575 765 1579 766
rect 1655 770 1659 771
rect 1655 765 1659 766
rect 1687 770 1691 771
rect 1687 765 1691 766
rect 1743 770 1747 771
rect 1743 765 1747 766
rect 1807 770 1811 771
rect 1807 765 1811 766
rect 1831 770 1835 771
rect 1831 765 1835 766
rect 1919 770 1923 771
rect 1919 765 1923 766
rect 1927 770 1931 771
rect 1927 765 1931 766
rect 2007 770 2011 771
rect 2007 765 2011 766
rect 2039 770 2043 771
rect 2039 765 2043 766
rect 2095 770 2099 771
rect 2095 765 2099 766
rect 2143 770 2147 771
rect 2143 765 2147 766
rect 2183 770 2187 771
rect 2183 765 2187 766
rect 2247 770 2251 771
rect 2247 765 2251 766
rect 2271 770 2275 771
rect 2271 765 2275 766
rect 2351 770 2355 771
rect 2351 765 2355 766
rect 2367 770 2371 771
rect 2367 765 2371 766
rect 2439 770 2443 771
rect 2439 765 2443 766
rect 2503 770 2507 771
rect 2503 765 2507 766
rect 1328 762 1330 765
rect 1350 764 1356 765
rect 1326 761 1332 762
rect 1326 757 1327 761
rect 1331 757 1332 761
rect 1350 760 1351 764
rect 1355 760 1356 764
rect 1350 759 1356 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1566 764 1572 765
rect 1566 760 1567 764
rect 1571 760 1572 764
rect 1566 759 1572 760
rect 1686 764 1692 765
rect 1686 760 1687 764
rect 1691 760 1692 764
rect 1686 759 1692 760
rect 1806 764 1812 765
rect 1806 760 1807 764
rect 1811 760 1812 764
rect 1806 759 1812 760
rect 1926 764 1932 765
rect 1926 760 1927 764
rect 1931 760 1932 764
rect 1926 759 1932 760
rect 2038 764 2044 765
rect 2038 760 2039 764
rect 2043 760 2044 764
rect 2038 759 2044 760
rect 2142 764 2148 765
rect 2142 760 2143 764
rect 2147 760 2148 764
rect 2142 759 2148 760
rect 2246 764 2252 765
rect 2246 760 2247 764
rect 2251 760 2252 764
rect 2246 759 2252 760
rect 2350 764 2356 765
rect 2350 760 2351 764
rect 2355 760 2356 764
rect 2350 759 2356 760
rect 2438 764 2444 765
rect 2438 760 2439 764
rect 2443 760 2444 764
rect 2504 762 2506 765
rect 2438 759 2444 760
rect 2502 761 2508 762
rect 110 756 116 757
rect 1286 756 1292 757
rect 1326 756 1332 757
rect 2502 757 2503 761
rect 2507 757 2508 761
rect 2502 756 2508 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 112 727 114 751
rect 166 750 172 751
rect 262 755 268 756
rect 262 751 263 755
rect 267 751 268 755
rect 262 750 268 751
rect 358 755 364 756
rect 358 751 359 755
rect 363 751 364 755
rect 358 750 364 751
rect 454 755 460 756
rect 454 751 455 755
rect 459 751 460 755
rect 454 750 460 751
rect 542 755 548 756
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 694 755 700 756
rect 694 751 695 755
rect 699 751 700 755
rect 694 750 700 751
rect 766 755 772 756
rect 766 751 767 755
rect 771 751 772 755
rect 766 750 772 751
rect 838 755 844 756
rect 838 751 839 755
rect 843 751 844 755
rect 838 750 844 751
rect 910 755 916 756
rect 910 751 911 755
rect 915 751 916 755
rect 910 750 916 751
rect 990 755 996 756
rect 990 751 991 755
rect 995 751 996 755
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 990 750 996 751
rect 168 727 170 750
rect 264 727 266 750
rect 360 727 362 750
rect 456 727 458 750
rect 544 727 546 750
rect 624 727 626 750
rect 696 727 698 750
rect 768 727 770 750
rect 840 727 842 750
rect 912 727 914 750
rect 992 727 994 750
rect 1288 727 1290 751
rect 1326 744 1332 745
rect 2502 744 2508 745
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 1326 739 1332 740
rect 1366 743 1372 744
rect 1366 739 1367 743
rect 1371 739 1372 743
rect 111 726 115 727
rect 111 721 115 722
rect 167 726 171 727
rect 167 721 171 722
rect 175 726 179 727
rect 175 721 179 722
rect 263 726 267 727
rect 263 721 267 722
rect 343 726 347 727
rect 343 721 347 722
rect 359 726 363 727
rect 359 721 363 722
rect 423 726 427 727
rect 423 721 427 722
rect 455 726 459 727
rect 455 721 459 722
rect 503 726 507 727
rect 503 721 507 722
rect 543 726 547 727
rect 543 721 547 722
rect 575 726 579 727
rect 575 721 579 722
rect 623 726 627 727
rect 623 721 627 722
rect 639 726 643 727
rect 639 721 643 722
rect 695 726 699 727
rect 695 721 699 722
rect 703 726 707 727
rect 703 721 707 722
rect 767 726 771 727
rect 767 721 771 722
rect 839 726 843 727
rect 839 721 843 722
rect 911 726 915 727
rect 911 721 915 722
rect 991 726 995 727
rect 991 721 995 722
rect 1287 726 1291 727
rect 1287 721 1291 722
rect 112 701 114 721
rect 176 702 178 721
rect 264 702 266 721
rect 344 702 346 721
rect 424 702 426 721
rect 504 702 506 721
rect 576 702 578 721
rect 640 702 642 721
rect 704 702 706 721
rect 768 702 770 721
rect 840 702 842 721
rect 912 702 914 721
rect 174 701 180 702
rect 110 700 116 701
rect 110 696 111 700
rect 115 696 116 700
rect 174 697 175 701
rect 179 697 180 701
rect 174 696 180 697
rect 262 701 268 702
rect 262 697 263 701
rect 267 697 268 701
rect 262 696 268 697
rect 342 701 348 702
rect 342 697 343 701
rect 347 697 348 701
rect 342 696 348 697
rect 422 701 428 702
rect 422 697 423 701
rect 427 697 428 701
rect 422 696 428 697
rect 502 701 508 702
rect 502 697 503 701
rect 507 697 508 701
rect 502 696 508 697
rect 574 701 580 702
rect 574 697 575 701
rect 579 697 580 701
rect 574 696 580 697
rect 638 701 644 702
rect 638 697 639 701
rect 643 697 644 701
rect 638 696 644 697
rect 702 701 708 702
rect 702 697 703 701
rect 707 697 708 701
rect 702 696 708 697
rect 766 701 772 702
rect 766 697 767 701
rect 771 697 772 701
rect 766 696 772 697
rect 838 701 844 702
rect 838 697 839 701
rect 843 697 844 701
rect 838 696 844 697
rect 910 701 916 702
rect 1288 701 1290 721
rect 1328 715 1330 739
rect 1366 738 1372 739
rect 1462 743 1468 744
rect 1462 739 1463 743
rect 1467 739 1468 743
rect 1462 738 1468 739
rect 1582 743 1588 744
rect 1582 739 1583 743
rect 1587 739 1588 743
rect 1582 738 1588 739
rect 1702 743 1708 744
rect 1702 739 1703 743
rect 1707 739 1708 743
rect 1702 738 1708 739
rect 1822 743 1828 744
rect 1822 739 1823 743
rect 1827 739 1828 743
rect 1822 738 1828 739
rect 1942 743 1948 744
rect 1942 739 1943 743
rect 1947 739 1948 743
rect 1942 738 1948 739
rect 2054 743 2060 744
rect 2054 739 2055 743
rect 2059 739 2060 743
rect 2054 738 2060 739
rect 2158 743 2164 744
rect 2158 739 2159 743
rect 2163 739 2164 743
rect 2158 738 2164 739
rect 2262 743 2268 744
rect 2262 739 2263 743
rect 2267 739 2268 743
rect 2262 738 2268 739
rect 2366 743 2372 744
rect 2366 739 2367 743
rect 2371 739 2372 743
rect 2366 738 2372 739
rect 2454 743 2460 744
rect 2454 739 2455 743
rect 2459 739 2460 743
rect 2502 740 2503 744
rect 2507 740 2508 744
rect 2502 739 2508 740
rect 2454 738 2460 739
rect 1368 715 1370 738
rect 1464 715 1466 738
rect 1584 715 1586 738
rect 1704 715 1706 738
rect 1824 715 1826 738
rect 1944 715 1946 738
rect 2056 715 2058 738
rect 2160 715 2162 738
rect 2264 715 2266 738
rect 2368 715 2370 738
rect 2456 715 2458 738
rect 2504 715 2506 739
rect 1327 714 1331 715
rect 1327 709 1331 710
rect 1367 714 1371 715
rect 1367 709 1371 710
rect 1431 714 1435 715
rect 1431 709 1435 710
rect 1463 714 1467 715
rect 1463 709 1467 710
rect 1535 714 1539 715
rect 1535 709 1539 710
rect 1583 714 1587 715
rect 1583 709 1587 710
rect 1639 714 1643 715
rect 1639 709 1643 710
rect 1703 714 1707 715
rect 1703 709 1707 710
rect 1751 714 1755 715
rect 1751 709 1755 710
rect 1823 714 1827 715
rect 1823 709 1827 710
rect 1863 714 1867 715
rect 1863 709 1867 710
rect 1943 714 1947 715
rect 1943 709 1947 710
rect 1967 714 1971 715
rect 1967 709 1971 710
rect 2055 714 2059 715
rect 2055 709 2059 710
rect 2063 714 2067 715
rect 2063 709 2067 710
rect 2151 714 2155 715
rect 2151 709 2155 710
rect 2159 714 2163 715
rect 2159 709 2163 710
rect 2231 714 2235 715
rect 2231 709 2235 710
rect 2263 714 2267 715
rect 2263 709 2267 710
rect 2311 714 2315 715
rect 2311 709 2315 710
rect 2367 714 2371 715
rect 2367 709 2371 710
rect 2391 714 2395 715
rect 2391 709 2395 710
rect 2455 714 2459 715
rect 2455 709 2459 710
rect 2503 714 2507 715
rect 2503 709 2507 710
rect 910 697 911 701
rect 915 697 916 701
rect 910 696 916 697
rect 1286 700 1292 701
rect 1286 696 1287 700
rect 1291 696 1292 700
rect 110 695 116 696
rect 1286 695 1292 696
rect 1328 689 1330 709
rect 1368 690 1370 709
rect 1432 690 1434 709
rect 1536 690 1538 709
rect 1640 690 1642 709
rect 1752 690 1754 709
rect 1864 690 1866 709
rect 1968 690 1970 709
rect 2064 690 2066 709
rect 2152 690 2154 709
rect 2232 690 2234 709
rect 2312 690 2314 709
rect 2392 690 2394 709
rect 2456 690 2458 709
rect 1366 689 1372 690
rect 1326 688 1332 689
rect 1326 684 1327 688
rect 1331 684 1332 688
rect 1366 685 1367 689
rect 1371 685 1372 689
rect 1366 684 1372 685
rect 1430 689 1436 690
rect 1430 685 1431 689
rect 1435 685 1436 689
rect 1430 684 1436 685
rect 1534 689 1540 690
rect 1534 685 1535 689
rect 1539 685 1540 689
rect 1534 684 1540 685
rect 1638 689 1644 690
rect 1638 685 1639 689
rect 1643 685 1644 689
rect 1638 684 1644 685
rect 1750 689 1756 690
rect 1750 685 1751 689
rect 1755 685 1756 689
rect 1750 684 1756 685
rect 1862 689 1868 690
rect 1862 685 1863 689
rect 1867 685 1868 689
rect 1862 684 1868 685
rect 1966 689 1972 690
rect 1966 685 1967 689
rect 1971 685 1972 689
rect 1966 684 1972 685
rect 2062 689 2068 690
rect 2062 685 2063 689
rect 2067 685 2068 689
rect 2062 684 2068 685
rect 2150 689 2156 690
rect 2150 685 2151 689
rect 2155 685 2156 689
rect 2150 684 2156 685
rect 2230 689 2236 690
rect 2230 685 2231 689
rect 2235 685 2236 689
rect 2230 684 2236 685
rect 2310 689 2316 690
rect 2310 685 2311 689
rect 2315 685 2316 689
rect 2310 684 2316 685
rect 2390 689 2396 690
rect 2390 685 2391 689
rect 2395 685 2396 689
rect 2390 684 2396 685
rect 2454 689 2460 690
rect 2504 689 2506 709
rect 2454 685 2455 689
rect 2459 685 2460 689
rect 2454 684 2460 685
rect 2502 688 2508 689
rect 2502 684 2503 688
rect 2507 684 2508 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1286 683 1292 684
rect 1326 683 1332 684
rect 2502 683 2508 684
rect 110 678 116 679
rect 158 680 164 681
rect 112 675 114 678
rect 158 676 159 680
rect 163 676 164 680
rect 158 675 164 676
rect 246 680 252 681
rect 246 676 247 680
rect 251 676 252 680
rect 246 675 252 676
rect 326 680 332 681
rect 326 676 327 680
rect 331 676 332 680
rect 326 675 332 676
rect 406 680 412 681
rect 406 676 407 680
rect 411 676 412 680
rect 406 675 412 676
rect 486 680 492 681
rect 486 676 487 680
rect 491 676 492 680
rect 486 675 492 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 686 680 692 681
rect 686 676 687 680
rect 691 676 692 680
rect 686 675 692 676
rect 750 680 756 681
rect 750 676 751 680
rect 755 676 756 680
rect 750 675 756 676
rect 822 680 828 681
rect 822 676 823 680
rect 827 676 828 680
rect 822 675 828 676
rect 894 680 900 681
rect 894 676 895 680
rect 899 676 900 680
rect 1286 679 1287 683
rect 1291 679 1292 683
rect 1286 678 1292 679
rect 894 675 900 676
rect 1288 675 1290 678
rect 111 674 115 675
rect 111 669 115 670
rect 159 674 163 675
rect 159 669 163 670
rect 215 674 219 675
rect 215 669 219 670
rect 247 674 251 675
rect 247 669 251 670
rect 295 674 299 675
rect 295 669 299 670
rect 327 674 331 675
rect 327 669 331 670
rect 375 674 379 675
rect 375 669 379 670
rect 407 674 411 675
rect 407 669 411 670
rect 455 674 459 675
rect 455 669 459 670
rect 487 674 491 675
rect 487 669 491 670
rect 527 674 531 675
rect 527 669 531 670
rect 559 674 563 675
rect 559 669 563 670
rect 591 674 595 675
rect 591 669 595 670
rect 623 674 627 675
rect 623 669 627 670
rect 655 674 659 675
rect 655 669 659 670
rect 687 674 691 675
rect 687 669 691 670
rect 719 674 723 675
rect 719 669 723 670
rect 751 674 755 675
rect 751 669 755 670
rect 783 674 787 675
rect 783 669 787 670
rect 823 674 827 675
rect 823 669 827 670
rect 847 674 851 675
rect 847 669 851 670
rect 895 674 899 675
rect 895 669 899 670
rect 919 674 923 675
rect 919 669 923 670
rect 1287 674 1291 675
rect 1287 669 1291 670
rect 1326 671 1332 672
rect 112 666 114 669
rect 214 668 220 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 214 664 215 668
rect 219 664 220 668
rect 214 663 220 664
rect 294 668 300 669
rect 294 664 295 668
rect 299 664 300 668
rect 294 663 300 664
rect 374 668 380 669
rect 374 664 375 668
rect 379 664 380 668
rect 374 663 380 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 526 668 532 669
rect 526 664 527 668
rect 531 664 532 668
rect 526 663 532 664
rect 590 668 596 669
rect 590 664 591 668
rect 595 664 596 668
rect 590 663 596 664
rect 654 668 660 669
rect 654 664 655 668
rect 659 664 660 668
rect 654 663 660 664
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 782 668 788 669
rect 782 664 783 668
rect 787 664 788 668
rect 782 663 788 664
rect 846 668 852 669
rect 846 664 847 668
rect 851 664 852 668
rect 846 663 852 664
rect 918 668 924 669
rect 918 664 919 668
rect 923 664 924 668
rect 1288 666 1290 669
rect 1326 667 1327 671
rect 1331 667 1332 671
rect 2502 671 2508 672
rect 1326 666 1332 667
rect 1350 668 1356 669
rect 918 663 924 664
rect 1286 665 1292 666
rect 110 660 116 661
rect 1286 661 1287 665
rect 1291 661 1292 665
rect 1286 660 1292 661
rect 1328 655 1330 666
rect 1350 664 1351 668
rect 1355 664 1356 668
rect 1350 663 1356 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1414 663 1420 664
rect 1518 668 1524 669
rect 1518 664 1519 668
rect 1523 664 1524 668
rect 1518 663 1524 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1734 668 1740 669
rect 1734 664 1735 668
rect 1739 664 1740 668
rect 1734 663 1740 664
rect 1846 668 1852 669
rect 1846 664 1847 668
rect 1851 664 1852 668
rect 1846 663 1852 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2134 668 2140 669
rect 2134 664 2135 668
rect 2139 664 2140 668
rect 2134 663 2140 664
rect 2214 668 2220 669
rect 2214 664 2215 668
rect 2219 664 2220 668
rect 2214 663 2220 664
rect 2294 668 2300 669
rect 2294 664 2295 668
rect 2299 664 2300 668
rect 2294 663 2300 664
rect 2374 668 2380 669
rect 2374 664 2375 668
rect 2379 664 2380 668
rect 2374 663 2380 664
rect 2438 668 2444 669
rect 2438 664 2439 668
rect 2443 664 2444 668
rect 2502 667 2503 671
rect 2507 667 2508 671
rect 2502 666 2508 667
rect 2438 663 2444 664
rect 1352 655 1354 663
rect 1416 655 1418 663
rect 1520 655 1522 663
rect 1624 655 1626 663
rect 1736 655 1738 663
rect 1848 655 1850 663
rect 1952 655 1954 663
rect 2048 655 2050 663
rect 2136 655 2138 663
rect 2216 655 2218 663
rect 2296 655 2298 663
rect 2376 655 2378 663
rect 2440 655 2442 663
rect 2504 655 2506 666
rect 1327 654 1331 655
rect 1327 649 1331 650
rect 1351 654 1355 655
rect 1351 649 1355 650
rect 1415 654 1419 655
rect 1415 649 1419 650
rect 1479 654 1483 655
rect 1479 649 1483 650
rect 1519 654 1523 655
rect 1519 649 1523 650
rect 1559 654 1563 655
rect 1559 649 1563 650
rect 1623 654 1627 655
rect 1623 649 1627 650
rect 1647 654 1651 655
rect 1647 649 1651 650
rect 1735 654 1739 655
rect 1735 649 1739 650
rect 1831 654 1835 655
rect 1831 649 1835 650
rect 1847 654 1851 655
rect 1847 649 1851 650
rect 1919 654 1923 655
rect 1919 649 1923 650
rect 1951 654 1955 655
rect 1951 649 1955 650
rect 2007 654 2011 655
rect 2007 649 2011 650
rect 2047 654 2051 655
rect 2047 649 2051 650
rect 2087 654 2091 655
rect 2087 649 2091 650
rect 2135 654 2139 655
rect 2135 649 2139 650
rect 2167 654 2171 655
rect 2167 649 2171 650
rect 2215 654 2219 655
rect 2215 649 2219 650
rect 2239 654 2243 655
rect 2239 649 2243 650
rect 2295 654 2299 655
rect 2295 649 2299 650
rect 2311 654 2315 655
rect 2311 649 2315 650
rect 2375 654 2379 655
rect 2375 649 2379 650
rect 2383 654 2387 655
rect 2383 649 2387 650
rect 2439 654 2443 655
rect 2439 649 2443 650
rect 2503 654 2507 655
rect 2503 649 2507 650
rect 110 648 116 649
rect 1286 648 1292 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 230 647 236 648
rect 230 643 231 647
rect 235 643 236 647
rect 112 619 114 643
rect 230 642 236 643
rect 310 647 316 648
rect 310 643 311 647
rect 315 643 316 647
rect 310 642 316 643
rect 390 647 396 648
rect 390 643 391 647
rect 395 643 396 647
rect 390 642 396 643
rect 470 647 476 648
rect 470 643 471 647
rect 475 643 476 647
rect 470 642 476 643
rect 542 647 548 648
rect 542 643 543 647
rect 547 643 548 647
rect 542 642 548 643
rect 606 647 612 648
rect 606 643 607 647
rect 611 643 612 647
rect 606 642 612 643
rect 670 647 676 648
rect 670 643 671 647
rect 675 643 676 647
rect 670 642 676 643
rect 734 647 740 648
rect 734 643 735 647
rect 739 643 740 647
rect 734 642 740 643
rect 798 647 804 648
rect 798 643 799 647
rect 803 643 804 647
rect 798 642 804 643
rect 862 647 868 648
rect 862 643 863 647
rect 867 643 868 647
rect 862 642 868 643
rect 934 647 940 648
rect 934 643 935 647
rect 939 643 940 647
rect 1286 644 1287 648
rect 1291 644 1292 648
rect 1328 646 1330 649
rect 1478 648 1484 649
rect 1286 643 1292 644
rect 1326 645 1332 646
rect 934 642 940 643
rect 232 619 234 642
rect 312 619 314 642
rect 392 619 394 642
rect 472 619 474 642
rect 544 619 546 642
rect 608 619 610 642
rect 672 619 674 642
rect 736 619 738 642
rect 800 619 802 642
rect 864 619 866 642
rect 936 619 938 642
rect 1288 619 1290 643
rect 1326 641 1327 645
rect 1331 641 1332 645
rect 1478 644 1479 648
rect 1483 644 1484 648
rect 1478 643 1484 644
rect 1558 648 1564 649
rect 1558 644 1559 648
rect 1563 644 1564 648
rect 1558 643 1564 644
rect 1646 648 1652 649
rect 1646 644 1647 648
rect 1651 644 1652 648
rect 1646 643 1652 644
rect 1734 648 1740 649
rect 1734 644 1735 648
rect 1739 644 1740 648
rect 1734 643 1740 644
rect 1830 648 1836 649
rect 1830 644 1831 648
rect 1835 644 1836 648
rect 1830 643 1836 644
rect 1918 648 1924 649
rect 1918 644 1919 648
rect 1923 644 1924 648
rect 1918 643 1924 644
rect 2006 648 2012 649
rect 2006 644 2007 648
rect 2011 644 2012 648
rect 2006 643 2012 644
rect 2086 648 2092 649
rect 2086 644 2087 648
rect 2091 644 2092 648
rect 2086 643 2092 644
rect 2166 648 2172 649
rect 2166 644 2167 648
rect 2171 644 2172 648
rect 2166 643 2172 644
rect 2238 648 2244 649
rect 2238 644 2239 648
rect 2243 644 2244 648
rect 2238 643 2244 644
rect 2310 648 2316 649
rect 2310 644 2311 648
rect 2315 644 2316 648
rect 2310 643 2316 644
rect 2382 648 2388 649
rect 2382 644 2383 648
rect 2387 644 2388 648
rect 2382 643 2388 644
rect 2438 648 2444 649
rect 2438 644 2439 648
rect 2443 644 2444 648
rect 2504 646 2506 649
rect 2438 643 2444 644
rect 2502 645 2508 646
rect 1326 640 1332 641
rect 2502 641 2503 645
rect 2507 641 2508 645
rect 2502 640 2508 641
rect 1326 628 1332 629
rect 2502 628 2508 629
rect 1326 624 1327 628
rect 1331 624 1332 628
rect 1326 623 1332 624
rect 1494 627 1500 628
rect 1494 623 1495 627
rect 1499 623 1500 627
rect 111 618 115 619
rect 111 613 115 614
rect 207 618 211 619
rect 207 613 211 614
rect 231 618 235 619
rect 231 613 235 614
rect 303 618 307 619
rect 303 613 307 614
rect 311 618 315 619
rect 311 613 315 614
rect 391 618 395 619
rect 391 613 395 614
rect 407 618 411 619
rect 407 613 411 614
rect 471 618 475 619
rect 471 613 475 614
rect 503 618 507 619
rect 503 613 507 614
rect 543 618 547 619
rect 543 613 547 614
rect 599 618 603 619
rect 599 613 603 614
rect 607 618 611 619
rect 607 613 611 614
rect 671 618 675 619
rect 671 613 675 614
rect 687 618 691 619
rect 687 613 691 614
rect 735 618 739 619
rect 735 613 739 614
rect 767 618 771 619
rect 767 613 771 614
rect 799 618 803 619
rect 799 613 803 614
rect 847 618 851 619
rect 847 613 851 614
rect 863 618 867 619
rect 863 613 867 614
rect 927 618 931 619
rect 927 613 931 614
rect 935 618 939 619
rect 935 613 939 614
rect 1007 618 1011 619
rect 1007 613 1011 614
rect 1087 618 1091 619
rect 1087 613 1091 614
rect 1287 618 1291 619
rect 1287 613 1291 614
rect 112 593 114 613
rect 208 594 210 613
rect 304 594 306 613
rect 408 594 410 613
rect 504 594 506 613
rect 600 594 602 613
rect 688 594 690 613
rect 768 594 770 613
rect 848 594 850 613
rect 928 594 930 613
rect 1008 594 1010 613
rect 1088 594 1090 613
rect 206 593 212 594
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 206 589 207 593
rect 211 589 212 593
rect 206 588 212 589
rect 302 593 308 594
rect 302 589 303 593
rect 307 589 308 593
rect 302 588 308 589
rect 406 593 412 594
rect 406 589 407 593
rect 411 589 412 593
rect 406 588 412 589
rect 502 593 508 594
rect 502 589 503 593
rect 507 589 508 593
rect 502 588 508 589
rect 598 593 604 594
rect 598 589 599 593
rect 603 589 604 593
rect 598 588 604 589
rect 686 593 692 594
rect 686 589 687 593
rect 691 589 692 593
rect 686 588 692 589
rect 766 593 772 594
rect 766 589 767 593
rect 771 589 772 593
rect 766 588 772 589
rect 846 593 852 594
rect 846 589 847 593
rect 851 589 852 593
rect 846 588 852 589
rect 926 593 932 594
rect 926 589 927 593
rect 931 589 932 593
rect 926 588 932 589
rect 1006 593 1012 594
rect 1006 589 1007 593
rect 1011 589 1012 593
rect 1006 588 1012 589
rect 1086 593 1092 594
rect 1288 593 1290 613
rect 1328 599 1330 623
rect 1494 622 1500 623
rect 1574 627 1580 628
rect 1574 623 1575 627
rect 1579 623 1580 627
rect 1574 622 1580 623
rect 1662 627 1668 628
rect 1662 623 1663 627
rect 1667 623 1668 627
rect 1662 622 1668 623
rect 1750 627 1756 628
rect 1750 623 1751 627
rect 1755 623 1756 627
rect 1750 622 1756 623
rect 1846 627 1852 628
rect 1846 623 1847 627
rect 1851 623 1852 627
rect 1846 622 1852 623
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 1934 622 1940 623
rect 2022 627 2028 628
rect 2022 623 2023 627
rect 2027 623 2028 627
rect 2022 622 2028 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2182 627 2188 628
rect 2182 623 2183 627
rect 2187 623 2188 627
rect 2182 622 2188 623
rect 2254 627 2260 628
rect 2254 623 2255 627
rect 2259 623 2260 627
rect 2254 622 2260 623
rect 2326 627 2332 628
rect 2326 623 2327 627
rect 2331 623 2332 627
rect 2326 622 2332 623
rect 2398 627 2404 628
rect 2398 623 2399 627
rect 2403 623 2404 627
rect 2398 622 2404 623
rect 2454 627 2460 628
rect 2454 623 2455 627
rect 2459 623 2460 627
rect 2502 624 2503 628
rect 2507 624 2508 628
rect 2502 623 2508 624
rect 2454 622 2460 623
rect 1496 599 1498 622
rect 1576 599 1578 622
rect 1664 599 1666 622
rect 1752 599 1754 622
rect 1848 599 1850 622
rect 1936 599 1938 622
rect 2024 599 2026 622
rect 2104 599 2106 622
rect 2184 599 2186 622
rect 2256 599 2258 622
rect 2328 599 2330 622
rect 2400 599 2402 622
rect 2456 599 2458 622
rect 2504 599 2506 623
rect 1327 598 1331 599
rect 1327 593 1331 594
rect 1455 598 1459 599
rect 1455 593 1459 594
rect 1495 598 1499 599
rect 1495 593 1499 594
rect 1559 598 1563 599
rect 1559 593 1563 594
rect 1575 598 1579 599
rect 1575 593 1579 594
rect 1663 598 1667 599
rect 1663 593 1667 594
rect 1671 598 1675 599
rect 1671 593 1675 594
rect 1751 598 1755 599
rect 1751 593 1755 594
rect 1775 598 1779 599
rect 1775 593 1779 594
rect 1847 598 1851 599
rect 1847 593 1851 594
rect 1879 598 1883 599
rect 1879 593 1883 594
rect 1935 598 1939 599
rect 1935 593 1939 594
rect 1983 598 1987 599
rect 1983 593 1987 594
rect 2023 598 2027 599
rect 2023 593 2027 594
rect 2087 598 2091 599
rect 2087 593 2091 594
rect 2103 598 2107 599
rect 2103 593 2107 594
rect 2183 598 2187 599
rect 2183 593 2187 594
rect 2255 598 2259 599
rect 2255 593 2259 594
rect 2279 598 2283 599
rect 2279 593 2283 594
rect 2327 598 2331 599
rect 2327 593 2331 594
rect 2375 598 2379 599
rect 2375 593 2379 594
rect 2399 598 2403 599
rect 2399 593 2403 594
rect 2455 598 2459 599
rect 2455 593 2459 594
rect 2503 598 2507 599
rect 2503 593 2507 594
rect 1086 589 1087 593
rect 1091 589 1092 593
rect 1086 588 1092 589
rect 1286 592 1292 593
rect 1286 588 1287 592
rect 1291 588 1292 592
rect 110 587 116 588
rect 1286 587 1292 588
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1286 575 1292 576
rect 110 570 116 571
rect 190 572 196 573
rect 112 563 114 570
rect 190 568 191 572
rect 195 568 196 572
rect 190 567 196 568
rect 286 572 292 573
rect 286 568 287 572
rect 291 568 292 572
rect 286 567 292 568
rect 390 572 396 573
rect 390 568 391 572
rect 395 568 396 572
rect 390 567 396 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 670 572 676 573
rect 670 568 671 572
rect 675 568 676 572
rect 670 567 676 568
rect 750 572 756 573
rect 750 568 751 572
rect 755 568 756 572
rect 750 567 756 568
rect 830 572 836 573
rect 830 568 831 572
rect 835 568 836 572
rect 830 567 836 568
rect 910 572 916 573
rect 910 568 911 572
rect 915 568 916 572
rect 910 567 916 568
rect 990 572 996 573
rect 990 568 991 572
rect 995 568 996 572
rect 990 567 996 568
rect 1070 572 1076 573
rect 1070 568 1071 572
rect 1075 568 1076 572
rect 1286 571 1287 575
rect 1291 571 1292 575
rect 1328 573 1330 593
rect 1456 574 1458 593
rect 1560 574 1562 593
rect 1672 574 1674 593
rect 1776 574 1778 593
rect 1880 574 1882 593
rect 1984 574 1986 593
rect 2088 574 2090 593
rect 2184 574 2186 593
rect 2280 574 2282 593
rect 2376 574 2378 593
rect 2456 574 2458 593
rect 1454 573 1460 574
rect 1286 570 1292 571
rect 1326 572 1332 573
rect 1070 567 1076 568
rect 192 563 194 567
rect 288 563 290 567
rect 392 563 394 567
rect 488 563 490 567
rect 584 563 586 567
rect 672 563 674 567
rect 752 563 754 567
rect 832 563 834 567
rect 912 563 914 567
rect 992 563 994 567
rect 1072 563 1074 567
rect 1288 563 1290 570
rect 1326 568 1327 572
rect 1331 568 1332 572
rect 1454 569 1455 573
rect 1459 569 1460 573
rect 1454 568 1460 569
rect 1558 573 1564 574
rect 1558 569 1559 573
rect 1563 569 1564 573
rect 1558 568 1564 569
rect 1670 573 1676 574
rect 1670 569 1671 573
rect 1675 569 1676 573
rect 1670 568 1676 569
rect 1774 573 1780 574
rect 1774 569 1775 573
rect 1779 569 1780 573
rect 1774 568 1780 569
rect 1878 573 1884 574
rect 1878 569 1879 573
rect 1883 569 1884 573
rect 1878 568 1884 569
rect 1982 573 1988 574
rect 1982 569 1983 573
rect 1987 569 1988 573
rect 1982 568 1988 569
rect 2086 573 2092 574
rect 2086 569 2087 573
rect 2091 569 2092 573
rect 2086 568 2092 569
rect 2182 573 2188 574
rect 2182 569 2183 573
rect 2187 569 2188 573
rect 2182 568 2188 569
rect 2278 573 2284 574
rect 2278 569 2279 573
rect 2283 569 2284 573
rect 2278 568 2284 569
rect 2374 573 2380 574
rect 2374 569 2375 573
rect 2379 569 2380 573
rect 2374 568 2380 569
rect 2454 573 2460 574
rect 2504 573 2506 593
rect 2454 569 2455 573
rect 2459 569 2460 573
rect 2454 568 2460 569
rect 2502 572 2508 573
rect 2502 568 2503 572
rect 2507 568 2508 572
rect 1326 567 1332 568
rect 2502 567 2508 568
rect 111 562 115 563
rect 111 557 115 558
rect 175 562 179 563
rect 175 557 179 558
rect 191 562 195 563
rect 191 557 195 558
rect 271 562 275 563
rect 271 557 275 558
rect 287 562 291 563
rect 287 557 291 558
rect 375 562 379 563
rect 375 557 379 558
rect 391 562 395 563
rect 391 557 395 558
rect 487 562 491 563
rect 487 557 491 558
rect 583 562 587 563
rect 583 557 587 558
rect 591 562 595 563
rect 591 557 595 558
rect 671 562 675 563
rect 671 557 675 558
rect 695 562 699 563
rect 695 557 699 558
rect 751 562 755 563
rect 751 557 755 558
rect 791 562 795 563
rect 791 557 795 558
rect 831 562 835 563
rect 831 557 835 558
rect 879 562 883 563
rect 879 557 883 558
rect 911 562 915 563
rect 911 557 915 558
rect 967 562 971 563
rect 967 557 971 558
rect 991 562 995 563
rect 991 557 995 558
rect 1055 562 1059 563
rect 1055 557 1059 558
rect 1071 562 1075 563
rect 1071 557 1075 558
rect 1151 562 1155 563
rect 1151 557 1155 558
rect 1287 562 1291 563
rect 1287 557 1291 558
rect 112 554 114 557
rect 174 556 180 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 270 556 276 557
rect 270 552 271 556
rect 275 552 276 556
rect 270 551 276 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 486 556 492 557
rect 486 552 487 556
rect 491 552 492 556
rect 486 551 492 552
rect 590 556 596 557
rect 590 552 591 556
rect 595 552 596 556
rect 590 551 596 552
rect 694 556 700 557
rect 694 552 695 556
rect 699 552 700 556
rect 694 551 700 552
rect 790 556 796 557
rect 790 552 791 556
rect 795 552 796 556
rect 790 551 796 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 966 556 972 557
rect 966 552 967 556
rect 971 552 972 556
rect 966 551 972 552
rect 1054 556 1060 557
rect 1054 552 1055 556
rect 1059 552 1060 556
rect 1054 551 1060 552
rect 1150 556 1156 557
rect 1150 552 1151 556
rect 1155 552 1156 556
rect 1288 554 1290 557
rect 1326 555 1332 556
rect 1150 551 1156 552
rect 1286 553 1292 554
rect 110 548 116 549
rect 1286 549 1287 553
rect 1291 549 1292 553
rect 1326 551 1327 555
rect 1331 551 1332 555
rect 2502 555 2508 556
rect 1326 550 1332 551
rect 1438 552 1444 553
rect 1286 548 1292 549
rect 1328 543 1330 550
rect 1438 548 1439 552
rect 1443 548 1444 552
rect 1438 547 1444 548
rect 1542 552 1548 553
rect 1542 548 1543 552
rect 1547 548 1548 552
rect 1542 547 1548 548
rect 1654 552 1660 553
rect 1654 548 1655 552
rect 1659 548 1660 552
rect 1654 547 1660 548
rect 1758 552 1764 553
rect 1758 548 1759 552
rect 1763 548 1764 552
rect 1758 547 1764 548
rect 1862 552 1868 553
rect 1862 548 1863 552
rect 1867 548 1868 552
rect 1862 547 1868 548
rect 1966 552 1972 553
rect 1966 548 1967 552
rect 1971 548 1972 552
rect 1966 547 1972 548
rect 2070 552 2076 553
rect 2070 548 2071 552
rect 2075 548 2076 552
rect 2070 547 2076 548
rect 2166 552 2172 553
rect 2166 548 2167 552
rect 2171 548 2172 552
rect 2166 547 2172 548
rect 2262 552 2268 553
rect 2262 548 2263 552
rect 2267 548 2268 552
rect 2262 547 2268 548
rect 2358 552 2364 553
rect 2358 548 2359 552
rect 2363 548 2364 552
rect 2358 547 2364 548
rect 2438 552 2444 553
rect 2438 548 2439 552
rect 2443 548 2444 552
rect 2502 551 2503 555
rect 2507 551 2508 555
rect 2502 550 2508 551
rect 2438 547 2444 548
rect 1440 543 1442 547
rect 1544 543 1546 547
rect 1656 543 1658 547
rect 1760 543 1762 547
rect 1864 543 1866 547
rect 1968 543 1970 547
rect 2072 543 2074 547
rect 2168 543 2170 547
rect 2264 543 2266 547
rect 2360 543 2362 547
rect 2440 543 2442 547
rect 2504 543 2506 550
rect 1327 542 1331 543
rect 1327 537 1331 538
rect 1367 542 1371 543
rect 1367 537 1371 538
rect 1439 542 1443 543
rect 1439 537 1443 538
rect 1447 542 1451 543
rect 1447 537 1451 538
rect 1527 542 1531 543
rect 1527 537 1531 538
rect 1543 542 1547 543
rect 1543 537 1547 538
rect 1615 542 1619 543
rect 1615 537 1619 538
rect 1655 542 1659 543
rect 1655 537 1659 538
rect 1711 542 1715 543
rect 1711 537 1715 538
rect 1759 542 1763 543
rect 1759 537 1763 538
rect 1799 542 1803 543
rect 1799 537 1803 538
rect 1863 542 1867 543
rect 1863 537 1867 538
rect 1887 542 1891 543
rect 1887 537 1891 538
rect 1967 542 1971 543
rect 1967 537 1971 538
rect 1975 542 1979 543
rect 1975 537 1979 538
rect 2063 542 2067 543
rect 2063 537 2067 538
rect 2071 542 2075 543
rect 2071 537 2075 538
rect 2151 542 2155 543
rect 2151 537 2155 538
rect 2167 542 2171 543
rect 2167 537 2171 538
rect 2247 542 2251 543
rect 2247 537 2251 538
rect 2263 542 2267 543
rect 2263 537 2267 538
rect 2343 542 2347 543
rect 2343 537 2347 538
rect 2359 542 2363 543
rect 2359 537 2363 538
rect 2439 542 2443 543
rect 2439 537 2443 538
rect 2503 542 2507 543
rect 2503 537 2507 538
rect 110 536 116 537
rect 1286 536 1292 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 190 535 196 536
rect 190 531 191 535
rect 195 531 196 535
rect 112 507 114 531
rect 190 530 196 531
rect 286 535 292 536
rect 286 531 287 535
rect 291 531 292 535
rect 286 530 292 531
rect 390 535 396 536
rect 390 531 391 535
rect 395 531 396 535
rect 390 530 396 531
rect 502 535 508 536
rect 502 531 503 535
rect 507 531 508 535
rect 502 530 508 531
rect 606 535 612 536
rect 606 531 607 535
rect 611 531 612 535
rect 606 530 612 531
rect 710 535 716 536
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 806 535 812 536
rect 806 531 807 535
rect 811 531 812 535
rect 806 530 812 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 982 535 988 536
rect 982 531 983 535
rect 987 531 988 535
rect 982 530 988 531
rect 1070 535 1076 536
rect 1070 531 1071 535
rect 1075 531 1076 535
rect 1070 530 1076 531
rect 1166 535 1172 536
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1286 532 1287 536
rect 1291 532 1292 536
rect 1328 534 1330 537
rect 1366 536 1372 537
rect 1286 531 1292 532
rect 1326 533 1332 534
rect 1166 530 1172 531
rect 192 507 194 530
rect 288 507 290 530
rect 392 507 394 530
rect 504 507 506 530
rect 608 507 610 530
rect 712 507 714 530
rect 808 507 810 530
rect 896 507 898 530
rect 984 507 986 530
rect 1072 507 1074 530
rect 1168 507 1170 530
rect 1288 507 1290 531
rect 1326 529 1327 533
rect 1331 529 1332 533
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1446 536 1452 537
rect 1446 532 1447 536
rect 1451 532 1452 536
rect 1446 531 1452 532
rect 1526 536 1532 537
rect 1526 532 1527 536
rect 1531 532 1532 536
rect 1526 531 1532 532
rect 1614 536 1620 537
rect 1614 532 1615 536
rect 1619 532 1620 536
rect 1614 531 1620 532
rect 1710 536 1716 537
rect 1710 532 1711 536
rect 1715 532 1716 536
rect 1710 531 1716 532
rect 1798 536 1804 537
rect 1798 532 1799 536
rect 1803 532 1804 536
rect 1798 531 1804 532
rect 1886 536 1892 537
rect 1886 532 1887 536
rect 1891 532 1892 536
rect 1886 531 1892 532
rect 1974 536 1980 537
rect 1974 532 1975 536
rect 1979 532 1980 536
rect 1974 531 1980 532
rect 2062 536 2068 537
rect 2062 532 2063 536
rect 2067 532 2068 536
rect 2062 531 2068 532
rect 2150 536 2156 537
rect 2150 532 2151 536
rect 2155 532 2156 536
rect 2150 531 2156 532
rect 2246 536 2252 537
rect 2246 532 2247 536
rect 2251 532 2252 536
rect 2246 531 2252 532
rect 2342 536 2348 537
rect 2342 532 2343 536
rect 2347 532 2348 536
rect 2342 531 2348 532
rect 2438 536 2444 537
rect 2438 532 2439 536
rect 2443 532 2444 536
rect 2504 534 2506 537
rect 2438 531 2444 532
rect 2502 533 2508 534
rect 1326 528 1332 529
rect 2502 529 2503 533
rect 2507 529 2508 533
rect 2502 528 2508 529
rect 1326 516 1332 517
rect 2502 516 2508 517
rect 1326 512 1327 516
rect 1331 512 1332 516
rect 1326 511 1332 512
rect 1382 515 1388 516
rect 1382 511 1383 515
rect 1387 511 1388 515
rect 111 506 115 507
rect 111 501 115 502
rect 151 506 155 507
rect 151 501 155 502
rect 191 506 195 507
rect 191 501 195 502
rect 247 506 251 507
rect 247 501 251 502
rect 287 506 291 507
rect 287 501 291 502
rect 367 506 371 507
rect 367 501 371 502
rect 391 506 395 507
rect 391 501 395 502
rect 487 506 491 507
rect 487 501 491 502
rect 503 506 507 507
rect 503 501 507 502
rect 607 506 611 507
rect 607 501 611 502
rect 615 506 619 507
rect 615 501 619 502
rect 711 506 715 507
rect 711 501 715 502
rect 735 506 739 507
rect 735 501 739 502
rect 807 506 811 507
rect 807 501 811 502
rect 847 506 851 507
rect 847 501 851 502
rect 895 506 899 507
rect 895 501 899 502
rect 951 506 955 507
rect 951 501 955 502
rect 983 506 987 507
rect 983 501 987 502
rect 1055 506 1059 507
rect 1055 501 1059 502
rect 1071 506 1075 507
rect 1071 501 1075 502
rect 1159 506 1163 507
rect 1159 501 1163 502
rect 1167 506 1171 507
rect 1167 501 1171 502
rect 1239 506 1243 507
rect 1239 501 1243 502
rect 1287 506 1291 507
rect 1287 501 1291 502
rect 112 481 114 501
rect 152 482 154 501
rect 248 482 250 501
rect 368 482 370 501
rect 488 482 490 501
rect 616 482 618 501
rect 736 482 738 501
rect 848 482 850 501
rect 952 482 954 501
rect 1056 482 1058 501
rect 1160 482 1162 501
rect 1240 482 1242 501
rect 150 481 156 482
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 150 477 151 481
rect 155 477 156 481
rect 150 476 156 477
rect 246 481 252 482
rect 246 477 247 481
rect 251 477 252 481
rect 246 476 252 477
rect 366 481 372 482
rect 366 477 367 481
rect 371 477 372 481
rect 366 476 372 477
rect 486 481 492 482
rect 486 477 487 481
rect 491 477 492 481
rect 486 476 492 477
rect 614 481 620 482
rect 614 477 615 481
rect 619 477 620 481
rect 614 476 620 477
rect 734 481 740 482
rect 734 477 735 481
rect 739 477 740 481
rect 734 476 740 477
rect 846 481 852 482
rect 846 477 847 481
rect 851 477 852 481
rect 846 476 852 477
rect 950 481 956 482
rect 950 477 951 481
rect 955 477 956 481
rect 950 476 956 477
rect 1054 481 1060 482
rect 1054 477 1055 481
rect 1059 477 1060 481
rect 1054 476 1060 477
rect 1158 481 1164 482
rect 1158 477 1159 481
rect 1163 477 1164 481
rect 1158 476 1164 477
rect 1238 481 1244 482
rect 1288 481 1290 501
rect 1328 487 1330 511
rect 1382 510 1388 511
rect 1462 515 1468 516
rect 1462 511 1463 515
rect 1467 511 1468 515
rect 1462 510 1468 511
rect 1542 515 1548 516
rect 1542 511 1543 515
rect 1547 511 1548 515
rect 1542 510 1548 511
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 1726 515 1732 516
rect 1726 511 1727 515
rect 1731 511 1732 515
rect 1726 510 1732 511
rect 1814 515 1820 516
rect 1814 511 1815 515
rect 1819 511 1820 515
rect 1814 510 1820 511
rect 1902 515 1908 516
rect 1902 511 1903 515
rect 1907 511 1908 515
rect 1902 510 1908 511
rect 1990 515 1996 516
rect 1990 511 1991 515
rect 1995 511 1996 515
rect 1990 510 1996 511
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2166 515 2172 516
rect 2166 511 2167 515
rect 2171 511 2172 515
rect 2166 510 2172 511
rect 2262 515 2268 516
rect 2262 511 2263 515
rect 2267 511 2268 515
rect 2262 510 2268 511
rect 2358 515 2364 516
rect 2358 511 2359 515
rect 2363 511 2364 515
rect 2358 510 2364 511
rect 2454 515 2460 516
rect 2454 511 2455 515
rect 2459 511 2460 515
rect 2502 512 2503 516
rect 2507 512 2508 516
rect 2502 511 2508 512
rect 2454 510 2460 511
rect 1384 487 1386 510
rect 1464 487 1466 510
rect 1544 487 1546 510
rect 1632 487 1634 510
rect 1728 487 1730 510
rect 1816 487 1818 510
rect 1904 487 1906 510
rect 1992 487 1994 510
rect 2080 487 2082 510
rect 2168 487 2170 510
rect 2264 487 2266 510
rect 2360 487 2362 510
rect 2456 487 2458 510
rect 2504 487 2506 511
rect 1327 486 1331 487
rect 1327 481 1331 482
rect 1367 486 1371 487
rect 1367 481 1371 482
rect 1383 486 1387 487
rect 1383 481 1387 482
rect 1431 486 1435 487
rect 1431 481 1435 482
rect 1463 486 1467 487
rect 1463 481 1467 482
rect 1519 486 1523 487
rect 1519 481 1523 482
rect 1543 486 1547 487
rect 1543 481 1547 482
rect 1615 486 1619 487
rect 1615 481 1619 482
rect 1631 486 1635 487
rect 1631 481 1635 482
rect 1711 486 1715 487
rect 1711 481 1715 482
rect 1727 486 1731 487
rect 1727 481 1731 482
rect 1815 486 1819 487
rect 1815 481 1819 482
rect 1903 486 1907 487
rect 1903 481 1907 482
rect 1927 486 1931 487
rect 1927 481 1931 482
rect 1991 486 1995 487
rect 1991 481 1995 482
rect 2055 486 2059 487
rect 2055 481 2059 482
rect 2079 486 2083 487
rect 2079 481 2083 482
rect 2167 486 2171 487
rect 2167 481 2171 482
rect 2191 486 2195 487
rect 2191 481 2195 482
rect 2263 486 2267 487
rect 2263 481 2267 482
rect 2335 486 2339 487
rect 2335 481 2339 482
rect 2359 486 2363 487
rect 2359 481 2363 482
rect 2455 486 2459 487
rect 2455 481 2459 482
rect 2503 486 2507 487
rect 2503 481 2507 482
rect 1238 477 1239 481
rect 1243 477 1244 481
rect 1238 476 1244 477
rect 1286 480 1292 481
rect 1286 476 1287 480
rect 1291 476 1292 480
rect 110 475 116 476
rect 1286 475 1292 476
rect 110 463 116 464
rect 110 459 111 463
rect 115 459 116 463
rect 1286 463 1292 464
rect 110 458 116 459
rect 134 460 140 461
rect 112 451 114 458
rect 134 456 135 460
rect 139 456 140 460
rect 134 455 140 456
rect 230 460 236 461
rect 230 456 231 460
rect 235 456 236 460
rect 230 455 236 456
rect 350 460 356 461
rect 350 456 351 460
rect 355 456 356 460
rect 350 455 356 456
rect 470 460 476 461
rect 470 456 471 460
rect 475 456 476 460
rect 470 455 476 456
rect 598 460 604 461
rect 598 456 599 460
rect 603 456 604 460
rect 598 455 604 456
rect 718 460 724 461
rect 718 456 719 460
rect 723 456 724 460
rect 718 455 724 456
rect 830 460 836 461
rect 830 456 831 460
rect 835 456 836 460
rect 830 455 836 456
rect 934 460 940 461
rect 934 456 935 460
rect 939 456 940 460
rect 934 455 940 456
rect 1038 460 1044 461
rect 1038 456 1039 460
rect 1043 456 1044 460
rect 1038 455 1044 456
rect 1142 460 1148 461
rect 1142 456 1143 460
rect 1147 456 1148 460
rect 1142 455 1148 456
rect 1222 460 1228 461
rect 1222 456 1223 460
rect 1227 456 1228 460
rect 1286 459 1287 463
rect 1291 459 1292 463
rect 1328 461 1330 481
rect 1368 462 1370 481
rect 1432 462 1434 481
rect 1520 462 1522 481
rect 1616 462 1618 481
rect 1712 462 1714 481
rect 1816 462 1818 481
rect 1928 462 1930 481
rect 2056 462 2058 481
rect 2192 462 2194 481
rect 2336 462 2338 481
rect 2456 462 2458 481
rect 1366 461 1372 462
rect 1286 458 1292 459
rect 1326 460 1332 461
rect 1222 455 1228 456
rect 136 451 138 455
rect 232 451 234 455
rect 352 451 354 455
rect 472 451 474 455
rect 600 451 602 455
rect 720 451 722 455
rect 832 451 834 455
rect 936 451 938 455
rect 1040 451 1042 455
rect 1144 451 1146 455
rect 1224 451 1226 455
rect 1288 451 1290 458
rect 1326 456 1327 460
rect 1331 456 1332 460
rect 1366 457 1367 461
rect 1371 457 1372 461
rect 1366 456 1372 457
rect 1430 461 1436 462
rect 1430 457 1431 461
rect 1435 457 1436 461
rect 1430 456 1436 457
rect 1518 461 1524 462
rect 1518 457 1519 461
rect 1523 457 1524 461
rect 1518 456 1524 457
rect 1614 461 1620 462
rect 1614 457 1615 461
rect 1619 457 1620 461
rect 1614 456 1620 457
rect 1710 461 1716 462
rect 1710 457 1711 461
rect 1715 457 1716 461
rect 1710 456 1716 457
rect 1814 461 1820 462
rect 1814 457 1815 461
rect 1819 457 1820 461
rect 1814 456 1820 457
rect 1926 461 1932 462
rect 1926 457 1927 461
rect 1931 457 1932 461
rect 1926 456 1932 457
rect 2054 461 2060 462
rect 2054 457 2055 461
rect 2059 457 2060 461
rect 2054 456 2060 457
rect 2190 461 2196 462
rect 2190 457 2191 461
rect 2195 457 2196 461
rect 2190 456 2196 457
rect 2334 461 2340 462
rect 2334 457 2335 461
rect 2339 457 2340 461
rect 2334 456 2340 457
rect 2454 461 2460 462
rect 2504 461 2506 481
rect 2454 457 2455 461
rect 2459 457 2460 461
rect 2454 456 2460 457
rect 2502 460 2508 461
rect 2502 456 2503 460
rect 2507 456 2508 460
rect 1326 455 1332 456
rect 2502 455 2508 456
rect 111 450 115 451
rect 111 445 115 446
rect 135 450 139 451
rect 135 445 139 446
rect 191 450 195 451
rect 191 445 195 446
rect 231 450 235 451
rect 231 445 235 446
rect 247 450 251 451
rect 247 445 251 446
rect 303 450 307 451
rect 303 445 307 446
rect 351 450 355 451
rect 351 445 355 446
rect 383 450 387 451
rect 383 445 387 446
rect 471 450 475 451
rect 471 445 475 446
rect 567 450 571 451
rect 567 445 571 446
rect 599 450 603 451
rect 599 445 603 446
rect 671 450 675 451
rect 671 445 675 446
rect 719 450 723 451
rect 719 445 723 446
rect 783 450 787 451
rect 783 445 787 446
rect 831 450 835 451
rect 831 445 835 446
rect 895 450 899 451
rect 895 445 899 446
rect 935 450 939 451
rect 935 445 939 446
rect 1007 450 1011 451
rect 1007 445 1011 446
rect 1039 450 1043 451
rect 1039 445 1043 446
rect 1127 450 1131 451
rect 1127 445 1131 446
rect 1143 450 1147 451
rect 1143 445 1147 446
rect 1223 450 1227 451
rect 1223 445 1227 446
rect 1287 450 1291 451
rect 1287 445 1291 446
rect 112 442 114 445
rect 134 444 140 445
rect 110 441 116 442
rect 110 437 111 441
rect 115 437 116 441
rect 134 440 135 444
rect 139 440 140 444
rect 134 439 140 440
rect 190 444 196 445
rect 190 440 191 444
rect 195 440 196 444
rect 190 439 196 440
rect 246 444 252 445
rect 246 440 247 444
rect 251 440 252 444
rect 246 439 252 440
rect 302 444 308 445
rect 302 440 303 444
rect 307 440 308 444
rect 302 439 308 440
rect 382 444 388 445
rect 382 440 383 444
rect 387 440 388 444
rect 382 439 388 440
rect 470 444 476 445
rect 470 440 471 444
rect 475 440 476 444
rect 470 439 476 440
rect 566 444 572 445
rect 566 440 567 444
rect 571 440 572 444
rect 566 439 572 440
rect 670 444 676 445
rect 670 440 671 444
rect 675 440 676 444
rect 670 439 676 440
rect 782 444 788 445
rect 782 440 783 444
rect 787 440 788 444
rect 782 439 788 440
rect 894 444 900 445
rect 894 440 895 444
rect 899 440 900 444
rect 894 439 900 440
rect 1006 444 1012 445
rect 1006 440 1007 444
rect 1011 440 1012 444
rect 1006 439 1012 440
rect 1126 444 1132 445
rect 1126 440 1127 444
rect 1131 440 1132 444
rect 1126 439 1132 440
rect 1222 444 1228 445
rect 1222 440 1223 444
rect 1227 440 1228 444
rect 1288 442 1290 445
rect 1326 443 1332 444
rect 1222 439 1228 440
rect 1286 441 1292 442
rect 110 436 116 437
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1326 439 1327 443
rect 1331 439 1332 443
rect 2502 443 2508 444
rect 1326 438 1332 439
rect 1350 440 1356 441
rect 1286 436 1292 437
rect 1328 431 1330 438
rect 1350 436 1351 440
rect 1355 436 1356 440
rect 1350 435 1356 436
rect 1414 440 1420 441
rect 1414 436 1415 440
rect 1419 436 1420 440
rect 1414 435 1420 436
rect 1502 440 1508 441
rect 1502 436 1503 440
rect 1507 436 1508 440
rect 1502 435 1508 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1694 440 1700 441
rect 1694 436 1695 440
rect 1699 436 1700 440
rect 1694 435 1700 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1910 440 1916 441
rect 1910 436 1911 440
rect 1915 436 1916 440
rect 1910 435 1916 436
rect 2038 440 2044 441
rect 2038 436 2039 440
rect 2043 436 2044 440
rect 2038 435 2044 436
rect 2174 440 2180 441
rect 2174 436 2175 440
rect 2179 436 2180 440
rect 2174 435 2180 436
rect 2318 440 2324 441
rect 2318 436 2319 440
rect 2323 436 2324 440
rect 2318 435 2324 436
rect 2438 440 2444 441
rect 2438 436 2439 440
rect 2443 436 2444 440
rect 2502 439 2503 443
rect 2507 439 2508 443
rect 2502 438 2508 439
rect 2438 435 2444 436
rect 1352 431 1354 435
rect 1416 431 1418 435
rect 1504 431 1506 435
rect 1600 431 1602 435
rect 1696 431 1698 435
rect 1800 431 1802 435
rect 1912 431 1914 435
rect 2040 431 2042 435
rect 2176 431 2178 435
rect 2320 431 2322 435
rect 2440 431 2442 435
rect 2504 431 2506 438
rect 1327 430 1331 431
rect 1327 425 1331 426
rect 1351 430 1355 431
rect 1351 425 1355 426
rect 1415 430 1419 431
rect 1415 425 1419 426
rect 1423 430 1427 431
rect 1423 425 1427 426
rect 1503 430 1507 431
rect 1503 425 1507 426
rect 1511 430 1515 431
rect 1511 425 1515 426
rect 1599 430 1603 431
rect 1599 425 1603 426
rect 1679 430 1683 431
rect 1679 425 1683 426
rect 1695 430 1699 431
rect 1695 425 1699 426
rect 1775 430 1779 431
rect 1775 425 1779 426
rect 1799 430 1803 431
rect 1799 425 1803 426
rect 1887 430 1891 431
rect 1887 425 1891 426
rect 1911 430 1915 431
rect 1911 425 1915 426
rect 2015 430 2019 431
rect 2015 425 2019 426
rect 2039 430 2043 431
rect 2039 425 2043 426
rect 2159 430 2163 431
rect 2159 425 2163 426
rect 2175 430 2179 431
rect 2175 425 2179 426
rect 2311 430 2315 431
rect 2311 425 2315 426
rect 2319 430 2323 431
rect 2319 425 2323 426
rect 2439 430 2443 431
rect 2439 425 2443 426
rect 2503 430 2507 431
rect 2503 425 2507 426
rect 110 424 116 425
rect 1286 424 1292 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 150 423 156 424
rect 150 419 151 423
rect 155 419 156 423
rect 112 391 114 419
rect 150 418 156 419
rect 206 423 212 424
rect 206 419 207 423
rect 211 419 212 423
rect 206 418 212 419
rect 262 423 268 424
rect 262 419 263 423
rect 267 419 268 423
rect 262 418 268 419
rect 318 423 324 424
rect 318 419 319 423
rect 323 419 324 423
rect 318 418 324 419
rect 398 423 404 424
rect 398 419 399 423
rect 403 419 404 423
rect 398 418 404 419
rect 486 423 492 424
rect 486 419 487 423
rect 491 419 492 423
rect 486 418 492 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 686 423 692 424
rect 686 419 687 423
rect 691 419 692 423
rect 686 418 692 419
rect 798 423 804 424
rect 798 419 799 423
rect 803 419 804 423
rect 798 418 804 419
rect 910 423 916 424
rect 910 419 911 423
rect 915 419 916 423
rect 910 418 916 419
rect 1022 423 1028 424
rect 1022 419 1023 423
rect 1027 419 1028 423
rect 1022 418 1028 419
rect 1142 423 1148 424
rect 1142 419 1143 423
rect 1147 419 1148 423
rect 1142 418 1148 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1286 420 1287 424
rect 1291 420 1292 424
rect 1328 422 1330 425
rect 1350 424 1356 425
rect 1286 419 1292 420
rect 1326 421 1332 422
rect 1238 418 1244 419
rect 152 391 154 418
rect 208 391 210 418
rect 264 391 266 418
rect 320 391 322 418
rect 400 391 402 418
rect 488 391 490 418
rect 584 391 586 418
rect 688 391 690 418
rect 800 391 802 418
rect 912 391 914 418
rect 1024 391 1026 418
rect 1144 391 1146 418
rect 1240 391 1242 418
rect 1288 391 1290 419
rect 1326 417 1327 421
rect 1331 417 1332 421
rect 1350 420 1351 424
rect 1355 420 1356 424
rect 1350 419 1356 420
rect 1422 424 1428 425
rect 1422 420 1423 424
rect 1427 420 1428 424
rect 1422 419 1428 420
rect 1510 424 1516 425
rect 1510 420 1511 424
rect 1515 420 1516 424
rect 1510 419 1516 420
rect 1598 424 1604 425
rect 1598 420 1599 424
rect 1603 420 1604 424
rect 1598 419 1604 420
rect 1678 424 1684 425
rect 1678 420 1679 424
rect 1683 420 1684 424
rect 1678 419 1684 420
rect 1774 424 1780 425
rect 1774 420 1775 424
rect 1779 420 1780 424
rect 1774 419 1780 420
rect 1886 424 1892 425
rect 1886 420 1887 424
rect 1891 420 1892 424
rect 1886 419 1892 420
rect 2014 424 2020 425
rect 2014 420 2015 424
rect 2019 420 2020 424
rect 2014 419 2020 420
rect 2158 424 2164 425
rect 2158 420 2159 424
rect 2163 420 2164 424
rect 2158 419 2164 420
rect 2310 424 2316 425
rect 2310 420 2311 424
rect 2315 420 2316 424
rect 2310 419 2316 420
rect 2438 424 2444 425
rect 2438 420 2439 424
rect 2443 420 2444 424
rect 2504 422 2506 425
rect 2438 419 2444 420
rect 2502 421 2508 422
rect 1326 416 1332 417
rect 2502 417 2503 421
rect 2507 417 2508 421
rect 2502 416 2508 417
rect 1326 404 1332 405
rect 2502 404 2508 405
rect 1326 400 1327 404
rect 1331 400 1332 404
rect 1326 399 1332 400
rect 1366 403 1372 404
rect 1366 399 1367 403
rect 1371 399 1372 403
rect 111 390 115 391
rect 111 385 115 386
rect 151 390 155 391
rect 151 385 155 386
rect 207 390 211 391
rect 207 385 211 386
rect 263 390 267 391
rect 263 385 267 386
rect 279 390 283 391
rect 279 385 283 386
rect 319 390 323 391
rect 319 385 323 386
rect 359 390 363 391
rect 359 385 363 386
rect 399 390 403 391
rect 399 385 403 386
rect 431 390 435 391
rect 431 385 435 386
rect 487 390 491 391
rect 487 385 491 386
rect 511 390 515 391
rect 511 385 515 386
rect 583 390 587 391
rect 583 385 587 386
rect 591 390 595 391
rect 591 385 595 386
rect 671 390 675 391
rect 671 385 675 386
rect 687 390 691 391
rect 687 385 691 386
rect 751 390 755 391
rect 751 385 755 386
rect 799 390 803 391
rect 799 385 803 386
rect 823 390 827 391
rect 823 385 827 386
rect 895 390 899 391
rect 895 385 899 386
rect 911 390 915 391
rect 911 385 915 386
rect 967 390 971 391
rect 967 385 971 386
rect 1023 390 1027 391
rect 1023 385 1027 386
rect 1039 390 1043 391
rect 1039 385 1043 386
rect 1111 390 1115 391
rect 1111 385 1115 386
rect 1143 390 1147 391
rect 1143 385 1147 386
rect 1183 390 1187 391
rect 1183 385 1187 386
rect 1239 390 1243 391
rect 1239 385 1243 386
rect 1287 390 1291 391
rect 1287 385 1291 386
rect 112 365 114 385
rect 152 366 154 385
rect 208 366 210 385
rect 280 366 282 385
rect 360 366 362 385
rect 432 366 434 385
rect 512 366 514 385
rect 592 366 594 385
rect 672 366 674 385
rect 752 366 754 385
rect 824 366 826 385
rect 896 366 898 385
rect 968 366 970 385
rect 1040 366 1042 385
rect 1112 366 1114 385
rect 1184 366 1186 385
rect 1240 366 1242 385
rect 150 365 156 366
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 150 361 151 365
rect 155 361 156 365
rect 150 360 156 361
rect 206 365 212 366
rect 206 361 207 365
rect 211 361 212 365
rect 206 360 212 361
rect 278 365 284 366
rect 278 361 279 365
rect 283 361 284 365
rect 278 360 284 361
rect 358 365 364 366
rect 358 361 359 365
rect 363 361 364 365
rect 358 360 364 361
rect 430 365 436 366
rect 430 361 431 365
rect 435 361 436 365
rect 430 360 436 361
rect 510 365 516 366
rect 510 361 511 365
rect 515 361 516 365
rect 510 360 516 361
rect 590 365 596 366
rect 590 361 591 365
rect 595 361 596 365
rect 590 360 596 361
rect 670 365 676 366
rect 670 361 671 365
rect 675 361 676 365
rect 670 360 676 361
rect 750 365 756 366
rect 750 361 751 365
rect 755 361 756 365
rect 750 360 756 361
rect 822 365 828 366
rect 822 361 823 365
rect 827 361 828 365
rect 822 360 828 361
rect 894 365 900 366
rect 894 361 895 365
rect 899 361 900 365
rect 894 360 900 361
rect 966 365 972 366
rect 966 361 967 365
rect 971 361 972 365
rect 966 360 972 361
rect 1038 365 1044 366
rect 1038 361 1039 365
rect 1043 361 1044 365
rect 1038 360 1044 361
rect 1110 365 1116 366
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 1182 365 1188 366
rect 1182 361 1183 365
rect 1187 361 1188 365
rect 1182 360 1188 361
rect 1238 365 1244 366
rect 1288 365 1290 385
rect 1328 375 1330 399
rect 1366 398 1372 399
rect 1438 403 1444 404
rect 1438 399 1439 403
rect 1443 399 1444 403
rect 1438 398 1444 399
rect 1526 403 1532 404
rect 1526 399 1527 403
rect 1531 399 1532 403
rect 1526 398 1532 399
rect 1614 403 1620 404
rect 1614 399 1615 403
rect 1619 399 1620 403
rect 1614 398 1620 399
rect 1694 403 1700 404
rect 1694 399 1695 403
rect 1699 399 1700 403
rect 1694 398 1700 399
rect 1790 403 1796 404
rect 1790 399 1791 403
rect 1795 399 1796 403
rect 1790 398 1796 399
rect 1902 403 1908 404
rect 1902 399 1903 403
rect 1907 399 1908 403
rect 1902 398 1908 399
rect 2030 403 2036 404
rect 2030 399 2031 403
rect 2035 399 2036 403
rect 2030 398 2036 399
rect 2174 403 2180 404
rect 2174 399 2175 403
rect 2179 399 2180 403
rect 2174 398 2180 399
rect 2326 403 2332 404
rect 2326 399 2327 403
rect 2331 399 2332 403
rect 2326 398 2332 399
rect 2454 403 2460 404
rect 2454 399 2455 403
rect 2459 399 2460 403
rect 2502 400 2503 404
rect 2507 400 2508 404
rect 2502 399 2508 400
rect 2454 398 2460 399
rect 1368 375 1370 398
rect 1440 375 1442 398
rect 1528 375 1530 398
rect 1616 375 1618 398
rect 1696 375 1698 398
rect 1792 375 1794 398
rect 1904 375 1906 398
rect 2032 375 2034 398
rect 2176 375 2178 398
rect 2328 375 2330 398
rect 2456 375 2458 398
rect 2504 375 2506 399
rect 1327 374 1331 375
rect 1327 369 1331 370
rect 1367 374 1371 375
rect 1367 369 1371 370
rect 1439 374 1443 375
rect 1439 369 1443 370
rect 1527 374 1531 375
rect 1527 369 1531 370
rect 1615 374 1619 375
rect 1615 369 1619 370
rect 1679 374 1683 375
rect 1679 369 1683 370
rect 1695 374 1699 375
rect 1695 369 1699 370
rect 1735 374 1739 375
rect 1735 369 1739 370
rect 1791 374 1795 375
rect 1791 369 1795 370
rect 1807 374 1811 375
rect 1807 369 1811 370
rect 1903 374 1907 375
rect 1903 369 1907 370
rect 2023 374 2027 375
rect 2023 369 2027 370
rect 2031 374 2035 375
rect 2031 369 2035 370
rect 2159 374 2163 375
rect 2159 369 2163 370
rect 2175 374 2179 375
rect 2175 369 2179 370
rect 2303 374 2307 375
rect 2303 369 2307 370
rect 2327 374 2331 375
rect 2327 369 2331 370
rect 2455 374 2459 375
rect 2455 369 2459 370
rect 2503 374 2507 375
rect 2503 369 2507 370
rect 1238 361 1239 365
rect 1243 361 1244 365
rect 1238 360 1244 361
rect 1286 364 1292 365
rect 1286 360 1287 364
rect 1291 360 1292 364
rect 110 359 116 360
rect 1286 359 1292 360
rect 1328 349 1330 369
rect 1680 350 1682 369
rect 1736 350 1738 369
rect 1808 350 1810 369
rect 1904 350 1906 369
rect 2024 350 2026 369
rect 2160 350 2162 369
rect 2304 350 2306 369
rect 2456 350 2458 369
rect 1678 349 1684 350
rect 1326 348 1332 349
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 1286 347 1292 348
rect 110 342 116 343
rect 134 344 140 345
rect 112 331 114 342
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 190 344 196 345
rect 190 340 191 344
rect 195 340 196 344
rect 190 339 196 340
rect 262 344 268 345
rect 262 340 263 344
rect 267 340 268 344
rect 262 339 268 340
rect 342 344 348 345
rect 342 340 343 344
rect 347 340 348 344
rect 342 339 348 340
rect 414 344 420 345
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 806 344 812 345
rect 806 340 807 344
rect 811 340 812 344
rect 806 339 812 340
rect 878 344 884 345
rect 878 340 879 344
rect 883 340 884 344
rect 878 339 884 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1022 344 1028 345
rect 1022 340 1023 344
rect 1027 340 1028 344
rect 1022 339 1028 340
rect 1094 344 1100 345
rect 1094 340 1095 344
rect 1099 340 1100 344
rect 1094 339 1100 340
rect 1166 344 1172 345
rect 1166 340 1167 344
rect 1171 340 1172 344
rect 1166 339 1172 340
rect 1222 344 1228 345
rect 1222 340 1223 344
rect 1227 340 1228 344
rect 1286 343 1287 347
rect 1291 343 1292 347
rect 1326 344 1327 348
rect 1331 344 1332 348
rect 1678 345 1679 349
rect 1683 345 1684 349
rect 1678 344 1684 345
rect 1734 349 1740 350
rect 1734 345 1735 349
rect 1739 345 1740 349
rect 1734 344 1740 345
rect 1806 349 1812 350
rect 1806 345 1807 349
rect 1811 345 1812 349
rect 1806 344 1812 345
rect 1902 349 1908 350
rect 1902 345 1903 349
rect 1907 345 1908 349
rect 1902 344 1908 345
rect 2022 349 2028 350
rect 2022 345 2023 349
rect 2027 345 2028 349
rect 2022 344 2028 345
rect 2158 349 2164 350
rect 2158 345 2159 349
rect 2163 345 2164 349
rect 2158 344 2164 345
rect 2302 349 2308 350
rect 2302 345 2303 349
rect 2307 345 2308 349
rect 2302 344 2308 345
rect 2454 349 2460 350
rect 2504 349 2506 369
rect 2454 345 2455 349
rect 2459 345 2460 349
rect 2454 344 2460 345
rect 2502 348 2508 349
rect 2502 344 2503 348
rect 2507 344 2508 348
rect 1326 343 1332 344
rect 2502 343 2508 344
rect 1286 342 1292 343
rect 1222 339 1228 340
rect 136 331 138 339
rect 192 331 194 339
rect 264 331 266 339
rect 344 331 346 339
rect 416 331 418 339
rect 496 331 498 339
rect 576 331 578 339
rect 656 331 658 339
rect 736 331 738 339
rect 808 331 810 339
rect 880 331 882 339
rect 952 331 954 339
rect 1024 331 1026 339
rect 1096 331 1098 339
rect 1168 331 1170 339
rect 1224 331 1226 339
rect 1288 331 1290 342
rect 1326 331 1332 332
rect 111 330 115 331
rect 111 325 115 326
rect 135 330 139 331
rect 135 325 139 326
rect 191 330 195 331
rect 191 325 195 326
rect 199 330 203 331
rect 199 325 203 326
rect 263 330 267 331
rect 263 325 267 326
rect 287 330 291 331
rect 287 325 291 326
rect 343 330 347 331
rect 343 325 347 326
rect 375 330 379 331
rect 375 325 379 326
rect 415 330 419 331
rect 415 325 419 326
rect 455 330 459 331
rect 455 325 459 326
rect 495 330 499 331
rect 495 325 499 326
rect 543 330 547 331
rect 543 325 547 326
rect 575 330 579 331
rect 575 325 579 326
rect 631 330 635 331
rect 631 325 635 326
rect 655 330 659 331
rect 655 325 659 326
rect 727 330 731 331
rect 727 325 731 326
rect 735 330 739 331
rect 735 325 739 326
rect 807 330 811 331
rect 807 325 811 326
rect 823 330 827 331
rect 823 325 827 326
rect 879 330 883 331
rect 879 325 883 326
rect 927 330 931 331
rect 927 325 931 326
rect 951 330 955 331
rect 951 325 955 326
rect 1023 330 1027 331
rect 1023 325 1027 326
rect 1031 330 1035 331
rect 1031 325 1035 326
rect 1095 330 1099 331
rect 1095 325 1099 326
rect 1135 330 1139 331
rect 1135 325 1139 326
rect 1167 330 1171 331
rect 1167 325 1171 326
rect 1223 330 1227 331
rect 1223 325 1227 326
rect 1287 330 1291 331
rect 1326 327 1327 331
rect 1331 327 1332 331
rect 2502 331 2508 332
rect 1326 326 1332 327
rect 1662 328 1668 329
rect 1287 325 1291 326
rect 112 322 114 325
rect 134 324 140 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 134 320 135 324
rect 139 320 140 324
rect 134 319 140 320
rect 198 324 204 325
rect 198 320 199 324
rect 203 320 204 324
rect 198 319 204 320
rect 286 324 292 325
rect 286 320 287 324
rect 291 320 292 324
rect 286 319 292 320
rect 374 324 380 325
rect 374 320 375 324
rect 379 320 380 324
rect 374 319 380 320
rect 454 324 460 325
rect 454 320 455 324
rect 459 320 460 324
rect 454 319 460 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 630 324 636 325
rect 630 320 631 324
rect 635 320 636 324
rect 630 319 636 320
rect 726 324 732 325
rect 726 320 727 324
rect 731 320 732 324
rect 726 319 732 320
rect 822 324 828 325
rect 822 320 823 324
rect 827 320 828 324
rect 822 319 828 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 1030 324 1036 325
rect 1030 320 1031 324
rect 1035 320 1036 324
rect 1030 319 1036 320
rect 1134 324 1140 325
rect 1134 320 1135 324
rect 1139 320 1140 324
rect 1134 319 1140 320
rect 1222 324 1228 325
rect 1222 320 1223 324
rect 1227 320 1228 324
rect 1288 322 1290 325
rect 1328 323 1330 326
rect 1662 324 1663 328
rect 1667 324 1668 328
rect 1662 323 1668 324
rect 1718 328 1724 329
rect 1718 324 1719 328
rect 1723 324 1724 328
rect 1718 323 1724 324
rect 1790 328 1796 329
rect 1790 324 1791 328
rect 1795 324 1796 328
rect 1790 323 1796 324
rect 1886 328 1892 329
rect 1886 324 1887 328
rect 1891 324 1892 328
rect 1886 323 1892 324
rect 2006 328 2012 329
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 2142 328 2148 329
rect 2142 324 2143 328
rect 2147 324 2148 328
rect 2142 323 2148 324
rect 2286 328 2292 329
rect 2286 324 2287 328
rect 2291 324 2292 328
rect 2286 323 2292 324
rect 2438 328 2444 329
rect 2438 324 2439 328
rect 2443 324 2444 328
rect 2502 327 2503 331
rect 2507 327 2508 331
rect 2502 326 2508 327
rect 2438 323 2444 324
rect 2504 323 2506 326
rect 1327 322 1331 323
rect 1222 319 1228 320
rect 1286 321 1292 322
rect 110 316 116 317
rect 1286 317 1287 321
rect 1291 317 1292 321
rect 1327 317 1331 318
rect 1351 322 1355 323
rect 1351 317 1355 318
rect 1431 322 1435 323
rect 1431 317 1435 318
rect 1527 322 1531 323
rect 1527 317 1531 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1663 322 1667 323
rect 1663 317 1667 318
rect 1711 322 1715 323
rect 1711 317 1715 318
rect 1719 322 1723 323
rect 1719 317 1723 318
rect 1791 322 1795 323
rect 1791 317 1795 318
rect 1807 322 1811 323
rect 1807 317 1811 318
rect 1887 322 1891 323
rect 1887 317 1891 318
rect 1911 322 1915 323
rect 1911 317 1915 318
rect 2007 322 2011 323
rect 2007 317 2011 318
rect 2023 322 2027 323
rect 2023 317 2027 318
rect 2143 322 2147 323
rect 2143 317 2147 318
rect 2151 322 2155 323
rect 2151 317 2155 318
rect 2287 322 2291 323
rect 2287 317 2291 318
rect 2423 322 2427 323
rect 2423 317 2427 318
rect 2439 322 2443 323
rect 2439 317 2443 318
rect 2503 322 2507 323
rect 2503 317 2507 318
rect 1286 316 1292 317
rect 1328 314 1330 317
rect 1350 316 1356 317
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1350 312 1351 316
rect 1355 312 1356 316
rect 1350 311 1356 312
rect 1430 316 1436 317
rect 1430 312 1431 316
rect 1435 312 1436 316
rect 1430 311 1436 312
rect 1526 316 1532 317
rect 1526 312 1527 316
rect 1531 312 1532 316
rect 1526 311 1532 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1710 316 1716 317
rect 1710 312 1711 316
rect 1715 312 1716 316
rect 1710 311 1716 312
rect 1806 316 1812 317
rect 1806 312 1807 316
rect 1811 312 1812 316
rect 1806 311 1812 312
rect 1910 316 1916 317
rect 1910 312 1911 316
rect 1915 312 1916 316
rect 1910 311 1916 312
rect 2022 316 2028 317
rect 2022 312 2023 316
rect 2027 312 2028 316
rect 2022 311 2028 312
rect 2150 316 2156 317
rect 2150 312 2151 316
rect 2155 312 2156 316
rect 2150 311 2156 312
rect 2286 316 2292 317
rect 2286 312 2287 316
rect 2291 312 2292 316
rect 2286 311 2292 312
rect 2422 316 2428 317
rect 2422 312 2423 316
rect 2427 312 2428 316
rect 2504 314 2506 317
rect 2422 311 2428 312
rect 2502 313 2508 314
rect 1326 308 1332 309
rect 2502 309 2503 313
rect 2507 309 2508 313
rect 2502 308 2508 309
rect 110 304 116 305
rect 1286 304 1292 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 150 303 156 304
rect 150 299 151 303
rect 155 299 156 303
rect 112 271 114 299
rect 150 298 156 299
rect 214 303 220 304
rect 214 299 215 303
rect 219 299 220 303
rect 214 298 220 299
rect 302 303 308 304
rect 302 299 303 303
rect 307 299 308 303
rect 302 298 308 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 470 303 476 304
rect 470 299 471 303
rect 475 299 476 303
rect 470 298 476 299
rect 558 303 564 304
rect 558 299 559 303
rect 563 299 564 303
rect 558 298 564 299
rect 646 303 652 304
rect 646 299 647 303
rect 651 299 652 303
rect 646 298 652 299
rect 742 303 748 304
rect 742 299 743 303
rect 747 299 748 303
rect 742 298 748 299
rect 838 303 844 304
rect 838 299 839 303
rect 843 299 844 303
rect 838 298 844 299
rect 942 303 948 304
rect 942 299 943 303
rect 947 299 948 303
rect 942 298 948 299
rect 1046 303 1052 304
rect 1046 299 1047 303
rect 1051 299 1052 303
rect 1046 298 1052 299
rect 1150 303 1156 304
rect 1150 299 1151 303
rect 1155 299 1156 303
rect 1150 298 1156 299
rect 1238 303 1244 304
rect 1238 299 1239 303
rect 1243 299 1244 303
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1238 298 1244 299
rect 152 271 154 298
rect 216 271 218 298
rect 304 271 306 298
rect 392 271 394 298
rect 472 271 474 298
rect 560 271 562 298
rect 648 271 650 298
rect 744 271 746 298
rect 840 271 842 298
rect 944 271 946 298
rect 1048 271 1050 298
rect 1152 271 1154 298
rect 1240 271 1242 298
rect 1288 271 1290 299
rect 1326 296 1332 297
rect 2502 296 2508 297
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1326 291 1332 292
rect 1366 295 1372 296
rect 1366 291 1367 295
rect 1371 291 1372 295
rect 111 270 115 271
rect 111 265 115 266
rect 151 270 155 271
rect 151 265 155 266
rect 215 270 219 271
rect 215 265 219 266
rect 231 270 235 271
rect 231 265 235 266
rect 303 270 307 271
rect 303 265 307 266
rect 327 270 331 271
rect 327 265 331 266
rect 391 270 395 271
rect 391 265 395 266
rect 423 270 427 271
rect 423 265 427 266
rect 471 270 475 271
rect 471 265 475 266
rect 519 270 523 271
rect 519 265 523 266
rect 559 270 563 271
rect 559 265 563 266
rect 615 270 619 271
rect 615 265 619 266
rect 647 270 651 271
rect 647 265 651 266
rect 711 270 715 271
rect 711 265 715 266
rect 743 270 747 271
rect 743 265 747 266
rect 807 270 811 271
rect 807 265 811 266
rect 839 270 843 271
rect 839 265 843 266
rect 903 270 907 271
rect 903 265 907 266
rect 943 270 947 271
rect 943 265 947 266
rect 1007 270 1011 271
rect 1007 265 1011 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1111 270 1115 271
rect 1111 265 1115 266
rect 1151 270 1155 271
rect 1151 265 1155 266
rect 1215 270 1219 271
rect 1215 265 1219 266
rect 1239 270 1243 271
rect 1239 265 1243 266
rect 1287 270 1291 271
rect 1328 267 1330 291
rect 1366 290 1372 291
rect 1446 295 1452 296
rect 1446 291 1447 295
rect 1451 291 1452 295
rect 1446 290 1452 291
rect 1542 295 1548 296
rect 1542 291 1543 295
rect 1547 291 1548 295
rect 1542 290 1548 291
rect 1638 295 1644 296
rect 1638 291 1639 295
rect 1643 291 1644 295
rect 1638 290 1644 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1822 295 1828 296
rect 1822 291 1823 295
rect 1827 291 1828 295
rect 1822 290 1828 291
rect 1926 295 1932 296
rect 1926 291 1927 295
rect 1931 291 1932 295
rect 1926 290 1932 291
rect 2038 295 2044 296
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2166 295 2172 296
rect 2166 291 2167 295
rect 2171 291 2172 295
rect 2166 290 2172 291
rect 2302 295 2308 296
rect 2302 291 2303 295
rect 2307 291 2308 295
rect 2302 290 2308 291
rect 2438 295 2444 296
rect 2438 291 2439 295
rect 2443 291 2444 295
rect 2502 292 2503 296
rect 2507 292 2508 296
rect 2502 291 2508 292
rect 2438 290 2444 291
rect 1368 267 1370 290
rect 1448 267 1450 290
rect 1544 267 1546 290
rect 1640 267 1642 290
rect 1728 267 1730 290
rect 1824 267 1826 290
rect 1928 267 1930 290
rect 2040 267 2042 290
rect 2168 267 2170 290
rect 2304 267 2306 290
rect 2440 267 2442 290
rect 2504 267 2506 291
rect 1287 265 1291 266
rect 1327 266 1331 267
rect 112 245 114 265
rect 152 246 154 265
rect 232 246 234 265
rect 328 246 330 265
rect 424 246 426 265
rect 520 246 522 265
rect 616 246 618 265
rect 712 246 714 265
rect 808 246 810 265
rect 904 246 906 265
rect 1008 246 1010 265
rect 1112 246 1114 265
rect 1216 246 1218 265
rect 150 245 156 246
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 150 241 151 245
rect 155 241 156 245
rect 150 240 156 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 230 240 236 241
rect 326 245 332 246
rect 326 241 327 245
rect 331 241 332 245
rect 326 240 332 241
rect 422 245 428 246
rect 422 241 423 245
rect 427 241 428 245
rect 422 240 428 241
rect 518 245 524 246
rect 518 241 519 245
rect 523 241 524 245
rect 518 240 524 241
rect 614 245 620 246
rect 614 241 615 245
rect 619 241 620 245
rect 614 240 620 241
rect 710 245 716 246
rect 710 241 711 245
rect 715 241 716 245
rect 710 240 716 241
rect 806 245 812 246
rect 806 241 807 245
rect 811 241 812 245
rect 806 240 812 241
rect 902 245 908 246
rect 902 241 903 245
rect 907 241 908 245
rect 902 240 908 241
rect 1006 245 1012 246
rect 1006 241 1007 245
rect 1011 241 1012 245
rect 1006 240 1012 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1214 245 1220 246
rect 1288 245 1290 265
rect 1327 261 1331 262
rect 1367 266 1371 267
rect 1367 261 1371 262
rect 1439 266 1443 267
rect 1439 261 1443 262
rect 1447 266 1451 267
rect 1447 261 1451 262
rect 1535 266 1539 267
rect 1535 261 1539 262
rect 1543 266 1547 267
rect 1543 261 1547 262
rect 1631 266 1635 267
rect 1631 261 1635 262
rect 1639 266 1643 267
rect 1639 261 1643 262
rect 1727 266 1731 267
rect 1727 261 1731 262
rect 1815 266 1819 267
rect 1815 261 1819 262
rect 1823 266 1827 267
rect 1823 261 1827 262
rect 1903 266 1907 267
rect 1903 261 1907 262
rect 1927 266 1931 267
rect 1927 261 1931 262
rect 1999 266 2003 267
rect 1999 261 2003 262
rect 2039 266 2043 267
rect 2039 261 2043 262
rect 2103 266 2107 267
rect 2103 261 2107 262
rect 2167 266 2171 267
rect 2167 261 2171 262
rect 2215 266 2219 267
rect 2215 261 2219 262
rect 2303 266 2307 267
rect 2303 261 2307 262
rect 2335 266 2339 267
rect 2335 261 2339 262
rect 2439 266 2443 267
rect 2439 261 2443 262
rect 2455 266 2459 267
rect 2455 261 2459 262
rect 2503 266 2507 267
rect 2503 261 2507 262
rect 1214 241 1215 245
rect 1219 241 1220 245
rect 1214 240 1220 241
rect 1286 244 1292 245
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1328 241 1330 261
rect 1368 242 1370 261
rect 1440 242 1442 261
rect 1536 242 1538 261
rect 1632 242 1634 261
rect 1728 242 1730 261
rect 1816 242 1818 261
rect 1904 242 1906 261
rect 2000 242 2002 261
rect 2104 242 2106 261
rect 2216 242 2218 261
rect 2336 242 2338 261
rect 2456 242 2458 261
rect 1366 241 1372 242
rect 110 239 116 240
rect 1286 239 1292 240
rect 1326 240 1332 241
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1438 241 1444 242
rect 1438 237 1439 241
rect 1443 237 1444 241
rect 1438 236 1444 237
rect 1534 241 1540 242
rect 1534 237 1535 241
rect 1539 237 1540 241
rect 1534 236 1540 237
rect 1630 241 1636 242
rect 1630 237 1631 241
rect 1635 237 1636 241
rect 1630 236 1636 237
rect 1726 241 1732 242
rect 1726 237 1727 241
rect 1731 237 1732 241
rect 1726 236 1732 237
rect 1814 241 1820 242
rect 1814 237 1815 241
rect 1819 237 1820 241
rect 1814 236 1820 237
rect 1902 241 1908 242
rect 1902 237 1903 241
rect 1907 237 1908 241
rect 1902 236 1908 237
rect 1998 241 2004 242
rect 1998 237 1999 241
rect 2003 237 2004 241
rect 1998 236 2004 237
rect 2102 241 2108 242
rect 2102 237 2103 241
rect 2107 237 2108 241
rect 2102 236 2108 237
rect 2214 241 2220 242
rect 2214 237 2215 241
rect 2219 237 2220 241
rect 2214 236 2220 237
rect 2334 241 2340 242
rect 2334 237 2335 241
rect 2339 237 2340 241
rect 2334 236 2340 237
rect 2454 241 2460 242
rect 2504 241 2506 261
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2454 236 2460 237
rect 2502 240 2508 241
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 1326 235 1332 236
rect 2502 235 2508 236
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1286 227 1292 228
rect 110 222 116 223
rect 134 224 140 225
rect 112 211 114 222
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 214 224 220 225
rect 214 220 215 224
rect 219 220 220 224
rect 214 219 220 220
rect 310 224 316 225
rect 310 220 311 224
rect 315 220 316 224
rect 310 219 316 220
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 502 224 508 225
rect 502 220 503 224
rect 507 220 508 224
rect 502 219 508 220
rect 598 224 604 225
rect 598 220 599 224
rect 603 220 604 224
rect 598 219 604 220
rect 694 224 700 225
rect 694 220 695 224
rect 699 220 700 224
rect 694 219 700 220
rect 790 224 796 225
rect 790 220 791 224
rect 795 220 796 224
rect 790 219 796 220
rect 886 224 892 225
rect 886 220 887 224
rect 891 220 892 224
rect 886 219 892 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1094 224 1100 225
rect 1094 220 1095 224
rect 1099 220 1100 224
rect 1094 219 1100 220
rect 1198 224 1204 225
rect 1198 220 1199 224
rect 1203 220 1204 224
rect 1286 223 1287 227
rect 1291 223 1292 227
rect 1286 222 1292 223
rect 1326 223 1332 224
rect 1198 219 1204 220
rect 136 211 138 219
rect 216 211 218 219
rect 312 211 314 219
rect 408 211 410 219
rect 504 211 506 219
rect 600 211 602 219
rect 696 211 698 219
rect 792 211 794 219
rect 888 211 890 219
rect 992 211 994 219
rect 1096 211 1098 219
rect 1200 211 1202 219
rect 1288 211 1290 222
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1328 211 1330 218
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1422 220 1428 221
rect 1422 216 1423 220
rect 1427 216 1428 220
rect 1422 215 1428 216
rect 1518 220 1524 221
rect 1518 216 1519 220
rect 1523 216 1524 220
rect 1518 215 1524 216
rect 1614 220 1620 221
rect 1614 216 1615 220
rect 1619 216 1620 220
rect 1614 215 1620 216
rect 1710 220 1716 221
rect 1710 216 1711 220
rect 1715 216 1716 220
rect 1710 215 1716 216
rect 1798 220 1804 221
rect 1798 216 1799 220
rect 1803 216 1804 220
rect 1798 215 1804 216
rect 1886 220 1892 221
rect 1886 216 1887 220
rect 1891 216 1892 220
rect 1886 215 1892 216
rect 1982 220 1988 221
rect 1982 216 1983 220
rect 1987 216 1988 220
rect 1982 215 1988 216
rect 2086 220 2092 221
rect 2086 216 2087 220
rect 2091 216 2092 220
rect 2086 215 2092 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2318 220 2324 221
rect 2318 216 2319 220
rect 2323 216 2324 220
rect 2318 215 2324 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 1352 211 1354 215
rect 1424 211 1426 215
rect 1520 211 1522 215
rect 1616 211 1618 215
rect 1712 211 1714 215
rect 1800 211 1802 215
rect 1888 211 1890 215
rect 1984 211 1986 215
rect 2088 211 2090 215
rect 2200 211 2202 215
rect 2320 211 2322 215
rect 2440 211 2442 215
rect 2504 211 2506 218
rect 111 210 115 211
rect 111 205 115 206
rect 135 210 139 211
rect 135 205 139 206
rect 159 210 163 211
rect 159 205 163 206
rect 215 210 219 211
rect 215 205 219 206
rect 239 210 243 211
rect 239 205 243 206
rect 311 210 315 211
rect 311 205 315 206
rect 327 210 331 211
rect 327 205 331 206
rect 407 210 411 211
rect 407 205 411 206
rect 415 210 419 211
rect 415 205 419 206
rect 503 210 507 211
rect 503 205 507 206
rect 511 210 515 211
rect 511 205 515 206
rect 599 210 603 211
rect 599 205 603 206
rect 607 210 611 211
rect 607 205 611 206
rect 695 210 699 211
rect 695 205 699 206
rect 783 210 787 211
rect 783 205 787 206
rect 791 210 795 211
rect 791 205 795 206
rect 871 210 875 211
rect 871 205 875 206
rect 887 210 891 211
rect 887 205 891 206
rect 959 210 963 211
rect 959 205 963 206
rect 991 210 995 211
rect 991 205 995 206
rect 1047 210 1051 211
rect 1047 205 1051 206
rect 1095 210 1099 211
rect 1095 205 1099 206
rect 1135 210 1139 211
rect 1135 205 1139 206
rect 1199 210 1203 211
rect 1199 205 1203 206
rect 1287 210 1291 211
rect 1287 205 1291 206
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1351 210 1355 211
rect 1351 205 1355 206
rect 1391 210 1395 211
rect 1391 205 1395 206
rect 1423 210 1427 211
rect 1423 205 1427 206
rect 1495 210 1499 211
rect 1495 205 1499 206
rect 1519 210 1523 211
rect 1519 205 1523 206
rect 1599 210 1603 211
rect 1599 205 1603 206
rect 1615 210 1619 211
rect 1615 205 1619 206
rect 1711 210 1715 211
rect 1711 205 1715 206
rect 1799 210 1803 211
rect 1799 205 1803 206
rect 1815 210 1819 211
rect 1815 205 1819 206
rect 1887 210 1891 211
rect 1887 205 1891 206
rect 1919 210 1923 211
rect 1919 205 1923 206
rect 1983 210 1987 211
rect 1983 205 1987 206
rect 2015 210 2019 211
rect 2015 205 2019 206
rect 2087 210 2091 211
rect 2087 205 2091 206
rect 2111 210 2115 211
rect 2111 205 2115 206
rect 2199 210 2203 211
rect 2199 205 2203 206
rect 2287 210 2291 211
rect 2287 205 2291 206
rect 2319 210 2323 211
rect 2319 205 2323 206
rect 2375 210 2379 211
rect 2375 205 2379 206
rect 2439 210 2443 211
rect 2439 205 2443 206
rect 2503 210 2507 211
rect 2503 205 2507 206
rect 112 202 114 205
rect 158 204 164 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 158 200 159 204
rect 163 200 164 204
rect 158 199 164 200
rect 238 204 244 205
rect 238 200 239 204
rect 243 200 244 204
rect 238 199 244 200
rect 326 204 332 205
rect 326 200 327 204
rect 331 200 332 204
rect 326 199 332 200
rect 414 204 420 205
rect 414 200 415 204
rect 419 200 420 204
rect 414 199 420 200
rect 510 204 516 205
rect 510 200 511 204
rect 515 200 516 204
rect 510 199 516 200
rect 606 204 612 205
rect 606 200 607 204
rect 611 200 612 204
rect 606 199 612 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 782 204 788 205
rect 782 200 783 204
rect 787 200 788 204
rect 782 199 788 200
rect 870 204 876 205
rect 870 200 871 204
rect 875 200 876 204
rect 870 199 876 200
rect 958 204 964 205
rect 958 200 959 204
rect 963 200 964 204
rect 958 199 964 200
rect 1046 204 1052 205
rect 1046 200 1047 204
rect 1051 200 1052 204
rect 1046 199 1052 200
rect 1134 204 1140 205
rect 1134 200 1135 204
rect 1139 200 1140 204
rect 1288 202 1290 205
rect 1328 202 1330 205
rect 1390 204 1396 205
rect 1134 199 1140 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1390 200 1391 204
rect 1395 200 1396 204
rect 1390 199 1396 200
rect 1494 204 1500 205
rect 1494 200 1495 204
rect 1499 200 1500 204
rect 1494 199 1500 200
rect 1598 204 1604 205
rect 1598 200 1599 204
rect 1603 200 1604 204
rect 1598 199 1604 200
rect 1710 204 1716 205
rect 1710 200 1711 204
rect 1715 200 1716 204
rect 1710 199 1716 200
rect 1814 204 1820 205
rect 1814 200 1815 204
rect 1819 200 1820 204
rect 1814 199 1820 200
rect 1918 204 1924 205
rect 1918 200 1919 204
rect 1923 200 1924 204
rect 1918 199 1924 200
rect 2014 204 2020 205
rect 2014 200 2015 204
rect 2019 200 2020 204
rect 2014 199 2020 200
rect 2110 204 2116 205
rect 2110 200 2111 204
rect 2115 200 2116 204
rect 2110 199 2116 200
rect 2198 204 2204 205
rect 2198 200 2199 204
rect 2203 200 2204 204
rect 2198 199 2204 200
rect 2286 204 2292 205
rect 2286 200 2287 204
rect 2291 200 2292 204
rect 2286 199 2292 200
rect 2374 204 2380 205
rect 2374 200 2375 204
rect 2379 200 2380 204
rect 2374 199 2380 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2504 202 2506 205
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 174 183 180 184
rect 174 179 175 183
rect 179 179 180 183
rect 112 139 114 179
rect 174 178 180 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 179 260 183
rect 254 178 260 179
rect 342 183 348 184
rect 342 179 343 183
rect 347 179 348 183
rect 342 178 348 179
rect 430 183 436 184
rect 430 179 431 183
rect 435 179 436 183
rect 430 178 436 179
rect 526 183 532 184
rect 526 179 527 183
rect 531 179 532 183
rect 526 178 532 179
rect 622 183 628 184
rect 622 179 623 183
rect 627 179 628 183
rect 622 178 628 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 798 183 804 184
rect 798 179 799 183
rect 803 179 804 183
rect 798 178 804 179
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 974 183 980 184
rect 974 179 975 183
rect 979 179 980 183
rect 974 178 980 179
rect 1062 183 1068 184
rect 1062 179 1063 183
rect 1067 179 1068 183
rect 1062 178 1068 179
rect 1150 183 1156 184
rect 1150 179 1151 183
rect 1155 179 1156 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1406 183 1412 184
rect 1406 179 1407 183
rect 1411 179 1412 183
rect 1150 178 1156 179
rect 176 139 178 178
rect 256 139 258 178
rect 344 139 346 178
rect 432 139 434 178
rect 528 139 530 178
rect 624 139 626 178
rect 712 139 714 178
rect 800 139 802 178
rect 888 139 890 178
rect 976 139 978 178
rect 1064 139 1066 178
rect 1152 139 1154 178
rect 1288 139 1290 179
rect 1328 139 1330 179
rect 1406 178 1412 179
rect 1510 183 1516 184
rect 1510 179 1511 183
rect 1515 179 1516 183
rect 1510 178 1516 179
rect 1614 183 1620 184
rect 1614 179 1615 183
rect 1619 179 1620 183
rect 1614 178 1620 179
rect 1726 183 1732 184
rect 1726 179 1727 183
rect 1731 179 1732 183
rect 1726 178 1732 179
rect 1830 183 1836 184
rect 1830 179 1831 183
rect 1835 179 1836 183
rect 1830 178 1836 179
rect 1934 183 1940 184
rect 1934 179 1935 183
rect 1939 179 1940 183
rect 1934 178 1940 179
rect 2030 183 2036 184
rect 2030 179 2031 183
rect 2035 179 2036 183
rect 2030 178 2036 179
rect 2126 183 2132 184
rect 2126 179 2127 183
rect 2131 179 2132 183
rect 2126 178 2132 179
rect 2214 183 2220 184
rect 2214 179 2215 183
rect 2219 179 2220 183
rect 2214 178 2220 179
rect 2302 183 2308 184
rect 2302 179 2303 183
rect 2307 179 2308 183
rect 2302 178 2308 179
rect 2390 183 2396 184
rect 2390 179 2391 183
rect 2395 179 2396 183
rect 2390 178 2396 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2454 178 2460 179
rect 1408 139 1410 178
rect 1512 139 1514 178
rect 1616 139 1618 178
rect 1728 139 1730 178
rect 1832 139 1834 178
rect 1936 139 1938 178
rect 2032 139 2034 178
rect 2128 139 2130 178
rect 2216 139 2218 178
rect 2304 139 2306 178
rect 2392 139 2394 178
rect 2456 139 2458 178
rect 2504 139 2506 179
rect 111 138 115 139
rect 111 133 115 134
rect 151 138 155 139
rect 151 133 155 134
rect 175 138 179 139
rect 175 133 179 134
rect 207 138 211 139
rect 207 133 211 134
rect 255 138 259 139
rect 255 133 259 134
rect 263 138 267 139
rect 263 133 267 134
rect 319 138 323 139
rect 319 133 323 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 431 138 435 139
rect 431 133 435 134
rect 487 138 491 139
rect 487 133 491 134
rect 527 138 531 139
rect 527 133 531 134
rect 551 138 555 139
rect 551 133 555 134
rect 623 138 627 139
rect 623 133 627 134
rect 687 138 691 139
rect 687 133 691 134
rect 711 138 715 139
rect 711 133 715 134
rect 751 138 755 139
rect 751 133 755 134
rect 799 138 803 139
rect 799 133 803 134
rect 815 138 819 139
rect 815 133 819 134
rect 879 138 883 139
rect 879 133 883 134
rect 887 138 891 139
rect 887 133 891 134
rect 943 138 947 139
rect 943 133 947 134
rect 975 138 979 139
rect 975 133 979 134
rect 1007 138 1011 139
rect 1007 133 1011 134
rect 1063 138 1067 139
rect 1063 133 1067 134
rect 1071 138 1075 139
rect 1071 133 1075 134
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1151 138 1155 139
rect 1151 133 1155 134
rect 1199 138 1203 139
rect 1199 133 1203 134
rect 1287 138 1291 139
rect 1287 133 1291 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1367 138 1371 139
rect 1367 133 1371 134
rect 1407 138 1411 139
rect 1407 133 1411 134
rect 1423 138 1427 139
rect 1423 133 1427 134
rect 1479 138 1483 139
rect 1479 133 1483 134
rect 1511 138 1515 139
rect 1511 133 1515 134
rect 1535 138 1539 139
rect 1535 133 1539 134
rect 1591 138 1595 139
rect 1591 133 1595 134
rect 1615 138 1619 139
rect 1615 133 1619 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1703 138 1707 139
rect 1703 133 1707 134
rect 1727 138 1731 139
rect 1727 133 1731 134
rect 1759 138 1763 139
rect 1759 133 1763 134
rect 1815 138 1819 139
rect 1815 133 1819 134
rect 1831 138 1835 139
rect 1831 133 1835 134
rect 1871 138 1875 139
rect 1871 133 1875 134
rect 1927 138 1931 139
rect 1927 133 1931 134
rect 1935 138 1939 139
rect 1935 133 1939 134
rect 1983 138 1987 139
rect 1983 133 1987 134
rect 2031 138 2035 139
rect 2031 133 2035 134
rect 2039 138 2043 139
rect 2039 133 2043 134
rect 2095 138 2099 139
rect 2095 133 2099 134
rect 2127 138 2131 139
rect 2127 133 2131 134
rect 2159 138 2163 139
rect 2159 133 2163 134
rect 2215 138 2219 139
rect 2215 133 2219 134
rect 2223 138 2227 139
rect 2223 133 2227 134
rect 2287 138 2291 139
rect 2287 133 2291 134
rect 2303 138 2307 139
rect 2303 133 2307 134
rect 2343 138 2347 139
rect 2343 133 2347 134
rect 2391 138 2395 139
rect 2391 133 2395 134
rect 2399 138 2403 139
rect 2399 133 2403 134
rect 2455 138 2459 139
rect 2455 133 2459 134
rect 2503 138 2507 139
rect 2503 133 2507 134
rect 112 113 114 133
rect 152 114 154 133
rect 208 114 210 133
rect 264 114 266 133
rect 320 114 322 133
rect 376 114 378 133
rect 432 114 434 133
rect 488 114 490 133
rect 552 114 554 133
rect 624 114 626 133
rect 688 114 690 133
rect 752 114 754 133
rect 816 114 818 133
rect 880 114 882 133
rect 944 114 946 133
rect 1008 114 1010 133
rect 1072 114 1074 133
rect 1136 114 1138 133
rect 1200 114 1202 133
rect 150 113 156 114
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 150 109 151 113
rect 155 109 156 113
rect 150 108 156 109
rect 206 113 212 114
rect 206 109 207 113
rect 211 109 212 113
rect 206 108 212 109
rect 262 113 268 114
rect 262 109 263 113
rect 267 109 268 113
rect 262 108 268 109
rect 318 113 324 114
rect 318 109 319 113
rect 323 109 324 113
rect 318 108 324 109
rect 374 113 380 114
rect 374 109 375 113
rect 379 109 380 113
rect 374 108 380 109
rect 430 113 436 114
rect 430 109 431 113
rect 435 109 436 113
rect 430 108 436 109
rect 486 113 492 114
rect 486 109 487 113
rect 491 109 492 113
rect 486 108 492 109
rect 550 113 556 114
rect 550 109 551 113
rect 555 109 556 113
rect 550 108 556 109
rect 622 113 628 114
rect 622 109 623 113
rect 627 109 628 113
rect 622 108 628 109
rect 686 113 692 114
rect 686 109 687 113
rect 691 109 692 113
rect 686 108 692 109
rect 750 113 756 114
rect 750 109 751 113
rect 755 109 756 113
rect 750 108 756 109
rect 814 113 820 114
rect 814 109 815 113
rect 819 109 820 113
rect 814 108 820 109
rect 878 113 884 114
rect 878 109 879 113
rect 883 109 884 113
rect 878 108 884 109
rect 942 113 948 114
rect 942 109 943 113
rect 947 109 948 113
rect 942 108 948 109
rect 1006 113 1012 114
rect 1006 109 1007 113
rect 1011 109 1012 113
rect 1006 108 1012 109
rect 1070 113 1076 114
rect 1070 109 1071 113
rect 1075 109 1076 113
rect 1070 108 1076 109
rect 1134 113 1140 114
rect 1134 109 1135 113
rect 1139 109 1140 113
rect 1134 108 1140 109
rect 1198 113 1204 114
rect 1288 113 1290 133
rect 1328 113 1330 133
rect 1368 114 1370 133
rect 1424 114 1426 133
rect 1480 114 1482 133
rect 1536 114 1538 133
rect 1592 114 1594 133
rect 1648 114 1650 133
rect 1704 114 1706 133
rect 1760 114 1762 133
rect 1816 114 1818 133
rect 1872 114 1874 133
rect 1928 114 1930 133
rect 1984 114 1986 133
rect 2040 114 2042 133
rect 2096 114 2098 133
rect 2160 114 2162 133
rect 2224 114 2226 133
rect 2288 114 2290 133
rect 2344 114 2346 133
rect 2400 114 2402 133
rect 2456 114 2458 133
rect 1366 113 1372 114
rect 1198 109 1199 113
rect 1203 109 1204 113
rect 1198 108 1204 109
rect 1286 112 1292 113
rect 1286 108 1287 112
rect 1291 108 1292 112
rect 110 107 116 108
rect 1286 107 1292 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1814 113 1820 114
rect 1814 109 1815 113
rect 1819 109 1820 113
rect 1814 108 1820 109
rect 1870 113 1876 114
rect 1870 109 1871 113
rect 1875 109 1876 113
rect 1870 108 1876 109
rect 1926 113 1932 114
rect 1926 109 1927 113
rect 1931 109 1932 113
rect 1926 108 1932 109
rect 1982 113 1988 114
rect 1982 109 1983 113
rect 1987 109 1988 113
rect 1982 108 1988 109
rect 2038 113 2044 114
rect 2038 109 2039 113
rect 2043 109 2044 113
rect 2038 108 2044 109
rect 2094 113 2100 114
rect 2094 109 2095 113
rect 2099 109 2100 113
rect 2094 108 2100 109
rect 2158 113 2164 114
rect 2158 109 2159 113
rect 2163 109 2164 113
rect 2158 108 2164 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2286 113 2292 114
rect 2286 109 2287 113
rect 2291 109 2292 113
rect 2286 108 2292 109
rect 2342 113 2348 114
rect 2342 109 2343 113
rect 2347 109 2348 113
rect 2342 108 2348 109
rect 2398 113 2404 114
rect 2398 109 2399 113
rect 2403 109 2404 113
rect 2398 108 2404 109
rect 2454 113 2460 114
rect 2504 113 2506 133
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 1326 107 1332 108
rect 2502 107 2508 108
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1286 95 1292 96
rect 110 90 116 91
rect 134 92 140 93
rect 112 87 114 90
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 246 92 252 93
rect 246 88 247 92
rect 251 88 252 92
rect 246 87 252 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 358 92 364 93
rect 358 88 359 92
rect 363 88 364 92
rect 358 87 364 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 606 92 612 93
rect 606 88 607 92
rect 611 88 612 92
rect 606 87 612 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 798 92 804 93
rect 798 88 799 92
rect 803 88 804 92
rect 798 87 804 88
rect 862 92 868 93
rect 862 88 863 92
rect 867 88 868 92
rect 862 87 868 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1054 92 1060 93
rect 1054 88 1055 92
rect 1059 88 1060 92
rect 1054 87 1060 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1182 92 1188 93
rect 1182 88 1183 92
rect 1187 88 1188 92
rect 1286 91 1287 95
rect 1291 91 1292 95
rect 1286 90 1292 91
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1182 87 1188 88
rect 1288 87 1290 90
rect 1328 87 1330 90
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1798 92 1804 93
rect 1798 88 1799 92
rect 1803 88 1804 92
rect 1798 87 1804 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1910 92 1916 93
rect 1910 88 1911 92
rect 1915 88 1916 92
rect 1910 87 1916 88
rect 1966 92 1972 93
rect 1966 88 1967 92
rect 1971 88 1972 92
rect 1966 87 1972 88
rect 2022 92 2028 93
rect 2022 88 2023 92
rect 2027 88 2028 92
rect 2022 87 2028 88
rect 2078 92 2084 93
rect 2078 88 2079 92
rect 2083 88 2084 92
rect 2078 87 2084 88
rect 2142 92 2148 93
rect 2142 88 2143 92
rect 2147 88 2148 92
rect 2142 87 2148 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2270 92 2276 93
rect 2270 88 2271 92
rect 2275 88 2276 92
rect 2270 87 2276 88
rect 2326 92 2332 93
rect 2326 88 2327 92
rect 2331 88 2332 92
rect 2326 87 2332 88
rect 2382 92 2388 93
rect 2382 88 2383 92
rect 2387 88 2388 92
rect 2382 87 2388 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
rect 2504 87 2506 90
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 191 86 195 87
rect 191 81 195 82
rect 247 86 251 87
rect 247 81 251 82
rect 303 86 307 87
rect 303 81 307 82
rect 359 86 363 87
rect 359 81 363 82
rect 415 86 419 87
rect 415 81 419 82
rect 471 86 475 87
rect 471 81 475 82
rect 535 86 539 87
rect 535 81 539 82
rect 607 86 611 87
rect 607 81 611 82
rect 671 86 675 87
rect 671 81 675 82
rect 735 86 739 87
rect 735 81 739 82
rect 799 86 803 87
rect 799 81 803 82
rect 863 86 867 87
rect 863 81 867 82
rect 927 86 931 87
rect 927 81 931 82
rect 991 86 995 87
rect 991 81 995 82
rect 1055 86 1059 87
rect 1055 81 1059 82
rect 1119 86 1123 87
rect 1119 81 1123 82
rect 1183 86 1187 87
rect 1183 81 1187 82
rect 1287 86 1291 87
rect 1287 81 1291 82
rect 1327 86 1331 87
rect 1327 81 1331 82
rect 1351 86 1355 87
rect 1351 81 1355 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1463 86 1467 87
rect 1463 81 1467 82
rect 1519 86 1523 87
rect 1519 81 1523 82
rect 1575 86 1579 87
rect 1575 81 1579 82
rect 1631 86 1635 87
rect 1631 81 1635 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1799 86 1803 87
rect 1799 81 1803 82
rect 1855 86 1859 87
rect 1855 81 1859 82
rect 1911 86 1915 87
rect 1911 81 1915 82
rect 1967 86 1971 87
rect 1967 81 1971 82
rect 2023 86 2027 87
rect 2023 81 2027 82
rect 2079 86 2083 87
rect 2079 81 2083 82
rect 2143 86 2147 87
rect 2143 81 2147 82
rect 2207 86 2211 87
rect 2207 81 2211 82
rect 2271 86 2275 87
rect 2271 81 2275 82
rect 2327 86 2331 87
rect 2327 81 2331 82
rect 2383 86 2387 87
rect 2383 81 2387 82
rect 2439 86 2443 87
rect 2439 81 2443 82
rect 2503 86 2507 87
rect 2503 81 2507 82
<< m4c >>
rect 111 2578 115 2582
rect 719 2578 723 2582
rect 775 2578 779 2582
rect 831 2578 835 2582
rect 887 2578 891 2582
rect 943 2578 947 2582
rect 1287 2578 1291 2582
rect 1327 2554 1331 2558
rect 1399 2554 1403 2558
rect 1455 2554 1459 2558
rect 1511 2554 1515 2558
rect 1567 2554 1571 2558
rect 1623 2554 1627 2558
rect 1679 2554 1683 2558
rect 1735 2554 1739 2558
rect 1791 2554 1795 2558
rect 1847 2554 1851 2558
rect 1903 2554 1907 2558
rect 1959 2554 1963 2558
rect 2015 2554 2019 2558
rect 2071 2554 2075 2558
rect 2127 2554 2131 2558
rect 2183 2554 2187 2558
rect 2503 2554 2507 2558
rect 111 2526 115 2530
rect 167 2526 171 2530
rect 223 2526 227 2530
rect 279 2526 283 2530
rect 343 2526 347 2530
rect 407 2526 411 2530
rect 479 2526 483 2530
rect 559 2526 563 2530
rect 639 2526 643 2530
rect 703 2526 707 2530
rect 719 2526 723 2530
rect 759 2526 763 2530
rect 799 2526 803 2530
rect 815 2526 819 2530
rect 871 2526 875 2530
rect 879 2526 883 2530
rect 927 2526 931 2530
rect 959 2526 963 2530
rect 1039 2526 1043 2530
rect 1287 2526 1291 2530
rect 1327 2494 1331 2498
rect 1351 2494 1355 2498
rect 1383 2494 1387 2498
rect 1423 2494 1427 2498
rect 1439 2494 1443 2498
rect 1495 2494 1499 2498
rect 1511 2494 1515 2498
rect 1551 2494 1555 2498
rect 1599 2494 1603 2498
rect 1607 2494 1611 2498
rect 1663 2494 1667 2498
rect 1687 2494 1691 2498
rect 1719 2494 1723 2498
rect 1775 2494 1779 2498
rect 1831 2494 1835 2498
rect 1863 2494 1867 2498
rect 1887 2494 1891 2498
rect 1943 2494 1947 2498
rect 1951 2494 1955 2498
rect 1999 2494 2003 2498
rect 2039 2494 2043 2498
rect 2055 2494 2059 2498
rect 2111 2494 2115 2498
rect 2127 2494 2131 2498
rect 2167 2494 2171 2498
rect 2503 2494 2507 2498
rect 111 2474 115 2478
rect 183 2474 187 2478
rect 239 2474 243 2478
rect 247 2474 251 2478
rect 295 2474 299 2478
rect 327 2474 331 2478
rect 359 2474 363 2478
rect 415 2474 419 2478
rect 423 2474 427 2478
rect 495 2474 499 2478
rect 503 2474 507 2478
rect 575 2474 579 2478
rect 599 2474 603 2478
rect 655 2474 659 2478
rect 695 2474 699 2478
rect 735 2474 739 2478
rect 791 2474 795 2478
rect 815 2474 819 2478
rect 879 2474 883 2478
rect 895 2474 899 2478
rect 967 2474 971 2478
rect 975 2474 979 2478
rect 1055 2474 1059 2478
rect 1063 2474 1067 2478
rect 1159 2474 1163 2478
rect 1287 2474 1291 2478
rect 1327 2434 1331 2438
rect 1367 2434 1371 2438
rect 1439 2434 1443 2438
rect 1527 2434 1531 2438
rect 1543 2434 1547 2438
rect 1615 2434 1619 2438
rect 1639 2434 1643 2438
rect 1703 2434 1707 2438
rect 1735 2434 1739 2438
rect 1791 2434 1795 2438
rect 1823 2434 1827 2438
rect 1879 2434 1883 2438
rect 1911 2434 1915 2438
rect 1967 2434 1971 2438
rect 2007 2434 2011 2438
rect 2055 2434 2059 2438
rect 2103 2434 2107 2438
rect 2143 2434 2147 2438
rect 2503 2434 2507 2438
rect 111 2418 115 2422
rect 151 2418 155 2422
rect 167 2418 171 2422
rect 231 2418 235 2422
rect 311 2418 315 2422
rect 319 2418 323 2422
rect 399 2418 403 2422
rect 415 2418 419 2422
rect 487 2418 491 2422
rect 519 2418 523 2422
rect 583 2418 587 2422
rect 623 2418 627 2422
rect 679 2418 683 2422
rect 727 2418 731 2422
rect 775 2418 779 2422
rect 831 2418 835 2422
rect 863 2418 867 2422
rect 935 2418 939 2422
rect 951 2418 955 2422
rect 1039 2418 1043 2422
rect 1047 2418 1051 2422
rect 1143 2418 1147 2422
rect 1151 2418 1155 2422
rect 1287 2418 1291 2422
rect 1327 2374 1331 2378
rect 1351 2374 1355 2378
rect 1407 2374 1411 2378
rect 1423 2374 1427 2378
rect 1495 2374 1499 2378
rect 1527 2374 1531 2378
rect 1583 2374 1587 2378
rect 1623 2374 1627 2378
rect 1671 2374 1675 2378
rect 1719 2374 1723 2378
rect 1751 2374 1755 2378
rect 1807 2374 1811 2378
rect 1831 2374 1835 2378
rect 1895 2374 1899 2378
rect 1919 2374 1923 2378
rect 1991 2374 1995 2378
rect 2007 2374 2011 2378
rect 2087 2374 2091 2378
rect 2095 2374 2099 2378
rect 2503 2374 2507 2378
rect 111 2366 115 2370
rect 167 2366 171 2370
rect 175 2366 179 2370
rect 247 2366 251 2370
rect 279 2366 283 2370
rect 335 2366 339 2370
rect 391 2366 395 2370
rect 431 2366 435 2370
rect 503 2366 507 2370
rect 535 2366 539 2370
rect 623 2366 627 2370
rect 639 2366 643 2370
rect 743 2366 747 2370
rect 847 2366 851 2370
rect 871 2366 875 2370
rect 951 2366 955 2370
rect 999 2366 1003 2370
rect 1055 2366 1059 2370
rect 1127 2366 1131 2370
rect 1167 2366 1171 2370
rect 1287 2366 1291 2370
rect 1327 2318 1331 2322
rect 1367 2318 1371 2322
rect 1423 2318 1427 2322
rect 1455 2318 1459 2322
rect 1511 2318 1515 2322
rect 1543 2318 1547 2322
rect 1599 2318 1603 2322
rect 1639 2318 1643 2322
rect 1687 2318 1691 2322
rect 1735 2318 1739 2322
rect 1767 2318 1771 2322
rect 1831 2318 1835 2322
rect 1847 2318 1851 2322
rect 1927 2318 1931 2322
rect 1935 2318 1939 2322
rect 2015 2318 2019 2322
rect 2023 2318 2027 2322
rect 2111 2318 2115 2322
rect 2207 2318 2211 2322
rect 2503 2318 2507 2322
rect 111 2310 115 2314
rect 159 2310 163 2314
rect 207 2310 211 2314
rect 263 2310 267 2314
rect 287 2310 291 2314
rect 375 2310 379 2314
rect 471 2310 475 2314
rect 487 2310 491 2314
rect 559 2310 563 2314
rect 607 2310 611 2314
rect 647 2310 651 2314
rect 727 2310 731 2314
rect 735 2310 739 2314
rect 815 2310 819 2314
rect 855 2310 859 2314
rect 903 2310 907 2314
rect 983 2310 987 2314
rect 991 2310 995 2314
rect 1079 2310 1083 2314
rect 1111 2310 1115 2314
rect 1287 2310 1291 2314
rect 1327 2266 1331 2270
rect 1351 2266 1355 2270
rect 1439 2266 1443 2270
rect 1455 2266 1459 2270
rect 1527 2266 1531 2270
rect 1543 2266 1547 2270
rect 1623 2266 1627 2270
rect 1639 2266 1643 2270
rect 1719 2266 1723 2270
rect 1735 2266 1739 2270
rect 1815 2266 1819 2270
rect 1839 2266 1843 2270
rect 1911 2266 1915 2270
rect 1935 2266 1939 2270
rect 1999 2266 2003 2270
rect 2031 2266 2035 2270
rect 2095 2266 2099 2270
rect 2119 2266 2123 2270
rect 2191 2266 2195 2270
rect 2215 2266 2219 2270
rect 2311 2266 2315 2270
rect 2503 2266 2507 2270
rect 111 2254 115 2258
rect 223 2254 227 2258
rect 263 2254 267 2258
rect 303 2254 307 2258
rect 319 2254 323 2258
rect 383 2254 387 2258
rect 391 2254 395 2258
rect 447 2254 451 2258
rect 487 2254 491 2258
rect 503 2254 507 2258
rect 559 2254 563 2258
rect 575 2254 579 2258
rect 615 2254 619 2258
rect 663 2254 667 2258
rect 671 2254 675 2258
rect 727 2254 731 2258
rect 751 2254 755 2258
rect 791 2254 795 2258
rect 831 2254 835 2258
rect 855 2254 859 2258
rect 919 2254 923 2258
rect 983 2254 987 2258
rect 1007 2254 1011 2258
rect 1047 2254 1051 2258
rect 1095 2254 1099 2258
rect 1111 2254 1115 2258
rect 1287 2254 1291 2258
rect 1327 2210 1331 2214
rect 1471 2210 1475 2214
rect 1559 2210 1563 2214
rect 1567 2210 1571 2214
rect 1623 2210 1627 2214
rect 1655 2210 1659 2214
rect 1679 2210 1683 2214
rect 1743 2210 1747 2214
rect 1751 2210 1755 2214
rect 1807 2210 1811 2214
rect 1855 2210 1859 2214
rect 1871 2210 1875 2214
rect 1927 2210 1931 2214
rect 1951 2210 1955 2214
rect 1983 2210 1987 2214
rect 2039 2210 2043 2214
rect 2047 2210 2051 2214
rect 2095 2210 2099 2214
rect 2135 2210 2139 2214
rect 2159 2210 2163 2214
rect 2223 2210 2227 2214
rect 2231 2210 2235 2214
rect 2287 2210 2291 2214
rect 2327 2210 2331 2214
rect 2343 2210 2347 2214
rect 2399 2210 2403 2214
rect 2455 2210 2459 2214
rect 2503 2210 2507 2214
rect 111 2198 115 2202
rect 247 2198 251 2202
rect 303 2198 307 2202
rect 335 2198 339 2202
rect 367 2198 371 2202
rect 391 2198 395 2202
rect 431 2198 435 2202
rect 447 2198 451 2202
rect 487 2198 491 2202
rect 503 2198 507 2202
rect 543 2198 547 2202
rect 559 2198 563 2202
rect 599 2198 603 2202
rect 655 2198 659 2202
rect 711 2198 715 2202
rect 775 2198 779 2202
rect 839 2198 843 2202
rect 903 2198 907 2202
rect 967 2198 971 2202
rect 1031 2198 1035 2202
rect 1095 2198 1099 2202
rect 1287 2198 1291 2202
rect 111 2146 115 2150
rect 351 2146 355 2150
rect 407 2146 411 2150
rect 415 2146 419 2150
rect 463 2146 467 2150
rect 511 2146 515 2150
rect 519 2146 523 2150
rect 575 2146 579 2150
rect 607 2146 611 2150
rect 711 2146 715 2150
rect 815 2146 819 2150
rect 927 2146 931 2150
rect 1039 2146 1043 2150
rect 1151 2146 1155 2150
rect 1239 2146 1243 2150
rect 1287 2146 1291 2150
rect 1327 2146 1331 2150
rect 1551 2146 1555 2150
rect 1607 2146 1611 2150
rect 1663 2146 1667 2150
rect 1719 2146 1723 2150
rect 1727 2146 1731 2150
rect 1791 2146 1795 2150
rect 1855 2146 1859 2150
rect 1871 2146 1875 2150
rect 1911 2146 1915 2150
rect 1967 2146 1971 2150
rect 2023 2146 2027 2150
rect 2079 2146 2083 2150
rect 2143 2146 2147 2150
rect 2199 2146 2203 2150
rect 2207 2146 2211 2150
rect 2271 2146 2275 2150
rect 2327 2146 2331 2150
rect 2383 2146 2387 2150
rect 2439 2146 2443 2150
rect 2503 2146 2507 2150
rect 111 2094 115 2098
rect 375 2094 379 2098
rect 399 2094 403 2098
rect 447 2094 451 2098
rect 495 2094 499 2098
rect 519 2094 523 2098
rect 591 2094 595 2098
rect 599 2094 603 2098
rect 679 2094 683 2098
rect 695 2094 699 2098
rect 759 2094 763 2098
rect 799 2094 803 2098
rect 831 2094 835 2098
rect 903 2094 907 2098
rect 911 2094 915 2098
rect 967 2094 971 2098
rect 1023 2094 1027 2098
rect 1031 2094 1035 2098
rect 1103 2094 1107 2098
rect 1135 2094 1139 2098
rect 1167 2094 1171 2098
rect 1223 2094 1227 2098
rect 1287 2094 1291 2098
rect 1327 2082 1331 2086
rect 1367 2082 1371 2086
rect 1423 2082 1427 2086
rect 1503 2082 1507 2086
rect 1591 2082 1595 2086
rect 1679 2082 1683 2086
rect 1735 2082 1739 2086
rect 1783 2082 1787 2086
rect 1807 2082 1811 2086
rect 1887 2082 1891 2086
rect 1895 2082 1899 2086
rect 1983 2082 1987 2086
rect 2023 2082 2027 2086
rect 2095 2082 2099 2086
rect 2167 2082 2171 2086
rect 2215 2082 2219 2086
rect 2319 2082 2323 2086
rect 2343 2082 2347 2086
rect 2455 2082 2459 2086
rect 2503 2082 2507 2086
rect 111 2038 115 2042
rect 295 2038 299 2042
rect 375 2038 379 2042
rect 391 2038 395 2042
rect 463 2038 467 2042
rect 535 2038 539 2042
rect 551 2038 555 2042
rect 615 2038 619 2042
rect 639 2038 643 2042
rect 695 2038 699 2042
rect 719 2038 723 2042
rect 775 2038 779 2042
rect 799 2038 803 2042
rect 847 2038 851 2042
rect 887 2038 891 2042
rect 919 2038 923 2042
rect 975 2038 979 2042
rect 983 2038 987 2042
rect 1047 2038 1051 2042
rect 1063 2038 1067 2042
rect 1119 2038 1123 2042
rect 1183 2038 1187 2042
rect 1239 2038 1243 2042
rect 1287 2038 1291 2042
rect 1327 2030 1331 2034
rect 1351 2030 1355 2034
rect 1407 2030 1411 2034
rect 1423 2030 1427 2034
rect 1487 2030 1491 2034
rect 1519 2030 1523 2034
rect 1575 2030 1579 2034
rect 1615 2030 1619 2034
rect 1663 2030 1667 2034
rect 1719 2030 1723 2034
rect 1767 2030 1771 2034
rect 1823 2030 1827 2034
rect 1879 2030 1883 2034
rect 1935 2030 1939 2034
rect 2007 2030 2011 2034
rect 2055 2030 2059 2034
rect 2151 2030 2155 2034
rect 2183 2030 2187 2034
rect 2303 2030 2307 2034
rect 2319 2030 2323 2034
rect 2439 2030 2443 2034
rect 2503 2030 2507 2034
rect 111 1982 115 1986
rect 135 1982 139 1986
rect 207 1982 211 1986
rect 279 1982 283 1986
rect 287 1982 291 1986
rect 359 1982 363 1986
rect 383 1982 387 1986
rect 447 1982 451 1986
rect 487 1982 491 1986
rect 535 1982 539 1986
rect 591 1982 595 1986
rect 623 1982 627 1986
rect 695 1982 699 1986
rect 703 1982 707 1986
rect 783 1982 787 1986
rect 799 1982 803 1986
rect 871 1982 875 1986
rect 903 1982 907 1986
rect 959 1982 963 1986
rect 1015 1982 1019 1986
rect 1047 1982 1051 1986
rect 1287 1982 1291 1986
rect 1327 1974 1331 1978
rect 1367 1974 1371 1978
rect 1439 1974 1443 1978
rect 1455 1974 1459 1978
rect 1535 1974 1539 1978
rect 1543 1974 1547 1978
rect 1631 1974 1635 1978
rect 1639 1974 1643 1978
rect 1735 1974 1739 1978
rect 1839 1974 1843 1978
rect 1943 1974 1947 1978
rect 1951 1974 1955 1978
rect 2047 1974 2051 1978
rect 2071 1974 2075 1978
rect 2151 1974 2155 1978
rect 2199 1974 2203 1978
rect 2255 1974 2259 1978
rect 2335 1974 2339 1978
rect 2367 1974 2371 1978
rect 2455 1974 2459 1978
rect 2503 1974 2507 1978
rect 111 1922 115 1926
rect 151 1922 155 1926
rect 223 1922 227 1926
rect 239 1922 243 1926
rect 303 1922 307 1926
rect 375 1922 379 1926
rect 399 1922 403 1926
rect 503 1922 507 1926
rect 527 1922 531 1926
rect 607 1922 611 1926
rect 687 1922 691 1926
rect 711 1922 715 1926
rect 815 1922 819 1926
rect 863 1922 867 1926
rect 919 1922 923 1926
rect 1031 1922 1035 1926
rect 1039 1922 1043 1926
rect 1287 1922 1291 1926
rect 1327 1918 1331 1922
rect 1439 1918 1443 1922
rect 1527 1918 1531 1922
rect 1615 1918 1619 1922
rect 1623 1918 1627 1922
rect 1711 1918 1715 1922
rect 1719 1918 1723 1922
rect 1815 1918 1819 1922
rect 1823 1918 1827 1922
rect 1919 1918 1923 1922
rect 1927 1918 1931 1922
rect 2015 1918 2019 1922
rect 2031 1918 2035 1922
rect 2111 1918 2115 1922
rect 2135 1918 2139 1922
rect 2199 1918 2203 1922
rect 2239 1918 2243 1922
rect 2287 1918 2291 1922
rect 2351 1918 2355 1922
rect 2375 1918 2379 1922
rect 2439 1918 2443 1922
rect 2503 1918 2507 1922
rect 111 1870 115 1874
rect 135 1870 139 1874
rect 191 1870 195 1874
rect 223 1870 227 1874
rect 263 1870 267 1874
rect 335 1870 339 1874
rect 359 1870 363 1874
rect 407 1870 411 1874
rect 479 1870 483 1874
rect 511 1870 515 1874
rect 551 1870 555 1874
rect 615 1870 619 1874
rect 671 1870 675 1874
rect 679 1870 683 1874
rect 743 1870 747 1874
rect 815 1870 819 1874
rect 847 1870 851 1874
rect 887 1870 891 1874
rect 959 1870 963 1874
rect 1023 1870 1027 1874
rect 1039 1870 1043 1874
rect 1287 1870 1291 1874
rect 1327 1866 1331 1870
rect 1535 1866 1539 1870
rect 1543 1866 1547 1870
rect 1607 1866 1611 1870
rect 1631 1866 1635 1870
rect 1687 1866 1691 1870
rect 1727 1866 1731 1870
rect 1783 1866 1787 1870
rect 1831 1866 1835 1870
rect 1879 1866 1883 1870
rect 1935 1866 1939 1870
rect 1983 1866 1987 1870
rect 2031 1866 2035 1870
rect 2079 1866 2083 1870
rect 2127 1866 2131 1870
rect 2175 1866 2179 1870
rect 2215 1866 2219 1870
rect 2271 1866 2275 1870
rect 2303 1866 2307 1870
rect 2367 1866 2371 1870
rect 2391 1866 2395 1870
rect 2455 1866 2459 1870
rect 2503 1866 2507 1870
rect 111 1810 115 1814
rect 151 1810 155 1814
rect 207 1810 211 1814
rect 231 1810 235 1814
rect 279 1810 283 1814
rect 335 1810 339 1814
rect 351 1810 355 1814
rect 423 1810 427 1814
rect 439 1810 443 1814
rect 495 1810 499 1814
rect 535 1810 539 1814
rect 567 1810 571 1814
rect 631 1810 635 1814
rect 695 1810 699 1814
rect 719 1810 723 1814
rect 759 1810 763 1814
rect 799 1810 803 1814
rect 831 1810 835 1814
rect 879 1810 883 1814
rect 903 1810 907 1814
rect 959 1810 963 1814
rect 975 1810 979 1814
rect 1039 1810 1043 1814
rect 1055 1810 1059 1814
rect 1119 1810 1123 1814
rect 1287 1810 1291 1814
rect 1327 1810 1331 1814
rect 1463 1810 1467 1814
rect 1519 1810 1523 1814
rect 1559 1810 1563 1814
rect 1591 1810 1595 1814
rect 1663 1810 1667 1814
rect 1671 1810 1675 1814
rect 1767 1810 1771 1814
rect 1863 1810 1867 1814
rect 1879 1810 1883 1814
rect 1967 1810 1971 1814
rect 1983 1810 1987 1814
rect 2063 1810 2067 1814
rect 2087 1810 2091 1814
rect 2159 1810 2163 1814
rect 2183 1810 2187 1814
rect 2255 1810 2259 1814
rect 2271 1810 2275 1814
rect 2351 1810 2355 1814
rect 2367 1810 2371 1814
rect 2439 1810 2443 1814
rect 2503 1810 2507 1814
rect 111 1754 115 1758
rect 135 1754 139 1758
rect 215 1754 219 1758
rect 239 1754 243 1758
rect 319 1754 323 1758
rect 351 1754 355 1758
rect 423 1754 427 1758
rect 463 1754 467 1758
rect 519 1754 523 1758
rect 575 1754 579 1758
rect 615 1754 619 1758
rect 679 1754 683 1758
rect 703 1754 707 1758
rect 783 1754 787 1758
rect 863 1754 867 1758
rect 887 1754 891 1758
rect 943 1754 947 1758
rect 991 1754 995 1758
rect 1023 1754 1027 1758
rect 1103 1754 1107 1758
rect 1287 1754 1291 1758
rect 1327 1754 1331 1758
rect 1375 1754 1379 1758
rect 1471 1754 1475 1758
rect 1479 1754 1483 1758
rect 1567 1754 1571 1758
rect 1575 1754 1579 1758
rect 1671 1754 1675 1758
rect 1679 1754 1683 1758
rect 1775 1754 1779 1758
rect 1783 1754 1787 1758
rect 1887 1754 1891 1758
rect 1895 1754 1899 1758
rect 1999 1754 2003 1758
rect 2103 1754 2107 1758
rect 2111 1754 2115 1758
rect 2199 1754 2203 1758
rect 2231 1754 2235 1758
rect 2287 1754 2291 1758
rect 2351 1754 2355 1758
rect 2383 1754 2387 1758
rect 2455 1754 2459 1758
rect 2503 1754 2507 1758
rect 111 1698 115 1702
rect 151 1698 155 1702
rect 191 1698 195 1702
rect 255 1698 259 1702
rect 271 1698 275 1702
rect 351 1698 355 1702
rect 367 1698 371 1702
rect 439 1698 443 1702
rect 479 1698 483 1702
rect 535 1698 539 1702
rect 591 1698 595 1702
rect 639 1698 643 1702
rect 695 1698 699 1702
rect 743 1698 747 1702
rect 799 1698 803 1702
rect 847 1698 851 1702
rect 903 1698 907 1702
rect 951 1698 955 1702
rect 1007 1698 1011 1702
rect 1063 1698 1067 1702
rect 1119 1698 1123 1702
rect 1175 1698 1179 1702
rect 1287 1698 1291 1702
rect 1327 1702 1331 1706
rect 1351 1702 1355 1706
rect 1359 1702 1363 1706
rect 1431 1702 1435 1706
rect 1455 1702 1459 1706
rect 1535 1702 1539 1706
rect 1551 1702 1555 1706
rect 1647 1702 1651 1706
rect 1655 1702 1659 1706
rect 1759 1702 1763 1706
rect 1871 1702 1875 1706
rect 1879 1702 1883 1706
rect 1983 1702 1987 1706
rect 2015 1702 2019 1706
rect 2095 1702 2099 1706
rect 2159 1702 2163 1706
rect 2215 1702 2219 1706
rect 2311 1702 2315 1706
rect 2335 1702 2339 1706
rect 2439 1702 2443 1706
rect 2503 1702 2507 1706
rect 111 1646 115 1650
rect 175 1646 179 1650
rect 215 1646 219 1650
rect 255 1646 259 1650
rect 271 1646 275 1650
rect 335 1646 339 1650
rect 407 1646 411 1650
rect 423 1646 427 1650
rect 479 1646 483 1650
rect 519 1646 523 1650
rect 559 1646 563 1650
rect 623 1646 627 1650
rect 647 1646 651 1650
rect 727 1646 731 1650
rect 743 1646 747 1650
rect 831 1646 835 1650
rect 839 1646 843 1650
rect 935 1646 939 1650
rect 943 1646 947 1650
rect 1047 1646 1051 1650
rect 1055 1646 1059 1650
rect 1159 1646 1163 1650
rect 1175 1646 1179 1650
rect 1287 1646 1291 1650
rect 1327 1642 1331 1646
rect 1367 1642 1371 1646
rect 1431 1642 1435 1646
rect 1447 1642 1451 1646
rect 1519 1642 1523 1646
rect 1551 1642 1555 1646
rect 1599 1642 1603 1646
rect 1663 1642 1667 1646
rect 1679 1642 1683 1646
rect 1751 1642 1755 1646
rect 1775 1642 1779 1646
rect 1839 1642 1843 1646
rect 1895 1642 1899 1646
rect 1935 1642 1939 1646
rect 2031 1642 2035 1646
rect 2055 1642 2059 1646
rect 2175 1642 2179 1646
rect 2183 1642 2187 1646
rect 2327 1642 2331 1646
rect 2455 1642 2459 1646
rect 2503 1642 2507 1646
rect 111 1594 115 1598
rect 231 1594 235 1598
rect 287 1594 291 1598
rect 351 1594 355 1598
rect 423 1594 427 1598
rect 495 1594 499 1598
rect 503 1594 507 1598
rect 575 1594 579 1598
rect 599 1594 603 1598
rect 663 1594 667 1598
rect 703 1594 707 1598
rect 759 1594 763 1598
rect 815 1594 819 1598
rect 855 1594 859 1598
rect 935 1594 939 1598
rect 959 1594 963 1598
rect 1063 1594 1067 1598
rect 1071 1594 1075 1598
rect 1191 1594 1195 1598
rect 1287 1594 1291 1598
rect 1327 1586 1331 1590
rect 1351 1586 1355 1590
rect 1415 1586 1419 1590
rect 1423 1586 1427 1590
rect 1503 1586 1507 1590
rect 1527 1586 1531 1590
rect 1583 1586 1587 1590
rect 1647 1586 1651 1590
rect 1663 1586 1667 1590
rect 1735 1586 1739 1590
rect 1783 1586 1787 1590
rect 1823 1586 1827 1590
rect 1919 1586 1923 1590
rect 1935 1586 1939 1590
rect 2039 1586 2043 1590
rect 2103 1586 2107 1590
rect 2167 1586 2171 1590
rect 2279 1586 2283 1590
rect 2311 1586 2315 1590
rect 2439 1586 2443 1590
rect 2503 1586 2507 1590
rect 111 1534 115 1538
rect 271 1534 275 1538
rect 335 1534 339 1538
rect 407 1534 411 1538
rect 471 1534 475 1538
rect 487 1534 491 1538
rect 551 1534 555 1538
rect 583 1534 587 1538
rect 639 1534 643 1538
rect 687 1534 691 1538
rect 735 1534 739 1538
rect 799 1534 803 1538
rect 839 1534 843 1538
rect 919 1534 923 1538
rect 951 1534 955 1538
rect 1047 1534 1051 1538
rect 1063 1534 1067 1538
rect 1175 1534 1179 1538
rect 1287 1534 1291 1538
rect 1327 1534 1331 1538
rect 1367 1534 1371 1538
rect 1439 1534 1443 1538
rect 1543 1534 1547 1538
rect 1647 1534 1651 1538
rect 1663 1534 1667 1538
rect 1751 1534 1755 1538
rect 1799 1534 1803 1538
rect 1855 1534 1859 1538
rect 1951 1534 1955 1538
rect 1959 1534 1963 1538
rect 2055 1534 2059 1538
rect 2119 1534 2123 1538
rect 2151 1534 2155 1538
rect 2247 1534 2251 1538
rect 2295 1534 2299 1538
rect 2343 1534 2347 1538
rect 2439 1534 2443 1538
rect 2455 1534 2459 1538
rect 2503 1534 2507 1538
rect 111 1482 115 1486
rect 375 1482 379 1486
rect 463 1482 467 1486
rect 487 1482 491 1486
rect 559 1482 563 1486
rect 567 1482 571 1486
rect 655 1482 659 1486
rect 751 1482 755 1486
rect 855 1482 859 1486
rect 959 1482 963 1486
rect 967 1482 971 1486
rect 1063 1482 1067 1486
rect 1079 1482 1083 1486
rect 1167 1482 1171 1486
rect 1191 1482 1195 1486
rect 1287 1482 1291 1486
rect 1327 1478 1331 1482
rect 1351 1478 1355 1482
rect 1423 1478 1427 1482
rect 1519 1478 1523 1482
rect 1527 1478 1531 1482
rect 1615 1478 1619 1482
rect 1631 1478 1635 1482
rect 1711 1478 1715 1482
rect 1735 1478 1739 1482
rect 1815 1478 1819 1482
rect 1839 1478 1843 1482
rect 1927 1478 1931 1482
rect 1943 1478 1947 1482
rect 2039 1478 2043 1482
rect 2047 1478 2051 1482
rect 2135 1478 2139 1482
rect 2175 1478 2179 1482
rect 2231 1478 2235 1482
rect 2303 1478 2307 1482
rect 2327 1478 2331 1482
rect 2423 1478 2427 1482
rect 2439 1478 2443 1482
rect 2503 1478 2507 1482
rect 111 1430 115 1434
rect 231 1430 235 1434
rect 319 1430 323 1434
rect 359 1430 363 1434
rect 415 1430 419 1434
rect 447 1430 451 1434
rect 511 1430 515 1434
rect 543 1430 547 1434
rect 615 1430 619 1434
rect 639 1430 643 1434
rect 711 1430 715 1434
rect 735 1430 739 1434
rect 807 1430 811 1434
rect 839 1430 843 1434
rect 895 1430 899 1434
rect 943 1430 947 1434
rect 991 1430 995 1434
rect 1047 1430 1051 1434
rect 1087 1430 1091 1434
rect 1151 1430 1155 1434
rect 1287 1430 1291 1434
rect 1327 1422 1331 1426
rect 1367 1422 1371 1426
rect 1423 1422 1427 1426
rect 1439 1422 1443 1426
rect 1503 1422 1507 1426
rect 1535 1422 1539 1426
rect 1591 1422 1595 1426
rect 1631 1422 1635 1426
rect 1679 1422 1683 1426
rect 1727 1422 1731 1426
rect 1775 1422 1779 1426
rect 1831 1422 1835 1426
rect 1879 1422 1883 1426
rect 1943 1422 1947 1426
rect 1991 1422 1995 1426
rect 2063 1422 2067 1426
rect 2111 1422 2115 1426
rect 2191 1422 2195 1426
rect 2231 1422 2235 1426
rect 2319 1422 2323 1426
rect 2351 1422 2355 1426
rect 2455 1422 2459 1426
rect 2503 1422 2507 1426
rect 111 1378 115 1382
rect 151 1378 155 1382
rect 215 1378 219 1382
rect 247 1378 251 1382
rect 311 1378 315 1382
rect 335 1378 339 1382
rect 407 1378 411 1382
rect 431 1378 435 1382
rect 511 1378 515 1382
rect 527 1378 531 1382
rect 607 1378 611 1382
rect 631 1378 635 1382
rect 703 1378 707 1382
rect 727 1378 731 1382
rect 799 1378 803 1382
rect 823 1378 827 1382
rect 895 1378 899 1382
rect 911 1378 915 1382
rect 999 1378 1003 1382
rect 1007 1378 1011 1382
rect 1103 1378 1107 1382
rect 1287 1378 1291 1382
rect 1327 1366 1331 1370
rect 1351 1366 1355 1370
rect 1407 1366 1411 1370
rect 1479 1366 1483 1370
rect 1487 1366 1491 1370
rect 1567 1366 1571 1370
rect 1575 1366 1579 1370
rect 1655 1366 1659 1370
rect 1663 1366 1667 1370
rect 1751 1366 1755 1370
rect 1759 1366 1763 1370
rect 1855 1366 1859 1370
rect 1863 1366 1867 1370
rect 1967 1366 1971 1370
rect 1975 1366 1979 1370
rect 2079 1366 2083 1370
rect 2095 1366 2099 1370
rect 2199 1366 2203 1370
rect 2215 1366 2219 1370
rect 2327 1366 2331 1370
rect 2335 1366 2339 1370
rect 2439 1366 2443 1370
rect 2503 1366 2507 1370
rect 111 1326 115 1330
rect 135 1326 139 1330
rect 199 1326 203 1330
rect 215 1326 219 1330
rect 295 1326 299 1330
rect 319 1326 323 1330
rect 391 1326 395 1330
rect 415 1326 419 1330
rect 495 1326 499 1330
rect 511 1326 515 1330
rect 591 1326 595 1330
rect 599 1326 603 1330
rect 687 1326 691 1330
rect 783 1326 787 1330
rect 879 1326 883 1330
rect 983 1326 987 1330
rect 1287 1326 1291 1330
rect 1327 1306 1331 1310
rect 1367 1306 1371 1310
rect 1423 1306 1427 1310
rect 1495 1306 1499 1310
rect 1519 1306 1523 1310
rect 1583 1306 1587 1310
rect 1615 1306 1619 1310
rect 1671 1306 1675 1310
rect 1719 1306 1723 1310
rect 1767 1306 1771 1310
rect 1823 1306 1827 1310
rect 1871 1306 1875 1310
rect 1919 1306 1923 1310
rect 1983 1306 1987 1310
rect 2015 1306 2019 1310
rect 2095 1306 2099 1310
rect 2103 1306 2107 1310
rect 2183 1306 2187 1310
rect 2215 1306 2219 1310
rect 2255 1306 2259 1310
rect 2327 1306 2331 1310
rect 2343 1306 2347 1310
rect 2399 1306 2403 1310
rect 2455 1306 2459 1310
rect 2503 1306 2507 1310
rect 111 1274 115 1278
rect 151 1274 155 1278
rect 191 1274 195 1278
rect 231 1274 235 1278
rect 247 1274 251 1278
rect 303 1274 307 1278
rect 335 1274 339 1278
rect 367 1274 371 1278
rect 431 1274 435 1278
rect 439 1274 443 1278
rect 527 1274 531 1278
rect 615 1274 619 1278
rect 639 1274 643 1278
rect 703 1274 707 1278
rect 775 1274 779 1278
rect 799 1274 803 1278
rect 895 1274 899 1278
rect 927 1274 931 1278
rect 1095 1274 1099 1278
rect 1239 1274 1243 1278
rect 1287 1274 1291 1278
rect 1327 1238 1331 1242
rect 1351 1238 1355 1242
rect 1407 1238 1411 1242
rect 1447 1238 1451 1242
rect 1503 1238 1507 1242
rect 1575 1238 1579 1242
rect 1599 1238 1603 1242
rect 1695 1238 1699 1242
rect 1703 1238 1707 1242
rect 1807 1238 1811 1242
rect 1815 1238 1819 1242
rect 1903 1238 1907 1242
rect 1927 1238 1931 1242
rect 1999 1238 2003 1242
rect 2031 1238 2035 1242
rect 2087 1238 2091 1242
rect 2127 1238 2131 1242
rect 2167 1238 2171 1242
rect 2215 1238 2219 1242
rect 2239 1238 2243 1242
rect 2295 1238 2299 1242
rect 2311 1238 2315 1242
rect 2375 1238 2379 1242
rect 2383 1238 2387 1242
rect 2439 1238 2443 1242
rect 2503 1238 2507 1242
rect 111 1222 115 1226
rect 175 1222 179 1226
rect 231 1222 235 1226
rect 287 1222 291 1226
rect 351 1222 355 1226
rect 407 1222 411 1226
rect 423 1222 427 1226
rect 463 1222 467 1226
rect 511 1222 515 1226
rect 519 1222 523 1226
rect 575 1222 579 1226
rect 623 1222 627 1226
rect 631 1222 635 1226
rect 687 1222 691 1226
rect 743 1222 747 1226
rect 759 1222 763 1226
rect 799 1222 803 1226
rect 855 1222 859 1226
rect 911 1222 915 1226
rect 1079 1222 1083 1226
rect 1223 1222 1227 1226
rect 1287 1222 1291 1226
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1463 1186 1467 1190
rect 1471 1186 1475 1190
rect 1591 1186 1595 1190
rect 1599 1186 1603 1190
rect 1711 1186 1715 1190
rect 1735 1186 1739 1190
rect 1831 1186 1835 1190
rect 1863 1186 1867 1190
rect 1943 1186 1947 1190
rect 1983 1186 1987 1190
rect 2047 1186 2051 1190
rect 2087 1186 2091 1190
rect 2143 1186 2147 1190
rect 2191 1186 2195 1190
rect 2231 1186 2235 1190
rect 2287 1186 2291 1190
rect 2311 1186 2315 1190
rect 2383 1186 2387 1190
rect 2391 1186 2395 1190
rect 2455 1186 2459 1190
rect 2503 1186 2507 1190
rect 111 1166 115 1170
rect 367 1166 371 1170
rect 423 1166 427 1170
rect 479 1166 483 1170
rect 535 1166 539 1170
rect 591 1166 595 1170
rect 647 1166 651 1170
rect 703 1166 707 1170
rect 759 1166 763 1170
rect 815 1166 819 1170
rect 871 1166 875 1170
rect 927 1166 931 1170
rect 983 1166 987 1170
rect 1287 1166 1291 1170
rect 1327 1130 1331 1134
rect 1351 1130 1355 1134
rect 1367 1130 1371 1134
rect 1447 1130 1451 1134
rect 1455 1130 1459 1134
rect 1535 1130 1539 1134
rect 1583 1130 1587 1134
rect 1631 1130 1635 1134
rect 1719 1130 1723 1134
rect 1807 1130 1811 1134
rect 1847 1130 1851 1134
rect 1895 1130 1899 1134
rect 1967 1130 1971 1134
rect 1983 1130 1987 1134
rect 2071 1130 2075 1134
rect 2159 1130 2163 1134
rect 2175 1130 2179 1134
rect 2255 1130 2259 1134
rect 2271 1130 2275 1134
rect 2359 1130 2363 1134
rect 2367 1130 2371 1134
rect 2439 1130 2443 1134
rect 2503 1130 2507 1134
rect 111 1110 115 1114
rect 223 1110 227 1114
rect 311 1110 315 1114
rect 399 1110 403 1114
rect 407 1110 411 1114
rect 463 1110 467 1114
rect 495 1110 499 1114
rect 519 1110 523 1114
rect 575 1110 579 1114
rect 591 1110 595 1114
rect 631 1110 635 1114
rect 679 1110 683 1114
rect 687 1110 691 1114
rect 743 1110 747 1114
rect 767 1110 771 1114
rect 799 1110 803 1114
rect 847 1110 851 1114
rect 855 1110 859 1114
rect 911 1110 915 1114
rect 927 1110 931 1114
rect 967 1110 971 1114
rect 1015 1110 1019 1114
rect 1103 1110 1107 1114
rect 1287 1110 1291 1114
rect 1327 1070 1331 1074
rect 1383 1070 1387 1074
rect 1431 1070 1435 1074
rect 1463 1070 1467 1074
rect 1495 1070 1499 1074
rect 1551 1070 1555 1074
rect 1567 1070 1571 1074
rect 1639 1070 1643 1074
rect 1647 1070 1651 1074
rect 1703 1070 1707 1074
rect 1735 1070 1739 1074
rect 1767 1070 1771 1074
rect 1823 1070 1827 1074
rect 1839 1070 1843 1074
rect 1911 1070 1915 1074
rect 1919 1070 1923 1074
rect 1999 1070 2003 1074
rect 2007 1070 2011 1074
rect 2087 1070 2091 1074
rect 2111 1070 2115 1074
rect 2175 1070 2179 1074
rect 2231 1070 2235 1074
rect 2271 1070 2275 1074
rect 2351 1070 2355 1074
rect 2375 1070 2379 1074
rect 2455 1070 2459 1074
rect 2503 1070 2507 1074
rect 111 1054 115 1058
rect 151 1054 155 1058
rect 207 1054 211 1058
rect 239 1054 243 1058
rect 303 1054 307 1058
rect 327 1054 331 1058
rect 415 1054 419 1058
rect 511 1054 515 1058
rect 535 1054 539 1058
rect 607 1054 611 1058
rect 655 1054 659 1058
rect 695 1054 699 1058
rect 767 1054 771 1058
rect 783 1054 787 1058
rect 863 1054 867 1058
rect 879 1054 883 1058
rect 943 1054 947 1058
rect 983 1054 987 1058
rect 1031 1054 1035 1058
rect 1095 1054 1099 1058
rect 1119 1054 1123 1058
rect 1207 1054 1211 1058
rect 1287 1054 1291 1058
rect 1327 1010 1331 1014
rect 1415 1010 1419 1014
rect 1479 1010 1483 1014
rect 1511 1010 1515 1014
rect 1551 1010 1555 1014
rect 1567 1010 1571 1014
rect 1623 1010 1627 1014
rect 1679 1010 1683 1014
rect 1687 1010 1691 1014
rect 1735 1010 1739 1014
rect 1751 1010 1755 1014
rect 1807 1010 1811 1014
rect 1823 1010 1827 1014
rect 1887 1010 1891 1014
rect 1903 1010 1907 1014
rect 1983 1010 1987 1014
rect 1991 1010 1995 1014
rect 2095 1010 2099 1014
rect 2215 1010 2219 1014
rect 2335 1010 2339 1014
rect 2439 1010 2443 1014
rect 2503 1010 2507 1014
rect 111 998 115 1002
rect 135 998 139 1002
rect 191 998 195 1002
rect 215 998 219 1002
rect 287 998 291 1002
rect 327 998 331 1002
rect 399 998 403 1002
rect 439 998 443 1002
rect 519 998 523 1002
rect 551 998 555 1002
rect 639 998 643 1002
rect 663 998 667 1002
rect 751 998 755 1002
rect 759 998 763 1002
rect 847 998 851 1002
rect 863 998 867 1002
rect 935 998 939 1002
rect 967 998 971 1002
rect 1015 998 1019 1002
rect 1079 998 1083 1002
rect 1087 998 1091 1002
rect 1167 998 1171 1002
rect 1191 998 1195 1002
rect 1223 998 1227 1002
rect 1287 998 1291 1002
rect 111 946 115 950
rect 151 946 155 950
rect 207 946 211 950
rect 231 946 235 950
rect 295 946 299 950
rect 343 946 347 950
rect 399 946 403 950
rect 455 946 459 950
rect 511 946 515 950
rect 567 946 571 950
rect 623 946 627 950
rect 679 946 683 950
rect 735 946 739 950
rect 775 946 779 950
rect 831 946 835 950
rect 863 946 867 950
rect 927 946 931 950
rect 951 946 955 950
rect 1015 946 1019 950
rect 1031 946 1035 950
rect 1095 946 1099 950
rect 1103 946 1107 950
rect 1175 946 1179 950
rect 1183 946 1187 950
rect 1239 946 1243 950
rect 1287 946 1291 950
rect 1327 942 1331 946
rect 1367 942 1371 946
rect 1439 942 1443 946
rect 1527 942 1531 946
rect 1583 942 1587 946
rect 1615 942 1619 946
rect 1639 942 1643 946
rect 1695 942 1699 946
rect 1751 942 1755 946
rect 1791 942 1795 946
rect 1823 942 1827 946
rect 1895 942 1899 946
rect 1903 942 1907 946
rect 1999 942 2003 946
rect 2015 942 2019 946
rect 2111 942 2115 946
rect 2151 942 2155 946
rect 2231 942 2235 946
rect 2295 942 2299 946
rect 2351 942 2355 946
rect 2439 942 2443 946
rect 2455 942 2459 946
rect 2503 942 2507 946
rect 111 890 115 894
rect 135 890 139 894
rect 191 890 195 894
rect 247 890 251 894
rect 279 890 283 894
rect 343 890 347 894
rect 383 890 387 894
rect 439 890 443 894
rect 495 890 499 894
rect 543 890 547 894
rect 607 890 611 894
rect 647 890 651 894
rect 719 890 723 894
rect 743 890 747 894
rect 815 890 819 894
rect 839 890 843 894
rect 911 890 915 894
rect 927 890 931 894
rect 999 890 1003 894
rect 1007 890 1011 894
rect 1079 890 1083 894
rect 1087 890 1091 894
rect 1159 890 1163 894
rect 1167 890 1171 894
rect 1223 890 1227 894
rect 1287 890 1291 894
rect 1327 882 1331 886
rect 1351 882 1355 886
rect 1423 882 1427 886
rect 1487 882 1491 886
rect 1511 882 1515 886
rect 1559 882 1563 886
rect 1599 882 1603 886
rect 1623 882 1627 886
rect 1679 882 1683 886
rect 1687 882 1691 886
rect 1751 882 1755 886
rect 1775 882 1779 886
rect 1815 882 1819 886
rect 1879 882 1883 886
rect 1887 882 1891 886
rect 1975 882 1979 886
rect 1999 882 2003 886
rect 2079 882 2083 886
rect 2135 882 2139 886
rect 2199 882 2203 886
rect 2279 882 2283 886
rect 2319 882 2323 886
rect 2423 882 2427 886
rect 2439 882 2443 886
rect 2503 882 2507 886
rect 111 834 115 838
rect 239 834 243 838
rect 263 834 267 838
rect 303 834 307 838
rect 359 834 363 838
rect 383 834 387 838
rect 455 834 459 838
rect 463 834 467 838
rect 551 834 555 838
rect 559 834 563 838
rect 639 834 643 838
rect 663 834 667 838
rect 727 834 731 838
rect 759 834 763 838
rect 807 834 811 838
rect 855 834 859 838
rect 895 834 899 838
rect 943 834 947 838
rect 983 834 987 838
rect 1023 834 1027 838
rect 1071 834 1075 838
rect 1103 834 1107 838
rect 1183 834 1187 838
rect 1239 834 1243 838
rect 1287 834 1291 838
rect 1327 822 1331 826
rect 1439 822 1443 826
rect 1503 822 1507 826
rect 1511 822 1515 826
rect 1575 822 1579 826
rect 1591 822 1595 826
rect 1639 822 1643 826
rect 1671 822 1675 826
rect 1703 822 1707 826
rect 1759 822 1763 826
rect 1767 822 1771 826
rect 1831 822 1835 826
rect 1847 822 1851 826
rect 1903 822 1907 826
rect 1935 822 1939 826
rect 1991 822 1995 826
rect 2023 822 2027 826
rect 2095 822 2099 826
rect 2111 822 2115 826
rect 2199 822 2203 826
rect 2215 822 2219 826
rect 2287 822 2291 826
rect 2335 822 2339 826
rect 2383 822 2387 826
rect 2455 822 2459 826
rect 2503 822 2507 826
rect 111 778 115 782
rect 151 778 155 782
rect 223 778 227 782
rect 247 778 251 782
rect 287 778 291 782
rect 343 778 347 782
rect 367 778 371 782
rect 439 778 443 782
rect 447 778 451 782
rect 527 778 531 782
rect 535 778 539 782
rect 607 778 611 782
rect 623 778 627 782
rect 679 778 683 782
rect 711 778 715 782
rect 751 778 755 782
rect 791 778 795 782
rect 823 778 827 782
rect 879 778 883 782
rect 895 778 899 782
rect 967 778 971 782
rect 975 778 979 782
rect 1055 778 1059 782
rect 1287 778 1291 782
rect 1327 766 1331 770
rect 1351 766 1355 770
rect 1423 766 1427 770
rect 1447 766 1451 770
rect 1495 766 1499 770
rect 1567 766 1571 770
rect 1575 766 1579 770
rect 1655 766 1659 770
rect 1687 766 1691 770
rect 1743 766 1747 770
rect 1807 766 1811 770
rect 1831 766 1835 770
rect 1919 766 1923 770
rect 1927 766 1931 770
rect 2007 766 2011 770
rect 2039 766 2043 770
rect 2095 766 2099 770
rect 2143 766 2147 770
rect 2183 766 2187 770
rect 2247 766 2251 770
rect 2271 766 2275 770
rect 2351 766 2355 770
rect 2367 766 2371 770
rect 2439 766 2443 770
rect 2503 766 2507 770
rect 111 722 115 726
rect 167 722 171 726
rect 175 722 179 726
rect 263 722 267 726
rect 343 722 347 726
rect 359 722 363 726
rect 423 722 427 726
rect 455 722 459 726
rect 503 722 507 726
rect 543 722 547 726
rect 575 722 579 726
rect 623 722 627 726
rect 639 722 643 726
rect 695 722 699 726
rect 703 722 707 726
rect 767 722 771 726
rect 839 722 843 726
rect 911 722 915 726
rect 991 722 995 726
rect 1287 722 1291 726
rect 1327 710 1331 714
rect 1367 710 1371 714
rect 1431 710 1435 714
rect 1463 710 1467 714
rect 1535 710 1539 714
rect 1583 710 1587 714
rect 1639 710 1643 714
rect 1703 710 1707 714
rect 1751 710 1755 714
rect 1823 710 1827 714
rect 1863 710 1867 714
rect 1943 710 1947 714
rect 1967 710 1971 714
rect 2055 710 2059 714
rect 2063 710 2067 714
rect 2151 710 2155 714
rect 2159 710 2163 714
rect 2231 710 2235 714
rect 2263 710 2267 714
rect 2311 710 2315 714
rect 2367 710 2371 714
rect 2391 710 2395 714
rect 2455 710 2459 714
rect 2503 710 2507 714
rect 111 670 115 674
rect 159 670 163 674
rect 215 670 219 674
rect 247 670 251 674
rect 295 670 299 674
rect 327 670 331 674
rect 375 670 379 674
rect 407 670 411 674
rect 455 670 459 674
rect 487 670 491 674
rect 527 670 531 674
rect 559 670 563 674
rect 591 670 595 674
rect 623 670 627 674
rect 655 670 659 674
rect 687 670 691 674
rect 719 670 723 674
rect 751 670 755 674
rect 783 670 787 674
rect 823 670 827 674
rect 847 670 851 674
rect 895 670 899 674
rect 919 670 923 674
rect 1287 670 1291 674
rect 1327 650 1331 654
rect 1351 650 1355 654
rect 1415 650 1419 654
rect 1479 650 1483 654
rect 1519 650 1523 654
rect 1559 650 1563 654
rect 1623 650 1627 654
rect 1647 650 1651 654
rect 1735 650 1739 654
rect 1831 650 1835 654
rect 1847 650 1851 654
rect 1919 650 1923 654
rect 1951 650 1955 654
rect 2007 650 2011 654
rect 2047 650 2051 654
rect 2087 650 2091 654
rect 2135 650 2139 654
rect 2167 650 2171 654
rect 2215 650 2219 654
rect 2239 650 2243 654
rect 2295 650 2299 654
rect 2311 650 2315 654
rect 2375 650 2379 654
rect 2383 650 2387 654
rect 2439 650 2443 654
rect 2503 650 2507 654
rect 111 614 115 618
rect 207 614 211 618
rect 231 614 235 618
rect 303 614 307 618
rect 311 614 315 618
rect 391 614 395 618
rect 407 614 411 618
rect 471 614 475 618
rect 503 614 507 618
rect 543 614 547 618
rect 599 614 603 618
rect 607 614 611 618
rect 671 614 675 618
rect 687 614 691 618
rect 735 614 739 618
rect 767 614 771 618
rect 799 614 803 618
rect 847 614 851 618
rect 863 614 867 618
rect 927 614 931 618
rect 935 614 939 618
rect 1007 614 1011 618
rect 1087 614 1091 618
rect 1287 614 1291 618
rect 1327 594 1331 598
rect 1455 594 1459 598
rect 1495 594 1499 598
rect 1559 594 1563 598
rect 1575 594 1579 598
rect 1663 594 1667 598
rect 1671 594 1675 598
rect 1751 594 1755 598
rect 1775 594 1779 598
rect 1847 594 1851 598
rect 1879 594 1883 598
rect 1935 594 1939 598
rect 1983 594 1987 598
rect 2023 594 2027 598
rect 2087 594 2091 598
rect 2103 594 2107 598
rect 2183 594 2187 598
rect 2255 594 2259 598
rect 2279 594 2283 598
rect 2327 594 2331 598
rect 2375 594 2379 598
rect 2399 594 2403 598
rect 2455 594 2459 598
rect 2503 594 2507 598
rect 111 558 115 562
rect 175 558 179 562
rect 191 558 195 562
rect 271 558 275 562
rect 287 558 291 562
rect 375 558 379 562
rect 391 558 395 562
rect 487 558 491 562
rect 583 558 587 562
rect 591 558 595 562
rect 671 558 675 562
rect 695 558 699 562
rect 751 558 755 562
rect 791 558 795 562
rect 831 558 835 562
rect 879 558 883 562
rect 911 558 915 562
rect 967 558 971 562
rect 991 558 995 562
rect 1055 558 1059 562
rect 1071 558 1075 562
rect 1151 558 1155 562
rect 1287 558 1291 562
rect 1327 538 1331 542
rect 1367 538 1371 542
rect 1439 538 1443 542
rect 1447 538 1451 542
rect 1527 538 1531 542
rect 1543 538 1547 542
rect 1615 538 1619 542
rect 1655 538 1659 542
rect 1711 538 1715 542
rect 1759 538 1763 542
rect 1799 538 1803 542
rect 1863 538 1867 542
rect 1887 538 1891 542
rect 1967 538 1971 542
rect 1975 538 1979 542
rect 2063 538 2067 542
rect 2071 538 2075 542
rect 2151 538 2155 542
rect 2167 538 2171 542
rect 2247 538 2251 542
rect 2263 538 2267 542
rect 2343 538 2347 542
rect 2359 538 2363 542
rect 2439 538 2443 542
rect 2503 538 2507 542
rect 111 502 115 506
rect 151 502 155 506
rect 191 502 195 506
rect 247 502 251 506
rect 287 502 291 506
rect 367 502 371 506
rect 391 502 395 506
rect 487 502 491 506
rect 503 502 507 506
rect 607 502 611 506
rect 615 502 619 506
rect 711 502 715 506
rect 735 502 739 506
rect 807 502 811 506
rect 847 502 851 506
rect 895 502 899 506
rect 951 502 955 506
rect 983 502 987 506
rect 1055 502 1059 506
rect 1071 502 1075 506
rect 1159 502 1163 506
rect 1167 502 1171 506
rect 1239 502 1243 506
rect 1287 502 1291 506
rect 1327 482 1331 486
rect 1367 482 1371 486
rect 1383 482 1387 486
rect 1431 482 1435 486
rect 1463 482 1467 486
rect 1519 482 1523 486
rect 1543 482 1547 486
rect 1615 482 1619 486
rect 1631 482 1635 486
rect 1711 482 1715 486
rect 1727 482 1731 486
rect 1815 482 1819 486
rect 1903 482 1907 486
rect 1927 482 1931 486
rect 1991 482 1995 486
rect 2055 482 2059 486
rect 2079 482 2083 486
rect 2167 482 2171 486
rect 2191 482 2195 486
rect 2263 482 2267 486
rect 2335 482 2339 486
rect 2359 482 2363 486
rect 2455 482 2459 486
rect 2503 482 2507 486
rect 111 446 115 450
rect 135 446 139 450
rect 191 446 195 450
rect 231 446 235 450
rect 247 446 251 450
rect 303 446 307 450
rect 351 446 355 450
rect 383 446 387 450
rect 471 446 475 450
rect 567 446 571 450
rect 599 446 603 450
rect 671 446 675 450
rect 719 446 723 450
rect 783 446 787 450
rect 831 446 835 450
rect 895 446 899 450
rect 935 446 939 450
rect 1007 446 1011 450
rect 1039 446 1043 450
rect 1127 446 1131 450
rect 1143 446 1147 450
rect 1223 446 1227 450
rect 1287 446 1291 450
rect 1327 426 1331 430
rect 1351 426 1355 430
rect 1415 426 1419 430
rect 1423 426 1427 430
rect 1503 426 1507 430
rect 1511 426 1515 430
rect 1599 426 1603 430
rect 1679 426 1683 430
rect 1695 426 1699 430
rect 1775 426 1779 430
rect 1799 426 1803 430
rect 1887 426 1891 430
rect 1911 426 1915 430
rect 2015 426 2019 430
rect 2039 426 2043 430
rect 2159 426 2163 430
rect 2175 426 2179 430
rect 2311 426 2315 430
rect 2319 426 2323 430
rect 2439 426 2443 430
rect 2503 426 2507 430
rect 111 386 115 390
rect 151 386 155 390
rect 207 386 211 390
rect 263 386 267 390
rect 279 386 283 390
rect 319 386 323 390
rect 359 386 363 390
rect 399 386 403 390
rect 431 386 435 390
rect 487 386 491 390
rect 511 386 515 390
rect 583 386 587 390
rect 591 386 595 390
rect 671 386 675 390
rect 687 386 691 390
rect 751 386 755 390
rect 799 386 803 390
rect 823 386 827 390
rect 895 386 899 390
rect 911 386 915 390
rect 967 386 971 390
rect 1023 386 1027 390
rect 1039 386 1043 390
rect 1111 386 1115 390
rect 1143 386 1147 390
rect 1183 386 1187 390
rect 1239 386 1243 390
rect 1287 386 1291 390
rect 1327 370 1331 374
rect 1367 370 1371 374
rect 1439 370 1443 374
rect 1527 370 1531 374
rect 1615 370 1619 374
rect 1679 370 1683 374
rect 1695 370 1699 374
rect 1735 370 1739 374
rect 1791 370 1795 374
rect 1807 370 1811 374
rect 1903 370 1907 374
rect 2023 370 2027 374
rect 2031 370 2035 374
rect 2159 370 2163 374
rect 2175 370 2179 374
rect 2303 370 2307 374
rect 2327 370 2331 374
rect 2455 370 2459 374
rect 2503 370 2507 374
rect 111 326 115 330
rect 135 326 139 330
rect 191 326 195 330
rect 199 326 203 330
rect 263 326 267 330
rect 287 326 291 330
rect 343 326 347 330
rect 375 326 379 330
rect 415 326 419 330
rect 455 326 459 330
rect 495 326 499 330
rect 543 326 547 330
rect 575 326 579 330
rect 631 326 635 330
rect 655 326 659 330
rect 727 326 731 330
rect 735 326 739 330
rect 807 326 811 330
rect 823 326 827 330
rect 879 326 883 330
rect 927 326 931 330
rect 951 326 955 330
rect 1023 326 1027 330
rect 1031 326 1035 330
rect 1095 326 1099 330
rect 1135 326 1139 330
rect 1167 326 1171 330
rect 1223 326 1227 330
rect 1287 326 1291 330
rect 1327 318 1331 322
rect 1351 318 1355 322
rect 1431 318 1435 322
rect 1527 318 1531 322
rect 1623 318 1627 322
rect 1663 318 1667 322
rect 1711 318 1715 322
rect 1719 318 1723 322
rect 1791 318 1795 322
rect 1807 318 1811 322
rect 1887 318 1891 322
rect 1911 318 1915 322
rect 2007 318 2011 322
rect 2023 318 2027 322
rect 2143 318 2147 322
rect 2151 318 2155 322
rect 2287 318 2291 322
rect 2423 318 2427 322
rect 2439 318 2443 322
rect 2503 318 2507 322
rect 111 266 115 270
rect 151 266 155 270
rect 215 266 219 270
rect 231 266 235 270
rect 303 266 307 270
rect 327 266 331 270
rect 391 266 395 270
rect 423 266 427 270
rect 471 266 475 270
rect 519 266 523 270
rect 559 266 563 270
rect 615 266 619 270
rect 647 266 651 270
rect 711 266 715 270
rect 743 266 747 270
rect 807 266 811 270
rect 839 266 843 270
rect 903 266 907 270
rect 943 266 947 270
rect 1007 266 1011 270
rect 1047 266 1051 270
rect 1111 266 1115 270
rect 1151 266 1155 270
rect 1215 266 1219 270
rect 1239 266 1243 270
rect 1287 266 1291 270
rect 1327 262 1331 266
rect 1367 262 1371 266
rect 1439 262 1443 266
rect 1447 262 1451 266
rect 1535 262 1539 266
rect 1543 262 1547 266
rect 1631 262 1635 266
rect 1639 262 1643 266
rect 1727 262 1731 266
rect 1815 262 1819 266
rect 1823 262 1827 266
rect 1903 262 1907 266
rect 1927 262 1931 266
rect 1999 262 2003 266
rect 2039 262 2043 266
rect 2103 262 2107 266
rect 2167 262 2171 266
rect 2215 262 2219 266
rect 2303 262 2307 266
rect 2335 262 2339 266
rect 2439 262 2443 266
rect 2455 262 2459 266
rect 2503 262 2507 266
rect 111 206 115 210
rect 135 206 139 210
rect 159 206 163 210
rect 215 206 219 210
rect 239 206 243 210
rect 311 206 315 210
rect 327 206 331 210
rect 407 206 411 210
rect 415 206 419 210
rect 503 206 507 210
rect 511 206 515 210
rect 599 206 603 210
rect 607 206 611 210
rect 695 206 699 210
rect 783 206 787 210
rect 791 206 795 210
rect 871 206 875 210
rect 887 206 891 210
rect 959 206 963 210
rect 991 206 995 210
rect 1047 206 1051 210
rect 1095 206 1099 210
rect 1135 206 1139 210
rect 1199 206 1203 210
rect 1287 206 1291 210
rect 1327 206 1331 210
rect 1351 206 1355 210
rect 1391 206 1395 210
rect 1423 206 1427 210
rect 1495 206 1499 210
rect 1519 206 1523 210
rect 1599 206 1603 210
rect 1615 206 1619 210
rect 1711 206 1715 210
rect 1799 206 1803 210
rect 1815 206 1819 210
rect 1887 206 1891 210
rect 1919 206 1923 210
rect 1983 206 1987 210
rect 2015 206 2019 210
rect 2087 206 2091 210
rect 2111 206 2115 210
rect 2199 206 2203 210
rect 2287 206 2291 210
rect 2319 206 2323 210
rect 2375 206 2379 210
rect 2439 206 2443 210
rect 2503 206 2507 210
rect 111 134 115 138
rect 151 134 155 138
rect 175 134 179 138
rect 207 134 211 138
rect 255 134 259 138
rect 263 134 267 138
rect 319 134 323 138
rect 343 134 347 138
rect 375 134 379 138
rect 431 134 435 138
rect 487 134 491 138
rect 527 134 531 138
rect 551 134 555 138
rect 623 134 627 138
rect 687 134 691 138
rect 711 134 715 138
rect 751 134 755 138
rect 799 134 803 138
rect 815 134 819 138
rect 879 134 883 138
rect 887 134 891 138
rect 943 134 947 138
rect 975 134 979 138
rect 1007 134 1011 138
rect 1063 134 1067 138
rect 1071 134 1075 138
rect 1135 134 1139 138
rect 1151 134 1155 138
rect 1199 134 1203 138
rect 1287 134 1291 138
rect 1327 134 1331 138
rect 1367 134 1371 138
rect 1407 134 1411 138
rect 1423 134 1427 138
rect 1479 134 1483 138
rect 1511 134 1515 138
rect 1535 134 1539 138
rect 1591 134 1595 138
rect 1615 134 1619 138
rect 1647 134 1651 138
rect 1703 134 1707 138
rect 1727 134 1731 138
rect 1759 134 1763 138
rect 1815 134 1819 138
rect 1831 134 1835 138
rect 1871 134 1875 138
rect 1927 134 1931 138
rect 1935 134 1939 138
rect 1983 134 1987 138
rect 2031 134 2035 138
rect 2039 134 2043 138
rect 2095 134 2099 138
rect 2127 134 2131 138
rect 2159 134 2163 138
rect 2215 134 2219 138
rect 2223 134 2227 138
rect 2287 134 2291 138
rect 2303 134 2307 138
rect 2343 134 2347 138
rect 2391 134 2395 138
rect 2399 134 2403 138
rect 2455 134 2459 138
rect 2503 134 2507 138
rect 111 82 115 86
rect 135 82 139 86
rect 191 82 195 86
rect 247 82 251 86
rect 303 82 307 86
rect 359 82 363 86
rect 415 82 419 86
rect 471 82 475 86
rect 535 82 539 86
rect 607 82 611 86
rect 671 82 675 86
rect 735 82 739 86
rect 799 82 803 86
rect 863 82 867 86
rect 927 82 931 86
rect 991 82 995 86
rect 1055 82 1059 86
rect 1119 82 1123 86
rect 1183 82 1187 86
rect 1287 82 1291 86
rect 1327 82 1331 86
rect 1351 82 1355 86
rect 1407 82 1411 86
rect 1463 82 1467 86
rect 1519 82 1523 86
rect 1575 82 1579 86
rect 1631 82 1635 86
rect 1687 82 1691 86
rect 1743 82 1747 86
rect 1799 82 1803 86
rect 1855 82 1859 86
rect 1911 82 1915 86
rect 1967 82 1971 86
rect 2023 82 2027 86
rect 2079 82 2083 86
rect 2143 82 2147 86
rect 2207 82 2211 86
rect 2271 82 2275 86
rect 2327 82 2331 86
rect 2383 82 2387 86
rect 2439 82 2443 86
rect 2503 82 2507 86
<< m4 >>
rect 96 2577 97 2583
rect 103 2582 1311 2583
rect 103 2578 111 2582
rect 115 2578 719 2582
rect 723 2578 775 2582
rect 779 2578 831 2582
rect 835 2578 887 2582
rect 891 2578 943 2582
rect 947 2578 1287 2582
rect 1291 2578 1311 2582
rect 103 2577 1311 2578
rect 1317 2577 1318 2583
rect 1310 2553 1311 2559
rect 1317 2558 2539 2559
rect 1317 2554 1327 2558
rect 1331 2554 1399 2558
rect 1403 2554 1455 2558
rect 1459 2554 1511 2558
rect 1515 2554 1567 2558
rect 1571 2554 1623 2558
rect 1627 2554 1679 2558
rect 1683 2554 1735 2558
rect 1739 2554 1791 2558
rect 1795 2554 1847 2558
rect 1851 2554 1903 2558
rect 1907 2554 1959 2558
rect 1963 2554 2015 2558
rect 2019 2554 2071 2558
rect 2075 2554 2127 2558
rect 2131 2554 2183 2558
rect 2187 2554 2503 2558
rect 2507 2554 2539 2558
rect 1317 2553 2539 2554
rect 2545 2553 2546 2559
rect 84 2525 85 2531
rect 91 2530 1299 2531
rect 91 2526 111 2530
rect 115 2526 167 2530
rect 171 2526 223 2530
rect 227 2526 279 2530
rect 283 2526 343 2530
rect 347 2526 407 2530
rect 411 2526 479 2530
rect 483 2526 559 2530
rect 563 2526 639 2530
rect 643 2526 703 2530
rect 707 2526 719 2530
rect 723 2526 759 2530
rect 763 2526 799 2530
rect 803 2526 815 2530
rect 819 2526 871 2530
rect 875 2526 879 2530
rect 883 2526 927 2530
rect 931 2526 959 2530
rect 963 2526 1039 2530
rect 1043 2526 1287 2530
rect 1291 2526 1299 2530
rect 91 2525 1299 2526
rect 1305 2525 1306 2531
rect 1298 2493 1299 2499
rect 1305 2498 2527 2499
rect 1305 2494 1327 2498
rect 1331 2494 1351 2498
rect 1355 2494 1383 2498
rect 1387 2494 1423 2498
rect 1427 2494 1439 2498
rect 1443 2494 1495 2498
rect 1499 2494 1511 2498
rect 1515 2494 1551 2498
rect 1555 2494 1599 2498
rect 1603 2494 1607 2498
rect 1611 2494 1663 2498
rect 1667 2494 1687 2498
rect 1691 2494 1719 2498
rect 1723 2494 1775 2498
rect 1779 2494 1831 2498
rect 1835 2494 1863 2498
rect 1867 2494 1887 2498
rect 1891 2494 1943 2498
rect 1947 2494 1951 2498
rect 1955 2494 1999 2498
rect 2003 2494 2039 2498
rect 2043 2494 2055 2498
rect 2059 2494 2111 2498
rect 2115 2494 2127 2498
rect 2131 2494 2167 2498
rect 2171 2494 2503 2498
rect 2507 2494 2527 2498
rect 1305 2493 2527 2494
rect 2533 2493 2534 2499
rect 96 2473 97 2479
rect 103 2478 1311 2479
rect 103 2474 111 2478
rect 115 2474 183 2478
rect 187 2474 239 2478
rect 243 2474 247 2478
rect 251 2474 295 2478
rect 299 2474 327 2478
rect 331 2474 359 2478
rect 363 2474 415 2478
rect 419 2474 423 2478
rect 427 2474 495 2478
rect 499 2474 503 2478
rect 507 2474 575 2478
rect 579 2474 599 2478
rect 603 2474 655 2478
rect 659 2474 695 2478
rect 699 2474 735 2478
rect 739 2474 791 2478
rect 795 2474 815 2478
rect 819 2474 879 2478
rect 883 2474 895 2478
rect 899 2474 967 2478
rect 971 2474 975 2478
rect 979 2474 1055 2478
rect 1059 2474 1063 2478
rect 1067 2474 1159 2478
rect 1163 2474 1287 2478
rect 1291 2474 1311 2478
rect 103 2473 1311 2474
rect 1317 2473 1318 2479
rect 1310 2433 1311 2439
rect 1317 2438 2539 2439
rect 1317 2434 1327 2438
rect 1331 2434 1367 2438
rect 1371 2434 1439 2438
rect 1443 2434 1527 2438
rect 1531 2434 1543 2438
rect 1547 2434 1615 2438
rect 1619 2434 1639 2438
rect 1643 2434 1703 2438
rect 1707 2434 1735 2438
rect 1739 2434 1791 2438
rect 1795 2434 1823 2438
rect 1827 2434 1879 2438
rect 1883 2434 1911 2438
rect 1915 2434 1967 2438
rect 1971 2434 2007 2438
rect 2011 2434 2055 2438
rect 2059 2434 2103 2438
rect 2107 2434 2143 2438
rect 2147 2434 2503 2438
rect 2507 2434 2539 2438
rect 1317 2433 2539 2434
rect 2545 2433 2546 2439
rect 84 2417 85 2423
rect 91 2422 1299 2423
rect 91 2418 111 2422
rect 115 2418 151 2422
rect 155 2418 167 2422
rect 171 2418 231 2422
rect 235 2418 311 2422
rect 315 2418 319 2422
rect 323 2418 399 2422
rect 403 2418 415 2422
rect 419 2418 487 2422
rect 491 2418 519 2422
rect 523 2418 583 2422
rect 587 2418 623 2422
rect 627 2418 679 2422
rect 683 2418 727 2422
rect 731 2418 775 2422
rect 779 2418 831 2422
rect 835 2418 863 2422
rect 867 2418 935 2422
rect 939 2418 951 2422
rect 955 2418 1039 2422
rect 1043 2418 1047 2422
rect 1051 2418 1143 2422
rect 1147 2418 1151 2422
rect 1155 2418 1287 2422
rect 1291 2418 1299 2422
rect 91 2417 1299 2418
rect 1305 2417 1306 2423
rect 1298 2375 1299 2381
rect 1305 2379 1330 2381
rect 1305 2378 2527 2379
rect 1305 2375 1327 2378
rect 1324 2374 1327 2375
rect 1331 2374 1351 2378
rect 1355 2374 1407 2378
rect 1411 2374 1423 2378
rect 1427 2374 1495 2378
rect 1499 2374 1527 2378
rect 1531 2374 1583 2378
rect 1587 2374 1623 2378
rect 1627 2374 1671 2378
rect 1675 2374 1719 2378
rect 1723 2374 1751 2378
rect 1755 2374 1807 2378
rect 1811 2374 1831 2378
rect 1835 2374 1895 2378
rect 1899 2374 1919 2378
rect 1923 2374 1991 2378
rect 1995 2374 2007 2378
rect 2011 2374 2087 2378
rect 2091 2374 2095 2378
rect 2099 2374 2503 2378
rect 2507 2374 2527 2378
rect 1324 2373 2527 2374
rect 2533 2373 2534 2379
rect 96 2365 97 2371
rect 103 2370 1311 2371
rect 103 2366 111 2370
rect 115 2366 167 2370
rect 171 2366 175 2370
rect 179 2366 247 2370
rect 251 2366 279 2370
rect 283 2366 335 2370
rect 339 2366 391 2370
rect 395 2366 431 2370
rect 435 2366 503 2370
rect 507 2366 535 2370
rect 539 2366 623 2370
rect 627 2366 639 2370
rect 643 2366 743 2370
rect 747 2366 847 2370
rect 851 2366 871 2370
rect 875 2366 951 2370
rect 955 2366 999 2370
rect 1003 2366 1055 2370
rect 1059 2366 1127 2370
rect 1131 2366 1167 2370
rect 1171 2366 1287 2370
rect 1291 2366 1311 2370
rect 103 2365 1311 2366
rect 1317 2365 1318 2371
rect 1310 2317 1311 2323
rect 1317 2322 2539 2323
rect 1317 2318 1327 2322
rect 1331 2318 1367 2322
rect 1371 2318 1423 2322
rect 1427 2318 1455 2322
rect 1459 2318 1511 2322
rect 1515 2318 1543 2322
rect 1547 2318 1599 2322
rect 1603 2318 1639 2322
rect 1643 2318 1687 2322
rect 1691 2318 1735 2322
rect 1739 2318 1767 2322
rect 1771 2318 1831 2322
rect 1835 2318 1847 2322
rect 1851 2318 1927 2322
rect 1931 2318 1935 2322
rect 1939 2318 2015 2322
rect 2019 2318 2023 2322
rect 2027 2318 2111 2322
rect 2115 2318 2207 2322
rect 2211 2318 2503 2322
rect 2507 2318 2539 2322
rect 1317 2317 2539 2318
rect 2545 2317 2546 2323
rect 84 2309 85 2315
rect 91 2314 1299 2315
rect 91 2310 111 2314
rect 115 2310 159 2314
rect 163 2310 207 2314
rect 211 2310 263 2314
rect 267 2310 287 2314
rect 291 2310 375 2314
rect 379 2310 471 2314
rect 475 2310 487 2314
rect 491 2310 559 2314
rect 563 2310 607 2314
rect 611 2310 647 2314
rect 651 2310 727 2314
rect 731 2310 735 2314
rect 739 2310 815 2314
rect 819 2310 855 2314
rect 859 2310 903 2314
rect 907 2310 983 2314
rect 987 2310 991 2314
rect 995 2310 1079 2314
rect 1083 2310 1111 2314
rect 1115 2310 1287 2314
rect 1291 2310 1299 2314
rect 91 2309 1299 2310
rect 1305 2309 1306 2315
rect 1298 2265 1299 2271
rect 1305 2270 2527 2271
rect 1305 2266 1327 2270
rect 1331 2266 1351 2270
rect 1355 2266 1439 2270
rect 1443 2266 1455 2270
rect 1459 2266 1527 2270
rect 1531 2266 1543 2270
rect 1547 2266 1623 2270
rect 1627 2266 1639 2270
rect 1643 2266 1719 2270
rect 1723 2266 1735 2270
rect 1739 2266 1815 2270
rect 1819 2266 1839 2270
rect 1843 2266 1911 2270
rect 1915 2266 1935 2270
rect 1939 2266 1999 2270
rect 2003 2266 2031 2270
rect 2035 2266 2095 2270
rect 2099 2266 2119 2270
rect 2123 2266 2191 2270
rect 2195 2266 2215 2270
rect 2219 2266 2311 2270
rect 2315 2266 2503 2270
rect 2507 2266 2527 2270
rect 1305 2265 2527 2266
rect 2533 2265 2534 2271
rect 96 2253 97 2259
rect 103 2258 1311 2259
rect 103 2254 111 2258
rect 115 2254 223 2258
rect 227 2254 263 2258
rect 267 2254 303 2258
rect 307 2254 319 2258
rect 323 2254 383 2258
rect 387 2254 391 2258
rect 395 2254 447 2258
rect 451 2254 487 2258
rect 491 2254 503 2258
rect 507 2254 559 2258
rect 563 2254 575 2258
rect 579 2254 615 2258
rect 619 2254 663 2258
rect 667 2254 671 2258
rect 675 2254 727 2258
rect 731 2254 751 2258
rect 755 2254 791 2258
rect 795 2254 831 2258
rect 835 2254 855 2258
rect 859 2254 919 2258
rect 923 2254 983 2258
rect 987 2254 1007 2258
rect 1011 2254 1047 2258
rect 1051 2254 1095 2258
rect 1099 2254 1111 2258
rect 1115 2254 1287 2258
rect 1291 2254 1311 2258
rect 103 2253 1311 2254
rect 1317 2253 1318 2259
rect 1310 2209 1311 2215
rect 1317 2214 2539 2215
rect 1317 2210 1327 2214
rect 1331 2210 1471 2214
rect 1475 2210 1559 2214
rect 1563 2210 1567 2214
rect 1571 2210 1623 2214
rect 1627 2210 1655 2214
rect 1659 2210 1679 2214
rect 1683 2210 1743 2214
rect 1747 2210 1751 2214
rect 1755 2210 1807 2214
rect 1811 2210 1855 2214
rect 1859 2210 1871 2214
rect 1875 2210 1927 2214
rect 1931 2210 1951 2214
rect 1955 2210 1983 2214
rect 1987 2210 2039 2214
rect 2043 2210 2047 2214
rect 2051 2210 2095 2214
rect 2099 2210 2135 2214
rect 2139 2210 2159 2214
rect 2163 2210 2223 2214
rect 2227 2210 2231 2214
rect 2235 2210 2287 2214
rect 2291 2210 2327 2214
rect 2331 2210 2343 2214
rect 2347 2210 2399 2214
rect 2403 2210 2455 2214
rect 2459 2210 2503 2214
rect 2507 2210 2539 2214
rect 1317 2209 2539 2210
rect 2545 2209 2546 2215
rect 84 2197 85 2203
rect 91 2202 1299 2203
rect 91 2198 111 2202
rect 115 2198 247 2202
rect 251 2198 303 2202
rect 307 2198 335 2202
rect 339 2198 367 2202
rect 371 2198 391 2202
rect 395 2198 431 2202
rect 435 2198 447 2202
rect 451 2198 487 2202
rect 491 2198 503 2202
rect 507 2198 543 2202
rect 547 2198 559 2202
rect 563 2198 599 2202
rect 603 2198 655 2202
rect 659 2198 711 2202
rect 715 2198 775 2202
rect 779 2198 839 2202
rect 843 2198 903 2202
rect 907 2198 967 2202
rect 971 2198 1031 2202
rect 1035 2198 1095 2202
rect 1099 2198 1287 2202
rect 1291 2198 1299 2202
rect 91 2197 1299 2198
rect 1305 2197 1306 2203
rect 1298 2155 1299 2161
rect 1305 2155 1330 2161
rect 1324 2151 1330 2155
rect 96 2145 97 2151
rect 103 2150 1311 2151
rect 103 2146 111 2150
rect 115 2146 351 2150
rect 355 2146 407 2150
rect 411 2146 415 2150
rect 419 2146 463 2150
rect 467 2146 511 2150
rect 515 2146 519 2150
rect 523 2146 575 2150
rect 579 2146 607 2150
rect 611 2146 711 2150
rect 715 2146 815 2150
rect 819 2146 927 2150
rect 931 2146 1039 2150
rect 1043 2146 1151 2150
rect 1155 2146 1239 2150
rect 1243 2146 1287 2150
rect 1291 2146 1311 2150
rect 103 2145 1311 2146
rect 1317 2145 1318 2151
rect 1324 2150 2527 2151
rect 1324 2146 1327 2150
rect 1331 2146 1551 2150
rect 1555 2146 1607 2150
rect 1611 2146 1663 2150
rect 1667 2146 1719 2150
rect 1723 2146 1727 2150
rect 1731 2146 1791 2150
rect 1795 2146 1855 2150
rect 1859 2146 1871 2150
rect 1875 2146 1911 2150
rect 1915 2146 1967 2150
rect 1971 2146 2023 2150
rect 2027 2146 2079 2150
rect 2083 2146 2143 2150
rect 2147 2146 2199 2150
rect 2203 2146 2207 2150
rect 2211 2146 2271 2150
rect 2275 2146 2327 2150
rect 2331 2146 2383 2150
rect 2387 2146 2439 2150
rect 2443 2146 2503 2150
rect 2507 2146 2527 2150
rect 1324 2145 2527 2146
rect 2533 2145 2534 2151
rect 84 2093 85 2099
rect 91 2098 1299 2099
rect 91 2094 111 2098
rect 115 2094 375 2098
rect 379 2094 399 2098
rect 403 2094 447 2098
rect 451 2094 495 2098
rect 499 2094 519 2098
rect 523 2094 591 2098
rect 595 2094 599 2098
rect 603 2094 679 2098
rect 683 2094 695 2098
rect 699 2094 759 2098
rect 763 2094 799 2098
rect 803 2094 831 2098
rect 835 2094 903 2098
rect 907 2094 911 2098
rect 915 2094 967 2098
rect 971 2094 1023 2098
rect 1027 2094 1031 2098
rect 1035 2094 1103 2098
rect 1107 2094 1135 2098
rect 1139 2094 1167 2098
rect 1171 2094 1223 2098
rect 1227 2094 1287 2098
rect 1291 2094 1299 2098
rect 91 2093 1299 2094
rect 1305 2093 1306 2099
rect 1310 2081 1311 2087
rect 1317 2086 2539 2087
rect 1317 2082 1327 2086
rect 1331 2082 1367 2086
rect 1371 2082 1423 2086
rect 1427 2082 1503 2086
rect 1507 2082 1591 2086
rect 1595 2082 1679 2086
rect 1683 2082 1735 2086
rect 1739 2082 1783 2086
rect 1787 2082 1807 2086
rect 1811 2082 1887 2086
rect 1891 2082 1895 2086
rect 1899 2082 1983 2086
rect 1987 2082 2023 2086
rect 2027 2082 2095 2086
rect 2099 2082 2167 2086
rect 2171 2082 2215 2086
rect 2219 2082 2319 2086
rect 2323 2082 2343 2086
rect 2347 2082 2455 2086
rect 2459 2082 2503 2086
rect 2507 2082 2539 2086
rect 1317 2081 2539 2082
rect 2545 2081 2546 2087
rect 1298 2047 1299 2053
rect 1305 2047 1330 2053
rect 96 2037 97 2043
rect 103 2042 1311 2043
rect 103 2038 111 2042
rect 115 2038 295 2042
rect 299 2038 375 2042
rect 379 2038 391 2042
rect 395 2038 463 2042
rect 467 2038 535 2042
rect 539 2038 551 2042
rect 555 2038 615 2042
rect 619 2038 639 2042
rect 643 2038 695 2042
rect 699 2038 719 2042
rect 723 2038 775 2042
rect 779 2038 799 2042
rect 803 2038 847 2042
rect 851 2038 887 2042
rect 891 2038 919 2042
rect 923 2038 975 2042
rect 979 2038 983 2042
rect 987 2038 1047 2042
rect 1051 2038 1063 2042
rect 1067 2038 1119 2042
rect 1123 2038 1183 2042
rect 1187 2038 1239 2042
rect 1243 2038 1287 2042
rect 1291 2038 1311 2042
rect 103 2037 1311 2038
rect 1317 2037 1318 2043
rect 1324 2035 1330 2047
rect 1324 2034 2527 2035
rect 1324 2030 1327 2034
rect 1331 2030 1351 2034
rect 1355 2030 1407 2034
rect 1411 2030 1423 2034
rect 1427 2030 1487 2034
rect 1491 2030 1519 2034
rect 1523 2030 1575 2034
rect 1579 2030 1615 2034
rect 1619 2030 1663 2034
rect 1667 2030 1719 2034
rect 1723 2030 1767 2034
rect 1771 2030 1823 2034
rect 1827 2030 1879 2034
rect 1883 2030 1935 2034
rect 1939 2030 2007 2034
rect 2011 2030 2055 2034
rect 2059 2030 2151 2034
rect 2155 2030 2183 2034
rect 2187 2030 2303 2034
rect 2307 2030 2319 2034
rect 2323 2030 2439 2034
rect 2443 2030 2503 2034
rect 2507 2030 2527 2034
rect 1324 2029 2527 2030
rect 2533 2029 2534 2035
rect 84 1981 85 1987
rect 91 1986 1299 1987
rect 91 1982 111 1986
rect 115 1982 135 1986
rect 139 1982 207 1986
rect 211 1982 279 1986
rect 283 1982 287 1986
rect 291 1982 359 1986
rect 363 1982 383 1986
rect 387 1982 447 1986
rect 451 1982 487 1986
rect 491 1982 535 1986
rect 539 1982 591 1986
rect 595 1982 623 1986
rect 627 1982 695 1986
rect 699 1982 703 1986
rect 707 1982 783 1986
rect 787 1982 799 1986
rect 803 1982 871 1986
rect 875 1982 903 1986
rect 907 1982 959 1986
rect 963 1982 1015 1986
rect 1019 1982 1047 1986
rect 1051 1982 1287 1986
rect 1291 1982 1299 1986
rect 91 1981 1299 1982
rect 1305 1981 1306 1987
rect 1310 1973 1311 1979
rect 1317 1978 2539 1979
rect 1317 1974 1327 1978
rect 1331 1974 1367 1978
rect 1371 1974 1439 1978
rect 1443 1974 1455 1978
rect 1459 1974 1535 1978
rect 1539 1974 1543 1978
rect 1547 1974 1631 1978
rect 1635 1974 1639 1978
rect 1643 1974 1735 1978
rect 1739 1974 1839 1978
rect 1843 1974 1943 1978
rect 1947 1974 1951 1978
rect 1955 1974 2047 1978
rect 2051 1974 2071 1978
rect 2075 1974 2151 1978
rect 2155 1974 2199 1978
rect 2203 1974 2255 1978
rect 2259 1974 2335 1978
rect 2339 1974 2367 1978
rect 2371 1974 2455 1978
rect 2459 1974 2503 1978
rect 2507 1974 2539 1978
rect 1317 1973 2539 1974
rect 2545 1973 2546 1979
rect 1298 1931 1299 1937
rect 1305 1931 1330 1937
rect 96 1921 97 1927
rect 103 1926 1311 1927
rect 103 1922 111 1926
rect 115 1922 151 1926
rect 155 1922 223 1926
rect 227 1922 239 1926
rect 243 1922 303 1926
rect 307 1922 375 1926
rect 379 1922 399 1926
rect 403 1922 503 1926
rect 507 1922 527 1926
rect 531 1922 607 1926
rect 611 1922 687 1926
rect 691 1922 711 1926
rect 715 1922 815 1926
rect 819 1922 863 1926
rect 867 1922 919 1926
rect 923 1922 1031 1926
rect 1035 1922 1039 1926
rect 1043 1922 1287 1926
rect 1291 1922 1311 1926
rect 103 1921 1311 1922
rect 1317 1921 1318 1927
rect 1324 1923 1330 1931
rect 1324 1922 2527 1923
rect 1324 1918 1327 1922
rect 1331 1918 1439 1922
rect 1443 1918 1527 1922
rect 1531 1918 1615 1922
rect 1619 1918 1623 1922
rect 1627 1918 1711 1922
rect 1715 1918 1719 1922
rect 1723 1918 1815 1922
rect 1819 1918 1823 1922
rect 1827 1918 1919 1922
rect 1923 1918 1927 1922
rect 1931 1918 2015 1922
rect 2019 1918 2031 1922
rect 2035 1918 2111 1922
rect 2115 1918 2135 1922
rect 2139 1918 2199 1922
rect 2203 1918 2239 1922
rect 2243 1918 2287 1922
rect 2291 1918 2351 1922
rect 2355 1918 2375 1922
rect 2379 1918 2439 1922
rect 2443 1918 2503 1922
rect 2507 1918 2527 1922
rect 1324 1917 2527 1918
rect 2533 1917 2534 1923
rect 84 1869 85 1875
rect 91 1874 1299 1875
rect 91 1870 111 1874
rect 115 1870 135 1874
rect 139 1870 191 1874
rect 195 1870 223 1874
rect 227 1870 263 1874
rect 267 1870 335 1874
rect 339 1870 359 1874
rect 363 1870 407 1874
rect 411 1870 479 1874
rect 483 1870 511 1874
rect 515 1870 551 1874
rect 555 1870 615 1874
rect 619 1870 671 1874
rect 675 1870 679 1874
rect 683 1870 743 1874
rect 747 1870 815 1874
rect 819 1870 847 1874
rect 851 1870 887 1874
rect 891 1870 959 1874
rect 963 1870 1023 1874
rect 1027 1870 1039 1874
rect 1043 1870 1287 1874
rect 1291 1870 1299 1874
rect 91 1869 1299 1870
rect 1305 1869 1306 1875
rect 1310 1865 1311 1871
rect 1317 1870 2539 1871
rect 1317 1866 1327 1870
rect 1331 1866 1535 1870
rect 1539 1866 1543 1870
rect 1547 1866 1607 1870
rect 1611 1866 1631 1870
rect 1635 1866 1687 1870
rect 1691 1866 1727 1870
rect 1731 1866 1783 1870
rect 1787 1866 1831 1870
rect 1835 1866 1879 1870
rect 1883 1866 1935 1870
rect 1939 1866 1983 1870
rect 1987 1866 2031 1870
rect 2035 1866 2079 1870
rect 2083 1866 2127 1870
rect 2131 1866 2175 1870
rect 2179 1866 2215 1870
rect 2219 1866 2271 1870
rect 2275 1866 2303 1870
rect 2307 1866 2367 1870
rect 2371 1866 2391 1870
rect 2395 1866 2455 1870
rect 2459 1866 2503 1870
rect 2507 1866 2539 1870
rect 1317 1865 2539 1866
rect 2545 1865 2546 1871
rect 1298 1819 1299 1825
rect 1305 1819 1330 1825
rect 1324 1815 1330 1819
rect 96 1809 97 1815
rect 103 1814 1311 1815
rect 103 1810 111 1814
rect 115 1810 151 1814
rect 155 1810 207 1814
rect 211 1810 231 1814
rect 235 1810 279 1814
rect 283 1810 335 1814
rect 339 1810 351 1814
rect 355 1810 423 1814
rect 427 1810 439 1814
rect 443 1810 495 1814
rect 499 1810 535 1814
rect 539 1810 567 1814
rect 571 1810 631 1814
rect 635 1810 695 1814
rect 699 1810 719 1814
rect 723 1810 759 1814
rect 763 1810 799 1814
rect 803 1810 831 1814
rect 835 1810 879 1814
rect 883 1810 903 1814
rect 907 1810 959 1814
rect 963 1810 975 1814
rect 979 1810 1039 1814
rect 1043 1810 1055 1814
rect 1059 1810 1119 1814
rect 1123 1810 1287 1814
rect 1291 1810 1311 1814
rect 103 1809 1311 1810
rect 1317 1809 1318 1815
rect 1324 1814 2527 1815
rect 1324 1810 1327 1814
rect 1331 1810 1463 1814
rect 1467 1810 1519 1814
rect 1523 1810 1559 1814
rect 1563 1810 1591 1814
rect 1595 1810 1663 1814
rect 1667 1810 1671 1814
rect 1675 1810 1767 1814
rect 1771 1810 1863 1814
rect 1867 1810 1879 1814
rect 1883 1810 1967 1814
rect 1971 1810 1983 1814
rect 1987 1810 2063 1814
rect 2067 1810 2087 1814
rect 2091 1810 2159 1814
rect 2163 1810 2183 1814
rect 2187 1810 2255 1814
rect 2259 1810 2271 1814
rect 2275 1810 2351 1814
rect 2355 1810 2367 1814
rect 2371 1810 2439 1814
rect 2443 1810 2503 1814
rect 2507 1810 2527 1814
rect 1324 1809 2527 1810
rect 2533 1809 2534 1815
rect 84 1753 85 1759
rect 91 1758 1299 1759
rect 91 1754 111 1758
rect 115 1754 135 1758
rect 139 1754 215 1758
rect 219 1754 239 1758
rect 243 1754 319 1758
rect 323 1754 351 1758
rect 355 1754 423 1758
rect 427 1754 463 1758
rect 467 1754 519 1758
rect 523 1754 575 1758
rect 579 1754 615 1758
rect 619 1754 679 1758
rect 683 1754 703 1758
rect 707 1754 783 1758
rect 787 1754 863 1758
rect 867 1754 887 1758
rect 891 1754 943 1758
rect 947 1754 991 1758
rect 995 1754 1023 1758
rect 1027 1754 1103 1758
rect 1107 1754 1287 1758
rect 1291 1754 1299 1758
rect 91 1753 1299 1754
rect 1305 1753 1306 1759
rect 1310 1753 1311 1759
rect 1317 1758 2539 1759
rect 1317 1754 1327 1758
rect 1331 1754 1375 1758
rect 1379 1754 1471 1758
rect 1475 1754 1479 1758
rect 1483 1754 1567 1758
rect 1571 1754 1575 1758
rect 1579 1754 1671 1758
rect 1675 1754 1679 1758
rect 1683 1754 1775 1758
rect 1779 1754 1783 1758
rect 1787 1754 1887 1758
rect 1891 1754 1895 1758
rect 1899 1754 1999 1758
rect 2003 1754 2103 1758
rect 2107 1754 2111 1758
rect 2115 1754 2199 1758
rect 2203 1754 2231 1758
rect 2235 1754 2287 1758
rect 2291 1754 2351 1758
rect 2355 1754 2383 1758
rect 2387 1754 2455 1758
rect 2459 1754 2503 1758
rect 2507 1754 2539 1758
rect 1317 1753 2539 1754
rect 2545 1753 2546 1759
rect 1298 1707 1299 1713
rect 1305 1707 1330 1713
rect 1324 1706 2527 1707
rect 96 1697 97 1703
rect 103 1702 1311 1703
rect 103 1698 111 1702
rect 115 1698 151 1702
rect 155 1698 191 1702
rect 195 1698 255 1702
rect 259 1698 271 1702
rect 275 1698 351 1702
rect 355 1698 367 1702
rect 371 1698 439 1702
rect 443 1698 479 1702
rect 483 1698 535 1702
rect 539 1698 591 1702
rect 595 1698 639 1702
rect 643 1698 695 1702
rect 699 1698 743 1702
rect 747 1698 799 1702
rect 803 1698 847 1702
rect 851 1698 903 1702
rect 907 1698 951 1702
rect 955 1698 1007 1702
rect 1011 1698 1063 1702
rect 1067 1698 1119 1702
rect 1123 1698 1175 1702
rect 1179 1698 1287 1702
rect 1291 1698 1311 1702
rect 103 1697 1311 1698
rect 1317 1697 1318 1703
rect 1324 1702 1327 1706
rect 1331 1702 1351 1706
rect 1355 1702 1359 1706
rect 1363 1702 1431 1706
rect 1435 1702 1455 1706
rect 1459 1702 1535 1706
rect 1539 1702 1551 1706
rect 1555 1702 1647 1706
rect 1651 1702 1655 1706
rect 1659 1702 1759 1706
rect 1763 1702 1871 1706
rect 1875 1702 1879 1706
rect 1883 1702 1983 1706
rect 1987 1702 2015 1706
rect 2019 1702 2095 1706
rect 2099 1702 2159 1706
rect 2163 1702 2215 1706
rect 2219 1702 2311 1706
rect 2315 1702 2335 1706
rect 2339 1702 2439 1706
rect 2443 1702 2503 1706
rect 2507 1702 2527 1706
rect 1324 1701 2527 1702
rect 2533 1701 2534 1707
rect 84 1645 85 1651
rect 91 1650 1299 1651
rect 91 1646 111 1650
rect 115 1646 175 1650
rect 179 1646 215 1650
rect 219 1646 255 1650
rect 259 1646 271 1650
rect 275 1646 335 1650
rect 339 1646 407 1650
rect 411 1646 423 1650
rect 427 1646 479 1650
rect 483 1646 519 1650
rect 523 1646 559 1650
rect 563 1646 623 1650
rect 627 1646 647 1650
rect 651 1646 727 1650
rect 731 1646 743 1650
rect 747 1646 831 1650
rect 835 1646 839 1650
rect 843 1646 935 1650
rect 939 1646 943 1650
rect 947 1646 1047 1650
rect 1051 1646 1055 1650
rect 1059 1646 1159 1650
rect 1163 1646 1175 1650
rect 1179 1646 1287 1650
rect 1291 1646 1299 1650
rect 91 1645 1299 1646
rect 1305 1645 1306 1651
rect 1310 1641 1311 1647
rect 1317 1646 2539 1647
rect 1317 1642 1327 1646
rect 1331 1642 1367 1646
rect 1371 1642 1431 1646
rect 1435 1642 1447 1646
rect 1451 1642 1519 1646
rect 1523 1642 1551 1646
rect 1555 1642 1599 1646
rect 1603 1642 1663 1646
rect 1667 1642 1679 1646
rect 1683 1642 1751 1646
rect 1755 1642 1775 1646
rect 1779 1642 1839 1646
rect 1843 1642 1895 1646
rect 1899 1642 1935 1646
rect 1939 1642 2031 1646
rect 2035 1642 2055 1646
rect 2059 1642 2175 1646
rect 2179 1642 2183 1646
rect 2187 1642 2327 1646
rect 2331 1642 2455 1646
rect 2459 1642 2503 1646
rect 2507 1642 2539 1646
rect 1317 1641 2539 1642
rect 2545 1641 2546 1647
rect 1298 1603 1299 1609
rect 1305 1603 1330 1609
rect 96 1593 97 1599
rect 103 1598 1311 1599
rect 103 1594 111 1598
rect 115 1594 231 1598
rect 235 1594 287 1598
rect 291 1594 351 1598
rect 355 1594 423 1598
rect 427 1594 495 1598
rect 499 1594 503 1598
rect 507 1594 575 1598
rect 579 1594 599 1598
rect 603 1594 663 1598
rect 667 1594 703 1598
rect 707 1594 759 1598
rect 763 1594 815 1598
rect 819 1594 855 1598
rect 859 1594 935 1598
rect 939 1594 959 1598
rect 963 1594 1063 1598
rect 1067 1594 1071 1598
rect 1075 1594 1191 1598
rect 1195 1594 1287 1598
rect 1291 1594 1311 1598
rect 103 1593 1311 1594
rect 1317 1593 1318 1599
rect 1324 1591 1330 1603
rect 1324 1590 2527 1591
rect 1324 1586 1327 1590
rect 1331 1586 1351 1590
rect 1355 1586 1415 1590
rect 1419 1586 1423 1590
rect 1427 1586 1503 1590
rect 1507 1586 1527 1590
rect 1531 1586 1583 1590
rect 1587 1586 1647 1590
rect 1651 1586 1663 1590
rect 1667 1586 1735 1590
rect 1739 1586 1783 1590
rect 1787 1586 1823 1590
rect 1827 1586 1919 1590
rect 1923 1586 1935 1590
rect 1939 1586 2039 1590
rect 2043 1586 2103 1590
rect 2107 1586 2167 1590
rect 2171 1586 2279 1590
rect 2283 1586 2311 1590
rect 2315 1586 2439 1590
rect 2443 1586 2503 1590
rect 2507 1586 2527 1590
rect 1324 1585 2527 1586
rect 2533 1585 2534 1591
rect 84 1533 85 1539
rect 91 1538 1299 1539
rect 91 1534 111 1538
rect 115 1534 271 1538
rect 275 1534 335 1538
rect 339 1534 407 1538
rect 411 1534 471 1538
rect 475 1534 487 1538
rect 491 1534 551 1538
rect 555 1534 583 1538
rect 587 1534 639 1538
rect 643 1534 687 1538
rect 691 1534 735 1538
rect 739 1534 799 1538
rect 803 1534 839 1538
rect 843 1534 919 1538
rect 923 1534 951 1538
rect 955 1534 1047 1538
rect 1051 1534 1063 1538
rect 1067 1534 1175 1538
rect 1179 1534 1287 1538
rect 1291 1534 1299 1538
rect 91 1533 1299 1534
rect 1305 1533 1306 1539
rect 1310 1533 1311 1539
rect 1317 1538 2539 1539
rect 1317 1534 1327 1538
rect 1331 1534 1367 1538
rect 1371 1534 1439 1538
rect 1443 1534 1543 1538
rect 1547 1534 1647 1538
rect 1651 1534 1663 1538
rect 1667 1534 1751 1538
rect 1755 1534 1799 1538
rect 1803 1534 1855 1538
rect 1859 1534 1951 1538
rect 1955 1534 1959 1538
rect 1963 1534 2055 1538
rect 2059 1534 2119 1538
rect 2123 1534 2151 1538
rect 2155 1534 2247 1538
rect 2251 1534 2295 1538
rect 2299 1534 2343 1538
rect 2347 1534 2439 1538
rect 2443 1534 2455 1538
rect 2459 1534 2503 1538
rect 2507 1534 2539 1538
rect 1317 1533 2539 1534
rect 2545 1533 2546 1539
rect 1298 1491 1299 1497
rect 1305 1491 1330 1497
rect 96 1481 97 1487
rect 103 1486 1311 1487
rect 103 1482 111 1486
rect 115 1482 375 1486
rect 379 1482 463 1486
rect 467 1482 487 1486
rect 491 1482 559 1486
rect 563 1482 567 1486
rect 571 1482 655 1486
rect 659 1482 751 1486
rect 755 1482 855 1486
rect 859 1482 959 1486
rect 963 1482 967 1486
rect 971 1482 1063 1486
rect 1067 1482 1079 1486
rect 1083 1482 1167 1486
rect 1171 1482 1191 1486
rect 1195 1482 1287 1486
rect 1291 1482 1311 1486
rect 103 1481 1311 1482
rect 1317 1481 1318 1487
rect 1324 1483 1330 1491
rect 1324 1482 2527 1483
rect 1324 1478 1327 1482
rect 1331 1478 1351 1482
rect 1355 1478 1423 1482
rect 1427 1478 1519 1482
rect 1523 1478 1527 1482
rect 1531 1478 1615 1482
rect 1619 1478 1631 1482
rect 1635 1478 1711 1482
rect 1715 1478 1735 1482
rect 1739 1478 1815 1482
rect 1819 1478 1839 1482
rect 1843 1478 1927 1482
rect 1931 1478 1943 1482
rect 1947 1478 2039 1482
rect 2043 1478 2047 1482
rect 2051 1478 2135 1482
rect 2139 1478 2175 1482
rect 2179 1478 2231 1482
rect 2235 1478 2303 1482
rect 2307 1478 2327 1482
rect 2331 1478 2423 1482
rect 2427 1478 2439 1482
rect 2443 1478 2503 1482
rect 2507 1478 2527 1482
rect 1324 1477 2527 1478
rect 2533 1477 2534 1483
rect 84 1429 85 1435
rect 91 1434 1299 1435
rect 91 1430 111 1434
rect 115 1430 231 1434
rect 235 1430 319 1434
rect 323 1430 359 1434
rect 363 1430 415 1434
rect 419 1430 447 1434
rect 451 1430 511 1434
rect 515 1430 543 1434
rect 547 1430 615 1434
rect 619 1430 639 1434
rect 643 1430 711 1434
rect 715 1430 735 1434
rect 739 1430 807 1434
rect 811 1430 839 1434
rect 843 1430 895 1434
rect 899 1430 943 1434
rect 947 1430 991 1434
rect 995 1430 1047 1434
rect 1051 1430 1087 1434
rect 1091 1430 1151 1434
rect 1155 1430 1287 1434
rect 1291 1430 1299 1434
rect 91 1429 1299 1430
rect 1305 1429 1306 1435
rect 1310 1421 1311 1427
rect 1317 1426 2539 1427
rect 1317 1422 1327 1426
rect 1331 1422 1367 1426
rect 1371 1422 1423 1426
rect 1427 1422 1439 1426
rect 1443 1422 1503 1426
rect 1507 1422 1535 1426
rect 1539 1422 1591 1426
rect 1595 1422 1631 1426
rect 1635 1422 1679 1426
rect 1683 1422 1727 1426
rect 1731 1422 1775 1426
rect 1779 1422 1831 1426
rect 1835 1422 1879 1426
rect 1883 1422 1943 1426
rect 1947 1422 1991 1426
rect 1995 1422 2063 1426
rect 2067 1422 2111 1426
rect 2115 1422 2191 1426
rect 2195 1422 2231 1426
rect 2235 1422 2319 1426
rect 2323 1422 2351 1426
rect 2355 1422 2455 1426
rect 2459 1422 2503 1426
rect 2507 1422 2539 1426
rect 1317 1421 2539 1422
rect 2545 1421 2546 1427
rect 96 1377 97 1383
rect 103 1382 1311 1383
rect 103 1378 111 1382
rect 115 1378 151 1382
rect 155 1378 215 1382
rect 219 1378 247 1382
rect 251 1378 311 1382
rect 315 1378 335 1382
rect 339 1378 407 1382
rect 411 1378 431 1382
rect 435 1378 511 1382
rect 515 1378 527 1382
rect 531 1378 607 1382
rect 611 1378 631 1382
rect 635 1378 703 1382
rect 707 1378 727 1382
rect 731 1378 799 1382
rect 803 1378 823 1382
rect 827 1378 895 1382
rect 899 1378 911 1382
rect 915 1378 999 1382
rect 1003 1378 1007 1382
rect 1011 1378 1103 1382
rect 1107 1378 1287 1382
rect 1291 1378 1311 1382
rect 103 1377 1311 1378
rect 1317 1377 1318 1383
rect 1298 1365 1299 1371
rect 1305 1370 2527 1371
rect 1305 1366 1327 1370
rect 1331 1366 1351 1370
rect 1355 1366 1407 1370
rect 1411 1366 1479 1370
rect 1483 1366 1487 1370
rect 1491 1366 1567 1370
rect 1571 1366 1575 1370
rect 1579 1366 1655 1370
rect 1659 1366 1663 1370
rect 1667 1366 1751 1370
rect 1755 1366 1759 1370
rect 1763 1366 1855 1370
rect 1859 1366 1863 1370
rect 1867 1366 1967 1370
rect 1971 1366 1975 1370
rect 1979 1366 2079 1370
rect 2083 1366 2095 1370
rect 2099 1366 2199 1370
rect 2203 1366 2215 1370
rect 2219 1366 2327 1370
rect 2331 1366 2335 1370
rect 2339 1366 2439 1370
rect 2443 1366 2503 1370
rect 2507 1366 2527 1370
rect 1305 1365 2527 1366
rect 2533 1365 2534 1371
rect 84 1325 85 1331
rect 91 1330 1299 1331
rect 91 1326 111 1330
rect 115 1326 135 1330
rect 139 1326 199 1330
rect 203 1326 215 1330
rect 219 1326 295 1330
rect 299 1326 319 1330
rect 323 1326 391 1330
rect 395 1326 415 1330
rect 419 1326 495 1330
rect 499 1326 511 1330
rect 515 1326 591 1330
rect 595 1326 599 1330
rect 603 1326 687 1330
rect 691 1326 783 1330
rect 787 1326 879 1330
rect 883 1326 983 1330
rect 987 1326 1287 1330
rect 1291 1326 1299 1330
rect 91 1325 1299 1326
rect 1305 1325 1306 1331
rect 1310 1305 1311 1311
rect 1317 1310 2539 1311
rect 1317 1306 1327 1310
rect 1331 1306 1367 1310
rect 1371 1306 1423 1310
rect 1427 1306 1495 1310
rect 1499 1306 1519 1310
rect 1523 1306 1583 1310
rect 1587 1306 1615 1310
rect 1619 1306 1671 1310
rect 1675 1306 1719 1310
rect 1723 1306 1767 1310
rect 1771 1306 1823 1310
rect 1827 1306 1871 1310
rect 1875 1306 1919 1310
rect 1923 1306 1983 1310
rect 1987 1306 2015 1310
rect 2019 1306 2095 1310
rect 2099 1306 2103 1310
rect 2107 1306 2183 1310
rect 2187 1306 2215 1310
rect 2219 1306 2255 1310
rect 2259 1306 2327 1310
rect 2331 1306 2343 1310
rect 2347 1306 2399 1310
rect 2403 1306 2455 1310
rect 2459 1306 2503 1310
rect 2507 1306 2539 1310
rect 1317 1305 2539 1306
rect 2545 1305 2546 1311
rect 96 1273 97 1279
rect 103 1278 1311 1279
rect 103 1274 111 1278
rect 115 1274 151 1278
rect 155 1274 191 1278
rect 195 1274 231 1278
rect 235 1274 247 1278
rect 251 1274 303 1278
rect 307 1274 335 1278
rect 339 1274 367 1278
rect 371 1274 431 1278
rect 435 1274 439 1278
rect 443 1274 527 1278
rect 531 1274 615 1278
rect 619 1274 639 1278
rect 643 1274 703 1278
rect 707 1274 775 1278
rect 779 1274 799 1278
rect 803 1274 895 1278
rect 899 1274 927 1278
rect 931 1274 1095 1278
rect 1099 1274 1239 1278
rect 1243 1274 1287 1278
rect 1291 1274 1311 1278
rect 103 1273 1311 1274
rect 1317 1273 1318 1279
rect 1298 1237 1299 1243
rect 1305 1242 2527 1243
rect 1305 1238 1327 1242
rect 1331 1238 1351 1242
rect 1355 1238 1407 1242
rect 1411 1238 1447 1242
rect 1451 1238 1503 1242
rect 1507 1238 1575 1242
rect 1579 1238 1599 1242
rect 1603 1238 1695 1242
rect 1699 1238 1703 1242
rect 1707 1238 1807 1242
rect 1811 1238 1815 1242
rect 1819 1238 1903 1242
rect 1907 1238 1927 1242
rect 1931 1238 1999 1242
rect 2003 1238 2031 1242
rect 2035 1238 2087 1242
rect 2091 1238 2127 1242
rect 2131 1238 2167 1242
rect 2171 1238 2215 1242
rect 2219 1238 2239 1242
rect 2243 1238 2295 1242
rect 2299 1238 2311 1242
rect 2315 1238 2375 1242
rect 2379 1238 2383 1242
rect 2387 1238 2439 1242
rect 2443 1238 2503 1242
rect 2507 1238 2527 1242
rect 1305 1237 2527 1238
rect 2533 1237 2534 1243
rect 84 1221 85 1227
rect 91 1226 1299 1227
rect 91 1222 111 1226
rect 115 1222 175 1226
rect 179 1222 231 1226
rect 235 1222 287 1226
rect 291 1222 351 1226
rect 355 1222 407 1226
rect 411 1222 423 1226
rect 427 1222 463 1226
rect 467 1222 511 1226
rect 515 1222 519 1226
rect 523 1222 575 1226
rect 579 1222 623 1226
rect 627 1222 631 1226
rect 635 1222 687 1226
rect 691 1222 743 1226
rect 747 1222 759 1226
rect 763 1222 799 1226
rect 803 1222 855 1226
rect 859 1222 911 1226
rect 915 1222 1079 1226
rect 1083 1222 1223 1226
rect 1227 1222 1287 1226
rect 1291 1222 1299 1226
rect 91 1221 1299 1222
rect 1305 1221 1306 1227
rect 1310 1185 1311 1191
rect 1317 1190 2539 1191
rect 1317 1186 1327 1190
rect 1331 1186 1367 1190
rect 1371 1186 1463 1190
rect 1467 1186 1471 1190
rect 1475 1186 1591 1190
rect 1595 1186 1599 1190
rect 1603 1186 1711 1190
rect 1715 1186 1735 1190
rect 1739 1186 1831 1190
rect 1835 1186 1863 1190
rect 1867 1186 1943 1190
rect 1947 1186 1983 1190
rect 1987 1186 2047 1190
rect 2051 1186 2087 1190
rect 2091 1186 2143 1190
rect 2147 1186 2191 1190
rect 2195 1186 2231 1190
rect 2235 1186 2287 1190
rect 2291 1186 2311 1190
rect 2315 1186 2383 1190
rect 2387 1186 2391 1190
rect 2395 1186 2455 1190
rect 2459 1186 2503 1190
rect 2507 1186 2539 1190
rect 1317 1185 2539 1186
rect 2545 1185 2546 1191
rect 96 1165 97 1171
rect 103 1170 1311 1171
rect 103 1166 111 1170
rect 115 1166 367 1170
rect 371 1166 423 1170
rect 427 1166 479 1170
rect 483 1166 535 1170
rect 539 1166 591 1170
rect 595 1166 647 1170
rect 651 1166 703 1170
rect 707 1166 759 1170
rect 763 1166 815 1170
rect 819 1166 871 1170
rect 875 1166 927 1170
rect 931 1166 983 1170
rect 987 1166 1287 1170
rect 1291 1166 1311 1170
rect 103 1165 1311 1166
rect 1317 1165 1318 1171
rect 1298 1129 1299 1135
rect 1305 1134 2527 1135
rect 1305 1130 1327 1134
rect 1331 1130 1351 1134
rect 1355 1130 1367 1134
rect 1371 1130 1447 1134
rect 1451 1130 1455 1134
rect 1459 1130 1535 1134
rect 1539 1130 1583 1134
rect 1587 1130 1631 1134
rect 1635 1130 1719 1134
rect 1723 1130 1807 1134
rect 1811 1130 1847 1134
rect 1851 1130 1895 1134
rect 1899 1130 1967 1134
rect 1971 1130 1983 1134
rect 1987 1130 2071 1134
rect 2075 1130 2159 1134
rect 2163 1130 2175 1134
rect 2179 1130 2255 1134
rect 2259 1130 2271 1134
rect 2275 1130 2359 1134
rect 2363 1130 2367 1134
rect 2371 1130 2439 1134
rect 2443 1130 2503 1134
rect 2507 1130 2527 1134
rect 1305 1129 2527 1130
rect 2533 1129 2534 1135
rect 84 1109 85 1115
rect 91 1114 1299 1115
rect 91 1110 111 1114
rect 115 1110 223 1114
rect 227 1110 311 1114
rect 315 1110 399 1114
rect 403 1110 407 1114
rect 411 1110 463 1114
rect 467 1110 495 1114
rect 499 1110 519 1114
rect 523 1110 575 1114
rect 579 1110 591 1114
rect 595 1110 631 1114
rect 635 1110 679 1114
rect 683 1110 687 1114
rect 691 1110 743 1114
rect 747 1110 767 1114
rect 771 1110 799 1114
rect 803 1110 847 1114
rect 851 1110 855 1114
rect 859 1110 911 1114
rect 915 1110 927 1114
rect 931 1110 967 1114
rect 971 1110 1015 1114
rect 1019 1110 1103 1114
rect 1107 1110 1287 1114
rect 1291 1110 1299 1114
rect 91 1109 1299 1110
rect 1305 1109 1306 1115
rect 1310 1069 1311 1075
rect 1317 1074 2539 1075
rect 1317 1070 1327 1074
rect 1331 1070 1383 1074
rect 1387 1070 1431 1074
rect 1435 1070 1463 1074
rect 1467 1070 1495 1074
rect 1499 1070 1551 1074
rect 1555 1070 1567 1074
rect 1571 1070 1639 1074
rect 1643 1070 1647 1074
rect 1651 1070 1703 1074
rect 1707 1070 1735 1074
rect 1739 1070 1767 1074
rect 1771 1070 1823 1074
rect 1827 1070 1839 1074
rect 1843 1070 1911 1074
rect 1915 1070 1919 1074
rect 1923 1070 1999 1074
rect 2003 1070 2007 1074
rect 2011 1070 2087 1074
rect 2091 1070 2111 1074
rect 2115 1070 2175 1074
rect 2179 1070 2231 1074
rect 2235 1070 2271 1074
rect 2275 1070 2351 1074
rect 2355 1070 2375 1074
rect 2379 1070 2455 1074
rect 2459 1070 2503 1074
rect 2507 1070 2539 1074
rect 1317 1069 2539 1070
rect 2545 1069 2546 1075
rect 96 1053 97 1059
rect 103 1058 1311 1059
rect 103 1054 111 1058
rect 115 1054 151 1058
rect 155 1054 207 1058
rect 211 1054 239 1058
rect 243 1054 303 1058
rect 307 1054 327 1058
rect 331 1054 415 1058
rect 419 1054 511 1058
rect 515 1054 535 1058
rect 539 1054 607 1058
rect 611 1054 655 1058
rect 659 1054 695 1058
rect 699 1054 767 1058
rect 771 1054 783 1058
rect 787 1054 863 1058
rect 867 1054 879 1058
rect 883 1054 943 1058
rect 947 1054 983 1058
rect 987 1054 1031 1058
rect 1035 1054 1095 1058
rect 1099 1054 1119 1058
rect 1123 1054 1207 1058
rect 1211 1054 1287 1058
rect 1291 1054 1311 1058
rect 103 1053 1311 1054
rect 1317 1053 1318 1059
rect 1298 1009 1299 1015
rect 1305 1014 2527 1015
rect 1305 1010 1327 1014
rect 1331 1010 1415 1014
rect 1419 1010 1479 1014
rect 1483 1010 1511 1014
rect 1515 1010 1551 1014
rect 1555 1010 1567 1014
rect 1571 1010 1623 1014
rect 1627 1010 1679 1014
rect 1683 1010 1687 1014
rect 1691 1010 1735 1014
rect 1739 1010 1751 1014
rect 1755 1010 1807 1014
rect 1811 1010 1823 1014
rect 1827 1010 1887 1014
rect 1891 1010 1903 1014
rect 1907 1010 1983 1014
rect 1987 1010 1991 1014
rect 1995 1010 2095 1014
rect 2099 1010 2215 1014
rect 2219 1010 2335 1014
rect 2339 1010 2439 1014
rect 2443 1010 2503 1014
rect 2507 1010 2527 1014
rect 1305 1009 2527 1010
rect 2533 1009 2534 1015
rect 84 997 85 1003
rect 91 1002 1299 1003
rect 91 998 111 1002
rect 115 998 135 1002
rect 139 998 191 1002
rect 195 998 215 1002
rect 219 998 287 1002
rect 291 998 327 1002
rect 331 998 399 1002
rect 403 998 439 1002
rect 443 998 519 1002
rect 523 998 551 1002
rect 555 998 639 1002
rect 643 998 663 1002
rect 667 998 751 1002
rect 755 998 759 1002
rect 763 998 847 1002
rect 851 998 863 1002
rect 867 998 935 1002
rect 939 998 967 1002
rect 971 998 1015 1002
rect 1019 998 1079 1002
rect 1083 998 1087 1002
rect 1091 998 1167 1002
rect 1171 998 1191 1002
rect 1195 998 1223 1002
rect 1227 998 1287 1002
rect 1291 998 1299 1002
rect 91 997 1299 998
rect 1305 997 1306 1003
rect 96 945 97 951
rect 103 950 1311 951
rect 103 946 111 950
rect 115 946 151 950
rect 155 946 207 950
rect 211 946 231 950
rect 235 946 295 950
rect 299 946 343 950
rect 347 946 399 950
rect 403 946 455 950
rect 459 946 511 950
rect 515 946 567 950
rect 571 946 623 950
rect 627 946 679 950
rect 683 946 735 950
rect 739 946 775 950
rect 779 946 831 950
rect 835 946 863 950
rect 867 946 927 950
rect 931 946 951 950
rect 955 946 1015 950
rect 1019 946 1031 950
rect 1035 946 1095 950
rect 1099 946 1103 950
rect 1107 946 1175 950
rect 1179 946 1183 950
rect 1187 946 1239 950
rect 1243 946 1287 950
rect 1291 946 1311 950
rect 103 945 1311 946
rect 1317 947 1318 951
rect 1317 946 2546 947
rect 1317 945 1327 946
rect 1310 942 1327 945
rect 1331 942 1367 946
rect 1371 942 1439 946
rect 1443 942 1527 946
rect 1531 942 1583 946
rect 1587 942 1615 946
rect 1619 942 1639 946
rect 1643 942 1695 946
rect 1699 942 1751 946
rect 1755 942 1791 946
rect 1795 942 1823 946
rect 1827 942 1895 946
rect 1899 942 1903 946
rect 1907 942 1999 946
rect 2003 942 2015 946
rect 2019 942 2111 946
rect 2115 942 2151 946
rect 2155 942 2231 946
rect 2235 942 2295 946
rect 2299 942 2351 946
rect 2355 942 2439 946
rect 2443 942 2455 946
rect 2459 942 2503 946
rect 2507 942 2546 946
rect 1310 941 2546 942
rect 84 889 85 895
rect 91 894 1299 895
rect 91 890 111 894
rect 115 890 135 894
rect 139 890 191 894
rect 195 890 247 894
rect 251 890 279 894
rect 283 890 343 894
rect 347 890 383 894
rect 387 890 439 894
rect 443 890 495 894
rect 499 890 543 894
rect 547 890 607 894
rect 611 890 647 894
rect 651 890 719 894
rect 723 890 743 894
rect 747 890 815 894
rect 819 890 839 894
rect 843 890 911 894
rect 915 890 927 894
rect 931 890 999 894
rect 1003 890 1007 894
rect 1011 890 1079 894
rect 1083 890 1087 894
rect 1091 890 1159 894
rect 1163 890 1167 894
rect 1171 890 1223 894
rect 1227 890 1287 894
rect 1291 890 1299 894
rect 91 889 1299 890
rect 1305 889 1306 895
rect 1298 887 1306 889
rect 1298 881 1299 887
rect 1305 886 2527 887
rect 1305 882 1327 886
rect 1331 882 1351 886
rect 1355 882 1423 886
rect 1427 882 1487 886
rect 1491 882 1511 886
rect 1515 882 1559 886
rect 1563 882 1599 886
rect 1603 882 1623 886
rect 1627 882 1679 886
rect 1683 882 1687 886
rect 1691 882 1751 886
rect 1755 882 1775 886
rect 1779 882 1815 886
rect 1819 882 1879 886
rect 1883 882 1887 886
rect 1891 882 1975 886
rect 1979 882 1999 886
rect 2003 882 2079 886
rect 2083 882 2135 886
rect 2139 882 2199 886
rect 2203 882 2279 886
rect 2283 882 2319 886
rect 2323 882 2423 886
rect 2427 882 2439 886
rect 2443 882 2503 886
rect 2507 882 2527 886
rect 1305 881 2527 882
rect 2533 881 2534 887
rect 96 833 97 839
rect 103 838 1311 839
rect 103 834 111 838
rect 115 834 239 838
rect 243 834 263 838
rect 267 834 303 838
rect 307 834 359 838
rect 363 834 383 838
rect 387 834 455 838
rect 459 834 463 838
rect 467 834 551 838
rect 555 834 559 838
rect 563 834 639 838
rect 643 834 663 838
rect 667 834 727 838
rect 731 834 759 838
rect 763 834 807 838
rect 811 834 855 838
rect 859 834 895 838
rect 899 834 943 838
rect 947 834 983 838
rect 987 834 1023 838
rect 1027 834 1071 838
rect 1075 834 1103 838
rect 1107 834 1183 838
rect 1187 834 1239 838
rect 1243 834 1287 838
rect 1291 834 1311 838
rect 103 833 1311 834
rect 1317 833 1318 839
rect 1310 821 1311 827
rect 1317 826 2539 827
rect 1317 822 1327 826
rect 1331 822 1439 826
rect 1443 822 1503 826
rect 1507 822 1511 826
rect 1515 822 1575 826
rect 1579 822 1591 826
rect 1595 822 1639 826
rect 1643 822 1671 826
rect 1675 822 1703 826
rect 1707 822 1759 826
rect 1763 822 1767 826
rect 1771 822 1831 826
rect 1835 822 1847 826
rect 1851 822 1903 826
rect 1907 822 1935 826
rect 1939 822 1991 826
rect 1995 822 2023 826
rect 2027 822 2095 826
rect 2099 822 2111 826
rect 2115 822 2199 826
rect 2203 822 2215 826
rect 2219 822 2287 826
rect 2291 822 2335 826
rect 2339 822 2383 826
rect 2387 822 2455 826
rect 2459 822 2503 826
rect 2507 822 2539 826
rect 1317 821 2539 822
rect 2545 821 2546 827
rect 84 777 85 783
rect 91 782 1299 783
rect 91 778 111 782
rect 115 778 151 782
rect 155 778 223 782
rect 227 778 247 782
rect 251 778 287 782
rect 291 778 343 782
rect 347 778 367 782
rect 371 778 439 782
rect 443 778 447 782
rect 451 778 527 782
rect 531 778 535 782
rect 539 778 607 782
rect 611 778 623 782
rect 627 778 679 782
rect 683 778 711 782
rect 715 778 751 782
rect 755 778 791 782
rect 795 778 823 782
rect 827 778 879 782
rect 883 778 895 782
rect 899 778 967 782
rect 971 778 975 782
rect 979 778 1055 782
rect 1059 778 1287 782
rect 1291 778 1299 782
rect 91 777 1299 778
rect 1305 777 1306 783
rect 1298 765 1299 771
rect 1305 770 2527 771
rect 1305 766 1327 770
rect 1331 766 1351 770
rect 1355 766 1423 770
rect 1427 766 1447 770
rect 1451 766 1495 770
rect 1499 766 1567 770
rect 1571 766 1575 770
rect 1579 766 1655 770
rect 1659 766 1687 770
rect 1691 766 1743 770
rect 1747 766 1807 770
rect 1811 766 1831 770
rect 1835 766 1919 770
rect 1923 766 1927 770
rect 1931 766 2007 770
rect 2011 766 2039 770
rect 2043 766 2095 770
rect 2099 766 2143 770
rect 2147 766 2183 770
rect 2187 766 2247 770
rect 2251 766 2271 770
rect 2275 766 2351 770
rect 2355 766 2367 770
rect 2371 766 2439 770
rect 2443 766 2503 770
rect 2507 766 2527 770
rect 1305 765 2527 766
rect 2533 765 2534 771
rect 96 721 97 727
rect 103 726 1311 727
rect 103 722 111 726
rect 115 722 167 726
rect 171 722 175 726
rect 179 722 263 726
rect 267 722 343 726
rect 347 722 359 726
rect 363 722 423 726
rect 427 722 455 726
rect 459 722 503 726
rect 507 722 543 726
rect 547 722 575 726
rect 579 722 623 726
rect 627 722 639 726
rect 643 722 695 726
rect 699 722 703 726
rect 707 722 767 726
rect 771 722 839 726
rect 843 722 911 726
rect 915 722 991 726
rect 995 722 1287 726
rect 1291 722 1311 726
rect 103 721 1311 722
rect 1317 721 1318 727
rect 1310 709 1311 715
rect 1317 714 2539 715
rect 1317 710 1327 714
rect 1331 710 1367 714
rect 1371 710 1431 714
rect 1435 710 1463 714
rect 1467 710 1535 714
rect 1539 710 1583 714
rect 1587 710 1639 714
rect 1643 710 1703 714
rect 1707 710 1751 714
rect 1755 710 1823 714
rect 1827 710 1863 714
rect 1867 710 1943 714
rect 1947 710 1967 714
rect 1971 710 2055 714
rect 2059 710 2063 714
rect 2067 710 2151 714
rect 2155 710 2159 714
rect 2163 710 2231 714
rect 2235 710 2263 714
rect 2267 710 2311 714
rect 2315 710 2367 714
rect 2371 710 2391 714
rect 2395 710 2455 714
rect 2459 710 2503 714
rect 2507 710 2539 714
rect 1317 709 2539 710
rect 2545 709 2546 715
rect 84 669 85 675
rect 91 674 1299 675
rect 91 670 111 674
rect 115 670 159 674
rect 163 670 215 674
rect 219 670 247 674
rect 251 670 295 674
rect 299 670 327 674
rect 331 670 375 674
rect 379 670 407 674
rect 411 670 455 674
rect 459 670 487 674
rect 491 670 527 674
rect 531 670 559 674
rect 563 670 591 674
rect 595 670 623 674
rect 627 670 655 674
rect 659 670 687 674
rect 691 670 719 674
rect 723 670 751 674
rect 755 670 783 674
rect 787 670 823 674
rect 827 670 847 674
rect 851 670 895 674
rect 899 670 919 674
rect 923 670 1287 674
rect 1291 670 1299 674
rect 91 669 1299 670
rect 1305 669 1306 675
rect 1298 649 1299 655
rect 1305 654 2527 655
rect 1305 650 1327 654
rect 1331 650 1351 654
rect 1355 650 1415 654
rect 1419 650 1479 654
rect 1483 650 1519 654
rect 1523 650 1559 654
rect 1563 650 1623 654
rect 1627 650 1647 654
rect 1651 650 1735 654
rect 1739 650 1831 654
rect 1835 650 1847 654
rect 1851 650 1919 654
rect 1923 650 1951 654
rect 1955 650 2007 654
rect 2011 650 2047 654
rect 2051 650 2087 654
rect 2091 650 2135 654
rect 2139 650 2167 654
rect 2171 650 2215 654
rect 2219 650 2239 654
rect 2243 650 2295 654
rect 2299 650 2311 654
rect 2315 650 2375 654
rect 2379 650 2383 654
rect 2387 650 2439 654
rect 2443 650 2503 654
rect 2507 650 2527 654
rect 1305 649 2527 650
rect 2533 649 2534 655
rect 96 613 97 619
rect 103 618 1311 619
rect 103 614 111 618
rect 115 614 207 618
rect 211 614 231 618
rect 235 614 303 618
rect 307 614 311 618
rect 315 614 391 618
rect 395 614 407 618
rect 411 614 471 618
rect 475 614 503 618
rect 507 614 543 618
rect 547 614 599 618
rect 603 614 607 618
rect 611 614 671 618
rect 675 614 687 618
rect 691 614 735 618
rect 739 614 767 618
rect 771 614 799 618
rect 803 614 847 618
rect 851 614 863 618
rect 867 614 927 618
rect 931 614 935 618
rect 939 614 1007 618
rect 1011 614 1087 618
rect 1091 614 1287 618
rect 1291 614 1311 618
rect 103 613 1311 614
rect 1317 613 1318 619
rect 1310 593 1311 599
rect 1317 598 2539 599
rect 1317 594 1327 598
rect 1331 594 1455 598
rect 1459 594 1495 598
rect 1499 594 1559 598
rect 1563 594 1575 598
rect 1579 594 1663 598
rect 1667 594 1671 598
rect 1675 594 1751 598
rect 1755 594 1775 598
rect 1779 594 1847 598
rect 1851 594 1879 598
rect 1883 594 1935 598
rect 1939 594 1983 598
rect 1987 594 2023 598
rect 2027 594 2087 598
rect 2091 594 2103 598
rect 2107 594 2183 598
rect 2187 594 2255 598
rect 2259 594 2279 598
rect 2283 594 2327 598
rect 2331 594 2375 598
rect 2379 594 2399 598
rect 2403 594 2455 598
rect 2459 594 2503 598
rect 2507 594 2539 598
rect 1317 593 2539 594
rect 2545 593 2546 599
rect 84 557 85 563
rect 91 562 1299 563
rect 91 558 111 562
rect 115 558 175 562
rect 179 558 191 562
rect 195 558 271 562
rect 275 558 287 562
rect 291 558 375 562
rect 379 558 391 562
rect 395 558 487 562
rect 491 558 583 562
rect 587 558 591 562
rect 595 558 671 562
rect 675 558 695 562
rect 699 558 751 562
rect 755 558 791 562
rect 795 558 831 562
rect 835 558 879 562
rect 883 558 911 562
rect 915 558 967 562
rect 971 558 991 562
rect 995 558 1055 562
rect 1059 558 1071 562
rect 1075 558 1151 562
rect 1155 558 1287 562
rect 1291 558 1299 562
rect 91 557 1299 558
rect 1305 557 1306 563
rect 1298 537 1299 543
rect 1305 542 2527 543
rect 1305 538 1327 542
rect 1331 538 1367 542
rect 1371 538 1439 542
rect 1443 538 1447 542
rect 1451 538 1527 542
rect 1531 538 1543 542
rect 1547 538 1615 542
rect 1619 538 1655 542
rect 1659 538 1711 542
rect 1715 538 1759 542
rect 1763 538 1799 542
rect 1803 538 1863 542
rect 1867 538 1887 542
rect 1891 538 1967 542
rect 1971 538 1975 542
rect 1979 538 2063 542
rect 2067 538 2071 542
rect 2075 538 2151 542
rect 2155 538 2167 542
rect 2171 538 2247 542
rect 2251 538 2263 542
rect 2267 538 2343 542
rect 2347 538 2359 542
rect 2363 538 2439 542
rect 2443 538 2503 542
rect 2507 538 2527 542
rect 1305 537 2527 538
rect 2533 537 2534 543
rect 96 501 97 507
rect 103 506 1311 507
rect 103 502 111 506
rect 115 502 151 506
rect 155 502 191 506
rect 195 502 247 506
rect 251 502 287 506
rect 291 502 367 506
rect 371 502 391 506
rect 395 502 487 506
rect 491 502 503 506
rect 507 502 607 506
rect 611 502 615 506
rect 619 502 711 506
rect 715 502 735 506
rect 739 502 807 506
rect 811 502 847 506
rect 851 502 895 506
rect 899 502 951 506
rect 955 502 983 506
rect 987 502 1055 506
rect 1059 502 1071 506
rect 1075 502 1159 506
rect 1163 502 1167 506
rect 1171 502 1239 506
rect 1243 502 1287 506
rect 1291 502 1311 506
rect 103 501 1311 502
rect 1317 501 1318 507
rect 1310 481 1311 487
rect 1317 486 2539 487
rect 1317 482 1327 486
rect 1331 482 1367 486
rect 1371 482 1383 486
rect 1387 482 1431 486
rect 1435 482 1463 486
rect 1467 482 1519 486
rect 1523 482 1543 486
rect 1547 482 1615 486
rect 1619 482 1631 486
rect 1635 482 1711 486
rect 1715 482 1727 486
rect 1731 482 1815 486
rect 1819 482 1903 486
rect 1907 482 1927 486
rect 1931 482 1991 486
rect 1995 482 2055 486
rect 2059 482 2079 486
rect 2083 482 2167 486
rect 2171 482 2191 486
rect 2195 482 2263 486
rect 2267 482 2335 486
rect 2339 482 2359 486
rect 2363 482 2455 486
rect 2459 482 2503 486
rect 2507 482 2539 486
rect 1317 481 2539 482
rect 2545 481 2546 487
rect 84 445 85 451
rect 91 450 1299 451
rect 91 446 111 450
rect 115 446 135 450
rect 139 446 191 450
rect 195 446 231 450
rect 235 446 247 450
rect 251 446 303 450
rect 307 446 351 450
rect 355 446 383 450
rect 387 446 471 450
rect 475 446 567 450
rect 571 446 599 450
rect 603 446 671 450
rect 675 446 719 450
rect 723 446 783 450
rect 787 446 831 450
rect 835 446 895 450
rect 899 446 935 450
rect 939 446 1007 450
rect 1011 446 1039 450
rect 1043 446 1127 450
rect 1131 446 1143 450
rect 1147 446 1223 450
rect 1227 446 1287 450
rect 1291 446 1299 450
rect 91 445 1299 446
rect 1305 445 1306 451
rect 1298 425 1299 431
rect 1305 430 2527 431
rect 1305 426 1327 430
rect 1331 426 1351 430
rect 1355 426 1415 430
rect 1419 426 1423 430
rect 1427 426 1503 430
rect 1507 426 1511 430
rect 1515 426 1599 430
rect 1603 426 1679 430
rect 1683 426 1695 430
rect 1699 426 1775 430
rect 1779 426 1799 430
rect 1803 426 1887 430
rect 1891 426 1911 430
rect 1915 426 2015 430
rect 2019 426 2039 430
rect 2043 426 2159 430
rect 2163 426 2175 430
rect 2179 426 2311 430
rect 2315 426 2319 430
rect 2323 426 2439 430
rect 2443 426 2503 430
rect 2507 426 2527 430
rect 1305 425 2527 426
rect 2533 425 2534 431
rect 96 385 97 391
rect 103 390 1311 391
rect 103 386 111 390
rect 115 386 151 390
rect 155 386 207 390
rect 211 386 263 390
rect 267 386 279 390
rect 283 386 319 390
rect 323 386 359 390
rect 363 386 399 390
rect 403 386 431 390
rect 435 386 487 390
rect 491 386 511 390
rect 515 386 583 390
rect 587 386 591 390
rect 595 386 671 390
rect 675 386 687 390
rect 691 386 751 390
rect 755 386 799 390
rect 803 386 823 390
rect 827 386 895 390
rect 899 386 911 390
rect 915 386 967 390
rect 971 386 1023 390
rect 1027 386 1039 390
rect 1043 386 1111 390
rect 1115 386 1143 390
rect 1147 386 1183 390
rect 1187 386 1239 390
rect 1243 386 1287 390
rect 1291 386 1311 390
rect 103 385 1311 386
rect 1317 385 1318 391
rect 1310 369 1311 375
rect 1317 374 2539 375
rect 1317 370 1327 374
rect 1331 370 1367 374
rect 1371 370 1439 374
rect 1443 370 1527 374
rect 1531 370 1615 374
rect 1619 370 1679 374
rect 1683 370 1695 374
rect 1699 370 1735 374
rect 1739 370 1791 374
rect 1795 370 1807 374
rect 1811 370 1903 374
rect 1907 370 2023 374
rect 2027 370 2031 374
rect 2035 370 2159 374
rect 2163 370 2175 374
rect 2179 370 2303 374
rect 2307 370 2327 374
rect 2331 370 2455 374
rect 2459 370 2503 374
rect 2507 370 2539 374
rect 1317 369 2539 370
rect 2545 369 2546 375
rect 84 325 85 331
rect 91 330 1299 331
rect 91 326 111 330
rect 115 326 135 330
rect 139 326 191 330
rect 195 326 199 330
rect 203 326 263 330
rect 267 326 287 330
rect 291 326 343 330
rect 347 326 375 330
rect 379 326 415 330
rect 419 326 455 330
rect 459 326 495 330
rect 499 326 543 330
rect 547 326 575 330
rect 579 326 631 330
rect 635 326 655 330
rect 659 326 727 330
rect 731 326 735 330
rect 739 326 807 330
rect 811 326 823 330
rect 827 326 879 330
rect 883 326 927 330
rect 931 326 951 330
rect 955 326 1023 330
rect 1027 326 1031 330
rect 1035 326 1095 330
rect 1099 326 1135 330
rect 1139 326 1167 330
rect 1171 326 1223 330
rect 1227 326 1287 330
rect 1291 326 1299 330
rect 91 325 1299 326
rect 1305 325 1306 331
rect 1298 323 1306 325
rect 1298 317 1299 323
rect 1305 322 2527 323
rect 1305 318 1327 322
rect 1331 318 1351 322
rect 1355 318 1431 322
rect 1435 318 1527 322
rect 1531 318 1623 322
rect 1627 318 1663 322
rect 1667 318 1711 322
rect 1715 318 1719 322
rect 1723 318 1791 322
rect 1795 318 1807 322
rect 1811 318 1887 322
rect 1891 318 1911 322
rect 1915 318 2007 322
rect 2011 318 2023 322
rect 2027 318 2143 322
rect 2147 318 2151 322
rect 2155 318 2287 322
rect 2291 318 2423 322
rect 2427 318 2439 322
rect 2443 318 2503 322
rect 2507 318 2527 322
rect 1305 317 2527 318
rect 2533 317 2534 323
rect 96 265 97 271
rect 103 270 1311 271
rect 103 266 111 270
rect 115 266 151 270
rect 155 266 215 270
rect 219 266 231 270
rect 235 266 303 270
rect 307 266 327 270
rect 331 266 391 270
rect 395 266 423 270
rect 427 266 471 270
rect 475 266 519 270
rect 523 266 559 270
rect 563 266 615 270
rect 619 266 647 270
rect 651 266 711 270
rect 715 266 743 270
rect 747 266 807 270
rect 811 266 839 270
rect 843 266 903 270
rect 907 266 943 270
rect 947 266 1007 270
rect 1011 266 1047 270
rect 1051 266 1111 270
rect 1115 266 1151 270
rect 1155 266 1215 270
rect 1219 266 1239 270
rect 1243 266 1287 270
rect 1291 266 1311 270
rect 103 265 1311 266
rect 1317 267 1318 271
rect 1317 266 2546 267
rect 1317 265 1327 266
rect 1310 262 1327 265
rect 1331 262 1367 266
rect 1371 262 1439 266
rect 1443 262 1447 266
rect 1451 262 1535 266
rect 1539 262 1543 266
rect 1547 262 1631 266
rect 1635 262 1639 266
rect 1643 262 1727 266
rect 1731 262 1815 266
rect 1819 262 1823 266
rect 1827 262 1903 266
rect 1907 262 1927 266
rect 1931 262 1999 266
rect 2003 262 2039 266
rect 2043 262 2103 266
rect 2107 262 2167 266
rect 2171 262 2215 266
rect 2219 262 2303 266
rect 2307 262 2335 266
rect 2339 262 2439 266
rect 2443 262 2455 266
rect 2459 262 2503 266
rect 2507 262 2546 266
rect 1310 261 2546 262
rect 84 205 85 211
rect 91 210 1299 211
rect 91 206 111 210
rect 115 206 135 210
rect 139 206 159 210
rect 163 206 215 210
rect 219 206 239 210
rect 243 206 311 210
rect 315 206 327 210
rect 331 206 407 210
rect 411 206 415 210
rect 419 206 503 210
rect 507 206 511 210
rect 515 206 599 210
rect 603 206 607 210
rect 611 206 695 210
rect 699 206 783 210
rect 787 206 791 210
rect 795 206 871 210
rect 875 206 887 210
rect 891 206 959 210
rect 963 206 991 210
rect 995 206 1047 210
rect 1051 206 1095 210
rect 1099 206 1135 210
rect 1139 206 1199 210
rect 1203 206 1287 210
rect 1291 206 1299 210
rect 91 205 1299 206
rect 1305 210 2534 211
rect 1305 206 1327 210
rect 1331 206 1351 210
rect 1355 206 1391 210
rect 1395 206 1423 210
rect 1427 206 1495 210
rect 1499 206 1519 210
rect 1523 206 1599 210
rect 1603 206 1615 210
rect 1619 206 1711 210
rect 1715 206 1799 210
rect 1803 206 1815 210
rect 1819 206 1887 210
rect 1891 206 1919 210
rect 1923 206 1983 210
rect 1987 206 2015 210
rect 2019 206 2087 210
rect 2091 206 2111 210
rect 2115 206 2199 210
rect 2203 206 2287 210
rect 2291 206 2319 210
rect 2323 206 2375 210
rect 2379 206 2439 210
rect 2443 206 2503 210
rect 2507 206 2534 210
rect 1305 205 2534 206
rect 96 133 97 139
rect 103 138 1311 139
rect 103 134 111 138
rect 115 134 151 138
rect 155 134 175 138
rect 179 134 207 138
rect 211 134 255 138
rect 259 134 263 138
rect 267 134 319 138
rect 323 134 343 138
rect 347 134 375 138
rect 379 134 431 138
rect 435 134 487 138
rect 491 134 527 138
rect 531 134 551 138
rect 555 134 623 138
rect 627 134 687 138
rect 691 134 711 138
rect 715 134 751 138
rect 755 134 799 138
rect 803 134 815 138
rect 819 134 879 138
rect 883 134 887 138
rect 891 134 943 138
rect 947 134 975 138
rect 979 134 1007 138
rect 1011 134 1063 138
rect 1067 134 1071 138
rect 1075 134 1135 138
rect 1139 134 1151 138
rect 1155 134 1199 138
rect 1203 134 1287 138
rect 1291 134 1311 138
rect 103 133 1311 134
rect 1317 138 2546 139
rect 1317 134 1327 138
rect 1331 134 1367 138
rect 1371 134 1407 138
rect 1411 134 1423 138
rect 1427 134 1479 138
rect 1483 134 1511 138
rect 1515 134 1535 138
rect 1539 134 1591 138
rect 1595 134 1615 138
rect 1619 134 1647 138
rect 1651 134 1703 138
rect 1707 134 1727 138
rect 1731 134 1759 138
rect 1763 134 1815 138
rect 1819 134 1831 138
rect 1835 134 1871 138
rect 1875 134 1927 138
rect 1931 134 1935 138
rect 1939 134 1983 138
rect 1987 134 2031 138
rect 2035 134 2039 138
rect 2043 134 2095 138
rect 2099 134 2127 138
rect 2131 134 2159 138
rect 2163 134 2215 138
rect 2219 134 2223 138
rect 2227 134 2287 138
rect 2291 134 2303 138
rect 2307 134 2343 138
rect 2347 134 2391 138
rect 2395 134 2399 138
rect 2403 134 2455 138
rect 2459 134 2503 138
rect 2507 134 2546 138
rect 1317 133 2546 134
rect 84 81 85 87
rect 91 86 1299 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 191 86
rect 195 82 247 86
rect 251 82 303 86
rect 307 82 359 86
rect 363 82 415 86
rect 419 82 471 86
rect 475 82 535 86
rect 539 82 607 86
rect 611 82 671 86
rect 675 82 735 86
rect 739 82 799 86
rect 803 82 863 86
rect 867 82 927 86
rect 931 82 991 86
rect 995 82 1055 86
rect 1059 82 1119 86
rect 1123 82 1183 86
rect 1187 82 1287 86
rect 1291 82 1299 86
rect 91 81 1299 82
rect 1305 86 2534 87
rect 1305 82 1327 86
rect 1331 82 1351 86
rect 1355 82 1407 86
rect 1411 82 1463 86
rect 1467 82 1519 86
rect 1523 82 1575 86
rect 1579 82 1631 86
rect 1635 82 1687 86
rect 1691 82 1743 86
rect 1747 82 1799 86
rect 1803 82 1855 86
rect 1859 82 1911 86
rect 1915 82 1967 86
rect 1971 82 2023 86
rect 2027 82 2079 86
rect 2083 82 2143 86
rect 2147 82 2207 86
rect 2211 82 2271 86
rect 2275 82 2327 86
rect 2331 82 2383 86
rect 2387 82 2439 86
rect 2443 82 2503 86
rect 2507 82 2534 86
rect 1305 81 2534 82
<< m5c >>
rect 97 2577 103 2583
rect 1311 2577 1317 2583
rect 1311 2553 1317 2559
rect 2539 2553 2545 2559
rect 85 2525 91 2531
rect 1299 2525 1305 2531
rect 1299 2493 1305 2499
rect 2527 2493 2533 2499
rect 97 2473 103 2479
rect 1311 2473 1317 2479
rect 1311 2433 1317 2439
rect 2539 2433 2545 2439
rect 85 2417 91 2423
rect 1299 2417 1305 2423
rect 1299 2375 1305 2381
rect 2527 2373 2533 2379
rect 97 2365 103 2371
rect 1311 2365 1317 2371
rect 1311 2317 1317 2323
rect 2539 2317 2545 2323
rect 85 2309 91 2315
rect 1299 2309 1305 2315
rect 1299 2265 1305 2271
rect 2527 2265 2533 2271
rect 97 2253 103 2259
rect 1311 2253 1317 2259
rect 1311 2209 1317 2215
rect 2539 2209 2545 2215
rect 85 2197 91 2203
rect 1299 2197 1305 2203
rect 1299 2155 1305 2161
rect 97 2145 103 2151
rect 1311 2145 1317 2151
rect 2527 2145 2533 2151
rect 85 2093 91 2099
rect 1299 2093 1305 2099
rect 1311 2081 1317 2087
rect 2539 2081 2545 2087
rect 1299 2047 1305 2053
rect 97 2037 103 2043
rect 1311 2037 1317 2043
rect 2527 2029 2533 2035
rect 85 1981 91 1987
rect 1299 1981 1305 1987
rect 1311 1973 1317 1979
rect 2539 1973 2545 1979
rect 1299 1931 1305 1937
rect 97 1921 103 1927
rect 1311 1921 1317 1927
rect 2527 1917 2533 1923
rect 85 1869 91 1875
rect 1299 1869 1305 1875
rect 1311 1865 1317 1871
rect 2539 1865 2545 1871
rect 1299 1819 1305 1825
rect 97 1809 103 1815
rect 1311 1809 1317 1815
rect 2527 1809 2533 1815
rect 85 1753 91 1759
rect 1299 1753 1305 1759
rect 1311 1753 1317 1759
rect 2539 1753 2545 1759
rect 1299 1707 1305 1713
rect 97 1697 103 1703
rect 1311 1697 1317 1703
rect 2527 1701 2533 1707
rect 85 1645 91 1651
rect 1299 1645 1305 1651
rect 1311 1641 1317 1647
rect 2539 1641 2545 1647
rect 1299 1603 1305 1609
rect 97 1593 103 1599
rect 1311 1593 1317 1599
rect 2527 1585 2533 1591
rect 85 1533 91 1539
rect 1299 1533 1305 1539
rect 1311 1533 1317 1539
rect 2539 1533 2545 1539
rect 1299 1491 1305 1497
rect 97 1481 103 1487
rect 1311 1481 1317 1487
rect 2527 1477 2533 1483
rect 85 1429 91 1435
rect 1299 1429 1305 1435
rect 1311 1421 1317 1427
rect 2539 1421 2545 1427
rect 97 1377 103 1383
rect 1311 1377 1317 1383
rect 1299 1365 1305 1371
rect 2527 1365 2533 1371
rect 85 1325 91 1331
rect 1299 1325 1305 1331
rect 1311 1305 1317 1311
rect 2539 1305 2545 1311
rect 97 1273 103 1279
rect 1311 1273 1317 1279
rect 1299 1237 1305 1243
rect 2527 1237 2533 1243
rect 85 1221 91 1227
rect 1299 1221 1305 1227
rect 1311 1185 1317 1191
rect 2539 1185 2545 1191
rect 97 1165 103 1171
rect 1311 1165 1317 1171
rect 1299 1129 1305 1135
rect 2527 1129 2533 1135
rect 85 1109 91 1115
rect 1299 1109 1305 1115
rect 1311 1069 1317 1075
rect 2539 1069 2545 1075
rect 97 1053 103 1059
rect 1311 1053 1317 1059
rect 1299 1009 1305 1015
rect 2527 1009 2533 1015
rect 85 997 91 1003
rect 1299 997 1305 1003
rect 97 945 103 951
rect 1311 945 1317 951
rect 85 889 91 895
rect 1299 889 1305 895
rect 1299 881 1305 887
rect 2527 881 2533 887
rect 97 833 103 839
rect 1311 833 1317 839
rect 1311 821 1317 827
rect 2539 821 2545 827
rect 85 777 91 783
rect 1299 777 1305 783
rect 1299 765 1305 771
rect 2527 765 2533 771
rect 97 721 103 727
rect 1311 721 1317 727
rect 1311 709 1317 715
rect 2539 709 2545 715
rect 85 669 91 675
rect 1299 669 1305 675
rect 1299 649 1305 655
rect 2527 649 2533 655
rect 97 613 103 619
rect 1311 613 1317 619
rect 1311 593 1317 599
rect 2539 593 2545 599
rect 85 557 91 563
rect 1299 557 1305 563
rect 1299 537 1305 543
rect 2527 537 2533 543
rect 97 501 103 507
rect 1311 501 1317 507
rect 1311 481 1317 487
rect 2539 481 2545 487
rect 85 445 91 451
rect 1299 445 1305 451
rect 1299 425 1305 431
rect 2527 425 2533 431
rect 97 385 103 391
rect 1311 385 1317 391
rect 1311 369 1317 375
rect 2539 369 2545 375
rect 85 325 91 331
rect 1299 325 1305 331
rect 1299 317 1305 323
rect 2527 317 2533 323
rect 97 265 103 271
rect 1311 265 1317 271
rect 85 205 91 211
rect 1299 205 1305 211
rect 97 133 103 139
rect 1311 133 1317 139
rect 85 81 91 87
rect 1299 81 1305 87
<< m5 >>
rect 84 2531 92 2592
rect 84 2525 85 2531
rect 91 2525 92 2531
rect 84 2423 92 2525
rect 84 2417 85 2423
rect 91 2417 92 2423
rect 84 2315 92 2417
rect 84 2309 85 2315
rect 91 2309 92 2315
rect 84 2203 92 2309
rect 84 2197 85 2203
rect 91 2197 92 2203
rect 84 2099 92 2197
rect 84 2093 85 2099
rect 91 2093 92 2099
rect 84 1987 92 2093
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1875 92 1981
rect 84 1869 85 1875
rect 91 1869 92 1875
rect 84 1759 92 1869
rect 84 1753 85 1759
rect 91 1753 92 1759
rect 84 1651 92 1753
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1539 92 1645
rect 84 1533 85 1539
rect 91 1533 92 1539
rect 84 1435 92 1533
rect 84 1429 85 1435
rect 91 1429 92 1435
rect 84 1331 92 1429
rect 84 1325 85 1331
rect 91 1325 92 1331
rect 84 1227 92 1325
rect 84 1221 85 1227
rect 91 1221 92 1227
rect 84 1115 92 1221
rect 84 1109 85 1115
rect 91 1109 92 1115
rect 84 1003 92 1109
rect 84 997 85 1003
rect 91 997 92 1003
rect 84 895 92 997
rect 84 889 85 895
rect 91 889 92 895
rect 84 783 92 889
rect 84 777 85 783
rect 91 777 92 783
rect 84 675 92 777
rect 84 669 85 675
rect 91 669 92 675
rect 84 563 92 669
rect 84 557 85 563
rect 91 557 92 563
rect 84 451 92 557
rect 84 445 85 451
rect 91 445 92 451
rect 84 331 92 445
rect 84 325 85 331
rect 91 325 92 331
rect 84 211 92 325
rect 84 205 85 211
rect 91 205 92 211
rect 84 87 92 205
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2583 104 2592
rect 96 2577 97 2583
rect 103 2577 104 2583
rect 96 2479 104 2577
rect 96 2473 97 2479
rect 103 2473 104 2479
rect 96 2371 104 2473
rect 96 2365 97 2371
rect 103 2365 104 2371
rect 96 2259 104 2365
rect 96 2253 97 2259
rect 103 2253 104 2259
rect 96 2151 104 2253
rect 96 2145 97 2151
rect 103 2145 104 2151
rect 96 2043 104 2145
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1927 104 2037
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1815 104 1921
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1703 104 1809
rect 96 1697 97 1703
rect 103 1697 104 1703
rect 96 1599 104 1697
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1487 104 1593
rect 96 1481 97 1487
rect 103 1481 104 1487
rect 96 1383 104 1481
rect 96 1377 97 1383
rect 103 1377 104 1383
rect 96 1279 104 1377
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1171 104 1273
rect 96 1165 97 1171
rect 103 1165 104 1171
rect 96 1059 104 1165
rect 96 1053 97 1059
rect 103 1053 104 1059
rect 96 951 104 1053
rect 96 945 97 951
rect 103 945 104 951
rect 96 839 104 945
rect 96 833 97 839
rect 103 833 104 839
rect 96 727 104 833
rect 96 721 97 727
rect 103 721 104 727
rect 96 619 104 721
rect 96 613 97 619
rect 103 613 104 619
rect 96 507 104 613
rect 96 501 97 507
rect 103 501 104 507
rect 96 391 104 501
rect 96 385 97 391
rect 103 385 104 391
rect 96 271 104 385
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1298 2531 1306 2592
rect 1298 2525 1299 2531
rect 1305 2525 1306 2531
rect 1298 2499 1306 2525
rect 1298 2493 1299 2499
rect 1305 2493 1306 2499
rect 1298 2423 1306 2493
rect 1298 2417 1299 2423
rect 1305 2417 1306 2423
rect 1298 2381 1306 2417
rect 1298 2375 1299 2381
rect 1305 2375 1306 2381
rect 1298 2315 1306 2375
rect 1298 2309 1299 2315
rect 1305 2309 1306 2315
rect 1298 2271 1306 2309
rect 1298 2265 1299 2271
rect 1305 2265 1306 2271
rect 1298 2203 1306 2265
rect 1298 2197 1299 2203
rect 1305 2197 1306 2203
rect 1298 2161 1306 2197
rect 1298 2155 1299 2161
rect 1305 2155 1306 2161
rect 1298 2099 1306 2155
rect 1298 2093 1299 2099
rect 1305 2093 1306 2099
rect 1298 2053 1306 2093
rect 1298 2047 1299 2053
rect 1305 2047 1306 2053
rect 1298 1987 1306 2047
rect 1298 1981 1299 1987
rect 1305 1981 1306 1987
rect 1298 1937 1306 1981
rect 1298 1931 1299 1937
rect 1305 1931 1306 1937
rect 1298 1875 1306 1931
rect 1298 1869 1299 1875
rect 1305 1869 1306 1875
rect 1298 1825 1306 1869
rect 1298 1819 1299 1825
rect 1305 1819 1306 1825
rect 1298 1759 1306 1819
rect 1298 1753 1299 1759
rect 1305 1753 1306 1759
rect 1298 1713 1306 1753
rect 1298 1707 1299 1713
rect 1305 1707 1306 1713
rect 1298 1651 1306 1707
rect 1298 1645 1299 1651
rect 1305 1645 1306 1651
rect 1298 1609 1306 1645
rect 1298 1603 1299 1609
rect 1305 1603 1306 1609
rect 1298 1539 1306 1603
rect 1298 1533 1299 1539
rect 1305 1533 1306 1539
rect 1298 1497 1306 1533
rect 1298 1491 1299 1497
rect 1305 1491 1306 1497
rect 1298 1435 1306 1491
rect 1298 1429 1299 1435
rect 1305 1429 1306 1435
rect 1298 1371 1306 1429
rect 1298 1365 1299 1371
rect 1305 1365 1306 1371
rect 1298 1331 1306 1365
rect 1298 1325 1299 1331
rect 1305 1325 1306 1331
rect 1298 1243 1306 1325
rect 1298 1237 1299 1243
rect 1305 1237 1306 1243
rect 1298 1227 1306 1237
rect 1298 1221 1299 1227
rect 1305 1221 1306 1227
rect 1298 1135 1306 1221
rect 1298 1129 1299 1135
rect 1305 1129 1306 1135
rect 1298 1115 1306 1129
rect 1298 1109 1299 1115
rect 1305 1109 1306 1115
rect 1298 1015 1306 1109
rect 1298 1009 1299 1015
rect 1305 1009 1306 1015
rect 1298 1003 1306 1009
rect 1298 997 1299 1003
rect 1305 997 1306 1003
rect 1298 895 1306 997
rect 1298 889 1299 895
rect 1305 889 1306 895
rect 1298 887 1306 889
rect 1298 881 1299 887
rect 1305 881 1306 887
rect 1298 783 1306 881
rect 1298 777 1299 783
rect 1305 777 1306 783
rect 1298 771 1306 777
rect 1298 765 1299 771
rect 1305 765 1306 771
rect 1298 675 1306 765
rect 1298 669 1299 675
rect 1305 669 1306 675
rect 1298 655 1306 669
rect 1298 649 1299 655
rect 1305 649 1306 655
rect 1298 563 1306 649
rect 1298 557 1299 563
rect 1305 557 1306 563
rect 1298 543 1306 557
rect 1298 537 1299 543
rect 1305 537 1306 543
rect 1298 451 1306 537
rect 1298 445 1299 451
rect 1305 445 1306 451
rect 1298 431 1306 445
rect 1298 425 1299 431
rect 1305 425 1306 431
rect 1298 331 1306 425
rect 1298 325 1299 331
rect 1305 325 1306 331
rect 1298 323 1306 325
rect 1298 317 1299 323
rect 1305 317 1306 323
rect 1298 211 1306 317
rect 1298 205 1299 211
rect 1305 205 1306 211
rect 1298 87 1306 205
rect 1298 81 1299 87
rect 1305 81 1306 87
rect 1298 72 1306 81
rect 1310 2583 1318 2592
rect 1310 2577 1311 2583
rect 1317 2577 1318 2583
rect 1310 2559 1318 2577
rect 1310 2553 1311 2559
rect 1317 2553 1318 2559
rect 1310 2479 1318 2553
rect 1310 2473 1311 2479
rect 1317 2473 1318 2479
rect 1310 2439 1318 2473
rect 1310 2433 1311 2439
rect 1317 2433 1318 2439
rect 1310 2371 1318 2433
rect 1310 2365 1311 2371
rect 1317 2365 1318 2371
rect 1310 2323 1318 2365
rect 1310 2317 1311 2323
rect 1317 2317 1318 2323
rect 1310 2259 1318 2317
rect 1310 2253 1311 2259
rect 1317 2253 1318 2259
rect 1310 2215 1318 2253
rect 1310 2209 1311 2215
rect 1317 2209 1318 2215
rect 1310 2151 1318 2209
rect 1310 2145 1311 2151
rect 1317 2145 1318 2151
rect 1310 2087 1318 2145
rect 1310 2081 1311 2087
rect 1317 2081 1318 2087
rect 1310 2043 1318 2081
rect 1310 2037 1311 2043
rect 1317 2037 1318 2043
rect 1310 1979 1318 2037
rect 1310 1973 1311 1979
rect 1317 1973 1318 1979
rect 1310 1927 1318 1973
rect 1310 1921 1311 1927
rect 1317 1921 1318 1927
rect 1310 1871 1318 1921
rect 1310 1865 1311 1871
rect 1317 1865 1318 1871
rect 1310 1815 1318 1865
rect 1310 1809 1311 1815
rect 1317 1809 1318 1815
rect 1310 1759 1318 1809
rect 1310 1753 1311 1759
rect 1317 1753 1318 1759
rect 1310 1703 1318 1753
rect 1310 1697 1311 1703
rect 1317 1697 1318 1703
rect 1310 1647 1318 1697
rect 1310 1641 1311 1647
rect 1317 1641 1318 1647
rect 1310 1599 1318 1641
rect 1310 1593 1311 1599
rect 1317 1593 1318 1599
rect 1310 1539 1318 1593
rect 1310 1533 1311 1539
rect 1317 1533 1318 1539
rect 1310 1487 1318 1533
rect 1310 1481 1311 1487
rect 1317 1481 1318 1487
rect 1310 1427 1318 1481
rect 1310 1421 1311 1427
rect 1317 1421 1318 1427
rect 1310 1383 1318 1421
rect 1310 1377 1311 1383
rect 1317 1377 1318 1383
rect 1310 1311 1318 1377
rect 1310 1305 1311 1311
rect 1317 1305 1318 1311
rect 1310 1279 1318 1305
rect 1310 1273 1311 1279
rect 1317 1273 1318 1279
rect 1310 1191 1318 1273
rect 1310 1185 1311 1191
rect 1317 1185 1318 1191
rect 1310 1171 1318 1185
rect 1310 1165 1311 1171
rect 1317 1165 1318 1171
rect 1310 1075 1318 1165
rect 1310 1069 1311 1075
rect 1317 1069 1318 1075
rect 1310 1059 1318 1069
rect 1310 1053 1311 1059
rect 1317 1053 1318 1059
rect 1310 951 1318 1053
rect 1310 945 1311 951
rect 1317 945 1318 951
rect 1310 839 1318 945
rect 1310 833 1311 839
rect 1317 833 1318 839
rect 1310 827 1318 833
rect 1310 821 1311 827
rect 1317 821 1318 827
rect 1310 727 1318 821
rect 1310 721 1311 727
rect 1317 721 1318 727
rect 1310 715 1318 721
rect 1310 709 1311 715
rect 1317 709 1318 715
rect 1310 619 1318 709
rect 1310 613 1311 619
rect 1317 613 1318 619
rect 1310 599 1318 613
rect 1310 593 1311 599
rect 1317 593 1318 599
rect 1310 507 1318 593
rect 1310 501 1311 507
rect 1317 501 1318 507
rect 1310 487 1318 501
rect 1310 481 1311 487
rect 1317 481 1318 487
rect 1310 391 1318 481
rect 1310 385 1311 391
rect 1317 385 1318 391
rect 1310 375 1318 385
rect 1310 369 1311 375
rect 1317 369 1318 375
rect 1310 271 1318 369
rect 1310 265 1311 271
rect 1317 265 1318 271
rect 1310 139 1318 265
rect 1310 133 1311 139
rect 1317 133 1318 139
rect 1310 72 1318 133
rect 2526 2499 2534 2592
rect 2526 2493 2527 2499
rect 2533 2493 2534 2499
rect 2526 2379 2534 2493
rect 2526 2373 2527 2379
rect 2533 2373 2534 2379
rect 2526 2271 2534 2373
rect 2526 2265 2527 2271
rect 2533 2265 2534 2271
rect 2526 2151 2534 2265
rect 2526 2145 2527 2151
rect 2533 2145 2534 2151
rect 2526 2035 2534 2145
rect 2526 2029 2527 2035
rect 2533 2029 2534 2035
rect 2526 1923 2534 2029
rect 2526 1917 2527 1923
rect 2533 1917 2534 1923
rect 2526 1815 2534 1917
rect 2526 1809 2527 1815
rect 2533 1809 2534 1815
rect 2526 1707 2534 1809
rect 2526 1701 2527 1707
rect 2533 1701 2534 1707
rect 2526 1591 2534 1701
rect 2526 1585 2527 1591
rect 2533 1585 2534 1591
rect 2526 1483 2534 1585
rect 2526 1477 2527 1483
rect 2533 1477 2534 1483
rect 2526 1371 2534 1477
rect 2526 1365 2527 1371
rect 2533 1365 2534 1371
rect 2526 1243 2534 1365
rect 2526 1237 2527 1243
rect 2533 1237 2534 1243
rect 2526 1135 2534 1237
rect 2526 1129 2527 1135
rect 2533 1129 2534 1135
rect 2526 1015 2534 1129
rect 2526 1009 2527 1015
rect 2533 1009 2534 1015
rect 2526 887 2534 1009
rect 2526 881 2527 887
rect 2533 881 2534 887
rect 2526 771 2534 881
rect 2526 765 2527 771
rect 2533 765 2534 771
rect 2526 655 2534 765
rect 2526 649 2527 655
rect 2533 649 2534 655
rect 2526 543 2534 649
rect 2526 537 2527 543
rect 2533 537 2534 543
rect 2526 431 2534 537
rect 2526 425 2527 431
rect 2533 425 2534 431
rect 2526 323 2534 425
rect 2526 317 2527 323
rect 2533 317 2534 323
rect 2526 72 2534 317
rect 2538 2559 2546 2592
rect 2538 2553 2539 2559
rect 2545 2553 2546 2559
rect 2538 2439 2546 2553
rect 2538 2433 2539 2439
rect 2545 2433 2546 2439
rect 2538 2323 2546 2433
rect 2538 2317 2539 2323
rect 2545 2317 2546 2323
rect 2538 2215 2546 2317
rect 2538 2209 2539 2215
rect 2545 2209 2546 2215
rect 2538 2087 2546 2209
rect 2538 2081 2539 2087
rect 2545 2081 2546 2087
rect 2538 1979 2546 2081
rect 2538 1973 2539 1979
rect 2545 1973 2546 1979
rect 2538 1871 2546 1973
rect 2538 1865 2539 1871
rect 2545 1865 2546 1871
rect 2538 1759 2546 1865
rect 2538 1753 2539 1759
rect 2545 1753 2546 1759
rect 2538 1647 2546 1753
rect 2538 1641 2539 1647
rect 2545 1641 2546 1647
rect 2538 1539 2546 1641
rect 2538 1533 2539 1539
rect 2545 1533 2546 1539
rect 2538 1427 2546 1533
rect 2538 1421 2539 1427
rect 2545 1421 2546 1427
rect 2538 1311 2546 1421
rect 2538 1305 2539 1311
rect 2545 1305 2546 1311
rect 2538 1191 2546 1305
rect 2538 1185 2539 1191
rect 2545 1185 2546 1191
rect 2538 1075 2546 1185
rect 2538 1069 2539 1075
rect 2545 1069 2546 1075
rect 2538 827 2546 1069
rect 2538 821 2539 827
rect 2545 821 2546 827
rect 2538 715 2546 821
rect 2538 709 2539 715
rect 2545 709 2546 715
rect 2538 599 2546 709
rect 2538 593 2539 599
rect 2545 593 2546 599
rect 2538 487 2546 593
rect 2538 481 2539 487
rect 2545 481 2546 487
rect 2538 375 2546 481
rect 2538 369 2539 375
rect 2545 369 2546 375
rect 2538 72 2546 369
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__175
timestamp 1731220652
transform 1 0 2496 0 1 2508
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220652
transform 1 0 1320 0 1 2508
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220652
transform 1 0 2496 0 -1 2492
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220652
transform 1 0 1320 0 -1 2492
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220652
transform 1 0 2496 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220652
transform 1 0 1320 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220652
transform 1 0 2496 0 -1 2372
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220652
transform 1 0 1320 0 -1 2372
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220652
transform 1 0 2496 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220652
transform 1 0 1320 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220652
transform 1 0 2496 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220652
transform 1 0 1320 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220652
transform 1 0 2496 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220652
transform 1 0 1320 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220652
transform 1 0 2496 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220652
transform 1 0 1320 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220652
transform 1 0 2496 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220652
transform 1 0 1320 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220652
transform 1 0 2496 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220652
transform 1 0 1320 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220652
transform 1 0 2496 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220652
transform 1 0 1320 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220652
transform 1 0 2496 0 -1 1916
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220652
transform 1 0 1320 0 -1 1916
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220652
transform 1 0 2496 0 1 1820
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220652
transform 1 0 1320 0 1 1820
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220652
transform 1 0 2496 0 -1 1808
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220652
transform 1 0 1320 0 -1 1808
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220652
transform 1 0 2496 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220652
transform 1 0 1320 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220652
transform 1 0 2496 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220652
transform 1 0 1320 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220652
transform 1 0 2496 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220652
transform 1 0 1320 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220652
transform 1 0 2496 0 -1 1584
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220652
transform 1 0 1320 0 -1 1584
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220652
transform 1 0 2496 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220652
transform 1 0 1320 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220652
transform 1 0 2496 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220652
transform 1 0 1320 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220652
transform 1 0 2496 0 1 1376
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220652
transform 1 0 1320 0 1 1376
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220652
transform 1 0 2496 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220652
transform 1 0 1320 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220652
transform 1 0 2496 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220652
transform 1 0 1320 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220652
transform 1 0 2496 0 -1 1236
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220652
transform 1 0 1320 0 -1 1236
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220652
transform 1 0 2496 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220652
transform 1 0 1320 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220652
transform 1 0 2496 0 -1 1128
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220652
transform 1 0 1320 0 -1 1128
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220652
transform 1 0 2496 0 1 1024
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220652
transform 1 0 1320 0 1 1024
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220652
transform 1 0 2496 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220652
transform 1 0 1320 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220652
transform 1 0 2496 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220652
transform 1 0 1320 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220652
transform 1 0 2496 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220652
transform 1 0 1320 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220652
transform 1 0 2496 0 1 776
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220652
transform 1 0 1320 0 1 776
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220652
transform 1 0 2496 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220652
transform 1 0 1320 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220652
transform 1 0 2496 0 1 664
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220652
transform 1 0 1320 0 1 664
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220652
transform 1 0 2496 0 -1 648
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220652
transform 1 0 1320 0 -1 648
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220652
transform 1 0 2496 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220652
transform 1 0 1320 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220652
transform 1 0 2496 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220652
transform 1 0 1320 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220652
transform 1 0 2496 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220652
transform 1 0 1320 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220652
transform 1 0 2496 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220652
transform 1 0 1320 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220652
transform 1 0 2496 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220652
transform 1 0 1320 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220652
transform 1 0 2496 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220652
transform 1 0 1320 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220652
transform 1 0 2496 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220652
transform 1 0 1320 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220652
transform 1 0 2496 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220652
transform 1 0 1320 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220652
transform 1 0 2496 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220652
transform 1 0 1320 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220652
transform 1 0 1280 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220652
transform 1 0 104 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220652
transform 1 0 1280 0 -1 2524
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220652
transform 1 0 104 0 -1 2524
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220652
transform 1 0 1280 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220652
transform 1 0 104 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220652
transform 1 0 1280 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220652
transform 1 0 104 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220652
transform 1 0 1280 0 1 2320
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220652
transform 1 0 104 0 1 2320
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220652
transform 1 0 1280 0 -1 2308
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220652
transform 1 0 104 0 -1 2308
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220652
transform 1 0 1280 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220652
transform 1 0 104 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220652
transform 1 0 1280 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220652
transform 1 0 104 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220652
transform 1 0 1280 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220652
transform 1 0 104 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220652
transform 1 0 1280 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220652
transform 1 0 104 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220652
transform 1 0 1280 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220652
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220652
transform 1 0 1280 0 -1 1980
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220652
transform 1 0 104 0 -1 1980
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220652
transform 1 0 1280 0 1 1876
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220652
transform 1 0 104 0 1 1876
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220652
transform 1 0 1280 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220652
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220652
transform 1 0 1280 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220652
transform 1 0 104 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220652
transform 1 0 1280 0 -1 1752
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220652
transform 1 0 104 0 -1 1752
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220652
transform 1 0 1280 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220652
transform 1 0 104 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220652
transform 1 0 1280 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220652
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220652
transform 1 0 1280 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220652
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220652
transform 1 0 1280 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220652
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220652
transform 1 0 1280 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220652
transform 1 0 104 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220652
transform 1 0 1280 0 -1 1428
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220652
transform 1 0 104 0 -1 1428
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220652
transform 1 0 1280 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220652
transform 1 0 104 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220652
transform 1 0 1280 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220652
transform 1 0 104 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220652
transform 1 0 1280 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220652
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220652
transform 1 0 1280 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220652
transform 1 0 104 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220652
transform 1 0 1280 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220652
transform 1 0 104 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220652
transform 1 0 1280 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220652
transform 1 0 104 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220652
transform 1 0 1280 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220652
transform 1 0 104 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220652
transform 1 0 1280 0 -1 996
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220652
transform 1 0 104 0 -1 996
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220652
transform 1 0 1280 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220652
transform 1 0 104 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220652
transform 1 0 1280 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220652
transform 1 0 104 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220652
transform 1 0 1280 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220652
transform 1 0 104 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220652
transform 1 0 1280 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220652
transform 1 0 104 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220652
transform 1 0 1280 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220652
transform 1 0 104 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220652
transform 1 0 1280 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220652
transform 1 0 104 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220652
transform 1 0 1280 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220652
transform 1 0 104 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220652
transform 1 0 1280 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220652
transform 1 0 104 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220652
transform 1 0 1280 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220652
transform 1 0 104 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220652
transform 1 0 1280 0 -1 444
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220652
transform 1 0 104 0 -1 444
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220652
transform 1 0 1280 0 1 340
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220652
transform 1 0 104 0 1 340
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220652
transform 1 0 1280 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220652
transform 1 0 104 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220652
transform 1 0 1280 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220652
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220652
transform 1 0 1280 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220652
transform 1 0 104 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220652
transform 1 0 1280 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220652
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0OR2X1  tst_5999_6
timestamp 1731220652
transform 1 0 2376 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5998_6
timestamp 1731220652
transform 1 0 2432 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5997_6
timestamp 1731220652
transform 1 0 2432 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5996_6
timestamp 1731220652
transform 1 0 2432 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5995_6
timestamp 1731220652
transform 1 0 2416 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5994_6
timestamp 1731220652
transform 1 0 2368 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5993_6
timestamp 1731220652
transform 1 0 2280 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5992_6
timestamp 1731220652
transform 1 0 2320 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5991_6
timestamp 1731220652
transform 1 0 2264 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5990_6
timestamp 1731220652
transform 1 0 2200 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5989_6
timestamp 1731220652
transform 1 0 2136 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5988_6
timestamp 1731220652
transform 1 0 2072 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5987_6
timestamp 1731220652
transform 1 0 2016 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5986_6
timestamp 1731220652
transform 1 0 1960 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5985_6
timestamp 1731220652
transform 1 0 1904 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5984_6
timestamp 1731220652
transform 1 0 1848 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5983_6
timestamp 1731220652
transform 1 0 2192 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5982_6
timestamp 1731220652
transform 1 0 2104 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5981_6
timestamp 1731220652
transform 1 0 2008 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5980_6
timestamp 1731220652
transform 1 0 1912 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5979_6
timestamp 1731220652
transform 1 0 2312 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5978_6
timestamp 1731220652
transform 1 0 2192 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5977_6
timestamp 1731220652
transform 1 0 2080 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5976_6
timestamp 1731220652
transform 1 0 1976 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5975_6
timestamp 1731220652
transform 1 0 1880 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5974_6
timestamp 1731220652
transform 1 0 2280 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5973_6
timestamp 1731220652
transform 1 0 2144 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5972_6
timestamp 1731220652
transform 1 0 2016 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5971_6
timestamp 1731220652
transform 1 0 1904 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5970_6
timestamp 1731220652
transform 1 0 1800 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5969_6
timestamp 1731220652
transform 1 0 2280 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5968_6
timestamp 1731220652
transform 1 0 2136 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5967_6
timestamp 1731220652
transform 1 0 2000 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5966_6
timestamp 1731220652
transform 1 0 1880 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5965_6
timestamp 1731220652
transform 1 0 1784 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5964_6
timestamp 1731220652
transform 1 0 1768 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5963_6
timestamp 1731220652
transform 1 0 1672 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5962_6
timestamp 1731220652
transform 1 0 1880 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5961_6
timestamp 1731220652
transform 1 0 2304 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5960_6
timestamp 1731220652
transform 1 0 2152 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5959_6
timestamp 1731220652
transform 1 0 2008 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5958_6
timestamp 1731220652
transform 1 0 1904 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5957_6
timestamp 1731220652
transform 1 0 1792 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5956_6
timestamp 1731220652
transform 1 0 2032 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5955_6
timestamp 1731220652
transform 1 0 2312 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5954_6
timestamp 1731220652
transform 1 0 2168 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5953_6
timestamp 1731220652
transform 1 0 2056 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5952_6
timestamp 1731220652
transform 1 0 1968 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5951_6
timestamp 1731220652
transform 1 0 1880 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5950_6
timestamp 1731220652
transform 1 0 2240 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5949_6
timestamp 1731220652
transform 1 0 2144 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5948_6
timestamp 1731220652
transform 1 0 2064 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5947_6
timestamp 1731220652
transform 1 0 1960 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5946_6
timestamp 1731220652
transform 1 0 2256 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5945_6
timestamp 1731220652
transform 1 0 2160 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5944_6
timestamp 1731220652
transform 1 0 2080 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5943_6
timestamp 1731220652
transform 1 0 2000 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5942_6
timestamp 1731220652
transform 1 0 2160 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5941_6
timestamp 1731220652
transform 1 0 2208 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5940_6
timestamp 1731220652
transform 1 0 2232 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5939_6
timestamp 1731220652
transform 1 0 2304 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5938_6
timestamp 1731220652
transform 1 0 2376 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5937_6
timestamp 1731220652
transform 1 0 2352 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5936_6
timestamp 1731220652
transform 1 0 2336 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5935_6
timestamp 1731220652
transform 1 0 2432 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5934_6
timestamp 1731220652
transform 1 0 2432 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5933_6
timestamp 1731220652
transform 1 0 2432 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5932_6
timestamp 1731220652
transform 1 0 2432 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5931_6
timestamp 1731220652
transform 1 0 2432 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5930_6
timestamp 1731220652
transform 1 0 2432 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5929_6
timestamp 1731220652
transform 1 0 2432 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5928_6
timestamp 1731220652
transform 1 0 2432 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5927_6
timestamp 1731220652
transform 1 0 2432 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5926_6
timestamp 1731220652
transform 1 0 2432 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5925_6
timestamp 1731220652
transform 1 0 2328 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5924_6
timestamp 1731220652
transform 1 0 2416 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5923_6
timestamp 1731220652
transform 1 0 2360 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5922_6
timestamp 1731220652
transform 1 0 2344 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5921_6
timestamp 1731220652
transform 1 0 2368 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5920_6
timestamp 1731220652
transform 1 0 2288 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5919_6
timestamp 1731220652
transform 1 0 2128 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5918_6
timestamp 1731220652
transform 1 0 2040 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5917_6
timestamp 1731220652
transform 1 0 1944 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5916_6
timestamp 1731220652
transform 1 0 2240 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5915_6
timestamp 1731220652
transform 1 0 2136 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5914_6
timestamp 1731220652
transform 1 0 2032 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5913_6
timestamp 1731220652
transform 1 0 1920 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5912_6
timestamp 1731220652
transform 1 0 2264 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5911_6
timestamp 1731220652
transform 1 0 2176 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5910_6
timestamp 1731220652
transform 1 0 2088 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5909_6
timestamp 1731220652
transform 1 0 2000 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5908_6
timestamp 1731220652
transform 1 0 1912 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5907_6
timestamp 1731220652
transform 1 0 2312 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5906_6
timestamp 1731220652
transform 1 0 2192 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5905_6
timestamp 1731220652
transform 1 0 2072 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5904_6
timestamp 1731220652
transform 1 0 1968 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5903_6
timestamp 1731220652
transform 1 0 1880 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5902_6
timestamp 1731220652
transform 1 0 1808 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5901_6
timestamp 1731220652
transform 1 0 2272 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5900_6
timestamp 1731220652
transform 1 0 2128 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5899_6
timestamp 1731220652
transform 1 0 1992 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5898_6
timestamp 1731220652
transform 1 0 1872 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5897_6
timestamp 1731220652
transform 1 0 1768 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5896_6
timestamp 1731220652
transform 1 0 1728 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5895_6
timestamp 1731220652
transform 1 0 1800 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5894_6
timestamp 1731220652
transform 1 0 1880 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5893_6
timestamp 1731220652
transform 1 0 2208 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5892_6
timestamp 1731220652
transform 1 0 2088 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5891_6
timestamp 1731220652
transform 1 0 1976 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5890_6
timestamp 1731220652
transform 1 0 1984 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5889_6
timestamp 1731220652
transform 1 0 1896 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5888_6
timestamp 1731220652
transform 1 0 1816 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5887_6
timestamp 1731220652
transform 1 0 2328 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5886_6
timestamp 1731220652
transform 1 0 2208 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5885_6
timestamp 1731220652
transform 1 0 2088 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5884_6
timestamp 1731220652
transform 1 0 2064 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5883_6
timestamp 1731220652
transform 1 0 1976 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5882_6
timestamp 1731220652
transform 1 0 1888 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5881_6
timestamp 1731220652
transform 1 0 2352 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5880_6
timestamp 1731220652
transform 1 0 2248 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5879_6
timestamp 1731220652
transform 1 0 2152 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5878_6
timestamp 1731220652
transform 1 0 2064 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5877_6
timestamp 1731220652
transform 1 0 1960 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5876_6
timestamp 1731220652
transform 1 0 2168 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5875_6
timestamp 1731220652
transform 1 0 2264 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5874_6
timestamp 1731220652
transform 1 0 2360 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5873_6
timestamp 1731220652
transform 1 0 2288 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5872_6
timestamp 1731220652
transform 1 0 2208 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5871_6
timestamp 1731220652
transform 1 0 2120 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5870_6
timestamp 1731220652
transform 1 0 2024 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5869_6
timestamp 1731220652
transform 1 0 1920 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5868_6
timestamp 1731220652
transform 1 0 2232 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5867_6
timestamp 1731220652
transform 1 0 2160 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5866_6
timestamp 1731220652
transform 1 0 2080 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5865_6
timestamp 1731220652
transform 1 0 1992 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5864_6
timestamp 1731220652
transform 1 0 1896 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5863_6
timestamp 1731220652
transform 1 0 2192 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5862_6
timestamp 1731220652
transform 1 0 2072 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5861_6
timestamp 1731220652
transform 1 0 1960 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5860_6
timestamp 1731220652
transform 1 0 1848 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5859_6
timestamp 1731220652
transform 1 0 2088 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5858_6
timestamp 1731220652
transform 1 0 1968 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5857_6
timestamp 1731220652
transform 1 0 1856 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5856_6
timestamp 1731220652
transform 1 0 1752 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5855_6
timestamp 1731220652
transform 1 0 1808 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5854_6
timestamp 1731220652
transform 1 0 1920 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5853_6
timestamp 1731220652
transform 1 0 2040 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5852_6
timestamp 1731220652
transform 1 0 2168 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5851_6
timestamp 1731220652
transform 1 0 2032 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5850_6
timestamp 1731220652
transform 1 0 1936 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5849_6
timestamp 1731220652
transform 1 0 2272 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5848_6
timestamp 1731220652
transform 1 0 2224 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5847_6
timestamp 1731220652
transform 1 0 2128 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5846_6
timestamp 1731220652
transform 1 0 2320 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5845_6
timestamp 1731220652
transform 1 0 2296 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5844_6
timestamp 1731220652
transform 1 0 2208 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5843_6
timestamp 1731220652
transform 1 0 2328 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5842_6
timestamp 1731220652
transform 1 0 2320 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5841_6
timestamp 1731220652
transform 1 0 2304 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5840_6
timestamp 1731220652
transform 1 0 2368 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5839_6
timestamp 1731220652
transform 1 0 2432 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5838_6
timestamp 1731220652
transform 1 0 2432 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5837_6
timestamp 1731220652
transform 1 0 2432 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5836_6
timestamp 1731220652
transform 1 0 2432 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5835_6
timestamp 1731220652
transform 1 0 2432 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5834_6
timestamp 1731220652
transform 1 0 2432 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5833_6
timestamp 1731220652
transform 1 0 2376 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5832_6
timestamp 1731220652
transform 1 0 2432 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5831_6
timestamp 1731220652
transform 1 0 2432 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5830_6
timestamp 1731220652
transform 1 0 2432 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5829_6
timestamp 1731220652
transform 1 0 2416 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5828_6
timestamp 1731220652
transform 1 0 2432 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5827_6
timestamp 1731220652
transform 1 0 2432 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5826_6
timestamp 1731220652
transform 1 0 2432 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5825_6
timestamp 1731220652
transform 1 0 2432 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5824_6
timestamp 1731220652
transform 1 0 2432 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5823_6
timestamp 1731220652
transform 1 0 2432 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5822_6
timestamp 1731220652
transform 1 0 2432 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5821_6
timestamp 1731220652
transform 1 0 2432 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5820_6
timestamp 1731220652
transform 1 0 2432 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5819_6
timestamp 1731220652
transform 1 0 2432 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5818_6
timestamp 1731220652
transform 1 0 2320 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5817_6
timestamp 1731220652
transform 1 0 2432 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5816_6
timestamp 1731220652
transform 1 0 2376 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5815_6
timestamp 1731220652
transform 1 0 2320 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5814_6
timestamp 1731220652
transform 1 0 2264 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5813_6
timestamp 1731220652
transform 1 0 2200 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5812_6
timestamp 1731220652
transform 1 0 2136 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5811_6
timestamp 1731220652
transform 1 0 2072 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5810_6
timestamp 1731220652
transform 1 0 2016 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5809_6
timestamp 1731220652
transform 1 0 1960 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5808_6
timestamp 1731220652
transform 1 0 1904 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5807_6
timestamp 1731220652
transform 1 0 2304 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5806_6
timestamp 1731220652
transform 1 0 2208 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5805_6
timestamp 1731220652
transform 1 0 2112 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5804_6
timestamp 1731220652
transform 1 0 2024 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5803_6
timestamp 1731220652
transform 1 0 1928 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5802_6
timestamp 1731220652
transform 1 0 2184 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5801_6
timestamp 1731220652
transform 1 0 2088 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5800_6
timestamp 1731220652
transform 1 0 1992 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5799_6
timestamp 1731220652
transform 1 0 1904 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5798_6
timestamp 1731220652
transform 1 0 1808 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5797_6
timestamp 1731220652
transform 1 0 2088 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5796_6
timestamp 1731220652
transform 1 0 2000 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5795_6
timestamp 1731220652
transform 1 0 1912 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5794_6
timestamp 1731220652
transform 1 0 1824 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5793_6
timestamp 1731220652
transform 1 0 1744 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5792_6
timestamp 1731220652
transform 1 0 1712 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5791_6
timestamp 1731220652
transform 1 0 1800 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5790_6
timestamp 1731220652
transform 1 0 1888 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5789_6
timestamp 1731220652
transform 1 0 1984 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5788_6
timestamp 1731220652
transform 1 0 2080 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5787_6
timestamp 1731220652
transform 1 0 2120 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5786_6
timestamp 1731220652
transform 1 0 2032 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5785_6
timestamp 1731220652
transform 1 0 1944 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5784_6
timestamp 1731220652
transform 1 0 1856 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5783_6
timestamp 1731220652
transform 1 0 1768 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5782_6
timestamp 1731220652
transform 1 0 2160 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5781_6
timestamp 1731220652
transform 1 0 2104 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5780_6
timestamp 1731220652
transform 1 0 2048 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5779_6
timestamp 1731220652
transform 1 0 1992 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5778_6
timestamp 1731220652
transform 1 0 1936 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5777_6
timestamp 1731220652
transform 1 0 1880 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5776_6
timestamp 1731220652
transform 1 0 1824 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5775_6
timestamp 1731220652
transform 1 0 1768 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5774_6
timestamp 1731220652
transform 1 0 1712 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5773_6
timestamp 1731220652
transform 1 0 1656 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5772_6
timestamp 1731220652
transform 1 0 1600 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5771_6
timestamp 1731220652
transform 1 0 1544 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5770_6
timestamp 1731220652
transform 1 0 1488 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5769_6
timestamp 1731220652
transform 1 0 1432 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5768_6
timestamp 1731220652
transform 1 0 1376 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5767_6
timestamp 1731220652
transform 1 0 1680 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5766_6
timestamp 1731220652
transform 1 0 1592 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5765_6
timestamp 1731220652
transform 1 0 1504 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5764_6
timestamp 1731220652
transform 1 0 1416 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5763_6
timestamp 1731220652
transform 1 0 1344 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5762_6
timestamp 1731220652
transform 1 0 1616 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5761_6
timestamp 1731220652
transform 1 0 1520 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5760_6
timestamp 1731220652
transform 1 0 1416 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5759_6
timestamp 1731220652
transform 1 0 1344 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5758_6
timestamp 1731220652
transform 1 0 1344 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5757_6
timestamp 1731220652
transform 1 0 1400 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5756_6
timestamp 1731220652
transform 1 0 1488 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5755_6
timestamp 1731220652
transform 1 0 1664 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5754_6
timestamp 1731220652
transform 1 0 1576 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5753_6
timestamp 1731220652
transform 1 0 1520 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5752_6
timestamp 1731220652
transform 1 0 1432 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5751_6
timestamp 1731220652
transform 1 0 1344 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5750_6
timestamp 1731220652
transform 1 0 1616 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5749_6
timestamp 1731220652
transform 1 0 1712 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5748_6
timestamp 1731220652
transform 1 0 1832 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5747_6
timestamp 1731220652
transform 1 0 1728 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5746_6
timestamp 1731220652
transform 1 0 1632 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5745_6
timestamp 1731220652
transform 1 0 1536 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5744_6
timestamp 1731220652
transform 1 0 1448 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5743_6
timestamp 1731220652
transform 1 0 1544 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5742_6
timestamp 1731220652
transform 1 0 1600 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5741_6
timestamp 1731220652
transform 1 0 1656 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5740_6
timestamp 1731220652
transform 1 0 1720 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5739_6
timestamp 1731220652
transform 1 0 1848 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5738_6
timestamp 1731220652
transform 1 0 1784 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5737_6
timestamp 1731220652
transform 1 0 1784 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5736_6
timestamp 1731220652
transform 1 0 1712 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5735_6
timestamp 1731220652
transform 1 0 1656 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5734_6
timestamp 1731220652
transform 1 0 1864 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5733_6
timestamp 1731220652
transform 1 0 1960 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5732_6
timestamp 1731220652
transform 1 0 2072 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5731_6
timestamp 1731220652
transform 1 0 2192 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5730_6
timestamp 1731220652
transform 1 0 2296 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5729_6
timestamp 1731220652
transform 1 0 2144 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5728_6
timestamp 1731220652
transform 1 0 2000 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5727_6
timestamp 1731220652
transform 1 0 1872 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5726_6
timestamp 1731220652
transform 1 0 1760 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5725_6
timestamp 1731220652
transform 1 0 1816 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5724_6
timestamp 1731220652
transform 1 0 1928 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5723_6
timestamp 1731220652
transform 1 0 2048 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5722_6
timestamp 1731220652
transform 1 0 2312 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5721_6
timestamp 1731220652
transform 1 0 2176 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5720_6
timestamp 1731220652
transform 1 0 2128 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5719_6
timestamp 1731220652
transform 1 0 2024 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5718_6
timestamp 1731220652
transform 1 0 1920 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5717_6
timestamp 1731220652
transform 1 0 2344 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5716_6
timestamp 1731220652
transform 1 0 2232 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5715_6
timestamp 1731220652
transform 1 0 2192 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5714_6
timestamp 1731220652
transform 1 0 2104 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5713_6
timestamp 1731220652
transform 1 0 2008 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5712_6
timestamp 1731220652
transform 1 0 2280 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5711_6
timestamp 1731220652
transform 1 0 2368 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5710_6
timestamp 1731220652
transform 1 0 2432 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5709_6
timestamp 1731220652
transform 1 0 2344 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5708_6
timestamp 1731220652
transform 1 0 2248 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5707_6
timestamp 1731220652
transform 1 0 2152 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5706_6
timestamp 1731220652
transform 1 0 2056 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5705_6
timestamp 1731220652
transform 1 0 2360 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5704_6
timestamp 1731220652
transform 1 0 2264 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5703_6
timestamp 1731220652
transform 1 0 2176 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5702_6
timestamp 1731220652
transform 1 0 2080 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5701_6
timestamp 1731220652
transform 1 0 1976 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5700_6
timestamp 1731220652
transform 1 0 2328 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5699_6
timestamp 1731220652
transform 1 0 2208 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5698_6
timestamp 1731220652
transform 1 0 2088 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5697_6
timestamp 1731220652
transform 1 0 1976 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5696_6
timestamp 1731220652
transform 1 0 1864 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5695_6
timestamp 1731220652
transform 1 0 2304 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5694_6
timestamp 1731220652
transform 1 0 2152 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5693_6
timestamp 1731220652
transform 1 0 2008 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5692_6
timestamp 1731220652
transform 1 0 1872 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5691_6
timestamp 1731220652
transform 1 0 1752 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5690_6
timestamp 1731220652
transform 1 0 2304 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5689_6
timestamp 1731220652
transform 1 0 2160 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5688_6
timestamp 1731220652
transform 1 0 2032 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5687_6
timestamp 1731220652
transform 1 0 1912 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5686_6
timestamp 1731220652
transform 1 0 1816 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5685_6
timestamp 1731220652
transform 1 0 1728 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5684_6
timestamp 1731220652
transform 1 0 1656 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5683_6
timestamp 1731220652
transform 1 0 1576 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5682_6
timestamp 1731220652
transform 1 0 2096 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5681_6
timestamp 1731220652
transform 1 0 1928 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5680_6
timestamp 1731220652
transform 1 0 1776 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5679_6
timestamp 1731220652
transform 1 0 1640 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5678_6
timestamp 1731220652
transform 1 0 1520 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5677_6
timestamp 1731220652
transform 1 0 1832 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5676_6
timestamp 1731220652
transform 1 0 1728 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5675_6
timestamp 1731220652
transform 1 0 1624 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5674_6
timestamp 1731220652
transform 1 0 1608 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5673_6
timestamp 1731220652
transform 1 0 1512 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5672_6
timestamp 1731220652
transform 1 0 1704 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5671_6
timestamp 1731220652
transform 1 0 1656 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5670_6
timestamp 1731220652
transform 1 0 1568 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5669_6
timestamp 1731220652
transform 1 0 1480 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5668_6
timestamp 1731220652
transform 1 0 1560 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5667_6
timestamp 1731220652
transform 1 0 1648 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5666_6
timestamp 1731220652
transform 1 0 1744 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5665_6
timestamp 1731220652
transform 1 0 1696 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5664_6
timestamp 1731220652
transform 1 0 1592 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5663_6
timestamp 1731220652
transform 1 0 1800 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5662_6
timestamp 1731220652
transform 1 0 1808 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5661_6
timestamp 1731220652
transform 1 0 1688 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5660_6
timestamp 1731220652
transform 1 0 1568 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5659_6
timestamp 1731220652
transform 1 0 1712 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5658_6
timestamp 1731220652
transform 1 0 1840 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5657_6
timestamp 1731220652
transform 1 0 1800 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5656_6
timestamp 1731220652
transform 1 0 1712 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5655_6
timestamp 1731220652
transform 1 0 1624 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5654_6
timestamp 1731220652
transform 1 0 1744 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5653_6
timestamp 1731220652
transform 1 0 1680 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5652_6
timestamp 1731220652
transform 1 0 1672 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5651_6
timestamp 1731220652
transform 1 0 1592 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5650_6
timestamp 1731220652
transform 1 0 1672 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5649_6
timestamp 1731220652
transform 1 0 1680 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5648_6
timestamp 1731220652
transform 1 0 1744 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5647_6
timestamp 1731220652
transform 1 0 1824 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5646_6
timestamp 1731220652
transform 1 0 1736 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5645_6
timestamp 1731220652
transform 1 0 1648 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5644_6
timestamp 1731220652
transform 1 0 1680 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5643_6
timestamp 1731220652
transform 1 0 1800 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5642_6
timestamp 1731220652
transform 1 0 1840 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5641_6
timestamp 1731220652
transform 1 0 1728 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5640_6
timestamp 1731220652
transform 1 0 1728 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5639_6
timestamp 1731220652
transform 1 0 1824 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5638_6
timestamp 1731220652
transform 1 0 1912 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5637_6
timestamp 1731220652
transform 1 0 1856 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5636_6
timestamp 1731220652
transform 1 0 1752 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5635_6
timestamp 1731220652
transform 1 0 1792 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5634_6
timestamp 1731220652
transform 1 0 1704 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5633_6
timestamp 1731220652
transform 1 0 1608 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5632_6
timestamp 1731220652
transform 1 0 1688 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5631_6
timestamp 1731220652
transform 1 0 1592 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5630_6
timestamp 1731220652
transform 1 0 1504 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5629_6
timestamp 1731220652
transform 1 0 1592 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5628_6
timestamp 1731220652
transform 1 0 1712 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5627_6
timestamp 1731220652
transform 1 0 1656 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5626_6
timestamp 1731220652
transform 1 0 1616 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5625_6
timestamp 1731220652
transform 1 0 1704 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5624_6
timestamp 1731220652
transform 1 0 1792 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5623_6
timestamp 1731220652
transform 1 0 1704 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5622_6
timestamp 1731220652
transform 1 0 1608 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5621_6
timestamp 1731220652
transform 1 0 1704 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5620_6
timestamp 1731220652
transform 1 0 1808 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5619_6
timestamp 1731220652
transform 1 0 1792 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5618_6
timestamp 1731220652
transform 1 0 1736 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5617_6
timestamp 1731220652
transform 1 0 1680 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5616_6
timestamp 1731220652
transform 1 0 1624 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5615_6
timestamp 1731220652
transform 1 0 1568 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5614_6
timestamp 1731220652
transform 1 0 1512 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5613_6
timestamp 1731220652
transform 1 0 1456 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5612_6
timestamp 1731220652
transform 1 0 1400 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5611_6
timestamp 1731220652
transform 1 0 1344 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5610_6
timestamp 1731220652
transform 1 0 1384 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5609_6
timestamp 1731220652
transform 1 0 1488 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5608_6
timestamp 1731220652
transform 1 0 1592 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5607_6
timestamp 1731220652
transform 1 0 1512 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5606_6
timestamp 1731220652
transform 1 0 1416 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5605_6
timestamp 1731220652
transform 1 0 1344 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5604_6
timestamp 1731220652
transform 1 0 1520 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5603_6
timestamp 1731220652
transform 1 0 1424 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5602_6
timestamp 1731220652
transform 1 0 1344 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5601_6
timestamp 1731220652
transform 1 0 1216 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5600_6
timestamp 1731220652
transform 1 0 1160 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5599_6
timestamp 1731220652
transform 1 0 1216 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5598_6
timestamp 1731220652
transform 1 0 1344 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5597_6
timestamp 1731220652
transform 1 0 1416 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5596_6
timestamp 1731220652
transform 1 0 1496 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5595_6
timestamp 1731220652
transform 1 0 1408 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5594_6
timestamp 1731220652
transform 1 0 1344 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5593_6
timestamp 1731220652
transform 1 0 1360 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5592_6
timestamp 1731220652
transform 1 0 1520 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5591_6
timestamp 1731220652
transform 1 0 1440 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5590_6
timestamp 1731220652
transform 1 0 1432 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5589_6
timestamp 1731220652
transform 1 0 1536 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5588_6
timestamp 1731220652
transform 1 0 1648 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5587_6
timestamp 1731220652
transform 1 0 1640 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5586_6
timestamp 1731220652
transform 1 0 1552 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5585_6
timestamp 1731220652
transform 1 0 1472 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5584_6
timestamp 1731220652
transform 1 0 1616 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5583_6
timestamp 1731220652
transform 1 0 1512 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5582_6
timestamp 1731220652
transform 1 0 1408 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5581_6
timestamp 1731220652
transform 1 0 1344 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5580_6
timestamp 1731220652
transform 1 0 1344 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5579_6
timestamp 1731220652
transform 1 0 1440 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5578_6
timestamp 1731220652
transform 1 0 1560 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5577_6
timestamp 1731220652
transform 1 0 1568 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5576_6
timestamp 1731220652
transform 1 0 1488 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5575_6
timestamp 1731220652
transform 1 0 1416 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5574_6
timestamp 1731220652
transform 1 0 1480 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5573_6
timestamp 1731220652
transform 1 0 1616 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5572_6
timestamp 1731220652
transform 1 0 1552 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5571_6
timestamp 1731220652
transform 1 0 1504 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5570_6
timestamp 1731220652
transform 1 0 1416 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5569_6
timestamp 1731220652
transform 1 0 1504 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5568_6
timestamp 1731220652
transform 1 0 1560 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5567_6
timestamp 1731220652
transform 1 0 1616 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5566_6
timestamp 1731220652
transform 1 0 1616 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5565_6
timestamp 1731220652
transform 1 0 1544 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5564_6
timestamp 1731220652
transform 1 0 1472 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5563_6
timestamp 1731220652
transform 1 0 1408 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5562_6
timestamp 1731220652
transform 1 0 1360 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5561_6
timestamp 1731220652
transform 1 0 1440 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5560_6
timestamp 1731220652
transform 1 0 1528 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5559_6
timestamp 1731220652
transform 1 0 1576 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5558_6
timestamp 1731220652
transform 1 0 1448 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5557_6
timestamp 1731220652
transform 1 0 1344 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5556_6
timestamp 1731220652
transform 1 0 1440 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5555_6
timestamp 1731220652
transform 1 0 1344 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5554_6
timestamp 1731220652
transform 1 0 1216 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5553_6
timestamp 1731220652
transform 1 0 1344 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5552_6
timestamp 1731220652
transform 1 0 1400 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5551_6
timestamp 1731220652
transform 1 0 1496 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5550_6
timestamp 1731220652
transform 1 0 1472 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5549_6
timestamp 1731220652
transform 1 0 1400 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5548_6
timestamp 1731220652
transform 1 0 1344 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5547_6
timestamp 1731220652
transform 1 0 1344 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5546_6
timestamp 1731220652
transform 1 0 1400 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5545_6
timestamp 1731220652
transform 1 0 1344 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5544_6
timestamp 1731220652
transform 1 0 1416 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5543_6
timestamp 1731220652
transform 1 0 1520 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5542_6
timestamp 1731220652
transform 1 0 1416 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5541_6
timestamp 1731220652
transform 1 0 1344 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5540_6
timestamp 1731220652
transform 1 0 1344 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5539_6
timestamp 1731220652
transform 1 0 1416 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5538_6
timestamp 1731220652
transform 1 0 1496 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5537_6
timestamp 1731220652
transform 1 0 1408 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5536_6
timestamp 1731220652
transform 1 0 1344 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5535_6
timestamp 1731220652
transform 1 0 1344 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5534_6
timestamp 1731220652
transform 1 0 1640 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5533_6
timestamp 1731220652
transform 1 0 1528 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5532_6
timestamp 1731220652
transform 1 0 1424 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5531_6
timestamp 1731220652
transform 1 0 1352 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5530_6
timestamp 1731220652
transform 1 0 1448 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5529_6
timestamp 1731220652
transform 1 0 1752 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5528_6
timestamp 1731220652
transform 1 0 1648 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5527_6
timestamp 1731220652
transform 1 0 1544 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5526_6
timestamp 1731220652
transform 1 0 1456 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5525_6
timestamp 1731220652
transform 1 0 1552 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5524_6
timestamp 1731220652
transform 1 0 1872 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5523_6
timestamp 1731220652
transform 1 0 1760 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5522_6
timestamp 1731220652
transform 1 0 1656 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5521_6
timestamp 1731220652
transform 1 0 1664 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5520_6
timestamp 1731220652
transform 1 0 1584 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5519_6
timestamp 1731220652
transform 1 0 1512 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5518_6
timestamp 1731220652
transform 1 0 1760 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5517_6
timestamp 1731220652
transform 1 0 1856 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5516_6
timestamp 1731220652
transform 1 0 1960 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5515_6
timestamp 1731220652
transform 1 0 1912 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5514_6
timestamp 1731220652
transform 1 0 1808 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5513_6
timestamp 1731220652
transform 1 0 1704 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5512_6
timestamp 1731220652
transform 1 0 1608 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5511_6
timestamp 1731220652
transform 1 0 1520 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5510_6
timestamp 1731220652
transform 1 0 1816 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5509_6
timestamp 1731220652
transform 1 0 1712 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5508_6
timestamp 1731220652
transform 1 0 1616 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5507_6
timestamp 1731220652
transform 1 0 1520 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5506_6
timestamp 1731220652
transform 1 0 1432 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5505_6
timestamp 1731220652
transform 1 0 1712 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5504_6
timestamp 1731220652
transform 1 0 1608 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5503_6
timestamp 1731220652
transform 1 0 1512 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5502_6
timestamp 1731220652
transform 1 0 1416 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5501_6
timestamp 1731220652
transform 1 0 1344 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5500_6
timestamp 1731220652
transform 1 0 1656 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5499_6
timestamp 1731220652
transform 1 0 1568 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5498_6
timestamp 1731220652
transform 1 0 1480 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5497_6
timestamp 1731220652
transform 1 0 1400 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5496_6
timestamp 1731220652
transform 1 0 1344 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5495_6
timestamp 1731220652
transform 1 0 1216 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5494_6
timestamp 1731220652
transform 1 0 1160 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5493_6
timestamp 1731220652
transform 1 0 1216 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5492_6
timestamp 1731220652
transform 1 0 1128 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5491_6
timestamp 1731220652
transform 1 0 1016 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5490_6
timestamp 1731220652
transform 1 0 904 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5489_6
timestamp 1731220652
transform 1 0 1096 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5488_6
timestamp 1731220652
transform 1 0 1024 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5487_6
timestamp 1731220652
transform 1 0 960 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5486_6
timestamp 1731220652
transform 1 0 896 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5485_6
timestamp 1731220652
transform 1 0 824 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5484_6
timestamp 1731220652
transform 1 0 752 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5483_6
timestamp 1731220652
transform 1 0 1040 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5482_6
timestamp 1731220652
transform 1 0 952 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5481_6
timestamp 1731220652
transform 1 0 864 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5480_6
timestamp 1731220652
transform 1 0 776 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5479_6
timestamp 1731220652
transform 1 0 696 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5478_6
timestamp 1731220652
transform 1 0 688 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5477_6
timestamp 1731220652
transform 1 0 792 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5476_6
timestamp 1731220652
transform 1 0 1008 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5475_6
timestamp 1731220652
transform 1 0 896 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5474_6
timestamp 1731220652
transform 1 0 840 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5473_6
timestamp 1731220652
transform 1 0 1016 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5472_6
timestamp 1731220652
transform 1 0 1032 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5471_6
timestamp 1731220652
transform 1 0 1016 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5470_6
timestamp 1731220652
transform 1 0 1096 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5469_6
timestamp 1731220652
transform 1 0 1096 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5468_6
timestamp 1731220652
transform 1 0 1152 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5467_6
timestamp 1731220652
transform 1 0 1040 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5466_6
timestamp 1731220652
transform 1 0 1048 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5465_6
timestamp 1731220652
transform 1 0 1168 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5464_6
timestamp 1731220652
transform 1 0 1168 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5463_6
timestamp 1731220652
transform 1 0 1040 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5462_6
timestamp 1731220652
transform 1 0 944 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5461_6
timestamp 1731220652
transform 1 0 1056 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5460_6
timestamp 1731220652
transform 1 0 1168 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5459_6
timestamp 1731220652
transform 1 0 1144 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5458_6
timestamp 1731220652
transform 1 0 1040 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5457_6
timestamp 1731220652
transform 1 0 936 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5456_6
timestamp 1731220652
transform 1 0 832 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5455_6
timestamp 1731220652
transform 1 0 1080 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5454_6
timestamp 1731220652
transform 1 0 984 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5453_6
timestamp 1731220652
transform 1 0 888 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5452_6
timestamp 1731220652
transform 1 0 800 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5451_6
timestamp 1731220652
transform 1 0 704 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5450_6
timestamp 1731220652
transform 1 0 976 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5449_6
timestamp 1731220652
transform 1 0 872 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5448_6
timestamp 1731220652
transform 1 0 776 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5447_6
timestamp 1731220652
transform 1 0 680 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5446_6
timestamp 1731220652
transform 1 0 584 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5445_6
timestamp 1731220652
transform 1 0 872 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5444_6
timestamp 1731220652
transform 1 0 776 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5443_6
timestamp 1731220652
transform 1 0 680 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5442_6
timestamp 1731220652
transform 1 0 592 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5441_6
timestamp 1731220652
transform 1 0 504 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5440_6
timestamp 1731220652
transform 1 0 1072 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5439_6
timestamp 1731220652
transform 1 0 904 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5438_6
timestamp 1731220652
transform 1 0 752 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5437_6
timestamp 1731220652
transform 1 0 616 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5436_6
timestamp 1731220652
transform 1 0 624 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5435_6
timestamp 1731220652
transform 1 0 680 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5434_6
timestamp 1731220652
transform 1 0 736 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5433_6
timestamp 1731220652
transform 1 0 792 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5432_6
timestamp 1731220652
transform 1 0 848 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5431_6
timestamp 1731220652
transform 1 0 904 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5430_6
timestamp 1731220652
transform 1 0 848 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5429_6
timestamp 1731220652
transform 1 0 792 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5428_6
timestamp 1731220652
transform 1 0 736 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5427_6
timestamp 1731220652
transform 1 0 960 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5426_6
timestamp 1731220652
transform 1 0 904 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5425_6
timestamp 1731220652
transform 1 0 840 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5424_6
timestamp 1731220652
transform 1 0 760 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5423_6
timestamp 1731220652
transform 1 0 672 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5422_6
timestamp 1731220652
transform 1 0 920 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5421_6
timestamp 1731220652
transform 1 0 1096 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5420_6
timestamp 1731220652
transform 1 0 1008 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5419_6
timestamp 1731220652
transform 1 0 960 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5418_6
timestamp 1731220652
transform 1 0 856 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5417_6
timestamp 1731220652
transform 1 0 744 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5416_6
timestamp 1731220652
transform 1 0 1184 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5415_6
timestamp 1731220652
transform 1 0 1072 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5414_6
timestamp 1731220652
transform 1 0 752 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5413_6
timestamp 1731220652
transform 1 0 656 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5412_6
timestamp 1731220652
transform 1 0 928 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5411_6
timestamp 1731220652
transform 1 0 1008 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5410_6
timestamp 1731220652
transform 1 0 1080 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5409_6
timestamp 1731220652
transform 1 0 1216 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5408_6
timestamp 1731220652
transform 1 0 1160 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5407_6
timestamp 1731220652
transform 1 0 1152 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5406_6
timestamp 1731220652
transform 1 0 1344 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5405_6
timestamp 1731220652
transform 1 0 1216 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5404_6
timestamp 1731220652
transform 1 0 1216 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5403_6
timestamp 1731220652
transform 1 0 1160 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5402_6
timestamp 1731220652
transform 1 0 1080 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5401_6
timestamp 1731220652
transform 1 0 1000 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5400_6
timestamp 1731220652
transform 1 0 920 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5399_6
timestamp 1731220652
transform 1 0 832 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5398_6
timestamp 1731220652
transform 1 0 1072 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5397_6
timestamp 1731220652
transform 1 0 992 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5396_6
timestamp 1731220652
transform 1 0 904 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5395_6
timestamp 1731220652
transform 1 0 840 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5394_6
timestamp 1731220652
transform 1 0 808 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5393_6
timestamp 1731220652
transform 1 0 712 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5392_6
timestamp 1731220652
transform 1 0 736 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5391_6
timestamp 1731220652
transform 1 0 1048 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5390_6
timestamp 1731220652
transform 1 0 960 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5389_6
timestamp 1731220652
transform 1 0 872 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5388_6
timestamp 1731220652
transform 1 0 784 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5387_6
timestamp 1731220652
transform 1 0 704 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5386_6
timestamp 1731220652
transform 1 0 968 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5385_6
timestamp 1731220652
transform 1 0 888 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5384_6
timestamp 1731220652
transform 1 0 816 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5383_6
timestamp 1731220652
transform 1 0 744 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5382_6
timestamp 1731220652
transform 1 0 672 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5381_6
timestamp 1731220652
transform 1 0 600 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5380_6
timestamp 1731220652
transform 1 0 888 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5379_6
timestamp 1731220652
transform 1 0 816 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5378_6
timestamp 1731220652
transform 1 0 744 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5377_6
timestamp 1731220652
transform 1 0 680 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5376_6
timestamp 1731220652
transform 1 0 616 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5375_6
timestamp 1731220652
transform 1 0 584 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5374_6
timestamp 1731220652
transform 1 0 648 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5373_6
timestamp 1731220652
transform 1 0 712 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5372_6
timestamp 1731220652
transform 1 0 776 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5371_6
timestamp 1731220652
transform 1 0 912 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5370_6
timestamp 1731220652
transform 1 0 840 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5369_6
timestamp 1731220652
transform 1 0 824 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5368_6
timestamp 1731220652
transform 1 0 744 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5367_6
timestamp 1731220652
transform 1 0 664 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5366_6
timestamp 1731220652
transform 1 0 904 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5365_6
timestamp 1731220652
transform 1 0 1064 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5364_6
timestamp 1731220652
transform 1 0 984 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5363_6
timestamp 1731220652
transform 1 0 960 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5362_6
timestamp 1731220652
transform 1 0 872 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5361_6
timestamp 1731220652
transform 1 0 784 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5360_6
timestamp 1731220652
transform 1 0 1144 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5359_6
timestamp 1731220652
transform 1 0 1048 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5358_6
timestamp 1731220652
transform 1 0 1032 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5357_6
timestamp 1731220652
transform 1 0 928 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5356_6
timestamp 1731220652
transform 1 0 824 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5355_6
timestamp 1731220652
transform 1 0 1136 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5354_6
timestamp 1731220652
transform 1 0 1216 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5353_6
timestamp 1731220652
transform 1 0 1216 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5352_6
timestamp 1731220652
transform 1 0 1120 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5351_6
timestamp 1731220652
transform 1 0 1000 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5350_6
timestamp 1731220652
transform 1 0 944 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5349_6
timestamp 1731220652
transform 1 0 1016 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5348_6
timestamp 1731220652
transform 1 0 1088 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5347_6
timestamp 1731220652
transform 1 0 1024 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5346_6
timestamp 1731220652
transform 1 0 1128 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5345_6
timestamp 1731220652
transform 1 0 1192 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5344_6
timestamp 1731220652
transform 1 0 1088 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5343_6
timestamp 1731220652
transform 1 0 984 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5342_6
timestamp 1731220652
transform 1 0 952 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5341_6
timestamp 1731220652
transform 1 0 1040 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5340_6
timestamp 1731220652
transform 1 0 1128 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5339_6
timestamp 1731220652
transform 1 0 1176 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5338_6
timestamp 1731220652
transform 1 0 1112 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5337_6
timestamp 1731220652
transform 1 0 1048 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5336_6
timestamp 1731220652
transform 1 0 984 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5335_6
timestamp 1731220652
transform 1 0 920 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5334_6
timestamp 1731220652
transform 1 0 856 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5333_6
timestamp 1731220652
transform 1 0 792 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5332_6
timestamp 1731220652
transform 1 0 728 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5331_6
timestamp 1731220652
transform 1 0 664 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5330_6
timestamp 1731220652
transform 1 0 688 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5329_6
timestamp 1731220652
transform 1 0 776 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5328_6
timestamp 1731220652
transform 1 0 864 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5327_6
timestamp 1731220652
transform 1 0 784 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5326_6
timestamp 1731220652
transform 1 0 688 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5325_6
timestamp 1731220652
transform 1 0 880 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5324_6
timestamp 1731220652
transform 1 0 920 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5323_6
timestamp 1731220652
transform 1 0 816 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5322_6
timestamp 1731220652
transform 1 0 720 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5321_6
timestamp 1731220652
transform 1 0 624 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5320_6
timestamp 1731220652
transform 1 0 568 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5319_6
timestamp 1731220652
transform 1 0 648 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5318_6
timestamp 1731220652
transform 1 0 728 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5317_6
timestamp 1731220652
transform 1 0 800 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5316_6
timestamp 1731220652
transform 1 0 872 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5315_6
timestamp 1731220652
transform 1 0 888 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5314_6
timestamp 1731220652
transform 1 0 776 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5313_6
timestamp 1731220652
transform 1 0 664 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5312_6
timestamp 1731220652
transform 1 0 560 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5311_6
timestamp 1731220652
transform 1 0 592 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5310_6
timestamp 1731220652
transform 1 0 712 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5309_6
timestamp 1731220652
transform 1 0 688 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5308_6
timestamp 1731220652
transform 1 0 584 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5307_6
timestamp 1731220652
transform 1 0 480 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5306_6
timestamp 1731220652
transform 1 0 576 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5305_6
timestamp 1731220652
transform 1 0 480 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5304_6
timestamp 1731220652
transform 1 0 448 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5303_6
timestamp 1731220652
transform 1 0 520 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5302_6
timestamp 1731220652
transform 1 0 480 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5301_6
timestamp 1731220652
transform 1 0 400 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5300_6
timestamp 1731220652
transform 1 0 552 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5299_6
timestamp 1731220652
transform 1 0 520 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5298_6
timestamp 1731220652
transform 1 0 432 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5297_6
timestamp 1731220652
transform 1 0 320 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5296_6
timestamp 1731220652
transform 1 0 240 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5295_6
timestamp 1731220652
transform 1 0 288 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5294_6
timestamp 1731220652
transform 1 0 368 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5293_6
timestamp 1731220652
transform 1 0 384 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5292_6
timestamp 1731220652
transform 1 0 368 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5291_6
timestamp 1731220652
transform 1 0 264 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5290_6
timestamp 1731220652
transform 1 0 464 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5289_6
timestamp 1731220652
transform 1 0 344 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5288_6
timestamp 1731220652
transform 1 0 296 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5287_6
timestamp 1731220652
transform 1 0 240 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5286_6
timestamp 1731220652
transform 1 0 376 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5285_6
timestamp 1731220652
transform 1 0 464 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5284_6
timestamp 1731220652
transform 1 0 488 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5283_6
timestamp 1731220652
transform 1 0 408 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5282_6
timestamp 1731220652
transform 1 0 336 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5281_6
timestamp 1731220652
transform 1 0 448 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5280_6
timestamp 1731220652
transform 1 0 368 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5279_6
timestamp 1731220652
transform 1 0 536 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5278_6
timestamp 1731220652
transform 1 0 496 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5277_6
timestamp 1731220652
transform 1 0 400 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5276_6
timestamp 1731220652
transform 1 0 592 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5275_6
timestamp 1731220652
transform 1 0 600 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5274_6
timestamp 1731220652
transform 1 0 504 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5273_6
timestamp 1731220652
transform 1 0 408 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5272_6
timestamp 1731220652
transform 1 0 600 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5271_6
timestamp 1731220652
transform 1 0 528 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5270_6
timestamp 1731220652
transform 1 0 464 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5269_6
timestamp 1731220652
transform 1 0 408 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5268_6
timestamp 1731220652
transform 1 0 352 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5267_6
timestamp 1731220652
transform 1 0 296 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5266_6
timestamp 1731220652
transform 1 0 240 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5265_6
timestamp 1731220652
transform 1 0 184 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5264_6
timestamp 1731220652
transform 1 0 128 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5263_6
timestamp 1731220652
transform 1 0 152 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5262_6
timestamp 1731220652
transform 1 0 320 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5261_6
timestamp 1731220652
transform 1 0 232 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5260_6
timestamp 1731220652
transform 1 0 208 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5259_6
timestamp 1731220652
transform 1 0 128 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5258_6
timestamp 1731220652
transform 1 0 304 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5257_6
timestamp 1731220652
transform 1 0 280 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5256_6
timestamp 1731220652
transform 1 0 192 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5255_6
timestamp 1731220652
transform 1 0 128 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5254_6
timestamp 1731220652
transform 1 0 128 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5253_6
timestamp 1731220652
transform 1 0 256 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5252_6
timestamp 1731220652
transform 1 0 184 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5251_6
timestamp 1731220652
transform 1 0 184 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5250_6
timestamp 1731220652
transform 1 0 128 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5249_6
timestamp 1731220652
transform 1 0 128 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5248_6
timestamp 1731220652
transform 1 0 224 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5247_6
timestamp 1731220652
transform 1 0 168 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5246_6
timestamp 1731220652
transform 1 0 184 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5245_6
timestamp 1731220652
transform 1 0 280 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5244_6
timestamp 1731220652
transform 1 0 208 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5243_6
timestamp 1731220652
transform 1 0 152 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5242_6
timestamp 1731220652
transform 1 0 144 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5241_6
timestamp 1731220652
transform 1 0 240 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5240_6
timestamp 1731220652
transform 1 0 336 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5239_6
timestamp 1731220652
transform 1 0 280 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5238_6
timestamp 1731220652
transform 1 0 216 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5237_6
timestamp 1731220652
transform 1 0 360 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5236_6
timestamp 1731220652
transform 1 0 440 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5235_6
timestamp 1731220652
transform 1 0 528 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5234_6
timestamp 1731220652
transform 1 0 616 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5233_6
timestamp 1731220652
transform 1 0 640 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5232_6
timestamp 1731220652
transform 1 0 536 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5231_6
timestamp 1731220652
transform 1 0 432 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5230_6
timestamp 1731220652
transform 1 0 336 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5229_6
timestamp 1731220652
transform 1 0 240 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5228_6
timestamp 1731220652
transform 1 0 600 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5227_6
timestamp 1731220652
transform 1 0 488 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5226_6
timestamp 1731220652
transform 1 0 376 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5225_6
timestamp 1731220652
transform 1 0 272 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5224_6
timestamp 1731220652
transform 1 0 184 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5223_6
timestamp 1731220652
transform 1 0 128 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5222_6
timestamp 1731220652
transform 1 0 128 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5221_6
timestamp 1731220652
transform 1 0 208 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5220_6
timestamp 1731220652
transform 1 0 544 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5219_6
timestamp 1731220652
transform 1 0 432 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5218_6
timestamp 1731220652
transform 1 0 320 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5217_6
timestamp 1731220652
transform 1 0 280 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5216_6
timestamp 1731220652
transform 1 0 184 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5215_6
timestamp 1731220652
transform 1 0 128 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5214_6
timestamp 1731220652
transform 1 0 632 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5213_6
timestamp 1731220652
transform 1 0 512 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5212_6
timestamp 1731220652
transform 1 0 392 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5211_6
timestamp 1731220652
transform 1 0 392 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5210_6
timestamp 1731220652
transform 1 0 304 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5209_6
timestamp 1731220652
transform 1 0 216 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5208_6
timestamp 1731220652
transform 1 0 488 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5207_6
timestamp 1731220652
transform 1 0 584 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5206_6
timestamp 1731220652
transform 1 0 512 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5205_6
timestamp 1731220652
transform 1 0 456 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5204_6
timestamp 1731220652
transform 1 0 400 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5203_6
timestamp 1731220652
transform 1 0 568 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5202_6
timestamp 1731220652
transform 1 0 680 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5201_6
timestamp 1731220652
transform 1 0 624 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5200_6
timestamp 1731220652
transform 1 0 568 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5199_6
timestamp 1731220652
transform 1 0 512 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5198_6
timestamp 1731220652
transform 1 0 456 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5197_6
timestamp 1731220652
transform 1 0 400 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5196_6
timestamp 1731220652
transform 1 0 344 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5195_6
timestamp 1731220652
transform 1 0 504 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5194_6
timestamp 1731220652
transform 1 0 416 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5193_6
timestamp 1731220652
transform 1 0 344 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5192_6
timestamp 1731220652
transform 1 0 280 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5191_6
timestamp 1731220652
transform 1 0 224 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5190_6
timestamp 1731220652
transform 1 0 168 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5189_6
timestamp 1731220652
transform 1 0 408 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5188_6
timestamp 1731220652
transform 1 0 312 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5187_6
timestamp 1731220652
transform 1 0 208 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5186_6
timestamp 1731220652
transform 1 0 128 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5185_6
timestamp 1731220652
transform 1 0 128 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5184_6
timestamp 1731220652
transform 1 0 192 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5183_6
timestamp 1731220652
transform 1 0 288 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5182_6
timestamp 1731220652
transform 1 0 384 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5181_6
timestamp 1731220652
transform 1 0 488 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5180_6
timestamp 1731220652
transform 1 0 408 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5179_6
timestamp 1731220652
transform 1 0 312 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5178_6
timestamp 1731220652
transform 1 0 224 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5177_6
timestamp 1731220652
transform 1 0 504 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5176_6
timestamp 1731220652
transform 1 0 608 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5175_6
timestamp 1731220652
transform 1 0 536 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5174_6
timestamp 1731220652
transform 1 0 440 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5173_6
timestamp 1731220652
transform 1 0 352 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5172_6
timestamp 1731220652
transform 1 0 728 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5171_6
timestamp 1731220652
transform 1 0 632 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5170_6
timestamp 1731220652
transform 1 0 632 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5169_6
timestamp 1731220652
transform 1 0 544 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5168_6
timestamp 1731220652
transform 1 0 464 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5167_6
timestamp 1731220652
transform 1 0 832 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5166_6
timestamp 1731220652
transform 1 0 728 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5165_6
timestamp 1731220652
transform 1 0 680 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5164_6
timestamp 1731220652
transform 1 0 576 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5163_6
timestamp 1731220652
transform 1 0 912 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5162_6
timestamp 1731220652
transform 1 0 792 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5161_6
timestamp 1731220652
transform 1 0 736 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5160_6
timestamp 1731220652
transform 1 0 640 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5159_6
timestamp 1731220652
transform 1 0 832 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5158_6
timestamp 1731220652
transform 1 0 936 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5157_6
timestamp 1731220652
transform 1 0 928 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5156_6
timestamp 1731220652
transform 1 0 824 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5155_6
timestamp 1731220652
transform 1 0 720 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5154_6
timestamp 1731220652
transform 1 0 672 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5153_6
timestamp 1731220652
transform 1 0 776 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5152_6
timestamp 1731220652
transform 1 0 880 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5151_6
timestamp 1731220652
transform 1 0 984 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5150_6
timestamp 1731220652
transform 1 0 936 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5149_6
timestamp 1731220652
transform 1 0 856 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5148_6
timestamp 1731220652
transform 1 0 776 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5147_6
timestamp 1731220652
transform 1 0 696 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5146_6
timestamp 1731220652
transform 1 0 952 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5145_6
timestamp 1731220652
transform 1 0 880 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5144_6
timestamp 1731220652
transform 1 0 808 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5143_6
timestamp 1731220652
transform 1 0 736 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5142_6
timestamp 1731220652
transform 1 0 672 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5141_6
timestamp 1731220652
transform 1 0 608 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5140_6
timestamp 1731220652
transform 1 0 544 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5139_6
timestamp 1731220652
transform 1 0 472 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5138_6
timestamp 1731220652
transform 1 0 400 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5137_6
timestamp 1731220652
transform 1 0 416 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5136_6
timestamp 1731220652
transform 1 0 608 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5135_6
timestamp 1731220652
transform 1 0 512 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5134_6
timestamp 1731220652
transform 1 0 456 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5133_6
timestamp 1731220652
transform 1 0 568 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5132_6
timestamp 1731220652
transform 1 0 616 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5131_6
timestamp 1731220652
transform 1 0 512 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5130_6
timestamp 1731220652
transform 1 0 416 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5129_6
timestamp 1731220652
transform 1 0 400 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5128_6
timestamp 1731220652
transform 1 0 472 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5127_6
timestamp 1731220652
transform 1 0 552 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5126_6
timestamp 1731220652
transform 1 0 480 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5125_6
timestamp 1731220652
transform 1 0 400 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5124_6
timestamp 1731220652
transform 1 0 328 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5123_6
timestamp 1731220652
transform 1 0 264 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5122_6
timestamp 1731220652
transform 1 0 264 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5121_6
timestamp 1731220652
transform 1 0 208 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5120_6
timestamp 1731220652
transform 1 0 328 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5119_6
timestamp 1731220652
transform 1 0 328 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5118_6
timestamp 1731220652
transform 1 0 248 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5117_6
timestamp 1731220652
transform 1 0 168 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5116_6
timestamp 1731220652
transform 1 0 128 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5115_6
timestamp 1731220652
transform 1 0 232 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5114_6
timestamp 1731220652
transform 1 0 344 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5113_6
timestamp 1731220652
transform 1 0 312 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5112_6
timestamp 1731220652
transform 1 0 208 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5111_6
timestamp 1731220652
transform 1 0 128 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5110_6
timestamp 1731220652
transform 1 0 128 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5109_6
timestamp 1731220652
transform 1 0 328 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5108_6
timestamp 1731220652
transform 1 0 256 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5107_6
timestamp 1731220652
transform 1 0 184 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5106_6
timestamp 1731220652
transform 1 0 128 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5105_6
timestamp 1731220652
transform 1 0 216 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5104_6
timestamp 1731220652
transform 1 0 664 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5103_6
timestamp 1731220652
transform 1 0 504 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5102_6
timestamp 1731220652
transform 1 0 352 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5101_6
timestamp 1731220652
transform 1 0 280 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5100_6
timestamp 1731220652
transform 1 0 200 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_599_6
timestamp 1731220652
transform 1 0 128 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_598_6
timestamp 1731220652
transform 1 0 584 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_597_6
timestamp 1731220652
transform 1 0 480 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_596_6
timestamp 1731220652
transform 1 0 376 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_595_6
timestamp 1731220652
transform 1 0 352 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_594_6
timestamp 1731220652
transform 1 0 272 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_593_6
timestamp 1731220652
transform 1 0 616 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_592_6
timestamp 1731220652
transform 1 0 528 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_591_6
timestamp 1731220652
transform 1 0 440 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_590_6
timestamp 1731220652
transform 1 0 368 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_589_6
timestamp 1731220652
transform 1 0 440 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_588_6
timestamp 1731220652
transform 1 0 512 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_587_6
timestamp 1731220652
transform 1 0 592 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_586_6
timestamp 1731220652
transform 1 0 672 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_585_6
timestamp 1731220652
transform 1 0 792 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_584_6
timestamp 1731220652
transform 1 0 688 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_583_6
timestamp 1731220652
transform 1 0 584 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_582_6
timestamp 1731220652
transform 1 0 488 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_581_6
timestamp 1731220652
transform 1 0 392 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_580_6
timestamp 1731220652
transform 1 0 552 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_579_6
timestamp 1731220652
transform 1 0 496 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_578_6
timestamp 1731220652
transform 1 0 440 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_577_6
timestamp 1731220652
transform 1 0 384 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_576_6
timestamp 1731220652
transform 1 0 328 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_575_6
timestamp 1731220652
transform 1 0 480 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_574_6
timestamp 1731220652
transform 1 0 424 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_573_6
timestamp 1731220652
transform 1 0 360 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_572_6
timestamp 1731220652
transform 1 0 296 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_571_6
timestamp 1731220652
transform 1 0 240 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_570_6
timestamp 1731220652
transform 1 0 464 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_569_6
timestamp 1731220652
transform 1 0 368 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_568_6
timestamp 1731220652
transform 1 0 280 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_567_6
timestamp 1731220652
transform 1 0 200 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_566_6
timestamp 1731220652
transform 1 0 480 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_565_6
timestamp 1731220652
transform 1 0 368 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_564_6
timestamp 1731220652
transform 1 0 256 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_563_6
timestamp 1731220652
transform 1 0 152 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_562_6
timestamp 1731220652
transform 1 0 408 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_561_6
timestamp 1731220652
transform 1 0 312 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_560_6
timestamp 1731220652
transform 1 0 224 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_559_6
timestamp 1731220652
transform 1 0 144 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_558_6
timestamp 1731220652
transform 1 0 160 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_557_6
timestamp 1731220652
transform 1 0 392 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_556_6
timestamp 1731220652
transform 1 0 304 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_555_6
timestamp 1731220652
transform 1 0 224 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_554_6
timestamp 1731220652
transform 1 0 216 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_553_6
timestamp 1731220652
transform 1 0 160 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_552_6
timestamp 1731220652
transform 1 0 272 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_551_6
timestamp 1731220652
transform 1 0 336 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_550_6
timestamp 1731220652
transform 1 0 400 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_549_6
timestamp 1731220652
transform 1 0 472 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_548_6
timestamp 1731220652
transform 1 0 552 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_547_6
timestamp 1731220652
transform 1 0 632 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_546_6
timestamp 1731220652
transform 1 0 576 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_545_6
timestamp 1731220652
transform 1 0 480 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_544_6
timestamp 1731220652
transform 1 0 672 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_543_6
timestamp 1731220652
transform 1 0 720 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_542_6
timestamp 1731220652
transform 1 0 616 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_541_6
timestamp 1731220652
transform 1 0 512 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_540_6
timestamp 1731220652
transform 1 0 600 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_539_6
timestamp 1731220652
transform 1 0 720 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_538_6
timestamp 1731220652
transform 1 0 728 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_537_6
timestamp 1731220652
transform 1 0 640 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_536_6
timestamp 1731220652
transform 1 0 552 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_535_6
timestamp 1731220652
transform 1 0 536 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_534_6
timestamp 1731220652
transform 1 0 592 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_533_6
timestamp 1731220652
transform 1 0 648 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_532_6
timestamp 1731220652
transform 1 0 704 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_531_6
timestamp 1731220652
transform 1 0 768 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_530_6
timestamp 1731220652
transform 1 0 832 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_529_6
timestamp 1731220652
transform 1 0 896 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_528_6
timestamp 1731220652
transform 1 0 1088 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_527_6
timestamp 1731220652
transform 1 0 1024 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_526_6
timestamp 1731220652
transform 1 0 960 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_525_6
timestamp 1731220652
transform 1 0 896 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_524_6
timestamp 1731220652
transform 1 0 808 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_523_6
timestamp 1731220652
transform 1 0 1072 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_522_6
timestamp 1731220652
transform 1 0 984 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_521_6
timestamp 1731220652
transform 1 0 976 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_520_6
timestamp 1731220652
transform 1 0 848 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_519_6
timestamp 1731220652
transform 1 0 1104 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_518_6
timestamp 1731220652
transform 1 0 1144 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_517_6
timestamp 1731220652
transform 1 0 1032 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_516_6
timestamp 1731220652
transform 1 0 928 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_515_6
timestamp 1731220652
transform 1 0 824 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_514_6
timestamp 1731220652
transform 1 0 1136 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_513_6
timestamp 1731220652
transform 1 0 1040 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_512_6
timestamp 1731220652
transform 1 0 944 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_511_6
timestamp 1731220652
transform 1 0 856 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_510_6
timestamp 1731220652
transform 1 0 768 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_59_6
timestamp 1731220652
transform 1 0 1032 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_58_6
timestamp 1731220652
transform 1 0 952 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_57_6
timestamp 1731220652
transform 1 0 872 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_56_6
timestamp 1731220652
transform 1 0 792 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_55_6
timestamp 1731220652
transform 1 0 712 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_54_6
timestamp 1731220652
transform 1 0 920 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_53_6
timestamp 1731220652
transform 1 0 864 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_52_6
timestamp 1731220652
transform 1 0 808 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_51_6
timestamp 1731220652
transform 1 0 752 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_50_6
timestamp 1731220652
transform 1 0 696 0 1 2528
box 4 4 48 48
<< end >>
