magic
tech sky130l
timestamp 1730953945
<< m1 >>
rect 728 1055 732 1071
rect 472 1019 476 1035
rect 512 943 516 1035
rect 400 895 404 939
rect 512 887 516 911
rect 1024 895 1028 911
rect 712 831 716 875
rect 1040 791 1044 875
rect 488 683 492 727
rect 648 683 652 727
rect 640 587 644 631
rect 712 431 716 475
rect 808 431 812 475
rect 440 283 444 327
rect 552 283 556 327
rect 672 283 676 327
rect 800 283 804 327
rect 536 243 540 271
rect 216 99 220 143
rect 304 99 308 143
<< m2c >>
rect 111 1249 115 1253
rect 1183 1249 1187 1253
rect 111 1231 115 1235
rect 1183 1231 1187 1235
rect 111 1181 115 1185
rect 1183 1181 1187 1185
rect 111 1163 115 1167
rect 1183 1163 1187 1167
rect 111 1089 115 1093
rect 1183 1089 1187 1093
rect 111 1071 115 1075
rect 496 1071 500 1075
rect 728 1071 732 1075
rect 792 1071 796 1075
rect 1088 1071 1092 1075
rect 1183 1071 1187 1075
rect 728 1051 732 1055
rect 472 1035 476 1039
rect 111 1013 115 1017
rect 384 1015 388 1019
rect 472 1015 476 1019
rect 512 1035 516 1039
rect 111 995 115 999
rect 536 1015 540 1019
rect 1183 1013 1187 1017
rect 1183 995 1187 999
rect 400 939 404 943
rect 512 939 516 943
rect 111 929 115 933
rect 111 911 115 915
rect 1183 929 1187 933
rect 400 891 404 895
rect 512 911 516 915
rect 552 911 556 915
rect 680 911 684 915
rect 1024 911 1028 915
rect 1080 911 1084 915
rect 1183 911 1187 915
rect 1024 891 1028 895
rect 512 883 516 887
rect 712 875 716 879
rect 111 853 115 857
rect 111 835 115 839
rect 1040 875 1044 879
rect 768 855 772 859
rect 712 827 716 831
rect 1183 853 1187 857
rect 1183 835 1187 839
rect 1040 787 1044 791
rect 111 777 115 781
rect 1183 777 1187 781
rect 111 759 115 763
rect 512 759 516 763
rect 656 759 660 763
rect 1088 759 1092 763
rect 1183 759 1187 763
rect 488 727 492 731
rect 111 705 115 709
rect 111 687 115 691
rect 488 679 492 683
rect 648 727 652 731
rect 720 707 724 711
rect 1183 705 1187 709
rect 1183 687 1187 691
rect 648 679 652 683
rect 640 631 644 635
rect 111 621 115 625
rect 111 603 115 607
rect 240 603 244 607
rect 384 603 388 607
rect 1183 621 1187 625
rect 712 603 716 607
rect 1183 603 1187 607
rect 640 583 644 587
rect 111 549 115 553
rect 624 551 628 555
rect 768 551 772 555
rect 1183 549 1187 553
rect 111 531 115 535
rect 1183 531 1187 535
rect 712 475 716 479
rect 111 465 115 469
rect 111 447 115 451
rect 712 427 716 431
rect 808 475 812 479
rect 1183 465 1187 469
rect 1088 447 1092 451
rect 1183 447 1187 451
rect 808 427 812 431
rect 111 393 115 397
rect 1183 393 1187 397
rect 648 383 652 387
rect 111 375 115 379
rect 1183 375 1187 379
rect 440 327 444 331
rect 111 317 115 321
rect 111 299 115 303
rect 440 279 444 283
rect 552 327 556 331
rect 552 279 556 283
rect 672 327 676 331
rect 672 279 676 283
rect 800 327 804 331
rect 1183 317 1187 321
rect 1183 299 1187 303
rect 800 279 804 283
rect 536 271 540 275
rect 111 237 115 241
rect 536 239 540 243
rect 544 239 548 243
rect 1183 237 1187 241
rect 111 219 115 223
rect 1183 219 1187 223
rect 216 143 220 147
rect 111 133 115 137
rect 111 115 115 119
rect 216 95 220 99
rect 304 143 308 147
rect 1183 133 1187 137
rect 1183 115 1187 119
rect 304 95 308 99
<< m2 >>
rect 574 1271 580 1272
rect 574 1267 575 1271
rect 579 1267 580 1271
rect 574 1266 580 1267
rect 682 1263 688 1264
rect 682 1262 683 1263
rect 625 1260 683 1262
rect 682 1259 683 1260
rect 687 1259 688 1263
rect 682 1258 688 1259
rect 110 1253 116 1254
rect 110 1249 111 1253
rect 115 1249 116 1253
rect 110 1248 116 1249
rect 1182 1253 1188 1254
rect 1182 1249 1183 1253
rect 1187 1249 1188 1253
rect 1182 1248 1188 1249
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1182 1235 1188 1236
rect 1182 1231 1183 1235
rect 1187 1231 1188 1235
rect 110 1230 116 1231
rect 578 1230 584 1231
rect 1182 1230 1188 1231
rect 578 1226 579 1230
rect 583 1226 584 1230
rect 578 1225 584 1226
rect 594 1215 600 1216
rect 594 1211 595 1215
rect 599 1211 600 1215
rect 594 1210 600 1211
rect 234 1207 240 1208
rect 234 1203 235 1207
rect 239 1203 240 1207
rect 234 1202 240 1203
rect 286 1207 292 1208
rect 286 1203 287 1207
rect 291 1206 292 1207
rect 374 1207 380 1208
rect 291 1204 325 1206
rect 291 1203 292 1204
rect 286 1202 292 1203
rect 374 1203 375 1207
rect 379 1206 380 1207
rect 462 1207 468 1208
rect 379 1204 413 1206
rect 379 1203 380 1204
rect 374 1202 380 1203
rect 462 1203 463 1207
rect 467 1206 468 1207
rect 550 1207 556 1208
rect 467 1204 501 1206
rect 467 1203 468 1204
rect 462 1202 468 1203
rect 550 1203 551 1207
rect 555 1206 556 1207
rect 682 1207 688 1208
rect 555 1204 589 1206
rect 555 1203 556 1204
rect 550 1202 556 1203
rect 682 1203 683 1207
rect 687 1203 688 1207
rect 682 1202 688 1203
rect 734 1207 740 1208
rect 734 1203 735 1207
rect 739 1206 740 1207
rect 838 1207 844 1208
rect 739 1204 789 1206
rect 739 1203 740 1204
rect 734 1202 740 1203
rect 838 1203 839 1207
rect 843 1206 844 1207
rect 1026 1207 1032 1208
rect 1026 1206 1027 1207
rect 843 1204 901 1206
rect 1021 1204 1027 1206
rect 843 1203 844 1204
rect 838 1202 844 1203
rect 1026 1203 1027 1204
rect 1031 1203 1032 1207
rect 1026 1202 1032 1203
rect 1070 1207 1076 1208
rect 1070 1203 1071 1207
rect 1075 1206 1076 1207
rect 1075 1204 1117 1206
rect 1075 1203 1076 1204
rect 1070 1202 1076 1203
rect 218 1190 224 1191
rect 218 1186 219 1190
rect 223 1186 224 1190
rect 110 1185 116 1186
rect 218 1185 224 1186
rect 306 1190 312 1191
rect 306 1186 307 1190
rect 311 1186 312 1190
rect 306 1185 312 1186
rect 394 1190 400 1191
rect 394 1186 395 1190
rect 399 1186 400 1190
rect 394 1185 400 1186
rect 482 1190 488 1191
rect 482 1186 483 1190
rect 487 1186 488 1190
rect 482 1185 488 1186
rect 570 1190 576 1191
rect 570 1186 571 1190
rect 575 1186 576 1190
rect 570 1185 576 1186
rect 666 1190 672 1191
rect 666 1186 667 1190
rect 671 1186 672 1190
rect 666 1185 672 1186
rect 770 1190 776 1191
rect 770 1186 771 1190
rect 775 1186 776 1190
rect 770 1185 776 1186
rect 882 1190 888 1191
rect 882 1186 883 1190
rect 887 1186 888 1190
rect 882 1185 888 1186
rect 1002 1190 1008 1191
rect 1002 1186 1003 1190
rect 1007 1186 1008 1190
rect 1002 1185 1008 1186
rect 1098 1190 1104 1191
rect 1098 1186 1099 1190
rect 1103 1186 1104 1190
rect 1098 1185 1104 1186
rect 1182 1185 1188 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 1182 1181 1183 1185
rect 1187 1181 1188 1185
rect 1182 1180 1188 1181
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 110 1162 116 1163
rect 1182 1167 1188 1168
rect 1182 1163 1183 1167
rect 1187 1163 1188 1167
rect 1182 1162 1188 1163
rect 286 1159 292 1160
rect 286 1158 287 1159
rect 265 1156 287 1158
rect 286 1155 287 1156
rect 291 1155 292 1159
rect 374 1159 380 1160
rect 374 1158 375 1159
rect 353 1156 375 1158
rect 286 1154 292 1155
rect 374 1155 375 1156
rect 379 1155 380 1159
rect 462 1159 468 1160
rect 462 1158 463 1159
rect 441 1156 463 1158
rect 374 1154 380 1155
rect 462 1155 463 1156
rect 467 1155 468 1159
rect 550 1159 556 1160
rect 550 1158 551 1159
rect 529 1156 551 1158
rect 462 1154 468 1155
rect 550 1155 551 1156
rect 555 1155 556 1159
rect 550 1154 556 1155
rect 590 1159 596 1160
rect 590 1155 591 1159
rect 595 1155 596 1159
rect 734 1159 740 1160
rect 734 1158 735 1159
rect 713 1156 735 1158
rect 590 1154 596 1155
rect 734 1155 735 1156
rect 739 1155 740 1159
rect 838 1159 844 1160
rect 838 1158 839 1159
rect 817 1156 839 1158
rect 734 1154 740 1155
rect 838 1155 839 1156
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 870 1159 876 1160
rect 870 1155 871 1159
rect 875 1155 876 1159
rect 1070 1159 1076 1160
rect 1070 1158 1071 1159
rect 1049 1156 1071 1158
rect 870 1154 876 1155
rect 1070 1155 1071 1156
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 214 1149 220 1150
rect 214 1145 215 1149
rect 219 1145 220 1149
rect 214 1144 220 1145
rect 302 1149 308 1150
rect 302 1145 303 1149
rect 307 1145 308 1149
rect 302 1144 308 1145
rect 390 1149 396 1150
rect 390 1145 391 1149
rect 395 1145 396 1149
rect 390 1144 396 1145
rect 478 1149 484 1150
rect 478 1145 479 1149
rect 483 1145 484 1149
rect 478 1144 484 1145
rect 566 1149 572 1150
rect 566 1145 567 1149
rect 571 1145 572 1149
rect 566 1144 572 1145
rect 662 1149 668 1150
rect 662 1145 663 1149
rect 667 1145 668 1149
rect 662 1144 668 1145
rect 766 1149 772 1150
rect 766 1145 767 1149
rect 771 1145 772 1149
rect 766 1144 772 1145
rect 878 1149 884 1150
rect 878 1145 879 1149
rect 883 1145 884 1149
rect 878 1144 884 1145
rect 998 1149 1004 1150
rect 998 1145 999 1149
rect 1003 1145 1004 1149
rect 998 1144 1004 1145
rect 1094 1149 1100 1150
rect 1094 1145 1095 1149
rect 1099 1145 1100 1149
rect 1094 1144 1100 1145
rect 214 1111 220 1112
rect 214 1107 215 1111
rect 219 1107 220 1111
rect 214 1106 220 1107
rect 358 1111 364 1112
rect 358 1107 359 1111
rect 363 1107 364 1111
rect 358 1106 364 1107
rect 502 1111 508 1112
rect 502 1107 503 1111
rect 507 1107 508 1111
rect 502 1106 508 1107
rect 646 1111 652 1112
rect 646 1107 647 1111
rect 651 1107 652 1111
rect 646 1106 652 1107
rect 798 1111 804 1112
rect 798 1107 799 1111
rect 803 1107 804 1111
rect 798 1106 804 1107
rect 950 1111 956 1112
rect 950 1107 951 1111
rect 955 1107 956 1111
rect 950 1106 956 1107
rect 1094 1111 1100 1112
rect 1094 1107 1095 1111
rect 1099 1107 1100 1111
rect 1094 1106 1100 1107
rect 438 1103 444 1104
rect 438 1102 439 1103
rect 409 1100 439 1102
rect 234 1099 240 1100
rect 234 1095 235 1099
rect 239 1095 240 1099
rect 438 1099 439 1100
rect 443 1099 444 1103
rect 722 1103 728 1104
rect 722 1102 723 1103
rect 697 1100 723 1102
rect 438 1098 444 1099
rect 722 1099 723 1100
rect 727 1099 728 1103
rect 1026 1103 1032 1104
rect 1026 1102 1027 1103
rect 1001 1100 1027 1102
rect 722 1098 728 1099
rect 1026 1099 1027 1100
rect 1031 1099 1032 1103
rect 1026 1098 1032 1099
rect 234 1094 240 1095
rect 110 1093 116 1094
rect 110 1089 111 1093
rect 115 1089 116 1093
rect 110 1088 116 1089
rect 1182 1093 1188 1094
rect 1182 1089 1183 1093
rect 1187 1089 1188 1093
rect 1182 1088 1188 1089
rect 110 1075 116 1076
rect 110 1071 111 1075
rect 115 1071 116 1075
rect 430 1075 436 1076
rect 430 1071 431 1075
rect 435 1074 436 1075
rect 495 1075 501 1076
rect 495 1074 496 1075
rect 435 1072 496 1074
rect 435 1071 436 1072
rect 110 1070 116 1071
rect 218 1070 224 1071
rect 218 1066 219 1070
rect 223 1066 224 1070
rect 218 1065 224 1066
rect 362 1070 368 1071
rect 430 1070 436 1071
rect 495 1071 496 1072
rect 500 1071 501 1075
rect 727 1075 733 1076
rect 727 1071 728 1075
rect 732 1074 733 1075
rect 791 1075 797 1076
rect 791 1074 792 1075
rect 732 1072 792 1074
rect 732 1071 733 1072
rect 495 1070 501 1071
rect 506 1070 512 1071
rect 362 1066 363 1070
rect 367 1066 368 1070
rect 362 1065 368 1066
rect 506 1066 507 1070
rect 511 1066 512 1070
rect 506 1065 512 1066
rect 650 1070 656 1071
rect 727 1070 733 1071
rect 791 1071 792 1072
rect 796 1071 797 1075
rect 1026 1075 1032 1076
rect 1026 1071 1027 1075
rect 1031 1074 1032 1075
rect 1087 1075 1093 1076
rect 1087 1074 1088 1075
rect 1031 1072 1088 1074
rect 1031 1071 1032 1072
rect 791 1070 797 1071
rect 802 1070 808 1071
rect 650 1066 651 1070
rect 655 1066 656 1070
rect 650 1065 656 1066
rect 802 1066 803 1070
rect 807 1066 808 1070
rect 802 1065 808 1066
rect 954 1070 960 1071
rect 1026 1070 1032 1071
rect 1087 1071 1088 1072
rect 1092 1071 1093 1075
rect 1182 1075 1188 1076
rect 1182 1071 1183 1075
rect 1187 1071 1188 1075
rect 1087 1070 1093 1071
rect 1098 1070 1104 1071
rect 1182 1070 1188 1071
rect 954 1066 955 1070
rect 959 1066 960 1070
rect 954 1065 960 1066
rect 1098 1066 1099 1070
rect 1103 1066 1104 1070
rect 1098 1065 1104 1066
rect 310 1055 316 1056
rect 310 1051 311 1055
rect 315 1054 316 1055
rect 438 1055 444 1056
rect 315 1052 381 1054
rect 315 1051 316 1052
rect 236 1046 238 1051
rect 310 1050 316 1051
rect 438 1051 439 1055
rect 443 1054 444 1055
rect 727 1055 733 1056
rect 727 1054 728 1055
rect 443 1052 525 1054
rect 669 1052 728 1054
rect 443 1051 444 1052
rect 438 1050 444 1051
rect 727 1051 728 1052
rect 732 1051 733 1055
rect 870 1055 876 1056
rect 870 1054 871 1055
rect 821 1052 871 1054
rect 727 1050 733 1051
rect 870 1051 871 1052
rect 875 1051 876 1055
rect 1026 1055 1032 1056
rect 1026 1054 1027 1055
rect 973 1052 1027 1054
rect 870 1050 876 1051
rect 1026 1051 1027 1052
rect 1031 1051 1032 1055
rect 1026 1050 1032 1051
rect 1114 1055 1120 1056
rect 1114 1051 1115 1055
rect 1119 1051 1120 1055
rect 1114 1050 1120 1051
rect 430 1047 436 1048
rect 430 1046 431 1047
rect 236 1044 431 1046
rect 430 1043 431 1044
rect 435 1043 436 1047
rect 430 1042 436 1043
rect 326 1039 332 1040
rect 326 1038 327 1039
rect 261 1036 327 1038
rect 326 1035 327 1036
rect 331 1035 332 1039
rect 471 1039 477 1040
rect 471 1038 472 1039
rect 413 1036 472 1038
rect 326 1034 332 1035
rect 471 1035 472 1036
rect 476 1035 477 1039
rect 471 1034 477 1035
rect 511 1039 517 1040
rect 511 1035 512 1039
rect 516 1038 517 1039
rect 722 1039 728 1040
rect 516 1036 565 1038
rect 516 1035 517 1036
rect 511 1034 517 1035
rect 722 1035 723 1039
rect 727 1035 728 1039
rect 722 1034 728 1035
rect 818 1039 824 1040
rect 818 1035 819 1039
rect 823 1038 824 1039
rect 1058 1039 1064 1040
rect 823 1036 893 1038
rect 823 1035 824 1036
rect 818 1034 824 1035
rect 1058 1035 1059 1039
rect 1063 1035 1064 1039
rect 1058 1034 1064 1035
rect 242 1022 248 1023
rect 242 1018 243 1022
rect 247 1018 248 1022
rect 394 1022 400 1023
rect 110 1017 116 1018
rect 242 1017 248 1018
rect 326 1019 332 1020
rect 110 1013 111 1017
rect 115 1013 116 1017
rect 326 1015 327 1019
rect 331 1018 332 1019
rect 383 1019 389 1020
rect 383 1018 384 1019
rect 331 1016 384 1018
rect 331 1015 332 1016
rect 326 1014 332 1015
rect 383 1015 384 1016
rect 388 1015 389 1019
rect 394 1018 395 1022
rect 399 1018 400 1022
rect 546 1022 552 1023
rect 394 1017 400 1018
rect 471 1019 477 1020
rect 383 1014 389 1015
rect 471 1015 472 1019
rect 476 1018 477 1019
rect 535 1019 541 1020
rect 535 1018 536 1019
rect 476 1016 536 1018
rect 476 1015 477 1016
rect 471 1014 477 1015
rect 535 1015 536 1016
rect 540 1015 541 1019
rect 546 1018 547 1022
rect 551 1018 552 1022
rect 546 1017 552 1018
rect 706 1022 712 1023
rect 706 1018 707 1022
rect 711 1018 712 1022
rect 706 1017 712 1018
rect 874 1022 880 1023
rect 874 1018 875 1022
rect 879 1018 880 1022
rect 874 1017 880 1018
rect 1042 1022 1048 1023
rect 1042 1018 1043 1022
rect 1047 1018 1048 1022
rect 1042 1017 1048 1018
rect 1182 1017 1188 1018
rect 535 1014 541 1015
rect 110 1012 116 1013
rect 1182 1013 1183 1017
rect 1187 1013 1188 1017
rect 1182 1012 1188 1013
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 110 994 116 995
rect 1182 999 1188 1000
rect 1182 995 1183 999
rect 1187 995 1188 999
rect 1182 994 1188 995
rect 310 991 316 992
rect 310 990 311 991
rect 289 988 311 990
rect 310 987 311 988
rect 315 987 316 991
rect 818 991 824 992
rect 818 990 819 991
rect 753 988 819 990
rect 310 986 316 987
rect 818 987 819 988
rect 823 987 824 991
rect 818 986 824 987
rect 834 991 840 992
rect 834 987 835 991
rect 839 990 840 991
rect 1114 991 1120 992
rect 1114 990 1115 991
rect 839 988 865 990
rect 1089 988 1115 990
rect 839 987 840 988
rect 834 986 840 987
rect 1114 987 1115 988
rect 1119 987 1120 991
rect 1114 986 1120 987
rect 238 981 244 982
rect 238 977 239 981
rect 243 977 244 981
rect 238 976 244 977
rect 390 981 396 982
rect 390 977 391 981
rect 395 977 396 981
rect 390 976 396 977
rect 542 981 548 982
rect 542 977 543 981
rect 547 977 548 981
rect 542 976 548 977
rect 702 981 708 982
rect 702 977 703 981
rect 707 977 708 981
rect 702 976 708 977
rect 870 981 876 982
rect 870 977 871 981
rect 875 977 876 981
rect 870 976 876 977
rect 1038 981 1044 982
rect 1038 977 1039 981
rect 1043 977 1044 981
rect 1038 976 1044 977
rect 326 951 332 952
rect 326 947 327 951
rect 331 947 332 951
rect 326 946 332 947
rect 438 951 444 952
rect 438 947 439 951
rect 443 947 444 951
rect 438 946 444 947
rect 558 951 564 952
rect 558 947 559 951
rect 563 947 564 951
rect 558 946 564 947
rect 686 951 692 952
rect 686 947 687 951
rect 691 947 692 951
rect 686 946 692 947
rect 814 951 820 952
rect 814 947 815 951
rect 819 947 820 951
rect 814 946 820 947
rect 950 951 956 952
rect 950 947 951 951
rect 955 947 956 951
rect 950 946 956 947
rect 1086 951 1092 952
rect 1086 947 1087 951
rect 1091 947 1092 951
rect 1086 946 1092 947
rect 399 943 405 944
rect 399 942 400 943
rect 377 940 400 942
rect 399 939 400 940
rect 404 939 405 943
rect 511 943 517 944
rect 511 942 512 943
rect 489 940 512 942
rect 399 938 405 939
rect 511 939 512 940
rect 516 939 517 943
rect 930 943 936 944
rect 930 942 931 943
rect 865 940 931 942
rect 511 938 517 939
rect 930 939 931 940
rect 935 939 936 943
rect 1058 943 1064 944
rect 1058 942 1059 943
rect 1001 940 1059 942
rect 930 938 936 939
rect 1058 939 1059 940
rect 1063 939 1064 943
rect 1058 938 1064 939
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 110 928 116 929
rect 1182 933 1188 934
rect 1182 929 1183 933
rect 1187 929 1188 933
rect 1182 928 1188 929
rect 110 915 116 916
rect 110 911 111 915
rect 115 911 116 915
rect 511 915 517 916
rect 511 911 512 915
rect 516 914 517 915
rect 551 915 557 916
rect 551 914 552 915
rect 516 912 552 914
rect 516 911 517 912
rect 110 910 116 911
rect 330 910 336 911
rect 330 906 331 910
rect 335 906 336 910
rect 330 905 336 906
rect 442 910 448 911
rect 511 910 517 911
rect 551 911 552 912
rect 556 911 557 915
rect 630 915 636 916
rect 630 911 631 915
rect 635 914 636 915
rect 679 915 685 916
rect 679 914 680 915
rect 635 912 680 914
rect 635 911 636 912
rect 551 910 557 911
rect 562 910 568 911
rect 630 910 636 911
rect 679 911 680 912
rect 684 911 685 915
rect 1023 915 1029 916
rect 1023 911 1024 915
rect 1028 914 1029 915
rect 1079 915 1085 916
rect 1079 914 1080 915
rect 1028 912 1080 914
rect 1028 911 1029 912
rect 679 910 685 911
rect 690 910 696 911
rect 442 906 443 910
rect 447 906 448 910
rect 442 905 448 906
rect 562 906 563 910
rect 567 906 568 910
rect 562 905 568 906
rect 690 906 691 910
rect 695 906 696 910
rect 690 905 696 906
rect 818 910 824 911
rect 818 906 819 910
rect 823 906 824 910
rect 818 905 824 906
rect 954 910 960 911
rect 1023 910 1029 911
rect 1079 911 1080 912
rect 1084 911 1085 915
rect 1182 915 1188 916
rect 1182 911 1183 915
rect 1187 911 1188 915
rect 1079 910 1085 911
rect 1090 910 1096 911
rect 1182 910 1188 911
rect 954 906 955 910
rect 959 906 960 910
rect 954 905 960 906
rect 1090 906 1091 910
rect 1095 906 1096 910
rect 1090 905 1096 906
rect 399 895 405 896
rect 399 891 400 895
rect 404 894 405 895
rect 630 895 636 896
rect 630 894 631 895
rect 404 892 461 894
rect 581 892 631 894
rect 404 891 405 892
rect 348 886 350 891
rect 399 890 405 891
rect 630 891 631 892
rect 635 891 636 895
rect 730 895 736 896
rect 730 894 731 895
rect 709 892 731 894
rect 630 890 636 891
rect 730 891 731 892
rect 735 891 736 895
rect 730 890 736 891
rect 834 895 840 896
rect 834 891 835 895
rect 839 891 840 895
rect 1023 895 1029 896
rect 1023 894 1024 895
rect 973 892 1024 894
rect 834 890 840 891
rect 1023 891 1024 892
rect 1028 891 1029 895
rect 1023 890 1029 891
rect 1070 895 1076 896
rect 1070 891 1071 895
rect 1075 894 1076 895
rect 1075 892 1109 894
rect 1075 891 1076 892
rect 1070 890 1076 891
rect 511 887 517 888
rect 511 886 512 887
rect 348 884 512 886
rect 511 883 512 884
rect 516 883 517 887
rect 511 882 517 883
rect 382 879 388 880
rect 382 875 383 879
rect 387 878 388 879
rect 474 879 480 880
rect 387 876 421 878
rect 387 875 388 876
rect 382 874 388 875
rect 474 875 475 879
rect 479 878 480 879
rect 582 879 588 880
rect 479 876 533 878
rect 479 875 480 876
rect 474 874 480 875
rect 582 875 583 879
rect 587 878 588 879
rect 711 879 717 880
rect 587 876 661 878
rect 587 875 588 876
rect 582 874 588 875
rect 711 875 712 879
rect 716 878 717 879
rect 930 879 936 880
rect 716 876 797 878
rect 716 875 717 876
rect 711 874 717 875
rect 930 875 931 879
rect 935 875 936 879
rect 930 874 936 875
rect 1039 879 1045 880
rect 1039 875 1040 879
rect 1044 878 1045 879
rect 1044 876 1077 878
rect 1044 875 1045 876
rect 1039 874 1045 875
rect 402 862 408 863
rect 402 858 403 862
rect 407 858 408 862
rect 110 857 116 858
rect 402 857 408 858
rect 514 862 520 863
rect 514 858 515 862
rect 519 858 520 862
rect 514 857 520 858
rect 642 862 648 863
rect 642 858 643 862
rect 647 858 648 862
rect 778 862 784 863
rect 642 857 648 858
rect 730 859 736 860
rect 110 853 111 857
rect 115 853 116 857
rect 730 855 731 859
rect 735 858 736 859
rect 767 859 773 860
rect 767 858 768 859
rect 735 856 768 858
rect 735 855 736 856
rect 730 854 736 855
rect 767 855 768 856
rect 772 855 773 859
rect 778 858 779 862
rect 783 858 784 862
rect 778 857 784 858
rect 914 862 920 863
rect 914 858 915 862
rect 919 858 920 862
rect 914 857 920 858
rect 1058 862 1064 863
rect 1058 858 1059 862
rect 1063 858 1064 862
rect 1058 857 1064 858
rect 1182 857 1188 858
rect 767 854 773 855
rect 110 852 116 853
rect 1182 853 1183 857
rect 1187 853 1188 857
rect 1182 852 1188 853
rect 110 839 116 840
rect 110 835 111 839
rect 115 835 116 839
rect 110 834 116 835
rect 1182 839 1188 840
rect 1182 835 1183 839
rect 1187 835 1188 839
rect 1182 834 1188 835
rect 474 831 480 832
rect 474 830 475 831
rect 449 828 475 830
rect 474 827 475 828
rect 479 827 480 831
rect 582 831 588 832
rect 582 830 583 831
rect 561 828 583 830
rect 474 826 480 827
rect 582 827 583 828
rect 587 827 588 831
rect 711 831 717 832
rect 711 830 712 831
rect 689 828 712 830
rect 582 826 588 827
rect 711 827 712 828
rect 716 827 717 831
rect 711 826 717 827
rect 902 831 908 832
rect 902 827 903 831
rect 907 827 908 831
rect 902 826 908 827
rect 1070 831 1076 832
rect 1070 827 1071 831
rect 1075 827 1076 831
rect 1070 826 1076 827
rect 398 821 404 822
rect 398 817 399 821
rect 403 817 404 821
rect 398 816 404 817
rect 510 821 516 822
rect 510 817 511 821
rect 515 817 516 821
rect 510 816 516 817
rect 638 821 644 822
rect 638 817 639 821
rect 643 817 644 821
rect 638 816 644 817
rect 774 821 780 822
rect 774 817 775 821
rect 779 817 780 821
rect 774 816 780 817
rect 910 821 916 822
rect 910 817 911 821
rect 915 817 916 821
rect 910 816 916 817
rect 1054 821 1060 822
rect 1054 817 1055 821
rect 1059 817 1060 821
rect 1054 816 1060 817
rect 374 799 380 800
rect 374 795 375 799
rect 379 795 380 799
rect 374 794 380 795
rect 518 799 524 800
rect 518 795 519 799
rect 523 795 524 799
rect 518 794 524 795
rect 662 799 668 800
rect 662 795 663 799
rect 667 795 668 799
rect 662 794 668 795
rect 814 799 820 800
rect 814 795 815 799
rect 819 795 820 799
rect 814 794 820 795
rect 966 799 972 800
rect 966 795 967 799
rect 971 795 972 799
rect 966 794 972 795
rect 1094 799 1100 800
rect 1094 795 1095 799
rect 1099 795 1100 799
rect 1094 794 1100 795
rect 922 791 928 792
rect 922 790 923 791
rect 865 788 923 790
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 922 787 923 788
rect 927 787 928 791
rect 1039 791 1045 792
rect 1039 790 1040 791
rect 1017 788 1040 790
rect 922 786 928 787
rect 1039 787 1040 788
rect 1044 787 1045 791
rect 1039 786 1045 787
rect 382 782 388 783
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 110 776 116 777
rect 1182 781 1188 782
rect 1182 777 1183 781
rect 1187 777 1188 781
rect 1182 776 1188 777
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 450 763 456 764
rect 450 759 451 763
rect 455 762 456 763
rect 511 763 517 764
rect 511 762 512 763
rect 455 760 512 762
rect 455 759 456 760
rect 110 758 116 759
rect 378 758 384 759
rect 450 758 456 759
rect 511 759 512 760
rect 516 759 517 763
rect 594 763 600 764
rect 594 759 595 763
rect 599 762 600 763
rect 655 763 661 764
rect 655 762 656 763
rect 599 760 656 762
rect 599 759 600 760
rect 511 758 517 759
rect 522 758 528 759
rect 594 758 600 759
rect 655 759 656 760
rect 660 759 661 763
rect 1038 763 1044 764
rect 1038 759 1039 763
rect 1043 762 1044 763
rect 1087 763 1093 764
rect 1087 762 1088 763
rect 1043 760 1088 762
rect 1043 759 1044 760
rect 655 758 661 759
rect 666 758 672 759
rect 378 754 379 758
rect 383 754 384 758
rect 378 753 384 754
rect 522 754 523 758
rect 527 754 528 758
rect 522 753 528 754
rect 666 754 667 758
rect 671 754 672 758
rect 666 753 672 754
rect 818 758 824 759
rect 818 754 819 758
rect 823 754 824 758
rect 818 753 824 754
rect 970 758 976 759
rect 1038 758 1044 759
rect 1087 759 1088 760
rect 1092 759 1093 763
rect 1182 763 1188 764
rect 1182 759 1183 763
rect 1187 759 1188 763
rect 1087 758 1093 759
rect 1098 758 1104 759
rect 1182 758 1188 759
rect 970 754 971 758
rect 975 754 976 758
rect 970 753 976 754
rect 1098 754 1099 758
rect 1103 754 1104 758
rect 1098 753 1104 754
rect 450 743 456 744
rect 450 742 451 743
rect 397 740 451 742
rect 450 739 451 740
rect 455 739 456 743
rect 594 743 600 744
rect 594 742 595 743
rect 541 740 595 742
rect 450 738 456 739
rect 594 739 595 740
rect 599 739 600 743
rect 594 738 600 739
rect 682 743 688 744
rect 682 739 683 743
rect 687 739 688 743
rect 902 743 908 744
rect 902 742 903 743
rect 837 740 903 742
rect 682 738 688 739
rect 902 739 903 740
rect 907 739 908 743
rect 1038 743 1044 744
rect 1038 742 1039 743
rect 989 740 1039 742
rect 902 738 908 739
rect 1038 739 1039 740
rect 1043 739 1044 743
rect 1038 738 1044 739
rect 1114 743 1120 744
rect 1114 739 1115 743
rect 1119 739 1120 743
rect 1114 738 1120 739
rect 162 731 168 732
rect 162 727 163 731
rect 167 727 168 731
rect 162 726 168 727
rect 214 731 220 732
rect 214 727 215 731
rect 219 730 220 731
rect 358 731 364 732
rect 219 728 285 730
rect 219 727 220 728
rect 214 726 220 727
rect 358 727 359 731
rect 363 730 364 731
rect 487 731 493 732
rect 363 728 429 730
rect 363 727 364 728
rect 358 726 364 727
rect 487 727 488 731
rect 492 730 493 731
rect 647 731 653 732
rect 492 728 581 730
rect 492 727 493 728
rect 487 726 493 727
rect 647 727 648 731
rect 652 730 653 731
rect 922 731 928 732
rect 652 728 749 730
rect 652 727 653 728
rect 647 726 653 727
rect 922 727 923 731
rect 927 727 928 731
rect 922 726 928 727
rect 1106 731 1112 732
rect 1106 727 1107 731
rect 1111 727 1112 731
rect 1106 726 1112 727
rect 146 714 152 715
rect 146 710 147 714
rect 151 710 152 714
rect 110 709 116 710
rect 146 709 152 710
rect 266 714 272 715
rect 266 710 267 714
rect 271 710 272 714
rect 266 709 272 710
rect 410 714 416 715
rect 410 710 411 714
rect 415 710 416 714
rect 410 709 416 710
rect 562 714 568 715
rect 562 710 563 714
rect 567 710 568 714
rect 730 714 736 715
rect 562 709 568 710
rect 682 711 688 712
rect 110 705 111 709
rect 115 705 116 709
rect 682 707 683 711
rect 687 710 688 711
rect 719 711 725 712
rect 719 710 720 711
rect 687 708 720 710
rect 687 707 688 708
rect 682 706 688 707
rect 719 707 720 708
rect 724 707 725 711
rect 730 710 731 714
rect 735 710 736 714
rect 730 709 736 710
rect 906 714 912 715
rect 906 710 907 714
rect 911 710 912 714
rect 906 709 912 710
rect 1090 714 1096 715
rect 1090 710 1091 714
rect 1095 710 1096 714
rect 1090 709 1096 710
rect 1182 709 1188 710
rect 719 706 725 707
rect 110 704 116 705
rect 1182 705 1183 709
rect 1187 705 1188 709
rect 1182 704 1188 705
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 110 686 116 687
rect 1182 691 1188 692
rect 1182 687 1183 691
rect 1187 687 1188 691
rect 1182 686 1188 687
rect 214 683 220 684
rect 214 682 215 683
rect 193 680 215 682
rect 214 679 215 680
rect 219 679 220 683
rect 358 683 364 684
rect 358 682 359 683
rect 313 680 359 682
rect 214 678 220 679
rect 358 679 359 680
rect 363 679 364 683
rect 487 683 493 684
rect 487 682 488 683
rect 457 680 488 682
rect 358 678 364 679
rect 487 679 488 680
rect 492 679 493 683
rect 647 683 653 684
rect 647 682 648 683
rect 609 680 648 682
rect 487 678 493 679
rect 647 679 648 680
rect 652 679 653 683
rect 647 678 653 679
rect 922 683 928 684
rect 922 679 923 683
rect 927 679 928 683
rect 922 678 928 679
rect 1110 683 1116 684
rect 1110 679 1111 683
rect 1115 679 1116 683
rect 1110 678 1116 679
rect 142 673 148 674
rect 142 669 143 673
rect 147 669 148 673
rect 142 668 148 669
rect 262 673 268 674
rect 262 669 263 673
rect 267 669 268 673
rect 262 668 268 669
rect 406 673 412 674
rect 406 669 407 673
rect 411 669 412 673
rect 406 668 412 669
rect 558 673 564 674
rect 558 669 559 673
rect 563 669 564 673
rect 558 668 564 669
rect 726 673 732 674
rect 726 669 727 673
rect 731 669 732 673
rect 726 668 732 669
rect 902 673 908 674
rect 902 669 903 673
rect 907 669 908 673
rect 902 668 908 669
rect 1086 673 1092 674
rect 1086 669 1087 673
rect 1091 669 1092 673
rect 1086 668 1092 669
rect 142 643 148 644
rect 142 639 143 643
rect 147 639 148 643
rect 142 638 148 639
rect 246 643 252 644
rect 246 639 247 643
rect 251 639 252 643
rect 246 638 252 639
rect 390 643 396 644
rect 390 639 391 643
rect 395 639 396 643
rect 390 638 396 639
rect 550 643 556 644
rect 550 639 551 643
rect 555 639 556 643
rect 550 638 556 639
rect 718 643 724 644
rect 718 639 719 643
rect 723 639 724 643
rect 718 638 724 639
rect 902 643 908 644
rect 902 639 903 643
rect 907 639 908 643
rect 902 638 908 639
rect 1086 643 1092 644
rect 1086 639 1087 643
rect 1091 639 1092 643
rect 1086 638 1092 639
rect 639 635 645 636
rect 639 634 640 635
rect 601 632 640 634
rect 162 631 168 632
rect 162 627 163 631
rect 167 627 168 631
rect 639 631 640 632
rect 644 631 645 635
rect 639 630 645 631
rect 914 631 920 632
rect 162 626 168 627
rect 914 627 915 631
rect 919 627 920 631
rect 914 626 920 627
rect 1102 631 1108 632
rect 1102 627 1103 631
rect 1107 627 1108 631
rect 1102 626 1108 627
rect 110 625 116 626
rect 110 621 111 625
rect 115 621 116 625
rect 110 620 116 621
rect 1182 625 1188 626
rect 1182 621 1183 625
rect 1187 621 1188 625
rect 1182 620 1188 621
rect 110 607 116 608
rect 110 603 111 607
rect 115 603 116 607
rect 214 607 220 608
rect 214 603 215 607
rect 219 606 220 607
rect 239 607 245 608
rect 239 606 240 607
rect 219 604 240 606
rect 219 603 220 604
rect 110 602 116 603
rect 146 602 152 603
rect 214 602 220 603
rect 239 603 240 604
rect 244 603 245 607
rect 330 607 336 608
rect 330 603 331 607
rect 335 606 336 607
rect 383 607 389 608
rect 383 606 384 607
rect 335 604 384 606
rect 335 603 336 604
rect 239 602 245 603
rect 250 602 256 603
rect 330 602 336 603
rect 383 603 384 604
rect 388 603 389 607
rect 622 607 628 608
rect 622 603 623 607
rect 627 606 628 607
rect 711 607 717 608
rect 711 606 712 607
rect 627 604 712 606
rect 627 603 628 604
rect 383 602 389 603
rect 394 602 400 603
rect 146 598 147 602
rect 151 598 152 602
rect 146 597 152 598
rect 250 598 251 602
rect 255 598 256 602
rect 250 597 256 598
rect 394 598 395 602
rect 399 598 400 602
rect 394 597 400 598
rect 554 602 560 603
rect 622 602 628 603
rect 711 603 712 604
rect 716 603 717 607
rect 1182 607 1188 608
rect 1182 603 1183 607
rect 1187 603 1188 607
rect 711 602 717 603
rect 722 602 728 603
rect 554 598 555 602
rect 559 598 560 602
rect 554 597 560 598
rect 722 598 723 602
rect 727 598 728 602
rect 722 597 728 598
rect 906 602 912 603
rect 906 598 907 602
rect 911 598 912 602
rect 906 597 912 598
rect 1090 602 1096 603
rect 1182 602 1188 603
rect 1090 598 1091 602
rect 1095 598 1096 602
rect 1090 597 1096 598
rect 214 587 220 588
rect 214 586 215 587
rect 165 584 215 586
rect 214 583 215 584
rect 219 583 220 587
rect 330 587 336 588
rect 330 586 331 587
rect 269 584 331 586
rect 214 582 220 583
rect 330 583 331 584
rect 335 583 336 587
rect 330 582 336 583
rect 410 587 416 588
rect 410 583 411 587
rect 415 583 416 587
rect 410 582 416 583
rect 570 587 576 588
rect 570 583 571 587
rect 575 583 576 587
rect 570 582 576 583
rect 639 587 645 588
rect 639 583 640 587
rect 644 586 645 587
rect 922 587 928 588
rect 644 584 741 586
rect 644 583 645 584
rect 639 582 645 583
rect 922 583 923 587
rect 927 583 928 587
rect 922 582 928 583
rect 1098 587 1104 588
rect 1098 583 1099 587
rect 1103 586 1104 587
rect 1103 584 1109 586
rect 1103 583 1104 584
rect 1098 582 1104 583
rect 282 575 288 576
rect 282 571 283 575
rect 287 571 288 575
rect 282 570 288 571
rect 354 575 360 576
rect 354 571 355 575
rect 359 574 360 575
rect 458 575 464 576
rect 359 572 397 574
rect 359 571 360 572
rect 354 570 360 571
rect 458 571 459 575
rect 463 574 464 575
rect 706 575 712 576
rect 706 574 707 575
rect 463 572 517 574
rect 653 572 707 574
rect 463 571 464 572
rect 458 570 464 571
rect 706 571 707 572
rect 711 571 712 575
rect 822 575 828 576
rect 822 574 823 575
rect 797 572 823 574
rect 706 570 712 571
rect 822 571 823 572
rect 827 571 828 575
rect 822 570 828 571
rect 914 575 920 576
rect 914 571 915 575
rect 919 574 920 575
rect 1078 575 1084 576
rect 919 572 949 574
rect 919 571 920 572
rect 914 570 920 571
rect 1078 571 1079 575
rect 1083 574 1084 575
rect 1083 572 1109 574
rect 1083 571 1084 572
rect 1078 570 1084 571
rect 266 558 272 559
rect 266 554 267 558
rect 271 554 272 558
rect 110 553 116 554
rect 266 553 272 554
rect 378 558 384 559
rect 378 554 379 558
rect 383 554 384 558
rect 378 553 384 554
rect 498 558 504 559
rect 498 554 499 558
rect 503 554 504 558
rect 634 558 640 559
rect 498 553 504 554
rect 578 555 584 556
rect 110 549 111 553
rect 115 549 116 553
rect 578 551 579 555
rect 583 554 584 555
rect 623 555 629 556
rect 623 554 624 555
rect 583 552 624 554
rect 583 551 584 552
rect 578 550 584 551
rect 623 551 624 552
rect 628 551 629 555
rect 634 554 635 558
rect 639 554 640 558
rect 778 558 784 559
rect 634 553 640 554
rect 706 555 712 556
rect 623 550 629 551
rect 706 551 707 555
rect 711 554 712 555
rect 767 555 773 556
rect 767 554 768 555
rect 711 552 768 554
rect 711 551 712 552
rect 706 550 712 551
rect 767 551 768 552
rect 772 551 773 555
rect 778 554 779 558
rect 783 554 784 558
rect 778 553 784 554
rect 930 558 936 559
rect 930 554 931 558
rect 935 554 936 558
rect 930 553 936 554
rect 1090 558 1096 559
rect 1090 554 1091 558
rect 1095 554 1096 558
rect 1090 553 1096 554
rect 1182 553 1188 554
rect 767 550 773 551
rect 110 548 116 549
rect 1182 549 1183 553
rect 1187 549 1188 553
rect 1182 548 1188 549
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 1182 535 1188 536
rect 1182 531 1183 535
rect 1187 531 1188 535
rect 1182 530 1188 531
rect 354 527 360 528
rect 354 526 355 527
rect 313 524 355 526
rect 354 523 355 524
rect 359 523 360 527
rect 458 527 464 528
rect 458 526 459 527
rect 425 524 459 526
rect 354 522 360 523
rect 458 523 459 524
rect 463 523 464 527
rect 570 527 576 528
rect 570 526 571 527
rect 545 524 571 526
rect 458 522 464 523
rect 570 523 571 524
rect 575 523 576 527
rect 570 522 576 523
rect 938 527 944 528
rect 938 523 939 527
rect 943 523 944 527
rect 938 522 944 523
rect 1098 527 1104 528
rect 1098 523 1099 527
rect 1103 523 1104 527
rect 1098 522 1104 523
rect 262 517 268 518
rect 262 513 263 517
rect 267 513 268 517
rect 262 512 268 513
rect 374 517 380 518
rect 374 513 375 517
rect 379 513 380 517
rect 374 512 380 513
rect 494 517 500 518
rect 494 513 495 517
rect 499 513 500 517
rect 494 512 500 513
rect 630 517 636 518
rect 630 513 631 517
rect 635 513 636 517
rect 630 512 636 513
rect 774 517 780 518
rect 774 513 775 517
rect 779 513 780 517
rect 774 512 780 513
rect 926 517 932 518
rect 926 513 927 517
rect 931 513 932 517
rect 926 512 932 513
rect 1086 517 1092 518
rect 1086 513 1087 517
rect 1091 513 1092 517
rect 1086 512 1092 513
rect 806 499 812 500
rect 806 495 807 499
rect 811 498 812 499
rect 910 499 916 500
rect 910 498 911 499
rect 811 496 911 498
rect 811 495 812 496
rect 806 494 812 495
rect 910 495 911 496
rect 915 495 916 499
rect 910 494 916 495
rect 462 487 468 488
rect 462 483 463 487
rect 467 483 468 487
rect 462 482 468 483
rect 550 487 556 488
rect 550 483 551 487
rect 555 483 556 487
rect 550 482 556 483
rect 638 487 644 488
rect 638 483 639 487
rect 643 483 644 487
rect 638 482 644 483
rect 734 487 740 488
rect 734 483 735 487
rect 739 483 740 487
rect 734 482 740 483
rect 830 487 836 488
rect 830 483 831 487
rect 835 483 836 487
rect 830 482 836 483
rect 918 487 924 488
rect 918 483 919 487
rect 923 483 924 487
rect 918 482 924 483
rect 1006 487 1012 488
rect 1006 483 1007 487
rect 1011 483 1012 487
rect 1006 482 1012 483
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 483 1100 487
rect 1094 482 1100 483
rect 711 479 717 480
rect 711 478 712 479
rect 513 476 538 478
rect 601 476 626 478
rect 689 476 712 478
rect 534 475 540 476
rect 534 471 535 475
rect 539 471 540 475
rect 534 470 540 471
rect 622 475 628 476
rect 622 471 623 475
rect 627 471 628 475
rect 711 475 712 476
rect 716 475 717 479
rect 807 479 813 480
rect 807 478 808 479
rect 785 476 808 478
rect 711 474 717 475
rect 807 475 808 476
rect 812 475 813 479
rect 807 474 813 475
rect 822 479 828 480
rect 822 475 823 479
rect 827 475 828 479
rect 822 474 828 475
rect 910 479 916 480
rect 910 475 911 479
rect 915 475 916 479
rect 1057 476 1082 478
rect 910 474 916 475
rect 1078 475 1084 476
rect 622 470 628 471
rect 1078 471 1079 475
rect 1083 471 1084 475
rect 1078 470 1084 471
rect 110 469 116 470
rect 110 465 111 469
rect 115 465 116 469
rect 110 464 116 465
rect 1182 469 1188 470
rect 1182 465 1183 469
rect 1187 465 1188 469
rect 1182 464 1188 465
rect 110 451 116 452
rect 110 447 111 451
rect 115 447 116 451
rect 1078 451 1084 452
rect 1078 447 1079 451
rect 1083 450 1084 451
rect 1087 451 1093 452
rect 1087 450 1088 451
rect 1083 448 1088 450
rect 1083 447 1084 448
rect 110 446 116 447
rect 466 446 472 447
rect 466 442 467 446
rect 471 442 472 446
rect 466 441 472 442
rect 554 446 560 447
rect 554 442 555 446
rect 559 442 560 446
rect 554 441 560 442
rect 642 446 648 447
rect 642 442 643 446
rect 647 442 648 446
rect 642 441 648 442
rect 738 446 744 447
rect 738 442 739 446
rect 743 442 744 446
rect 738 441 744 442
rect 834 446 840 447
rect 834 442 835 446
rect 839 442 840 446
rect 834 441 840 442
rect 922 446 928 447
rect 922 442 923 446
rect 927 442 928 446
rect 922 441 928 442
rect 1010 446 1016 447
rect 1078 446 1084 447
rect 1087 447 1088 448
rect 1092 447 1093 451
rect 1182 451 1188 452
rect 1182 447 1183 451
rect 1187 447 1188 451
rect 1087 446 1093 447
rect 1098 446 1104 447
rect 1182 446 1188 447
rect 1010 442 1011 446
rect 1015 442 1016 446
rect 1010 441 1016 442
rect 1098 442 1099 446
rect 1103 442 1104 446
rect 1098 441 1104 442
rect 534 431 540 432
rect 534 427 535 431
rect 539 430 540 431
rect 622 431 628 432
rect 539 428 573 430
rect 539 427 540 428
rect 484 422 486 427
rect 534 426 540 427
rect 622 427 623 431
rect 627 430 628 431
rect 711 431 717 432
rect 627 428 661 430
rect 627 427 628 428
rect 622 426 628 427
rect 711 427 712 431
rect 716 430 717 431
rect 807 431 813 432
rect 716 428 757 430
rect 716 427 717 428
rect 711 426 717 427
rect 807 427 808 431
rect 812 430 813 431
rect 938 431 944 432
rect 812 428 853 430
rect 812 427 813 428
rect 807 426 813 427
rect 938 427 939 431
rect 943 427 944 431
rect 1078 431 1084 432
rect 1078 430 1079 431
rect 1029 428 1079 430
rect 938 426 944 427
rect 1078 427 1079 428
rect 1083 427 1084 431
rect 1078 426 1084 427
rect 1106 431 1112 432
rect 1106 427 1107 431
rect 1111 430 1112 431
rect 1111 428 1117 430
rect 1111 427 1112 428
rect 1106 426 1112 427
rect 622 423 628 424
rect 622 422 623 423
rect 484 420 623 422
rect 454 419 460 420
rect 454 418 455 419
rect 413 416 455 418
rect 454 415 455 416
rect 459 415 460 419
rect 622 419 623 420
rect 627 419 628 423
rect 622 418 628 419
rect 806 419 812 420
rect 806 418 807 419
rect 454 414 460 415
rect 464 416 501 418
rect 552 416 589 418
rect 640 416 677 418
rect 765 416 807 418
rect 464 412 466 416
rect 552 412 554 416
rect 640 412 642 416
rect 806 415 807 416
rect 811 415 812 419
rect 806 414 812 415
rect 814 419 820 420
rect 814 415 815 419
rect 819 418 820 419
rect 938 419 944 420
rect 819 416 853 418
rect 819 415 820 416
rect 814 414 820 415
rect 938 415 939 419
rect 943 415 944 419
rect 938 414 944 415
rect 990 419 996 420
rect 990 415 991 419
rect 995 418 996 419
rect 1078 419 1084 420
rect 995 416 1029 418
rect 995 415 996 416
rect 990 414 996 415
rect 1078 415 1079 419
rect 1083 418 1084 419
rect 1083 416 1117 418
rect 1083 415 1084 416
rect 1078 414 1084 415
rect 462 411 468 412
rect 462 407 463 411
rect 467 407 468 411
rect 462 406 468 407
rect 550 411 556 412
rect 550 407 551 411
rect 555 407 556 411
rect 550 406 556 407
rect 638 411 644 412
rect 638 407 639 411
rect 643 407 644 411
rect 638 406 644 407
rect 394 402 400 403
rect 394 398 395 402
rect 399 398 400 402
rect 110 397 116 398
rect 394 397 400 398
rect 482 402 488 403
rect 482 398 483 402
rect 487 398 488 402
rect 482 397 488 398
rect 570 402 576 403
rect 570 398 571 402
rect 575 398 576 402
rect 570 397 576 398
rect 658 402 664 403
rect 658 398 659 402
rect 663 398 664 402
rect 658 397 664 398
rect 746 402 752 403
rect 746 398 747 402
rect 751 398 752 402
rect 746 397 752 398
rect 834 402 840 403
rect 834 398 835 402
rect 839 398 840 402
rect 834 397 840 398
rect 922 402 928 403
rect 922 398 923 402
rect 927 398 928 402
rect 922 397 928 398
rect 1010 402 1016 403
rect 1010 398 1011 402
rect 1015 398 1016 402
rect 1010 397 1016 398
rect 1098 402 1104 403
rect 1098 398 1099 402
rect 1103 398 1104 402
rect 1098 397 1104 398
rect 1182 397 1188 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 1182 393 1183 397
rect 1187 393 1188 397
rect 1182 392 1188 393
rect 622 387 628 388
rect 622 383 623 387
rect 627 386 628 387
rect 647 387 653 388
rect 647 386 648 387
rect 627 384 648 386
rect 627 383 628 384
rect 622 382 628 383
rect 647 383 648 384
rect 652 383 653 387
rect 647 382 653 383
rect 110 379 116 380
rect 110 375 111 379
rect 115 375 116 379
rect 110 374 116 375
rect 1182 379 1188 380
rect 1182 375 1183 379
rect 1187 375 1188 379
rect 1182 374 1188 375
rect 462 371 468 372
rect 462 370 463 371
rect 441 368 463 370
rect 462 367 463 368
rect 467 367 468 371
rect 550 371 556 372
rect 550 370 551 371
rect 529 368 551 370
rect 462 366 468 367
rect 550 367 551 368
rect 555 367 556 371
rect 638 371 644 372
rect 638 370 639 371
rect 617 368 639 370
rect 550 366 556 367
rect 638 367 639 368
rect 643 367 644 371
rect 814 371 820 372
rect 814 370 815 371
rect 793 368 815 370
rect 638 366 644 367
rect 814 367 815 368
rect 819 367 820 371
rect 902 371 908 372
rect 902 370 903 371
rect 881 368 903 370
rect 814 366 820 367
rect 902 367 903 368
rect 907 367 908 371
rect 990 371 996 372
rect 990 370 991 371
rect 969 368 991 370
rect 902 366 908 367
rect 990 367 991 368
rect 995 367 996 371
rect 1078 371 1084 372
rect 1078 370 1079 371
rect 1057 368 1079 370
rect 990 366 996 367
rect 1078 367 1079 368
rect 1083 367 1084 371
rect 1078 366 1084 367
rect 1106 371 1112 372
rect 1106 367 1107 371
rect 1111 367 1112 371
rect 1106 366 1112 367
rect 390 361 396 362
rect 390 357 391 361
rect 395 357 396 361
rect 390 356 396 357
rect 478 361 484 362
rect 478 357 479 361
rect 483 357 484 361
rect 478 356 484 357
rect 566 361 572 362
rect 566 357 567 361
rect 571 357 572 361
rect 566 356 572 357
rect 654 361 660 362
rect 654 357 655 361
rect 659 357 660 361
rect 654 356 660 357
rect 742 361 748 362
rect 742 357 743 361
rect 747 357 748 361
rect 742 356 748 357
rect 830 361 836 362
rect 830 357 831 361
rect 835 357 836 361
rect 830 356 836 357
rect 918 361 924 362
rect 918 357 919 361
rect 923 357 924 361
rect 918 356 924 357
rect 1006 361 1012 362
rect 1006 357 1007 361
rect 1011 357 1012 361
rect 1006 356 1012 357
rect 1094 361 1100 362
rect 1094 357 1095 361
rect 1099 357 1100 361
rect 1094 356 1100 357
rect 366 339 372 340
rect 366 335 367 339
rect 371 335 372 339
rect 366 334 372 335
rect 478 339 484 340
rect 478 335 479 339
rect 483 335 484 339
rect 478 334 484 335
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 726 339 732 340
rect 726 335 727 339
rect 731 335 732 339
rect 726 334 732 335
rect 862 339 868 340
rect 862 335 863 339
rect 867 335 868 339
rect 862 334 868 335
rect 1006 339 1012 340
rect 1006 335 1007 339
rect 1011 335 1012 339
rect 1006 334 1012 335
rect 439 331 445 332
rect 439 330 440 331
rect 417 328 440 330
rect 439 327 440 328
rect 444 327 445 331
rect 551 331 557 332
rect 551 330 552 331
rect 529 328 552 330
rect 439 326 445 327
rect 551 327 552 328
rect 556 327 557 331
rect 671 331 677 332
rect 671 330 672 331
rect 649 328 672 330
rect 551 326 557 327
rect 671 327 672 328
rect 676 327 677 331
rect 799 331 805 332
rect 799 330 800 331
rect 777 328 800 330
rect 671 326 677 327
rect 799 327 800 328
rect 804 327 805 331
rect 799 326 805 327
rect 854 331 860 332
rect 854 327 855 331
rect 859 327 860 331
rect 854 326 860 327
rect 938 331 944 332
rect 938 327 939 331
rect 943 330 944 331
rect 943 328 1001 330
rect 943 327 944 328
rect 938 326 944 327
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 110 316 116 317
rect 1182 321 1188 322
rect 1182 317 1183 321
rect 1187 317 1188 321
rect 1182 316 1188 317
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 1182 303 1188 304
rect 1182 299 1183 303
rect 1187 299 1188 303
rect 110 298 116 299
rect 370 298 376 299
rect 370 294 371 298
rect 375 294 376 298
rect 370 293 376 294
rect 482 298 488 299
rect 482 294 483 298
rect 487 294 488 298
rect 482 293 488 294
rect 602 298 608 299
rect 602 294 603 298
rect 607 294 608 298
rect 602 293 608 294
rect 730 298 736 299
rect 730 294 731 298
rect 735 294 736 298
rect 730 293 736 294
rect 866 298 872 299
rect 866 294 867 298
rect 871 294 872 298
rect 866 293 872 294
rect 1010 298 1016 299
rect 1182 298 1188 299
rect 1010 294 1011 298
rect 1015 294 1016 298
rect 1010 293 1016 294
rect 439 283 445 284
rect 439 279 440 283
rect 444 282 445 283
rect 551 283 557 284
rect 444 280 501 282
rect 444 279 445 280
rect 388 274 390 279
rect 439 278 445 279
rect 551 279 552 283
rect 556 282 557 283
rect 671 283 677 284
rect 556 280 621 282
rect 556 279 557 280
rect 551 278 557 279
rect 671 279 672 283
rect 676 282 677 283
rect 799 283 805 284
rect 676 280 749 282
rect 676 279 677 280
rect 671 278 677 279
rect 799 279 800 283
rect 804 282 805 283
rect 902 283 908 284
rect 804 280 885 282
rect 804 279 805 280
rect 799 278 805 279
rect 902 279 903 283
rect 907 282 908 283
rect 907 280 1029 282
rect 907 279 908 280
rect 902 278 908 279
rect 535 275 541 276
rect 535 274 536 275
rect 388 272 536 274
rect 535 271 536 272
rect 540 271 541 275
rect 535 270 541 271
rect 218 263 224 264
rect 218 259 219 263
rect 223 259 224 263
rect 218 258 224 259
rect 270 263 276 264
rect 270 259 271 263
rect 275 262 276 263
rect 358 263 364 264
rect 275 260 309 262
rect 275 259 276 260
rect 270 258 276 259
rect 358 259 359 263
rect 363 262 364 263
rect 446 263 452 264
rect 363 260 397 262
rect 363 259 364 260
rect 358 258 364 259
rect 446 259 447 263
rect 451 262 452 263
rect 534 263 540 264
rect 451 260 485 262
rect 451 259 452 260
rect 446 258 452 259
rect 534 259 535 263
rect 539 262 540 263
rect 539 260 573 262
rect 539 259 540 260
rect 534 258 540 259
rect 202 246 208 247
rect 202 242 203 246
rect 207 242 208 246
rect 110 241 116 242
rect 202 241 208 242
rect 290 246 296 247
rect 290 242 291 246
rect 295 242 296 246
rect 290 241 296 242
rect 378 246 384 247
rect 378 242 379 246
rect 383 242 384 246
rect 378 241 384 242
rect 466 246 472 247
rect 466 242 467 246
rect 471 242 472 246
rect 554 246 560 247
rect 466 241 472 242
rect 535 243 541 244
rect 110 237 111 241
rect 115 237 116 241
rect 535 239 536 243
rect 540 242 541 243
rect 543 243 549 244
rect 543 242 544 243
rect 540 240 544 242
rect 540 239 541 240
rect 535 238 541 239
rect 543 239 544 240
rect 548 239 549 243
rect 554 242 555 246
rect 559 242 560 246
rect 554 241 560 242
rect 1182 241 1188 242
rect 543 238 549 239
rect 110 236 116 237
rect 1182 237 1183 241
rect 1187 237 1188 241
rect 1182 236 1188 237
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 110 218 116 219
rect 1182 223 1188 224
rect 1182 219 1183 223
rect 1187 219 1188 223
rect 1182 218 1188 219
rect 270 215 276 216
rect 270 214 271 215
rect 249 212 271 214
rect 270 211 271 212
rect 275 211 276 215
rect 358 215 364 216
rect 358 214 359 215
rect 337 212 359 214
rect 270 210 276 211
rect 358 211 359 212
rect 363 211 364 215
rect 446 215 452 216
rect 446 214 447 215
rect 425 212 447 214
rect 358 210 364 211
rect 446 211 447 212
rect 451 211 452 215
rect 534 215 540 216
rect 534 214 535 215
rect 513 212 535 214
rect 446 210 452 211
rect 534 211 535 212
rect 539 211 540 215
rect 534 210 540 211
rect 198 205 204 206
rect 198 201 199 205
rect 203 201 204 205
rect 198 200 204 201
rect 286 205 292 206
rect 286 201 287 205
rect 291 201 292 205
rect 286 200 292 201
rect 374 205 380 206
rect 374 201 375 205
rect 379 201 380 205
rect 374 200 380 201
rect 462 205 468 206
rect 462 201 463 205
rect 467 201 468 205
rect 462 200 468 201
rect 550 205 556 206
rect 550 201 551 205
rect 555 201 556 205
rect 550 200 556 201
rect 218 191 224 192
rect 218 187 219 191
rect 223 190 224 191
rect 750 191 756 192
rect 750 190 751 191
rect 223 188 751 190
rect 223 187 224 188
rect 218 186 224 187
rect 750 187 751 188
rect 755 187 756 191
rect 750 186 756 187
rect 142 155 148 156
rect 142 151 143 155
rect 147 151 148 155
rect 142 150 148 151
rect 230 155 236 156
rect 230 151 231 155
rect 235 151 236 155
rect 230 150 236 151
rect 318 155 324 156
rect 318 151 319 155
rect 323 151 324 155
rect 318 150 324 151
rect 406 155 412 156
rect 406 151 407 155
rect 411 151 412 155
rect 406 150 412 151
rect 494 155 500 156
rect 494 151 495 155
rect 499 151 500 155
rect 494 150 500 151
rect 582 155 588 156
rect 582 151 583 155
rect 587 151 588 155
rect 582 150 588 151
rect 670 155 676 156
rect 670 151 671 155
rect 675 151 676 155
rect 670 150 676 151
rect 758 155 764 156
rect 758 151 759 155
rect 763 151 764 155
rect 758 150 764 151
rect 215 147 221 148
rect 215 146 216 147
rect 193 144 216 146
rect 215 143 216 144
rect 220 143 221 147
rect 303 147 309 148
rect 303 146 304 147
rect 281 144 304 146
rect 215 142 221 143
rect 303 143 304 144
rect 308 143 309 147
rect 750 147 756 148
rect 369 144 394 146
rect 457 144 482 146
rect 545 144 570 146
rect 633 144 658 146
rect 721 144 746 146
rect 303 142 309 143
rect 390 143 396 144
rect 390 139 391 143
rect 395 139 396 143
rect 390 138 396 139
rect 478 143 484 144
rect 478 139 479 143
rect 483 139 484 143
rect 478 138 484 139
rect 566 143 572 144
rect 566 139 567 143
rect 571 139 572 143
rect 566 138 572 139
rect 654 143 660 144
rect 654 139 655 143
rect 659 139 660 143
rect 654 138 660 139
rect 742 143 748 144
rect 742 139 743 143
rect 747 139 748 143
rect 750 143 751 147
rect 755 143 756 147
rect 750 142 756 143
rect 742 138 748 139
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 110 132 116 133
rect 1182 137 1188 138
rect 1182 133 1183 137
rect 1187 133 1188 137
rect 1182 132 1188 133
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 1182 119 1188 120
rect 1182 115 1183 119
rect 1187 115 1188 119
rect 110 114 116 115
rect 146 114 152 115
rect 146 110 147 114
rect 151 110 152 114
rect 146 109 152 110
rect 234 114 240 115
rect 234 110 235 114
rect 239 110 240 114
rect 234 109 240 110
rect 322 114 328 115
rect 322 110 323 114
rect 327 110 328 114
rect 322 109 328 110
rect 410 114 416 115
rect 410 110 411 114
rect 415 110 416 114
rect 410 109 416 110
rect 498 114 504 115
rect 498 110 499 114
rect 503 110 504 114
rect 498 109 504 110
rect 586 114 592 115
rect 586 110 587 114
rect 591 110 592 114
rect 586 109 592 110
rect 674 114 680 115
rect 674 110 675 114
rect 679 110 680 114
rect 674 109 680 110
rect 762 114 768 115
rect 1182 114 1188 115
rect 762 110 763 114
rect 767 110 768 114
rect 762 109 768 110
rect 215 99 221 100
rect 215 95 216 99
rect 220 98 221 99
rect 303 99 309 100
rect 220 96 253 98
rect 220 95 221 96
rect 215 94 221 95
rect 303 95 304 99
rect 308 98 309 99
rect 390 99 396 100
rect 308 96 341 98
rect 308 95 309 96
rect 303 94 309 95
rect 390 95 391 99
rect 395 98 396 99
rect 478 99 484 100
rect 395 96 429 98
rect 395 95 396 96
rect 390 94 396 95
rect 478 95 479 99
rect 483 98 484 99
rect 566 99 572 100
rect 483 96 517 98
rect 483 95 484 96
rect 478 94 484 95
rect 566 95 567 99
rect 571 98 572 99
rect 654 99 660 100
rect 571 96 605 98
rect 571 95 572 96
rect 566 94 572 95
rect 654 95 655 99
rect 659 98 660 99
rect 742 99 748 100
rect 659 96 693 98
rect 659 95 660 96
rect 654 94 660 95
rect 742 95 743 99
rect 747 98 748 99
rect 747 96 781 98
rect 747 95 748 96
rect 742 94 748 95
<< m3c >>
rect 575 1267 579 1271
rect 683 1259 687 1263
rect 111 1249 115 1253
rect 1183 1249 1187 1253
rect 111 1231 115 1235
rect 1183 1231 1187 1235
rect 579 1226 583 1230
rect 595 1211 599 1215
rect 235 1203 239 1207
rect 287 1203 291 1207
rect 375 1203 379 1207
rect 463 1203 467 1207
rect 551 1203 555 1207
rect 683 1203 687 1207
rect 735 1203 739 1207
rect 839 1203 843 1207
rect 1027 1203 1031 1207
rect 1071 1203 1075 1207
rect 219 1186 223 1190
rect 307 1186 311 1190
rect 395 1186 399 1190
rect 483 1186 487 1190
rect 571 1186 575 1190
rect 667 1186 671 1190
rect 771 1186 775 1190
rect 883 1186 887 1190
rect 1003 1186 1007 1190
rect 1099 1186 1103 1190
rect 111 1181 115 1185
rect 1183 1181 1187 1185
rect 111 1163 115 1167
rect 1183 1163 1187 1167
rect 287 1155 291 1159
rect 375 1155 379 1159
rect 463 1155 467 1159
rect 551 1155 555 1159
rect 591 1155 595 1159
rect 735 1155 739 1159
rect 839 1155 843 1159
rect 871 1155 875 1159
rect 1071 1155 1075 1159
rect 215 1145 219 1149
rect 303 1145 307 1149
rect 391 1145 395 1149
rect 479 1145 483 1149
rect 567 1145 571 1149
rect 663 1145 667 1149
rect 767 1145 771 1149
rect 879 1145 883 1149
rect 999 1145 1003 1149
rect 1095 1145 1099 1149
rect 215 1107 219 1111
rect 359 1107 363 1111
rect 503 1107 507 1111
rect 647 1107 651 1111
rect 799 1107 803 1111
rect 951 1107 955 1111
rect 1095 1107 1099 1111
rect 235 1095 239 1099
rect 439 1099 443 1103
rect 723 1099 727 1103
rect 1027 1099 1031 1103
rect 111 1089 115 1093
rect 1183 1089 1187 1093
rect 111 1071 115 1075
rect 431 1071 435 1075
rect 219 1066 223 1070
rect 363 1066 367 1070
rect 507 1066 511 1070
rect 1027 1071 1031 1075
rect 651 1066 655 1070
rect 803 1066 807 1070
rect 1183 1071 1187 1075
rect 955 1066 959 1070
rect 1099 1066 1103 1070
rect 311 1051 315 1055
rect 439 1051 443 1055
rect 871 1051 875 1055
rect 1027 1051 1031 1055
rect 1115 1051 1119 1055
rect 431 1043 435 1047
rect 327 1035 331 1039
rect 723 1035 727 1039
rect 819 1035 823 1039
rect 1059 1035 1063 1039
rect 243 1018 247 1022
rect 111 1013 115 1017
rect 327 1015 331 1019
rect 395 1018 399 1022
rect 547 1018 551 1022
rect 707 1018 711 1022
rect 875 1018 879 1022
rect 1043 1018 1047 1022
rect 1183 1013 1187 1017
rect 111 995 115 999
rect 1183 995 1187 999
rect 311 987 315 991
rect 819 987 823 991
rect 835 987 839 991
rect 1115 987 1119 991
rect 239 977 243 981
rect 391 977 395 981
rect 543 977 547 981
rect 703 977 707 981
rect 871 977 875 981
rect 1039 977 1043 981
rect 327 947 331 951
rect 439 947 443 951
rect 559 947 563 951
rect 687 947 691 951
rect 815 947 819 951
rect 951 947 955 951
rect 1087 947 1091 951
rect 931 939 935 943
rect 1059 939 1063 943
rect 111 929 115 933
rect 1183 929 1187 933
rect 111 911 115 915
rect 331 906 335 910
rect 631 911 635 915
rect 443 906 447 910
rect 563 906 567 910
rect 691 906 695 910
rect 819 906 823 910
rect 1183 911 1187 915
rect 955 906 959 910
rect 1091 906 1095 910
rect 631 891 635 895
rect 731 891 735 895
rect 835 891 839 895
rect 1071 891 1075 895
rect 383 875 387 879
rect 475 875 479 879
rect 583 875 587 879
rect 931 875 935 879
rect 403 858 407 862
rect 515 858 519 862
rect 643 858 647 862
rect 111 853 115 857
rect 731 855 735 859
rect 779 858 783 862
rect 915 858 919 862
rect 1059 858 1063 862
rect 1183 853 1187 857
rect 111 835 115 839
rect 1183 835 1187 839
rect 475 827 479 831
rect 583 827 587 831
rect 903 827 907 831
rect 1071 827 1075 831
rect 399 817 403 821
rect 511 817 515 821
rect 639 817 643 821
rect 775 817 779 821
rect 911 817 915 821
rect 1055 817 1059 821
rect 375 795 379 799
rect 519 795 523 799
rect 663 795 667 799
rect 815 795 819 799
rect 967 795 971 799
rect 1095 795 1099 799
rect 383 783 387 787
rect 923 787 927 791
rect 111 777 115 781
rect 1183 777 1187 781
rect 111 759 115 763
rect 451 759 455 763
rect 595 759 599 763
rect 1039 759 1043 763
rect 379 754 383 758
rect 523 754 527 758
rect 667 754 671 758
rect 819 754 823 758
rect 1183 759 1187 763
rect 971 754 975 758
rect 1099 754 1103 758
rect 451 739 455 743
rect 595 739 599 743
rect 683 739 687 743
rect 903 739 907 743
rect 1039 739 1043 743
rect 1115 739 1119 743
rect 163 727 167 731
rect 215 727 219 731
rect 359 727 363 731
rect 923 727 927 731
rect 1107 727 1111 731
rect 147 710 151 714
rect 267 710 271 714
rect 411 710 415 714
rect 563 710 567 714
rect 111 705 115 709
rect 683 707 687 711
rect 731 710 735 714
rect 907 710 911 714
rect 1091 710 1095 714
rect 1183 705 1187 709
rect 111 687 115 691
rect 1183 687 1187 691
rect 215 679 219 683
rect 359 679 363 683
rect 923 679 927 683
rect 1111 679 1115 683
rect 143 669 147 673
rect 263 669 267 673
rect 407 669 411 673
rect 559 669 563 673
rect 727 669 731 673
rect 903 669 907 673
rect 1087 669 1091 673
rect 143 639 147 643
rect 247 639 251 643
rect 391 639 395 643
rect 551 639 555 643
rect 719 639 723 643
rect 903 639 907 643
rect 1087 639 1091 643
rect 163 627 167 631
rect 915 627 919 631
rect 1103 627 1107 631
rect 111 621 115 625
rect 1183 621 1187 625
rect 111 603 115 607
rect 215 603 219 607
rect 331 603 335 607
rect 623 603 627 607
rect 147 598 151 602
rect 251 598 255 602
rect 395 598 399 602
rect 1183 603 1187 607
rect 555 598 559 602
rect 723 598 727 602
rect 907 598 911 602
rect 1091 598 1095 602
rect 215 583 219 587
rect 331 583 335 587
rect 411 583 415 587
rect 571 583 575 587
rect 923 583 927 587
rect 1099 583 1103 587
rect 283 571 287 575
rect 355 571 359 575
rect 459 571 463 575
rect 707 571 711 575
rect 823 571 827 575
rect 915 571 919 575
rect 1079 571 1083 575
rect 267 554 271 558
rect 379 554 383 558
rect 499 554 503 558
rect 111 549 115 553
rect 579 551 583 555
rect 635 554 639 558
rect 707 551 711 555
rect 779 554 783 558
rect 931 554 935 558
rect 1091 554 1095 558
rect 1183 549 1187 553
rect 111 531 115 535
rect 1183 531 1187 535
rect 355 523 359 527
rect 459 523 463 527
rect 571 523 575 527
rect 939 523 943 527
rect 1099 523 1103 527
rect 263 513 267 517
rect 375 513 379 517
rect 495 513 499 517
rect 631 513 635 517
rect 775 513 779 517
rect 927 513 931 517
rect 1087 513 1091 517
rect 807 495 811 499
rect 911 495 915 499
rect 463 483 467 487
rect 551 483 555 487
rect 639 483 643 487
rect 735 483 739 487
rect 831 483 835 487
rect 919 483 923 487
rect 1007 483 1011 487
rect 1095 483 1099 487
rect 535 471 539 475
rect 623 471 627 475
rect 823 475 827 479
rect 911 475 915 479
rect 1079 471 1083 475
rect 111 465 115 469
rect 1183 465 1187 469
rect 111 447 115 451
rect 1079 447 1083 451
rect 467 442 471 446
rect 555 442 559 446
rect 643 442 647 446
rect 739 442 743 446
rect 835 442 839 446
rect 923 442 927 446
rect 1183 447 1187 451
rect 1011 442 1015 446
rect 1099 442 1103 446
rect 535 427 539 431
rect 623 427 627 431
rect 939 427 943 431
rect 1079 427 1083 431
rect 1107 427 1111 431
rect 455 415 459 419
rect 623 419 627 423
rect 807 415 811 419
rect 815 415 819 419
rect 939 415 943 419
rect 991 415 995 419
rect 1079 415 1083 419
rect 463 407 467 411
rect 551 407 555 411
rect 639 407 643 411
rect 395 398 399 402
rect 483 398 487 402
rect 571 398 575 402
rect 659 398 663 402
rect 747 398 751 402
rect 835 398 839 402
rect 923 398 927 402
rect 1011 398 1015 402
rect 1099 398 1103 402
rect 111 393 115 397
rect 1183 393 1187 397
rect 623 383 627 387
rect 111 375 115 379
rect 1183 375 1187 379
rect 463 367 467 371
rect 551 367 555 371
rect 639 367 643 371
rect 815 367 819 371
rect 903 367 907 371
rect 991 367 995 371
rect 1079 367 1083 371
rect 1107 367 1111 371
rect 391 357 395 361
rect 479 357 483 361
rect 567 357 571 361
rect 655 357 659 361
rect 743 357 747 361
rect 831 357 835 361
rect 919 357 923 361
rect 1007 357 1011 361
rect 1095 357 1099 361
rect 367 335 371 339
rect 479 335 483 339
rect 599 335 603 339
rect 727 335 731 339
rect 863 335 867 339
rect 1007 335 1011 339
rect 855 327 859 331
rect 939 327 943 331
rect 111 317 115 321
rect 1183 317 1187 321
rect 111 299 115 303
rect 1183 299 1187 303
rect 371 294 375 298
rect 483 294 487 298
rect 603 294 607 298
rect 731 294 735 298
rect 867 294 871 298
rect 1011 294 1015 298
rect 903 279 907 283
rect 219 259 223 263
rect 271 259 275 263
rect 359 259 363 263
rect 447 259 451 263
rect 535 259 539 263
rect 203 242 207 246
rect 291 242 295 246
rect 379 242 383 246
rect 467 242 471 246
rect 111 237 115 241
rect 555 242 559 246
rect 1183 237 1187 241
rect 111 219 115 223
rect 1183 219 1187 223
rect 271 211 275 215
rect 359 211 363 215
rect 447 211 451 215
rect 535 211 539 215
rect 199 201 203 205
rect 287 201 291 205
rect 375 201 379 205
rect 463 201 467 205
rect 551 201 555 205
rect 219 187 223 191
rect 751 187 755 191
rect 143 151 147 155
rect 231 151 235 155
rect 319 151 323 155
rect 407 151 411 155
rect 495 151 499 155
rect 583 151 587 155
rect 671 151 675 155
rect 759 151 763 155
rect 391 139 395 143
rect 479 139 483 143
rect 567 139 571 143
rect 655 139 659 143
rect 743 139 747 143
rect 751 143 755 147
rect 111 133 115 137
rect 1183 133 1187 137
rect 111 115 115 119
rect 1183 115 1187 119
rect 147 110 151 114
rect 235 110 239 114
rect 323 110 327 114
rect 411 110 415 114
rect 499 110 503 114
rect 587 110 591 114
rect 675 110 679 114
rect 763 110 767 114
rect 391 95 395 99
rect 479 95 483 99
rect 567 95 571 99
rect 655 95 659 99
rect 743 95 747 99
<< m3 >>
rect 111 1282 115 1283
rect 111 1277 115 1278
rect 575 1282 579 1283
rect 575 1277 579 1278
rect 1183 1282 1187 1283
rect 1183 1277 1187 1278
rect 112 1254 114 1277
rect 576 1272 578 1277
rect 574 1271 580 1272
rect 574 1267 575 1271
rect 579 1267 580 1271
rect 574 1266 580 1267
rect 682 1263 688 1264
rect 682 1259 683 1263
rect 687 1259 688 1263
rect 682 1258 688 1259
rect 110 1253 116 1254
rect 110 1249 111 1253
rect 115 1249 116 1253
rect 110 1248 116 1249
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 578 1230 584 1231
rect 112 1211 114 1230
rect 578 1226 579 1230
rect 583 1226 584 1230
rect 578 1225 584 1226
rect 580 1211 582 1225
rect 594 1215 600 1216
rect 594 1211 595 1215
rect 599 1211 600 1215
rect 111 1210 115 1211
rect 111 1205 115 1206
rect 219 1210 223 1211
rect 307 1210 311 1211
rect 219 1205 223 1206
rect 234 1207 240 1208
rect 112 1186 114 1205
rect 220 1191 222 1205
rect 234 1203 235 1207
rect 239 1203 240 1207
rect 234 1202 240 1203
rect 286 1207 292 1208
rect 286 1203 287 1207
rect 291 1203 292 1207
rect 395 1210 399 1211
rect 307 1205 311 1206
rect 374 1207 380 1208
rect 286 1202 292 1203
rect 218 1190 224 1191
rect 218 1186 219 1190
rect 223 1186 224 1190
rect 110 1185 116 1186
rect 218 1185 224 1186
rect 110 1181 111 1185
rect 115 1181 116 1185
rect 110 1180 116 1181
rect 110 1167 116 1168
rect 110 1163 111 1167
rect 115 1163 116 1167
rect 110 1162 116 1163
rect 112 1123 114 1162
rect 214 1149 220 1150
rect 214 1145 215 1149
rect 219 1145 220 1149
rect 214 1144 220 1145
rect 216 1123 218 1144
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 215 1122 219 1123
rect 215 1117 219 1118
rect 112 1094 114 1117
rect 216 1112 218 1117
rect 214 1111 220 1112
rect 214 1107 215 1111
rect 219 1107 220 1111
rect 214 1106 220 1107
rect 236 1100 238 1202
rect 288 1160 290 1202
rect 308 1191 310 1205
rect 374 1203 375 1207
rect 379 1203 380 1207
rect 483 1210 487 1211
rect 395 1205 399 1206
rect 462 1207 468 1208
rect 374 1202 380 1203
rect 306 1190 312 1191
rect 306 1186 307 1190
rect 311 1186 312 1190
rect 306 1185 312 1186
rect 376 1160 378 1202
rect 396 1191 398 1205
rect 462 1203 463 1207
rect 467 1203 468 1207
rect 571 1210 575 1211
rect 483 1205 487 1206
rect 550 1207 556 1208
rect 462 1202 468 1203
rect 394 1190 400 1191
rect 394 1186 395 1190
rect 399 1186 400 1190
rect 394 1185 400 1186
rect 464 1160 466 1202
rect 484 1191 486 1205
rect 550 1203 551 1207
rect 555 1203 556 1207
rect 571 1205 575 1206
rect 579 1210 583 1211
rect 594 1210 600 1211
rect 667 1210 671 1211
rect 579 1205 583 1206
rect 550 1202 556 1203
rect 482 1190 488 1191
rect 482 1186 483 1190
rect 487 1186 488 1190
rect 482 1185 488 1186
rect 552 1160 554 1202
rect 572 1191 574 1205
rect 570 1190 576 1191
rect 570 1186 571 1190
rect 575 1186 576 1190
rect 596 1187 598 1210
rect 684 1208 686 1258
rect 1184 1254 1186 1277
rect 1182 1253 1188 1254
rect 1182 1249 1183 1253
rect 1187 1249 1188 1253
rect 1182 1248 1188 1249
rect 1182 1235 1188 1236
rect 1182 1231 1183 1235
rect 1187 1231 1188 1235
rect 1182 1230 1188 1231
rect 1184 1211 1186 1230
rect 771 1210 775 1211
rect 667 1205 671 1206
rect 682 1207 688 1208
rect 668 1191 670 1205
rect 682 1203 683 1207
rect 687 1203 688 1207
rect 682 1202 688 1203
rect 734 1207 740 1208
rect 734 1203 735 1207
rect 739 1203 740 1207
rect 883 1210 887 1211
rect 771 1205 775 1206
rect 838 1207 844 1208
rect 734 1202 740 1203
rect 570 1185 576 1186
rect 592 1185 598 1187
rect 666 1190 672 1191
rect 666 1186 667 1190
rect 671 1186 672 1190
rect 666 1185 672 1186
rect 592 1160 594 1185
rect 736 1160 738 1202
rect 772 1191 774 1205
rect 838 1203 839 1207
rect 843 1203 844 1207
rect 883 1205 887 1206
rect 1003 1210 1007 1211
rect 1099 1210 1103 1211
rect 1003 1205 1007 1206
rect 1026 1207 1032 1208
rect 838 1202 844 1203
rect 770 1190 776 1191
rect 770 1186 771 1190
rect 775 1186 776 1190
rect 770 1185 776 1186
rect 840 1160 842 1202
rect 884 1191 886 1205
rect 1004 1191 1006 1205
rect 1026 1203 1027 1207
rect 1031 1203 1032 1207
rect 1026 1202 1032 1203
rect 1070 1207 1076 1208
rect 1070 1203 1071 1207
rect 1075 1203 1076 1207
rect 1099 1205 1103 1206
rect 1183 1210 1187 1211
rect 1183 1205 1187 1206
rect 1070 1202 1076 1203
rect 882 1190 888 1191
rect 882 1186 883 1190
rect 887 1186 888 1190
rect 882 1185 888 1186
rect 1002 1190 1008 1191
rect 1002 1186 1003 1190
rect 1007 1186 1008 1190
rect 1002 1185 1008 1186
rect 286 1159 292 1160
rect 286 1155 287 1159
rect 291 1155 292 1159
rect 286 1154 292 1155
rect 374 1159 380 1160
rect 374 1155 375 1159
rect 379 1155 380 1159
rect 374 1154 380 1155
rect 462 1159 468 1160
rect 462 1155 463 1159
rect 467 1155 468 1159
rect 462 1154 468 1155
rect 550 1159 556 1160
rect 550 1155 551 1159
rect 555 1155 556 1159
rect 550 1154 556 1155
rect 590 1159 596 1160
rect 590 1155 591 1159
rect 595 1155 596 1159
rect 590 1154 596 1155
rect 734 1159 740 1160
rect 734 1155 735 1159
rect 739 1155 740 1159
rect 734 1154 740 1155
rect 838 1159 844 1160
rect 838 1155 839 1159
rect 843 1155 844 1159
rect 838 1154 844 1155
rect 870 1159 876 1160
rect 870 1155 871 1159
rect 875 1155 876 1159
rect 870 1154 876 1155
rect 302 1149 308 1150
rect 302 1145 303 1149
rect 307 1145 308 1149
rect 302 1144 308 1145
rect 390 1149 396 1150
rect 390 1145 391 1149
rect 395 1145 396 1149
rect 390 1144 396 1145
rect 478 1149 484 1150
rect 478 1145 479 1149
rect 483 1145 484 1149
rect 478 1144 484 1145
rect 566 1149 572 1150
rect 566 1145 567 1149
rect 571 1145 572 1149
rect 566 1144 572 1145
rect 662 1149 668 1150
rect 662 1145 663 1149
rect 667 1145 668 1149
rect 662 1144 668 1145
rect 766 1149 772 1150
rect 766 1145 767 1149
rect 771 1145 772 1149
rect 766 1144 772 1145
rect 304 1123 306 1144
rect 392 1123 394 1144
rect 480 1123 482 1144
rect 568 1123 570 1144
rect 664 1123 666 1144
rect 768 1123 770 1144
rect 303 1122 307 1123
rect 303 1117 307 1118
rect 359 1122 363 1123
rect 359 1117 363 1118
rect 391 1122 395 1123
rect 391 1117 395 1118
rect 479 1122 483 1123
rect 479 1117 483 1118
rect 503 1122 507 1123
rect 503 1117 507 1118
rect 567 1122 571 1123
rect 567 1117 571 1118
rect 647 1122 651 1123
rect 647 1117 651 1118
rect 663 1122 667 1123
rect 663 1117 667 1118
rect 767 1122 771 1123
rect 767 1117 771 1118
rect 799 1122 803 1123
rect 799 1117 803 1118
rect 360 1112 362 1117
rect 504 1112 506 1117
rect 648 1112 650 1117
rect 800 1112 802 1117
rect 358 1111 364 1112
rect 358 1107 359 1111
rect 363 1107 364 1111
rect 358 1106 364 1107
rect 502 1111 508 1112
rect 502 1107 503 1111
rect 507 1107 508 1111
rect 502 1106 508 1107
rect 646 1111 652 1112
rect 646 1107 647 1111
rect 651 1107 652 1111
rect 646 1106 652 1107
rect 798 1111 804 1112
rect 798 1107 799 1111
rect 803 1107 804 1111
rect 798 1106 804 1107
rect 438 1103 444 1104
rect 234 1099 240 1100
rect 234 1095 235 1099
rect 239 1095 240 1099
rect 438 1099 439 1103
rect 443 1099 444 1103
rect 438 1098 444 1099
rect 722 1103 728 1104
rect 722 1099 723 1103
rect 727 1099 728 1103
rect 722 1098 728 1099
rect 234 1094 240 1095
rect 110 1093 116 1094
rect 110 1089 111 1093
rect 115 1089 116 1093
rect 110 1088 116 1089
rect 110 1075 116 1076
rect 110 1071 111 1075
rect 115 1071 116 1075
rect 430 1075 436 1076
rect 430 1071 431 1075
rect 435 1071 436 1075
rect 110 1070 116 1071
rect 218 1070 224 1071
rect 112 1043 114 1070
rect 218 1066 219 1070
rect 223 1066 224 1070
rect 218 1065 224 1066
rect 362 1070 368 1071
rect 430 1070 436 1071
rect 362 1066 363 1070
rect 367 1066 368 1070
rect 362 1065 368 1066
rect 220 1043 222 1065
rect 310 1055 316 1056
rect 310 1051 311 1055
rect 315 1051 316 1055
rect 310 1050 316 1051
rect 111 1042 115 1043
rect 111 1037 115 1038
rect 219 1042 223 1043
rect 219 1037 223 1038
rect 243 1042 247 1043
rect 243 1037 247 1038
rect 112 1018 114 1037
rect 244 1023 246 1037
rect 242 1022 248 1023
rect 242 1018 243 1022
rect 247 1018 248 1022
rect 110 1017 116 1018
rect 242 1017 248 1018
rect 110 1013 111 1017
rect 115 1013 116 1017
rect 110 1012 116 1013
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 110 994 116 995
rect 112 963 114 994
rect 312 992 314 1050
rect 364 1043 366 1065
rect 432 1048 434 1070
rect 440 1056 442 1098
rect 506 1070 512 1071
rect 506 1066 507 1070
rect 511 1066 512 1070
rect 506 1065 512 1066
rect 650 1070 656 1071
rect 650 1066 651 1070
rect 655 1066 656 1070
rect 650 1065 656 1066
rect 438 1055 444 1056
rect 438 1051 439 1055
rect 443 1051 444 1055
rect 438 1050 444 1051
rect 430 1047 436 1048
rect 430 1043 431 1047
rect 435 1043 436 1047
rect 508 1043 510 1065
rect 652 1043 654 1065
rect 363 1042 367 1043
rect 326 1039 332 1040
rect 326 1035 327 1039
rect 331 1035 332 1039
rect 363 1037 367 1038
rect 395 1042 399 1043
rect 430 1042 436 1043
rect 507 1042 511 1043
rect 395 1037 399 1038
rect 507 1037 511 1038
rect 547 1042 551 1043
rect 547 1037 551 1038
rect 651 1042 655 1043
rect 651 1037 655 1038
rect 707 1042 711 1043
rect 724 1040 726 1098
rect 802 1070 808 1071
rect 802 1066 803 1070
rect 807 1066 808 1070
rect 802 1065 808 1066
rect 804 1043 806 1065
rect 872 1056 874 1154
rect 878 1149 884 1150
rect 878 1145 879 1149
rect 883 1145 884 1149
rect 878 1144 884 1145
rect 998 1149 1004 1150
rect 998 1145 999 1149
rect 1003 1145 1004 1149
rect 998 1144 1004 1145
rect 880 1123 882 1144
rect 1000 1123 1002 1144
rect 879 1122 883 1123
rect 879 1117 883 1118
rect 951 1122 955 1123
rect 951 1117 955 1118
rect 999 1122 1003 1123
rect 999 1117 1003 1118
rect 952 1112 954 1117
rect 950 1111 956 1112
rect 950 1107 951 1111
rect 955 1107 956 1111
rect 950 1106 956 1107
rect 1028 1104 1030 1202
rect 1072 1160 1074 1202
rect 1100 1191 1102 1205
rect 1098 1190 1104 1191
rect 1098 1186 1099 1190
rect 1103 1186 1104 1190
rect 1184 1186 1186 1205
rect 1098 1185 1104 1186
rect 1182 1185 1188 1186
rect 1182 1181 1183 1185
rect 1187 1181 1188 1185
rect 1182 1180 1188 1181
rect 1182 1167 1188 1168
rect 1182 1163 1183 1167
rect 1187 1163 1188 1167
rect 1182 1162 1188 1163
rect 1070 1159 1076 1160
rect 1070 1155 1071 1159
rect 1075 1155 1076 1159
rect 1070 1154 1076 1155
rect 1094 1149 1100 1150
rect 1094 1145 1095 1149
rect 1099 1145 1100 1149
rect 1094 1144 1100 1145
rect 1096 1123 1098 1144
rect 1184 1123 1186 1162
rect 1095 1122 1099 1123
rect 1095 1117 1099 1118
rect 1183 1122 1187 1123
rect 1183 1117 1187 1118
rect 1096 1112 1098 1117
rect 1094 1111 1100 1112
rect 1094 1107 1095 1111
rect 1099 1107 1100 1111
rect 1094 1106 1100 1107
rect 1026 1103 1032 1104
rect 1026 1099 1027 1103
rect 1031 1099 1032 1103
rect 1026 1098 1032 1099
rect 1184 1094 1186 1117
rect 1182 1093 1188 1094
rect 1182 1089 1183 1093
rect 1187 1089 1188 1093
rect 1182 1088 1188 1089
rect 1026 1075 1032 1076
rect 1026 1071 1027 1075
rect 1031 1071 1032 1075
rect 1182 1075 1188 1076
rect 1182 1071 1183 1075
rect 1187 1071 1188 1075
rect 954 1070 960 1071
rect 1026 1070 1032 1071
rect 1098 1070 1104 1071
rect 1182 1070 1188 1071
rect 954 1066 955 1070
rect 959 1066 960 1070
rect 954 1065 960 1066
rect 870 1055 876 1056
rect 870 1051 871 1055
rect 875 1051 876 1055
rect 870 1050 876 1051
rect 956 1043 958 1065
rect 1028 1056 1030 1070
rect 1098 1066 1099 1070
rect 1103 1066 1104 1070
rect 1098 1065 1104 1066
rect 1026 1055 1032 1056
rect 1026 1051 1027 1055
rect 1031 1051 1032 1055
rect 1026 1050 1032 1051
rect 1100 1043 1102 1065
rect 1114 1055 1120 1056
rect 1114 1051 1115 1055
rect 1119 1051 1120 1055
rect 1114 1050 1120 1051
rect 803 1042 807 1043
rect 707 1037 711 1038
rect 722 1039 728 1040
rect 326 1034 332 1035
rect 328 1020 330 1034
rect 396 1023 398 1037
rect 548 1023 550 1037
rect 708 1023 710 1037
rect 722 1035 723 1039
rect 727 1035 728 1039
rect 875 1042 879 1043
rect 803 1037 807 1038
rect 818 1039 824 1040
rect 722 1034 728 1035
rect 818 1035 819 1039
rect 823 1035 824 1039
rect 875 1037 879 1038
rect 955 1042 959 1043
rect 955 1037 959 1038
rect 1043 1042 1047 1043
rect 1099 1042 1103 1043
rect 1043 1037 1047 1038
rect 1058 1039 1064 1040
rect 818 1034 824 1035
rect 394 1022 400 1023
rect 326 1019 332 1020
rect 326 1015 327 1019
rect 331 1015 332 1019
rect 394 1018 395 1022
rect 399 1018 400 1022
rect 394 1017 400 1018
rect 546 1022 552 1023
rect 546 1018 547 1022
rect 551 1018 552 1022
rect 546 1017 552 1018
rect 706 1022 712 1023
rect 706 1018 707 1022
rect 711 1018 712 1022
rect 706 1017 712 1018
rect 326 1014 332 1015
rect 820 992 822 1034
rect 876 1023 878 1037
rect 1044 1023 1046 1037
rect 1058 1035 1059 1039
rect 1063 1035 1064 1039
rect 1099 1037 1103 1038
rect 1058 1034 1064 1035
rect 874 1022 880 1023
rect 874 1018 875 1022
rect 879 1018 880 1022
rect 874 1017 880 1018
rect 1042 1022 1048 1023
rect 1042 1018 1043 1022
rect 1047 1018 1048 1022
rect 1042 1017 1048 1018
rect 310 991 316 992
rect 310 987 311 991
rect 315 987 316 991
rect 310 986 316 987
rect 818 991 824 992
rect 818 987 819 991
rect 823 987 824 991
rect 818 986 824 987
rect 834 991 840 992
rect 834 987 835 991
rect 839 987 840 991
rect 834 986 840 987
rect 238 981 244 982
rect 238 977 239 981
rect 243 977 244 981
rect 238 976 244 977
rect 390 981 396 982
rect 390 977 391 981
rect 395 977 396 981
rect 390 976 396 977
rect 542 981 548 982
rect 542 977 543 981
rect 547 977 548 981
rect 542 976 548 977
rect 702 981 708 982
rect 702 977 703 981
rect 707 977 708 981
rect 702 976 708 977
rect 240 963 242 976
rect 392 963 394 976
rect 544 963 546 976
rect 704 963 706 976
rect 111 962 115 963
rect 111 957 115 958
rect 239 962 243 963
rect 239 957 243 958
rect 327 962 331 963
rect 327 957 331 958
rect 391 962 395 963
rect 391 957 395 958
rect 439 962 443 963
rect 439 957 443 958
rect 543 962 547 963
rect 543 957 547 958
rect 559 962 563 963
rect 559 957 563 958
rect 687 962 691 963
rect 687 957 691 958
rect 703 962 707 963
rect 703 957 707 958
rect 815 962 819 963
rect 815 957 819 958
rect 112 934 114 957
rect 328 952 330 957
rect 440 952 442 957
rect 560 952 562 957
rect 688 952 690 957
rect 816 952 818 957
rect 326 951 332 952
rect 326 947 327 951
rect 331 947 332 951
rect 326 946 332 947
rect 438 951 444 952
rect 438 947 439 951
rect 443 947 444 951
rect 438 946 444 947
rect 558 951 564 952
rect 558 947 559 951
rect 563 947 564 951
rect 558 946 564 947
rect 686 951 692 952
rect 686 947 687 951
rect 691 947 692 951
rect 686 946 692 947
rect 814 951 820 952
rect 814 947 815 951
rect 819 947 820 951
rect 814 946 820 947
rect 110 933 116 934
rect 110 929 111 933
rect 115 929 116 933
rect 110 928 116 929
rect 110 915 116 916
rect 110 911 111 915
rect 115 911 116 915
rect 630 915 636 916
rect 630 911 631 915
rect 635 911 636 915
rect 110 910 116 911
rect 330 910 336 911
rect 112 883 114 910
rect 330 906 331 910
rect 335 906 336 910
rect 330 905 336 906
rect 442 910 448 911
rect 442 906 443 910
rect 447 906 448 910
rect 442 905 448 906
rect 562 910 568 911
rect 630 910 636 911
rect 690 910 696 911
rect 562 906 563 910
rect 567 906 568 910
rect 562 905 568 906
rect 332 883 334 905
rect 444 883 446 905
rect 564 883 566 905
rect 632 896 634 910
rect 690 906 691 910
rect 695 906 696 910
rect 690 905 696 906
rect 818 910 824 911
rect 818 906 819 910
rect 823 906 824 910
rect 818 905 824 906
rect 630 895 636 896
rect 630 891 631 895
rect 635 891 636 895
rect 630 890 636 891
rect 692 883 694 905
rect 730 895 736 896
rect 730 891 731 895
rect 735 891 736 895
rect 730 890 736 891
rect 111 882 115 883
rect 111 877 115 878
rect 331 882 335 883
rect 403 882 407 883
rect 331 877 335 878
rect 382 879 388 880
rect 112 858 114 877
rect 382 875 383 879
rect 387 875 388 879
rect 403 877 407 878
rect 443 882 447 883
rect 515 882 519 883
rect 443 877 447 878
rect 474 879 480 880
rect 382 874 388 875
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 110 852 116 853
rect 110 839 116 840
rect 110 835 111 839
rect 115 835 116 839
rect 110 834 116 835
rect 112 811 114 834
rect 111 810 115 811
rect 111 805 115 806
rect 375 810 379 811
rect 375 805 379 806
rect 112 782 114 805
rect 376 800 378 805
rect 374 799 380 800
rect 374 795 375 799
rect 379 795 380 799
rect 374 794 380 795
rect 384 788 386 874
rect 404 863 406 877
rect 474 875 475 879
rect 479 875 480 879
rect 515 877 519 878
rect 563 882 567 883
rect 643 882 647 883
rect 563 877 567 878
rect 582 879 588 880
rect 474 874 480 875
rect 402 862 408 863
rect 402 858 403 862
rect 407 858 408 862
rect 402 857 408 858
rect 476 832 478 874
rect 516 863 518 877
rect 582 875 583 879
rect 587 875 588 879
rect 643 877 647 878
rect 691 882 695 883
rect 691 877 695 878
rect 582 874 588 875
rect 514 862 520 863
rect 514 858 515 862
rect 519 858 520 862
rect 514 857 520 858
rect 584 832 586 874
rect 644 863 646 877
rect 642 862 648 863
rect 642 858 643 862
rect 647 858 648 862
rect 732 860 734 890
rect 820 883 822 905
rect 836 896 838 986
rect 870 981 876 982
rect 870 977 871 981
rect 875 977 876 981
rect 870 976 876 977
rect 1038 981 1044 982
rect 1038 977 1039 981
rect 1043 977 1044 981
rect 1038 976 1044 977
rect 872 963 874 976
rect 1040 963 1042 976
rect 871 962 875 963
rect 871 957 875 958
rect 951 962 955 963
rect 951 957 955 958
rect 1039 962 1043 963
rect 1039 957 1043 958
rect 952 952 954 957
rect 950 951 956 952
rect 950 947 951 951
rect 955 947 956 951
rect 950 946 956 947
rect 1060 944 1062 1034
rect 1116 992 1118 1050
rect 1184 1043 1186 1070
rect 1183 1042 1187 1043
rect 1183 1037 1187 1038
rect 1184 1018 1186 1037
rect 1182 1017 1188 1018
rect 1182 1013 1183 1017
rect 1187 1013 1188 1017
rect 1182 1012 1188 1013
rect 1182 999 1188 1000
rect 1182 995 1183 999
rect 1187 995 1188 999
rect 1182 994 1188 995
rect 1114 991 1120 992
rect 1114 987 1115 991
rect 1119 987 1120 991
rect 1114 986 1120 987
rect 1184 963 1186 994
rect 1087 962 1091 963
rect 1087 957 1091 958
rect 1183 962 1187 963
rect 1183 957 1187 958
rect 1088 952 1090 957
rect 1086 951 1092 952
rect 1086 947 1087 951
rect 1091 947 1092 951
rect 1086 946 1092 947
rect 930 943 936 944
rect 930 939 931 943
rect 935 939 936 943
rect 930 938 936 939
rect 1058 943 1064 944
rect 1058 939 1059 943
rect 1063 939 1064 943
rect 1058 938 1064 939
rect 834 895 840 896
rect 834 891 835 895
rect 839 891 840 895
rect 834 890 840 891
rect 779 882 783 883
rect 779 877 783 878
rect 819 882 823 883
rect 819 877 823 878
rect 915 882 919 883
rect 932 880 934 938
rect 1184 934 1186 957
rect 1182 933 1188 934
rect 1182 929 1183 933
rect 1187 929 1188 933
rect 1182 928 1188 929
rect 1182 915 1188 916
rect 1182 911 1183 915
rect 1187 911 1188 915
rect 954 910 960 911
rect 954 906 955 910
rect 959 906 960 910
rect 954 905 960 906
rect 1090 910 1096 911
rect 1182 910 1188 911
rect 1090 906 1091 910
rect 1095 906 1096 910
rect 1090 905 1096 906
rect 956 883 958 905
rect 1070 895 1076 896
rect 1070 891 1071 895
rect 1075 891 1076 895
rect 1070 890 1076 891
rect 955 882 959 883
rect 915 877 919 878
rect 930 879 936 880
rect 780 863 782 877
rect 916 863 918 877
rect 930 875 931 879
rect 935 875 936 879
rect 955 877 959 878
rect 1059 882 1063 883
rect 1059 877 1063 878
rect 930 874 936 875
rect 1060 863 1062 877
rect 778 862 784 863
rect 642 857 648 858
rect 730 859 736 860
rect 730 855 731 859
rect 735 855 736 859
rect 778 858 779 862
rect 783 858 784 862
rect 778 857 784 858
rect 914 862 920 863
rect 914 858 915 862
rect 919 858 920 862
rect 914 857 920 858
rect 1058 862 1064 863
rect 1058 858 1059 862
rect 1063 858 1064 862
rect 1058 857 1064 858
rect 730 854 736 855
rect 1072 832 1074 890
rect 1092 883 1094 905
rect 1184 883 1186 910
rect 1091 882 1095 883
rect 1091 877 1095 878
rect 1183 882 1187 883
rect 1183 877 1187 878
rect 1184 858 1186 877
rect 1182 857 1188 858
rect 1182 853 1183 857
rect 1187 853 1188 857
rect 1182 852 1188 853
rect 1182 839 1188 840
rect 1182 835 1183 839
rect 1187 835 1188 839
rect 1182 834 1188 835
rect 474 831 480 832
rect 474 827 475 831
rect 479 827 480 831
rect 474 826 480 827
rect 582 831 588 832
rect 582 827 583 831
rect 587 827 588 831
rect 582 826 588 827
rect 902 831 908 832
rect 902 827 903 831
rect 907 827 908 831
rect 902 826 908 827
rect 1070 831 1076 832
rect 1070 827 1071 831
rect 1075 827 1076 831
rect 1070 826 1076 827
rect 398 821 404 822
rect 398 817 399 821
rect 403 817 404 821
rect 398 816 404 817
rect 510 821 516 822
rect 510 817 511 821
rect 515 817 516 821
rect 510 816 516 817
rect 638 821 644 822
rect 638 817 639 821
rect 643 817 644 821
rect 638 816 644 817
rect 774 821 780 822
rect 774 817 775 821
rect 779 817 780 821
rect 774 816 780 817
rect 400 811 402 816
rect 512 811 514 816
rect 640 811 642 816
rect 776 811 778 816
rect 399 810 403 811
rect 399 805 403 806
rect 511 810 515 811
rect 511 805 515 806
rect 519 810 523 811
rect 519 805 523 806
rect 639 810 643 811
rect 639 805 643 806
rect 663 810 667 811
rect 663 805 667 806
rect 775 810 779 811
rect 775 805 779 806
rect 815 810 819 811
rect 815 805 819 806
rect 520 800 522 805
rect 664 800 666 805
rect 816 800 818 805
rect 518 799 524 800
rect 518 795 519 799
rect 523 795 524 799
rect 518 794 524 795
rect 662 799 668 800
rect 662 795 663 799
rect 667 795 668 799
rect 662 794 668 795
rect 814 799 820 800
rect 814 795 815 799
rect 819 795 820 799
rect 814 794 820 795
rect 382 787 388 788
rect 382 783 383 787
rect 387 783 388 787
rect 382 782 388 783
rect 110 781 116 782
rect 110 777 111 781
rect 115 777 116 781
rect 110 776 116 777
rect 110 763 116 764
rect 110 759 111 763
rect 115 759 116 763
rect 450 763 456 764
rect 450 759 451 763
rect 455 759 456 763
rect 594 763 600 764
rect 594 759 595 763
rect 599 759 600 763
rect 110 758 116 759
rect 378 758 384 759
rect 450 758 456 759
rect 522 758 528 759
rect 594 758 600 759
rect 666 758 672 759
rect 112 735 114 758
rect 378 754 379 758
rect 383 754 384 758
rect 378 753 384 754
rect 380 735 382 753
rect 452 744 454 758
rect 522 754 523 758
rect 527 754 528 758
rect 522 753 528 754
rect 450 743 456 744
rect 450 739 451 743
rect 455 739 456 743
rect 450 738 456 739
rect 524 735 526 753
rect 596 744 598 758
rect 666 754 667 758
rect 671 754 672 758
rect 666 753 672 754
rect 818 758 824 759
rect 818 754 819 758
rect 823 754 824 758
rect 818 753 824 754
rect 594 743 600 744
rect 594 739 595 743
rect 599 739 600 743
rect 594 738 600 739
rect 668 735 670 753
rect 682 743 688 744
rect 682 739 683 743
rect 687 739 688 743
rect 682 738 688 739
rect 111 734 115 735
rect 111 729 115 730
rect 147 734 151 735
rect 267 734 271 735
rect 147 729 151 730
rect 162 731 168 732
rect 112 710 114 729
rect 148 715 150 729
rect 162 727 163 731
rect 167 727 168 731
rect 162 726 168 727
rect 214 731 220 732
rect 214 727 215 731
rect 219 727 220 731
rect 379 734 383 735
rect 267 729 271 730
rect 358 731 364 732
rect 214 726 220 727
rect 146 714 152 715
rect 146 710 147 714
rect 151 710 152 714
rect 110 709 116 710
rect 146 709 152 710
rect 110 705 111 709
rect 115 705 116 709
rect 110 704 116 705
rect 110 691 116 692
rect 110 687 111 691
rect 115 687 116 691
rect 110 686 116 687
rect 112 655 114 686
rect 142 673 148 674
rect 142 669 143 673
rect 147 669 148 673
rect 142 668 148 669
rect 144 655 146 668
rect 111 654 115 655
rect 111 649 115 650
rect 143 654 147 655
rect 143 649 147 650
rect 112 626 114 649
rect 144 644 146 649
rect 142 643 148 644
rect 142 639 143 643
rect 147 639 148 643
rect 142 638 148 639
rect 164 632 166 726
rect 216 684 218 726
rect 268 715 270 729
rect 358 727 359 731
rect 363 727 364 731
rect 379 729 383 730
rect 411 734 415 735
rect 411 729 415 730
rect 523 734 527 735
rect 523 729 527 730
rect 563 734 567 735
rect 563 729 567 730
rect 667 734 671 735
rect 667 729 671 730
rect 358 726 364 727
rect 266 714 272 715
rect 266 710 267 714
rect 271 710 272 714
rect 266 709 272 710
rect 360 684 362 726
rect 412 715 414 729
rect 564 715 566 729
rect 410 714 416 715
rect 410 710 411 714
rect 415 710 416 714
rect 410 709 416 710
rect 562 714 568 715
rect 562 710 563 714
rect 567 710 568 714
rect 684 712 686 738
rect 820 735 822 753
rect 904 744 906 826
rect 910 821 916 822
rect 910 817 911 821
rect 915 817 916 821
rect 910 816 916 817
rect 1054 821 1060 822
rect 1054 817 1055 821
rect 1059 817 1060 821
rect 1054 816 1060 817
rect 912 811 914 816
rect 1056 811 1058 816
rect 1184 811 1186 834
rect 911 810 915 811
rect 911 805 915 806
rect 967 810 971 811
rect 967 805 971 806
rect 1055 810 1059 811
rect 1055 805 1059 806
rect 1095 810 1099 811
rect 1095 805 1099 806
rect 1183 810 1187 811
rect 1183 805 1187 806
rect 968 800 970 805
rect 1096 800 1098 805
rect 966 799 972 800
rect 966 795 967 799
rect 971 795 972 799
rect 966 794 972 795
rect 1094 799 1100 800
rect 1094 795 1095 799
rect 1099 795 1100 799
rect 1094 794 1100 795
rect 922 791 928 792
rect 922 787 923 791
rect 927 787 928 791
rect 922 786 928 787
rect 902 743 908 744
rect 902 739 903 743
rect 907 739 908 743
rect 902 738 908 739
rect 731 734 735 735
rect 731 729 735 730
rect 819 734 823 735
rect 819 729 823 730
rect 907 734 911 735
rect 924 732 926 786
rect 1184 782 1186 805
rect 1182 781 1188 782
rect 1182 777 1183 781
rect 1187 777 1188 781
rect 1182 776 1188 777
rect 1038 763 1044 764
rect 1038 759 1039 763
rect 1043 759 1044 763
rect 1182 763 1188 764
rect 1182 759 1183 763
rect 1187 759 1188 763
rect 970 758 976 759
rect 1038 758 1044 759
rect 1098 758 1104 759
rect 1182 758 1188 759
rect 970 754 971 758
rect 975 754 976 758
rect 970 753 976 754
rect 972 735 974 753
rect 1040 744 1042 758
rect 1098 754 1099 758
rect 1103 754 1104 758
rect 1098 753 1104 754
rect 1038 743 1044 744
rect 1038 739 1039 743
rect 1043 739 1044 743
rect 1038 738 1044 739
rect 1100 735 1102 753
rect 1114 743 1120 744
rect 1114 739 1115 743
rect 1119 739 1120 743
rect 1114 738 1120 739
rect 971 734 975 735
rect 907 729 911 730
rect 922 731 928 732
rect 732 715 734 729
rect 908 715 910 729
rect 922 727 923 731
rect 927 727 928 731
rect 971 729 975 730
rect 1091 734 1095 735
rect 1091 729 1095 730
rect 1099 734 1103 735
rect 1099 729 1103 730
rect 1106 731 1112 732
rect 922 726 928 727
rect 1092 715 1094 729
rect 1106 727 1107 731
rect 1111 727 1112 731
rect 1106 726 1112 727
rect 730 714 736 715
rect 562 709 568 710
rect 682 711 688 712
rect 682 707 683 711
rect 687 707 688 711
rect 730 710 731 714
rect 735 710 736 714
rect 730 709 736 710
rect 906 714 912 715
rect 906 710 907 714
rect 911 710 912 714
rect 906 709 912 710
rect 1090 714 1096 715
rect 1090 710 1091 714
rect 1095 710 1096 714
rect 1090 709 1096 710
rect 682 706 688 707
rect 1108 691 1110 726
rect 1116 715 1118 738
rect 1184 735 1186 758
rect 1183 734 1187 735
rect 1183 729 1187 730
rect 1104 689 1110 691
rect 1112 713 1118 715
rect 214 683 220 684
rect 214 679 215 683
rect 219 679 220 683
rect 214 678 220 679
rect 358 683 364 684
rect 358 679 359 683
rect 363 679 364 683
rect 358 678 364 679
rect 922 683 928 684
rect 922 679 923 683
rect 927 679 928 683
rect 922 678 928 679
rect 262 673 268 674
rect 262 669 263 673
rect 267 669 268 673
rect 262 668 268 669
rect 406 673 412 674
rect 406 669 407 673
rect 411 669 412 673
rect 406 668 412 669
rect 558 673 564 674
rect 558 669 559 673
rect 563 669 564 673
rect 558 668 564 669
rect 726 673 732 674
rect 726 669 727 673
rect 731 669 732 673
rect 726 668 732 669
rect 902 673 908 674
rect 902 669 903 673
rect 907 669 908 673
rect 902 668 908 669
rect 264 655 266 668
rect 408 655 410 668
rect 560 655 562 668
rect 728 655 730 668
rect 904 655 906 668
rect 247 654 251 655
rect 247 649 251 650
rect 263 654 267 655
rect 263 649 267 650
rect 391 654 395 655
rect 391 649 395 650
rect 407 654 411 655
rect 407 649 411 650
rect 551 654 555 655
rect 551 649 555 650
rect 559 654 563 655
rect 559 649 563 650
rect 719 654 723 655
rect 719 649 723 650
rect 727 654 731 655
rect 727 649 731 650
rect 903 654 907 655
rect 903 649 907 650
rect 248 644 250 649
rect 392 644 394 649
rect 552 644 554 649
rect 720 644 722 649
rect 904 644 906 649
rect 246 643 252 644
rect 246 639 247 643
rect 251 639 252 643
rect 246 638 252 639
rect 390 643 396 644
rect 390 639 391 643
rect 395 639 396 643
rect 390 638 396 639
rect 550 643 556 644
rect 550 639 551 643
rect 555 639 556 643
rect 550 638 556 639
rect 718 643 724 644
rect 718 639 719 643
rect 723 639 724 643
rect 718 638 724 639
rect 902 643 908 644
rect 902 639 903 643
rect 907 639 908 643
rect 902 638 908 639
rect 162 631 168 632
rect 162 627 163 631
rect 167 627 168 631
rect 162 626 168 627
rect 914 631 920 632
rect 914 627 915 631
rect 919 627 920 631
rect 914 626 920 627
rect 110 625 116 626
rect 110 621 111 625
rect 115 621 116 625
rect 110 620 116 621
rect 110 607 116 608
rect 110 603 111 607
rect 115 603 116 607
rect 214 607 220 608
rect 214 603 215 607
rect 219 603 220 607
rect 330 607 336 608
rect 330 603 331 607
rect 335 603 336 607
rect 622 607 628 608
rect 622 603 623 607
rect 627 603 628 607
rect 110 602 116 603
rect 146 602 152 603
rect 214 602 220 603
rect 250 602 256 603
rect 330 602 336 603
rect 394 602 400 603
rect 112 579 114 602
rect 146 598 147 602
rect 151 598 152 602
rect 146 597 152 598
rect 148 579 150 597
rect 216 588 218 602
rect 250 598 251 602
rect 255 598 256 602
rect 250 597 256 598
rect 214 587 220 588
rect 214 583 215 587
rect 219 583 220 587
rect 214 582 220 583
rect 252 579 254 597
rect 332 588 334 602
rect 394 598 395 602
rect 399 598 400 602
rect 394 597 400 598
rect 554 602 560 603
rect 622 602 628 603
rect 722 602 728 603
rect 554 598 555 602
rect 559 598 560 602
rect 554 597 560 598
rect 624 597 626 602
rect 722 598 723 602
rect 727 598 728 602
rect 722 597 728 598
rect 906 602 912 603
rect 906 598 907 602
rect 911 598 912 602
rect 906 597 912 598
rect 330 587 336 588
rect 330 583 331 587
rect 335 583 336 587
rect 330 582 336 583
rect 396 579 398 597
rect 411 596 415 597
rect 411 591 415 592
rect 412 588 414 591
rect 410 587 416 588
rect 410 583 411 587
rect 415 583 416 587
rect 410 582 416 583
rect 556 579 558 597
rect 623 596 627 597
rect 623 591 627 592
rect 570 587 576 588
rect 570 583 571 587
rect 575 583 576 587
rect 570 582 576 583
rect 111 578 115 579
rect 111 573 115 574
rect 147 578 151 579
rect 147 573 151 574
rect 251 578 255 579
rect 251 573 255 574
rect 267 578 271 579
rect 379 578 383 579
rect 267 573 271 574
rect 282 575 288 576
rect 112 554 114 573
rect 268 559 270 573
rect 282 571 283 575
rect 287 571 288 575
rect 282 570 288 571
rect 354 575 360 576
rect 354 571 355 575
rect 359 571 360 575
rect 379 573 383 574
rect 395 578 399 579
rect 499 578 503 579
rect 395 573 399 574
rect 458 575 464 576
rect 354 570 360 571
rect 284 565 286 570
rect 283 564 287 565
rect 283 559 287 560
rect 266 558 272 559
rect 266 554 267 558
rect 271 554 272 558
rect 110 553 116 554
rect 266 553 272 554
rect 110 549 111 553
rect 115 549 116 553
rect 110 548 116 549
rect 110 535 116 536
rect 110 531 111 535
rect 115 531 116 535
rect 110 530 116 531
rect 112 499 114 530
rect 356 528 358 570
rect 380 559 382 573
rect 458 571 459 575
rect 463 571 464 575
rect 499 573 503 574
rect 555 578 559 579
rect 555 573 559 574
rect 458 570 464 571
rect 378 558 384 559
rect 378 554 379 558
rect 383 554 384 558
rect 378 553 384 554
rect 460 528 462 570
rect 500 559 502 573
rect 498 558 504 559
rect 498 554 499 558
rect 503 554 504 558
rect 498 553 504 554
rect 572 528 574 582
rect 724 579 726 597
rect 908 579 910 597
rect 635 578 639 579
rect 723 578 727 579
rect 635 573 639 574
rect 706 575 712 576
rect 579 564 583 565
rect 579 559 583 560
rect 636 559 638 573
rect 706 571 707 575
rect 711 571 712 575
rect 723 573 727 574
rect 779 578 783 579
rect 907 578 911 579
rect 779 573 783 574
rect 822 575 828 576
rect 706 570 712 571
rect 580 556 582 559
rect 634 558 640 559
rect 578 555 584 556
rect 578 551 579 555
rect 583 551 584 555
rect 634 554 635 558
rect 639 554 640 558
rect 708 556 710 570
rect 780 559 782 573
rect 822 571 823 575
rect 827 571 828 575
rect 916 576 918 626
rect 924 588 926 678
rect 1086 673 1092 674
rect 1086 669 1087 673
rect 1091 669 1092 673
rect 1086 668 1092 669
rect 1088 655 1090 668
rect 1087 654 1091 655
rect 1087 649 1091 650
rect 1088 644 1090 649
rect 1086 643 1092 644
rect 1086 639 1087 643
rect 1091 639 1092 643
rect 1086 638 1092 639
rect 1104 632 1106 689
rect 1112 684 1114 713
rect 1184 710 1186 729
rect 1182 709 1188 710
rect 1182 705 1183 709
rect 1187 705 1188 709
rect 1182 704 1188 705
rect 1182 691 1188 692
rect 1182 687 1183 691
rect 1187 687 1188 691
rect 1182 686 1188 687
rect 1110 683 1116 684
rect 1110 679 1111 683
rect 1115 679 1116 683
rect 1110 678 1116 679
rect 1184 655 1186 686
rect 1183 654 1187 655
rect 1183 649 1187 650
rect 1102 631 1108 632
rect 1102 627 1103 631
rect 1107 627 1108 631
rect 1102 626 1108 627
rect 1184 626 1186 649
rect 1182 625 1188 626
rect 1182 621 1183 625
rect 1187 621 1188 625
rect 1182 620 1188 621
rect 1182 607 1188 608
rect 1182 603 1183 607
rect 1187 603 1188 607
rect 1090 602 1096 603
rect 1182 602 1188 603
rect 1090 598 1091 602
rect 1095 598 1096 602
rect 1090 597 1096 598
rect 922 587 928 588
rect 922 583 923 587
rect 927 583 928 587
rect 922 582 928 583
rect 1092 579 1094 597
rect 1098 587 1104 588
rect 1098 583 1099 587
rect 1103 583 1104 587
rect 1098 582 1104 583
rect 931 578 935 579
rect 907 573 911 574
rect 914 575 920 576
rect 822 570 828 571
rect 914 571 915 575
rect 919 571 920 575
rect 1091 578 1095 579
rect 931 573 935 574
rect 1078 575 1084 576
rect 914 570 920 571
rect 778 558 784 559
rect 634 553 640 554
rect 706 555 712 556
rect 578 550 584 551
rect 706 551 707 555
rect 711 551 712 555
rect 778 554 779 558
rect 783 554 784 558
rect 778 553 784 554
rect 706 550 712 551
rect 354 527 360 528
rect 354 523 355 527
rect 359 523 360 527
rect 354 522 360 523
rect 458 527 464 528
rect 458 523 459 527
rect 463 523 464 527
rect 458 522 464 523
rect 570 527 576 528
rect 570 523 571 527
rect 575 523 576 527
rect 570 522 576 523
rect 262 517 268 518
rect 262 513 263 517
rect 267 513 268 517
rect 262 512 268 513
rect 374 517 380 518
rect 374 513 375 517
rect 379 513 380 517
rect 374 512 380 513
rect 494 517 500 518
rect 494 513 495 517
rect 499 513 500 517
rect 494 512 500 513
rect 630 517 636 518
rect 630 513 631 517
rect 635 513 636 517
rect 630 512 636 513
rect 774 517 780 518
rect 774 513 775 517
rect 779 513 780 517
rect 774 512 780 513
rect 264 499 266 512
rect 376 499 378 512
rect 496 499 498 512
rect 632 499 634 512
rect 776 499 778 512
rect 806 499 812 500
rect 111 498 115 499
rect 111 493 115 494
rect 263 498 267 499
rect 263 493 267 494
rect 375 498 379 499
rect 375 493 379 494
rect 463 498 467 499
rect 463 493 467 494
rect 495 498 499 499
rect 495 493 499 494
rect 551 498 555 499
rect 551 493 555 494
rect 631 498 635 499
rect 631 493 635 494
rect 639 498 643 499
rect 639 493 643 494
rect 735 498 739 499
rect 735 493 739 494
rect 775 498 779 499
rect 806 495 807 499
rect 811 495 812 499
rect 806 494 812 495
rect 775 493 779 494
rect 112 470 114 493
rect 464 488 466 493
rect 552 488 554 493
rect 640 488 642 493
rect 736 488 738 493
rect 462 487 468 488
rect 462 483 463 487
rect 467 483 468 487
rect 462 482 468 483
rect 550 487 556 488
rect 550 483 551 487
rect 555 483 556 487
rect 550 482 556 483
rect 638 487 644 488
rect 638 483 639 487
rect 643 483 644 487
rect 638 482 644 483
rect 734 487 740 488
rect 734 483 735 487
rect 739 483 740 487
rect 734 482 740 483
rect 534 475 540 476
rect 534 471 535 475
rect 539 471 540 475
rect 534 470 540 471
rect 622 475 628 476
rect 622 471 623 475
rect 627 471 628 475
rect 622 470 628 471
rect 110 469 116 470
rect 110 465 111 469
rect 115 465 116 469
rect 110 464 116 465
rect 110 451 116 452
rect 110 447 111 451
rect 115 447 116 451
rect 110 446 116 447
rect 466 446 472 447
rect 112 423 114 446
rect 466 442 467 446
rect 471 442 472 446
rect 466 441 472 442
rect 468 423 470 441
rect 536 432 538 470
rect 554 446 560 447
rect 554 442 555 446
rect 559 442 560 446
rect 554 441 560 442
rect 534 431 540 432
rect 534 427 535 431
rect 539 427 540 431
rect 534 426 540 427
rect 556 423 558 441
rect 624 432 626 470
rect 642 446 648 447
rect 642 442 643 446
rect 647 442 648 446
rect 642 441 648 442
rect 738 446 744 447
rect 738 442 739 446
rect 743 442 744 446
rect 738 441 744 442
rect 622 431 628 432
rect 622 427 623 431
rect 627 427 628 431
rect 622 426 628 427
rect 622 423 628 424
rect 644 423 646 441
rect 740 423 742 441
rect 111 422 115 423
rect 111 417 115 418
rect 395 422 399 423
rect 467 422 471 423
rect 395 417 399 418
rect 454 419 460 420
rect 112 398 114 417
rect 396 403 398 417
rect 454 415 455 419
rect 459 415 460 419
rect 467 417 471 418
rect 483 422 487 423
rect 483 417 487 418
rect 555 422 559 423
rect 555 417 559 418
rect 571 422 575 423
rect 622 419 623 423
rect 627 419 628 423
rect 622 418 628 419
rect 643 422 647 423
rect 571 417 575 418
rect 454 414 460 415
rect 394 402 400 403
rect 394 398 395 402
rect 399 398 400 402
rect 110 397 116 398
rect 394 397 400 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 110 379 116 380
rect 110 375 111 379
rect 115 375 116 379
rect 110 374 116 375
rect 112 351 114 374
rect 456 373 458 414
rect 462 411 468 412
rect 462 407 463 411
rect 467 407 468 411
rect 462 406 468 407
rect 455 372 459 373
rect 464 372 466 406
rect 484 403 486 417
rect 550 411 556 412
rect 550 407 551 411
rect 555 407 556 411
rect 550 406 556 407
rect 482 402 488 403
rect 482 398 483 402
rect 487 398 488 402
rect 482 397 488 398
rect 552 372 554 406
rect 572 403 574 417
rect 570 402 576 403
rect 570 398 571 402
rect 575 398 576 402
rect 570 397 576 398
rect 624 388 626 418
rect 643 417 647 418
rect 659 422 663 423
rect 659 417 663 418
rect 739 422 743 423
rect 739 417 743 418
rect 747 422 751 423
rect 808 420 810 494
rect 824 480 826 570
rect 932 559 934 573
rect 1078 571 1079 575
rect 1083 571 1084 575
rect 1091 573 1095 574
rect 1078 570 1084 571
rect 930 558 936 559
rect 930 554 931 558
rect 935 554 936 558
rect 930 553 936 554
rect 938 527 944 528
rect 938 523 939 527
rect 943 523 944 527
rect 938 522 944 523
rect 926 517 932 518
rect 926 513 927 517
rect 931 513 932 517
rect 926 512 932 513
rect 910 499 916 500
rect 928 499 930 512
rect 831 498 835 499
rect 910 495 911 499
rect 915 495 916 499
rect 910 494 916 495
rect 919 498 923 499
rect 831 493 835 494
rect 832 488 834 493
rect 830 487 836 488
rect 830 483 831 487
rect 835 483 836 487
rect 830 482 836 483
rect 912 480 914 494
rect 919 493 923 494
rect 927 498 931 499
rect 927 493 931 494
rect 920 488 922 493
rect 918 487 924 488
rect 918 483 919 487
rect 923 483 924 487
rect 918 482 924 483
rect 822 479 828 480
rect 822 475 823 479
rect 827 475 828 479
rect 822 474 828 475
rect 910 479 916 480
rect 910 475 911 479
rect 915 475 916 479
rect 910 474 916 475
rect 834 446 840 447
rect 834 442 835 446
rect 839 442 840 446
rect 834 441 840 442
rect 922 446 928 447
rect 922 442 923 446
rect 927 442 928 446
rect 922 441 928 442
rect 836 423 838 441
rect 924 423 926 441
rect 940 432 942 522
rect 1007 498 1011 499
rect 1007 493 1011 494
rect 1008 488 1010 493
rect 1006 487 1012 488
rect 1006 483 1007 487
rect 1011 483 1012 487
rect 1006 482 1012 483
rect 1080 476 1082 570
rect 1092 559 1094 573
rect 1090 558 1096 559
rect 1090 554 1091 558
rect 1095 554 1096 558
rect 1090 553 1096 554
rect 1100 528 1102 582
rect 1184 579 1186 602
rect 1183 578 1187 579
rect 1183 573 1187 574
rect 1184 554 1186 573
rect 1182 553 1188 554
rect 1182 549 1183 553
rect 1187 549 1188 553
rect 1182 548 1188 549
rect 1182 535 1188 536
rect 1182 531 1183 535
rect 1187 531 1188 535
rect 1182 530 1188 531
rect 1098 527 1104 528
rect 1098 523 1099 527
rect 1103 523 1104 527
rect 1098 522 1104 523
rect 1086 517 1092 518
rect 1086 513 1087 517
rect 1091 513 1092 517
rect 1086 512 1092 513
rect 1088 499 1090 512
rect 1184 499 1186 530
rect 1087 498 1091 499
rect 1087 493 1091 494
rect 1095 498 1099 499
rect 1095 493 1099 494
rect 1183 498 1187 499
rect 1183 493 1187 494
rect 1096 488 1098 493
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 483 1100 487
rect 1094 482 1100 483
rect 1078 475 1084 476
rect 1078 471 1079 475
rect 1083 471 1084 475
rect 1078 470 1084 471
rect 1184 470 1186 493
rect 1182 469 1188 470
rect 1182 465 1183 469
rect 1187 465 1188 469
rect 1182 464 1188 465
rect 1078 451 1084 452
rect 1078 447 1079 451
rect 1083 447 1084 451
rect 1182 451 1188 452
rect 1182 447 1183 451
rect 1187 447 1188 451
rect 1010 446 1016 447
rect 1078 446 1084 447
rect 1098 446 1104 447
rect 1182 446 1188 447
rect 1010 442 1011 446
rect 1015 442 1016 446
rect 1010 441 1016 442
rect 938 431 944 432
rect 938 427 939 431
rect 943 427 944 431
rect 938 426 944 427
rect 1012 423 1014 441
rect 1080 432 1082 446
rect 1098 442 1099 446
rect 1103 442 1104 446
rect 1098 441 1104 442
rect 1078 431 1084 432
rect 1078 427 1079 431
rect 1083 427 1084 431
rect 1078 426 1084 427
rect 1100 423 1102 441
rect 1106 431 1112 432
rect 1106 427 1107 431
rect 1111 427 1112 431
rect 1106 426 1112 427
rect 835 422 839 423
rect 747 417 751 418
rect 806 419 812 420
rect 638 411 644 412
rect 638 407 639 411
rect 643 407 644 411
rect 638 406 644 407
rect 622 387 628 388
rect 622 383 623 387
rect 627 383 628 387
rect 622 382 628 383
rect 640 372 642 406
rect 660 403 662 417
rect 748 403 750 417
rect 806 415 807 419
rect 811 415 812 419
rect 806 414 812 415
rect 814 419 820 420
rect 814 415 815 419
rect 819 415 820 419
rect 835 417 839 418
rect 923 422 927 423
rect 1011 422 1015 423
rect 923 417 927 418
rect 938 419 944 420
rect 814 414 820 415
rect 658 402 664 403
rect 658 398 659 402
rect 663 398 664 402
rect 658 397 664 398
rect 746 402 752 403
rect 746 398 747 402
rect 751 398 752 402
rect 746 397 752 398
rect 816 372 818 414
rect 836 403 838 417
rect 924 403 926 417
rect 938 415 939 419
rect 943 415 944 419
rect 938 414 944 415
rect 990 419 996 420
rect 990 415 991 419
rect 995 415 996 419
rect 1099 422 1103 423
rect 1011 417 1015 418
rect 1078 419 1084 420
rect 990 414 996 415
rect 834 402 840 403
rect 834 398 835 402
rect 839 398 840 402
rect 834 397 840 398
rect 922 402 928 403
rect 922 398 923 402
rect 927 398 928 402
rect 922 397 928 398
rect 855 372 859 373
rect 455 367 459 368
rect 462 371 468 372
rect 462 367 463 371
rect 467 367 468 371
rect 462 366 468 367
rect 550 371 556 372
rect 550 367 551 371
rect 555 367 556 371
rect 550 366 556 367
rect 638 371 644 372
rect 638 367 639 371
rect 643 367 644 371
rect 638 366 644 367
rect 814 371 820 372
rect 814 367 815 371
rect 819 367 820 371
rect 855 367 859 368
rect 902 371 908 372
rect 902 367 903 371
rect 907 367 908 371
rect 814 366 820 367
rect 390 361 396 362
rect 390 357 391 361
rect 395 357 396 361
rect 390 356 396 357
rect 478 361 484 362
rect 478 357 479 361
rect 483 357 484 361
rect 478 356 484 357
rect 566 361 572 362
rect 566 357 567 361
rect 571 357 572 361
rect 566 356 572 357
rect 654 361 660 362
rect 654 357 655 361
rect 659 357 660 361
rect 654 356 660 357
rect 742 361 748 362
rect 742 357 743 361
rect 747 357 748 361
rect 742 356 748 357
rect 830 361 836 362
rect 830 357 831 361
rect 835 357 836 361
rect 830 356 836 357
rect 392 351 394 356
rect 480 351 482 356
rect 568 351 570 356
rect 656 351 658 356
rect 744 351 746 356
rect 832 351 834 356
rect 111 350 115 351
rect 111 345 115 346
rect 367 350 371 351
rect 367 345 371 346
rect 391 350 395 351
rect 391 345 395 346
rect 479 350 483 351
rect 479 345 483 346
rect 567 350 571 351
rect 567 345 571 346
rect 599 350 603 351
rect 599 345 603 346
rect 655 350 659 351
rect 655 345 659 346
rect 727 350 731 351
rect 727 345 731 346
rect 743 350 747 351
rect 743 345 747 346
rect 831 350 835 351
rect 831 345 835 346
rect 112 322 114 345
rect 368 340 370 345
rect 480 340 482 345
rect 600 340 602 345
rect 728 340 730 345
rect 366 339 372 340
rect 366 335 367 339
rect 371 335 372 339
rect 366 334 372 335
rect 478 339 484 340
rect 478 335 479 339
rect 483 335 484 339
rect 478 334 484 335
rect 598 339 604 340
rect 598 335 599 339
rect 603 335 604 339
rect 598 334 604 335
rect 726 339 732 340
rect 726 335 727 339
rect 731 335 732 339
rect 726 334 732 335
rect 856 332 858 367
rect 902 366 908 367
rect 863 350 867 351
rect 863 345 867 346
rect 864 340 866 345
rect 862 339 868 340
rect 862 335 863 339
rect 867 335 868 339
rect 862 334 868 335
rect 854 331 860 332
rect 854 327 855 331
rect 859 327 860 331
rect 854 326 860 327
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 110 316 116 317
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 110 298 116 299
rect 370 298 376 299
rect 112 267 114 298
rect 370 294 371 298
rect 375 294 376 298
rect 370 293 376 294
rect 482 298 488 299
rect 482 294 483 298
rect 487 294 488 298
rect 482 293 488 294
rect 602 298 608 299
rect 602 294 603 298
rect 607 294 608 298
rect 602 293 608 294
rect 730 298 736 299
rect 730 294 731 298
rect 735 294 736 298
rect 730 293 736 294
rect 866 298 872 299
rect 866 294 867 298
rect 871 294 872 298
rect 866 293 872 294
rect 372 267 374 293
rect 484 267 486 293
rect 604 267 606 293
rect 732 267 734 293
rect 868 267 870 293
rect 904 284 906 366
rect 918 361 924 362
rect 918 357 919 361
rect 923 357 924 361
rect 918 356 924 357
rect 920 351 922 356
rect 919 350 923 351
rect 919 345 923 346
rect 940 332 942 414
rect 992 372 994 414
rect 1012 403 1014 417
rect 1078 415 1079 419
rect 1083 415 1084 419
rect 1099 417 1103 418
rect 1078 414 1084 415
rect 1010 402 1016 403
rect 1010 398 1011 402
rect 1015 398 1016 402
rect 1010 397 1016 398
rect 1080 372 1082 414
rect 1100 403 1102 417
rect 1098 402 1104 403
rect 1098 398 1099 402
rect 1103 398 1104 402
rect 1098 397 1104 398
rect 1108 372 1110 426
rect 1184 423 1186 446
rect 1183 422 1187 423
rect 1183 417 1187 418
rect 1184 398 1186 417
rect 1182 397 1188 398
rect 1182 393 1183 397
rect 1187 393 1188 397
rect 1182 392 1188 393
rect 1182 379 1188 380
rect 1182 375 1183 379
rect 1187 375 1188 379
rect 1182 374 1188 375
rect 990 371 996 372
rect 990 367 991 371
rect 995 367 996 371
rect 990 366 996 367
rect 1078 371 1084 372
rect 1078 367 1079 371
rect 1083 367 1084 371
rect 1078 366 1084 367
rect 1106 371 1112 372
rect 1106 367 1107 371
rect 1111 367 1112 371
rect 1106 366 1112 367
rect 1006 361 1012 362
rect 1006 357 1007 361
rect 1011 357 1012 361
rect 1006 356 1012 357
rect 1094 361 1100 362
rect 1094 357 1095 361
rect 1099 357 1100 361
rect 1094 356 1100 357
rect 1008 351 1010 356
rect 1096 351 1098 356
rect 1184 351 1186 374
rect 1007 350 1011 351
rect 1007 345 1011 346
rect 1095 350 1099 351
rect 1095 345 1099 346
rect 1183 350 1187 351
rect 1183 345 1187 346
rect 1008 340 1010 345
rect 1006 339 1012 340
rect 1006 335 1007 339
rect 1011 335 1012 339
rect 1006 334 1012 335
rect 938 331 944 332
rect 938 327 939 331
rect 943 327 944 331
rect 938 326 944 327
rect 1184 322 1186 345
rect 1182 321 1188 322
rect 1182 317 1183 321
rect 1187 317 1188 321
rect 1182 316 1188 317
rect 1182 303 1188 304
rect 1182 299 1183 303
rect 1187 299 1188 303
rect 1010 298 1016 299
rect 1182 298 1188 299
rect 1010 294 1011 298
rect 1015 294 1016 298
rect 1010 293 1016 294
rect 902 283 908 284
rect 902 279 903 283
rect 907 279 908 283
rect 902 278 908 279
rect 1012 267 1014 293
rect 1184 267 1186 298
rect 111 266 115 267
rect 111 261 115 262
rect 203 266 207 267
rect 291 266 295 267
rect 203 261 207 262
rect 218 263 224 264
rect 112 242 114 261
rect 204 247 206 261
rect 218 259 219 263
rect 223 259 224 263
rect 218 258 224 259
rect 270 263 276 264
rect 270 259 271 263
rect 275 259 276 263
rect 371 266 375 267
rect 291 261 295 262
rect 358 263 364 264
rect 270 258 276 259
rect 202 246 208 247
rect 202 242 203 246
rect 207 242 208 246
rect 110 241 116 242
rect 202 241 208 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 110 223 116 224
rect 110 219 111 223
rect 115 219 116 223
rect 110 218 116 219
rect 112 167 114 218
rect 198 205 204 206
rect 198 201 199 205
rect 203 201 204 205
rect 198 200 204 201
rect 200 167 202 200
rect 220 192 222 258
rect 272 216 274 258
rect 292 247 294 261
rect 358 259 359 263
rect 363 259 364 263
rect 371 261 375 262
rect 379 266 383 267
rect 467 266 471 267
rect 379 261 383 262
rect 446 263 452 264
rect 358 258 364 259
rect 290 246 296 247
rect 290 242 291 246
rect 295 242 296 246
rect 290 241 296 242
rect 360 216 362 258
rect 380 247 382 261
rect 446 259 447 263
rect 451 259 452 263
rect 467 261 471 262
rect 483 266 487 267
rect 555 266 559 267
rect 483 261 487 262
rect 534 263 540 264
rect 446 258 452 259
rect 378 246 384 247
rect 378 242 379 246
rect 383 242 384 246
rect 378 241 384 242
rect 448 216 450 258
rect 468 247 470 261
rect 534 259 535 263
rect 539 259 540 263
rect 555 261 559 262
rect 603 266 607 267
rect 603 261 607 262
rect 731 266 735 267
rect 731 261 735 262
rect 867 266 871 267
rect 867 261 871 262
rect 1011 266 1015 267
rect 1011 261 1015 262
rect 1183 266 1187 267
rect 1183 261 1187 262
rect 534 258 540 259
rect 466 246 472 247
rect 466 242 467 246
rect 471 242 472 246
rect 466 241 472 242
rect 536 216 538 258
rect 556 247 558 261
rect 554 246 560 247
rect 554 242 555 246
rect 559 242 560 246
rect 1184 242 1186 261
rect 554 241 560 242
rect 1182 241 1188 242
rect 1182 237 1183 241
rect 1187 237 1188 241
rect 1182 236 1188 237
rect 1182 223 1188 224
rect 1182 219 1183 223
rect 1187 219 1188 223
rect 1182 218 1188 219
rect 270 215 276 216
rect 270 211 271 215
rect 275 211 276 215
rect 270 210 276 211
rect 358 215 364 216
rect 358 211 359 215
rect 363 211 364 215
rect 358 210 364 211
rect 446 215 452 216
rect 446 211 447 215
rect 451 211 452 215
rect 446 210 452 211
rect 534 215 540 216
rect 534 211 535 215
rect 539 211 540 215
rect 534 210 540 211
rect 286 205 292 206
rect 286 201 287 205
rect 291 201 292 205
rect 286 200 292 201
rect 374 205 380 206
rect 374 201 375 205
rect 379 201 380 205
rect 374 200 380 201
rect 462 205 468 206
rect 462 201 463 205
rect 467 201 468 205
rect 462 200 468 201
rect 550 205 556 206
rect 550 201 551 205
rect 555 201 556 205
rect 550 200 556 201
rect 218 191 224 192
rect 218 187 219 191
rect 223 187 224 191
rect 218 186 224 187
rect 288 167 290 200
rect 376 167 378 200
rect 464 167 466 200
rect 552 167 554 200
rect 750 191 756 192
rect 750 187 751 191
rect 755 187 756 191
rect 750 186 756 187
rect 111 166 115 167
rect 111 161 115 162
rect 143 166 147 167
rect 143 161 147 162
rect 199 166 203 167
rect 199 161 203 162
rect 231 166 235 167
rect 231 161 235 162
rect 287 166 291 167
rect 287 161 291 162
rect 319 166 323 167
rect 319 161 323 162
rect 375 166 379 167
rect 375 161 379 162
rect 407 166 411 167
rect 407 161 411 162
rect 463 166 467 167
rect 463 161 467 162
rect 495 166 499 167
rect 495 161 499 162
rect 551 166 555 167
rect 551 161 555 162
rect 583 166 587 167
rect 583 161 587 162
rect 671 166 675 167
rect 671 161 675 162
rect 112 138 114 161
rect 144 156 146 161
rect 232 156 234 161
rect 320 156 322 161
rect 408 156 410 161
rect 496 156 498 161
rect 584 156 586 161
rect 672 156 674 161
rect 142 155 148 156
rect 142 151 143 155
rect 147 151 148 155
rect 142 150 148 151
rect 230 155 236 156
rect 230 151 231 155
rect 235 151 236 155
rect 230 150 236 151
rect 318 155 324 156
rect 318 151 319 155
rect 323 151 324 155
rect 318 150 324 151
rect 406 155 412 156
rect 406 151 407 155
rect 411 151 412 155
rect 406 150 412 151
rect 494 155 500 156
rect 494 151 495 155
rect 499 151 500 155
rect 494 150 500 151
rect 582 155 588 156
rect 582 151 583 155
rect 587 151 588 155
rect 582 150 588 151
rect 670 155 676 156
rect 670 151 671 155
rect 675 151 676 155
rect 670 150 676 151
rect 752 148 754 186
rect 1184 167 1186 218
rect 759 166 763 167
rect 759 161 763 162
rect 1183 166 1187 167
rect 1183 161 1187 162
rect 760 156 762 161
rect 758 155 764 156
rect 758 151 759 155
rect 763 151 764 155
rect 758 150 764 151
rect 750 147 756 148
rect 390 143 396 144
rect 390 139 391 143
rect 395 139 396 143
rect 390 138 396 139
rect 478 143 484 144
rect 478 139 479 143
rect 483 139 484 143
rect 478 138 484 139
rect 566 143 572 144
rect 566 139 567 143
rect 571 139 572 143
rect 566 138 572 139
rect 654 143 660 144
rect 654 139 655 143
rect 659 139 660 143
rect 654 138 660 139
rect 742 143 748 144
rect 742 139 743 143
rect 747 139 748 143
rect 750 143 751 147
rect 755 143 756 147
rect 750 142 756 143
rect 742 138 748 139
rect 1184 138 1186 161
rect 110 137 116 138
rect 110 133 111 137
rect 115 133 116 137
rect 110 132 116 133
rect 110 119 116 120
rect 110 115 111 119
rect 115 115 116 119
rect 110 114 116 115
rect 146 114 152 115
rect 112 95 114 114
rect 146 110 147 114
rect 151 110 152 114
rect 146 109 152 110
rect 234 114 240 115
rect 234 110 235 114
rect 239 110 240 114
rect 234 109 240 110
rect 322 114 328 115
rect 322 110 323 114
rect 327 110 328 114
rect 322 109 328 110
rect 148 95 150 109
rect 236 95 238 109
rect 324 95 326 109
rect 392 100 394 138
rect 410 114 416 115
rect 410 110 411 114
rect 415 110 416 114
rect 410 109 416 110
rect 390 99 396 100
rect 390 95 391 99
rect 395 95 396 99
rect 412 95 414 109
rect 480 100 482 138
rect 498 114 504 115
rect 498 110 499 114
rect 503 110 504 114
rect 498 109 504 110
rect 478 99 484 100
rect 478 95 479 99
rect 483 95 484 99
rect 500 95 502 109
rect 568 100 570 138
rect 586 114 592 115
rect 586 110 587 114
rect 591 110 592 114
rect 586 109 592 110
rect 566 99 572 100
rect 566 95 567 99
rect 571 95 572 99
rect 588 95 590 109
rect 656 100 658 138
rect 674 114 680 115
rect 674 110 675 114
rect 679 110 680 114
rect 674 109 680 110
rect 654 99 660 100
rect 654 95 655 99
rect 659 95 660 99
rect 676 95 678 109
rect 744 100 746 138
rect 1182 137 1188 138
rect 1182 133 1183 137
rect 1187 133 1188 137
rect 1182 132 1188 133
rect 1182 119 1188 120
rect 1182 115 1183 119
rect 1187 115 1188 119
rect 762 114 768 115
rect 1182 114 1188 115
rect 762 110 763 114
rect 767 110 768 114
rect 762 109 768 110
rect 742 99 748 100
rect 742 95 743 99
rect 747 95 748 99
rect 764 95 766 109
rect 1184 95 1186 114
rect 111 94 115 95
rect 111 89 115 90
rect 147 94 151 95
rect 147 89 151 90
rect 235 94 239 95
rect 235 89 239 90
rect 323 94 327 95
rect 390 94 396 95
rect 411 94 415 95
rect 478 94 484 95
rect 499 94 503 95
rect 566 94 572 95
rect 587 94 591 95
rect 654 94 660 95
rect 675 94 679 95
rect 742 94 748 95
rect 763 94 767 95
rect 323 89 327 90
rect 411 89 415 90
rect 499 89 503 90
rect 587 89 591 90
rect 675 89 679 90
rect 763 89 767 90
rect 1183 94 1187 95
rect 1183 89 1187 90
<< m4c >>
rect 111 1278 115 1282
rect 575 1278 579 1282
rect 1183 1278 1187 1282
rect 111 1206 115 1210
rect 219 1206 223 1210
rect 307 1206 311 1210
rect 111 1118 115 1122
rect 215 1118 219 1122
rect 395 1206 399 1210
rect 483 1206 487 1210
rect 571 1206 575 1210
rect 579 1206 583 1210
rect 667 1206 671 1210
rect 771 1206 775 1210
rect 883 1206 887 1210
rect 1003 1206 1007 1210
rect 1099 1206 1103 1210
rect 1183 1206 1187 1210
rect 303 1118 307 1122
rect 359 1118 363 1122
rect 391 1118 395 1122
rect 479 1118 483 1122
rect 503 1118 507 1122
rect 567 1118 571 1122
rect 647 1118 651 1122
rect 663 1118 667 1122
rect 767 1118 771 1122
rect 799 1118 803 1122
rect 111 1038 115 1042
rect 219 1038 223 1042
rect 243 1038 247 1042
rect 363 1038 367 1042
rect 395 1038 399 1042
rect 507 1038 511 1042
rect 547 1038 551 1042
rect 651 1038 655 1042
rect 707 1038 711 1042
rect 879 1118 883 1122
rect 951 1118 955 1122
rect 999 1118 1003 1122
rect 1095 1118 1099 1122
rect 1183 1118 1187 1122
rect 803 1038 807 1042
rect 875 1038 879 1042
rect 955 1038 959 1042
rect 1043 1038 1047 1042
rect 1099 1038 1103 1042
rect 111 958 115 962
rect 239 958 243 962
rect 327 958 331 962
rect 391 958 395 962
rect 439 958 443 962
rect 543 958 547 962
rect 559 958 563 962
rect 687 958 691 962
rect 703 958 707 962
rect 815 958 819 962
rect 111 878 115 882
rect 331 878 335 882
rect 403 878 407 882
rect 443 878 447 882
rect 111 806 115 810
rect 375 806 379 810
rect 515 878 519 882
rect 563 878 567 882
rect 643 878 647 882
rect 691 878 695 882
rect 871 958 875 962
rect 951 958 955 962
rect 1039 958 1043 962
rect 1183 1038 1187 1042
rect 1087 958 1091 962
rect 1183 958 1187 962
rect 779 878 783 882
rect 819 878 823 882
rect 915 878 919 882
rect 955 878 959 882
rect 1059 878 1063 882
rect 1091 878 1095 882
rect 1183 878 1187 882
rect 399 806 403 810
rect 511 806 515 810
rect 519 806 523 810
rect 639 806 643 810
rect 663 806 667 810
rect 775 806 779 810
rect 815 806 819 810
rect 111 730 115 734
rect 147 730 151 734
rect 267 730 271 734
rect 111 650 115 654
rect 143 650 147 654
rect 379 730 383 734
rect 411 730 415 734
rect 523 730 527 734
rect 563 730 567 734
rect 667 730 671 734
rect 911 806 915 810
rect 967 806 971 810
rect 1055 806 1059 810
rect 1095 806 1099 810
rect 1183 806 1187 810
rect 731 730 735 734
rect 819 730 823 734
rect 907 730 911 734
rect 971 730 975 734
rect 1091 730 1095 734
rect 1099 730 1103 734
rect 1183 730 1187 734
rect 247 650 251 654
rect 263 650 267 654
rect 391 650 395 654
rect 407 650 411 654
rect 551 650 555 654
rect 559 650 563 654
rect 719 650 723 654
rect 727 650 731 654
rect 903 650 907 654
rect 411 592 415 596
rect 623 592 627 596
rect 111 574 115 578
rect 147 574 151 578
rect 251 574 255 578
rect 267 574 271 578
rect 379 574 383 578
rect 395 574 399 578
rect 283 560 287 564
rect 499 574 503 578
rect 555 574 559 578
rect 635 574 639 578
rect 579 560 583 564
rect 723 574 727 578
rect 779 574 783 578
rect 907 574 911 578
rect 1087 650 1091 654
rect 1183 650 1187 654
rect 931 574 935 578
rect 111 494 115 498
rect 263 494 267 498
rect 375 494 379 498
rect 463 494 467 498
rect 495 494 499 498
rect 551 494 555 498
rect 631 494 635 498
rect 639 494 643 498
rect 735 494 739 498
rect 775 494 779 498
rect 111 418 115 422
rect 395 418 399 422
rect 467 418 471 422
rect 483 418 487 422
rect 555 418 559 422
rect 571 418 575 422
rect 643 418 647 422
rect 659 418 663 422
rect 739 418 743 422
rect 747 418 751 422
rect 1091 574 1095 578
rect 831 494 835 498
rect 919 494 923 498
rect 927 494 931 498
rect 1007 494 1011 498
rect 1183 574 1187 578
rect 1087 494 1091 498
rect 1095 494 1099 498
rect 1183 494 1187 498
rect 835 418 839 422
rect 923 418 927 422
rect 1011 418 1015 422
rect 455 368 459 372
rect 855 368 859 372
rect 111 346 115 350
rect 367 346 371 350
rect 391 346 395 350
rect 479 346 483 350
rect 567 346 571 350
rect 599 346 603 350
rect 655 346 659 350
rect 727 346 731 350
rect 743 346 747 350
rect 831 346 835 350
rect 863 346 867 350
rect 919 346 923 350
rect 1099 418 1103 422
rect 1183 418 1187 422
rect 1007 346 1011 350
rect 1095 346 1099 350
rect 1183 346 1187 350
rect 111 262 115 266
rect 203 262 207 266
rect 291 262 295 266
rect 371 262 375 266
rect 379 262 383 266
rect 467 262 471 266
rect 483 262 487 266
rect 555 262 559 266
rect 603 262 607 266
rect 731 262 735 266
rect 867 262 871 266
rect 1011 262 1015 266
rect 1183 262 1187 266
rect 111 162 115 166
rect 143 162 147 166
rect 199 162 203 166
rect 231 162 235 166
rect 287 162 291 166
rect 319 162 323 166
rect 375 162 379 166
rect 407 162 411 166
rect 463 162 467 166
rect 495 162 499 166
rect 551 162 555 166
rect 583 162 587 166
rect 671 162 675 166
rect 759 162 763 166
rect 1183 162 1187 166
rect 111 90 115 94
rect 147 90 151 94
rect 235 90 239 94
rect 323 90 327 94
rect 411 90 415 94
rect 499 90 503 94
rect 587 90 591 94
rect 675 90 679 94
rect 763 90 767 94
rect 1183 90 1187 94
<< m4 >>
rect 96 1277 97 1283
rect 103 1282 1219 1283
rect 103 1278 111 1282
rect 115 1278 575 1282
rect 579 1278 1183 1282
rect 1187 1278 1219 1282
rect 103 1277 1219 1278
rect 1225 1277 1226 1283
rect 84 1205 85 1211
rect 91 1210 1207 1211
rect 91 1206 111 1210
rect 115 1206 219 1210
rect 223 1206 307 1210
rect 311 1206 395 1210
rect 399 1206 483 1210
rect 487 1206 571 1210
rect 575 1206 579 1210
rect 583 1206 667 1210
rect 671 1206 771 1210
rect 775 1206 883 1210
rect 887 1206 1003 1210
rect 1007 1206 1099 1210
rect 1103 1206 1183 1210
rect 1187 1206 1207 1210
rect 91 1205 1207 1206
rect 1213 1205 1214 1211
rect 96 1117 97 1123
rect 103 1122 1219 1123
rect 103 1118 111 1122
rect 115 1118 215 1122
rect 219 1118 303 1122
rect 307 1118 359 1122
rect 363 1118 391 1122
rect 395 1118 479 1122
rect 483 1118 503 1122
rect 507 1118 567 1122
rect 571 1118 647 1122
rect 651 1118 663 1122
rect 667 1118 767 1122
rect 771 1118 799 1122
rect 803 1118 879 1122
rect 883 1118 951 1122
rect 955 1118 999 1122
rect 1003 1118 1095 1122
rect 1099 1118 1183 1122
rect 1187 1118 1219 1122
rect 103 1117 1219 1118
rect 1225 1117 1226 1123
rect 84 1037 85 1043
rect 91 1042 1207 1043
rect 91 1038 111 1042
rect 115 1038 219 1042
rect 223 1038 243 1042
rect 247 1038 363 1042
rect 367 1038 395 1042
rect 399 1038 507 1042
rect 511 1038 547 1042
rect 551 1038 651 1042
rect 655 1038 707 1042
rect 711 1038 803 1042
rect 807 1038 875 1042
rect 879 1038 955 1042
rect 959 1038 1043 1042
rect 1047 1038 1099 1042
rect 1103 1038 1183 1042
rect 1187 1038 1207 1042
rect 91 1037 1207 1038
rect 1213 1037 1214 1043
rect 96 957 97 963
rect 103 962 1219 963
rect 103 958 111 962
rect 115 958 239 962
rect 243 958 327 962
rect 331 958 391 962
rect 395 958 439 962
rect 443 958 543 962
rect 547 958 559 962
rect 563 958 687 962
rect 691 958 703 962
rect 707 958 815 962
rect 819 958 871 962
rect 875 958 951 962
rect 955 958 1039 962
rect 1043 958 1087 962
rect 1091 958 1183 962
rect 1187 958 1219 962
rect 103 957 1219 958
rect 1225 957 1226 963
rect 84 877 85 883
rect 91 882 1207 883
rect 91 878 111 882
rect 115 878 331 882
rect 335 878 403 882
rect 407 878 443 882
rect 447 878 515 882
rect 519 878 563 882
rect 567 878 643 882
rect 647 878 691 882
rect 695 878 779 882
rect 783 878 819 882
rect 823 878 915 882
rect 919 878 955 882
rect 959 878 1059 882
rect 1063 878 1091 882
rect 1095 878 1183 882
rect 1187 878 1207 882
rect 91 877 1207 878
rect 1213 877 1214 883
rect 96 805 97 811
rect 103 810 1219 811
rect 103 806 111 810
rect 115 806 375 810
rect 379 806 399 810
rect 403 806 511 810
rect 515 806 519 810
rect 523 806 639 810
rect 643 806 663 810
rect 667 806 775 810
rect 779 806 815 810
rect 819 806 911 810
rect 915 806 967 810
rect 971 806 1055 810
rect 1059 806 1095 810
rect 1099 806 1183 810
rect 1187 806 1219 810
rect 103 805 1219 806
rect 1225 805 1226 811
rect 84 729 85 735
rect 91 734 1207 735
rect 91 730 111 734
rect 115 730 147 734
rect 151 730 267 734
rect 271 730 379 734
rect 383 730 411 734
rect 415 730 523 734
rect 527 730 563 734
rect 567 730 667 734
rect 671 730 731 734
rect 735 730 819 734
rect 823 730 907 734
rect 911 730 971 734
rect 975 730 1091 734
rect 1095 730 1099 734
rect 1103 730 1183 734
rect 1187 730 1207 734
rect 91 729 1207 730
rect 1213 729 1214 735
rect 96 649 97 655
rect 103 654 1219 655
rect 103 650 111 654
rect 115 650 143 654
rect 147 650 247 654
rect 251 650 263 654
rect 267 650 391 654
rect 395 650 407 654
rect 411 650 551 654
rect 555 650 559 654
rect 563 650 719 654
rect 723 650 727 654
rect 731 650 903 654
rect 907 650 1087 654
rect 1091 650 1183 654
rect 1187 650 1219 654
rect 103 649 1219 650
rect 1225 649 1226 655
rect 410 596 416 597
rect 622 596 628 597
rect 410 592 411 596
rect 415 592 623 596
rect 627 592 628 596
rect 410 591 416 592
rect 622 591 628 592
rect 84 573 85 579
rect 91 578 1207 579
rect 91 574 111 578
rect 115 574 147 578
rect 151 574 251 578
rect 255 574 267 578
rect 271 574 379 578
rect 383 574 395 578
rect 399 574 499 578
rect 503 574 555 578
rect 559 574 635 578
rect 639 574 723 578
rect 727 574 779 578
rect 783 574 907 578
rect 911 574 931 578
rect 935 574 1091 578
rect 1095 574 1183 578
rect 1187 574 1207 578
rect 91 573 1207 574
rect 1213 573 1214 579
rect 282 564 288 565
rect 578 564 584 565
rect 282 560 283 564
rect 287 560 579 564
rect 583 560 584 564
rect 282 559 288 560
rect 578 559 584 560
rect 96 493 97 499
rect 103 498 1219 499
rect 103 494 111 498
rect 115 494 263 498
rect 267 494 375 498
rect 379 494 463 498
rect 467 494 495 498
rect 499 494 551 498
rect 555 494 631 498
rect 635 494 639 498
rect 643 494 735 498
rect 739 494 775 498
rect 779 494 831 498
rect 835 494 919 498
rect 923 494 927 498
rect 931 494 1007 498
rect 1011 494 1087 498
rect 1091 494 1095 498
rect 1099 494 1183 498
rect 1187 494 1219 498
rect 103 493 1219 494
rect 1225 493 1226 499
rect 84 417 85 423
rect 91 422 1207 423
rect 91 418 111 422
rect 115 418 395 422
rect 399 418 467 422
rect 471 418 483 422
rect 487 418 555 422
rect 559 418 571 422
rect 575 418 643 422
rect 647 418 659 422
rect 663 418 739 422
rect 743 418 747 422
rect 751 418 835 422
rect 839 418 923 422
rect 927 418 1011 422
rect 1015 418 1099 422
rect 1103 418 1183 422
rect 1187 418 1207 422
rect 91 417 1207 418
rect 1213 417 1214 423
rect 454 372 460 373
rect 854 372 860 373
rect 454 368 455 372
rect 459 368 855 372
rect 859 368 860 372
rect 454 367 460 368
rect 854 367 860 368
rect 96 345 97 351
rect 103 350 1219 351
rect 103 346 111 350
rect 115 346 367 350
rect 371 346 391 350
rect 395 346 479 350
rect 483 346 567 350
rect 571 346 599 350
rect 603 346 655 350
rect 659 346 727 350
rect 731 346 743 350
rect 747 346 831 350
rect 835 346 863 350
rect 867 346 919 350
rect 923 346 1007 350
rect 1011 346 1095 350
rect 1099 346 1183 350
rect 1187 346 1219 350
rect 103 345 1219 346
rect 1225 345 1226 351
rect 84 261 85 267
rect 91 266 1207 267
rect 91 262 111 266
rect 115 262 203 266
rect 207 262 291 266
rect 295 262 371 266
rect 375 262 379 266
rect 383 262 467 266
rect 471 262 483 266
rect 487 262 555 266
rect 559 262 603 266
rect 607 262 731 266
rect 735 262 867 266
rect 871 262 1011 266
rect 1015 262 1183 266
rect 1187 262 1207 266
rect 91 261 1207 262
rect 1213 261 1214 267
rect 96 161 97 167
rect 103 166 1219 167
rect 103 162 111 166
rect 115 162 143 166
rect 147 162 199 166
rect 203 162 231 166
rect 235 162 287 166
rect 291 162 319 166
rect 323 162 375 166
rect 379 162 407 166
rect 411 162 463 166
rect 467 162 495 166
rect 499 162 551 166
rect 555 162 583 166
rect 587 162 671 166
rect 675 162 759 166
rect 763 162 1183 166
rect 1187 162 1219 166
rect 103 161 1219 162
rect 1225 161 1226 167
rect 84 89 85 95
rect 91 94 1207 95
rect 91 90 111 94
rect 115 90 147 94
rect 151 90 235 94
rect 239 90 323 94
rect 327 90 411 94
rect 415 90 499 94
rect 503 90 587 94
rect 591 90 675 94
rect 679 90 763 94
rect 767 90 1183 94
rect 1187 90 1207 94
rect 91 89 1207 90
rect 1213 89 1214 95
<< m5c >>
rect 97 1277 103 1283
rect 1219 1277 1225 1283
rect 85 1205 91 1211
rect 1207 1205 1213 1211
rect 97 1117 103 1123
rect 1219 1117 1225 1123
rect 85 1037 91 1043
rect 1207 1037 1213 1043
rect 97 957 103 963
rect 1219 957 1225 963
rect 85 877 91 883
rect 1207 877 1213 883
rect 97 805 103 811
rect 1219 805 1225 811
rect 85 729 91 735
rect 1207 729 1213 735
rect 97 649 103 655
rect 1219 649 1225 655
rect 85 573 91 579
rect 1207 573 1213 579
rect 97 493 103 499
rect 1219 493 1225 499
rect 85 417 91 423
rect 1207 417 1213 423
rect 97 345 103 351
rect 1219 345 1225 351
rect 85 261 91 267
rect 1207 261 1213 267
rect 97 161 103 167
rect 1219 161 1225 167
rect 85 89 91 95
rect 1207 89 1213 95
<< m5 >>
rect 84 1211 92 1296
rect 84 1205 85 1211
rect 91 1205 92 1211
rect 84 1043 92 1205
rect 84 1037 85 1043
rect 91 1037 92 1043
rect 84 883 92 1037
rect 84 877 85 883
rect 91 877 92 883
rect 84 735 92 877
rect 84 729 85 735
rect 91 729 92 735
rect 84 579 92 729
rect 84 573 85 579
rect 91 573 92 579
rect 84 423 92 573
rect 84 417 85 423
rect 91 417 92 423
rect 84 267 92 417
rect 84 261 85 267
rect 91 261 92 267
rect 84 95 92 261
rect 84 89 85 95
rect 91 89 92 95
rect 84 72 92 89
rect 96 1283 104 1296
rect 96 1277 97 1283
rect 103 1277 104 1283
rect 96 1123 104 1277
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 963 104 1117
rect 96 957 97 963
rect 103 957 104 963
rect 96 811 104 957
rect 96 805 97 811
rect 103 805 104 811
rect 96 655 104 805
rect 96 649 97 655
rect 103 649 104 655
rect 96 499 104 649
rect 96 493 97 499
rect 103 493 104 499
rect 96 351 104 493
rect 96 345 97 351
rect 103 345 104 351
rect 96 167 104 345
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 1206 1211 1214 1296
rect 1206 1205 1207 1211
rect 1213 1205 1214 1211
rect 1206 1043 1214 1205
rect 1206 1037 1207 1043
rect 1213 1037 1214 1043
rect 1206 883 1214 1037
rect 1206 877 1207 883
rect 1213 877 1214 883
rect 1206 735 1214 877
rect 1206 729 1207 735
rect 1213 729 1214 735
rect 1206 579 1214 729
rect 1206 573 1207 579
rect 1213 573 1214 579
rect 1206 423 1214 573
rect 1206 417 1207 423
rect 1213 417 1214 423
rect 1206 267 1214 417
rect 1206 261 1207 267
rect 1213 261 1214 267
rect 1206 95 1214 261
rect 1206 89 1207 95
rect 1213 89 1214 95
rect 1206 72 1214 89
rect 1218 1283 1226 1296
rect 1218 1277 1219 1283
rect 1225 1277 1226 1283
rect 1218 1123 1226 1277
rect 1218 1117 1219 1123
rect 1225 1117 1226 1123
rect 1218 963 1226 1117
rect 1218 957 1219 963
rect 1225 957 1226 963
rect 1218 811 1226 957
rect 1218 805 1219 811
rect 1225 805 1226 811
rect 1218 655 1226 805
rect 1218 649 1219 655
rect 1225 649 1226 655
rect 1218 499 1226 649
rect 1218 493 1219 499
rect 1225 493 1226 499
rect 1218 351 1226 493
rect 1218 345 1219 351
rect 1225 345 1226 351
rect 1218 167 1226 345
rect 1218 161 1219 167
rect 1225 161 1226 167
rect 1218 72 1226 161
use _0_0std_0_0cells_0_0LATCH  latch_50_6
timestamp 1730953945
transform 1 0 128 0 1 92
box 7 3 85 69
use welltap_svt  __well_tap__0
timestamp 1730953945
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0LATCH  latch_50_6
timestamp 1730953945
transform 1 0 128 0 1 92
box 7 3 85 69
use welltap_svt  __well_tap__0
timestamp 1730953945
transform 1 0 104 0 1 112
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0LATCH  latch_51_6
timestamp 1730953945
transform 1 0 216 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_51_6
timestamp 1730953945
transform 1 0 216 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_52_6
timestamp 1730953945
transform 1 0 304 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_52_6
timestamp 1730953945
transform 1 0 304 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_53_6
timestamp 1730953945
transform 1 0 392 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_53_6
timestamp 1730953945
transform 1 0 392 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_54_6
timestamp 1730953945
transform 1 0 480 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_54_6
timestamp 1730953945
transform 1 0 480 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_55_6
timestamp 1730953945
transform 1 0 568 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_55_6
timestamp 1730953945
transform 1 0 568 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_56_6
timestamp 1730953945
transform 1 0 656 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_56_6
timestamp 1730953945
transform 1 0 656 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_57_6
timestamp 1730953945
transform 1 0 744 0 1 92
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_57_6
timestamp 1730953945
transform 1 0 744 0 1 92
box 7 3 85 69
use welltap_svt  __well_tap__1
timestamp 1730953945
transform 1 0 1176 0 1 112
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730953945
transform 1 0 1176 0 1 112
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_58_6
timestamp 1730953945
transform 1 0 184 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_58_6
timestamp 1730953945
transform 1 0 184 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_59_6
timestamp 1730953945
transform 1 0 272 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_59_6
timestamp 1730953945
transform 1 0 272 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_510_6
timestamp 1730953945
transform 1 0 360 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_510_6
timestamp 1730953945
transform 1 0 360 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_511_6
timestamp 1730953945
transform 1 0 448 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_511_6
timestamp 1730953945
transform 1 0 448 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_512_6
timestamp 1730953945
transform 1 0 536 0 -1 264
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_512_6
timestamp 1730953945
transform 1 0 536 0 -1 264
box 7 3 85 69
use welltap_svt  __well_tap__2
timestamp 1730953945
transform 1 0 104 0 -1 244
box 8 4 12 24
use welltap_svt  __well_tap__2
timestamp 1730953945
transform 1 0 104 0 -1 244
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_513_6
timestamp 1730953945
transform 1 0 352 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_513_6
timestamp 1730953945
transform 1 0 352 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_514_6
timestamp 1730953945
transform 1 0 464 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_514_6
timestamp 1730953945
transform 1 0 464 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_515_6
timestamp 1730953945
transform 1 0 584 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_515_6
timestamp 1730953945
transform 1 0 584 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_516_6
timestamp 1730953945
transform 1 0 712 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_516_6
timestamp 1730953945
transform 1 0 712 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_517_6
timestamp 1730953945
transform 1 0 848 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_517_6
timestamp 1730953945
transform 1 0 848 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_581_6
timestamp 1730953945
transform 1 0 992 0 1 276
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_581_6
timestamp 1730953945
transform 1 0 992 0 1 276
box 7 3 85 69
use welltap_svt  __well_tap__3
timestamp 1730953945
transform 1 0 1176 0 -1 244
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730953945
transform 1 0 1176 0 -1 244
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730953945
transform 1 0 104 0 1 296
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730953945
transform 1 0 104 0 1 296
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_518_6
timestamp 1730953945
transform 1 0 376 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_518_6
timestamp 1730953945
transform 1 0 376 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_519_6
timestamp 1730953945
transform 1 0 464 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_519_6
timestamp 1730953945
transform 1 0 464 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_520_6
timestamp 1730953945
transform 1 0 552 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_520_6
timestamp 1730953945
transform 1 0 552 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_521_6
timestamp 1730953945
transform 1 0 640 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_521_6
timestamp 1730953945
transform 1 0 640 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_579_6
timestamp 1730953945
transform 1 0 728 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_579_6
timestamp 1730953945
transform 1 0 728 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_580_6
timestamp 1730953945
transform 1 0 816 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_580_6
timestamp 1730953945
transform 1 0 816 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_582_6
timestamp 1730953945
transform 1 0 904 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_582_6
timestamp 1730953945
transform 1 0 904 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_583_6
timestamp 1730953945
transform 1 0 992 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_583_6
timestamp 1730953945
transform 1 0 992 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_584_6
timestamp 1730953945
transform 1 0 1080 0 -1 420
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_584_6
timestamp 1730953945
transform 1 0 1080 0 -1 420
box 7 3 85 69
use welltap_svt  __well_tap__5
timestamp 1730953945
transform 1 0 1176 0 1 296
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730953945
transform 1 0 1176 0 1 296
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730953945
transform 1 0 104 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__6
timestamp 1730953945
transform 1 0 104 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730953945
transform 1 0 1176 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730953945
transform 1 0 1176 0 -1 400
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730953945
transform 1 0 104 0 1 444
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730953945
transform 1 0 104 0 1 444
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_522_6
timestamp 1730953945
transform 1 0 448 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_522_6
timestamp 1730953945
transform 1 0 448 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_523_6
timestamp 1730953945
transform 1 0 536 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_523_6
timestamp 1730953945
transform 1 0 536 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_524_6
timestamp 1730953945
transform 1 0 624 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_524_6
timestamp 1730953945
transform 1 0 624 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_525_6
timestamp 1730953945
transform 1 0 720 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_525_6
timestamp 1730953945
transform 1 0 720 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_526_6
timestamp 1730953945
transform 1 0 816 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_526_6
timestamp 1730953945
transform 1 0 816 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_578_6
timestamp 1730953945
transform 1 0 904 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_578_6
timestamp 1730953945
transform 1 0 904 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_586_6
timestamp 1730953945
transform 1 0 992 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_586_6
timestamp 1730953945
transform 1 0 992 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_585_6
timestamp 1730953945
transform 1 0 1080 0 1 424
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_585_6
timestamp 1730953945
transform 1 0 1080 0 1 424
box 7 3 85 69
use welltap_svt  __well_tap__9
timestamp 1730953945
transform 1 0 1176 0 1 444
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730953945
transform 1 0 1176 0 1 444
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730953945
transform 1 0 104 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730953945
transform 1 0 104 0 -1 556
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_529_6
timestamp 1730953945
transform 1 0 248 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_529_6
timestamp 1730953945
transform 1 0 248 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_530_6
timestamp 1730953945
transform 1 0 360 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_530_6
timestamp 1730953945
transform 1 0 360 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_531_6
timestamp 1730953945
transform 1 0 480 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_531_6
timestamp 1730953945
transform 1 0 480 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_528_6
timestamp 1730953945
transform 1 0 616 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_528_6
timestamp 1730953945
transform 1 0 616 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_527_6
timestamp 1730953945
transform 1 0 760 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_527_6
timestamp 1730953945
transform 1 0 760 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_577_6
timestamp 1730953945
transform 1 0 912 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_577_6
timestamp 1730953945
transform 1 0 912 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_587_6
timestamp 1730953945
transform 1 0 1072 0 -1 576
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_587_6
timestamp 1730953945
transform 1 0 1072 0 -1 576
box 7 3 85 69
use welltap_svt  __well_tap__11
timestamp 1730953945
transform 1 0 1176 0 -1 556
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730953945
transform 1 0 1176 0 -1 556
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_536_6
timestamp 1730953945
transform 1 0 128 0 1 580
box 7 3 85 69
use welltap_svt  __well_tap__12
timestamp 1730953945
transform 1 0 104 0 1 600
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_536_6
timestamp 1730953945
transform 1 0 128 0 1 580
box 7 3 85 69
use welltap_svt  __well_tap__12
timestamp 1730953945
transform 1 0 104 0 1 600
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_535_6
timestamp 1730953945
transform 1 0 232 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_535_6
timestamp 1730953945
transform 1 0 232 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_534_6
timestamp 1730953945
transform 1 0 376 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_534_6
timestamp 1730953945
transform 1 0 376 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_532_6
timestamp 1730953945
transform 1 0 536 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_532_6
timestamp 1730953945
transform 1 0 536 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_533_6
timestamp 1730953945
transform 1 0 704 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_533_6
timestamp 1730953945
transform 1 0 704 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_576_6
timestamp 1730953945
transform 1 0 888 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_576_6
timestamp 1730953945
transform 1 0 888 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_588_6
timestamp 1730953945
transform 1 0 1072 0 1 580
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_588_6
timestamp 1730953945
transform 1 0 1072 0 1 580
box 7 3 85 69
use welltap_svt  __well_tap__13
timestamp 1730953945
transform 1 0 1176 0 1 600
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730953945
transform 1 0 1176 0 1 600
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_537_6
timestamp 1730953945
transform 1 0 128 0 -1 732
box 7 3 85 69
use welltap_svt  __well_tap__14
timestamp 1730953945
transform 1 0 104 0 -1 712
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_537_6
timestamp 1730953945
transform 1 0 128 0 -1 732
box 7 3 85 69
use welltap_svt  __well_tap__14
timestamp 1730953945
transform 1 0 104 0 -1 712
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_538_6
timestamp 1730953945
transform 1 0 248 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_538_6
timestamp 1730953945
transform 1 0 248 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_539_6
timestamp 1730953945
transform 1 0 392 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_539_6
timestamp 1730953945
transform 1 0 392 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_540_6
timestamp 1730953945
transform 1 0 544 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_540_6
timestamp 1730953945
transform 1 0 544 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_541_6
timestamp 1730953945
transform 1 0 712 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_541_6
timestamp 1730953945
transform 1 0 712 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_575_6
timestamp 1730953945
transform 1 0 888 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_575_6
timestamp 1730953945
transform 1 0 888 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_589_6
timestamp 1730953945
transform 1 0 1072 0 -1 732
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_589_6
timestamp 1730953945
transform 1 0 1072 0 -1 732
box 7 3 85 69
use welltap_svt  __well_tap__15
timestamp 1730953945
transform 1 0 1176 0 -1 712
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730953945
transform 1 0 1176 0 -1 712
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730953945
transform 1 0 104 0 1 756
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730953945
transform 1 0 104 0 1 756
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_544_6
timestamp 1730953945
transform 1 0 360 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_544_6
timestamp 1730953945
transform 1 0 360 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_543_6
timestamp 1730953945
transform 1 0 504 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_543_6
timestamp 1730953945
transform 1 0 504 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_542_6
timestamp 1730953945
transform 1 0 648 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_542_6
timestamp 1730953945
transform 1 0 648 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_574_6
timestamp 1730953945
transform 1 0 800 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_574_6
timestamp 1730953945
transform 1 0 800 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_591_6
timestamp 1730953945
transform 1 0 952 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_591_6
timestamp 1730953945
transform 1 0 952 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_590_6
timestamp 1730953945
transform 1 0 1080 0 1 736
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_590_6
timestamp 1730953945
transform 1 0 1080 0 1 736
box 7 3 85 69
use welltap_svt  __well_tap__17
timestamp 1730953945
transform 1 0 1176 0 1 756
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730953945
transform 1 0 1176 0 1 756
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730953945
transform 1 0 104 0 -1 860
box 8 4 12 24
use welltap_svt  __well_tap__18
timestamp 1730953945
transform 1 0 104 0 -1 860
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_545_6
timestamp 1730953945
transform 1 0 384 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_545_6
timestamp 1730953945
transform 1 0 384 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_546_6
timestamp 1730953945
transform 1 0 496 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_546_6
timestamp 1730953945
transform 1 0 496 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_547_6
timestamp 1730953945
transform 1 0 624 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_547_6
timestamp 1730953945
transform 1 0 624 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_548_6
timestamp 1730953945
transform 1 0 760 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_548_6
timestamp 1730953945
transform 1 0 760 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_573_6
timestamp 1730953945
transform 1 0 896 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_573_6
timestamp 1730953945
transform 1 0 896 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_592_6
timestamp 1730953945
transform 1 0 1040 0 -1 880
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_592_6
timestamp 1730953945
transform 1 0 1040 0 -1 880
box 7 3 85 69
use welltap_svt  __well_tap__19
timestamp 1730953945
transform 1 0 1176 0 -1 860
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730953945
transform 1 0 1176 0 -1 860
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_551_6
timestamp 1730953945
transform 1 0 312 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_551_6
timestamp 1730953945
transform 1 0 312 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_552_6
timestamp 1730953945
transform 1 0 424 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_552_6
timestamp 1730953945
transform 1 0 424 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_550_6
timestamp 1730953945
transform 1 0 544 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_550_6
timestamp 1730953945
transform 1 0 544 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_549_6
timestamp 1730953945
transform 1 0 672 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_549_6
timestamp 1730953945
transform 1 0 672 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_572_6
timestamp 1730953945
transform 1 0 800 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_572_6
timestamp 1730953945
transform 1 0 800 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_594_6
timestamp 1730953945
transform 1 0 936 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_594_6
timestamp 1730953945
transform 1 0 936 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_593_6
timestamp 1730953945
transform 1 0 1072 0 1 888
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_593_6
timestamp 1730953945
transform 1 0 1072 0 1 888
box 7 3 85 69
use welltap_svt  __well_tap__20
timestamp 1730953945
transform 1 0 104 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__20
timestamp 1730953945
transform 1 0 104 0 1 908
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_555_6
timestamp 1730953945
transform 1 0 224 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_555_6
timestamp 1730953945
transform 1 0 224 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_554_6
timestamp 1730953945
transform 1 0 376 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_554_6
timestamp 1730953945
transform 1 0 376 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_553_6
timestamp 1730953945
transform 1 0 528 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_553_6
timestamp 1730953945
transform 1 0 528 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_570_6
timestamp 1730953945
transform 1 0 688 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_570_6
timestamp 1730953945
transform 1 0 688 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_571_6
timestamp 1730953945
transform 1 0 856 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_571_6
timestamp 1730953945
transform 1 0 856 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_595_6
timestamp 1730953945
transform 1 0 1024 0 -1 1040
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_595_6
timestamp 1730953945
transform 1 0 1024 0 -1 1040
box 7 3 85 69
use welltap_svt  __well_tap__21
timestamp 1730953945
transform 1 0 1176 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730953945
transform 1 0 1176 0 1 908
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730953945
transform 1 0 104 0 -1 1020
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730953945
transform 1 0 104 0 -1 1020
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_558_6
timestamp 1730953945
transform 1 0 200 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_558_6
timestamp 1730953945
transform 1 0 200 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_556_6
timestamp 1730953945
transform 1 0 344 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_556_6
timestamp 1730953945
transform 1 0 344 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_557_6
timestamp 1730953945
transform 1 0 488 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_557_6
timestamp 1730953945
transform 1 0 488 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_569_6
timestamp 1730953945
transform 1 0 632 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_569_6
timestamp 1730953945
transform 1 0 632 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_568_6
timestamp 1730953945
transform 1 0 784 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_568_6
timestamp 1730953945
transform 1 0 784 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_597_6
timestamp 1730953945
transform 1 0 936 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_597_6
timestamp 1730953945
transform 1 0 936 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_596_6
timestamp 1730953945
transform 1 0 1080 0 1 1048
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_596_6
timestamp 1730953945
transform 1 0 1080 0 1 1048
box 7 3 85 69
use welltap_svt  __well_tap__23
timestamp 1730953945
transform 1 0 1176 0 -1 1020
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730953945
transform 1 0 1176 0 -1 1020
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730953945
transform 1 0 104 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730953945
transform 1 0 104 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730953945
transform 1 0 1176 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730953945
transform 1 0 1176 0 1 1068
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730953945
transform 1 0 104 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730953945
transform 1 0 104 0 -1 1188
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_559_6
timestamp 1730953945
transform 1 0 200 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_559_6
timestamp 1730953945
transform 1 0 200 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_560_6
timestamp 1730953945
transform 1 0 288 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_560_6
timestamp 1730953945
transform 1 0 288 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_561_6
timestamp 1730953945
transform 1 0 376 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_561_6
timestamp 1730953945
transform 1 0 376 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_562_6
timestamp 1730953945
transform 1 0 464 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_562_6
timestamp 1730953945
transform 1 0 464 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_563_6
timestamp 1730953945
transform 1 0 552 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_563_6
timestamp 1730953945
transform 1 0 552 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_565_6
timestamp 1730953945
transform 1 0 648 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_565_6
timestamp 1730953945
transform 1 0 648 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_566_6
timestamp 1730953945
transform 1 0 752 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_566_6
timestamp 1730953945
transform 1 0 752 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_567_6
timestamp 1730953945
transform 1 0 864 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_567_6
timestamp 1730953945
transform 1 0 864 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_598_6
timestamp 1730953945
transform 1 0 984 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_598_6
timestamp 1730953945
transform 1 0 984 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_599_6
timestamp 1730953945
transform 1 0 1080 0 -1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_599_6
timestamp 1730953945
transform 1 0 1080 0 -1 1208
box 7 3 85 69
use welltap_svt  __well_tap__27
timestamp 1730953945
transform 1 0 1176 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730953945
transform 1 0 1176 0 -1 1188
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730953945
transform 1 0 104 0 1 1228
box 8 4 12 24
use welltap_svt  __well_tap__28
timestamp 1730953945
transform 1 0 104 0 1 1228
box 8 4 12 24
use _0_0std_0_0cells_0_0LATCH  latch_564_6
timestamp 1730953945
transform 1 0 560 0 1 1208
box 7 3 85 69
use _0_0std_0_0cells_0_0LATCH  latch_564_6
timestamp 1730953945
transform 1 0 560 0 1 1208
box 7 3 85 69
use welltap_svt  __well_tap__29
timestamp 1730953945
transform 1 0 1176 0 1 1228
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730953945
transform 1 0 1176 0 1 1228
box 8 4 12 24
<< end >>
