magic
tech TSMC180
timestamp 1734143631
<< m1 >>
rect 6 97 9 100
rect 18 97 21 100
rect 30 97 33 100
rect 6 18 29 91
rect 6 10 9 13
<< labels >>
rlabel m1 s 6 97 9 100 6 in_50_6
port 1 nsew signal input
rlabel m1 s 6 10 9 13 6 out
port 2 nsew signal output
rlabel m1 s 18 97 21 100 6 Vdd
port 3 nsew power input
rlabel m1 s 30 97 33 100 6 GND
port 4 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 36 110
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
