magic
tech sky130l
timestamp 1731220321
<< m2 >>
rect 1806 3500 1812 3501
rect 3462 3500 3468 3501
rect 1806 3496 1807 3500
rect 1811 3496 1812 3500
rect 1806 3495 1812 3496
rect 2006 3499 2012 3500
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 2238 3499 2244 3500
rect 2238 3495 2239 3499
rect 2243 3495 2244 3499
rect 2238 3494 2244 3495
rect 2454 3499 2460 3500
rect 2454 3495 2455 3499
rect 2459 3495 2460 3499
rect 2454 3494 2460 3495
rect 2654 3499 2660 3500
rect 2654 3495 2655 3499
rect 2659 3495 2660 3499
rect 2654 3494 2660 3495
rect 2854 3499 2860 3500
rect 2854 3495 2855 3499
rect 2859 3495 2860 3499
rect 2854 3494 2860 3495
rect 3046 3499 3052 3500
rect 3046 3495 3047 3499
rect 3051 3495 3052 3499
rect 3046 3494 3052 3495
rect 3246 3499 3252 3500
rect 3246 3495 3247 3499
rect 3251 3495 3252 3499
rect 3462 3496 3463 3500
rect 3467 3496 3468 3500
rect 3462 3495 3468 3496
rect 3246 3494 3252 3495
rect 1806 3483 1812 3484
rect 1806 3479 1807 3483
rect 1811 3479 1812 3483
rect 3462 3483 3468 3484
rect 1806 3478 1812 3479
rect 2006 3480 2012 3481
rect 2006 3476 2007 3480
rect 2011 3476 2012 3480
rect 2006 3475 2012 3476
rect 2238 3480 2244 3481
rect 2238 3476 2239 3480
rect 2243 3476 2244 3480
rect 2238 3475 2244 3476
rect 2454 3480 2460 3481
rect 2454 3476 2455 3480
rect 2459 3476 2460 3480
rect 2454 3475 2460 3476
rect 2654 3480 2660 3481
rect 2654 3476 2655 3480
rect 2659 3476 2660 3480
rect 2654 3475 2660 3476
rect 2854 3480 2860 3481
rect 2854 3476 2855 3480
rect 2859 3476 2860 3480
rect 2854 3475 2860 3476
rect 3046 3480 3052 3481
rect 3046 3476 3047 3480
rect 3051 3476 3052 3480
rect 3046 3475 3052 3476
rect 3246 3480 3252 3481
rect 3246 3476 3247 3480
rect 3251 3476 3252 3480
rect 3462 3479 3463 3483
rect 3467 3479 3468 3483
rect 3462 3478 3468 3479
rect 3246 3475 3252 3476
rect 110 3464 116 3465
rect 1766 3464 1772 3465
rect 110 3460 111 3464
rect 115 3460 116 3464
rect 110 3459 116 3460
rect 454 3463 460 3464
rect 454 3459 455 3463
rect 459 3459 460 3463
rect 454 3458 460 3459
rect 542 3463 548 3464
rect 542 3459 543 3463
rect 547 3459 548 3463
rect 542 3458 548 3459
rect 630 3463 636 3464
rect 630 3459 631 3463
rect 635 3459 636 3463
rect 630 3458 636 3459
rect 718 3463 724 3464
rect 718 3459 719 3463
rect 723 3459 724 3463
rect 718 3458 724 3459
rect 806 3463 812 3464
rect 806 3459 807 3463
rect 811 3459 812 3463
rect 806 3458 812 3459
rect 894 3463 900 3464
rect 894 3459 895 3463
rect 899 3459 900 3463
rect 894 3458 900 3459
rect 982 3463 988 3464
rect 982 3459 983 3463
rect 987 3459 988 3463
rect 982 3458 988 3459
rect 1070 3463 1076 3464
rect 1070 3459 1071 3463
rect 1075 3459 1076 3463
rect 1070 3458 1076 3459
rect 1158 3463 1164 3464
rect 1158 3459 1159 3463
rect 1163 3459 1164 3463
rect 1766 3460 1767 3464
rect 1771 3460 1772 3464
rect 1766 3459 1772 3460
rect 1158 3458 1164 3459
rect 110 3447 116 3448
rect 110 3443 111 3447
rect 115 3443 116 3447
rect 1766 3447 1772 3448
rect 110 3442 116 3443
rect 454 3444 460 3445
rect 454 3440 455 3444
rect 459 3440 460 3444
rect 454 3439 460 3440
rect 542 3444 548 3445
rect 542 3440 543 3444
rect 547 3440 548 3444
rect 542 3439 548 3440
rect 630 3444 636 3445
rect 630 3440 631 3444
rect 635 3440 636 3444
rect 630 3439 636 3440
rect 718 3444 724 3445
rect 718 3440 719 3444
rect 723 3440 724 3444
rect 718 3439 724 3440
rect 806 3444 812 3445
rect 806 3440 807 3444
rect 811 3440 812 3444
rect 806 3439 812 3440
rect 894 3444 900 3445
rect 894 3440 895 3444
rect 899 3440 900 3444
rect 894 3439 900 3440
rect 982 3444 988 3445
rect 982 3440 983 3444
rect 987 3440 988 3444
rect 982 3439 988 3440
rect 1070 3444 1076 3445
rect 1070 3440 1071 3444
rect 1075 3440 1076 3444
rect 1070 3439 1076 3440
rect 1158 3444 1164 3445
rect 1158 3440 1159 3444
rect 1163 3440 1164 3444
rect 1766 3443 1767 3447
rect 1771 3443 1772 3447
rect 1766 3442 1772 3443
rect 1158 3439 1164 3440
rect 1830 3436 1836 3437
rect 1806 3433 1812 3434
rect 1806 3429 1807 3433
rect 1811 3429 1812 3433
rect 1830 3432 1831 3436
rect 1835 3432 1836 3436
rect 1830 3431 1836 3432
rect 1942 3436 1948 3437
rect 1942 3432 1943 3436
rect 1947 3432 1948 3436
rect 1942 3431 1948 3432
rect 2078 3436 2084 3437
rect 2078 3432 2079 3436
rect 2083 3432 2084 3436
rect 2078 3431 2084 3432
rect 2214 3436 2220 3437
rect 2214 3432 2215 3436
rect 2219 3432 2220 3436
rect 2214 3431 2220 3432
rect 2350 3436 2356 3437
rect 2350 3432 2351 3436
rect 2355 3432 2356 3436
rect 2350 3431 2356 3432
rect 2478 3436 2484 3437
rect 2478 3432 2479 3436
rect 2483 3432 2484 3436
rect 2478 3431 2484 3432
rect 2598 3436 2604 3437
rect 2598 3432 2599 3436
rect 2603 3432 2604 3436
rect 2598 3431 2604 3432
rect 2718 3436 2724 3437
rect 2718 3432 2719 3436
rect 2723 3432 2724 3436
rect 2718 3431 2724 3432
rect 2846 3436 2852 3437
rect 2846 3432 2847 3436
rect 2851 3432 2852 3436
rect 2846 3431 2852 3432
rect 2974 3436 2980 3437
rect 2974 3432 2975 3436
rect 2979 3432 2980 3436
rect 2974 3431 2980 3432
rect 3462 3433 3468 3434
rect 1806 3428 1812 3429
rect 3462 3429 3463 3433
rect 3467 3429 3468 3433
rect 3462 3428 3468 3429
rect 1830 3417 1836 3418
rect 1806 3416 1812 3417
rect 1806 3412 1807 3416
rect 1811 3412 1812 3416
rect 1830 3413 1831 3417
rect 1835 3413 1836 3417
rect 1830 3412 1836 3413
rect 1942 3417 1948 3418
rect 1942 3413 1943 3417
rect 1947 3413 1948 3417
rect 1942 3412 1948 3413
rect 2078 3417 2084 3418
rect 2078 3413 2079 3417
rect 2083 3413 2084 3417
rect 2078 3412 2084 3413
rect 2214 3417 2220 3418
rect 2214 3413 2215 3417
rect 2219 3413 2220 3417
rect 2214 3412 2220 3413
rect 2350 3417 2356 3418
rect 2350 3413 2351 3417
rect 2355 3413 2356 3417
rect 2350 3412 2356 3413
rect 2478 3417 2484 3418
rect 2478 3413 2479 3417
rect 2483 3413 2484 3417
rect 2478 3412 2484 3413
rect 2598 3417 2604 3418
rect 2598 3413 2599 3417
rect 2603 3413 2604 3417
rect 2598 3412 2604 3413
rect 2718 3417 2724 3418
rect 2718 3413 2719 3417
rect 2723 3413 2724 3417
rect 2718 3412 2724 3413
rect 2846 3417 2852 3418
rect 2846 3413 2847 3417
rect 2851 3413 2852 3417
rect 2846 3412 2852 3413
rect 2974 3417 2980 3418
rect 2974 3413 2975 3417
rect 2979 3413 2980 3417
rect 2974 3412 2980 3413
rect 3462 3416 3468 3417
rect 3462 3412 3463 3416
rect 3467 3412 3468 3416
rect 1806 3411 1812 3412
rect 3462 3411 3468 3412
rect 414 3400 420 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 414 3396 415 3400
rect 419 3396 420 3400
rect 414 3395 420 3396
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 590 3400 596 3401
rect 590 3396 591 3400
rect 595 3396 596 3400
rect 590 3395 596 3396
rect 678 3400 684 3401
rect 678 3396 679 3400
rect 683 3396 684 3400
rect 678 3395 684 3396
rect 766 3400 772 3401
rect 766 3396 767 3400
rect 771 3396 772 3400
rect 766 3395 772 3396
rect 854 3400 860 3401
rect 854 3396 855 3400
rect 859 3396 860 3400
rect 854 3395 860 3396
rect 942 3400 948 3401
rect 942 3396 943 3400
rect 947 3396 948 3400
rect 942 3395 948 3396
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 1118 3400 1124 3401
rect 1118 3396 1119 3400
rect 1123 3396 1124 3400
rect 1118 3395 1124 3396
rect 1206 3400 1212 3401
rect 1206 3396 1207 3400
rect 1211 3396 1212 3400
rect 1206 3395 1212 3396
rect 1302 3400 1308 3401
rect 1302 3396 1303 3400
rect 1307 3396 1308 3400
rect 1302 3395 1308 3396
rect 1766 3397 1772 3398
rect 110 3392 116 3393
rect 1766 3393 1767 3397
rect 1771 3393 1772 3397
rect 1766 3392 1772 3393
rect 414 3381 420 3382
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 414 3377 415 3381
rect 419 3377 420 3381
rect 414 3376 420 3377
rect 502 3381 508 3382
rect 502 3377 503 3381
rect 507 3377 508 3381
rect 502 3376 508 3377
rect 590 3381 596 3382
rect 590 3377 591 3381
rect 595 3377 596 3381
rect 590 3376 596 3377
rect 678 3381 684 3382
rect 678 3377 679 3381
rect 683 3377 684 3381
rect 678 3376 684 3377
rect 766 3381 772 3382
rect 766 3377 767 3381
rect 771 3377 772 3381
rect 766 3376 772 3377
rect 854 3381 860 3382
rect 854 3377 855 3381
rect 859 3377 860 3381
rect 854 3376 860 3377
rect 942 3381 948 3382
rect 942 3377 943 3381
rect 947 3377 948 3381
rect 942 3376 948 3377
rect 1030 3381 1036 3382
rect 1030 3377 1031 3381
rect 1035 3377 1036 3381
rect 1030 3376 1036 3377
rect 1118 3381 1124 3382
rect 1118 3377 1119 3381
rect 1123 3377 1124 3381
rect 1118 3376 1124 3377
rect 1206 3381 1212 3382
rect 1206 3377 1207 3381
rect 1211 3377 1212 3381
rect 1206 3376 1212 3377
rect 1302 3381 1308 3382
rect 1302 3377 1303 3381
rect 1307 3377 1308 3381
rect 1302 3376 1308 3377
rect 1766 3380 1772 3381
rect 1766 3376 1767 3380
rect 1771 3376 1772 3380
rect 110 3375 116 3376
rect 1766 3375 1772 3376
rect 1806 3364 1812 3365
rect 3462 3364 3468 3365
rect 1806 3360 1807 3364
rect 1811 3360 1812 3364
rect 1806 3359 1812 3360
rect 1830 3363 1836 3364
rect 1830 3359 1831 3363
rect 1835 3359 1836 3363
rect 1830 3358 1836 3359
rect 1950 3363 1956 3364
rect 1950 3359 1951 3363
rect 1955 3359 1956 3363
rect 1950 3358 1956 3359
rect 2094 3363 2100 3364
rect 2094 3359 2095 3363
rect 2099 3359 2100 3363
rect 2094 3358 2100 3359
rect 2238 3363 2244 3364
rect 2238 3359 2239 3363
rect 2243 3359 2244 3363
rect 2238 3358 2244 3359
rect 2382 3363 2388 3364
rect 2382 3359 2383 3363
rect 2387 3359 2388 3363
rect 2382 3358 2388 3359
rect 2518 3363 2524 3364
rect 2518 3359 2519 3363
rect 2523 3359 2524 3363
rect 2518 3358 2524 3359
rect 2646 3363 2652 3364
rect 2646 3359 2647 3363
rect 2651 3359 2652 3363
rect 2646 3358 2652 3359
rect 2774 3363 2780 3364
rect 2774 3359 2775 3363
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2902 3363 2908 3364
rect 2902 3359 2903 3363
rect 2907 3359 2908 3363
rect 2902 3358 2908 3359
rect 3038 3363 3044 3364
rect 3038 3359 3039 3363
rect 3043 3359 3044 3363
rect 3462 3360 3463 3364
rect 3467 3360 3468 3364
rect 3462 3359 3468 3360
rect 3038 3358 3044 3359
rect 1806 3347 1812 3348
rect 1806 3343 1807 3347
rect 1811 3343 1812 3347
rect 3462 3347 3468 3348
rect 1806 3342 1812 3343
rect 1830 3344 1836 3345
rect 1830 3340 1831 3344
rect 1835 3340 1836 3344
rect 1830 3339 1836 3340
rect 1950 3344 1956 3345
rect 1950 3340 1951 3344
rect 1955 3340 1956 3344
rect 1950 3339 1956 3340
rect 2094 3344 2100 3345
rect 2094 3340 2095 3344
rect 2099 3340 2100 3344
rect 2094 3339 2100 3340
rect 2238 3344 2244 3345
rect 2238 3340 2239 3344
rect 2243 3340 2244 3344
rect 2238 3339 2244 3340
rect 2382 3344 2388 3345
rect 2382 3340 2383 3344
rect 2387 3340 2388 3344
rect 2382 3339 2388 3340
rect 2518 3344 2524 3345
rect 2518 3340 2519 3344
rect 2523 3340 2524 3344
rect 2518 3339 2524 3340
rect 2646 3344 2652 3345
rect 2646 3340 2647 3344
rect 2651 3340 2652 3344
rect 2646 3339 2652 3340
rect 2774 3344 2780 3345
rect 2774 3340 2775 3344
rect 2779 3340 2780 3344
rect 2774 3339 2780 3340
rect 2902 3344 2908 3345
rect 2902 3340 2903 3344
rect 2907 3340 2908 3344
rect 2902 3339 2908 3340
rect 3038 3344 3044 3345
rect 3038 3340 3039 3344
rect 3043 3340 3044 3344
rect 3462 3343 3463 3347
rect 3467 3343 3468 3347
rect 3462 3342 3468 3343
rect 3038 3339 3044 3340
rect 110 3332 116 3333
rect 1766 3332 1772 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 398 3331 404 3332
rect 398 3327 399 3331
rect 403 3327 404 3331
rect 398 3326 404 3327
rect 494 3331 500 3332
rect 494 3327 495 3331
rect 499 3327 500 3331
rect 494 3326 500 3327
rect 598 3331 604 3332
rect 598 3327 599 3331
rect 603 3327 604 3331
rect 598 3326 604 3327
rect 702 3331 708 3332
rect 702 3327 703 3331
rect 707 3327 708 3331
rect 702 3326 708 3327
rect 806 3331 812 3332
rect 806 3327 807 3331
rect 811 3327 812 3331
rect 806 3326 812 3327
rect 910 3331 916 3332
rect 910 3327 911 3331
rect 915 3327 916 3331
rect 910 3326 916 3327
rect 1014 3331 1020 3332
rect 1014 3327 1015 3331
rect 1019 3327 1020 3331
rect 1014 3326 1020 3327
rect 1118 3331 1124 3332
rect 1118 3327 1119 3331
rect 1123 3327 1124 3331
rect 1118 3326 1124 3327
rect 1222 3331 1228 3332
rect 1222 3327 1223 3331
rect 1227 3327 1228 3331
rect 1222 3326 1228 3327
rect 1326 3331 1332 3332
rect 1326 3327 1327 3331
rect 1331 3327 1332 3331
rect 1766 3328 1767 3332
rect 1771 3328 1772 3332
rect 1766 3327 1772 3328
rect 1326 3326 1332 3327
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 1766 3315 1772 3316
rect 110 3310 116 3311
rect 398 3312 404 3313
rect 398 3308 399 3312
rect 403 3308 404 3312
rect 398 3307 404 3308
rect 494 3312 500 3313
rect 494 3308 495 3312
rect 499 3308 500 3312
rect 494 3307 500 3308
rect 598 3312 604 3313
rect 598 3308 599 3312
rect 603 3308 604 3312
rect 598 3307 604 3308
rect 702 3312 708 3313
rect 702 3308 703 3312
rect 707 3308 708 3312
rect 702 3307 708 3308
rect 806 3312 812 3313
rect 806 3308 807 3312
rect 811 3308 812 3312
rect 806 3307 812 3308
rect 910 3312 916 3313
rect 910 3308 911 3312
rect 915 3308 916 3312
rect 910 3307 916 3308
rect 1014 3312 1020 3313
rect 1014 3308 1015 3312
rect 1019 3308 1020 3312
rect 1014 3307 1020 3308
rect 1118 3312 1124 3313
rect 1118 3308 1119 3312
rect 1123 3308 1124 3312
rect 1118 3307 1124 3308
rect 1222 3312 1228 3313
rect 1222 3308 1223 3312
rect 1227 3308 1228 3312
rect 1222 3307 1228 3308
rect 1326 3312 1332 3313
rect 1326 3308 1327 3312
rect 1331 3308 1332 3312
rect 1766 3311 1767 3315
rect 1771 3311 1772 3315
rect 1766 3310 1772 3311
rect 1326 3307 1332 3308
rect 1830 3292 1836 3293
rect 1806 3289 1812 3290
rect 1806 3285 1807 3289
rect 1811 3285 1812 3289
rect 1830 3288 1831 3292
rect 1835 3288 1836 3292
rect 1830 3287 1836 3288
rect 1974 3292 1980 3293
rect 1974 3288 1975 3292
rect 1979 3288 1980 3292
rect 1974 3287 1980 3288
rect 2150 3292 2156 3293
rect 2150 3288 2151 3292
rect 2155 3288 2156 3292
rect 2150 3287 2156 3288
rect 2334 3292 2340 3293
rect 2334 3288 2335 3292
rect 2339 3288 2340 3292
rect 2334 3287 2340 3288
rect 2510 3292 2516 3293
rect 2510 3288 2511 3292
rect 2515 3288 2516 3292
rect 2510 3287 2516 3288
rect 2678 3292 2684 3293
rect 2678 3288 2679 3292
rect 2683 3288 2684 3292
rect 2678 3287 2684 3288
rect 2830 3292 2836 3293
rect 2830 3288 2831 3292
rect 2835 3288 2836 3292
rect 2830 3287 2836 3288
rect 2974 3292 2980 3293
rect 2974 3288 2975 3292
rect 2979 3288 2980 3292
rect 2974 3287 2980 3288
rect 3110 3292 3116 3293
rect 3110 3288 3111 3292
rect 3115 3288 3116 3292
rect 3110 3287 3116 3288
rect 3246 3292 3252 3293
rect 3246 3288 3247 3292
rect 3251 3288 3252 3292
rect 3246 3287 3252 3288
rect 3366 3292 3372 3293
rect 3366 3288 3367 3292
rect 3371 3288 3372 3292
rect 3366 3287 3372 3288
rect 3462 3289 3468 3290
rect 1806 3284 1812 3285
rect 3462 3285 3463 3289
rect 3467 3285 3468 3289
rect 3462 3284 3468 3285
rect 1830 3273 1836 3274
rect 1806 3272 1812 3273
rect 1806 3268 1807 3272
rect 1811 3268 1812 3272
rect 1830 3269 1831 3273
rect 1835 3269 1836 3273
rect 1830 3268 1836 3269
rect 1974 3273 1980 3274
rect 1974 3269 1975 3273
rect 1979 3269 1980 3273
rect 1974 3268 1980 3269
rect 2150 3273 2156 3274
rect 2150 3269 2151 3273
rect 2155 3269 2156 3273
rect 2150 3268 2156 3269
rect 2334 3273 2340 3274
rect 2334 3269 2335 3273
rect 2339 3269 2340 3273
rect 2334 3268 2340 3269
rect 2510 3273 2516 3274
rect 2510 3269 2511 3273
rect 2515 3269 2516 3273
rect 2510 3268 2516 3269
rect 2678 3273 2684 3274
rect 2678 3269 2679 3273
rect 2683 3269 2684 3273
rect 2678 3268 2684 3269
rect 2830 3273 2836 3274
rect 2830 3269 2831 3273
rect 2835 3269 2836 3273
rect 2830 3268 2836 3269
rect 2974 3273 2980 3274
rect 2974 3269 2975 3273
rect 2979 3269 2980 3273
rect 2974 3268 2980 3269
rect 3110 3273 3116 3274
rect 3110 3269 3111 3273
rect 3115 3269 3116 3273
rect 3110 3268 3116 3269
rect 3246 3273 3252 3274
rect 3246 3269 3247 3273
rect 3251 3269 3252 3273
rect 3246 3268 3252 3269
rect 3366 3273 3372 3274
rect 3366 3269 3367 3273
rect 3371 3269 3372 3273
rect 3366 3268 3372 3269
rect 3462 3272 3468 3273
rect 3462 3268 3463 3272
rect 3467 3268 3468 3272
rect 1806 3267 1812 3268
rect 3462 3267 3468 3268
rect 382 3264 388 3265
rect 110 3261 116 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 382 3260 383 3264
rect 387 3260 388 3264
rect 382 3259 388 3260
rect 494 3264 500 3265
rect 494 3260 495 3264
rect 499 3260 500 3264
rect 494 3259 500 3260
rect 606 3264 612 3265
rect 606 3260 607 3264
rect 611 3260 612 3264
rect 606 3259 612 3260
rect 726 3264 732 3265
rect 726 3260 727 3264
rect 731 3260 732 3264
rect 726 3259 732 3260
rect 846 3264 852 3265
rect 846 3260 847 3264
rect 851 3260 852 3264
rect 846 3259 852 3260
rect 966 3264 972 3265
rect 966 3260 967 3264
rect 971 3260 972 3264
rect 966 3259 972 3260
rect 1086 3264 1092 3265
rect 1086 3260 1087 3264
rect 1091 3260 1092 3264
rect 1086 3259 1092 3260
rect 1206 3264 1212 3265
rect 1206 3260 1207 3264
rect 1211 3260 1212 3264
rect 1206 3259 1212 3260
rect 1334 3264 1340 3265
rect 1334 3260 1335 3264
rect 1339 3260 1340 3264
rect 1334 3259 1340 3260
rect 1766 3261 1772 3262
rect 110 3256 116 3257
rect 1766 3257 1767 3261
rect 1771 3257 1772 3261
rect 1766 3256 1772 3257
rect 382 3245 388 3246
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 382 3241 383 3245
rect 387 3241 388 3245
rect 382 3240 388 3241
rect 494 3245 500 3246
rect 494 3241 495 3245
rect 499 3241 500 3245
rect 494 3240 500 3241
rect 606 3245 612 3246
rect 606 3241 607 3245
rect 611 3241 612 3245
rect 606 3240 612 3241
rect 726 3245 732 3246
rect 726 3241 727 3245
rect 731 3241 732 3245
rect 726 3240 732 3241
rect 846 3245 852 3246
rect 846 3241 847 3245
rect 851 3241 852 3245
rect 846 3240 852 3241
rect 966 3245 972 3246
rect 966 3241 967 3245
rect 971 3241 972 3245
rect 966 3240 972 3241
rect 1086 3245 1092 3246
rect 1086 3241 1087 3245
rect 1091 3241 1092 3245
rect 1086 3240 1092 3241
rect 1206 3245 1212 3246
rect 1206 3241 1207 3245
rect 1211 3241 1212 3245
rect 1206 3240 1212 3241
rect 1334 3245 1340 3246
rect 1334 3241 1335 3245
rect 1339 3241 1340 3245
rect 1334 3240 1340 3241
rect 1766 3244 1772 3245
rect 1766 3240 1767 3244
rect 1771 3240 1772 3244
rect 110 3239 116 3240
rect 1766 3239 1772 3240
rect 1806 3220 1812 3221
rect 3462 3220 3468 3221
rect 1806 3216 1807 3220
rect 1811 3216 1812 3220
rect 1806 3215 1812 3216
rect 1830 3219 1836 3220
rect 1830 3215 1831 3219
rect 1835 3215 1836 3219
rect 1830 3214 1836 3215
rect 2030 3219 2036 3220
rect 2030 3215 2031 3219
rect 2035 3215 2036 3219
rect 2030 3214 2036 3215
rect 2246 3219 2252 3220
rect 2246 3215 2247 3219
rect 2251 3215 2252 3219
rect 2246 3214 2252 3215
rect 2454 3219 2460 3220
rect 2454 3215 2455 3219
rect 2459 3215 2460 3219
rect 2454 3214 2460 3215
rect 2654 3219 2660 3220
rect 2654 3215 2655 3219
rect 2659 3215 2660 3219
rect 2654 3214 2660 3215
rect 2838 3219 2844 3220
rect 2838 3215 2839 3219
rect 2843 3215 2844 3219
rect 2838 3214 2844 3215
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3215 3028 3219
rect 3022 3214 3028 3215
rect 3206 3219 3212 3220
rect 3206 3215 3207 3219
rect 3211 3215 3212 3219
rect 3206 3214 3212 3215
rect 3366 3219 3372 3220
rect 3366 3215 3367 3219
rect 3371 3215 3372 3219
rect 3462 3216 3463 3220
rect 3467 3216 3468 3220
rect 3462 3215 3468 3216
rect 3366 3214 3372 3215
rect 1806 3203 1812 3204
rect 1806 3199 1807 3203
rect 1811 3199 1812 3203
rect 3462 3203 3468 3204
rect 1806 3198 1812 3199
rect 1830 3200 1836 3201
rect 110 3196 116 3197
rect 1766 3196 1772 3197
rect 110 3192 111 3196
rect 115 3192 116 3196
rect 110 3191 116 3192
rect 302 3195 308 3196
rect 302 3191 303 3195
rect 307 3191 308 3195
rect 302 3190 308 3191
rect 422 3195 428 3196
rect 422 3191 423 3195
rect 427 3191 428 3195
rect 422 3190 428 3191
rect 542 3195 548 3196
rect 542 3191 543 3195
rect 547 3191 548 3195
rect 542 3190 548 3191
rect 670 3195 676 3196
rect 670 3191 671 3195
rect 675 3191 676 3195
rect 670 3190 676 3191
rect 798 3195 804 3196
rect 798 3191 799 3195
rect 803 3191 804 3195
rect 798 3190 804 3191
rect 926 3195 932 3196
rect 926 3191 927 3195
rect 931 3191 932 3195
rect 926 3190 932 3191
rect 1054 3195 1060 3196
rect 1054 3191 1055 3195
rect 1059 3191 1060 3195
rect 1054 3190 1060 3191
rect 1174 3195 1180 3196
rect 1174 3191 1175 3195
rect 1179 3191 1180 3195
rect 1174 3190 1180 3191
rect 1302 3195 1308 3196
rect 1302 3191 1303 3195
rect 1307 3191 1308 3195
rect 1302 3190 1308 3191
rect 1430 3195 1436 3196
rect 1430 3191 1431 3195
rect 1435 3191 1436 3195
rect 1766 3192 1767 3196
rect 1771 3192 1772 3196
rect 1830 3196 1831 3200
rect 1835 3196 1836 3200
rect 1830 3195 1836 3196
rect 2030 3200 2036 3201
rect 2030 3196 2031 3200
rect 2035 3196 2036 3200
rect 2030 3195 2036 3196
rect 2246 3200 2252 3201
rect 2246 3196 2247 3200
rect 2251 3196 2252 3200
rect 2246 3195 2252 3196
rect 2454 3200 2460 3201
rect 2454 3196 2455 3200
rect 2459 3196 2460 3200
rect 2454 3195 2460 3196
rect 2654 3200 2660 3201
rect 2654 3196 2655 3200
rect 2659 3196 2660 3200
rect 2654 3195 2660 3196
rect 2838 3200 2844 3201
rect 2838 3196 2839 3200
rect 2843 3196 2844 3200
rect 2838 3195 2844 3196
rect 3022 3200 3028 3201
rect 3022 3196 3023 3200
rect 3027 3196 3028 3200
rect 3022 3195 3028 3196
rect 3206 3200 3212 3201
rect 3206 3196 3207 3200
rect 3211 3196 3212 3200
rect 3206 3195 3212 3196
rect 3366 3200 3372 3201
rect 3366 3196 3367 3200
rect 3371 3196 3372 3200
rect 3462 3199 3463 3203
rect 3467 3199 3468 3203
rect 3462 3198 3468 3199
rect 3366 3195 3372 3196
rect 1766 3191 1772 3192
rect 1430 3190 1436 3191
rect 110 3179 116 3180
rect 110 3175 111 3179
rect 115 3175 116 3179
rect 1766 3179 1772 3180
rect 110 3174 116 3175
rect 302 3176 308 3177
rect 302 3172 303 3176
rect 307 3172 308 3176
rect 302 3171 308 3172
rect 422 3176 428 3177
rect 422 3172 423 3176
rect 427 3172 428 3176
rect 422 3171 428 3172
rect 542 3176 548 3177
rect 542 3172 543 3176
rect 547 3172 548 3176
rect 542 3171 548 3172
rect 670 3176 676 3177
rect 670 3172 671 3176
rect 675 3172 676 3176
rect 670 3171 676 3172
rect 798 3176 804 3177
rect 798 3172 799 3176
rect 803 3172 804 3176
rect 798 3171 804 3172
rect 926 3176 932 3177
rect 926 3172 927 3176
rect 931 3172 932 3176
rect 926 3171 932 3172
rect 1054 3176 1060 3177
rect 1054 3172 1055 3176
rect 1059 3172 1060 3176
rect 1054 3171 1060 3172
rect 1174 3176 1180 3177
rect 1174 3172 1175 3176
rect 1179 3172 1180 3176
rect 1174 3171 1180 3172
rect 1302 3176 1308 3177
rect 1302 3172 1303 3176
rect 1307 3172 1308 3176
rect 1302 3171 1308 3172
rect 1430 3176 1436 3177
rect 1430 3172 1431 3176
rect 1435 3172 1436 3176
rect 1766 3175 1767 3179
rect 1771 3175 1772 3179
rect 1766 3174 1772 3175
rect 1430 3171 1436 3172
rect 1838 3156 1844 3157
rect 1806 3153 1812 3154
rect 1806 3149 1807 3153
rect 1811 3149 1812 3153
rect 1838 3152 1839 3156
rect 1843 3152 1844 3156
rect 1838 3151 1844 3152
rect 2030 3156 2036 3157
rect 2030 3152 2031 3156
rect 2035 3152 2036 3156
rect 2030 3151 2036 3152
rect 2222 3156 2228 3157
rect 2222 3152 2223 3156
rect 2227 3152 2228 3156
rect 2222 3151 2228 3152
rect 2406 3156 2412 3157
rect 2406 3152 2407 3156
rect 2411 3152 2412 3156
rect 2406 3151 2412 3152
rect 2574 3156 2580 3157
rect 2574 3152 2575 3156
rect 2579 3152 2580 3156
rect 2574 3151 2580 3152
rect 2734 3156 2740 3157
rect 2734 3152 2735 3156
rect 2739 3152 2740 3156
rect 2734 3151 2740 3152
rect 2878 3156 2884 3157
rect 2878 3152 2879 3156
rect 2883 3152 2884 3156
rect 2878 3151 2884 3152
rect 3006 3156 3012 3157
rect 3006 3152 3007 3156
rect 3011 3152 3012 3156
rect 3006 3151 3012 3152
rect 3134 3156 3140 3157
rect 3134 3152 3135 3156
rect 3139 3152 3140 3156
rect 3134 3151 3140 3152
rect 3262 3156 3268 3157
rect 3262 3152 3263 3156
rect 3267 3152 3268 3156
rect 3262 3151 3268 3152
rect 3366 3156 3372 3157
rect 3366 3152 3367 3156
rect 3371 3152 3372 3156
rect 3366 3151 3372 3152
rect 3462 3153 3468 3154
rect 1806 3148 1812 3149
rect 3462 3149 3463 3153
rect 3467 3149 3468 3153
rect 3462 3148 3468 3149
rect 1838 3137 1844 3138
rect 1806 3136 1812 3137
rect 1806 3132 1807 3136
rect 1811 3132 1812 3136
rect 1838 3133 1839 3137
rect 1843 3133 1844 3137
rect 1838 3132 1844 3133
rect 2030 3137 2036 3138
rect 2030 3133 2031 3137
rect 2035 3133 2036 3137
rect 2030 3132 2036 3133
rect 2222 3137 2228 3138
rect 2222 3133 2223 3137
rect 2227 3133 2228 3137
rect 2222 3132 2228 3133
rect 2406 3137 2412 3138
rect 2406 3133 2407 3137
rect 2411 3133 2412 3137
rect 2406 3132 2412 3133
rect 2574 3137 2580 3138
rect 2574 3133 2575 3137
rect 2579 3133 2580 3137
rect 2574 3132 2580 3133
rect 2734 3137 2740 3138
rect 2734 3133 2735 3137
rect 2739 3133 2740 3137
rect 2734 3132 2740 3133
rect 2878 3137 2884 3138
rect 2878 3133 2879 3137
rect 2883 3133 2884 3137
rect 2878 3132 2884 3133
rect 3006 3137 3012 3138
rect 3006 3133 3007 3137
rect 3011 3133 3012 3137
rect 3006 3132 3012 3133
rect 3134 3137 3140 3138
rect 3134 3133 3135 3137
rect 3139 3133 3140 3137
rect 3134 3132 3140 3133
rect 3262 3137 3268 3138
rect 3262 3133 3263 3137
rect 3267 3133 3268 3137
rect 3262 3132 3268 3133
rect 3366 3137 3372 3138
rect 3366 3133 3367 3137
rect 3371 3133 3372 3137
rect 3366 3132 3372 3133
rect 3462 3136 3468 3137
rect 3462 3132 3463 3136
rect 3467 3132 3468 3136
rect 1806 3131 1812 3132
rect 3462 3131 3468 3132
rect 174 3120 180 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 174 3116 175 3120
rect 179 3116 180 3120
rect 174 3115 180 3116
rect 318 3120 324 3121
rect 318 3116 319 3120
rect 323 3116 324 3120
rect 318 3115 324 3116
rect 470 3120 476 3121
rect 470 3116 471 3120
rect 475 3116 476 3120
rect 470 3115 476 3116
rect 622 3120 628 3121
rect 622 3116 623 3120
rect 627 3116 628 3120
rect 622 3115 628 3116
rect 774 3120 780 3121
rect 774 3116 775 3120
rect 779 3116 780 3120
rect 774 3115 780 3116
rect 918 3120 924 3121
rect 918 3116 919 3120
rect 923 3116 924 3120
rect 918 3115 924 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1198 3120 1204 3121
rect 1198 3116 1199 3120
rect 1203 3116 1204 3120
rect 1198 3115 1204 3116
rect 1342 3120 1348 3121
rect 1342 3116 1343 3120
rect 1347 3116 1348 3120
rect 1342 3115 1348 3116
rect 1486 3120 1492 3121
rect 1486 3116 1487 3120
rect 1491 3116 1492 3120
rect 1486 3115 1492 3116
rect 1766 3117 1772 3118
rect 110 3112 116 3113
rect 1766 3113 1767 3117
rect 1771 3113 1772 3117
rect 1766 3112 1772 3113
rect 174 3101 180 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 174 3097 175 3101
rect 179 3097 180 3101
rect 174 3096 180 3097
rect 318 3101 324 3102
rect 318 3097 319 3101
rect 323 3097 324 3101
rect 318 3096 324 3097
rect 470 3101 476 3102
rect 470 3097 471 3101
rect 475 3097 476 3101
rect 470 3096 476 3097
rect 622 3101 628 3102
rect 622 3097 623 3101
rect 627 3097 628 3101
rect 622 3096 628 3097
rect 774 3101 780 3102
rect 774 3097 775 3101
rect 779 3097 780 3101
rect 774 3096 780 3097
rect 918 3101 924 3102
rect 918 3097 919 3101
rect 923 3097 924 3101
rect 918 3096 924 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1198 3101 1204 3102
rect 1198 3097 1199 3101
rect 1203 3097 1204 3101
rect 1198 3096 1204 3097
rect 1342 3101 1348 3102
rect 1342 3097 1343 3101
rect 1347 3097 1348 3101
rect 1342 3096 1348 3097
rect 1486 3101 1492 3102
rect 1486 3097 1487 3101
rect 1491 3097 1492 3101
rect 1486 3096 1492 3097
rect 1766 3100 1772 3101
rect 1766 3096 1767 3100
rect 1771 3096 1772 3100
rect 110 3095 116 3096
rect 1766 3095 1772 3096
rect 1806 3088 1812 3089
rect 3462 3088 3468 3089
rect 1806 3084 1807 3088
rect 1811 3084 1812 3088
rect 1806 3083 1812 3084
rect 1934 3087 1940 3088
rect 1934 3083 1935 3087
rect 1939 3083 1940 3087
rect 1934 3082 1940 3083
rect 2054 3087 2060 3088
rect 2054 3083 2055 3087
rect 2059 3083 2060 3087
rect 2054 3082 2060 3083
rect 2174 3087 2180 3088
rect 2174 3083 2175 3087
rect 2179 3083 2180 3087
rect 2174 3082 2180 3083
rect 2302 3087 2308 3088
rect 2302 3083 2303 3087
rect 2307 3083 2308 3087
rect 2302 3082 2308 3083
rect 2430 3087 2436 3088
rect 2430 3083 2431 3087
rect 2435 3083 2436 3087
rect 2430 3082 2436 3083
rect 2566 3087 2572 3088
rect 2566 3083 2567 3087
rect 2571 3083 2572 3087
rect 2566 3082 2572 3083
rect 2718 3087 2724 3088
rect 2718 3083 2719 3087
rect 2723 3083 2724 3087
rect 2718 3082 2724 3083
rect 2870 3087 2876 3088
rect 2870 3083 2871 3087
rect 2875 3083 2876 3087
rect 2870 3082 2876 3083
rect 3030 3087 3036 3088
rect 3030 3083 3031 3087
rect 3035 3083 3036 3087
rect 3030 3082 3036 3083
rect 3198 3087 3204 3088
rect 3198 3083 3199 3087
rect 3203 3083 3204 3087
rect 3198 3082 3204 3083
rect 3366 3087 3372 3088
rect 3366 3083 3367 3087
rect 3371 3083 3372 3087
rect 3462 3084 3463 3088
rect 3467 3084 3468 3088
rect 3462 3083 3468 3084
rect 3366 3082 3372 3083
rect 1806 3071 1812 3072
rect 1806 3067 1807 3071
rect 1811 3067 1812 3071
rect 3462 3071 3468 3072
rect 1806 3066 1812 3067
rect 1934 3068 1940 3069
rect 1934 3064 1935 3068
rect 1939 3064 1940 3068
rect 1934 3063 1940 3064
rect 2054 3068 2060 3069
rect 2054 3064 2055 3068
rect 2059 3064 2060 3068
rect 2054 3063 2060 3064
rect 2174 3068 2180 3069
rect 2174 3064 2175 3068
rect 2179 3064 2180 3068
rect 2174 3063 2180 3064
rect 2302 3068 2308 3069
rect 2302 3064 2303 3068
rect 2307 3064 2308 3068
rect 2302 3063 2308 3064
rect 2430 3068 2436 3069
rect 2430 3064 2431 3068
rect 2435 3064 2436 3068
rect 2430 3063 2436 3064
rect 2566 3068 2572 3069
rect 2566 3064 2567 3068
rect 2571 3064 2572 3068
rect 2566 3063 2572 3064
rect 2718 3068 2724 3069
rect 2718 3064 2719 3068
rect 2723 3064 2724 3068
rect 2718 3063 2724 3064
rect 2870 3068 2876 3069
rect 2870 3064 2871 3068
rect 2875 3064 2876 3068
rect 2870 3063 2876 3064
rect 3030 3068 3036 3069
rect 3030 3064 3031 3068
rect 3035 3064 3036 3068
rect 3030 3063 3036 3064
rect 3198 3068 3204 3069
rect 3198 3064 3199 3068
rect 3203 3064 3204 3068
rect 3198 3063 3204 3064
rect 3366 3068 3372 3069
rect 3366 3064 3367 3068
rect 3371 3064 3372 3068
rect 3462 3067 3463 3071
rect 3467 3067 3468 3071
rect 3462 3066 3468 3067
rect 3366 3063 3372 3064
rect 110 3048 116 3049
rect 1766 3048 1772 3049
rect 110 3044 111 3048
rect 115 3044 116 3048
rect 110 3043 116 3044
rect 134 3047 140 3048
rect 134 3043 135 3047
rect 139 3043 140 3047
rect 134 3042 140 3043
rect 262 3047 268 3048
rect 262 3043 263 3047
rect 267 3043 268 3047
rect 262 3042 268 3043
rect 430 3047 436 3048
rect 430 3043 431 3047
rect 435 3043 436 3047
rect 430 3042 436 3043
rect 606 3047 612 3048
rect 606 3043 607 3047
rect 611 3043 612 3047
rect 606 3042 612 3043
rect 790 3047 796 3048
rect 790 3043 791 3047
rect 795 3043 796 3047
rect 790 3042 796 3043
rect 966 3047 972 3048
rect 966 3043 967 3047
rect 971 3043 972 3047
rect 966 3042 972 3043
rect 1142 3047 1148 3048
rect 1142 3043 1143 3047
rect 1147 3043 1148 3047
rect 1142 3042 1148 3043
rect 1326 3047 1332 3048
rect 1326 3043 1327 3047
rect 1331 3043 1332 3047
rect 1326 3042 1332 3043
rect 1510 3047 1516 3048
rect 1510 3043 1511 3047
rect 1515 3043 1516 3047
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 1766 3043 1772 3044
rect 1510 3042 1516 3043
rect 110 3031 116 3032
rect 110 3027 111 3031
rect 115 3027 116 3031
rect 1766 3031 1772 3032
rect 110 3026 116 3027
rect 134 3028 140 3029
rect 134 3024 135 3028
rect 139 3024 140 3028
rect 134 3023 140 3024
rect 262 3028 268 3029
rect 262 3024 263 3028
rect 267 3024 268 3028
rect 262 3023 268 3024
rect 430 3028 436 3029
rect 430 3024 431 3028
rect 435 3024 436 3028
rect 430 3023 436 3024
rect 606 3028 612 3029
rect 606 3024 607 3028
rect 611 3024 612 3028
rect 606 3023 612 3024
rect 790 3028 796 3029
rect 790 3024 791 3028
rect 795 3024 796 3028
rect 790 3023 796 3024
rect 966 3028 972 3029
rect 966 3024 967 3028
rect 971 3024 972 3028
rect 966 3023 972 3024
rect 1142 3028 1148 3029
rect 1142 3024 1143 3028
rect 1147 3024 1148 3028
rect 1142 3023 1148 3024
rect 1326 3028 1332 3029
rect 1326 3024 1327 3028
rect 1331 3024 1332 3028
rect 1326 3023 1332 3024
rect 1510 3028 1516 3029
rect 1510 3024 1511 3028
rect 1515 3024 1516 3028
rect 1766 3027 1767 3031
rect 1771 3027 1772 3031
rect 1766 3026 1772 3027
rect 1510 3023 1516 3024
rect 2022 3016 2028 3017
rect 1806 3013 1812 3014
rect 1806 3009 1807 3013
rect 1811 3009 1812 3013
rect 2022 3012 2023 3016
rect 2027 3012 2028 3016
rect 2022 3011 2028 3012
rect 2126 3016 2132 3017
rect 2126 3012 2127 3016
rect 2131 3012 2132 3016
rect 2126 3011 2132 3012
rect 2230 3016 2236 3017
rect 2230 3012 2231 3016
rect 2235 3012 2236 3016
rect 2230 3011 2236 3012
rect 2334 3016 2340 3017
rect 2334 3012 2335 3016
rect 2339 3012 2340 3016
rect 2334 3011 2340 3012
rect 2438 3016 2444 3017
rect 2438 3012 2439 3016
rect 2443 3012 2444 3016
rect 2438 3011 2444 3012
rect 2542 3016 2548 3017
rect 2542 3012 2543 3016
rect 2547 3012 2548 3016
rect 2542 3011 2548 3012
rect 2646 3016 2652 3017
rect 2646 3012 2647 3016
rect 2651 3012 2652 3016
rect 2646 3011 2652 3012
rect 2758 3016 2764 3017
rect 2758 3012 2759 3016
rect 2763 3012 2764 3016
rect 2758 3011 2764 3012
rect 3462 3013 3468 3014
rect 1806 3008 1812 3009
rect 3462 3009 3463 3013
rect 3467 3009 3468 3013
rect 3462 3008 3468 3009
rect 2022 2997 2028 2998
rect 1806 2996 1812 2997
rect 1806 2992 1807 2996
rect 1811 2992 1812 2996
rect 2022 2993 2023 2997
rect 2027 2993 2028 2997
rect 2022 2992 2028 2993
rect 2126 2997 2132 2998
rect 2126 2993 2127 2997
rect 2131 2993 2132 2997
rect 2126 2992 2132 2993
rect 2230 2997 2236 2998
rect 2230 2993 2231 2997
rect 2235 2993 2236 2997
rect 2230 2992 2236 2993
rect 2334 2997 2340 2998
rect 2334 2993 2335 2997
rect 2339 2993 2340 2997
rect 2334 2992 2340 2993
rect 2438 2997 2444 2998
rect 2438 2993 2439 2997
rect 2443 2993 2444 2997
rect 2438 2992 2444 2993
rect 2542 2997 2548 2998
rect 2542 2993 2543 2997
rect 2547 2993 2548 2997
rect 2542 2992 2548 2993
rect 2646 2997 2652 2998
rect 2646 2993 2647 2997
rect 2651 2993 2652 2997
rect 2646 2992 2652 2993
rect 2758 2997 2764 2998
rect 2758 2993 2759 2997
rect 2763 2993 2764 2997
rect 2758 2992 2764 2993
rect 3462 2996 3468 2997
rect 3462 2992 3463 2996
rect 3467 2992 3468 2996
rect 1806 2991 1812 2992
rect 3462 2991 3468 2992
rect 134 2980 140 2981
rect 110 2977 116 2978
rect 110 2973 111 2977
rect 115 2973 116 2977
rect 134 2976 135 2980
rect 139 2976 140 2980
rect 134 2975 140 2976
rect 326 2980 332 2981
rect 326 2976 327 2980
rect 331 2976 332 2980
rect 326 2975 332 2976
rect 534 2980 540 2981
rect 534 2976 535 2980
rect 539 2976 540 2980
rect 534 2975 540 2976
rect 734 2980 740 2981
rect 734 2976 735 2980
rect 739 2976 740 2980
rect 734 2975 740 2976
rect 926 2980 932 2981
rect 926 2976 927 2980
rect 931 2976 932 2980
rect 926 2975 932 2976
rect 1102 2980 1108 2981
rect 1102 2976 1103 2980
rect 1107 2976 1108 2980
rect 1102 2975 1108 2976
rect 1278 2980 1284 2981
rect 1278 2976 1279 2980
rect 1283 2976 1284 2980
rect 1278 2975 1284 2976
rect 1446 2980 1452 2981
rect 1446 2976 1447 2980
rect 1451 2976 1452 2980
rect 1446 2975 1452 2976
rect 1622 2980 1628 2981
rect 1622 2976 1623 2980
rect 1627 2976 1628 2980
rect 1622 2975 1628 2976
rect 1766 2977 1772 2978
rect 110 2972 116 2973
rect 1766 2973 1767 2977
rect 1771 2973 1772 2977
rect 1766 2972 1772 2973
rect 134 2961 140 2962
rect 110 2960 116 2961
rect 110 2956 111 2960
rect 115 2956 116 2960
rect 134 2957 135 2961
rect 139 2957 140 2961
rect 134 2956 140 2957
rect 326 2961 332 2962
rect 326 2957 327 2961
rect 331 2957 332 2961
rect 326 2956 332 2957
rect 534 2961 540 2962
rect 534 2957 535 2961
rect 539 2957 540 2961
rect 534 2956 540 2957
rect 734 2961 740 2962
rect 734 2957 735 2961
rect 739 2957 740 2961
rect 734 2956 740 2957
rect 926 2961 932 2962
rect 926 2957 927 2961
rect 931 2957 932 2961
rect 926 2956 932 2957
rect 1102 2961 1108 2962
rect 1102 2957 1103 2961
rect 1107 2957 1108 2961
rect 1102 2956 1108 2957
rect 1278 2961 1284 2962
rect 1278 2957 1279 2961
rect 1283 2957 1284 2961
rect 1278 2956 1284 2957
rect 1446 2961 1452 2962
rect 1446 2957 1447 2961
rect 1451 2957 1452 2961
rect 1446 2956 1452 2957
rect 1622 2961 1628 2962
rect 1622 2957 1623 2961
rect 1627 2957 1628 2961
rect 1622 2956 1628 2957
rect 1766 2960 1772 2961
rect 1766 2956 1767 2960
rect 1771 2956 1772 2960
rect 110 2955 116 2956
rect 1766 2955 1772 2956
rect 1806 2952 1812 2953
rect 3462 2952 3468 2953
rect 1806 2948 1807 2952
rect 1811 2948 1812 2952
rect 1806 2947 1812 2948
rect 2054 2951 2060 2952
rect 2054 2947 2055 2951
rect 2059 2947 2060 2951
rect 2054 2946 2060 2947
rect 2142 2951 2148 2952
rect 2142 2947 2143 2951
rect 2147 2947 2148 2951
rect 2142 2946 2148 2947
rect 2230 2951 2236 2952
rect 2230 2947 2231 2951
rect 2235 2947 2236 2951
rect 2230 2946 2236 2947
rect 2318 2951 2324 2952
rect 2318 2947 2319 2951
rect 2323 2947 2324 2951
rect 2318 2946 2324 2947
rect 2406 2951 2412 2952
rect 2406 2947 2407 2951
rect 2411 2947 2412 2951
rect 2406 2946 2412 2947
rect 2494 2951 2500 2952
rect 2494 2947 2495 2951
rect 2499 2947 2500 2951
rect 2494 2946 2500 2947
rect 2582 2951 2588 2952
rect 2582 2947 2583 2951
rect 2587 2947 2588 2951
rect 2582 2946 2588 2947
rect 2670 2951 2676 2952
rect 2670 2947 2671 2951
rect 2675 2947 2676 2951
rect 2670 2946 2676 2947
rect 2758 2951 2764 2952
rect 2758 2947 2759 2951
rect 2763 2947 2764 2951
rect 2758 2946 2764 2947
rect 2846 2951 2852 2952
rect 2846 2947 2847 2951
rect 2851 2947 2852 2951
rect 3462 2948 3463 2952
rect 3467 2948 3468 2952
rect 3462 2947 3468 2948
rect 2846 2946 2852 2947
rect 1806 2935 1812 2936
rect 1806 2931 1807 2935
rect 1811 2931 1812 2935
rect 3462 2935 3468 2936
rect 1806 2930 1812 2931
rect 2054 2932 2060 2933
rect 2054 2928 2055 2932
rect 2059 2928 2060 2932
rect 2054 2927 2060 2928
rect 2142 2932 2148 2933
rect 2142 2928 2143 2932
rect 2147 2928 2148 2932
rect 2142 2927 2148 2928
rect 2230 2932 2236 2933
rect 2230 2928 2231 2932
rect 2235 2928 2236 2932
rect 2230 2927 2236 2928
rect 2318 2932 2324 2933
rect 2318 2928 2319 2932
rect 2323 2928 2324 2932
rect 2318 2927 2324 2928
rect 2406 2932 2412 2933
rect 2406 2928 2407 2932
rect 2411 2928 2412 2932
rect 2406 2927 2412 2928
rect 2494 2932 2500 2933
rect 2494 2928 2495 2932
rect 2499 2928 2500 2932
rect 2494 2927 2500 2928
rect 2582 2932 2588 2933
rect 2582 2928 2583 2932
rect 2587 2928 2588 2932
rect 2582 2927 2588 2928
rect 2670 2932 2676 2933
rect 2670 2928 2671 2932
rect 2675 2928 2676 2932
rect 2670 2927 2676 2928
rect 2758 2932 2764 2933
rect 2758 2928 2759 2932
rect 2763 2928 2764 2932
rect 2758 2927 2764 2928
rect 2846 2932 2852 2933
rect 2846 2928 2847 2932
rect 2851 2928 2852 2932
rect 3462 2931 3463 2935
rect 3467 2931 3468 2935
rect 3462 2930 3468 2931
rect 2846 2927 2852 2928
rect 110 2908 116 2909
rect 1766 2908 1772 2909
rect 110 2904 111 2908
rect 115 2904 116 2908
rect 110 2903 116 2904
rect 134 2907 140 2908
rect 134 2903 135 2907
rect 139 2903 140 2907
rect 134 2902 140 2903
rect 262 2907 268 2908
rect 262 2903 263 2907
rect 267 2903 268 2907
rect 262 2902 268 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 606 2907 612 2908
rect 606 2903 607 2907
rect 611 2903 612 2907
rect 606 2902 612 2903
rect 782 2907 788 2908
rect 782 2903 783 2907
rect 787 2903 788 2907
rect 782 2902 788 2903
rect 950 2907 956 2908
rect 950 2903 951 2907
rect 955 2903 956 2907
rect 950 2902 956 2903
rect 1110 2907 1116 2908
rect 1110 2903 1111 2907
rect 1115 2903 1116 2907
rect 1110 2902 1116 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1430 2907 1436 2908
rect 1430 2903 1431 2907
rect 1435 2903 1436 2907
rect 1430 2902 1436 2903
rect 1590 2907 1596 2908
rect 1590 2903 1591 2907
rect 1595 2903 1596 2907
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1590 2902 1596 2903
rect 110 2891 116 2892
rect 110 2887 111 2891
rect 115 2887 116 2891
rect 1766 2891 1772 2892
rect 110 2886 116 2887
rect 134 2888 140 2889
rect 134 2884 135 2888
rect 139 2884 140 2888
rect 134 2883 140 2884
rect 262 2888 268 2889
rect 262 2884 263 2888
rect 267 2884 268 2888
rect 262 2883 268 2884
rect 430 2888 436 2889
rect 430 2884 431 2888
rect 435 2884 436 2888
rect 430 2883 436 2884
rect 606 2888 612 2889
rect 606 2884 607 2888
rect 611 2884 612 2888
rect 606 2883 612 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 950 2888 956 2889
rect 950 2884 951 2888
rect 955 2884 956 2888
rect 950 2883 956 2884
rect 1110 2888 1116 2889
rect 1110 2884 1111 2888
rect 1115 2884 1116 2888
rect 1110 2883 1116 2884
rect 1270 2888 1276 2889
rect 1270 2884 1271 2888
rect 1275 2884 1276 2888
rect 1270 2883 1276 2884
rect 1430 2888 1436 2889
rect 1430 2884 1431 2888
rect 1435 2884 1436 2888
rect 1430 2883 1436 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1766 2887 1767 2891
rect 1771 2887 1772 2891
rect 1766 2886 1772 2887
rect 1590 2883 1596 2884
rect 2070 2880 2076 2881
rect 1806 2877 1812 2878
rect 1806 2873 1807 2877
rect 1811 2873 1812 2877
rect 2070 2876 2071 2880
rect 2075 2876 2076 2880
rect 2070 2875 2076 2876
rect 2174 2880 2180 2881
rect 2174 2876 2175 2880
rect 2179 2876 2180 2880
rect 2174 2875 2180 2876
rect 2270 2880 2276 2881
rect 2270 2876 2271 2880
rect 2275 2876 2276 2880
rect 2270 2875 2276 2876
rect 2366 2880 2372 2881
rect 2366 2876 2367 2880
rect 2371 2876 2372 2880
rect 2366 2875 2372 2876
rect 2470 2880 2476 2881
rect 2470 2876 2471 2880
rect 2475 2876 2476 2880
rect 2470 2875 2476 2876
rect 2574 2880 2580 2881
rect 2574 2876 2575 2880
rect 2579 2876 2580 2880
rect 2574 2875 2580 2876
rect 2678 2880 2684 2881
rect 2678 2876 2679 2880
rect 2683 2876 2684 2880
rect 2678 2875 2684 2876
rect 2782 2880 2788 2881
rect 2782 2876 2783 2880
rect 2787 2876 2788 2880
rect 2782 2875 2788 2876
rect 3462 2877 3468 2878
rect 1806 2872 1812 2873
rect 3462 2873 3463 2877
rect 3467 2873 3468 2877
rect 3462 2872 3468 2873
rect 2070 2861 2076 2862
rect 1806 2860 1812 2861
rect 1806 2856 1807 2860
rect 1811 2856 1812 2860
rect 2070 2857 2071 2861
rect 2075 2857 2076 2861
rect 2070 2856 2076 2857
rect 2174 2861 2180 2862
rect 2174 2857 2175 2861
rect 2179 2857 2180 2861
rect 2174 2856 2180 2857
rect 2270 2861 2276 2862
rect 2270 2857 2271 2861
rect 2275 2857 2276 2861
rect 2270 2856 2276 2857
rect 2366 2861 2372 2862
rect 2366 2857 2367 2861
rect 2371 2857 2372 2861
rect 2366 2856 2372 2857
rect 2470 2861 2476 2862
rect 2470 2857 2471 2861
rect 2475 2857 2476 2861
rect 2470 2856 2476 2857
rect 2574 2861 2580 2862
rect 2574 2857 2575 2861
rect 2579 2857 2580 2861
rect 2574 2856 2580 2857
rect 2678 2861 2684 2862
rect 2678 2857 2679 2861
rect 2683 2857 2684 2861
rect 2678 2856 2684 2857
rect 2782 2861 2788 2862
rect 2782 2857 2783 2861
rect 2787 2857 2788 2861
rect 2782 2856 2788 2857
rect 3462 2860 3468 2861
rect 3462 2856 3463 2860
rect 3467 2856 3468 2860
rect 1806 2855 1812 2856
rect 3462 2855 3468 2856
rect 134 2840 140 2841
rect 110 2837 116 2838
rect 110 2833 111 2837
rect 115 2833 116 2837
rect 134 2836 135 2840
rect 139 2836 140 2840
rect 134 2835 140 2836
rect 254 2840 260 2841
rect 254 2836 255 2840
rect 259 2836 260 2840
rect 254 2835 260 2836
rect 406 2840 412 2841
rect 406 2836 407 2840
rect 411 2836 412 2840
rect 406 2835 412 2836
rect 566 2840 572 2841
rect 566 2836 567 2840
rect 571 2836 572 2840
rect 566 2835 572 2836
rect 726 2840 732 2841
rect 726 2836 727 2840
rect 731 2836 732 2840
rect 726 2835 732 2836
rect 878 2840 884 2841
rect 878 2836 879 2840
rect 883 2836 884 2840
rect 878 2835 884 2836
rect 1022 2840 1028 2841
rect 1022 2836 1023 2840
rect 1027 2836 1028 2840
rect 1022 2835 1028 2836
rect 1166 2840 1172 2841
rect 1166 2836 1167 2840
rect 1171 2836 1172 2840
rect 1166 2835 1172 2836
rect 1310 2840 1316 2841
rect 1310 2836 1311 2840
rect 1315 2836 1316 2840
rect 1310 2835 1316 2836
rect 1462 2840 1468 2841
rect 1462 2836 1463 2840
rect 1467 2836 1468 2840
rect 1462 2835 1468 2836
rect 1766 2837 1772 2838
rect 110 2832 116 2833
rect 1766 2833 1767 2837
rect 1771 2833 1772 2837
rect 1766 2832 1772 2833
rect 134 2821 140 2822
rect 110 2820 116 2821
rect 110 2816 111 2820
rect 115 2816 116 2820
rect 134 2817 135 2821
rect 139 2817 140 2821
rect 134 2816 140 2817
rect 254 2821 260 2822
rect 254 2817 255 2821
rect 259 2817 260 2821
rect 254 2816 260 2817
rect 406 2821 412 2822
rect 406 2817 407 2821
rect 411 2817 412 2821
rect 406 2816 412 2817
rect 566 2821 572 2822
rect 566 2817 567 2821
rect 571 2817 572 2821
rect 566 2816 572 2817
rect 726 2821 732 2822
rect 726 2817 727 2821
rect 731 2817 732 2821
rect 726 2816 732 2817
rect 878 2821 884 2822
rect 878 2817 879 2821
rect 883 2817 884 2821
rect 878 2816 884 2817
rect 1022 2821 1028 2822
rect 1022 2817 1023 2821
rect 1027 2817 1028 2821
rect 1022 2816 1028 2817
rect 1166 2821 1172 2822
rect 1166 2817 1167 2821
rect 1171 2817 1172 2821
rect 1166 2816 1172 2817
rect 1310 2821 1316 2822
rect 1310 2817 1311 2821
rect 1315 2817 1316 2821
rect 1310 2816 1316 2817
rect 1462 2821 1468 2822
rect 1462 2817 1463 2821
rect 1467 2817 1468 2821
rect 1462 2816 1468 2817
rect 1766 2820 1772 2821
rect 1766 2816 1767 2820
rect 1771 2816 1772 2820
rect 110 2815 116 2816
rect 1766 2815 1772 2816
rect 1806 2812 1812 2813
rect 3462 2812 3468 2813
rect 1806 2808 1807 2812
rect 1811 2808 1812 2812
rect 1806 2807 1812 2808
rect 1982 2811 1988 2812
rect 1982 2807 1983 2811
rect 1987 2807 1988 2811
rect 1982 2806 1988 2807
rect 2110 2811 2116 2812
rect 2110 2807 2111 2811
rect 2115 2807 2116 2811
rect 2110 2806 2116 2807
rect 2238 2811 2244 2812
rect 2238 2807 2239 2811
rect 2243 2807 2244 2811
rect 2238 2806 2244 2807
rect 2366 2811 2372 2812
rect 2366 2807 2367 2811
rect 2371 2807 2372 2811
rect 2366 2806 2372 2807
rect 2486 2811 2492 2812
rect 2486 2807 2487 2811
rect 2491 2807 2492 2811
rect 2486 2806 2492 2807
rect 2606 2811 2612 2812
rect 2606 2807 2607 2811
rect 2611 2807 2612 2811
rect 2606 2806 2612 2807
rect 2718 2811 2724 2812
rect 2718 2807 2719 2811
rect 2723 2807 2724 2811
rect 2718 2806 2724 2807
rect 2838 2811 2844 2812
rect 2838 2807 2839 2811
rect 2843 2807 2844 2811
rect 2838 2806 2844 2807
rect 2958 2811 2964 2812
rect 2958 2807 2959 2811
rect 2963 2807 2964 2811
rect 3462 2808 3463 2812
rect 3467 2808 3468 2812
rect 3462 2807 3468 2808
rect 2958 2806 2964 2807
rect 1806 2795 1812 2796
rect 1806 2791 1807 2795
rect 1811 2791 1812 2795
rect 3462 2795 3468 2796
rect 1806 2790 1812 2791
rect 1982 2792 1988 2793
rect 1982 2788 1983 2792
rect 1987 2788 1988 2792
rect 1982 2787 1988 2788
rect 2110 2792 2116 2793
rect 2110 2788 2111 2792
rect 2115 2788 2116 2792
rect 2110 2787 2116 2788
rect 2238 2792 2244 2793
rect 2238 2788 2239 2792
rect 2243 2788 2244 2792
rect 2238 2787 2244 2788
rect 2366 2792 2372 2793
rect 2366 2788 2367 2792
rect 2371 2788 2372 2792
rect 2366 2787 2372 2788
rect 2486 2792 2492 2793
rect 2486 2788 2487 2792
rect 2491 2788 2492 2792
rect 2486 2787 2492 2788
rect 2606 2792 2612 2793
rect 2606 2788 2607 2792
rect 2611 2788 2612 2792
rect 2606 2787 2612 2788
rect 2718 2792 2724 2793
rect 2718 2788 2719 2792
rect 2723 2788 2724 2792
rect 2718 2787 2724 2788
rect 2838 2792 2844 2793
rect 2838 2788 2839 2792
rect 2843 2788 2844 2792
rect 2838 2787 2844 2788
rect 2958 2792 2964 2793
rect 2958 2788 2959 2792
rect 2963 2788 2964 2792
rect 3462 2791 3463 2795
rect 3467 2791 3468 2795
rect 3462 2790 3468 2791
rect 2958 2787 2964 2788
rect 110 2768 116 2769
rect 1766 2768 1772 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 286 2767 292 2768
rect 286 2763 287 2767
rect 291 2763 292 2767
rect 286 2762 292 2763
rect 390 2767 396 2768
rect 390 2763 391 2767
rect 395 2763 396 2767
rect 390 2762 396 2763
rect 502 2767 508 2768
rect 502 2763 503 2767
rect 507 2763 508 2767
rect 502 2762 508 2763
rect 622 2767 628 2768
rect 622 2763 623 2767
rect 627 2763 628 2767
rect 622 2762 628 2763
rect 742 2767 748 2768
rect 742 2763 743 2767
rect 747 2763 748 2767
rect 742 2762 748 2763
rect 854 2767 860 2768
rect 854 2763 855 2767
rect 859 2763 860 2767
rect 854 2762 860 2763
rect 966 2767 972 2768
rect 966 2763 967 2767
rect 971 2763 972 2767
rect 966 2762 972 2763
rect 1078 2767 1084 2768
rect 1078 2763 1079 2767
rect 1083 2763 1084 2767
rect 1078 2762 1084 2763
rect 1198 2767 1204 2768
rect 1198 2763 1199 2767
rect 1203 2763 1204 2767
rect 1198 2762 1204 2763
rect 1318 2767 1324 2768
rect 1318 2763 1319 2767
rect 1323 2763 1324 2767
rect 1766 2764 1767 2768
rect 1771 2764 1772 2768
rect 1766 2763 1772 2764
rect 1318 2762 1324 2763
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 1766 2751 1772 2752
rect 110 2746 116 2747
rect 286 2748 292 2749
rect 286 2744 287 2748
rect 291 2744 292 2748
rect 286 2743 292 2744
rect 390 2748 396 2749
rect 390 2744 391 2748
rect 395 2744 396 2748
rect 390 2743 396 2744
rect 502 2748 508 2749
rect 502 2744 503 2748
rect 507 2744 508 2748
rect 502 2743 508 2744
rect 622 2748 628 2749
rect 622 2744 623 2748
rect 627 2744 628 2748
rect 622 2743 628 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 854 2748 860 2749
rect 854 2744 855 2748
rect 859 2744 860 2748
rect 854 2743 860 2744
rect 966 2748 972 2749
rect 966 2744 967 2748
rect 971 2744 972 2748
rect 966 2743 972 2744
rect 1078 2748 1084 2749
rect 1078 2744 1079 2748
rect 1083 2744 1084 2748
rect 1078 2743 1084 2744
rect 1198 2748 1204 2749
rect 1198 2744 1199 2748
rect 1203 2744 1204 2748
rect 1198 2743 1204 2744
rect 1318 2748 1324 2749
rect 1318 2744 1319 2748
rect 1323 2744 1324 2748
rect 1766 2747 1767 2751
rect 1771 2747 1772 2751
rect 1766 2746 1772 2747
rect 1318 2743 1324 2744
rect 1886 2744 1892 2745
rect 1806 2741 1812 2742
rect 1806 2737 1807 2741
rect 1811 2737 1812 2741
rect 1886 2740 1887 2744
rect 1891 2740 1892 2744
rect 1886 2739 1892 2740
rect 2030 2744 2036 2745
rect 2030 2740 2031 2744
rect 2035 2740 2036 2744
rect 2030 2739 2036 2740
rect 2182 2744 2188 2745
rect 2182 2740 2183 2744
rect 2187 2740 2188 2744
rect 2182 2739 2188 2740
rect 2334 2744 2340 2745
rect 2334 2740 2335 2744
rect 2339 2740 2340 2744
rect 2334 2739 2340 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2622 2744 2628 2745
rect 2622 2740 2623 2744
rect 2627 2740 2628 2744
rect 2622 2739 2628 2740
rect 2766 2744 2772 2745
rect 2766 2740 2767 2744
rect 2771 2740 2772 2744
rect 2766 2739 2772 2740
rect 2910 2744 2916 2745
rect 2910 2740 2911 2744
rect 2915 2740 2916 2744
rect 2910 2739 2916 2740
rect 3054 2744 3060 2745
rect 3054 2740 3055 2744
rect 3059 2740 3060 2744
rect 3054 2739 3060 2740
rect 3462 2741 3468 2742
rect 1806 2736 1812 2737
rect 3462 2737 3463 2741
rect 3467 2737 3468 2741
rect 3462 2736 3468 2737
rect 1886 2725 1892 2726
rect 1806 2724 1812 2725
rect 1806 2720 1807 2724
rect 1811 2720 1812 2724
rect 1886 2721 1887 2725
rect 1891 2721 1892 2725
rect 1886 2720 1892 2721
rect 2030 2725 2036 2726
rect 2030 2721 2031 2725
rect 2035 2721 2036 2725
rect 2030 2720 2036 2721
rect 2182 2725 2188 2726
rect 2182 2721 2183 2725
rect 2187 2721 2188 2725
rect 2182 2720 2188 2721
rect 2334 2725 2340 2726
rect 2334 2721 2335 2725
rect 2339 2721 2340 2725
rect 2334 2720 2340 2721
rect 2478 2725 2484 2726
rect 2478 2721 2479 2725
rect 2483 2721 2484 2725
rect 2478 2720 2484 2721
rect 2622 2725 2628 2726
rect 2622 2721 2623 2725
rect 2627 2721 2628 2725
rect 2622 2720 2628 2721
rect 2766 2725 2772 2726
rect 2766 2721 2767 2725
rect 2771 2721 2772 2725
rect 2766 2720 2772 2721
rect 2910 2725 2916 2726
rect 2910 2721 2911 2725
rect 2915 2721 2916 2725
rect 2910 2720 2916 2721
rect 3054 2725 3060 2726
rect 3054 2721 3055 2725
rect 3059 2721 3060 2725
rect 3054 2720 3060 2721
rect 3462 2724 3468 2725
rect 3462 2720 3463 2724
rect 3467 2720 3468 2724
rect 1806 2719 1812 2720
rect 3462 2719 3468 2720
rect 478 2700 484 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 566 2700 572 2701
rect 566 2696 567 2700
rect 571 2696 572 2700
rect 566 2695 572 2696
rect 654 2700 660 2701
rect 654 2696 655 2700
rect 659 2696 660 2700
rect 654 2695 660 2696
rect 742 2700 748 2701
rect 742 2696 743 2700
rect 747 2696 748 2700
rect 742 2695 748 2696
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 918 2700 924 2701
rect 918 2696 919 2700
rect 923 2696 924 2700
rect 918 2695 924 2696
rect 1006 2700 1012 2701
rect 1006 2696 1007 2700
rect 1011 2696 1012 2700
rect 1006 2695 1012 2696
rect 1094 2700 1100 2701
rect 1094 2696 1095 2700
rect 1099 2696 1100 2700
rect 1094 2695 1100 2696
rect 1182 2700 1188 2701
rect 1182 2696 1183 2700
rect 1187 2696 1188 2700
rect 1182 2695 1188 2696
rect 1766 2697 1772 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1766 2692 1772 2693
rect 478 2681 484 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 566 2681 572 2682
rect 566 2677 567 2681
rect 571 2677 572 2681
rect 566 2676 572 2677
rect 654 2681 660 2682
rect 654 2677 655 2681
rect 659 2677 660 2681
rect 654 2676 660 2677
rect 742 2681 748 2682
rect 742 2677 743 2681
rect 747 2677 748 2681
rect 742 2676 748 2677
rect 830 2681 836 2682
rect 830 2677 831 2681
rect 835 2677 836 2681
rect 830 2676 836 2677
rect 918 2681 924 2682
rect 918 2677 919 2681
rect 923 2677 924 2681
rect 918 2676 924 2677
rect 1006 2681 1012 2682
rect 1006 2677 1007 2681
rect 1011 2677 1012 2681
rect 1006 2676 1012 2677
rect 1094 2681 1100 2682
rect 1094 2677 1095 2681
rect 1099 2677 1100 2681
rect 1094 2676 1100 2677
rect 1182 2681 1188 2682
rect 1182 2677 1183 2681
rect 1187 2677 1188 2681
rect 1182 2676 1188 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 110 2675 116 2676
rect 1766 2675 1772 2676
rect 1806 2680 1812 2681
rect 3462 2680 3468 2681
rect 1806 2676 1807 2680
rect 1811 2676 1812 2680
rect 1806 2675 1812 2676
rect 1830 2679 1836 2680
rect 1830 2675 1831 2679
rect 1835 2675 1836 2679
rect 1830 2674 1836 2675
rect 2022 2679 2028 2680
rect 2022 2675 2023 2679
rect 2027 2675 2028 2679
rect 2022 2674 2028 2675
rect 2230 2679 2236 2680
rect 2230 2675 2231 2679
rect 2235 2675 2236 2679
rect 2230 2674 2236 2675
rect 2430 2679 2436 2680
rect 2430 2675 2431 2679
rect 2435 2675 2436 2679
rect 2430 2674 2436 2675
rect 2614 2679 2620 2680
rect 2614 2675 2615 2679
rect 2619 2675 2620 2679
rect 2614 2674 2620 2675
rect 2782 2679 2788 2680
rect 2782 2675 2783 2679
rect 2787 2675 2788 2679
rect 2782 2674 2788 2675
rect 2942 2679 2948 2680
rect 2942 2675 2943 2679
rect 2947 2675 2948 2679
rect 2942 2674 2948 2675
rect 3094 2679 3100 2680
rect 3094 2675 3095 2679
rect 3099 2675 3100 2679
rect 3094 2674 3100 2675
rect 3238 2679 3244 2680
rect 3238 2675 3239 2679
rect 3243 2675 3244 2679
rect 3238 2674 3244 2675
rect 3366 2679 3372 2680
rect 3366 2675 3367 2679
rect 3371 2675 3372 2679
rect 3462 2676 3463 2680
rect 3467 2676 3468 2680
rect 3462 2675 3468 2676
rect 3366 2674 3372 2675
rect 1806 2663 1812 2664
rect 1806 2659 1807 2663
rect 1811 2659 1812 2663
rect 3462 2663 3468 2664
rect 1806 2658 1812 2659
rect 1830 2660 1836 2661
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 2022 2660 2028 2661
rect 2022 2656 2023 2660
rect 2027 2656 2028 2660
rect 2022 2655 2028 2656
rect 2230 2660 2236 2661
rect 2230 2656 2231 2660
rect 2235 2656 2236 2660
rect 2230 2655 2236 2656
rect 2430 2660 2436 2661
rect 2430 2656 2431 2660
rect 2435 2656 2436 2660
rect 2430 2655 2436 2656
rect 2614 2660 2620 2661
rect 2614 2656 2615 2660
rect 2619 2656 2620 2660
rect 2614 2655 2620 2656
rect 2782 2660 2788 2661
rect 2782 2656 2783 2660
rect 2787 2656 2788 2660
rect 2782 2655 2788 2656
rect 2942 2660 2948 2661
rect 2942 2656 2943 2660
rect 2947 2656 2948 2660
rect 2942 2655 2948 2656
rect 3094 2660 3100 2661
rect 3094 2656 3095 2660
rect 3099 2656 3100 2660
rect 3094 2655 3100 2656
rect 3238 2660 3244 2661
rect 3238 2656 3239 2660
rect 3243 2656 3244 2660
rect 3238 2655 3244 2656
rect 3366 2660 3372 2661
rect 3366 2656 3367 2660
rect 3371 2656 3372 2660
rect 3462 2659 3463 2663
rect 3467 2659 3468 2663
rect 3462 2658 3468 2659
rect 3366 2655 3372 2656
rect 110 2628 116 2629
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 470 2627 476 2628
rect 470 2623 471 2627
rect 475 2623 476 2627
rect 470 2622 476 2623
rect 558 2627 564 2628
rect 558 2623 559 2627
rect 563 2623 564 2627
rect 558 2622 564 2623
rect 646 2627 652 2628
rect 646 2623 647 2627
rect 651 2623 652 2627
rect 646 2622 652 2623
rect 734 2627 740 2628
rect 734 2623 735 2627
rect 739 2623 740 2627
rect 734 2622 740 2623
rect 822 2627 828 2628
rect 822 2623 823 2627
rect 827 2623 828 2627
rect 822 2622 828 2623
rect 910 2627 916 2628
rect 910 2623 911 2627
rect 915 2623 916 2627
rect 910 2622 916 2623
rect 998 2627 1004 2628
rect 998 2623 999 2627
rect 1003 2623 1004 2627
rect 998 2622 1004 2623
rect 1086 2627 1092 2628
rect 1086 2623 1087 2627
rect 1091 2623 1092 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1086 2622 1092 2623
rect 1830 2612 1836 2613
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 470 2608 476 2609
rect 470 2604 471 2608
rect 475 2604 476 2608
rect 470 2603 476 2604
rect 558 2608 564 2609
rect 558 2604 559 2608
rect 563 2604 564 2608
rect 558 2603 564 2604
rect 646 2608 652 2609
rect 646 2604 647 2608
rect 651 2604 652 2608
rect 646 2603 652 2604
rect 734 2608 740 2609
rect 734 2604 735 2608
rect 739 2604 740 2608
rect 734 2603 740 2604
rect 822 2608 828 2609
rect 822 2604 823 2608
rect 827 2604 828 2608
rect 822 2603 828 2604
rect 910 2608 916 2609
rect 910 2604 911 2608
rect 915 2604 916 2608
rect 910 2603 916 2604
rect 998 2608 1004 2609
rect 998 2604 999 2608
rect 1003 2604 1004 2608
rect 998 2603 1004 2604
rect 1086 2608 1092 2609
rect 1086 2604 1087 2608
rect 1091 2604 1092 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1766 2606 1772 2607
rect 1806 2609 1812 2610
rect 1806 2605 1807 2609
rect 1811 2605 1812 2609
rect 1830 2608 1831 2612
rect 1835 2608 1836 2612
rect 1830 2607 1836 2608
rect 1998 2612 2004 2613
rect 1998 2608 1999 2612
rect 2003 2608 2004 2612
rect 1998 2607 2004 2608
rect 2182 2612 2188 2613
rect 2182 2608 2183 2612
rect 2187 2608 2188 2612
rect 2182 2607 2188 2608
rect 2358 2612 2364 2613
rect 2358 2608 2359 2612
rect 2363 2608 2364 2612
rect 2358 2607 2364 2608
rect 2518 2612 2524 2613
rect 2518 2608 2519 2612
rect 2523 2608 2524 2612
rect 2518 2607 2524 2608
rect 2670 2612 2676 2613
rect 2670 2608 2671 2612
rect 2675 2608 2676 2612
rect 2670 2607 2676 2608
rect 2806 2612 2812 2613
rect 2806 2608 2807 2612
rect 2811 2608 2812 2612
rect 2806 2607 2812 2608
rect 2926 2612 2932 2613
rect 2926 2608 2927 2612
rect 2931 2608 2932 2612
rect 2926 2607 2932 2608
rect 3046 2612 3052 2613
rect 3046 2608 3047 2612
rect 3051 2608 3052 2612
rect 3046 2607 3052 2608
rect 3158 2612 3164 2613
rect 3158 2608 3159 2612
rect 3163 2608 3164 2612
rect 3158 2607 3164 2608
rect 3270 2612 3276 2613
rect 3270 2608 3271 2612
rect 3275 2608 3276 2612
rect 3270 2607 3276 2608
rect 3366 2612 3372 2613
rect 3366 2608 3367 2612
rect 3371 2608 3372 2612
rect 3366 2607 3372 2608
rect 3462 2609 3468 2610
rect 1806 2604 1812 2605
rect 3462 2605 3463 2609
rect 3467 2605 3468 2609
rect 3462 2604 3468 2605
rect 1086 2603 1092 2604
rect 1830 2593 1836 2594
rect 1806 2592 1812 2593
rect 1806 2588 1807 2592
rect 1811 2588 1812 2592
rect 1830 2589 1831 2593
rect 1835 2589 1836 2593
rect 1830 2588 1836 2589
rect 1998 2593 2004 2594
rect 1998 2589 1999 2593
rect 2003 2589 2004 2593
rect 1998 2588 2004 2589
rect 2182 2593 2188 2594
rect 2182 2589 2183 2593
rect 2187 2589 2188 2593
rect 2182 2588 2188 2589
rect 2358 2593 2364 2594
rect 2358 2589 2359 2593
rect 2363 2589 2364 2593
rect 2358 2588 2364 2589
rect 2518 2593 2524 2594
rect 2518 2589 2519 2593
rect 2523 2589 2524 2593
rect 2518 2588 2524 2589
rect 2670 2593 2676 2594
rect 2670 2589 2671 2593
rect 2675 2589 2676 2593
rect 2670 2588 2676 2589
rect 2806 2593 2812 2594
rect 2806 2589 2807 2593
rect 2811 2589 2812 2593
rect 2806 2588 2812 2589
rect 2926 2593 2932 2594
rect 2926 2589 2927 2593
rect 2931 2589 2932 2593
rect 2926 2588 2932 2589
rect 3046 2593 3052 2594
rect 3046 2589 3047 2593
rect 3051 2589 3052 2593
rect 3046 2588 3052 2589
rect 3158 2593 3164 2594
rect 3158 2589 3159 2593
rect 3163 2589 3164 2593
rect 3158 2588 3164 2589
rect 3270 2593 3276 2594
rect 3270 2589 3271 2593
rect 3275 2589 3276 2593
rect 3270 2588 3276 2589
rect 3366 2593 3372 2594
rect 3366 2589 3367 2593
rect 3371 2589 3372 2593
rect 3366 2588 3372 2589
rect 3462 2592 3468 2593
rect 3462 2588 3463 2592
rect 3467 2588 3468 2592
rect 1806 2587 1812 2588
rect 3462 2587 3468 2588
rect 222 2552 228 2553
rect 110 2549 116 2550
rect 110 2545 111 2549
rect 115 2545 116 2549
rect 222 2548 223 2552
rect 227 2548 228 2552
rect 222 2547 228 2548
rect 310 2552 316 2553
rect 310 2548 311 2552
rect 315 2548 316 2552
rect 310 2547 316 2548
rect 406 2552 412 2553
rect 406 2548 407 2552
rect 411 2548 412 2552
rect 406 2547 412 2548
rect 502 2552 508 2553
rect 502 2548 503 2552
rect 507 2548 508 2552
rect 502 2547 508 2548
rect 590 2552 596 2553
rect 590 2548 591 2552
rect 595 2548 596 2552
rect 590 2547 596 2548
rect 678 2552 684 2553
rect 678 2548 679 2552
rect 683 2548 684 2552
rect 678 2547 684 2548
rect 766 2552 772 2553
rect 766 2548 767 2552
rect 771 2548 772 2552
rect 766 2547 772 2548
rect 854 2552 860 2553
rect 854 2548 855 2552
rect 859 2548 860 2552
rect 854 2547 860 2548
rect 942 2552 948 2553
rect 942 2548 943 2552
rect 947 2548 948 2552
rect 942 2547 948 2548
rect 1030 2552 1036 2553
rect 1030 2548 1031 2552
rect 1035 2548 1036 2552
rect 1030 2547 1036 2548
rect 1118 2552 1124 2553
rect 1118 2548 1119 2552
rect 1123 2548 1124 2552
rect 1118 2547 1124 2548
rect 1214 2552 1220 2553
rect 1214 2548 1215 2552
rect 1219 2548 1220 2552
rect 1214 2547 1220 2548
rect 1310 2552 1316 2553
rect 1310 2548 1311 2552
rect 1315 2548 1316 2552
rect 1310 2547 1316 2548
rect 1406 2552 1412 2553
rect 1406 2548 1407 2552
rect 1411 2548 1412 2552
rect 1406 2547 1412 2548
rect 1494 2552 1500 2553
rect 1494 2548 1495 2552
rect 1499 2548 1500 2552
rect 1494 2547 1500 2548
rect 1582 2552 1588 2553
rect 1582 2548 1583 2552
rect 1587 2548 1588 2552
rect 1582 2547 1588 2548
rect 1670 2552 1676 2553
rect 1670 2548 1671 2552
rect 1675 2548 1676 2552
rect 1670 2547 1676 2548
rect 1766 2549 1772 2550
rect 110 2544 116 2545
rect 1766 2545 1767 2549
rect 1771 2545 1772 2549
rect 1766 2544 1772 2545
rect 1806 2540 1812 2541
rect 3462 2540 3468 2541
rect 1806 2536 1807 2540
rect 1811 2536 1812 2540
rect 1806 2535 1812 2536
rect 2206 2539 2212 2540
rect 2206 2535 2207 2539
rect 2211 2535 2212 2539
rect 2206 2534 2212 2535
rect 2798 2539 2804 2540
rect 2798 2535 2799 2539
rect 2803 2535 2804 2539
rect 2798 2534 2804 2535
rect 3366 2539 3372 2540
rect 3366 2535 3367 2539
rect 3371 2535 3372 2539
rect 3462 2536 3463 2540
rect 3467 2536 3468 2540
rect 3462 2535 3468 2536
rect 3366 2534 3372 2535
rect 222 2533 228 2534
rect 110 2532 116 2533
rect 110 2528 111 2532
rect 115 2528 116 2532
rect 222 2529 223 2533
rect 227 2529 228 2533
rect 222 2528 228 2529
rect 310 2533 316 2534
rect 310 2529 311 2533
rect 315 2529 316 2533
rect 310 2528 316 2529
rect 406 2533 412 2534
rect 406 2529 407 2533
rect 411 2529 412 2533
rect 406 2528 412 2529
rect 502 2533 508 2534
rect 502 2529 503 2533
rect 507 2529 508 2533
rect 502 2528 508 2529
rect 590 2533 596 2534
rect 590 2529 591 2533
rect 595 2529 596 2533
rect 590 2528 596 2529
rect 678 2533 684 2534
rect 678 2529 679 2533
rect 683 2529 684 2533
rect 678 2528 684 2529
rect 766 2533 772 2534
rect 766 2529 767 2533
rect 771 2529 772 2533
rect 766 2528 772 2529
rect 854 2533 860 2534
rect 854 2529 855 2533
rect 859 2529 860 2533
rect 854 2528 860 2529
rect 942 2533 948 2534
rect 942 2529 943 2533
rect 947 2529 948 2533
rect 942 2528 948 2529
rect 1030 2533 1036 2534
rect 1030 2529 1031 2533
rect 1035 2529 1036 2533
rect 1030 2528 1036 2529
rect 1118 2533 1124 2534
rect 1118 2529 1119 2533
rect 1123 2529 1124 2533
rect 1118 2528 1124 2529
rect 1214 2533 1220 2534
rect 1214 2529 1215 2533
rect 1219 2529 1220 2533
rect 1214 2528 1220 2529
rect 1310 2533 1316 2534
rect 1310 2529 1311 2533
rect 1315 2529 1316 2533
rect 1310 2528 1316 2529
rect 1406 2533 1412 2534
rect 1406 2529 1407 2533
rect 1411 2529 1412 2533
rect 1406 2528 1412 2529
rect 1494 2533 1500 2534
rect 1494 2529 1495 2533
rect 1499 2529 1500 2533
rect 1494 2528 1500 2529
rect 1582 2533 1588 2534
rect 1582 2529 1583 2533
rect 1587 2529 1588 2533
rect 1582 2528 1588 2529
rect 1670 2533 1676 2534
rect 1670 2529 1671 2533
rect 1675 2529 1676 2533
rect 1670 2528 1676 2529
rect 1766 2532 1772 2533
rect 1766 2528 1767 2532
rect 1771 2528 1772 2532
rect 110 2527 116 2528
rect 1766 2527 1772 2528
rect 1806 2523 1812 2524
rect 1806 2519 1807 2523
rect 1811 2519 1812 2523
rect 3462 2523 3468 2524
rect 1806 2518 1812 2519
rect 2206 2520 2212 2521
rect 2206 2516 2207 2520
rect 2211 2516 2212 2520
rect 2206 2515 2212 2516
rect 2798 2520 2804 2521
rect 2798 2516 2799 2520
rect 2803 2516 2804 2520
rect 2798 2515 2804 2516
rect 3366 2520 3372 2521
rect 3366 2516 3367 2520
rect 3371 2516 3372 2520
rect 3462 2519 3463 2523
rect 3467 2519 3468 2523
rect 3462 2518 3468 2519
rect 3366 2515 3372 2516
rect 110 2488 116 2489
rect 1766 2488 1772 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 246 2487 252 2488
rect 246 2483 247 2487
rect 251 2483 252 2487
rect 246 2482 252 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 542 2487 548 2488
rect 542 2483 543 2487
rect 547 2483 548 2487
rect 542 2482 548 2483
rect 694 2487 700 2488
rect 694 2483 695 2487
rect 699 2483 700 2487
rect 694 2482 700 2483
rect 838 2487 844 2488
rect 838 2483 839 2487
rect 843 2483 844 2487
rect 838 2482 844 2483
rect 974 2487 980 2488
rect 974 2483 975 2487
rect 979 2483 980 2487
rect 974 2482 980 2483
rect 1102 2487 1108 2488
rect 1102 2483 1103 2487
rect 1107 2483 1108 2487
rect 1102 2482 1108 2483
rect 1230 2487 1236 2488
rect 1230 2483 1231 2487
rect 1235 2483 1236 2487
rect 1230 2482 1236 2483
rect 1350 2487 1356 2488
rect 1350 2483 1351 2487
rect 1355 2483 1356 2487
rect 1350 2482 1356 2483
rect 1462 2487 1468 2488
rect 1462 2483 1463 2487
rect 1467 2483 1468 2487
rect 1462 2482 1468 2483
rect 1574 2487 1580 2488
rect 1574 2483 1575 2487
rect 1579 2483 1580 2487
rect 1574 2482 1580 2483
rect 1670 2487 1676 2488
rect 1670 2483 1671 2487
rect 1675 2483 1676 2487
rect 1766 2484 1767 2488
rect 1771 2484 1772 2488
rect 1766 2483 1772 2484
rect 1670 2482 1676 2483
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 1766 2471 1772 2472
rect 110 2466 116 2467
rect 134 2468 140 2469
rect 134 2464 135 2468
rect 139 2464 140 2468
rect 134 2463 140 2464
rect 246 2468 252 2469
rect 246 2464 247 2468
rect 251 2464 252 2468
rect 246 2463 252 2464
rect 390 2468 396 2469
rect 390 2464 391 2468
rect 395 2464 396 2468
rect 390 2463 396 2464
rect 542 2468 548 2469
rect 542 2464 543 2468
rect 547 2464 548 2468
rect 542 2463 548 2464
rect 694 2468 700 2469
rect 694 2464 695 2468
rect 699 2464 700 2468
rect 694 2463 700 2464
rect 838 2468 844 2469
rect 838 2464 839 2468
rect 843 2464 844 2468
rect 838 2463 844 2464
rect 974 2468 980 2469
rect 974 2464 975 2468
rect 979 2464 980 2468
rect 974 2463 980 2464
rect 1102 2468 1108 2469
rect 1102 2464 1103 2468
rect 1107 2464 1108 2468
rect 1102 2463 1108 2464
rect 1230 2468 1236 2469
rect 1230 2464 1231 2468
rect 1235 2464 1236 2468
rect 1230 2463 1236 2464
rect 1350 2468 1356 2469
rect 1350 2464 1351 2468
rect 1355 2464 1356 2468
rect 1350 2463 1356 2464
rect 1462 2468 1468 2469
rect 1462 2464 1463 2468
rect 1467 2464 1468 2468
rect 1462 2463 1468 2464
rect 1574 2468 1580 2469
rect 1574 2464 1575 2468
rect 1579 2464 1580 2468
rect 1574 2463 1580 2464
rect 1670 2468 1676 2469
rect 1670 2464 1671 2468
rect 1675 2464 1676 2468
rect 1766 2467 1767 2471
rect 1771 2467 1772 2471
rect 1766 2466 1772 2467
rect 1670 2463 1676 2464
rect 2014 2460 2020 2461
rect 1806 2457 1812 2458
rect 1806 2453 1807 2457
rect 1811 2453 1812 2457
rect 2014 2456 2015 2460
rect 2019 2456 2020 2460
rect 2014 2455 2020 2456
rect 2198 2460 2204 2461
rect 2198 2456 2199 2460
rect 2203 2456 2204 2460
rect 2198 2455 2204 2456
rect 2366 2460 2372 2461
rect 2366 2456 2367 2460
rect 2371 2456 2372 2460
rect 2366 2455 2372 2456
rect 2526 2460 2532 2461
rect 2526 2456 2527 2460
rect 2531 2456 2532 2460
rect 2526 2455 2532 2456
rect 2670 2460 2676 2461
rect 2670 2456 2671 2460
rect 2675 2456 2676 2460
rect 2670 2455 2676 2456
rect 2806 2460 2812 2461
rect 2806 2456 2807 2460
rect 2811 2456 2812 2460
rect 2806 2455 2812 2456
rect 2926 2460 2932 2461
rect 2926 2456 2927 2460
rect 2931 2456 2932 2460
rect 2926 2455 2932 2456
rect 3046 2460 3052 2461
rect 3046 2456 3047 2460
rect 3051 2456 3052 2460
rect 3046 2455 3052 2456
rect 3158 2460 3164 2461
rect 3158 2456 3159 2460
rect 3163 2456 3164 2460
rect 3158 2455 3164 2456
rect 3270 2460 3276 2461
rect 3270 2456 3271 2460
rect 3275 2456 3276 2460
rect 3270 2455 3276 2456
rect 3366 2460 3372 2461
rect 3366 2456 3367 2460
rect 3371 2456 3372 2460
rect 3366 2455 3372 2456
rect 3462 2457 3468 2458
rect 1806 2452 1812 2453
rect 3462 2453 3463 2457
rect 3467 2453 3468 2457
rect 3462 2452 3468 2453
rect 2014 2441 2020 2442
rect 1806 2440 1812 2441
rect 1806 2436 1807 2440
rect 1811 2436 1812 2440
rect 2014 2437 2015 2441
rect 2019 2437 2020 2441
rect 2014 2436 2020 2437
rect 2198 2441 2204 2442
rect 2198 2437 2199 2441
rect 2203 2437 2204 2441
rect 2198 2436 2204 2437
rect 2366 2441 2372 2442
rect 2366 2437 2367 2441
rect 2371 2437 2372 2441
rect 2366 2436 2372 2437
rect 2526 2441 2532 2442
rect 2526 2437 2527 2441
rect 2531 2437 2532 2441
rect 2526 2436 2532 2437
rect 2670 2441 2676 2442
rect 2670 2437 2671 2441
rect 2675 2437 2676 2441
rect 2670 2436 2676 2437
rect 2806 2441 2812 2442
rect 2806 2437 2807 2441
rect 2811 2437 2812 2441
rect 2806 2436 2812 2437
rect 2926 2441 2932 2442
rect 2926 2437 2927 2441
rect 2931 2437 2932 2441
rect 2926 2436 2932 2437
rect 3046 2441 3052 2442
rect 3046 2437 3047 2441
rect 3051 2437 3052 2441
rect 3046 2436 3052 2437
rect 3158 2441 3164 2442
rect 3158 2437 3159 2441
rect 3163 2437 3164 2441
rect 3158 2436 3164 2437
rect 3270 2441 3276 2442
rect 3270 2437 3271 2441
rect 3275 2437 3276 2441
rect 3270 2436 3276 2437
rect 3366 2441 3372 2442
rect 3366 2437 3367 2441
rect 3371 2437 3372 2441
rect 3366 2436 3372 2437
rect 3462 2440 3468 2441
rect 3462 2436 3463 2440
rect 3467 2436 3468 2440
rect 1806 2435 1812 2436
rect 3462 2435 3468 2436
rect 134 2408 140 2409
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 134 2404 135 2408
rect 139 2404 140 2408
rect 134 2403 140 2404
rect 238 2408 244 2409
rect 238 2404 239 2408
rect 243 2404 244 2408
rect 238 2403 244 2404
rect 390 2408 396 2409
rect 390 2404 391 2408
rect 395 2404 396 2408
rect 390 2403 396 2404
rect 550 2408 556 2409
rect 550 2404 551 2408
rect 555 2404 556 2408
rect 550 2403 556 2404
rect 718 2408 724 2409
rect 718 2404 719 2408
rect 723 2404 724 2408
rect 718 2403 724 2404
rect 894 2408 900 2409
rect 894 2404 895 2408
rect 899 2404 900 2408
rect 894 2403 900 2404
rect 1062 2408 1068 2409
rect 1062 2404 1063 2408
rect 1067 2404 1068 2408
rect 1062 2403 1068 2404
rect 1238 2408 1244 2409
rect 1238 2404 1239 2408
rect 1243 2404 1244 2408
rect 1238 2403 1244 2404
rect 1414 2408 1420 2409
rect 1414 2404 1415 2408
rect 1419 2404 1420 2408
rect 1414 2403 1420 2404
rect 1590 2408 1596 2409
rect 1590 2404 1591 2408
rect 1595 2404 1596 2408
rect 1590 2403 1596 2404
rect 1766 2405 1772 2406
rect 110 2400 116 2401
rect 1766 2401 1767 2405
rect 1771 2401 1772 2405
rect 1766 2400 1772 2401
rect 1806 2392 1812 2393
rect 3462 2392 3468 2393
rect 134 2389 140 2390
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 134 2385 135 2389
rect 139 2385 140 2389
rect 134 2384 140 2385
rect 238 2389 244 2390
rect 238 2385 239 2389
rect 243 2385 244 2389
rect 238 2384 244 2385
rect 390 2389 396 2390
rect 390 2385 391 2389
rect 395 2385 396 2389
rect 390 2384 396 2385
rect 550 2389 556 2390
rect 550 2385 551 2389
rect 555 2385 556 2389
rect 550 2384 556 2385
rect 718 2389 724 2390
rect 718 2385 719 2389
rect 723 2385 724 2389
rect 718 2384 724 2385
rect 894 2389 900 2390
rect 894 2385 895 2389
rect 899 2385 900 2389
rect 894 2384 900 2385
rect 1062 2389 1068 2390
rect 1062 2385 1063 2389
rect 1067 2385 1068 2389
rect 1062 2384 1068 2385
rect 1238 2389 1244 2390
rect 1238 2385 1239 2389
rect 1243 2385 1244 2389
rect 1238 2384 1244 2385
rect 1414 2389 1420 2390
rect 1414 2385 1415 2389
rect 1419 2385 1420 2389
rect 1414 2384 1420 2385
rect 1590 2389 1596 2390
rect 1590 2385 1591 2389
rect 1595 2385 1596 2389
rect 1590 2384 1596 2385
rect 1766 2388 1772 2389
rect 1766 2384 1767 2388
rect 1771 2384 1772 2388
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1838 2391 1844 2392
rect 1838 2387 1839 2391
rect 1843 2387 1844 2391
rect 1838 2386 1844 2387
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2387 2012 2391
rect 2006 2386 2012 2387
rect 2182 2391 2188 2392
rect 2182 2387 2183 2391
rect 2187 2387 2188 2391
rect 2182 2386 2188 2387
rect 2366 2391 2372 2392
rect 2366 2387 2367 2391
rect 2371 2387 2372 2391
rect 2366 2386 2372 2387
rect 2558 2391 2564 2392
rect 2558 2387 2559 2391
rect 2563 2387 2564 2391
rect 2558 2386 2564 2387
rect 2758 2391 2764 2392
rect 2758 2387 2759 2391
rect 2763 2387 2764 2391
rect 2758 2386 2764 2387
rect 2966 2391 2972 2392
rect 2966 2387 2967 2391
rect 2971 2387 2972 2391
rect 2966 2386 2972 2387
rect 3174 2391 3180 2392
rect 3174 2387 3175 2391
rect 3179 2387 3180 2391
rect 3174 2386 3180 2387
rect 3366 2391 3372 2392
rect 3366 2387 3367 2391
rect 3371 2387 3372 2391
rect 3462 2388 3463 2392
rect 3467 2388 3468 2392
rect 3462 2387 3468 2388
rect 3366 2386 3372 2387
rect 110 2383 116 2384
rect 1766 2383 1772 2384
rect 1806 2375 1812 2376
rect 1806 2371 1807 2375
rect 1811 2371 1812 2375
rect 3462 2375 3468 2376
rect 1806 2370 1812 2371
rect 1838 2372 1844 2373
rect 1838 2368 1839 2372
rect 1843 2368 1844 2372
rect 1838 2367 1844 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2182 2372 2188 2373
rect 2182 2368 2183 2372
rect 2187 2368 2188 2372
rect 2182 2367 2188 2368
rect 2366 2372 2372 2373
rect 2366 2368 2367 2372
rect 2371 2368 2372 2372
rect 2366 2367 2372 2368
rect 2558 2372 2564 2373
rect 2558 2368 2559 2372
rect 2563 2368 2564 2372
rect 2558 2367 2564 2368
rect 2758 2372 2764 2373
rect 2758 2368 2759 2372
rect 2763 2368 2764 2372
rect 2758 2367 2764 2368
rect 2966 2372 2972 2373
rect 2966 2368 2967 2372
rect 2971 2368 2972 2372
rect 2966 2367 2972 2368
rect 3174 2372 3180 2373
rect 3174 2368 3175 2372
rect 3179 2368 3180 2372
rect 3174 2367 3180 2368
rect 3366 2372 3372 2373
rect 3366 2368 3367 2372
rect 3371 2368 3372 2372
rect 3462 2371 3463 2375
rect 3467 2371 3468 2375
rect 3462 2370 3468 2371
rect 3366 2367 3372 2368
rect 110 2336 116 2337
rect 1766 2336 1772 2337
rect 110 2332 111 2336
rect 115 2332 116 2336
rect 110 2331 116 2332
rect 374 2335 380 2336
rect 374 2331 375 2335
rect 379 2331 380 2335
rect 374 2330 380 2331
rect 478 2335 484 2336
rect 478 2331 479 2335
rect 483 2331 484 2335
rect 478 2330 484 2331
rect 598 2335 604 2336
rect 598 2331 599 2335
rect 603 2331 604 2335
rect 598 2330 604 2331
rect 718 2335 724 2336
rect 718 2331 719 2335
rect 723 2331 724 2335
rect 718 2330 724 2331
rect 846 2335 852 2336
rect 846 2331 847 2335
rect 851 2331 852 2335
rect 846 2330 852 2331
rect 974 2335 980 2336
rect 974 2331 975 2335
rect 979 2331 980 2335
rect 974 2330 980 2331
rect 1102 2335 1108 2336
rect 1102 2331 1103 2335
rect 1107 2331 1108 2335
rect 1102 2330 1108 2331
rect 1238 2335 1244 2336
rect 1238 2331 1239 2335
rect 1243 2331 1244 2335
rect 1238 2330 1244 2331
rect 1374 2335 1380 2336
rect 1374 2331 1375 2335
rect 1379 2331 1380 2335
rect 1374 2330 1380 2331
rect 1510 2335 1516 2336
rect 1510 2331 1511 2335
rect 1515 2331 1516 2335
rect 1766 2332 1767 2336
rect 1771 2332 1772 2336
rect 1766 2331 1772 2332
rect 1510 2330 1516 2331
rect 1886 2328 1892 2329
rect 1806 2325 1812 2326
rect 1806 2321 1807 2325
rect 1811 2321 1812 2325
rect 1886 2324 1887 2328
rect 1891 2324 1892 2328
rect 1886 2323 1892 2324
rect 2014 2328 2020 2329
rect 2014 2324 2015 2328
rect 2019 2324 2020 2328
rect 2014 2323 2020 2324
rect 2150 2328 2156 2329
rect 2150 2324 2151 2328
rect 2155 2324 2156 2328
rect 2150 2323 2156 2324
rect 2302 2328 2308 2329
rect 2302 2324 2303 2328
rect 2307 2324 2308 2328
rect 2302 2323 2308 2324
rect 2462 2328 2468 2329
rect 2462 2324 2463 2328
rect 2467 2324 2468 2328
rect 2462 2323 2468 2324
rect 2646 2328 2652 2329
rect 2646 2324 2647 2328
rect 2651 2324 2652 2328
rect 2646 2323 2652 2324
rect 2838 2328 2844 2329
rect 2838 2324 2839 2328
rect 2843 2324 2844 2328
rect 2838 2323 2844 2324
rect 3046 2328 3052 2329
rect 3046 2324 3047 2328
rect 3051 2324 3052 2328
rect 3046 2323 3052 2324
rect 3254 2328 3260 2329
rect 3254 2324 3255 2328
rect 3259 2324 3260 2328
rect 3254 2323 3260 2324
rect 3462 2325 3468 2326
rect 1806 2320 1812 2321
rect 3462 2321 3463 2325
rect 3467 2321 3468 2325
rect 3462 2320 3468 2321
rect 110 2319 116 2320
rect 110 2315 111 2319
rect 115 2315 116 2319
rect 1766 2319 1772 2320
rect 110 2314 116 2315
rect 374 2316 380 2317
rect 374 2312 375 2316
rect 379 2312 380 2316
rect 374 2311 380 2312
rect 478 2316 484 2317
rect 478 2312 479 2316
rect 483 2312 484 2316
rect 478 2311 484 2312
rect 598 2316 604 2317
rect 598 2312 599 2316
rect 603 2312 604 2316
rect 598 2311 604 2312
rect 718 2316 724 2317
rect 718 2312 719 2316
rect 723 2312 724 2316
rect 718 2311 724 2312
rect 846 2316 852 2317
rect 846 2312 847 2316
rect 851 2312 852 2316
rect 846 2311 852 2312
rect 974 2316 980 2317
rect 974 2312 975 2316
rect 979 2312 980 2316
rect 974 2311 980 2312
rect 1102 2316 1108 2317
rect 1102 2312 1103 2316
rect 1107 2312 1108 2316
rect 1102 2311 1108 2312
rect 1238 2316 1244 2317
rect 1238 2312 1239 2316
rect 1243 2312 1244 2316
rect 1238 2311 1244 2312
rect 1374 2316 1380 2317
rect 1374 2312 1375 2316
rect 1379 2312 1380 2316
rect 1374 2311 1380 2312
rect 1510 2316 1516 2317
rect 1510 2312 1511 2316
rect 1515 2312 1516 2316
rect 1766 2315 1767 2319
rect 1771 2315 1772 2319
rect 1766 2314 1772 2315
rect 1510 2311 1516 2312
rect 1886 2309 1892 2310
rect 1806 2308 1812 2309
rect 1806 2304 1807 2308
rect 1811 2304 1812 2308
rect 1886 2305 1887 2309
rect 1891 2305 1892 2309
rect 1886 2304 1892 2305
rect 2014 2309 2020 2310
rect 2014 2305 2015 2309
rect 2019 2305 2020 2309
rect 2014 2304 2020 2305
rect 2150 2309 2156 2310
rect 2150 2305 2151 2309
rect 2155 2305 2156 2309
rect 2150 2304 2156 2305
rect 2302 2309 2308 2310
rect 2302 2305 2303 2309
rect 2307 2305 2308 2309
rect 2302 2304 2308 2305
rect 2462 2309 2468 2310
rect 2462 2305 2463 2309
rect 2467 2305 2468 2309
rect 2462 2304 2468 2305
rect 2646 2309 2652 2310
rect 2646 2305 2647 2309
rect 2651 2305 2652 2309
rect 2646 2304 2652 2305
rect 2838 2309 2844 2310
rect 2838 2305 2839 2309
rect 2843 2305 2844 2309
rect 2838 2304 2844 2305
rect 3046 2309 3052 2310
rect 3046 2305 3047 2309
rect 3051 2305 3052 2309
rect 3046 2304 3052 2305
rect 3254 2309 3260 2310
rect 3254 2305 3255 2309
rect 3259 2305 3260 2309
rect 3254 2304 3260 2305
rect 3462 2308 3468 2309
rect 3462 2304 3463 2308
rect 3467 2304 3468 2308
rect 1806 2303 1812 2304
rect 3462 2303 3468 2304
rect 574 2264 580 2265
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 574 2260 575 2264
rect 579 2260 580 2264
rect 574 2259 580 2260
rect 662 2264 668 2265
rect 662 2260 663 2264
rect 667 2260 668 2264
rect 662 2259 668 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 862 2264 868 2265
rect 862 2260 863 2264
rect 867 2260 868 2264
rect 862 2259 868 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1078 2264 1084 2265
rect 1078 2260 1079 2264
rect 1083 2260 1084 2264
rect 1078 2259 1084 2260
rect 1190 2264 1196 2265
rect 1190 2260 1191 2264
rect 1195 2260 1196 2264
rect 1190 2259 1196 2260
rect 1302 2264 1308 2265
rect 1302 2260 1303 2264
rect 1307 2260 1308 2264
rect 1302 2259 1308 2260
rect 1414 2264 1420 2265
rect 1414 2260 1415 2264
rect 1419 2260 1420 2264
rect 1414 2259 1420 2260
rect 1766 2261 1772 2262
rect 110 2256 116 2257
rect 1766 2257 1767 2261
rect 1771 2257 1772 2261
rect 1766 2256 1772 2257
rect 1806 2260 1812 2261
rect 3462 2260 3468 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1806 2255 1812 2256
rect 2038 2259 2044 2260
rect 2038 2255 2039 2259
rect 2043 2255 2044 2259
rect 2038 2254 2044 2255
rect 2134 2259 2140 2260
rect 2134 2255 2135 2259
rect 2139 2255 2140 2259
rect 2134 2254 2140 2255
rect 2238 2259 2244 2260
rect 2238 2255 2239 2259
rect 2243 2255 2244 2259
rect 2238 2254 2244 2255
rect 2342 2259 2348 2260
rect 2342 2255 2343 2259
rect 2347 2255 2348 2259
rect 2342 2254 2348 2255
rect 2462 2259 2468 2260
rect 2462 2255 2463 2259
rect 2467 2255 2468 2259
rect 2462 2254 2468 2255
rect 2590 2259 2596 2260
rect 2590 2255 2591 2259
rect 2595 2255 2596 2259
rect 2590 2254 2596 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2886 2259 2892 2260
rect 2886 2255 2887 2259
rect 2891 2255 2892 2259
rect 2886 2254 2892 2255
rect 3046 2259 3052 2260
rect 3046 2255 3047 2259
rect 3051 2255 3052 2259
rect 3046 2254 3052 2255
rect 3214 2259 3220 2260
rect 3214 2255 3215 2259
rect 3219 2255 3220 2259
rect 3214 2254 3220 2255
rect 3366 2259 3372 2260
rect 3366 2255 3367 2259
rect 3371 2255 3372 2259
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 3462 2255 3468 2256
rect 3366 2254 3372 2255
rect 574 2245 580 2246
rect 110 2244 116 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 574 2241 575 2245
rect 579 2241 580 2245
rect 574 2240 580 2241
rect 662 2245 668 2246
rect 662 2241 663 2245
rect 667 2241 668 2245
rect 662 2240 668 2241
rect 758 2245 764 2246
rect 758 2241 759 2245
rect 763 2241 764 2245
rect 758 2240 764 2241
rect 862 2245 868 2246
rect 862 2241 863 2245
rect 867 2241 868 2245
rect 862 2240 868 2241
rect 966 2245 972 2246
rect 966 2241 967 2245
rect 971 2241 972 2245
rect 966 2240 972 2241
rect 1078 2245 1084 2246
rect 1078 2241 1079 2245
rect 1083 2241 1084 2245
rect 1078 2240 1084 2241
rect 1190 2245 1196 2246
rect 1190 2241 1191 2245
rect 1195 2241 1196 2245
rect 1190 2240 1196 2241
rect 1302 2245 1308 2246
rect 1302 2241 1303 2245
rect 1307 2241 1308 2245
rect 1302 2240 1308 2241
rect 1414 2245 1420 2246
rect 1414 2241 1415 2245
rect 1419 2241 1420 2245
rect 1414 2240 1420 2241
rect 1766 2244 1772 2245
rect 1766 2240 1767 2244
rect 1771 2240 1772 2244
rect 110 2239 116 2240
rect 1766 2239 1772 2240
rect 1806 2243 1812 2244
rect 1806 2239 1807 2243
rect 1811 2239 1812 2243
rect 3462 2243 3468 2244
rect 1806 2238 1812 2239
rect 2038 2240 2044 2241
rect 2038 2236 2039 2240
rect 2043 2236 2044 2240
rect 2038 2235 2044 2236
rect 2134 2240 2140 2241
rect 2134 2236 2135 2240
rect 2139 2236 2140 2240
rect 2134 2235 2140 2236
rect 2238 2240 2244 2241
rect 2238 2236 2239 2240
rect 2243 2236 2244 2240
rect 2238 2235 2244 2236
rect 2342 2240 2348 2241
rect 2342 2236 2343 2240
rect 2347 2236 2348 2240
rect 2342 2235 2348 2236
rect 2462 2240 2468 2241
rect 2462 2236 2463 2240
rect 2467 2236 2468 2240
rect 2462 2235 2468 2236
rect 2590 2240 2596 2241
rect 2590 2236 2591 2240
rect 2595 2236 2596 2240
rect 2590 2235 2596 2236
rect 2734 2240 2740 2241
rect 2734 2236 2735 2240
rect 2739 2236 2740 2240
rect 2734 2235 2740 2236
rect 2886 2240 2892 2241
rect 2886 2236 2887 2240
rect 2891 2236 2892 2240
rect 2886 2235 2892 2236
rect 3046 2240 3052 2241
rect 3046 2236 3047 2240
rect 3051 2236 3052 2240
rect 3046 2235 3052 2236
rect 3214 2240 3220 2241
rect 3214 2236 3215 2240
rect 3219 2236 3220 2240
rect 3214 2235 3220 2236
rect 3366 2240 3372 2241
rect 3366 2236 3367 2240
rect 3371 2236 3372 2240
rect 3462 2239 3463 2243
rect 3467 2239 3468 2243
rect 3462 2238 3468 2239
rect 3366 2235 3372 2236
rect 110 2200 116 2201
rect 1766 2200 1772 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 438 2199 444 2200
rect 438 2195 439 2199
rect 443 2195 444 2199
rect 438 2194 444 2195
rect 526 2199 532 2200
rect 526 2195 527 2199
rect 531 2195 532 2199
rect 526 2194 532 2195
rect 614 2199 620 2200
rect 614 2195 615 2199
rect 619 2195 620 2199
rect 614 2194 620 2195
rect 702 2199 708 2200
rect 702 2195 703 2199
rect 707 2195 708 2199
rect 702 2194 708 2195
rect 790 2199 796 2200
rect 790 2195 791 2199
rect 795 2195 796 2199
rect 790 2194 796 2195
rect 878 2199 884 2200
rect 878 2195 879 2199
rect 883 2195 884 2199
rect 878 2194 884 2195
rect 966 2199 972 2200
rect 966 2195 967 2199
rect 971 2195 972 2199
rect 966 2194 972 2195
rect 1054 2199 1060 2200
rect 1054 2195 1055 2199
rect 1059 2195 1060 2199
rect 1054 2194 1060 2195
rect 1142 2199 1148 2200
rect 1142 2195 1143 2199
rect 1147 2195 1148 2199
rect 1142 2194 1148 2195
rect 1230 2199 1236 2200
rect 1230 2195 1231 2199
rect 1235 2195 1236 2199
rect 1230 2194 1236 2195
rect 1318 2199 1324 2200
rect 1318 2195 1319 2199
rect 1323 2195 1324 2199
rect 1766 2196 1767 2200
rect 1771 2196 1772 2200
rect 1766 2195 1772 2196
rect 1318 2194 1324 2195
rect 2182 2184 2188 2185
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 1766 2183 1772 2184
rect 110 2178 116 2179
rect 438 2180 444 2181
rect 438 2176 439 2180
rect 443 2176 444 2180
rect 438 2175 444 2176
rect 526 2180 532 2181
rect 526 2176 527 2180
rect 531 2176 532 2180
rect 526 2175 532 2176
rect 614 2180 620 2181
rect 614 2176 615 2180
rect 619 2176 620 2180
rect 614 2175 620 2176
rect 702 2180 708 2181
rect 702 2176 703 2180
rect 707 2176 708 2180
rect 702 2175 708 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 878 2180 884 2181
rect 878 2176 879 2180
rect 883 2176 884 2180
rect 878 2175 884 2176
rect 966 2180 972 2181
rect 966 2176 967 2180
rect 971 2176 972 2180
rect 966 2175 972 2176
rect 1054 2180 1060 2181
rect 1054 2176 1055 2180
rect 1059 2176 1060 2180
rect 1054 2175 1060 2176
rect 1142 2180 1148 2181
rect 1142 2176 1143 2180
rect 1147 2176 1148 2180
rect 1142 2175 1148 2176
rect 1230 2180 1236 2181
rect 1230 2176 1231 2180
rect 1235 2176 1236 2180
rect 1230 2175 1236 2176
rect 1318 2180 1324 2181
rect 1318 2176 1319 2180
rect 1323 2176 1324 2180
rect 1766 2179 1767 2183
rect 1771 2179 1772 2183
rect 1766 2178 1772 2179
rect 1806 2181 1812 2182
rect 1806 2177 1807 2181
rect 1811 2177 1812 2181
rect 2182 2180 2183 2184
rect 2187 2180 2188 2184
rect 2182 2179 2188 2180
rect 2278 2184 2284 2185
rect 2278 2180 2279 2184
rect 2283 2180 2284 2184
rect 2278 2179 2284 2180
rect 2382 2184 2388 2185
rect 2382 2180 2383 2184
rect 2387 2180 2388 2184
rect 2382 2179 2388 2180
rect 2494 2184 2500 2185
rect 2494 2180 2495 2184
rect 2499 2180 2500 2184
rect 2494 2179 2500 2180
rect 2606 2184 2612 2185
rect 2606 2180 2607 2184
rect 2611 2180 2612 2184
rect 2606 2179 2612 2180
rect 2718 2184 2724 2185
rect 2718 2180 2719 2184
rect 2723 2180 2724 2184
rect 2718 2179 2724 2180
rect 2838 2184 2844 2185
rect 2838 2180 2839 2184
rect 2843 2180 2844 2184
rect 2838 2179 2844 2180
rect 2966 2184 2972 2185
rect 2966 2180 2967 2184
rect 2971 2180 2972 2184
rect 2966 2179 2972 2180
rect 3102 2184 3108 2185
rect 3102 2180 3103 2184
rect 3107 2180 3108 2184
rect 3102 2179 3108 2180
rect 3246 2184 3252 2185
rect 3246 2180 3247 2184
rect 3251 2180 3252 2184
rect 3246 2179 3252 2180
rect 3366 2184 3372 2185
rect 3366 2180 3367 2184
rect 3371 2180 3372 2184
rect 3366 2179 3372 2180
rect 3462 2181 3468 2182
rect 1806 2176 1812 2177
rect 3462 2177 3463 2181
rect 3467 2177 3468 2181
rect 3462 2176 3468 2177
rect 1318 2175 1324 2176
rect 2182 2165 2188 2166
rect 1806 2164 1812 2165
rect 1806 2160 1807 2164
rect 1811 2160 1812 2164
rect 2182 2161 2183 2165
rect 2187 2161 2188 2165
rect 2182 2160 2188 2161
rect 2278 2165 2284 2166
rect 2278 2161 2279 2165
rect 2283 2161 2284 2165
rect 2278 2160 2284 2161
rect 2382 2165 2388 2166
rect 2382 2161 2383 2165
rect 2387 2161 2388 2165
rect 2382 2160 2388 2161
rect 2494 2165 2500 2166
rect 2494 2161 2495 2165
rect 2499 2161 2500 2165
rect 2494 2160 2500 2161
rect 2606 2165 2612 2166
rect 2606 2161 2607 2165
rect 2611 2161 2612 2165
rect 2606 2160 2612 2161
rect 2718 2165 2724 2166
rect 2718 2161 2719 2165
rect 2723 2161 2724 2165
rect 2718 2160 2724 2161
rect 2838 2165 2844 2166
rect 2838 2161 2839 2165
rect 2843 2161 2844 2165
rect 2838 2160 2844 2161
rect 2966 2165 2972 2166
rect 2966 2161 2967 2165
rect 2971 2161 2972 2165
rect 2966 2160 2972 2161
rect 3102 2165 3108 2166
rect 3102 2161 3103 2165
rect 3107 2161 3108 2165
rect 3102 2160 3108 2161
rect 3246 2165 3252 2166
rect 3246 2161 3247 2165
rect 3251 2161 3252 2165
rect 3246 2160 3252 2161
rect 3366 2165 3372 2166
rect 3366 2161 3367 2165
rect 3371 2161 3372 2165
rect 3366 2160 3372 2161
rect 3462 2164 3468 2165
rect 3462 2160 3463 2164
rect 3467 2160 3468 2164
rect 1806 2159 1812 2160
rect 3462 2159 3468 2160
rect 302 2120 308 2121
rect 110 2117 116 2118
rect 110 2113 111 2117
rect 115 2113 116 2117
rect 302 2116 303 2120
rect 307 2116 308 2120
rect 302 2115 308 2116
rect 406 2120 412 2121
rect 406 2116 407 2120
rect 411 2116 412 2120
rect 406 2115 412 2116
rect 518 2120 524 2121
rect 518 2116 519 2120
rect 523 2116 524 2120
rect 518 2115 524 2116
rect 630 2120 636 2121
rect 630 2116 631 2120
rect 635 2116 636 2120
rect 630 2115 636 2116
rect 742 2120 748 2121
rect 742 2116 743 2120
rect 747 2116 748 2120
rect 742 2115 748 2116
rect 862 2120 868 2121
rect 862 2116 863 2120
rect 867 2116 868 2120
rect 862 2115 868 2116
rect 982 2120 988 2121
rect 982 2116 983 2120
rect 987 2116 988 2120
rect 982 2115 988 2116
rect 1766 2117 1772 2118
rect 110 2112 116 2113
rect 1766 2113 1767 2117
rect 1771 2113 1772 2117
rect 1766 2112 1772 2113
rect 1806 2112 1812 2113
rect 3462 2112 3468 2113
rect 1806 2108 1807 2112
rect 1811 2108 1812 2112
rect 1806 2107 1812 2108
rect 2134 2111 2140 2112
rect 2134 2107 2135 2111
rect 2139 2107 2140 2111
rect 2134 2106 2140 2107
rect 2254 2111 2260 2112
rect 2254 2107 2255 2111
rect 2259 2107 2260 2111
rect 2254 2106 2260 2107
rect 2382 2111 2388 2112
rect 2382 2107 2383 2111
rect 2387 2107 2388 2111
rect 2382 2106 2388 2107
rect 2518 2111 2524 2112
rect 2518 2107 2519 2111
rect 2523 2107 2524 2111
rect 2518 2106 2524 2107
rect 2654 2111 2660 2112
rect 2654 2107 2655 2111
rect 2659 2107 2660 2111
rect 2654 2106 2660 2107
rect 2782 2111 2788 2112
rect 2782 2107 2783 2111
rect 2787 2107 2788 2111
rect 2782 2106 2788 2107
rect 2910 2111 2916 2112
rect 2910 2107 2911 2111
rect 2915 2107 2916 2111
rect 2910 2106 2916 2107
rect 3030 2111 3036 2112
rect 3030 2107 3031 2111
rect 3035 2107 3036 2111
rect 3030 2106 3036 2107
rect 3150 2111 3156 2112
rect 3150 2107 3151 2111
rect 3155 2107 3156 2111
rect 3150 2106 3156 2107
rect 3270 2111 3276 2112
rect 3270 2107 3271 2111
rect 3275 2107 3276 2111
rect 3270 2106 3276 2107
rect 3366 2111 3372 2112
rect 3366 2107 3367 2111
rect 3371 2107 3372 2111
rect 3462 2108 3463 2112
rect 3467 2108 3468 2112
rect 3462 2107 3468 2108
rect 3366 2106 3372 2107
rect 302 2101 308 2102
rect 110 2100 116 2101
rect 110 2096 111 2100
rect 115 2096 116 2100
rect 302 2097 303 2101
rect 307 2097 308 2101
rect 302 2096 308 2097
rect 406 2101 412 2102
rect 406 2097 407 2101
rect 411 2097 412 2101
rect 406 2096 412 2097
rect 518 2101 524 2102
rect 518 2097 519 2101
rect 523 2097 524 2101
rect 518 2096 524 2097
rect 630 2101 636 2102
rect 630 2097 631 2101
rect 635 2097 636 2101
rect 630 2096 636 2097
rect 742 2101 748 2102
rect 742 2097 743 2101
rect 747 2097 748 2101
rect 742 2096 748 2097
rect 862 2101 868 2102
rect 862 2097 863 2101
rect 867 2097 868 2101
rect 862 2096 868 2097
rect 982 2101 988 2102
rect 982 2097 983 2101
rect 987 2097 988 2101
rect 982 2096 988 2097
rect 1766 2100 1772 2101
rect 1766 2096 1767 2100
rect 1771 2096 1772 2100
rect 110 2095 116 2096
rect 1766 2095 1772 2096
rect 1806 2095 1812 2096
rect 1806 2091 1807 2095
rect 1811 2091 1812 2095
rect 3462 2095 3468 2096
rect 1806 2090 1812 2091
rect 2134 2092 2140 2093
rect 2134 2088 2135 2092
rect 2139 2088 2140 2092
rect 2134 2087 2140 2088
rect 2254 2092 2260 2093
rect 2254 2088 2255 2092
rect 2259 2088 2260 2092
rect 2254 2087 2260 2088
rect 2382 2092 2388 2093
rect 2382 2088 2383 2092
rect 2387 2088 2388 2092
rect 2382 2087 2388 2088
rect 2518 2092 2524 2093
rect 2518 2088 2519 2092
rect 2523 2088 2524 2092
rect 2518 2087 2524 2088
rect 2654 2092 2660 2093
rect 2654 2088 2655 2092
rect 2659 2088 2660 2092
rect 2654 2087 2660 2088
rect 2782 2092 2788 2093
rect 2782 2088 2783 2092
rect 2787 2088 2788 2092
rect 2782 2087 2788 2088
rect 2910 2092 2916 2093
rect 2910 2088 2911 2092
rect 2915 2088 2916 2092
rect 2910 2087 2916 2088
rect 3030 2092 3036 2093
rect 3030 2088 3031 2092
rect 3035 2088 3036 2092
rect 3030 2087 3036 2088
rect 3150 2092 3156 2093
rect 3150 2088 3151 2092
rect 3155 2088 3156 2092
rect 3150 2087 3156 2088
rect 3270 2092 3276 2093
rect 3270 2088 3271 2092
rect 3275 2088 3276 2092
rect 3270 2087 3276 2088
rect 3366 2092 3372 2093
rect 3366 2088 3367 2092
rect 3371 2088 3372 2092
rect 3462 2091 3463 2095
rect 3467 2091 3468 2095
rect 3462 2090 3468 2091
rect 3366 2087 3372 2088
rect 110 2056 116 2057
rect 1766 2056 1772 2057
rect 110 2052 111 2056
rect 115 2052 116 2056
rect 110 2051 116 2052
rect 254 2055 260 2056
rect 254 2051 255 2055
rect 259 2051 260 2055
rect 254 2050 260 2051
rect 374 2055 380 2056
rect 374 2051 375 2055
rect 379 2051 380 2055
rect 374 2050 380 2051
rect 494 2055 500 2056
rect 494 2051 495 2055
rect 499 2051 500 2055
rect 494 2050 500 2051
rect 614 2055 620 2056
rect 614 2051 615 2055
rect 619 2051 620 2055
rect 614 2050 620 2051
rect 726 2055 732 2056
rect 726 2051 727 2055
rect 731 2051 732 2055
rect 726 2050 732 2051
rect 830 2055 836 2056
rect 830 2051 831 2055
rect 835 2051 836 2055
rect 830 2050 836 2051
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 1254 2055 1260 2056
rect 1254 2051 1255 2055
rect 1259 2051 1260 2055
rect 1766 2052 1767 2056
rect 1771 2052 1772 2056
rect 1766 2051 1772 2052
rect 1254 2050 1260 2051
rect 2246 2040 2252 2041
rect 110 2039 116 2040
rect 110 2035 111 2039
rect 115 2035 116 2039
rect 1766 2039 1772 2040
rect 110 2034 116 2035
rect 254 2036 260 2037
rect 254 2032 255 2036
rect 259 2032 260 2036
rect 254 2031 260 2032
rect 374 2036 380 2037
rect 374 2032 375 2036
rect 379 2032 380 2036
rect 374 2031 380 2032
rect 494 2036 500 2037
rect 494 2032 495 2036
rect 499 2032 500 2036
rect 494 2031 500 2032
rect 614 2036 620 2037
rect 614 2032 615 2036
rect 619 2032 620 2036
rect 614 2031 620 2032
rect 726 2036 732 2037
rect 726 2032 727 2036
rect 731 2032 732 2036
rect 726 2031 732 2032
rect 830 2036 836 2037
rect 830 2032 831 2036
rect 835 2032 836 2036
rect 830 2031 836 2032
rect 934 2036 940 2037
rect 934 2032 935 2036
rect 939 2032 940 2036
rect 934 2031 940 2032
rect 1038 2036 1044 2037
rect 1038 2032 1039 2036
rect 1043 2032 1044 2036
rect 1038 2031 1044 2032
rect 1142 2036 1148 2037
rect 1142 2032 1143 2036
rect 1147 2032 1148 2036
rect 1142 2031 1148 2032
rect 1254 2036 1260 2037
rect 1254 2032 1255 2036
rect 1259 2032 1260 2036
rect 1766 2035 1767 2039
rect 1771 2035 1772 2039
rect 1766 2034 1772 2035
rect 1806 2037 1812 2038
rect 1806 2033 1807 2037
rect 1811 2033 1812 2037
rect 2246 2036 2247 2040
rect 2251 2036 2252 2040
rect 2246 2035 2252 2036
rect 2414 2040 2420 2041
rect 2414 2036 2415 2040
rect 2419 2036 2420 2040
rect 2414 2035 2420 2036
rect 2574 2040 2580 2041
rect 2574 2036 2575 2040
rect 2579 2036 2580 2040
rect 2574 2035 2580 2036
rect 2726 2040 2732 2041
rect 2726 2036 2727 2040
rect 2731 2036 2732 2040
rect 2726 2035 2732 2036
rect 2870 2040 2876 2041
rect 2870 2036 2871 2040
rect 2875 2036 2876 2040
rect 2870 2035 2876 2036
rect 3006 2040 3012 2041
rect 3006 2036 3007 2040
rect 3011 2036 3012 2040
rect 3006 2035 3012 2036
rect 3134 2040 3140 2041
rect 3134 2036 3135 2040
rect 3139 2036 3140 2040
rect 3134 2035 3140 2036
rect 3262 2040 3268 2041
rect 3262 2036 3263 2040
rect 3267 2036 3268 2040
rect 3262 2035 3268 2036
rect 3366 2040 3372 2041
rect 3366 2036 3367 2040
rect 3371 2036 3372 2040
rect 3366 2035 3372 2036
rect 3462 2037 3468 2038
rect 1806 2032 1812 2033
rect 3462 2033 3463 2037
rect 3467 2033 3468 2037
rect 3462 2032 3468 2033
rect 1254 2031 1260 2032
rect 2246 2021 2252 2022
rect 1806 2020 1812 2021
rect 1806 2016 1807 2020
rect 1811 2016 1812 2020
rect 2246 2017 2247 2021
rect 2251 2017 2252 2021
rect 2246 2016 2252 2017
rect 2414 2021 2420 2022
rect 2414 2017 2415 2021
rect 2419 2017 2420 2021
rect 2414 2016 2420 2017
rect 2574 2021 2580 2022
rect 2574 2017 2575 2021
rect 2579 2017 2580 2021
rect 2574 2016 2580 2017
rect 2726 2021 2732 2022
rect 2726 2017 2727 2021
rect 2731 2017 2732 2021
rect 2726 2016 2732 2017
rect 2870 2021 2876 2022
rect 2870 2017 2871 2021
rect 2875 2017 2876 2021
rect 2870 2016 2876 2017
rect 3006 2021 3012 2022
rect 3006 2017 3007 2021
rect 3011 2017 3012 2021
rect 3006 2016 3012 2017
rect 3134 2021 3140 2022
rect 3134 2017 3135 2021
rect 3139 2017 3140 2021
rect 3134 2016 3140 2017
rect 3262 2021 3268 2022
rect 3262 2017 3263 2021
rect 3267 2017 3268 2021
rect 3262 2016 3268 2017
rect 3366 2021 3372 2022
rect 3366 2017 3367 2021
rect 3371 2017 3372 2021
rect 3366 2016 3372 2017
rect 3462 2020 3468 2021
rect 3462 2016 3463 2020
rect 3467 2016 3468 2020
rect 1806 2015 1812 2016
rect 3462 2015 3468 2016
rect 358 1992 364 1993
rect 110 1989 116 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 358 1988 359 1992
rect 363 1988 364 1992
rect 358 1987 364 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 622 1992 628 1993
rect 622 1988 623 1992
rect 627 1988 628 1992
rect 622 1987 628 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 894 1992 900 1993
rect 894 1988 895 1992
rect 899 1988 900 1992
rect 894 1987 900 1988
rect 1022 1992 1028 1993
rect 1022 1988 1023 1992
rect 1027 1988 1028 1992
rect 1022 1987 1028 1988
rect 1150 1992 1156 1993
rect 1150 1988 1151 1992
rect 1155 1988 1156 1992
rect 1150 1987 1156 1988
rect 1270 1992 1276 1993
rect 1270 1988 1271 1992
rect 1275 1988 1276 1992
rect 1270 1987 1276 1988
rect 1398 1992 1404 1993
rect 1398 1988 1399 1992
rect 1403 1988 1404 1992
rect 1398 1987 1404 1988
rect 1526 1992 1532 1993
rect 1526 1988 1527 1992
rect 1531 1988 1532 1992
rect 1526 1987 1532 1988
rect 1766 1989 1772 1990
rect 110 1984 116 1985
rect 1766 1985 1767 1989
rect 1771 1985 1772 1989
rect 1766 1984 1772 1985
rect 358 1973 364 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 358 1969 359 1973
rect 363 1969 364 1973
rect 358 1968 364 1969
rect 486 1973 492 1974
rect 486 1969 487 1973
rect 491 1969 492 1973
rect 486 1968 492 1969
rect 622 1973 628 1974
rect 622 1969 623 1973
rect 627 1969 628 1973
rect 622 1968 628 1969
rect 758 1973 764 1974
rect 758 1969 759 1973
rect 763 1969 764 1973
rect 758 1968 764 1969
rect 894 1973 900 1974
rect 894 1969 895 1973
rect 899 1969 900 1973
rect 894 1968 900 1969
rect 1022 1973 1028 1974
rect 1022 1969 1023 1973
rect 1027 1969 1028 1973
rect 1022 1968 1028 1969
rect 1150 1973 1156 1974
rect 1150 1969 1151 1973
rect 1155 1969 1156 1973
rect 1150 1968 1156 1969
rect 1270 1973 1276 1974
rect 1270 1969 1271 1973
rect 1275 1969 1276 1973
rect 1270 1968 1276 1969
rect 1398 1973 1404 1974
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1526 1973 1532 1974
rect 1526 1969 1527 1973
rect 1531 1969 1532 1973
rect 1526 1968 1532 1969
rect 1766 1972 1772 1973
rect 1766 1968 1767 1972
rect 1771 1968 1772 1972
rect 110 1967 116 1968
rect 1766 1967 1772 1968
rect 1806 1960 1812 1961
rect 3462 1960 3468 1961
rect 1806 1956 1807 1960
rect 1811 1956 1812 1960
rect 1806 1955 1812 1956
rect 1830 1959 1836 1960
rect 1830 1955 1831 1959
rect 1835 1955 1836 1959
rect 1830 1954 1836 1955
rect 1918 1959 1924 1960
rect 1918 1955 1919 1959
rect 1923 1955 1924 1959
rect 1918 1954 1924 1955
rect 2046 1959 2052 1960
rect 2046 1955 2047 1959
rect 2051 1955 2052 1959
rect 2046 1954 2052 1955
rect 2182 1959 2188 1960
rect 2182 1955 2183 1959
rect 2187 1955 2188 1959
rect 2182 1954 2188 1955
rect 2326 1959 2332 1960
rect 2326 1955 2327 1959
rect 2331 1955 2332 1959
rect 2326 1954 2332 1955
rect 2470 1959 2476 1960
rect 2470 1955 2471 1959
rect 2475 1955 2476 1959
rect 2470 1954 2476 1955
rect 2614 1959 2620 1960
rect 2614 1955 2615 1959
rect 2619 1955 2620 1959
rect 2614 1954 2620 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2886 1959 2892 1960
rect 2886 1955 2887 1959
rect 2891 1955 2892 1959
rect 2886 1954 2892 1955
rect 3030 1959 3036 1960
rect 3030 1955 3031 1959
rect 3035 1955 3036 1959
rect 3030 1954 3036 1955
rect 3174 1959 3180 1960
rect 3174 1955 3175 1959
rect 3179 1955 3180 1959
rect 3174 1954 3180 1955
rect 3318 1959 3324 1960
rect 3318 1955 3319 1959
rect 3323 1955 3324 1959
rect 3462 1956 3463 1960
rect 3467 1956 3468 1960
rect 3462 1955 3468 1956
rect 3318 1954 3324 1955
rect 1806 1943 1812 1944
rect 1806 1939 1807 1943
rect 1811 1939 1812 1943
rect 3462 1943 3468 1944
rect 1806 1938 1812 1939
rect 1830 1940 1836 1941
rect 1830 1936 1831 1940
rect 1835 1936 1836 1940
rect 1830 1935 1836 1936
rect 1918 1940 1924 1941
rect 1918 1936 1919 1940
rect 1923 1936 1924 1940
rect 1918 1935 1924 1936
rect 2046 1940 2052 1941
rect 2046 1936 2047 1940
rect 2051 1936 2052 1940
rect 2046 1935 2052 1936
rect 2182 1940 2188 1941
rect 2182 1936 2183 1940
rect 2187 1936 2188 1940
rect 2182 1935 2188 1936
rect 2326 1940 2332 1941
rect 2326 1936 2327 1940
rect 2331 1936 2332 1940
rect 2326 1935 2332 1936
rect 2470 1940 2476 1941
rect 2470 1936 2471 1940
rect 2475 1936 2476 1940
rect 2470 1935 2476 1936
rect 2614 1940 2620 1941
rect 2614 1936 2615 1940
rect 2619 1936 2620 1940
rect 2614 1935 2620 1936
rect 2750 1940 2756 1941
rect 2750 1936 2751 1940
rect 2755 1936 2756 1940
rect 2750 1935 2756 1936
rect 2886 1940 2892 1941
rect 2886 1936 2887 1940
rect 2891 1936 2892 1940
rect 2886 1935 2892 1936
rect 3030 1940 3036 1941
rect 3030 1936 3031 1940
rect 3035 1936 3036 1940
rect 3030 1935 3036 1936
rect 3174 1940 3180 1941
rect 3174 1936 3175 1940
rect 3179 1936 3180 1940
rect 3174 1935 3180 1936
rect 3318 1940 3324 1941
rect 3318 1936 3319 1940
rect 3323 1936 3324 1940
rect 3462 1939 3463 1943
rect 3467 1939 3468 1943
rect 3462 1938 3468 1939
rect 3318 1935 3324 1936
rect 110 1928 116 1929
rect 1766 1928 1772 1929
rect 110 1924 111 1928
rect 115 1924 116 1928
rect 110 1923 116 1924
rect 446 1927 452 1928
rect 446 1923 447 1927
rect 451 1923 452 1927
rect 446 1922 452 1923
rect 574 1927 580 1928
rect 574 1923 575 1927
rect 579 1923 580 1927
rect 574 1922 580 1923
rect 710 1927 716 1928
rect 710 1923 711 1927
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 846 1927 852 1928
rect 846 1923 847 1927
rect 851 1923 852 1927
rect 846 1922 852 1923
rect 982 1927 988 1928
rect 982 1923 983 1927
rect 987 1923 988 1927
rect 982 1922 988 1923
rect 1118 1927 1124 1928
rect 1118 1923 1119 1927
rect 1123 1923 1124 1927
rect 1118 1922 1124 1923
rect 1254 1927 1260 1928
rect 1254 1923 1255 1927
rect 1259 1923 1260 1927
rect 1254 1922 1260 1923
rect 1382 1927 1388 1928
rect 1382 1923 1383 1927
rect 1387 1923 1388 1927
rect 1382 1922 1388 1923
rect 1518 1927 1524 1928
rect 1518 1923 1519 1927
rect 1523 1923 1524 1927
rect 1518 1922 1524 1923
rect 1654 1927 1660 1928
rect 1654 1923 1655 1927
rect 1659 1923 1660 1927
rect 1766 1924 1767 1928
rect 1771 1924 1772 1928
rect 1766 1923 1772 1924
rect 1654 1922 1660 1923
rect 110 1911 116 1912
rect 110 1907 111 1911
rect 115 1907 116 1911
rect 1766 1911 1772 1912
rect 110 1906 116 1907
rect 446 1908 452 1909
rect 446 1904 447 1908
rect 451 1904 452 1908
rect 446 1903 452 1904
rect 574 1908 580 1909
rect 574 1904 575 1908
rect 579 1904 580 1908
rect 574 1903 580 1904
rect 710 1908 716 1909
rect 710 1904 711 1908
rect 715 1904 716 1908
rect 710 1903 716 1904
rect 846 1908 852 1909
rect 846 1904 847 1908
rect 851 1904 852 1908
rect 846 1903 852 1904
rect 982 1908 988 1909
rect 982 1904 983 1908
rect 987 1904 988 1908
rect 982 1903 988 1904
rect 1118 1908 1124 1909
rect 1118 1904 1119 1908
rect 1123 1904 1124 1908
rect 1118 1903 1124 1904
rect 1254 1908 1260 1909
rect 1254 1904 1255 1908
rect 1259 1904 1260 1908
rect 1254 1903 1260 1904
rect 1382 1908 1388 1909
rect 1382 1904 1383 1908
rect 1387 1904 1388 1908
rect 1382 1903 1388 1904
rect 1518 1908 1524 1909
rect 1518 1904 1519 1908
rect 1523 1904 1524 1908
rect 1518 1903 1524 1904
rect 1654 1908 1660 1909
rect 1654 1904 1655 1908
rect 1659 1904 1660 1908
rect 1766 1907 1767 1911
rect 1771 1907 1772 1911
rect 1766 1906 1772 1907
rect 1654 1903 1660 1904
rect 1830 1892 1836 1893
rect 1806 1889 1812 1890
rect 1806 1885 1807 1889
rect 1811 1885 1812 1889
rect 1830 1888 1831 1892
rect 1835 1888 1836 1892
rect 1830 1887 1836 1888
rect 1918 1892 1924 1893
rect 1918 1888 1919 1892
rect 1923 1888 1924 1892
rect 1918 1887 1924 1888
rect 2038 1892 2044 1893
rect 2038 1888 2039 1892
rect 2043 1888 2044 1892
rect 2038 1887 2044 1888
rect 2166 1892 2172 1893
rect 2166 1888 2167 1892
rect 2171 1888 2172 1892
rect 2166 1887 2172 1888
rect 2302 1892 2308 1893
rect 2302 1888 2303 1892
rect 2307 1888 2308 1892
rect 2302 1887 2308 1888
rect 2454 1892 2460 1893
rect 2454 1888 2455 1892
rect 2459 1888 2460 1892
rect 2454 1887 2460 1888
rect 2614 1892 2620 1893
rect 2614 1888 2615 1892
rect 2619 1888 2620 1892
rect 2614 1887 2620 1888
rect 2790 1892 2796 1893
rect 2790 1888 2791 1892
rect 2795 1888 2796 1892
rect 2790 1887 2796 1888
rect 2982 1892 2988 1893
rect 2982 1888 2983 1892
rect 2987 1888 2988 1892
rect 2982 1887 2988 1888
rect 3182 1892 3188 1893
rect 3182 1888 3183 1892
rect 3187 1888 3188 1892
rect 3182 1887 3188 1888
rect 3366 1892 3372 1893
rect 3366 1888 3367 1892
rect 3371 1888 3372 1892
rect 3366 1887 3372 1888
rect 3462 1889 3468 1890
rect 1806 1884 1812 1885
rect 3462 1885 3463 1889
rect 3467 1885 3468 1889
rect 3462 1884 3468 1885
rect 1830 1873 1836 1874
rect 1806 1872 1812 1873
rect 1806 1868 1807 1872
rect 1811 1868 1812 1872
rect 1830 1869 1831 1873
rect 1835 1869 1836 1873
rect 1830 1868 1836 1869
rect 1918 1873 1924 1874
rect 1918 1869 1919 1873
rect 1923 1869 1924 1873
rect 1918 1868 1924 1869
rect 2038 1873 2044 1874
rect 2038 1869 2039 1873
rect 2043 1869 2044 1873
rect 2038 1868 2044 1869
rect 2166 1873 2172 1874
rect 2166 1869 2167 1873
rect 2171 1869 2172 1873
rect 2166 1868 2172 1869
rect 2302 1873 2308 1874
rect 2302 1869 2303 1873
rect 2307 1869 2308 1873
rect 2302 1868 2308 1869
rect 2454 1873 2460 1874
rect 2454 1869 2455 1873
rect 2459 1869 2460 1873
rect 2454 1868 2460 1869
rect 2614 1873 2620 1874
rect 2614 1869 2615 1873
rect 2619 1869 2620 1873
rect 2614 1868 2620 1869
rect 2790 1873 2796 1874
rect 2790 1869 2791 1873
rect 2795 1869 2796 1873
rect 2790 1868 2796 1869
rect 2982 1873 2988 1874
rect 2982 1869 2983 1873
rect 2987 1869 2988 1873
rect 2982 1868 2988 1869
rect 3182 1873 3188 1874
rect 3182 1869 3183 1873
rect 3187 1869 3188 1873
rect 3182 1868 3188 1869
rect 3366 1873 3372 1874
rect 3366 1869 3367 1873
rect 3371 1869 3372 1873
rect 3366 1868 3372 1869
rect 3462 1872 3468 1873
rect 3462 1868 3463 1872
rect 3467 1868 3468 1872
rect 1806 1867 1812 1868
rect 3462 1867 3468 1868
rect 558 1864 564 1865
rect 110 1861 116 1862
rect 110 1857 111 1861
rect 115 1857 116 1861
rect 558 1860 559 1864
rect 563 1860 564 1864
rect 558 1859 564 1860
rect 694 1864 700 1865
rect 694 1860 695 1864
rect 699 1860 700 1864
rect 694 1859 700 1860
rect 830 1864 836 1865
rect 830 1860 831 1864
rect 835 1860 836 1864
rect 830 1859 836 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1078 1864 1084 1865
rect 1078 1860 1079 1864
rect 1083 1860 1084 1864
rect 1078 1859 1084 1860
rect 1198 1864 1204 1865
rect 1198 1860 1199 1864
rect 1203 1860 1204 1864
rect 1198 1859 1204 1860
rect 1326 1864 1332 1865
rect 1326 1860 1327 1864
rect 1331 1860 1332 1864
rect 1326 1859 1332 1860
rect 1454 1864 1460 1865
rect 1454 1860 1455 1864
rect 1459 1860 1460 1864
rect 1454 1859 1460 1860
rect 1766 1861 1772 1862
rect 110 1856 116 1857
rect 1766 1857 1767 1861
rect 1771 1857 1772 1861
rect 1766 1856 1772 1857
rect 558 1845 564 1846
rect 110 1844 116 1845
rect 110 1840 111 1844
rect 115 1840 116 1844
rect 558 1841 559 1845
rect 563 1841 564 1845
rect 558 1840 564 1841
rect 694 1845 700 1846
rect 694 1841 695 1845
rect 699 1841 700 1845
rect 694 1840 700 1841
rect 830 1845 836 1846
rect 830 1841 831 1845
rect 835 1841 836 1845
rect 830 1840 836 1841
rect 958 1845 964 1846
rect 958 1841 959 1845
rect 963 1841 964 1845
rect 958 1840 964 1841
rect 1078 1845 1084 1846
rect 1078 1841 1079 1845
rect 1083 1841 1084 1845
rect 1078 1840 1084 1841
rect 1198 1845 1204 1846
rect 1198 1841 1199 1845
rect 1203 1841 1204 1845
rect 1198 1840 1204 1841
rect 1326 1845 1332 1846
rect 1326 1841 1327 1845
rect 1331 1841 1332 1845
rect 1326 1840 1332 1841
rect 1454 1845 1460 1846
rect 1454 1841 1455 1845
rect 1459 1841 1460 1845
rect 1454 1840 1460 1841
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 110 1839 116 1840
rect 1766 1839 1772 1840
rect 1806 1824 1812 1825
rect 3462 1824 3468 1825
rect 1806 1820 1807 1824
rect 1811 1820 1812 1824
rect 1806 1819 1812 1820
rect 1830 1823 1836 1824
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1958 1823 1964 1824
rect 1958 1819 1959 1823
rect 1963 1819 1964 1823
rect 1958 1818 1964 1819
rect 2110 1823 2116 1824
rect 2110 1819 2111 1823
rect 2115 1819 2116 1823
rect 2110 1818 2116 1819
rect 2254 1823 2260 1824
rect 2254 1819 2255 1823
rect 2259 1819 2260 1823
rect 2254 1818 2260 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 2566 1823 2572 1824
rect 2566 1819 2567 1823
rect 2571 1819 2572 1823
rect 2566 1818 2572 1819
rect 2742 1823 2748 1824
rect 2742 1819 2743 1823
rect 2747 1819 2748 1823
rect 2742 1818 2748 1819
rect 2934 1823 2940 1824
rect 2934 1819 2935 1823
rect 2939 1819 2940 1823
rect 2934 1818 2940 1819
rect 3134 1823 3140 1824
rect 3134 1819 3135 1823
rect 3139 1819 3140 1823
rect 3134 1818 3140 1819
rect 3342 1823 3348 1824
rect 3342 1819 3343 1823
rect 3347 1819 3348 1823
rect 3462 1820 3463 1824
rect 3467 1820 3468 1824
rect 3462 1819 3468 1820
rect 3342 1818 3348 1819
rect 1806 1807 1812 1808
rect 1806 1803 1807 1807
rect 1811 1803 1812 1807
rect 3462 1807 3468 1808
rect 1806 1802 1812 1803
rect 1830 1804 1836 1805
rect 1830 1800 1831 1804
rect 1835 1800 1836 1804
rect 1830 1799 1836 1800
rect 1958 1804 1964 1805
rect 1958 1800 1959 1804
rect 1963 1800 1964 1804
rect 1958 1799 1964 1800
rect 2110 1804 2116 1805
rect 2110 1800 2111 1804
rect 2115 1800 2116 1804
rect 2110 1799 2116 1800
rect 2254 1804 2260 1805
rect 2254 1800 2255 1804
rect 2259 1800 2260 1804
rect 2254 1799 2260 1800
rect 2406 1804 2412 1805
rect 2406 1800 2407 1804
rect 2411 1800 2412 1804
rect 2406 1799 2412 1800
rect 2566 1804 2572 1805
rect 2566 1800 2567 1804
rect 2571 1800 2572 1804
rect 2566 1799 2572 1800
rect 2742 1804 2748 1805
rect 2742 1800 2743 1804
rect 2747 1800 2748 1804
rect 2742 1799 2748 1800
rect 2934 1804 2940 1805
rect 2934 1800 2935 1804
rect 2939 1800 2940 1804
rect 2934 1799 2940 1800
rect 3134 1804 3140 1805
rect 3134 1800 3135 1804
rect 3139 1800 3140 1804
rect 3134 1799 3140 1800
rect 3342 1804 3348 1805
rect 3342 1800 3343 1804
rect 3347 1800 3348 1804
rect 3462 1803 3463 1807
rect 3467 1803 3468 1807
rect 3462 1802 3468 1803
rect 3342 1799 3348 1800
rect 110 1792 116 1793
rect 1766 1792 1772 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 222 1791 228 1792
rect 222 1787 223 1791
rect 227 1787 228 1791
rect 222 1786 228 1787
rect 310 1791 316 1792
rect 310 1787 311 1791
rect 315 1787 316 1791
rect 310 1786 316 1787
rect 406 1791 412 1792
rect 406 1787 407 1791
rect 411 1787 412 1791
rect 406 1786 412 1787
rect 526 1791 532 1792
rect 526 1787 527 1791
rect 531 1787 532 1791
rect 526 1786 532 1787
rect 654 1791 660 1792
rect 654 1787 655 1791
rect 659 1787 660 1791
rect 654 1786 660 1787
rect 798 1791 804 1792
rect 798 1787 799 1791
rect 803 1787 804 1791
rect 798 1786 804 1787
rect 942 1791 948 1792
rect 942 1787 943 1791
rect 947 1787 948 1791
rect 942 1786 948 1787
rect 1086 1791 1092 1792
rect 1086 1787 1087 1791
rect 1091 1787 1092 1791
rect 1086 1786 1092 1787
rect 1238 1791 1244 1792
rect 1238 1787 1239 1791
rect 1243 1787 1244 1791
rect 1238 1786 1244 1787
rect 1390 1791 1396 1792
rect 1390 1787 1391 1791
rect 1395 1787 1396 1791
rect 1390 1786 1396 1787
rect 1542 1791 1548 1792
rect 1542 1787 1543 1791
rect 1547 1787 1548 1791
rect 1542 1786 1548 1787
rect 1670 1791 1676 1792
rect 1670 1787 1671 1791
rect 1675 1787 1676 1791
rect 1766 1788 1767 1792
rect 1771 1788 1772 1792
rect 1766 1787 1772 1788
rect 1670 1786 1676 1787
rect 110 1775 116 1776
rect 110 1771 111 1775
rect 115 1771 116 1775
rect 1766 1775 1772 1776
rect 110 1770 116 1771
rect 134 1772 140 1773
rect 134 1768 135 1772
rect 139 1768 140 1772
rect 134 1767 140 1768
rect 222 1772 228 1773
rect 222 1768 223 1772
rect 227 1768 228 1772
rect 222 1767 228 1768
rect 310 1772 316 1773
rect 310 1768 311 1772
rect 315 1768 316 1772
rect 310 1767 316 1768
rect 406 1772 412 1773
rect 406 1768 407 1772
rect 411 1768 412 1772
rect 406 1767 412 1768
rect 526 1772 532 1773
rect 526 1768 527 1772
rect 531 1768 532 1772
rect 526 1767 532 1768
rect 654 1772 660 1773
rect 654 1768 655 1772
rect 659 1768 660 1772
rect 654 1767 660 1768
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 942 1772 948 1773
rect 942 1768 943 1772
rect 947 1768 948 1772
rect 942 1767 948 1768
rect 1086 1772 1092 1773
rect 1086 1768 1087 1772
rect 1091 1768 1092 1772
rect 1086 1767 1092 1768
rect 1238 1772 1244 1773
rect 1238 1768 1239 1772
rect 1243 1768 1244 1772
rect 1238 1767 1244 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1542 1772 1548 1773
rect 1542 1768 1543 1772
rect 1547 1768 1548 1772
rect 1542 1767 1548 1768
rect 1670 1772 1676 1773
rect 1670 1768 1671 1772
rect 1675 1768 1676 1772
rect 1766 1771 1767 1775
rect 1771 1771 1772 1775
rect 1766 1770 1772 1771
rect 1670 1767 1676 1768
rect 1878 1748 1884 1749
rect 1806 1745 1812 1746
rect 1806 1741 1807 1745
rect 1811 1741 1812 1745
rect 1878 1744 1879 1748
rect 1883 1744 1884 1748
rect 1878 1743 1884 1744
rect 2014 1748 2020 1749
rect 2014 1744 2015 1748
rect 2019 1744 2020 1748
rect 2014 1743 2020 1744
rect 2150 1748 2156 1749
rect 2150 1744 2151 1748
rect 2155 1744 2156 1748
rect 2150 1743 2156 1744
rect 2302 1748 2308 1749
rect 2302 1744 2303 1748
rect 2307 1744 2308 1748
rect 2302 1743 2308 1744
rect 2478 1748 2484 1749
rect 2478 1744 2479 1748
rect 2483 1744 2484 1748
rect 2478 1743 2484 1744
rect 2686 1748 2692 1749
rect 2686 1744 2687 1748
rect 2691 1744 2692 1748
rect 2686 1743 2692 1744
rect 2910 1748 2916 1749
rect 2910 1744 2911 1748
rect 2915 1744 2916 1748
rect 2910 1743 2916 1744
rect 3150 1748 3156 1749
rect 3150 1744 3151 1748
rect 3155 1744 3156 1748
rect 3150 1743 3156 1744
rect 3366 1748 3372 1749
rect 3366 1744 3367 1748
rect 3371 1744 3372 1748
rect 3366 1743 3372 1744
rect 3462 1745 3468 1746
rect 1806 1740 1812 1741
rect 3462 1741 3463 1745
rect 3467 1741 3468 1745
rect 3462 1740 3468 1741
rect 1878 1729 1884 1730
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1878 1725 1879 1729
rect 1883 1725 1884 1729
rect 1878 1724 1884 1725
rect 2014 1729 2020 1730
rect 2014 1725 2015 1729
rect 2019 1725 2020 1729
rect 2014 1724 2020 1725
rect 2150 1729 2156 1730
rect 2150 1725 2151 1729
rect 2155 1725 2156 1729
rect 2150 1724 2156 1725
rect 2302 1729 2308 1730
rect 2302 1725 2303 1729
rect 2307 1725 2308 1729
rect 2302 1724 2308 1725
rect 2478 1729 2484 1730
rect 2478 1725 2479 1729
rect 2483 1725 2484 1729
rect 2478 1724 2484 1725
rect 2686 1729 2692 1730
rect 2686 1725 2687 1729
rect 2691 1725 2692 1729
rect 2686 1724 2692 1725
rect 2910 1729 2916 1730
rect 2910 1725 2911 1729
rect 2915 1725 2916 1729
rect 2910 1724 2916 1725
rect 3150 1729 3156 1730
rect 3150 1725 3151 1729
rect 3155 1725 3156 1729
rect 3150 1724 3156 1725
rect 3366 1729 3372 1730
rect 3366 1725 3367 1729
rect 3371 1725 3372 1729
rect 3366 1724 3372 1725
rect 3462 1728 3468 1729
rect 3462 1724 3463 1728
rect 3467 1724 3468 1728
rect 1806 1723 1812 1724
rect 3462 1723 3468 1724
rect 134 1716 140 1717
rect 110 1713 116 1714
rect 110 1709 111 1713
rect 115 1709 116 1713
rect 134 1712 135 1716
rect 139 1712 140 1716
rect 134 1711 140 1712
rect 246 1716 252 1717
rect 246 1712 247 1716
rect 251 1712 252 1716
rect 246 1711 252 1712
rect 398 1716 404 1717
rect 398 1712 399 1716
rect 403 1712 404 1716
rect 398 1711 404 1712
rect 566 1716 572 1717
rect 566 1712 567 1716
rect 571 1712 572 1716
rect 566 1711 572 1712
rect 750 1716 756 1717
rect 750 1712 751 1716
rect 755 1712 756 1716
rect 750 1711 756 1712
rect 934 1716 940 1717
rect 934 1712 935 1716
rect 939 1712 940 1716
rect 934 1711 940 1712
rect 1118 1716 1124 1717
rect 1118 1712 1119 1716
rect 1123 1712 1124 1716
rect 1118 1711 1124 1712
rect 1310 1716 1316 1717
rect 1310 1712 1311 1716
rect 1315 1712 1316 1716
rect 1310 1711 1316 1712
rect 1502 1716 1508 1717
rect 1502 1712 1503 1716
rect 1507 1712 1508 1716
rect 1502 1711 1508 1712
rect 1670 1716 1676 1717
rect 1670 1712 1671 1716
rect 1675 1712 1676 1716
rect 1670 1711 1676 1712
rect 1766 1713 1772 1714
rect 110 1708 116 1709
rect 1766 1709 1767 1713
rect 1771 1709 1772 1713
rect 1766 1708 1772 1709
rect 134 1697 140 1698
rect 110 1696 116 1697
rect 110 1692 111 1696
rect 115 1692 116 1696
rect 134 1693 135 1697
rect 139 1693 140 1697
rect 134 1692 140 1693
rect 246 1697 252 1698
rect 246 1693 247 1697
rect 251 1693 252 1697
rect 246 1692 252 1693
rect 398 1697 404 1698
rect 398 1693 399 1697
rect 403 1693 404 1697
rect 398 1692 404 1693
rect 566 1697 572 1698
rect 566 1693 567 1697
rect 571 1693 572 1697
rect 566 1692 572 1693
rect 750 1697 756 1698
rect 750 1693 751 1697
rect 755 1693 756 1697
rect 750 1692 756 1693
rect 934 1697 940 1698
rect 934 1693 935 1697
rect 939 1693 940 1697
rect 934 1692 940 1693
rect 1118 1697 1124 1698
rect 1118 1693 1119 1697
rect 1123 1693 1124 1697
rect 1118 1692 1124 1693
rect 1310 1697 1316 1698
rect 1310 1693 1311 1697
rect 1315 1693 1316 1697
rect 1310 1692 1316 1693
rect 1502 1697 1508 1698
rect 1502 1693 1503 1697
rect 1507 1693 1508 1697
rect 1502 1692 1508 1693
rect 1670 1697 1676 1698
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 1766 1696 1772 1697
rect 1766 1692 1767 1696
rect 1771 1692 1772 1696
rect 110 1691 116 1692
rect 1766 1691 1772 1692
rect 1806 1676 1812 1677
rect 3462 1676 3468 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1830 1675 1836 1676
rect 1830 1671 1831 1675
rect 1835 1671 1836 1675
rect 1830 1670 1836 1671
rect 1934 1675 1940 1676
rect 1934 1671 1935 1675
rect 1939 1671 1940 1675
rect 1934 1670 1940 1671
rect 2062 1675 2068 1676
rect 2062 1671 2063 1675
rect 2067 1671 2068 1675
rect 2062 1670 2068 1671
rect 2182 1675 2188 1676
rect 2182 1671 2183 1675
rect 2187 1671 2188 1675
rect 2182 1670 2188 1671
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2310 1670 2316 1671
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1671 2444 1675
rect 2438 1670 2444 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1671 2580 1675
rect 2574 1670 2580 1671
rect 2726 1675 2732 1676
rect 2726 1671 2727 1675
rect 2731 1671 2732 1675
rect 2726 1670 2732 1671
rect 2886 1675 2892 1676
rect 2886 1671 2887 1675
rect 2891 1671 2892 1675
rect 2886 1670 2892 1671
rect 3046 1675 3052 1676
rect 3046 1671 3047 1675
rect 3051 1671 3052 1675
rect 3046 1670 3052 1671
rect 3214 1675 3220 1676
rect 3214 1671 3215 1675
rect 3219 1671 3220 1675
rect 3214 1670 3220 1671
rect 3366 1675 3372 1676
rect 3366 1671 3367 1675
rect 3371 1671 3372 1675
rect 3462 1672 3463 1676
rect 3467 1672 3468 1676
rect 3462 1671 3468 1672
rect 3366 1670 3372 1671
rect 1806 1659 1812 1660
rect 1806 1655 1807 1659
rect 1811 1655 1812 1659
rect 3462 1659 3468 1660
rect 1806 1654 1812 1655
rect 1830 1656 1836 1657
rect 1830 1652 1831 1656
rect 1835 1652 1836 1656
rect 1830 1651 1836 1652
rect 1934 1656 1940 1657
rect 1934 1652 1935 1656
rect 1939 1652 1940 1656
rect 1934 1651 1940 1652
rect 2062 1656 2068 1657
rect 2062 1652 2063 1656
rect 2067 1652 2068 1656
rect 2062 1651 2068 1652
rect 2182 1656 2188 1657
rect 2182 1652 2183 1656
rect 2187 1652 2188 1656
rect 2182 1651 2188 1652
rect 2310 1656 2316 1657
rect 2310 1652 2311 1656
rect 2315 1652 2316 1656
rect 2310 1651 2316 1652
rect 2438 1656 2444 1657
rect 2438 1652 2439 1656
rect 2443 1652 2444 1656
rect 2438 1651 2444 1652
rect 2574 1656 2580 1657
rect 2574 1652 2575 1656
rect 2579 1652 2580 1656
rect 2574 1651 2580 1652
rect 2726 1656 2732 1657
rect 2726 1652 2727 1656
rect 2731 1652 2732 1656
rect 2726 1651 2732 1652
rect 2886 1656 2892 1657
rect 2886 1652 2887 1656
rect 2891 1652 2892 1656
rect 2886 1651 2892 1652
rect 3046 1656 3052 1657
rect 3046 1652 3047 1656
rect 3051 1652 3052 1656
rect 3046 1651 3052 1652
rect 3214 1656 3220 1657
rect 3214 1652 3215 1656
rect 3219 1652 3220 1656
rect 3214 1651 3220 1652
rect 3366 1656 3372 1657
rect 3366 1652 3367 1656
rect 3371 1652 3372 1656
rect 3462 1655 3463 1659
rect 3467 1655 3468 1659
rect 3462 1654 3468 1655
rect 3366 1651 3372 1652
rect 110 1648 116 1649
rect 1766 1648 1772 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 190 1647 196 1648
rect 190 1643 191 1647
rect 195 1643 196 1647
rect 190 1642 196 1643
rect 294 1647 300 1648
rect 294 1643 295 1647
rect 299 1643 300 1647
rect 294 1642 300 1643
rect 406 1647 412 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 406 1642 412 1643
rect 534 1647 540 1648
rect 534 1643 535 1647
rect 539 1643 540 1647
rect 534 1642 540 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 854 1647 860 1648
rect 854 1643 855 1647
rect 859 1643 860 1647
rect 854 1642 860 1643
rect 1038 1647 1044 1648
rect 1038 1643 1039 1647
rect 1043 1643 1044 1647
rect 1038 1642 1044 1643
rect 1230 1647 1236 1648
rect 1230 1643 1231 1647
rect 1235 1643 1236 1647
rect 1230 1642 1236 1643
rect 1430 1647 1436 1648
rect 1430 1643 1431 1647
rect 1435 1643 1436 1647
rect 1430 1642 1436 1643
rect 1638 1647 1644 1648
rect 1638 1643 1639 1647
rect 1643 1643 1644 1647
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 1766 1643 1772 1644
rect 1638 1642 1644 1643
rect 110 1631 116 1632
rect 110 1627 111 1631
rect 115 1627 116 1631
rect 1766 1631 1772 1632
rect 110 1626 116 1627
rect 190 1628 196 1629
rect 190 1624 191 1628
rect 195 1624 196 1628
rect 190 1623 196 1624
rect 294 1628 300 1629
rect 294 1624 295 1628
rect 299 1624 300 1628
rect 294 1623 300 1624
rect 406 1628 412 1629
rect 406 1624 407 1628
rect 411 1624 412 1628
rect 406 1623 412 1624
rect 534 1628 540 1629
rect 534 1624 535 1628
rect 539 1624 540 1628
rect 534 1623 540 1624
rect 686 1628 692 1629
rect 686 1624 687 1628
rect 691 1624 692 1628
rect 686 1623 692 1624
rect 854 1628 860 1629
rect 854 1624 855 1628
rect 859 1624 860 1628
rect 854 1623 860 1624
rect 1038 1628 1044 1629
rect 1038 1624 1039 1628
rect 1043 1624 1044 1628
rect 1038 1623 1044 1624
rect 1230 1628 1236 1629
rect 1230 1624 1231 1628
rect 1235 1624 1236 1628
rect 1230 1623 1236 1624
rect 1430 1628 1436 1629
rect 1430 1624 1431 1628
rect 1435 1624 1436 1628
rect 1430 1623 1436 1624
rect 1638 1628 1644 1629
rect 1638 1624 1639 1628
rect 1643 1624 1644 1628
rect 1766 1627 1767 1631
rect 1771 1627 1772 1631
rect 1766 1626 1772 1627
rect 1638 1623 1644 1624
rect 1830 1604 1836 1605
rect 1806 1601 1812 1602
rect 1806 1597 1807 1601
rect 1811 1597 1812 1601
rect 1830 1600 1831 1604
rect 1835 1600 1836 1604
rect 1830 1599 1836 1600
rect 1942 1604 1948 1605
rect 1942 1600 1943 1604
rect 1947 1600 1948 1604
rect 1942 1599 1948 1600
rect 2086 1604 2092 1605
rect 2086 1600 2087 1604
rect 2091 1600 2092 1604
rect 2086 1599 2092 1600
rect 2230 1604 2236 1605
rect 2230 1600 2231 1604
rect 2235 1600 2236 1604
rect 2230 1599 2236 1600
rect 2366 1604 2372 1605
rect 2366 1600 2367 1604
rect 2371 1600 2372 1604
rect 2366 1599 2372 1600
rect 2502 1604 2508 1605
rect 2502 1600 2503 1604
rect 2507 1600 2508 1604
rect 2502 1599 2508 1600
rect 2638 1604 2644 1605
rect 2638 1600 2639 1604
rect 2643 1600 2644 1604
rect 2638 1599 2644 1600
rect 2766 1604 2772 1605
rect 2766 1600 2767 1604
rect 2771 1600 2772 1604
rect 2766 1599 2772 1600
rect 2894 1604 2900 1605
rect 2894 1600 2895 1604
rect 2899 1600 2900 1604
rect 2894 1599 2900 1600
rect 3014 1604 3020 1605
rect 3014 1600 3015 1604
rect 3019 1600 3020 1604
rect 3014 1599 3020 1600
rect 3134 1604 3140 1605
rect 3134 1600 3135 1604
rect 3139 1600 3140 1604
rect 3134 1599 3140 1600
rect 3262 1604 3268 1605
rect 3262 1600 3263 1604
rect 3267 1600 3268 1604
rect 3262 1599 3268 1600
rect 3366 1604 3372 1605
rect 3366 1600 3367 1604
rect 3371 1600 3372 1604
rect 3366 1599 3372 1600
rect 3462 1601 3468 1602
rect 1806 1596 1812 1597
rect 3462 1597 3463 1601
rect 3467 1597 3468 1601
rect 3462 1596 3468 1597
rect 1830 1585 1836 1586
rect 1806 1584 1812 1585
rect 326 1580 332 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 326 1576 327 1580
rect 331 1576 332 1580
rect 326 1575 332 1576
rect 430 1580 436 1581
rect 430 1576 431 1580
rect 435 1576 436 1580
rect 430 1575 436 1576
rect 542 1580 548 1581
rect 542 1576 543 1580
rect 547 1576 548 1580
rect 542 1575 548 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 966 1580 972 1581
rect 966 1576 967 1580
rect 971 1576 972 1580
rect 966 1575 972 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1278 1580 1284 1581
rect 1278 1576 1279 1580
rect 1283 1576 1284 1580
rect 1278 1575 1284 1576
rect 1438 1580 1444 1581
rect 1438 1576 1439 1580
rect 1443 1576 1444 1580
rect 1438 1575 1444 1576
rect 1606 1580 1612 1581
rect 1606 1576 1607 1580
rect 1611 1576 1612 1580
rect 1806 1580 1807 1584
rect 1811 1580 1812 1584
rect 1830 1581 1831 1585
rect 1835 1581 1836 1585
rect 1830 1580 1836 1581
rect 1942 1585 1948 1586
rect 1942 1581 1943 1585
rect 1947 1581 1948 1585
rect 1942 1580 1948 1581
rect 2086 1585 2092 1586
rect 2086 1581 2087 1585
rect 2091 1581 2092 1585
rect 2086 1580 2092 1581
rect 2230 1585 2236 1586
rect 2230 1581 2231 1585
rect 2235 1581 2236 1585
rect 2230 1580 2236 1581
rect 2366 1585 2372 1586
rect 2366 1581 2367 1585
rect 2371 1581 2372 1585
rect 2366 1580 2372 1581
rect 2502 1585 2508 1586
rect 2502 1581 2503 1585
rect 2507 1581 2508 1585
rect 2502 1580 2508 1581
rect 2638 1585 2644 1586
rect 2638 1581 2639 1585
rect 2643 1581 2644 1585
rect 2638 1580 2644 1581
rect 2766 1585 2772 1586
rect 2766 1581 2767 1585
rect 2771 1581 2772 1585
rect 2766 1580 2772 1581
rect 2894 1585 2900 1586
rect 2894 1581 2895 1585
rect 2899 1581 2900 1585
rect 2894 1580 2900 1581
rect 3014 1585 3020 1586
rect 3014 1581 3015 1585
rect 3019 1581 3020 1585
rect 3014 1580 3020 1581
rect 3134 1585 3140 1586
rect 3134 1581 3135 1585
rect 3139 1581 3140 1585
rect 3134 1580 3140 1581
rect 3262 1585 3268 1586
rect 3262 1581 3263 1585
rect 3267 1581 3268 1585
rect 3262 1580 3268 1581
rect 3366 1585 3372 1586
rect 3366 1581 3367 1585
rect 3371 1581 3372 1585
rect 3366 1580 3372 1581
rect 3462 1584 3468 1585
rect 3462 1580 3463 1584
rect 3467 1580 3468 1584
rect 1806 1579 1812 1580
rect 3462 1579 3468 1580
rect 1606 1575 1612 1576
rect 1766 1577 1772 1578
rect 110 1572 116 1573
rect 1766 1573 1767 1577
rect 1771 1573 1772 1577
rect 1766 1572 1772 1573
rect 326 1561 332 1562
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 326 1557 327 1561
rect 331 1557 332 1561
rect 326 1556 332 1557
rect 430 1561 436 1562
rect 430 1557 431 1561
rect 435 1557 436 1561
rect 430 1556 436 1557
rect 542 1561 548 1562
rect 542 1557 543 1561
rect 547 1557 548 1561
rect 542 1556 548 1557
rect 670 1561 676 1562
rect 670 1557 671 1561
rect 675 1557 676 1561
rect 670 1556 676 1557
rect 814 1561 820 1562
rect 814 1557 815 1561
rect 819 1557 820 1561
rect 814 1556 820 1557
rect 966 1561 972 1562
rect 966 1557 967 1561
rect 971 1557 972 1561
rect 966 1556 972 1557
rect 1118 1561 1124 1562
rect 1118 1557 1119 1561
rect 1123 1557 1124 1561
rect 1118 1556 1124 1557
rect 1278 1561 1284 1562
rect 1278 1557 1279 1561
rect 1283 1557 1284 1561
rect 1278 1556 1284 1557
rect 1438 1561 1444 1562
rect 1438 1557 1439 1561
rect 1443 1557 1444 1561
rect 1438 1556 1444 1557
rect 1606 1561 1612 1562
rect 1606 1557 1607 1561
rect 1611 1557 1612 1561
rect 1606 1556 1612 1557
rect 1766 1560 1772 1561
rect 1766 1556 1767 1560
rect 1771 1556 1772 1560
rect 110 1555 116 1556
rect 1766 1555 1772 1556
rect 1806 1532 1812 1533
rect 3462 1532 3468 1533
rect 1806 1528 1807 1532
rect 1811 1528 1812 1532
rect 1806 1527 1812 1528
rect 1838 1531 1844 1532
rect 1838 1527 1839 1531
rect 1843 1527 1844 1531
rect 1838 1526 1844 1527
rect 1990 1531 1996 1532
rect 1990 1527 1991 1531
rect 1995 1527 1996 1531
rect 1990 1526 1996 1527
rect 2150 1531 2156 1532
rect 2150 1527 2151 1531
rect 2155 1527 2156 1531
rect 2150 1526 2156 1527
rect 2302 1531 2308 1532
rect 2302 1527 2303 1531
rect 2307 1527 2308 1531
rect 2302 1526 2308 1527
rect 2454 1531 2460 1532
rect 2454 1527 2455 1531
rect 2459 1527 2460 1531
rect 2454 1526 2460 1527
rect 2598 1531 2604 1532
rect 2598 1527 2599 1531
rect 2603 1527 2604 1531
rect 2598 1526 2604 1527
rect 2734 1531 2740 1532
rect 2734 1527 2735 1531
rect 2739 1527 2740 1531
rect 2734 1526 2740 1527
rect 2870 1531 2876 1532
rect 2870 1527 2871 1531
rect 2875 1527 2876 1531
rect 2870 1526 2876 1527
rect 3006 1531 3012 1532
rect 3006 1527 3007 1531
rect 3011 1527 3012 1531
rect 3006 1526 3012 1527
rect 3142 1531 3148 1532
rect 3142 1527 3143 1531
rect 3147 1527 3148 1531
rect 3462 1528 3463 1532
rect 3467 1528 3468 1532
rect 3462 1527 3468 1528
rect 3142 1526 3148 1527
rect 1806 1515 1812 1516
rect 110 1512 116 1513
rect 1766 1512 1772 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 222 1511 228 1512
rect 222 1507 223 1511
rect 227 1507 228 1511
rect 222 1506 228 1507
rect 342 1511 348 1512
rect 342 1507 343 1511
rect 347 1507 348 1511
rect 342 1506 348 1507
rect 470 1511 476 1512
rect 470 1507 471 1511
rect 475 1507 476 1511
rect 470 1506 476 1507
rect 606 1511 612 1512
rect 606 1507 607 1511
rect 611 1507 612 1511
rect 606 1506 612 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 894 1511 900 1512
rect 894 1507 895 1511
rect 899 1507 900 1511
rect 894 1506 900 1507
rect 1046 1511 1052 1512
rect 1046 1507 1047 1511
rect 1051 1507 1052 1511
rect 1046 1506 1052 1507
rect 1198 1511 1204 1512
rect 1198 1507 1199 1511
rect 1203 1507 1204 1511
rect 1198 1506 1204 1507
rect 1350 1511 1356 1512
rect 1350 1507 1351 1511
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1502 1511 1508 1512
rect 1502 1507 1503 1511
rect 1507 1507 1508 1511
rect 1766 1508 1767 1512
rect 1771 1508 1772 1512
rect 1806 1511 1807 1515
rect 1811 1511 1812 1515
rect 3462 1515 3468 1516
rect 1806 1510 1812 1511
rect 1838 1512 1844 1513
rect 1766 1507 1772 1508
rect 1838 1508 1839 1512
rect 1843 1508 1844 1512
rect 1838 1507 1844 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2150 1512 2156 1513
rect 2150 1508 2151 1512
rect 2155 1508 2156 1512
rect 2150 1507 2156 1508
rect 2302 1512 2308 1513
rect 2302 1508 2303 1512
rect 2307 1508 2308 1512
rect 2302 1507 2308 1508
rect 2454 1512 2460 1513
rect 2454 1508 2455 1512
rect 2459 1508 2460 1512
rect 2454 1507 2460 1508
rect 2598 1512 2604 1513
rect 2598 1508 2599 1512
rect 2603 1508 2604 1512
rect 2598 1507 2604 1508
rect 2734 1512 2740 1513
rect 2734 1508 2735 1512
rect 2739 1508 2740 1512
rect 2734 1507 2740 1508
rect 2870 1512 2876 1513
rect 2870 1508 2871 1512
rect 2875 1508 2876 1512
rect 2870 1507 2876 1508
rect 3006 1512 3012 1513
rect 3006 1508 3007 1512
rect 3011 1508 3012 1512
rect 3006 1507 3012 1508
rect 3142 1512 3148 1513
rect 3142 1508 3143 1512
rect 3147 1508 3148 1512
rect 3462 1511 3463 1515
rect 3467 1511 3468 1515
rect 3462 1510 3468 1511
rect 3142 1507 3148 1508
rect 1502 1506 1508 1507
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 1766 1495 1772 1496
rect 110 1490 116 1491
rect 222 1492 228 1493
rect 222 1488 223 1492
rect 227 1488 228 1492
rect 222 1487 228 1488
rect 342 1492 348 1493
rect 342 1488 343 1492
rect 347 1488 348 1492
rect 342 1487 348 1488
rect 470 1492 476 1493
rect 470 1488 471 1492
rect 475 1488 476 1492
rect 470 1487 476 1488
rect 606 1492 612 1493
rect 606 1488 607 1492
rect 611 1488 612 1492
rect 606 1487 612 1488
rect 750 1492 756 1493
rect 750 1488 751 1492
rect 755 1488 756 1492
rect 750 1487 756 1488
rect 894 1492 900 1493
rect 894 1488 895 1492
rect 899 1488 900 1492
rect 894 1487 900 1488
rect 1046 1492 1052 1493
rect 1046 1488 1047 1492
rect 1051 1488 1052 1492
rect 1046 1487 1052 1488
rect 1198 1492 1204 1493
rect 1198 1488 1199 1492
rect 1203 1488 1204 1492
rect 1198 1487 1204 1488
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1502 1492 1508 1493
rect 1502 1488 1503 1492
rect 1507 1488 1508 1492
rect 1766 1491 1767 1495
rect 1771 1491 1772 1495
rect 1766 1490 1772 1491
rect 1502 1487 1508 1488
rect 1942 1460 1948 1461
rect 1806 1457 1812 1458
rect 1806 1453 1807 1457
rect 1811 1453 1812 1457
rect 1942 1456 1943 1460
rect 1947 1456 1948 1460
rect 1942 1455 1948 1456
rect 2054 1460 2060 1461
rect 2054 1456 2055 1460
rect 2059 1456 2060 1460
rect 2054 1455 2060 1456
rect 2190 1460 2196 1461
rect 2190 1456 2191 1460
rect 2195 1456 2196 1460
rect 2190 1455 2196 1456
rect 2334 1460 2340 1461
rect 2334 1456 2335 1460
rect 2339 1456 2340 1460
rect 2334 1455 2340 1456
rect 2478 1460 2484 1461
rect 2478 1456 2479 1460
rect 2483 1456 2484 1460
rect 2478 1455 2484 1456
rect 2630 1460 2636 1461
rect 2630 1456 2631 1460
rect 2635 1456 2636 1460
rect 2630 1455 2636 1456
rect 2782 1460 2788 1461
rect 2782 1456 2783 1460
rect 2787 1456 2788 1460
rect 2782 1455 2788 1456
rect 2934 1460 2940 1461
rect 2934 1456 2935 1460
rect 2939 1456 2940 1460
rect 2934 1455 2940 1456
rect 3086 1460 3092 1461
rect 3086 1456 3087 1460
rect 3091 1456 3092 1460
rect 3086 1455 3092 1456
rect 3238 1460 3244 1461
rect 3238 1456 3239 1460
rect 3243 1456 3244 1460
rect 3238 1455 3244 1456
rect 3462 1457 3468 1458
rect 1806 1452 1812 1453
rect 3462 1453 3463 1457
rect 3467 1453 3468 1457
rect 3462 1452 3468 1453
rect 1942 1441 1948 1442
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 302 1440 308 1441
rect 302 1436 303 1440
rect 307 1436 308 1440
rect 302 1435 308 1436
rect 470 1440 476 1441
rect 470 1436 471 1440
rect 475 1436 476 1440
rect 470 1435 476 1436
rect 630 1440 636 1441
rect 630 1436 631 1440
rect 635 1436 636 1440
rect 630 1435 636 1436
rect 782 1440 788 1441
rect 782 1436 783 1440
rect 787 1436 788 1440
rect 782 1435 788 1436
rect 926 1440 932 1441
rect 926 1436 927 1440
rect 931 1436 932 1440
rect 926 1435 932 1436
rect 1062 1440 1068 1441
rect 1062 1436 1063 1440
rect 1067 1436 1068 1440
rect 1062 1435 1068 1436
rect 1198 1440 1204 1441
rect 1198 1436 1199 1440
rect 1203 1436 1204 1440
rect 1198 1435 1204 1436
rect 1334 1440 1340 1441
rect 1334 1436 1335 1440
rect 1339 1436 1340 1440
rect 1334 1435 1340 1436
rect 1470 1440 1476 1441
rect 1470 1436 1471 1440
rect 1475 1436 1476 1440
rect 1806 1440 1812 1441
rect 1470 1435 1476 1436
rect 1766 1437 1772 1438
rect 110 1432 116 1433
rect 1766 1433 1767 1437
rect 1771 1433 1772 1437
rect 1806 1436 1807 1440
rect 1811 1436 1812 1440
rect 1942 1437 1943 1441
rect 1947 1437 1948 1441
rect 1942 1436 1948 1437
rect 2054 1441 2060 1442
rect 2054 1437 2055 1441
rect 2059 1437 2060 1441
rect 2054 1436 2060 1437
rect 2190 1441 2196 1442
rect 2190 1437 2191 1441
rect 2195 1437 2196 1441
rect 2190 1436 2196 1437
rect 2334 1441 2340 1442
rect 2334 1437 2335 1441
rect 2339 1437 2340 1441
rect 2334 1436 2340 1437
rect 2478 1441 2484 1442
rect 2478 1437 2479 1441
rect 2483 1437 2484 1441
rect 2478 1436 2484 1437
rect 2630 1441 2636 1442
rect 2630 1437 2631 1441
rect 2635 1437 2636 1441
rect 2630 1436 2636 1437
rect 2782 1441 2788 1442
rect 2782 1437 2783 1441
rect 2787 1437 2788 1441
rect 2782 1436 2788 1437
rect 2934 1441 2940 1442
rect 2934 1437 2935 1441
rect 2939 1437 2940 1441
rect 2934 1436 2940 1437
rect 3086 1441 3092 1442
rect 3086 1437 3087 1441
rect 3091 1437 3092 1441
rect 3086 1436 3092 1437
rect 3238 1441 3244 1442
rect 3238 1437 3239 1441
rect 3243 1437 3244 1441
rect 3238 1436 3244 1437
rect 3462 1440 3468 1441
rect 3462 1436 3463 1440
rect 3467 1436 3468 1440
rect 1806 1435 1812 1436
rect 3462 1435 3468 1436
rect 1766 1432 1772 1433
rect 134 1421 140 1422
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 134 1417 135 1421
rect 139 1417 140 1421
rect 134 1416 140 1417
rect 302 1421 308 1422
rect 302 1417 303 1421
rect 307 1417 308 1421
rect 302 1416 308 1417
rect 470 1421 476 1422
rect 470 1417 471 1421
rect 475 1417 476 1421
rect 470 1416 476 1417
rect 630 1421 636 1422
rect 630 1417 631 1421
rect 635 1417 636 1421
rect 630 1416 636 1417
rect 782 1421 788 1422
rect 782 1417 783 1421
rect 787 1417 788 1421
rect 782 1416 788 1417
rect 926 1421 932 1422
rect 926 1417 927 1421
rect 931 1417 932 1421
rect 926 1416 932 1417
rect 1062 1421 1068 1422
rect 1062 1417 1063 1421
rect 1067 1417 1068 1421
rect 1062 1416 1068 1417
rect 1198 1421 1204 1422
rect 1198 1417 1199 1421
rect 1203 1417 1204 1421
rect 1198 1416 1204 1417
rect 1334 1421 1340 1422
rect 1334 1417 1335 1421
rect 1339 1417 1340 1421
rect 1334 1416 1340 1417
rect 1470 1421 1476 1422
rect 1470 1417 1471 1421
rect 1475 1417 1476 1421
rect 1470 1416 1476 1417
rect 1766 1420 1772 1421
rect 1766 1416 1767 1420
rect 1771 1416 1772 1420
rect 110 1415 116 1416
rect 1766 1415 1772 1416
rect 1806 1388 1812 1389
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 2094 1387 2100 1388
rect 2094 1383 2095 1387
rect 2099 1383 2100 1387
rect 2094 1382 2100 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2318 1387 2324 1388
rect 2318 1383 2319 1387
rect 2323 1383 2324 1387
rect 2318 1382 2324 1383
rect 2454 1387 2460 1388
rect 2454 1383 2455 1387
rect 2459 1383 2460 1387
rect 2454 1382 2460 1383
rect 2598 1387 2604 1388
rect 2598 1383 2599 1387
rect 2603 1383 2604 1387
rect 2598 1382 2604 1383
rect 2742 1387 2748 1388
rect 2742 1383 2743 1387
rect 2747 1383 2748 1387
rect 2742 1382 2748 1383
rect 2886 1387 2892 1388
rect 2886 1383 2887 1387
rect 2891 1383 2892 1387
rect 2886 1382 2892 1383
rect 3030 1387 3036 1388
rect 3030 1383 3031 1387
rect 3035 1383 3036 1387
rect 3030 1382 3036 1383
rect 3174 1387 3180 1388
rect 3174 1383 3175 1387
rect 3179 1383 3180 1387
rect 3174 1382 3180 1383
rect 3326 1387 3332 1388
rect 3326 1383 3327 1387
rect 3331 1383 3332 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3326 1382 3332 1383
rect 110 1372 116 1373
rect 1766 1372 1772 1373
rect 110 1368 111 1372
rect 115 1368 116 1372
rect 110 1367 116 1368
rect 134 1371 140 1372
rect 134 1367 135 1371
rect 139 1367 140 1371
rect 134 1366 140 1367
rect 278 1371 284 1372
rect 278 1367 279 1371
rect 283 1367 284 1371
rect 278 1366 284 1367
rect 446 1371 452 1372
rect 446 1367 447 1371
rect 451 1367 452 1371
rect 446 1366 452 1367
rect 606 1371 612 1372
rect 606 1367 607 1371
rect 611 1367 612 1371
rect 606 1366 612 1367
rect 758 1371 764 1372
rect 758 1367 759 1371
rect 763 1367 764 1371
rect 758 1366 764 1367
rect 902 1371 908 1372
rect 902 1367 903 1371
rect 907 1367 908 1371
rect 902 1366 908 1367
rect 1030 1371 1036 1372
rect 1030 1367 1031 1371
rect 1035 1367 1036 1371
rect 1030 1366 1036 1367
rect 1158 1371 1164 1372
rect 1158 1367 1159 1371
rect 1163 1367 1164 1371
rect 1158 1366 1164 1367
rect 1286 1371 1292 1372
rect 1286 1367 1287 1371
rect 1291 1367 1292 1371
rect 1286 1366 1292 1367
rect 1414 1371 1420 1372
rect 1414 1367 1415 1371
rect 1419 1367 1420 1371
rect 1766 1368 1767 1372
rect 1771 1368 1772 1372
rect 1766 1367 1772 1368
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 3462 1371 3468 1372
rect 1414 1366 1420 1367
rect 1806 1366 1812 1367
rect 2094 1368 2100 1369
rect 2094 1364 2095 1368
rect 2099 1364 2100 1368
rect 2094 1363 2100 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2318 1368 2324 1369
rect 2318 1364 2319 1368
rect 2323 1364 2324 1368
rect 2318 1363 2324 1364
rect 2454 1368 2460 1369
rect 2454 1364 2455 1368
rect 2459 1364 2460 1368
rect 2454 1363 2460 1364
rect 2598 1368 2604 1369
rect 2598 1364 2599 1368
rect 2603 1364 2604 1368
rect 2598 1363 2604 1364
rect 2742 1368 2748 1369
rect 2742 1364 2743 1368
rect 2747 1364 2748 1368
rect 2742 1363 2748 1364
rect 2886 1368 2892 1369
rect 2886 1364 2887 1368
rect 2891 1364 2892 1368
rect 2886 1363 2892 1364
rect 3030 1368 3036 1369
rect 3030 1364 3031 1368
rect 3035 1364 3036 1368
rect 3030 1363 3036 1364
rect 3174 1368 3180 1369
rect 3174 1364 3175 1368
rect 3179 1364 3180 1368
rect 3174 1363 3180 1364
rect 3326 1368 3332 1369
rect 3326 1364 3327 1368
rect 3331 1364 3332 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3326 1363 3332 1364
rect 110 1355 116 1356
rect 110 1351 111 1355
rect 115 1351 116 1355
rect 1766 1355 1772 1356
rect 110 1350 116 1351
rect 134 1352 140 1353
rect 134 1348 135 1352
rect 139 1348 140 1352
rect 134 1347 140 1348
rect 278 1352 284 1353
rect 278 1348 279 1352
rect 283 1348 284 1352
rect 278 1347 284 1348
rect 446 1352 452 1353
rect 446 1348 447 1352
rect 451 1348 452 1352
rect 446 1347 452 1348
rect 606 1352 612 1353
rect 606 1348 607 1352
rect 611 1348 612 1352
rect 606 1347 612 1348
rect 758 1352 764 1353
rect 758 1348 759 1352
rect 763 1348 764 1352
rect 758 1347 764 1348
rect 902 1352 908 1353
rect 902 1348 903 1352
rect 907 1348 908 1352
rect 902 1347 908 1348
rect 1030 1352 1036 1353
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 1158 1352 1164 1353
rect 1158 1348 1159 1352
rect 1163 1348 1164 1352
rect 1158 1347 1164 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1414 1352 1420 1353
rect 1414 1348 1415 1352
rect 1419 1348 1420 1352
rect 1766 1351 1767 1355
rect 1771 1351 1772 1355
rect 1766 1350 1772 1351
rect 1414 1347 1420 1348
rect 2102 1320 2108 1321
rect 1806 1317 1812 1318
rect 1806 1313 1807 1317
rect 1811 1313 1812 1317
rect 2102 1316 2103 1320
rect 2107 1316 2108 1320
rect 2102 1315 2108 1316
rect 2238 1320 2244 1321
rect 2238 1316 2239 1320
rect 2243 1316 2244 1320
rect 2238 1315 2244 1316
rect 2382 1320 2388 1321
rect 2382 1316 2383 1320
rect 2387 1316 2388 1320
rect 2382 1315 2388 1316
rect 2534 1320 2540 1321
rect 2534 1316 2535 1320
rect 2539 1316 2540 1320
rect 2534 1315 2540 1316
rect 2686 1320 2692 1321
rect 2686 1316 2687 1320
rect 2691 1316 2692 1320
rect 2686 1315 2692 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2990 1320 2996 1321
rect 2990 1316 2991 1320
rect 2995 1316 2996 1320
rect 2990 1315 2996 1316
rect 3142 1320 3148 1321
rect 3142 1316 3143 1320
rect 3147 1316 3148 1320
rect 3142 1315 3148 1316
rect 3302 1320 3308 1321
rect 3302 1316 3303 1320
rect 3307 1316 3308 1320
rect 3302 1315 3308 1316
rect 3462 1317 3468 1318
rect 1806 1312 1812 1313
rect 3462 1313 3463 1317
rect 3467 1313 3468 1317
rect 3462 1312 3468 1313
rect 134 1304 140 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 134 1300 135 1304
rect 139 1300 140 1304
rect 134 1299 140 1300
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 438 1304 444 1305
rect 438 1300 439 1304
rect 443 1300 444 1304
rect 438 1299 444 1300
rect 582 1304 588 1305
rect 582 1300 583 1304
rect 587 1300 588 1304
rect 582 1299 588 1300
rect 718 1304 724 1305
rect 718 1300 719 1304
rect 723 1300 724 1304
rect 718 1299 724 1300
rect 846 1304 852 1305
rect 846 1300 847 1304
rect 851 1300 852 1304
rect 846 1299 852 1300
rect 966 1304 972 1305
rect 966 1300 967 1304
rect 971 1300 972 1304
rect 966 1299 972 1300
rect 1078 1304 1084 1305
rect 1078 1300 1079 1304
rect 1083 1300 1084 1304
rect 1078 1299 1084 1300
rect 1190 1304 1196 1305
rect 1190 1300 1191 1304
rect 1195 1300 1196 1304
rect 1190 1299 1196 1300
rect 1310 1304 1316 1305
rect 1310 1300 1311 1304
rect 1315 1300 1316 1304
rect 1310 1299 1316 1300
rect 1766 1301 1772 1302
rect 2102 1301 2108 1302
rect 110 1296 116 1297
rect 1766 1297 1767 1301
rect 1771 1297 1772 1301
rect 1766 1296 1772 1297
rect 1806 1300 1812 1301
rect 1806 1296 1807 1300
rect 1811 1296 1812 1300
rect 2102 1297 2103 1301
rect 2107 1297 2108 1301
rect 2102 1296 2108 1297
rect 2238 1301 2244 1302
rect 2238 1297 2239 1301
rect 2243 1297 2244 1301
rect 2238 1296 2244 1297
rect 2382 1301 2388 1302
rect 2382 1297 2383 1301
rect 2387 1297 2388 1301
rect 2382 1296 2388 1297
rect 2534 1301 2540 1302
rect 2534 1297 2535 1301
rect 2539 1297 2540 1301
rect 2534 1296 2540 1297
rect 2686 1301 2692 1302
rect 2686 1297 2687 1301
rect 2691 1297 2692 1301
rect 2686 1296 2692 1297
rect 2838 1301 2844 1302
rect 2838 1297 2839 1301
rect 2843 1297 2844 1301
rect 2838 1296 2844 1297
rect 2990 1301 2996 1302
rect 2990 1297 2991 1301
rect 2995 1297 2996 1301
rect 2990 1296 2996 1297
rect 3142 1301 3148 1302
rect 3142 1297 3143 1301
rect 3147 1297 3148 1301
rect 3142 1296 3148 1297
rect 3302 1301 3308 1302
rect 3302 1297 3303 1301
rect 3307 1297 3308 1301
rect 3302 1296 3308 1297
rect 3462 1300 3468 1301
rect 3462 1296 3463 1300
rect 3467 1296 3468 1300
rect 1806 1295 1812 1296
rect 3462 1295 3468 1296
rect 134 1285 140 1286
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 134 1281 135 1285
rect 139 1281 140 1285
rect 134 1280 140 1281
rect 278 1285 284 1286
rect 278 1281 279 1285
rect 283 1281 284 1285
rect 278 1280 284 1281
rect 438 1285 444 1286
rect 438 1281 439 1285
rect 443 1281 444 1285
rect 438 1280 444 1281
rect 582 1285 588 1286
rect 582 1281 583 1285
rect 587 1281 588 1285
rect 582 1280 588 1281
rect 718 1285 724 1286
rect 718 1281 719 1285
rect 723 1281 724 1285
rect 718 1280 724 1281
rect 846 1285 852 1286
rect 846 1281 847 1285
rect 851 1281 852 1285
rect 846 1280 852 1281
rect 966 1285 972 1286
rect 966 1281 967 1285
rect 971 1281 972 1285
rect 966 1280 972 1281
rect 1078 1285 1084 1286
rect 1078 1281 1079 1285
rect 1083 1281 1084 1285
rect 1078 1280 1084 1281
rect 1190 1285 1196 1286
rect 1190 1281 1191 1285
rect 1195 1281 1196 1285
rect 1190 1280 1196 1281
rect 1310 1285 1316 1286
rect 1310 1281 1311 1285
rect 1315 1281 1316 1285
rect 1310 1280 1316 1281
rect 1766 1284 1772 1285
rect 1766 1280 1767 1284
rect 1771 1280 1772 1284
rect 110 1279 116 1280
rect 1766 1279 1772 1280
rect 1806 1256 1812 1257
rect 3462 1256 3468 1257
rect 1806 1252 1807 1256
rect 1811 1252 1812 1256
rect 1806 1251 1812 1252
rect 1934 1255 1940 1256
rect 1934 1251 1935 1255
rect 1939 1251 1940 1255
rect 1934 1250 1940 1251
rect 2062 1255 2068 1256
rect 2062 1251 2063 1255
rect 2067 1251 2068 1255
rect 2062 1250 2068 1251
rect 2198 1255 2204 1256
rect 2198 1251 2199 1255
rect 2203 1251 2204 1255
rect 2198 1250 2204 1251
rect 2342 1255 2348 1256
rect 2342 1251 2343 1255
rect 2347 1251 2348 1255
rect 2342 1250 2348 1251
rect 2494 1255 2500 1256
rect 2494 1251 2495 1255
rect 2499 1251 2500 1255
rect 2494 1250 2500 1251
rect 2654 1255 2660 1256
rect 2654 1251 2655 1255
rect 2659 1251 2660 1255
rect 2654 1250 2660 1251
rect 2814 1255 2820 1256
rect 2814 1251 2815 1255
rect 2819 1251 2820 1255
rect 2814 1250 2820 1251
rect 2974 1255 2980 1256
rect 2974 1251 2975 1255
rect 2979 1251 2980 1255
rect 2974 1250 2980 1251
rect 3142 1255 3148 1256
rect 3142 1251 3143 1255
rect 3147 1251 3148 1255
rect 3462 1252 3463 1256
rect 3467 1252 3468 1256
rect 3462 1251 3468 1252
rect 3142 1250 3148 1251
rect 1806 1239 1812 1240
rect 110 1236 116 1237
rect 1766 1236 1772 1237
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 110 1231 116 1232
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 238 1235 244 1236
rect 238 1231 239 1235
rect 243 1231 244 1235
rect 238 1230 244 1231
rect 366 1235 372 1236
rect 366 1231 367 1235
rect 371 1231 372 1235
rect 366 1230 372 1231
rect 494 1235 500 1236
rect 494 1231 495 1235
rect 499 1231 500 1235
rect 494 1230 500 1231
rect 614 1235 620 1236
rect 614 1231 615 1235
rect 619 1231 620 1235
rect 614 1230 620 1231
rect 734 1235 740 1236
rect 734 1231 735 1235
rect 739 1231 740 1235
rect 734 1230 740 1231
rect 846 1235 852 1236
rect 846 1231 847 1235
rect 851 1231 852 1235
rect 846 1230 852 1231
rect 958 1235 964 1236
rect 958 1231 959 1235
rect 963 1231 964 1235
rect 958 1230 964 1231
rect 1070 1235 1076 1236
rect 1070 1231 1071 1235
rect 1075 1231 1076 1235
rect 1070 1230 1076 1231
rect 1190 1235 1196 1236
rect 1190 1231 1191 1235
rect 1195 1231 1196 1235
rect 1766 1232 1767 1236
rect 1771 1232 1772 1236
rect 1806 1235 1807 1239
rect 1811 1235 1812 1239
rect 3462 1239 3468 1240
rect 1806 1234 1812 1235
rect 1934 1236 1940 1237
rect 1766 1231 1772 1232
rect 1934 1232 1935 1236
rect 1939 1232 1940 1236
rect 1934 1231 1940 1232
rect 2062 1236 2068 1237
rect 2062 1232 2063 1236
rect 2067 1232 2068 1236
rect 2062 1231 2068 1232
rect 2198 1236 2204 1237
rect 2198 1232 2199 1236
rect 2203 1232 2204 1236
rect 2198 1231 2204 1232
rect 2342 1236 2348 1237
rect 2342 1232 2343 1236
rect 2347 1232 2348 1236
rect 2342 1231 2348 1232
rect 2494 1236 2500 1237
rect 2494 1232 2495 1236
rect 2499 1232 2500 1236
rect 2494 1231 2500 1232
rect 2654 1236 2660 1237
rect 2654 1232 2655 1236
rect 2659 1232 2660 1236
rect 2654 1231 2660 1232
rect 2814 1236 2820 1237
rect 2814 1232 2815 1236
rect 2819 1232 2820 1236
rect 2814 1231 2820 1232
rect 2974 1236 2980 1237
rect 2974 1232 2975 1236
rect 2979 1232 2980 1236
rect 2974 1231 2980 1232
rect 3142 1236 3148 1237
rect 3142 1232 3143 1236
rect 3147 1232 3148 1236
rect 3462 1235 3463 1239
rect 3467 1235 3468 1239
rect 3462 1234 3468 1235
rect 3142 1231 3148 1232
rect 1190 1230 1196 1231
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 1766 1219 1772 1220
rect 110 1214 116 1215
rect 134 1216 140 1217
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 238 1216 244 1217
rect 238 1212 239 1216
rect 243 1212 244 1216
rect 238 1211 244 1212
rect 366 1216 372 1217
rect 366 1212 367 1216
rect 371 1212 372 1216
rect 366 1211 372 1212
rect 494 1216 500 1217
rect 494 1212 495 1216
rect 499 1212 500 1216
rect 494 1211 500 1212
rect 614 1216 620 1217
rect 614 1212 615 1216
rect 619 1212 620 1216
rect 614 1211 620 1212
rect 734 1216 740 1217
rect 734 1212 735 1216
rect 739 1212 740 1216
rect 734 1211 740 1212
rect 846 1216 852 1217
rect 846 1212 847 1216
rect 851 1212 852 1216
rect 846 1211 852 1212
rect 958 1216 964 1217
rect 958 1212 959 1216
rect 963 1212 964 1216
rect 958 1211 964 1212
rect 1070 1216 1076 1217
rect 1070 1212 1071 1216
rect 1075 1212 1076 1216
rect 1070 1211 1076 1212
rect 1190 1216 1196 1217
rect 1190 1212 1191 1216
rect 1195 1212 1196 1216
rect 1766 1215 1767 1219
rect 1771 1215 1772 1219
rect 1766 1214 1772 1215
rect 1190 1211 1196 1212
rect 1830 1192 1836 1193
rect 1806 1189 1812 1190
rect 1806 1185 1807 1189
rect 1811 1185 1812 1189
rect 1830 1188 1831 1192
rect 1835 1188 1836 1192
rect 1830 1187 1836 1188
rect 1934 1192 1940 1193
rect 1934 1188 1935 1192
rect 1939 1188 1940 1192
rect 1934 1187 1940 1188
rect 2078 1192 2084 1193
rect 2078 1188 2079 1192
rect 2083 1188 2084 1192
rect 2078 1187 2084 1188
rect 2230 1192 2236 1193
rect 2230 1188 2231 1192
rect 2235 1188 2236 1192
rect 2230 1187 2236 1188
rect 2390 1192 2396 1193
rect 2390 1188 2391 1192
rect 2395 1188 2396 1192
rect 2390 1187 2396 1188
rect 2542 1192 2548 1193
rect 2542 1188 2543 1192
rect 2547 1188 2548 1192
rect 2542 1187 2548 1188
rect 2694 1192 2700 1193
rect 2694 1188 2695 1192
rect 2699 1188 2700 1192
rect 2694 1187 2700 1188
rect 2846 1192 2852 1193
rect 2846 1188 2847 1192
rect 2851 1188 2852 1192
rect 2846 1187 2852 1188
rect 2998 1192 3004 1193
rect 2998 1188 2999 1192
rect 3003 1188 3004 1192
rect 2998 1187 3004 1188
rect 3158 1192 3164 1193
rect 3158 1188 3159 1192
rect 3163 1188 3164 1192
rect 3158 1187 3164 1188
rect 3462 1189 3468 1190
rect 1806 1184 1812 1185
rect 3462 1185 3463 1189
rect 3467 1185 3468 1189
rect 3462 1184 3468 1185
rect 1830 1173 1836 1174
rect 1806 1172 1812 1173
rect 134 1168 140 1169
rect 110 1165 116 1166
rect 110 1161 111 1165
rect 115 1161 116 1165
rect 134 1164 135 1168
rect 139 1164 140 1168
rect 134 1163 140 1164
rect 238 1168 244 1169
rect 238 1164 239 1168
rect 243 1164 244 1168
rect 238 1163 244 1164
rect 374 1168 380 1169
rect 374 1164 375 1168
rect 379 1164 380 1168
rect 374 1163 380 1164
rect 510 1168 516 1169
rect 510 1164 511 1168
rect 515 1164 516 1168
rect 510 1163 516 1164
rect 654 1168 660 1169
rect 654 1164 655 1168
rect 659 1164 660 1168
rect 654 1163 660 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 926 1168 932 1169
rect 926 1164 927 1168
rect 931 1164 932 1168
rect 926 1163 932 1164
rect 1062 1168 1068 1169
rect 1062 1164 1063 1168
rect 1067 1164 1068 1168
rect 1062 1163 1068 1164
rect 1198 1168 1204 1169
rect 1198 1164 1199 1168
rect 1203 1164 1204 1168
rect 1198 1163 1204 1164
rect 1334 1168 1340 1169
rect 1334 1164 1335 1168
rect 1339 1164 1340 1168
rect 1806 1168 1807 1172
rect 1811 1168 1812 1172
rect 1830 1169 1831 1173
rect 1835 1169 1836 1173
rect 1830 1168 1836 1169
rect 1934 1173 1940 1174
rect 1934 1169 1935 1173
rect 1939 1169 1940 1173
rect 1934 1168 1940 1169
rect 2078 1173 2084 1174
rect 2078 1169 2079 1173
rect 2083 1169 2084 1173
rect 2078 1168 2084 1169
rect 2230 1173 2236 1174
rect 2230 1169 2231 1173
rect 2235 1169 2236 1173
rect 2230 1168 2236 1169
rect 2390 1173 2396 1174
rect 2390 1169 2391 1173
rect 2395 1169 2396 1173
rect 2390 1168 2396 1169
rect 2542 1173 2548 1174
rect 2542 1169 2543 1173
rect 2547 1169 2548 1173
rect 2542 1168 2548 1169
rect 2694 1173 2700 1174
rect 2694 1169 2695 1173
rect 2699 1169 2700 1173
rect 2694 1168 2700 1169
rect 2846 1173 2852 1174
rect 2846 1169 2847 1173
rect 2851 1169 2852 1173
rect 2846 1168 2852 1169
rect 2998 1173 3004 1174
rect 2998 1169 2999 1173
rect 3003 1169 3004 1173
rect 2998 1168 3004 1169
rect 3158 1173 3164 1174
rect 3158 1169 3159 1173
rect 3163 1169 3164 1173
rect 3158 1168 3164 1169
rect 3462 1172 3468 1173
rect 3462 1168 3463 1172
rect 3467 1168 3468 1172
rect 1806 1167 1812 1168
rect 3462 1167 3468 1168
rect 1334 1163 1340 1164
rect 1766 1165 1772 1166
rect 110 1160 116 1161
rect 1766 1161 1767 1165
rect 1771 1161 1772 1165
rect 1766 1160 1772 1161
rect 134 1149 140 1150
rect 110 1148 116 1149
rect 110 1144 111 1148
rect 115 1144 116 1148
rect 134 1145 135 1149
rect 139 1145 140 1149
rect 134 1144 140 1145
rect 238 1149 244 1150
rect 238 1145 239 1149
rect 243 1145 244 1149
rect 238 1144 244 1145
rect 374 1149 380 1150
rect 374 1145 375 1149
rect 379 1145 380 1149
rect 374 1144 380 1145
rect 510 1149 516 1150
rect 510 1145 511 1149
rect 515 1145 516 1149
rect 510 1144 516 1145
rect 654 1149 660 1150
rect 654 1145 655 1149
rect 659 1145 660 1149
rect 654 1144 660 1145
rect 790 1149 796 1150
rect 790 1145 791 1149
rect 795 1145 796 1149
rect 790 1144 796 1145
rect 926 1149 932 1150
rect 926 1145 927 1149
rect 931 1145 932 1149
rect 926 1144 932 1145
rect 1062 1149 1068 1150
rect 1062 1145 1063 1149
rect 1067 1145 1068 1149
rect 1062 1144 1068 1145
rect 1198 1149 1204 1150
rect 1198 1145 1199 1149
rect 1203 1145 1204 1149
rect 1198 1144 1204 1145
rect 1334 1149 1340 1150
rect 1334 1145 1335 1149
rect 1339 1145 1340 1149
rect 1334 1144 1340 1145
rect 1766 1148 1772 1149
rect 1766 1144 1767 1148
rect 1771 1144 1772 1148
rect 110 1143 116 1144
rect 1766 1143 1772 1144
rect 1806 1116 1812 1117
rect 3462 1116 3468 1117
rect 1806 1112 1807 1116
rect 1811 1112 1812 1116
rect 1806 1111 1812 1112
rect 1862 1115 1868 1116
rect 1862 1111 1863 1115
rect 1867 1111 1868 1115
rect 1862 1110 1868 1111
rect 1982 1115 1988 1116
rect 1982 1111 1983 1115
rect 1987 1111 1988 1115
rect 1982 1110 1988 1111
rect 2110 1115 2116 1116
rect 2110 1111 2111 1115
rect 2115 1111 2116 1115
rect 2110 1110 2116 1111
rect 2246 1115 2252 1116
rect 2246 1111 2247 1115
rect 2251 1111 2252 1115
rect 2246 1110 2252 1111
rect 2382 1115 2388 1116
rect 2382 1111 2383 1115
rect 2387 1111 2388 1115
rect 2382 1110 2388 1111
rect 2510 1115 2516 1116
rect 2510 1111 2511 1115
rect 2515 1111 2516 1115
rect 2510 1110 2516 1111
rect 2638 1115 2644 1116
rect 2638 1111 2639 1115
rect 2643 1111 2644 1115
rect 2638 1110 2644 1111
rect 2758 1115 2764 1116
rect 2758 1111 2759 1115
rect 2763 1111 2764 1115
rect 2758 1110 2764 1111
rect 2870 1115 2876 1116
rect 2870 1111 2871 1115
rect 2875 1111 2876 1115
rect 2870 1110 2876 1111
rect 2974 1115 2980 1116
rect 2974 1111 2975 1115
rect 2979 1111 2980 1115
rect 2974 1110 2980 1111
rect 3078 1115 3084 1116
rect 3078 1111 3079 1115
rect 3083 1111 3084 1115
rect 3078 1110 3084 1111
rect 3182 1115 3188 1116
rect 3182 1111 3183 1115
rect 3187 1111 3188 1115
rect 3182 1110 3188 1111
rect 3278 1115 3284 1116
rect 3278 1111 3279 1115
rect 3283 1111 3284 1115
rect 3278 1110 3284 1111
rect 3366 1115 3372 1116
rect 3366 1111 3367 1115
rect 3371 1111 3372 1115
rect 3462 1112 3463 1116
rect 3467 1112 3468 1116
rect 3462 1111 3468 1112
rect 3366 1110 3372 1111
rect 110 1100 116 1101
rect 1766 1100 1772 1101
rect 110 1096 111 1100
rect 115 1096 116 1100
rect 110 1095 116 1096
rect 190 1099 196 1100
rect 190 1095 191 1099
rect 195 1095 196 1099
rect 190 1094 196 1095
rect 334 1099 340 1100
rect 334 1095 335 1099
rect 339 1095 340 1099
rect 334 1094 340 1095
rect 494 1099 500 1100
rect 494 1095 495 1099
rect 499 1095 500 1099
rect 494 1094 500 1095
rect 654 1099 660 1100
rect 654 1095 655 1099
rect 659 1095 660 1099
rect 654 1094 660 1095
rect 814 1099 820 1100
rect 814 1095 815 1099
rect 819 1095 820 1099
rect 814 1094 820 1095
rect 966 1099 972 1100
rect 966 1095 967 1099
rect 971 1095 972 1099
rect 966 1094 972 1095
rect 1118 1099 1124 1100
rect 1118 1095 1119 1099
rect 1123 1095 1124 1099
rect 1118 1094 1124 1095
rect 1262 1099 1268 1100
rect 1262 1095 1263 1099
rect 1267 1095 1268 1099
rect 1262 1094 1268 1095
rect 1406 1099 1412 1100
rect 1406 1095 1407 1099
rect 1411 1095 1412 1099
rect 1406 1094 1412 1095
rect 1558 1099 1564 1100
rect 1558 1095 1559 1099
rect 1563 1095 1564 1099
rect 1766 1096 1767 1100
rect 1771 1096 1772 1100
rect 1766 1095 1772 1096
rect 1806 1099 1812 1100
rect 1806 1095 1807 1099
rect 1811 1095 1812 1099
rect 3462 1099 3468 1100
rect 1558 1094 1564 1095
rect 1806 1094 1812 1095
rect 1862 1096 1868 1097
rect 1862 1092 1863 1096
rect 1867 1092 1868 1096
rect 1862 1091 1868 1092
rect 1982 1096 1988 1097
rect 1982 1092 1983 1096
rect 1987 1092 1988 1096
rect 1982 1091 1988 1092
rect 2110 1096 2116 1097
rect 2110 1092 2111 1096
rect 2115 1092 2116 1096
rect 2110 1091 2116 1092
rect 2246 1096 2252 1097
rect 2246 1092 2247 1096
rect 2251 1092 2252 1096
rect 2246 1091 2252 1092
rect 2382 1096 2388 1097
rect 2382 1092 2383 1096
rect 2387 1092 2388 1096
rect 2382 1091 2388 1092
rect 2510 1096 2516 1097
rect 2510 1092 2511 1096
rect 2515 1092 2516 1096
rect 2510 1091 2516 1092
rect 2638 1096 2644 1097
rect 2638 1092 2639 1096
rect 2643 1092 2644 1096
rect 2638 1091 2644 1092
rect 2758 1096 2764 1097
rect 2758 1092 2759 1096
rect 2763 1092 2764 1096
rect 2758 1091 2764 1092
rect 2870 1096 2876 1097
rect 2870 1092 2871 1096
rect 2875 1092 2876 1096
rect 2870 1091 2876 1092
rect 2974 1096 2980 1097
rect 2974 1092 2975 1096
rect 2979 1092 2980 1096
rect 2974 1091 2980 1092
rect 3078 1096 3084 1097
rect 3078 1092 3079 1096
rect 3083 1092 3084 1096
rect 3078 1091 3084 1092
rect 3182 1096 3188 1097
rect 3182 1092 3183 1096
rect 3187 1092 3188 1096
rect 3182 1091 3188 1092
rect 3278 1096 3284 1097
rect 3278 1092 3279 1096
rect 3283 1092 3284 1096
rect 3278 1091 3284 1092
rect 3366 1096 3372 1097
rect 3366 1092 3367 1096
rect 3371 1092 3372 1096
rect 3462 1095 3463 1099
rect 3467 1095 3468 1099
rect 3462 1094 3468 1095
rect 3366 1091 3372 1092
rect 110 1083 116 1084
rect 110 1079 111 1083
rect 115 1079 116 1083
rect 1766 1083 1772 1084
rect 110 1078 116 1079
rect 190 1080 196 1081
rect 190 1076 191 1080
rect 195 1076 196 1080
rect 190 1075 196 1076
rect 334 1080 340 1081
rect 334 1076 335 1080
rect 339 1076 340 1080
rect 334 1075 340 1076
rect 494 1080 500 1081
rect 494 1076 495 1080
rect 499 1076 500 1080
rect 494 1075 500 1076
rect 654 1080 660 1081
rect 654 1076 655 1080
rect 659 1076 660 1080
rect 654 1075 660 1076
rect 814 1080 820 1081
rect 814 1076 815 1080
rect 819 1076 820 1080
rect 814 1075 820 1076
rect 966 1080 972 1081
rect 966 1076 967 1080
rect 971 1076 972 1080
rect 966 1075 972 1076
rect 1118 1080 1124 1081
rect 1118 1076 1119 1080
rect 1123 1076 1124 1080
rect 1118 1075 1124 1076
rect 1262 1080 1268 1081
rect 1262 1076 1263 1080
rect 1267 1076 1268 1080
rect 1262 1075 1268 1076
rect 1406 1080 1412 1081
rect 1406 1076 1407 1080
rect 1411 1076 1412 1080
rect 1406 1075 1412 1076
rect 1558 1080 1564 1081
rect 1558 1076 1559 1080
rect 1563 1076 1564 1080
rect 1766 1079 1767 1083
rect 1771 1079 1772 1083
rect 1766 1078 1772 1079
rect 1558 1075 1564 1076
rect 2102 1044 2108 1045
rect 1806 1041 1812 1042
rect 1806 1037 1807 1041
rect 1811 1037 1812 1041
rect 2102 1040 2103 1044
rect 2107 1040 2108 1044
rect 2102 1039 2108 1040
rect 2190 1044 2196 1045
rect 2190 1040 2191 1044
rect 2195 1040 2196 1044
rect 2190 1039 2196 1040
rect 2278 1044 2284 1045
rect 2278 1040 2279 1044
rect 2283 1040 2284 1044
rect 2278 1039 2284 1040
rect 2366 1044 2372 1045
rect 2366 1040 2367 1044
rect 2371 1040 2372 1044
rect 2366 1039 2372 1040
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2542 1044 2548 1045
rect 2542 1040 2543 1044
rect 2547 1040 2548 1044
rect 2542 1039 2548 1040
rect 2630 1044 2636 1045
rect 2630 1040 2631 1044
rect 2635 1040 2636 1044
rect 2630 1039 2636 1040
rect 2718 1044 2724 1045
rect 2718 1040 2719 1044
rect 2723 1040 2724 1044
rect 2718 1039 2724 1040
rect 2806 1044 2812 1045
rect 2806 1040 2807 1044
rect 2811 1040 2812 1044
rect 2806 1039 2812 1040
rect 3462 1041 3468 1042
rect 1806 1036 1812 1037
rect 3462 1037 3463 1041
rect 3467 1037 3468 1041
rect 3462 1036 3468 1037
rect 326 1028 332 1029
rect 110 1025 116 1026
rect 110 1021 111 1025
rect 115 1021 116 1025
rect 326 1024 327 1028
rect 331 1024 332 1028
rect 326 1023 332 1024
rect 462 1028 468 1029
rect 462 1024 463 1028
rect 467 1024 468 1028
rect 462 1023 468 1024
rect 606 1028 612 1029
rect 606 1024 607 1028
rect 611 1024 612 1028
rect 606 1023 612 1024
rect 766 1028 772 1029
rect 766 1024 767 1028
rect 771 1024 772 1028
rect 766 1023 772 1024
rect 926 1028 932 1029
rect 926 1024 927 1028
rect 931 1024 932 1028
rect 926 1023 932 1024
rect 1078 1028 1084 1029
rect 1078 1024 1079 1028
rect 1083 1024 1084 1028
rect 1078 1023 1084 1024
rect 1230 1028 1236 1029
rect 1230 1024 1231 1028
rect 1235 1024 1236 1028
rect 1230 1023 1236 1024
rect 1382 1028 1388 1029
rect 1382 1024 1383 1028
rect 1387 1024 1388 1028
rect 1382 1023 1388 1024
rect 1534 1028 1540 1029
rect 1534 1024 1535 1028
rect 1539 1024 1540 1028
rect 1534 1023 1540 1024
rect 1670 1028 1676 1029
rect 1670 1024 1671 1028
rect 1675 1024 1676 1028
rect 1670 1023 1676 1024
rect 1766 1025 1772 1026
rect 2102 1025 2108 1026
rect 110 1020 116 1021
rect 1766 1021 1767 1025
rect 1771 1021 1772 1025
rect 1766 1020 1772 1021
rect 1806 1024 1812 1025
rect 1806 1020 1807 1024
rect 1811 1020 1812 1024
rect 2102 1021 2103 1025
rect 2107 1021 2108 1025
rect 2102 1020 2108 1021
rect 2190 1025 2196 1026
rect 2190 1021 2191 1025
rect 2195 1021 2196 1025
rect 2190 1020 2196 1021
rect 2278 1025 2284 1026
rect 2278 1021 2279 1025
rect 2283 1021 2284 1025
rect 2278 1020 2284 1021
rect 2366 1025 2372 1026
rect 2366 1021 2367 1025
rect 2371 1021 2372 1025
rect 2366 1020 2372 1021
rect 2454 1025 2460 1026
rect 2454 1021 2455 1025
rect 2459 1021 2460 1025
rect 2454 1020 2460 1021
rect 2542 1025 2548 1026
rect 2542 1021 2543 1025
rect 2547 1021 2548 1025
rect 2542 1020 2548 1021
rect 2630 1025 2636 1026
rect 2630 1021 2631 1025
rect 2635 1021 2636 1025
rect 2630 1020 2636 1021
rect 2718 1025 2724 1026
rect 2718 1021 2719 1025
rect 2723 1021 2724 1025
rect 2718 1020 2724 1021
rect 2806 1025 2812 1026
rect 2806 1021 2807 1025
rect 2811 1021 2812 1025
rect 2806 1020 2812 1021
rect 3462 1024 3468 1025
rect 3462 1020 3463 1024
rect 3467 1020 3468 1024
rect 1806 1019 1812 1020
rect 3462 1019 3468 1020
rect 326 1009 332 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 326 1005 327 1009
rect 331 1005 332 1009
rect 326 1004 332 1005
rect 462 1009 468 1010
rect 462 1005 463 1009
rect 467 1005 468 1009
rect 462 1004 468 1005
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 926 1009 932 1010
rect 926 1005 927 1009
rect 931 1005 932 1009
rect 926 1004 932 1005
rect 1078 1009 1084 1010
rect 1078 1005 1079 1009
rect 1083 1005 1084 1009
rect 1078 1004 1084 1005
rect 1230 1009 1236 1010
rect 1230 1005 1231 1009
rect 1235 1005 1236 1009
rect 1230 1004 1236 1005
rect 1382 1009 1388 1010
rect 1382 1005 1383 1009
rect 1387 1005 1388 1009
rect 1382 1004 1388 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1670 1009 1676 1010
rect 1670 1005 1671 1009
rect 1675 1005 1676 1009
rect 1670 1004 1676 1005
rect 1766 1008 1772 1009
rect 1766 1004 1767 1008
rect 1771 1004 1772 1008
rect 110 1003 116 1004
rect 1766 1003 1772 1004
rect 1806 980 1812 981
rect 3462 980 3468 981
rect 1806 976 1807 980
rect 1811 976 1812 980
rect 1806 975 1812 976
rect 2310 979 2316 980
rect 2310 975 2311 979
rect 2315 975 2316 979
rect 2310 974 2316 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 2510 979 2516 980
rect 2510 975 2511 979
rect 2515 975 2516 979
rect 2510 974 2516 975
rect 2622 979 2628 980
rect 2622 975 2623 979
rect 2627 975 2628 979
rect 2622 974 2628 975
rect 2750 979 2756 980
rect 2750 975 2751 979
rect 2755 975 2756 979
rect 2750 974 2756 975
rect 2894 979 2900 980
rect 2894 975 2895 979
rect 2899 975 2900 979
rect 2894 974 2900 975
rect 3054 979 3060 980
rect 3054 975 3055 979
rect 3059 975 3060 979
rect 3054 974 3060 975
rect 3222 979 3228 980
rect 3222 975 3223 979
rect 3227 975 3228 979
rect 3222 974 3228 975
rect 3366 979 3372 980
rect 3366 975 3367 979
rect 3371 975 3372 979
rect 3462 976 3463 980
rect 3467 976 3468 980
rect 3462 975 3468 976
rect 3366 974 3372 975
rect 1806 963 1812 964
rect 110 960 116 961
rect 1766 960 1772 961
rect 110 956 111 960
rect 115 956 116 960
rect 110 955 116 956
rect 470 959 476 960
rect 470 955 471 959
rect 475 955 476 959
rect 470 954 476 955
rect 566 959 572 960
rect 566 955 567 959
rect 571 955 572 959
rect 566 954 572 955
rect 670 959 676 960
rect 670 955 671 959
rect 675 955 676 959
rect 670 954 676 955
rect 782 959 788 960
rect 782 955 783 959
rect 787 955 788 959
rect 782 954 788 955
rect 886 959 892 960
rect 886 955 887 959
rect 891 955 892 959
rect 886 954 892 955
rect 990 959 996 960
rect 990 955 991 959
rect 995 955 996 959
rect 990 954 996 955
rect 1094 959 1100 960
rect 1094 955 1095 959
rect 1099 955 1100 959
rect 1094 954 1100 955
rect 1198 959 1204 960
rect 1198 955 1199 959
rect 1203 955 1204 959
rect 1198 954 1204 955
rect 1294 959 1300 960
rect 1294 955 1295 959
rect 1299 955 1300 959
rect 1294 954 1300 955
rect 1390 959 1396 960
rect 1390 955 1391 959
rect 1395 955 1396 959
rect 1390 954 1396 955
rect 1486 959 1492 960
rect 1486 955 1487 959
rect 1491 955 1492 959
rect 1486 954 1492 955
rect 1582 959 1588 960
rect 1582 955 1583 959
rect 1587 955 1588 959
rect 1582 954 1588 955
rect 1670 959 1676 960
rect 1670 955 1671 959
rect 1675 955 1676 959
rect 1766 956 1767 960
rect 1771 956 1772 960
rect 1806 959 1807 963
rect 1811 959 1812 963
rect 3462 963 3468 964
rect 1806 958 1812 959
rect 2310 960 2316 961
rect 1766 955 1772 956
rect 2310 956 2311 960
rect 2315 956 2316 960
rect 2310 955 2316 956
rect 2406 960 2412 961
rect 2406 956 2407 960
rect 2411 956 2412 960
rect 2406 955 2412 956
rect 2510 960 2516 961
rect 2510 956 2511 960
rect 2515 956 2516 960
rect 2510 955 2516 956
rect 2622 960 2628 961
rect 2622 956 2623 960
rect 2627 956 2628 960
rect 2622 955 2628 956
rect 2750 960 2756 961
rect 2750 956 2751 960
rect 2755 956 2756 960
rect 2750 955 2756 956
rect 2894 960 2900 961
rect 2894 956 2895 960
rect 2899 956 2900 960
rect 2894 955 2900 956
rect 3054 960 3060 961
rect 3054 956 3055 960
rect 3059 956 3060 960
rect 3054 955 3060 956
rect 3222 960 3228 961
rect 3222 956 3223 960
rect 3227 956 3228 960
rect 3222 955 3228 956
rect 3366 960 3372 961
rect 3366 956 3367 960
rect 3371 956 3372 960
rect 3462 959 3463 963
rect 3467 959 3468 963
rect 3462 958 3468 959
rect 3366 955 3372 956
rect 1670 954 1676 955
rect 110 943 116 944
rect 110 939 111 943
rect 115 939 116 943
rect 1766 943 1772 944
rect 110 938 116 939
rect 470 940 476 941
rect 470 936 471 940
rect 475 936 476 940
rect 470 935 476 936
rect 566 940 572 941
rect 566 936 567 940
rect 571 936 572 940
rect 566 935 572 936
rect 670 940 676 941
rect 670 936 671 940
rect 675 936 676 940
rect 670 935 676 936
rect 782 940 788 941
rect 782 936 783 940
rect 787 936 788 940
rect 782 935 788 936
rect 886 940 892 941
rect 886 936 887 940
rect 891 936 892 940
rect 886 935 892 936
rect 990 940 996 941
rect 990 936 991 940
rect 995 936 996 940
rect 990 935 996 936
rect 1094 940 1100 941
rect 1094 936 1095 940
rect 1099 936 1100 940
rect 1094 935 1100 936
rect 1198 940 1204 941
rect 1198 936 1199 940
rect 1203 936 1204 940
rect 1198 935 1204 936
rect 1294 940 1300 941
rect 1294 936 1295 940
rect 1299 936 1300 940
rect 1294 935 1300 936
rect 1390 940 1396 941
rect 1390 936 1391 940
rect 1395 936 1396 940
rect 1390 935 1396 936
rect 1486 940 1492 941
rect 1486 936 1487 940
rect 1491 936 1492 940
rect 1486 935 1492 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1670 940 1676 941
rect 1670 936 1671 940
rect 1675 936 1676 940
rect 1766 939 1767 943
rect 1771 939 1772 943
rect 1766 938 1772 939
rect 1670 935 1676 936
rect 1830 904 1836 905
rect 1806 901 1812 902
rect 1806 897 1807 901
rect 1811 897 1812 901
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1982 904 1988 905
rect 1982 900 1983 904
rect 1987 900 1988 904
rect 1982 899 1988 900
rect 2150 904 2156 905
rect 2150 900 2151 904
rect 2155 900 2156 904
rect 2150 899 2156 900
rect 2326 904 2332 905
rect 2326 900 2327 904
rect 2331 900 2332 904
rect 2326 899 2332 900
rect 2518 904 2524 905
rect 2518 900 2519 904
rect 2523 900 2524 904
rect 2518 899 2524 900
rect 2718 904 2724 905
rect 2718 900 2719 904
rect 2723 900 2724 904
rect 2718 899 2724 900
rect 2934 904 2940 905
rect 2934 900 2935 904
rect 2939 900 2940 904
rect 2934 899 2940 900
rect 3158 904 3164 905
rect 3158 900 3159 904
rect 3163 900 3164 904
rect 3158 899 3164 900
rect 3366 904 3372 905
rect 3366 900 3367 904
rect 3371 900 3372 904
rect 3366 899 3372 900
rect 3462 901 3468 902
rect 1806 896 1812 897
rect 3462 897 3463 901
rect 3467 897 3468 901
rect 3462 896 3468 897
rect 606 892 612 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 606 888 607 892
rect 611 888 612 892
rect 606 887 612 888
rect 694 892 700 893
rect 694 888 695 892
rect 699 888 700 892
rect 694 887 700 888
rect 790 892 796 893
rect 790 888 791 892
rect 795 888 796 892
rect 790 887 796 888
rect 894 892 900 893
rect 894 888 895 892
rect 899 888 900 892
rect 894 887 900 888
rect 998 892 1004 893
rect 998 888 999 892
rect 1003 888 1004 892
rect 998 887 1004 888
rect 1110 892 1116 893
rect 1110 888 1111 892
rect 1115 888 1116 892
rect 1110 887 1116 888
rect 1222 892 1228 893
rect 1222 888 1223 892
rect 1227 888 1228 892
rect 1222 887 1228 888
rect 1342 892 1348 893
rect 1342 888 1343 892
rect 1347 888 1348 892
rect 1342 887 1348 888
rect 1462 892 1468 893
rect 1462 888 1463 892
rect 1467 888 1468 892
rect 1462 887 1468 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1582 887 1588 888
rect 1766 889 1772 890
rect 110 884 116 885
rect 1766 885 1767 889
rect 1771 885 1772 889
rect 1830 885 1836 886
rect 1766 884 1772 885
rect 1806 884 1812 885
rect 1806 880 1807 884
rect 1811 880 1812 884
rect 1830 881 1831 885
rect 1835 881 1836 885
rect 1830 880 1836 881
rect 1982 885 1988 886
rect 1982 881 1983 885
rect 1987 881 1988 885
rect 1982 880 1988 881
rect 2150 885 2156 886
rect 2150 881 2151 885
rect 2155 881 2156 885
rect 2150 880 2156 881
rect 2326 885 2332 886
rect 2326 881 2327 885
rect 2331 881 2332 885
rect 2326 880 2332 881
rect 2518 885 2524 886
rect 2518 881 2519 885
rect 2523 881 2524 885
rect 2518 880 2524 881
rect 2718 885 2724 886
rect 2718 881 2719 885
rect 2723 881 2724 885
rect 2718 880 2724 881
rect 2934 885 2940 886
rect 2934 881 2935 885
rect 2939 881 2940 885
rect 2934 880 2940 881
rect 3158 885 3164 886
rect 3158 881 3159 885
rect 3163 881 3164 885
rect 3158 880 3164 881
rect 3366 885 3372 886
rect 3366 881 3367 885
rect 3371 881 3372 885
rect 3366 880 3372 881
rect 3462 884 3468 885
rect 3462 880 3463 884
rect 3467 880 3468 884
rect 1806 879 1812 880
rect 3462 879 3468 880
rect 606 873 612 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 606 869 607 873
rect 611 869 612 873
rect 606 868 612 869
rect 694 873 700 874
rect 694 869 695 873
rect 699 869 700 873
rect 694 868 700 869
rect 790 873 796 874
rect 790 869 791 873
rect 795 869 796 873
rect 790 868 796 869
rect 894 873 900 874
rect 894 869 895 873
rect 899 869 900 873
rect 894 868 900 869
rect 998 873 1004 874
rect 998 869 999 873
rect 1003 869 1004 873
rect 998 868 1004 869
rect 1110 873 1116 874
rect 1110 869 1111 873
rect 1115 869 1116 873
rect 1110 868 1116 869
rect 1222 873 1228 874
rect 1222 869 1223 873
rect 1227 869 1228 873
rect 1222 868 1228 869
rect 1342 873 1348 874
rect 1342 869 1343 873
rect 1347 869 1348 873
rect 1342 868 1348 869
rect 1462 873 1468 874
rect 1462 869 1463 873
rect 1467 869 1468 873
rect 1462 868 1468 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1766 872 1772 873
rect 1766 868 1767 872
rect 1771 868 1772 872
rect 110 867 116 868
rect 1766 867 1772 868
rect 1806 836 1812 837
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 1830 835 1836 836
rect 1830 831 1831 835
rect 1835 831 1836 835
rect 1830 830 1836 831
rect 1958 835 1964 836
rect 1958 831 1959 835
rect 1963 831 1964 835
rect 1958 830 1964 831
rect 2086 835 2092 836
rect 2086 831 2087 835
rect 2091 831 2092 835
rect 2086 830 2092 831
rect 2206 835 2212 836
rect 2206 831 2207 835
rect 2211 831 2212 835
rect 2206 830 2212 831
rect 2326 835 2332 836
rect 2326 831 2327 835
rect 2331 831 2332 835
rect 2326 830 2332 831
rect 2462 835 2468 836
rect 2462 831 2463 835
rect 2467 831 2468 835
rect 2462 830 2468 831
rect 2614 835 2620 836
rect 2614 831 2615 835
rect 2619 831 2620 835
rect 2614 830 2620 831
rect 2790 835 2796 836
rect 2790 831 2791 835
rect 2795 831 2796 835
rect 2790 830 2796 831
rect 2982 835 2988 836
rect 2982 831 2983 835
rect 2987 831 2988 835
rect 2982 830 2988 831
rect 3182 835 3188 836
rect 3182 831 3183 835
rect 3187 831 3188 835
rect 3182 830 3188 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 110 824 116 825
rect 1766 824 1772 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 518 823 524 824
rect 518 819 519 823
rect 523 819 524 823
rect 518 818 524 819
rect 614 823 620 824
rect 614 819 615 823
rect 619 819 620 823
rect 614 818 620 819
rect 718 823 724 824
rect 718 819 719 823
rect 723 819 724 823
rect 718 818 724 819
rect 830 823 836 824
rect 830 819 831 823
rect 835 819 836 823
rect 830 818 836 819
rect 950 823 956 824
rect 950 819 951 823
rect 955 819 956 823
rect 950 818 956 819
rect 1070 823 1076 824
rect 1070 819 1071 823
rect 1075 819 1076 823
rect 1070 818 1076 819
rect 1190 823 1196 824
rect 1190 819 1191 823
rect 1195 819 1196 823
rect 1190 818 1196 819
rect 1310 823 1316 824
rect 1310 819 1311 823
rect 1315 819 1316 823
rect 1310 818 1316 819
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1558 823 1564 824
rect 1558 819 1559 823
rect 1563 819 1564 823
rect 1766 820 1767 824
rect 1771 820 1772 824
rect 1766 819 1772 820
rect 1806 819 1812 820
rect 1558 818 1564 819
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 1830 816 1836 817
rect 1830 812 1831 816
rect 1835 812 1836 816
rect 1830 811 1836 812
rect 1958 816 1964 817
rect 1958 812 1959 816
rect 1963 812 1964 816
rect 1958 811 1964 812
rect 2086 816 2092 817
rect 2086 812 2087 816
rect 2091 812 2092 816
rect 2086 811 2092 812
rect 2206 816 2212 817
rect 2206 812 2207 816
rect 2211 812 2212 816
rect 2206 811 2212 812
rect 2326 816 2332 817
rect 2326 812 2327 816
rect 2331 812 2332 816
rect 2326 811 2332 812
rect 2462 816 2468 817
rect 2462 812 2463 816
rect 2467 812 2468 816
rect 2462 811 2468 812
rect 2614 816 2620 817
rect 2614 812 2615 816
rect 2619 812 2620 816
rect 2614 811 2620 812
rect 2790 816 2796 817
rect 2790 812 2791 816
rect 2795 812 2796 816
rect 2790 811 2796 812
rect 2982 816 2988 817
rect 2982 812 2983 816
rect 2987 812 2988 816
rect 2982 811 2988 812
rect 3182 816 3188 817
rect 3182 812 3183 816
rect 3187 812 3188 816
rect 3182 811 3188 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 1766 807 1772 808
rect 110 802 116 803
rect 518 804 524 805
rect 518 800 519 804
rect 523 800 524 804
rect 518 799 524 800
rect 614 804 620 805
rect 614 800 615 804
rect 619 800 620 804
rect 614 799 620 800
rect 718 804 724 805
rect 718 800 719 804
rect 723 800 724 804
rect 718 799 724 800
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 950 804 956 805
rect 950 800 951 804
rect 955 800 956 804
rect 950 799 956 800
rect 1070 804 1076 805
rect 1070 800 1071 804
rect 1075 800 1076 804
rect 1070 799 1076 800
rect 1190 804 1196 805
rect 1190 800 1191 804
rect 1195 800 1196 804
rect 1190 799 1196 800
rect 1310 804 1316 805
rect 1310 800 1311 804
rect 1315 800 1316 804
rect 1310 799 1316 800
rect 1430 804 1436 805
rect 1430 800 1431 804
rect 1435 800 1436 804
rect 1430 799 1436 800
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1766 803 1767 807
rect 1771 803 1772 807
rect 1766 802 1772 803
rect 1558 799 1564 800
rect 1878 768 1884 769
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 1878 764 1879 768
rect 1883 764 1884 768
rect 1878 763 1884 764
rect 2014 768 2020 769
rect 2014 764 2015 768
rect 2019 764 2020 768
rect 2014 763 2020 764
rect 2150 768 2156 769
rect 2150 764 2151 768
rect 2155 764 2156 768
rect 2150 763 2156 764
rect 2286 768 2292 769
rect 2286 764 2287 768
rect 2291 764 2292 768
rect 2286 763 2292 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 1806 760 1812 761
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 382 756 388 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 470 756 476 757
rect 470 752 471 756
rect 475 752 476 756
rect 470 751 476 752
rect 574 756 580 757
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 678 756 684 757
rect 678 752 679 756
rect 683 752 684 756
rect 678 751 684 752
rect 790 756 796 757
rect 790 752 791 756
rect 795 752 796 756
rect 790 751 796 752
rect 910 756 916 757
rect 910 752 911 756
rect 915 752 916 756
rect 910 751 916 752
rect 1030 756 1036 757
rect 1030 752 1031 756
rect 1035 752 1036 756
rect 1030 751 1036 752
rect 1158 756 1164 757
rect 1158 752 1159 756
rect 1163 752 1164 756
rect 1158 751 1164 752
rect 1286 756 1292 757
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1414 756 1420 757
rect 1414 752 1415 756
rect 1419 752 1420 756
rect 1414 751 1420 752
rect 1766 753 1772 754
rect 110 748 116 749
rect 1766 749 1767 753
rect 1771 749 1772 753
rect 1878 749 1884 750
rect 1766 748 1772 749
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1878 745 1879 749
rect 1883 745 1884 749
rect 1878 744 1884 745
rect 2014 749 2020 750
rect 2014 745 2015 749
rect 2019 745 2020 749
rect 2014 744 2020 745
rect 2150 749 2156 750
rect 2150 745 2151 749
rect 2155 745 2156 749
rect 2150 744 2156 745
rect 2286 749 2292 750
rect 2286 745 2287 749
rect 2291 745 2292 749
rect 2286 744 2292 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1806 743 1812 744
rect 3462 743 3468 744
rect 382 737 388 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 382 733 383 737
rect 387 733 388 737
rect 382 732 388 733
rect 470 737 476 738
rect 470 733 471 737
rect 475 733 476 737
rect 470 732 476 733
rect 574 737 580 738
rect 574 733 575 737
rect 579 733 580 737
rect 574 732 580 733
rect 678 737 684 738
rect 678 733 679 737
rect 683 733 684 737
rect 678 732 684 733
rect 790 737 796 738
rect 790 733 791 737
rect 795 733 796 737
rect 790 732 796 733
rect 910 737 916 738
rect 910 733 911 737
rect 915 733 916 737
rect 910 732 916 733
rect 1030 737 1036 738
rect 1030 733 1031 737
rect 1035 733 1036 737
rect 1030 732 1036 733
rect 1158 737 1164 738
rect 1158 733 1159 737
rect 1163 733 1164 737
rect 1158 732 1164 733
rect 1286 737 1292 738
rect 1286 733 1287 737
rect 1291 733 1292 737
rect 1286 732 1292 733
rect 1414 737 1420 738
rect 1414 733 1415 737
rect 1419 733 1420 737
rect 1414 732 1420 733
rect 1766 736 1772 737
rect 1766 732 1767 736
rect 1771 732 1772 736
rect 110 731 116 732
rect 1766 731 1772 732
rect 1806 700 1812 701
rect 3462 700 3468 701
rect 1806 696 1807 700
rect 1811 696 1812 700
rect 1806 695 1812 696
rect 1830 699 1836 700
rect 1830 695 1831 699
rect 1835 695 1836 699
rect 1830 694 1836 695
rect 1950 699 1956 700
rect 1950 695 1951 699
rect 1955 695 1956 699
rect 1950 694 1956 695
rect 2102 699 2108 700
rect 2102 695 2103 699
rect 2107 695 2108 699
rect 2102 694 2108 695
rect 2262 699 2268 700
rect 2262 695 2263 699
rect 2267 695 2268 699
rect 2262 694 2268 695
rect 2414 699 2420 700
rect 2414 695 2415 699
rect 2419 695 2420 699
rect 2414 694 2420 695
rect 2566 699 2572 700
rect 2566 695 2567 699
rect 2571 695 2572 699
rect 2566 694 2572 695
rect 2718 699 2724 700
rect 2718 695 2719 699
rect 2723 695 2724 699
rect 2718 694 2724 695
rect 2878 699 2884 700
rect 2878 695 2879 699
rect 2883 695 2884 699
rect 2878 694 2884 695
rect 3038 699 3044 700
rect 3038 695 3039 699
rect 3043 695 3044 699
rect 3038 694 3044 695
rect 3198 699 3204 700
rect 3198 695 3199 699
rect 3203 695 3204 699
rect 3462 696 3463 700
rect 3467 696 3468 700
rect 3462 695 3468 696
rect 3198 694 3204 695
rect 110 684 116 685
rect 1766 684 1772 685
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 246 683 252 684
rect 246 679 247 683
rect 251 679 252 683
rect 246 678 252 679
rect 342 683 348 684
rect 342 679 343 683
rect 347 679 348 683
rect 342 678 348 679
rect 454 683 460 684
rect 454 679 455 683
rect 459 679 460 683
rect 454 678 460 679
rect 566 683 572 684
rect 566 679 567 683
rect 571 679 572 683
rect 566 678 572 679
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 830 683 836 684
rect 830 679 831 683
rect 835 679 836 683
rect 830 678 836 679
rect 982 683 988 684
rect 982 679 983 683
rect 987 679 988 683
rect 982 678 988 679
rect 1150 683 1156 684
rect 1150 679 1151 683
rect 1155 679 1156 683
rect 1150 678 1156 679
rect 1326 683 1332 684
rect 1326 679 1327 683
rect 1331 679 1332 683
rect 1326 678 1332 679
rect 1510 683 1516 684
rect 1510 679 1511 683
rect 1515 679 1516 683
rect 1510 678 1516 679
rect 1670 683 1676 684
rect 1670 679 1671 683
rect 1675 679 1676 683
rect 1766 680 1767 684
rect 1771 680 1772 684
rect 1766 679 1772 680
rect 1806 683 1812 684
rect 1806 679 1807 683
rect 1811 679 1812 683
rect 3462 683 3468 684
rect 1670 678 1676 679
rect 1806 678 1812 679
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1950 680 1956 681
rect 1950 676 1951 680
rect 1955 676 1956 680
rect 1950 675 1956 676
rect 2102 680 2108 681
rect 2102 676 2103 680
rect 2107 676 2108 680
rect 2102 675 2108 676
rect 2262 680 2268 681
rect 2262 676 2263 680
rect 2267 676 2268 680
rect 2262 675 2268 676
rect 2414 680 2420 681
rect 2414 676 2415 680
rect 2419 676 2420 680
rect 2414 675 2420 676
rect 2566 680 2572 681
rect 2566 676 2567 680
rect 2571 676 2572 680
rect 2566 675 2572 676
rect 2718 680 2724 681
rect 2718 676 2719 680
rect 2723 676 2724 680
rect 2718 675 2724 676
rect 2878 680 2884 681
rect 2878 676 2879 680
rect 2883 676 2884 680
rect 2878 675 2884 676
rect 3038 680 3044 681
rect 3038 676 3039 680
rect 3043 676 3044 680
rect 3038 675 3044 676
rect 3198 680 3204 681
rect 3198 676 3199 680
rect 3203 676 3204 680
rect 3462 679 3463 683
rect 3467 679 3468 683
rect 3462 678 3468 679
rect 3198 675 3204 676
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 1766 667 1772 668
rect 110 662 116 663
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 342 664 348 665
rect 342 660 343 664
rect 347 660 348 664
rect 342 659 348 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 566 664 572 665
rect 566 660 567 664
rect 571 660 572 664
rect 566 659 572 660
rect 694 664 700 665
rect 694 660 695 664
rect 699 660 700 664
rect 694 659 700 660
rect 830 664 836 665
rect 830 660 831 664
rect 835 660 836 664
rect 830 659 836 660
rect 982 664 988 665
rect 982 660 983 664
rect 987 660 988 664
rect 982 659 988 660
rect 1150 664 1156 665
rect 1150 660 1151 664
rect 1155 660 1156 664
rect 1150 659 1156 660
rect 1326 664 1332 665
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1510 664 1516 665
rect 1510 660 1511 664
rect 1515 660 1516 664
rect 1510 659 1516 660
rect 1670 664 1676 665
rect 1670 660 1671 664
rect 1675 660 1676 664
rect 1766 663 1767 667
rect 1771 663 1772 667
rect 1766 662 1772 663
rect 1670 659 1676 660
rect 1974 636 1980 637
rect 1806 633 1812 634
rect 1806 629 1807 633
rect 1811 629 1812 633
rect 1974 632 1975 636
rect 1979 632 1980 636
rect 1974 631 1980 632
rect 2238 636 2244 637
rect 2238 632 2239 636
rect 2243 632 2244 636
rect 2238 631 2244 632
rect 2478 636 2484 637
rect 2478 632 2479 636
rect 2483 632 2484 636
rect 2478 631 2484 632
rect 2686 636 2692 637
rect 2686 632 2687 636
rect 2691 632 2692 636
rect 2686 631 2692 632
rect 2878 636 2884 637
rect 2878 632 2879 636
rect 2883 632 2884 636
rect 2878 631 2884 632
rect 3054 636 3060 637
rect 3054 632 3055 636
rect 3059 632 3060 636
rect 3054 631 3060 632
rect 3222 636 3228 637
rect 3222 632 3223 636
rect 3227 632 3228 636
rect 3222 631 3228 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3366 631 3372 632
rect 3462 633 3468 634
rect 1806 628 1812 629
rect 3462 629 3463 633
rect 3467 629 3468 633
rect 3462 628 3468 629
rect 1974 617 1980 618
rect 134 616 140 617
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 134 612 135 616
rect 139 612 140 616
rect 134 611 140 612
rect 230 616 236 617
rect 230 612 231 616
rect 235 612 236 616
rect 230 611 236 612
rect 358 616 364 617
rect 358 612 359 616
rect 363 612 364 616
rect 358 611 364 612
rect 486 616 492 617
rect 486 612 487 616
rect 491 612 492 616
rect 486 611 492 612
rect 622 616 628 617
rect 622 612 623 616
rect 627 612 628 616
rect 622 611 628 612
rect 766 616 772 617
rect 766 612 767 616
rect 771 612 772 616
rect 766 611 772 612
rect 910 616 916 617
rect 910 612 911 616
rect 915 612 916 616
rect 910 611 916 612
rect 1054 616 1060 617
rect 1054 612 1055 616
rect 1059 612 1060 616
rect 1054 611 1060 612
rect 1206 616 1212 617
rect 1206 612 1207 616
rect 1211 612 1212 616
rect 1206 611 1212 612
rect 1366 616 1372 617
rect 1366 612 1367 616
rect 1371 612 1372 616
rect 1366 611 1372 612
rect 1526 616 1532 617
rect 1526 612 1527 616
rect 1531 612 1532 616
rect 1526 611 1532 612
rect 1670 616 1676 617
rect 1670 612 1671 616
rect 1675 612 1676 616
rect 1806 616 1812 617
rect 1670 611 1676 612
rect 1766 613 1772 614
rect 110 608 116 609
rect 1766 609 1767 613
rect 1771 609 1772 613
rect 1806 612 1807 616
rect 1811 612 1812 616
rect 1974 613 1975 617
rect 1979 613 1980 617
rect 1974 612 1980 613
rect 2238 617 2244 618
rect 2238 613 2239 617
rect 2243 613 2244 617
rect 2238 612 2244 613
rect 2478 617 2484 618
rect 2478 613 2479 617
rect 2483 613 2484 617
rect 2478 612 2484 613
rect 2686 617 2692 618
rect 2686 613 2687 617
rect 2691 613 2692 617
rect 2686 612 2692 613
rect 2878 617 2884 618
rect 2878 613 2879 617
rect 2883 613 2884 617
rect 2878 612 2884 613
rect 3054 617 3060 618
rect 3054 613 3055 617
rect 3059 613 3060 617
rect 3054 612 3060 613
rect 3222 617 3228 618
rect 3222 613 3223 617
rect 3227 613 3228 617
rect 3222 612 3228 613
rect 3366 617 3372 618
rect 3366 613 3367 617
rect 3371 613 3372 617
rect 3366 612 3372 613
rect 3462 616 3468 617
rect 3462 612 3463 616
rect 3467 612 3468 616
rect 1806 611 1812 612
rect 3462 611 3468 612
rect 1766 608 1772 609
rect 134 597 140 598
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 134 593 135 597
rect 139 593 140 597
rect 134 592 140 593
rect 230 597 236 598
rect 230 593 231 597
rect 235 593 236 597
rect 230 592 236 593
rect 358 597 364 598
rect 358 593 359 597
rect 363 593 364 597
rect 358 592 364 593
rect 486 597 492 598
rect 486 593 487 597
rect 491 593 492 597
rect 486 592 492 593
rect 622 597 628 598
rect 622 593 623 597
rect 627 593 628 597
rect 622 592 628 593
rect 766 597 772 598
rect 766 593 767 597
rect 771 593 772 597
rect 766 592 772 593
rect 910 597 916 598
rect 910 593 911 597
rect 915 593 916 597
rect 910 592 916 593
rect 1054 597 1060 598
rect 1054 593 1055 597
rect 1059 593 1060 597
rect 1054 592 1060 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1366 597 1372 598
rect 1366 593 1367 597
rect 1371 593 1372 597
rect 1366 592 1372 593
rect 1526 597 1532 598
rect 1526 593 1527 597
rect 1531 593 1532 597
rect 1526 592 1532 593
rect 1670 597 1676 598
rect 1670 593 1671 597
rect 1675 593 1676 597
rect 1670 592 1676 593
rect 1766 596 1772 597
rect 1766 592 1767 596
rect 1771 592 1772 596
rect 110 591 116 592
rect 1766 591 1772 592
rect 1806 564 1812 565
rect 3462 564 3468 565
rect 1806 560 1807 564
rect 1811 560 1812 564
rect 1806 559 1812 560
rect 1894 563 1900 564
rect 1894 559 1895 563
rect 1899 559 1900 563
rect 1894 558 1900 559
rect 2014 563 2020 564
rect 2014 559 2015 563
rect 2019 559 2020 563
rect 2014 558 2020 559
rect 2142 563 2148 564
rect 2142 559 2143 563
rect 2147 559 2148 563
rect 2142 558 2148 559
rect 2278 563 2284 564
rect 2278 559 2279 563
rect 2283 559 2284 563
rect 2278 558 2284 559
rect 2422 563 2428 564
rect 2422 559 2423 563
rect 2427 559 2428 563
rect 2422 558 2428 559
rect 2566 563 2572 564
rect 2566 559 2567 563
rect 2571 559 2572 563
rect 2566 558 2572 559
rect 2718 563 2724 564
rect 2718 559 2719 563
rect 2723 559 2724 563
rect 2718 558 2724 559
rect 2870 563 2876 564
rect 2870 559 2871 563
rect 2875 559 2876 563
rect 2870 558 2876 559
rect 3030 563 3036 564
rect 3030 559 3031 563
rect 3035 559 3036 563
rect 3030 558 3036 559
rect 3198 563 3204 564
rect 3198 559 3199 563
rect 3203 559 3204 563
rect 3198 558 3204 559
rect 3366 563 3372 564
rect 3366 559 3367 563
rect 3371 559 3372 563
rect 3462 560 3463 564
rect 3467 560 3468 564
rect 3462 559 3468 560
rect 3366 558 3372 559
rect 110 548 116 549
rect 1766 548 1772 549
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 134 547 140 548
rect 134 543 135 547
rect 139 543 140 547
rect 134 542 140 543
rect 246 547 252 548
rect 246 543 247 547
rect 251 543 252 547
rect 246 542 252 543
rect 406 547 412 548
rect 406 543 407 547
rect 411 543 412 547
rect 406 542 412 543
rect 582 547 588 548
rect 582 543 583 547
rect 587 543 588 547
rect 582 542 588 543
rect 766 547 772 548
rect 766 543 767 547
rect 771 543 772 547
rect 766 542 772 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 1134 542 1140 543
rect 1318 547 1324 548
rect 1318 543 1319 547
rect 1323 543 1324 547
rect 1318 542 1324 543
rect 1502 547 1508 548
rect 1502 543 1503 547
rect 1507 543 1508 547
rect 1502 542 1508 543
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1766 544 1767 548
rect 1771 544 1772 548
rect 1766 543 1772 544
rect 1806 547 1812 548
rect 1806 543 1807 547
rect 1811 543 1812 547
rect 3462 547 3468 548
rect 1670 542 1676 543
rect 1806 542 1812 543
rect 1894 544 1900 545
rect 1894 540 1895 544
rect 1899 540 1900 544
rect 1894 539 1900 540
rect 2014 544 2020 545
rect 2014 540 2015 544
rect 2019 540 2020 544
rect 2014 539 2020 540
rect 2142 544 2148 545
rect 2142 540 2143 544
rect 2147 540 2148 544
rect 2142 539 2148 540
rect 2278 544 2284 545
rect 2278 540 2279 544
rect 2283 540 2284 544
rect 2278 539 2284 540
rect 2422 544 2428 545
rect 2422 540 2423 544
rect 2427 540 2428 544
rect 2422 539 2428 540
rect 2566 544 2572 545
rect 2566 540 2567 544
rect 2571 540 2572 544
rect 2566 539 2572 540
rect 2718 544 2724 545
rect 2718 540 2719 544
rect 2723 540 2724 544
rect 2718 539 2724 540
rect 2870 544 2876 545
rect 2870 540 2871 544
rect 2875 540 2876 544
rect 2870 539 2876 540
rect 3030 544 3036 545
rect 3030 540 3031 544
rect 3035 540 3036 544
rect 3030 539 3036 540
rect 3198 544 3204 545
rect 3198 540 3199 544
rect 3203 540 3204 544
rect 3198 539 3204 540
rect 3366 544 3372 545
rect 3366 540 3367 544
rect 3371 540 3372 544
rect 3462 543 3463 547
rect 3467 543 3468 547
rect 3462 542 3468 543
rect 3366 539 3372 540
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 1766 531 1772 532
rect 110 526 116 527
rect 134 528 140 529
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 246 528 252 529
rect 246 524 247 528
rect 251 524 252 528
rect 246 523 252 524
rect 406 528 412 529
rect 406 524 407 528
rect 411 524 412 528
rect 406 523 412 524
rect 582 528 588 529
rect 582 524 583 528
rect 587 524 588 528
rect 582 523 588 524
rect 766 528 772 529
rect 766 524 767 528
rect 771 524 772 528
rect 766 523 772 524
rect 950 528 956 529
rect 950 524 951 528
rect 955 524 956 528
rect 950 523 956 524
rect 1134 528 1140 529
rect 1134 524 1135 528
rect 1139 524 1140 528
rect 1134 523 1140 524
rect 1318 528 1324 529
rect 1318 524 1319 528
rect 1323 524 1324 528
rect 1318 523 1324 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1670 528 1676 529
rect 1670 524 1671 528
rect 1675 524 1676 528
rect 1766 527 1767 531
rect 1771 527 1772 531
rect 1766 526 1772 527
rect 1670 523 1676 524
rect 2134 496 2140 497
rect 1806 493 1812 494
rect 1806 489 1807 493
rect 1811 489 1812 493
rect 2134 492 2135 496
rect 2139 492 2140 496
rect 2134 491 2140 492
rect 2238 496 2244 497
rect 2238 492 2239 496
rect 2243 492 2244 496
rect 2238 491 2244 492
rect 2358 496 2364 497
rect 2358 492 2359 496
rect 2363 492 2364 496
rect 2358 491 2364 492
rect 2486 496 2492 497
rect 2486 492 2487 496
rect 2491 492 2492 496
rect 2486 491 2492 492
rect 2614 496 2620 497
rect 2614 492 2615 496
rect 2619 492 2620 496
rect 2614 491 2620 492
rect 2750 496 2756 497
rect 2750 492 2751 496
rect 2755 492 2756 496
rect 2750 491 2756 492
rect 2878 496 2884 497
rect 2878 492 2879 496
rect 2883 492 2884 496
rect 2878 491 2884 492
rect 3006 496 3012 497
rect 3006 492 3007 496
rect 3011 492 3012 496
rect 3006 491 3012 492
rect 3134 496 3140 497
rect 3134 492 3135 496
rect 3139 492 3140 496
rect 3134 491 3140 492
rect 3262 496 3268 497
rect 3262 492 3263 496
rect 3267 492 3268 496
rect 3262 491 3268 492
rect 3366 496 3372 497
rect 3366 492 3367 496
rect 3371 492 3372 496
rect 3366 491 3372 492
rect 3462 493 3468 494
rect 1806 488 1812 489
rect 3462 489 3463 493
rect 3467 489 3468 493
rect 3462 488 3468 489
rect 246 480 252 481
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 246 476 247 480
rect 251 476 252 480
rect 246 475 252 476
rect 398 480 404 481
rect 398 476 399 480
rect 403 476 404 480
rect 398 475 404 476
rect 566 480 572 481
rect 566 476 567 480
rect 571 476 572 480
rect 566 475 572 476
rect 734 480 740 481
rect 734 476 735 480
rect 739 476 740 480
rect 734 475 740 476
rect 902 480 908 481
rect 902 476 903 480
rect 907 476 908 480
rect 902 475 908 476
rect 1062 480 1068 481
rect 1062 476 1063 480
rect 1067 476 1068 480
rect 1062 475 1068 476
rect 1222 480 1228 481
rect 1222 476 1223 480
rect 1227 476 1228 480
rect 1222 475 1228 476
rect 1374 480 1380 481
rect 1374 476 1375 480
rect 1379 476 1380 480
rect 1374 475 1380 476
rect 1526 480 1532 481
rect 1526 476 1527 480
rect 1531 476 1532 480
rect 1526 475 1532 476
rect 1670 480 1676 481
rect 1670 476 1671 480
rect 1675 476 1676 480
rect 1670 475 1676 476
rect 1766 477 1772 478
rect 2134 477 2140 478
rect 110 472 116 473
rect 1766 473 1767 477
rect 1771 473 1772 477
rect 1766 472 1772 473
rect 1806 476 1812 477
rect 1806 472 1807 476
rect 1811 472 1812 476
rect 2134 473 2135 477
rect 2139 473 2140 477
rect 2134 472 2140 473
rect 2238 477 2244 478
rect 2238 473 2239 477
rect 2243 473 2244 477
rect 2238 472 2244 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 2486 477 2492 478
rect 2486 473 2487 477
rect 2491 473 2492 477
rect 2486 472 2492 473
rect 2614 477 2620 478
rect 2614 473 2615 477
rect 2619 473 2620 477
rect 2614 472 2620 473
rect 2750 477 2756 478
rect 2750 473 2751 477
rect 2755 473 2756 477
rect 2750 472 2756 473
rect 2878 477 2884 478
rect 2878 473 2879 477
rect 2883 473 2884 477
rect 2878 472 2884 473
rect 3006 477 3012 478
rect 3006 473 3007 477
rect 3011 473 3012 477
rect 3006 472 3012 473
rect 3134 477 3140 478
rect 3134 473 3135 477
rect 3139 473 3140 477
rect 3134 472 3140 473
rect 3262 477 3268 478
rect 3262 473 3263 477
rect 3267 473 3268 477
rect 3262 472 3268 473
rect 3366 477 3372 478
rect 3366 473 3367 477
rect 3371 473 3372 477
rect 3366 472 3372 473
rect 3462 476 3468 477
rect 3462 472 3463 476
rect 3467 472 3468 476
rect 1806 471 1812 472
rect 3462 471 3468 472
rect 246 461 252 462
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 246 457 247 461
rect 251 457 252 461
rect 246 456 252 457
rect 398 461 404 462
rect 398 457 399 461
rect 403 457 404 461
rect 398 456 404 457
rect 566 461 572 462
rect 566 457 567 461
rect 571 457 572 461
rect 566 456 572 457
rect 734 461 740 462
rect 734 457 735 461
rect 739 457 740 461
rect 734 456 740 457
rect 902 461 908 462
rect 902 457 903 461
rect 907 457 908 461
rect 902 456 908 457
rect 1062 461 1068 462
rect 1062 457 1063 461
rect 1067 457 1068 461
rect 1062 456 1068 457
rect 1222 461 1228 462
rect 1222 457 1223 461
rect 1227 457 1228 461
rect 1222 456 1228 457
rect 1374 461 1380 462
rect 1374 457 1375 461
rect 1379 457 1380 461
rect 1374 456 1380 457
rect 1526 461 1532 462
rect 1526 457 1527 461
rect 1531 457 1532 461
rect 1526 456 1532 457
rect 1670 461 1676 462
rect 1670 457 1671 461
rect 1675 457 1676 461
rect 1670 456 1676 457
rect 1766 460 1772 461
rect 1766 456 1767 460
rect 1771 456 1772 460
rect 110 455 116 456
rect 1766 455 1772 456
rect 1806 424 1812 425
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 2238 423 2244 424
rect 2238 419 2239 423
rect 2243 419 2244 423
rect 2238 418 2244 419
rect 2334 423 2340 424
rect 2334 419 2335 423
rect 2339 419 2340 423
rect 2334 418 2340 419
rect 2446 423 2452 424
rect 2446 419 2447 423
rect 2451 419 2452 423
rect 2446 418 2452 419
rect 2558 423 2564 424
rect 2558 419 2559 423
rect 2563 419 2564 423
rect 2558 418 2564 419
rect 2678 423 2684 424
rect 2678 419 2679 423
rect 2683 419 2684 423
rect 2678 418 2684 419
rect 2798 423 2804 424
rect 2798 419 2799 423
rect 2803 419 2804 423
rect 2798 418 2804 419
rect 2910 423 2916 424
rect 2910 419 2911 423
rect 2915 419 2916 423
rect 2910 418 2916 419
rect 3022 423 3028 424
rect 3022 419 3023 423
rect 3027 419 3028 423
rect 3022 418 3028 419
rect 3142 423 3148 424
rect 3142 419 3143 423
rect 3147 419 3148 423
rect 3142 418 3148 419
rect 3262 423 3268 424
rect 3262 419 3263 423
rect 3267 419 3268 423
rect 3262 418 3268 419
rect 3366 423 3372 424
rect 3366 419 3367 423
rect 3371 419 3372 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3366 418 3372 419
rect 110 412 116 413
rect 1766 412 1772 413
rect 110 408 111 412
rect 115 408 116 412
rect 110 407 116 408
rect 518 411 524 412
rect 518 407 519 411
rect 523 407 524 411
rect 518 406 524 407
rect 614 411 620 412
rect 614 407 615 411
rect 619 407 620 411
rect 614 406 620 407
rect 718 411 724 412
rect 718 407 719 411
rect 723 407 724 411
rect 718 406 724 407
rect 822 411 828 412
rect 822 407 823 411
rect 827 407 828 411
rect 822 406 828 407
rect 926 411 932 412
rect 926 407 927 411
rect 931 407 932 411
rect 926 406 932 407
rect 1022 411 1028 412
rect 1022 407 1023 411
rect 1027 407 1028 411
rect 1022 406 1028 407
rect 1126 411 1132 412
rect 1126 407 1127 411
rect 1131 407 1132 411
rect 1126 406 1132 407
rect 1230 411 1236 412
rect 1230 407 1231 411
rect 1235 407 1236 411
rect 1230 406 1236 407
rect 1334 411 1340 412
rect 1334 407 1335 411
rect 1339 407 1340 411
rect 1334 406 1340 407
rect 1438 411 1444 412
rect 1438 407 1439 411
rect 1443 407 1444 411
rect 1766 408 1767 412
rect 1771 408 1772 412
rect 1766 407 1772 408
rect 1806 407 1812 408
rect 1438 406 1444 407
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 3462 407 3468 408
rect 1806 402 1812 403
rect 2238 404 2244 405
rect 2238 400 2239 404
rect 2243 400 2244 404
rect 2238 399 2244 400
rect 2334 404 2340 405
rect 2334 400 2335 404
rect 2339 400 2340 404
rect 2334 399 2340 400
rect 2446 404 2452 405
rect 2446 400 2447 404
rect 2451 400 2452 404
rect 2446 399 2452 400
rect 2558 404 2564 405
rect 2558 400 2559 404
rect 2563 400 2564 404
rect 2558 399 2564 400
rect 2678 404 2684 405
rect 2678 400 2679 404
rect 2683 400 2684 404
rect 2678 399 2684 400
rect 2798 404 2804 405
rect 2798 400 2799 404
rect 2803 400 2804 404
rect 2798 399 2804 400
rect 2910 404 2916 405
rect 2910 400 2911 404
rect 2915 400 2916 404
rect 2910 399 2916 400
rect 3022 404 3028 405
rect 3022 400 3023 404
rect 3027 400 3028 404
rect 3022 399 3028 400
rect 3142 404 3148 405
rect 3142 400 3143 404
rect 3147 400 3148 404
rect 3142 399 3148 400
rect 3262 404 3268 405
rect 3262 400 3263 404
rect 3267 400 3268 404
rect 3262 399 3268 400
rect 3366 404 3372 405
rect 3366 400 3367 404
rect 3371 400 3372 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3366 399 3372 400
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 1766 395 1772 396
rect 110 390 116 391
rect 518 392 524 393
rect 518 388 519 392
rect 523 388 524 392
rect 518 387 524 388
rect 614 392 620 393
rect 614 388 615 392
rect 619 388 620 392
rect 614 387 620 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 822 392 828 393
rect 822 388 823 392
rect 827 388 828 392
rect 822 387 828 388
rect 926 392 932 393
rect 926 388 927 392
rect 931 388 932 392
rect 926 387 932 388
rect 1022 392 1028 393
rect 1022 388 1023 392
rect 1027 388 1028 392
rect 1022 387 1028 388
rect 1126 392 1132 393
rect 1126 388 1127 392
rect 1131 388 1132 392
rect 1126 387 1132 388
rect 1230 392 1236 393
rect 1230 388 1231 392
rect 1235 388 1236 392
rect 1230 387 1236 388
rect 1334 392 1340 393
rect 1334 388 1335 392
rect 1339 388 1340 392
rect 1334 387 1340 388
rect 1438 392 1444 393
rect 1438 388 1439 392
rect 1443 388 1444 392
rect 1766 391 1767 395
rect 1771 391 1772 395
rect 1766 390 1772 391
rect 1438 387 1444 388
rect 2062 356 2068 357
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 2062 352 2063 356
rect 2067 352 2068 356
rect 2062 351 2068 352
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2246 356 2252 357
rect 2246 352 2247 356
rect 2251 352 2252 356
rect 2246 351 2252 352
rect 2358 356 2364 357
rect 2358 352 2359 356
rect 2363 352 2364 356
rect 2358 351 2364 352
rect 2478 356 2484 357
rect 2478 352 2479 356
rect 2483 352 2484 356
rect 2478 351 2484 352
rect 2614 356 2620 357
rect 2614 352 2615 356
rect 2619 352 2620 356
rect 2614 351 2620 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2910 356 2916 357
rect 2910 352 2911 356
rect 2915 352 2916 356
rect 2910 351 2916 352
rect 3062 356 3068 357
rect 3062 352 3063 356
rect 3067 352 3068 356
rect 3062 351 3068 352
rect 3222 356 3228 357
rect 3222 352 3223 356
rect 3227 352 3228 356
rect 3222 351 3228 352
rect 3366 356 3372 357
rect 3366 352 3367 356
rect 3371 352 3372 356
rect 3366 351 3372 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 470 344 476 345
rect 110 341 116 342
rect 110 337 111 341
rect 115 337 116 341
rect 470 340 471 344
rect 475 340 476 344
rect 470 339 476 340
rect 558 344 564 345
rect 558 340 559 344
rect 563 340 564 344
rect 558 339 564 340
rect 646 344 652 345
rect 646 340 647 344
rect 651 340 652 344
rect 646 339 652 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 822 344 828 345
rect 822 340 823 344
rect 827 340 828 344
rect 822 339 828 340
rect 910 344 916 345
rect 910 340 911 344
rect 915 340 916 344
rect 910 339 916 340
rect 998 344 1004 345
rect 998 340 999 344
rect 1003 340 1004 344
rect 998 339 1004 340
rect 1086 344 1092 345
rect 1086 340 1087 344
rect 1091 340 1092 344
rect 1086 339 1092 340
rect 1174 344 1180 345
rect 1174 340 1175 344
rect 1179 340 1180 344
rect 1174 339 1180 340
rect 1262 344 1268 345
rect 1262 340 1263 344
rect 1267 340 1268 344
rect 1262 339 1268 340
rect 1766 341 1772 342
rect 110 336 116 337
rect 1766 337 1767 341
rect 1771 337 1772 341
rect 2062 337 2068 338
rect 1766 336 1772 337
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 2062 333 2063 337
rect 2067 333 2068 337
rect 2062 332 2068 333
rect 2150 337 2156 338
rect 2150 333 2151 337
rect 2155 333 2156 337
rect 2150 332 2156 333
rect 2246 337 2252 338
rect 2246 333 2247 337
rect 2251 333 2252 337
rect 2246 332 2252 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 2478 337 2484 338
rect 2478 333 2479 337
rect 2483 333 2484 337
rect 2478 332 2484 333
rect 2614 337 2620 338
rect 2614 333 2615 337
rect 2619 333 2620 337
rect 2614 332 2620 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2910 337 2916 338
rect 2910 333 2911 337
rect 2915 333 2916 337
rect 2910 332 2916 333
rect 3062 337 3068 338
rect 3062 333 3063 337
rect 3067 333 3068 337
rect 3062 332 3068 333
rect 3222 337 3228 338
rect 3222 333 3223 337
rect 3227 333 3228 337
rect 3222 332 3228 333
rect 3366 337 3372 338
rect 3366 333 3367 337
rect 3371 333 3372 337
rect 3366 332 3372 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 3462 331 3468 332
rect 470 325 476 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 470 321 471 325
rect 475 321 476 325
rect 470 320 476 321
rect 558 325 564 326
rect 558 321 559 325
rect 563 321 564 325
rect 558 320 564 321
rect 646 325 652 326
rect 646 321 647 325
rect 651 321 652 325
rect 646 320 652 321
rect 734 325 740 326
rect 734 321 735 325
rect 739 321 740 325
rect 734 320 740 321
rect 822 325 828 326
rect 822 321 823 325
rect 827 321 828 325
rect 822 320 828 321
rect 910 325 916 326
rect 910 321 911 325
rect 915 321 916 325
rect 910 320 916 321
rect 998 325 1004 326
rect 998 321 999 325
rect 1003 321 1004 325
rect 998 320 1004 321
rect 1086 325 1092 326
rect 1086 321 1087 325
rect 1091 321 1092 325
rect 1086 320 1092 321
rect 1174 325 1180 326
rect 1174 321 1175 325
rect 1179 321 1180 325
rect 1174 320 1180 321
rect 1262 325 1268 326
rect 1262 321 1263 325
rect 1267 321 1268 325
rect 1262 320 1268 321
rect 1766 324 1772 325
rect 1766 320 1767 324
rect 1771 320 1772 324
rect 110 319 116 320
rect 1766 319 1772 320
rect 1806 288 1812 289
rect 3462 288 3468 289
rect 1806 284 1807 288
rect 1811 284 1812 288
rect 1806 283 1812 284
rect 1926 287 1932 288
rect 1926 283 1927 287
rect 1931 283 1932 287
rect 1926 282 1932 283
rect 2038 287 2044 288
rect 2038 283 2039 287
rect 2043 283 2044 287
rect 2038 282 2044 283
rect 2166 287 2172 288
rect 2166 283 2167 287
rect 2171 283 2172 287
rect 2166 282 2172 283
rect 2302 287 2308 288
rect 2302 283 2303 287
rect 2307 283 2308 287
rect 2302 282 2308 283
rect 2446 287 2452 288
rect 2446 283 2447 287
rect 2451 283 2452 287
rect 2446 282 2452 283
rect 2598 287 2604 288
rect 2598 283 2599 287
rect 2603 283 2604 287
rect 2598 282 2604 283
rect 2758 287 2764 288
rect 2758 283 2759 287
rect 2763 283 2764 287
rect 2758 282 2764 283
rect 2918 287 2924 288
rect 2918 283 2919 287
rect 2923 283 2924 287
rect 2918 282 2924 283
rect 3086 287 3092 288
rect 3086 283 3087 287
rect 3091 283 3092 287
rect 3086 282 3092 283
rect 3254 287 3260 288
rect 3254 283 3255 287
rect 3259 283 3260 287
rect 3462 284 3463 288
rect 3467 284 3468 288
rect 3462 283 3468 284
rect 3254 282 3260 283
rect 110 276 116 277
rect 1766 276 1772 277
rect 110 272 111 276
rect 115 272 116 276
rect 110 271 116 272
rect 278 275 284 276
rect 278 271 279 275
rect 283 271 284 275
rect 278 270 284 271
rect 366 275 372 276
rect 366 271 367 275
rect 371 271 372 275
rect 366 270 372 271
rect 462 275 468 276
rect 462 271 463 275
rect 467 271 468 275
rect 462 270 468 271
rect 558 275 564 276
rect 558 271 559 275
rect 563 271 564 275
rect 558 270 564 271
rect 654 275 660 276
rect 654 271 655 275
rect 659 271 660 275
rect 654 270 660 271
rect 750 275 756 276
rect 750 271 751 275
rect 755 271 756 275
rect 750 270 756 271
rect 846 275 852 276
rect 846 271 847 275
rect 851 271 852 275
rect 846 270 852 271
rect 942 275 948 276
rect 942 271 943 275
rect 947 271 948 275
rect 942 270 948 271
rect 1046 275 1052 276
rect 1046 271 1047 275
rect 1051 271 1052 275
rect 1046 270 1052 271
rect 1150 275 1156 276
rect 1150 271 1151 275
rect 1155 271 1156 275
rect 1766 272 1767 276
rect 1771 272 1772 276
rect 1766 271 1772 272
rect 1806 271 1812 272
rect 1150 270 1156 271
rect 1806 267 1807 271
rect 1811 267 1812 271
rect 3462 271 3468 272
rect 1806 266 1812 267
rect 1926 268 1932 269
rect 1926 264 1927 268
rect 1931 264 1932 268
rect 1926 263 1932 264
rect 2038 268 2044 269
rect 2038 264 2039 268
rect 2043 264 2044 268
rect 2038 263 2044 264
rect 2166 268 2172 269
rect 2166 264 2167 268
rect 2171 264 2172 268
rect 2166 263 2172 264
rect 2302 268 2308 269
rect 2302 264 2303 268
rect 2307 264 2308 268
rect 2302 263 2308 264
rect 2446 268 2452 269
rect 2446 264 2447 268
rect 2451 264 2452 268
rect 2446 263 2452 264
rect 2598 268 2604 269
rect 2598 264 2599 268
rect 2603 264 2604 268
rect 2598 263 2604 264
rect 2758 268 2764 269
rect 2758 264 2759 268
rect 2763 264 2764 268
rect 2758 263 2764 264
rect 2918 268 2924 269
rect 2918 264 2919 268
rect 2923 264 2924 268
rect 2918 263 2924 264
rect 3086 268 3092 269
rect 3086 264 3087 268
rect 3091 264 3092 268
rect 3086 263 3092 264
rect 3254 268 3260 269
rect 3254 264 3255 268
rect 3259 264 3260 268
rect 3462 267 3463 271
rect 3467 267 3468 271
rect 3462 266 3468 267
rect 3254 263 3260 264
rect 110 259 116 260
rect 110 255 111 259
rect 115 255 116 259
rect 1766 259 1772 260
rect 110 254 116 255
rect 278 256 284 257
rect 278 252 279 256
rect 283 252 284 256
rect 278 251 284 252
rect 366 256 372 257
rect 366 252 367 256
rect 371 252 372 256
rect 366 251 372 252
rect 462 256 468 257
rect 462 252 463 256
rect 467 252 468 256
rect 462 251 468 252
rect 558 256 564 257
rect 558 252 559 256
rect 563 252 564 256
rect 558 251 564 252
rect 654 256 660 257
rect 654 252 655 256
rect 659 252 660 256
rect 654 251 660 252
rect 750 256 756 257
rect 750 252 751 256
rect 755 252 756 256
rect 750 251 756 252
rect 846 256 852 257
rect 846 252 847 256
rect 851 252 852 256
rect 846 251 852 252
rect 942 256 948 257
rect 942 252 943 256
rect 947 252 948 256
rect 942 251 948 252
rect 1046 256 1052 257
rect 1046 252 1047 256
rect 1051 252 1052 256
rect 1046 251 1052 252
rect 1150 256 1156 257
rect 1150 252 1151 256
rect 1155 252 1156 256
rect 1766 255 1767 259
rect 1771 255 1772 259
rect 1766 254 1772 255
rect 1150 251 1156 252
rect 1830 220 1836 221
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 1830 216 1831 220
rect 1835 216 1836 220
rect 1830 215 1836 216
rect 1926 220 1932 221
rect 1926 216 1927 220
rect 1931 216 1932 220
rect 1926 215 1932 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2350 220 2356 221
rect 2350 216 2351 220
rect 2355 216 2356 220
rect 2350 215 2356 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2678 220 2684 221
rect 2678 216 2679 220
rect 2683 216 2684 220
rect 2678 215 2684 216
rect 2846 220 2852 221
rect 2846 216 2847 220
rect 2851 216 2852 220
rect 2846 215 2852 216
rect 3022 220 3028 221
rect 3022 216 3023 220
rect 3027 216 3028 220
rect 3022 215 3028 216
rect 3206 220 3212 221
rect 3206 216 3207 220
rect 3211 216 3212 220
rect 3206 215 3212 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 166 208 172 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 166 204 167 208
rect 171 204 172 208
rect 166 203 172 204
rect 342 208 348 209
rect 342 204 343 208
rect 347 204 348 208
rect 342 203 348 204
rect 510 208 516 209
rect 510 204 511 208
rect 515 204 516 208
rect 510 203 516 204
rect 678 208 684 209
rect 678 204 679 208
rect 683 204 684 208
rect 678 203 684 204
rect 838 208 844 209
rect 838 204 839 208
rect 843 204 844 208
rect 838 203 844 204
rect 990 208 996 209
rect 990 204 991 208
rect 995 204 996 208
rect 990 203 996 204
rect 1134 208 1140 209
rect 1134 204 1135 208
rect 1139 204 1140 208
rect 1134 203 1140 204
rect 1278 208 1284 209
rect 1278 204 1279 208
rect 1283 204 1284 208
rect 1278 203 1284 204
rect 1430 208 1436 209
rect 1430 204 1431 208
rect 1435 204 1436 208
rect 1430 203 1436 204
rect 1766 205 1772 206
rect 110 200 116 201
rect 1766 201 1767 205
rect 1771 201 1772 205
rect 1830 201 1836 202
rect 1766 200 1772 201
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1830 197 1831 201
rect 1835 197 1836 201
rect 1830 196 1836 197
rect 1926 201 1932 202
rect 1926 197 1927 201
rect 1931 197 1932 201
rect 1926 196 1932 197
rect 2054 201 2060 202
rect 2054 197 2055 201
rect 2059 197 2060 201
rect 2054 196 2060 197
rect 2198 201 2204 202
rect 2198 197 2199 201
rect 2203 197 2204 201
rect 2198 196 2204 197
rect 2350 201 2356 202
rect 2350 197 2351 201
rect 2355 197 2356 201
rect 2350 196 2356 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2678 201 2684 202
rect 2678 197 2679 201
rect 2683 197 2684 201
rect 2678 196 2684 197
rect 2846 201 2852 202
rect 2846 197 2847 201
rect 2851 197 2852 201
rect 2846 196 2852 197
rect 3022 201 3028 202
rect 3022 197 3023 201
rect 3027 197 3028 201
rect 3022 196 3028 197
rect 3206 201 3212 202
rect 3206 197 3207 201
rect 3211 197 3212 201
rect 3206 196 3212 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1806 195 1812 196
rect 3462 195 3468 196
rect 166 189 172 190
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 166 185 167 189
rect 171 185 172 189
rect 166 184 172 185
rect 342 189 348 190
rect 342 185 343 189
rect 347 185 348 189
rect 342 184 348 185
rect 510 189 516 190
rect 510 185 511 189
rect 515 185 516 189
rect 510 184 516 185
rect 678 189 684 190
rect 678 185 679 189
rect 683 185 684 189
rect 678 184 684 185
rect 838 189 844 190
rect 838 185 839 189
rect 843 185 844 189
rect 838 184 844 185
rect 990 189 996 190
rect 990 185 991 189
rect 995 185 996 189
rect 990 184 996 185
rect 1134 189 1140 190
rect 1134 185 1135 189
rect 1139 185 1140 189
rect 1134 184 1140 185
rect 1278 189 1284 190
rect 1278 185 1279 189
rect 1283 185 1284 189
rect 1278 184 1284 185
rect 1430 189 1436 190
rect 1430 185 1431 189
rect 1435 185 1436 189
rect 1430 184 1436 185
rect 1766 188 1772 189
rect 1766 184 1767 188
rect 1771 184 1772 188
rect 110 183 116 184
rect 1766 183 1772 184
rect 1806 136 1812 137
rect 3462 136 3468 137
rect 1806 132 1807 136
rect 1811 132 1812 136
rect 1806 131 1812 132
rect 1830 135 1836 136
rect 1830 131 1831 135
rect 1835 131 1836 135
rect 1830 130 1836 131
rect 1918 135 1924 136
rect 1918 131 1919 135
rect 1923 131 1924 135
rect 1918 130 1924 131
rect 2038 135 2044 136
rect 2038 131 2039 135
rect 2043 131 2044 135
rect 2038 130 2044 131
rect 2158 135 2164 136
rect 2158 131 2159 135
rect 2163 131 2164 135
rect 2158 130 2164 131
rect 2278 135 2284 136
rect 2278 131 2279 135
rect 2283 131 2284 135
rect 2278 130 2284 131
rect 2398 135 2404 136
rect 2398 131 2399 135
rect 2403 131 2404 135
rect 2398 130 2404 131
rect 2510 135 2516 136
rect 2510 131 2511 135
rect 2515 131 2516 135
rect 2510 130 2516 131
rect 2622 135 2628 136
rect 2622 131 2623 135
rect 2627 131 2628 135
rect 2622 130 2628 131
rect 2734 135 2740 136
rect 2734 131 2735 135
rect 2739 131 2740 135
rect 2734 130 2740 131
rect 2838 135 2844 136
rect 2838 131 2839 135
rect 2843 131 2844 135
rect 2838 130 2844 131
rect 2942 135 2948 136
rect 2942 131 2943 135
rect 2947 131 2948 135
rect 2942 130 2948 131
rect 3054 135 3060 136
rect 3054 131 3055 135
rect 3059 131 3060 135
rect 3054 130 3060 131
rect 3166 135 3172 136
rect 3166 131 3167 135
rect 3171 131 3172 135
rect 3166 130 3172 131
rect 3278 135 3284 136
rect 3278 131 3279 135
rect 3283 131 3284 135
rect 3278 130 3284 131
rect 3366 135 3372 136
rect 3366 131 3367 135
rect 3371 131 3372 135
rect 3462 132 3463 136
rect 3467 132 3468 136
rect 3462 131 3468 132
rect 3366 130 3372 131
rect 110 120 116 121
rect 1766 120 1772 121
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 134 119 140 120
rect 134 115 135 119
rect 139 115 140 119
rect 134 114 140 115
rect 222 119 228 120
rect 222 115 223 119
rect 227 115 228 119
rect 222 114 228 115
rect 310 119 316 120
rect 310 115 311 119
rect 315 115 316 119
rect 310 114 316 115
rect 398 119 404 120
rect 398 115 399 119
rect 403 115 404 119
rect 398 114 404 115
rect 486 119 492 120
rect 486 115 487 119
rect 491 115 492 119
rect 486 114 492 115
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 662 119 668 120
rect 662 115 663 119
rect 667 115 668 119
rect 662 114 668 115
rect 750 119 756 120
rect 750 115 751 119
rect 755 115 756 119
rect 750 114 756 115
rect 846 119 852 120
rect 846 115 847 119
rect 851 115 852 119
rect 846 114 852 115
rect 942 119 948 120
rect 942 115 943 119
rect 947 115 948 119
rect 942 114 948 115
rect 1030 119 1036 120
rect 1030 115 1031 119
rect 1035 115 1036 119
rect 1030 114 1036 115
rect 1118 119 1124 120
rect 1118 115 1119 119
rect 1123 115 1124 119
rect 1118 114 1124 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1310 119 1316 120
rect 1310 115 1311 119
rect 1315 115 1316 119
rect 1310 114 1316 115
rect 1406 119 1412 120
rect 1406 115 1407 119
rect 1411 115 1412 119
rect 1406 114 1412 115
rect 1494 119 1500 120
rect 1494 115 1495 119
rect 1499 115 1500 119
rect 1494 114 1500 115
rect 1582 119 1588 120
rect 1582 115 1583 119
rect 1587 115 1588 119
rect 1582 114 1588 115
rect 1670 119 1676 120
rect 1670 115 1671 119
rect 1675 115 1676 119
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 119 1812 120
rect 1806 115 1807 119
rect 1811 115 1812 119
rect 3462 119 3468 120
rect 1670 114 1676 115
rect 1806 114 1812 115
rect 1830 116 1836 117
rect 1830 112 1831 116
rect 1835 112 1836 116
rect 1830 111 1836 112
rect 1918 116 1924 117
rect 1918 112 1919 116
rect 1923 112 1924 116
rect 1918 111 1924 112
rect 2038 116 2044 117
rect 2038 112 2039 116
rect 2043 112 2044 116
rect 2038 111 2044 112
rect 2158 116 2164 117
rect 2158 112 2159 116
rect 2163 112 2164 116
rect 2158 111 2164 112
rect 2278 116 2284 117
rect 2278 112 2279 116
rect 2283 112 2284 116
rect 2278 111 2284 112
rect 2398 116 2404 117
rect 2398 112 2399 116
rect 2403 112 2404 116
rect 2398 111 2404 112
rect 2510 116 2516 117
rect 2510 112 2511 116
rect 2515 112 2516 116
rect 2510 111 2516 112
rect 2622 116 2628 117
rect 2622 112 2623 116
rect 2627 112 2628 116
rect 2622 111 2628 112
rect 2734 116 2740 117
rect 2734 112 2735 116
rect 2739 112 2740 116
rect 2734 111 2740 112
rect 2838 116 2844 117
rect 2838 112 2839 116
rect 2843 112 2844 116
rect 2838 111 2844 112
rect 2942 116 2948 117
rect 2942 112 2943 116
rect 2947 112 2948 116
rect 2942 111 2948 112
rect 3054 116 3060 117
rect 3054 112 3055 116
rect 3059 112 3060 116
rect 3054 111 3060 112
rect 3166 116 3172 117
rect 3166 112 3167 116
rect 3171 112 3172 116
rect 3166 111 3172 112
rect 3278 116 3284 117
rect 3278 112 3279 116
rect 3283 112 3284 116
rect 3278 111 3284 112
rect 3366 116 3372 117
rect 3366 112 3367 116
rect 3371 112 3372 116
rect 3462 115 3463 119
rect 3467 115 3468 119
rect 3462 114 3468 115
rect 3366 111 3372 112
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 1766 103 1772 104
rect 110 98 116 99
rect 134 100 140 101
rect 134 96 135 100
rect 139 96 140 100
rect 134 95 140 96
rect 222 100 228 101
rect 222 96 223 100
rect 227 96 228 100
rect 222 95 228 96
rect 310 100 316 101
rect 310 96 311 100
rect 315 96 316 100
rect 310 95 316 96
rect 398 100 404 101
rect 398 96 399 100
rect 403 96 404 100
rect 398 95 404 96
rect 486 100 492 101
rect 486 96 487 100
rect 491 96 492 100
rect 486 95 492 96
rect 574 100 580 101
rect 574 96 575 100
rect 579 96 580 100
rect 574 95 580 96
rect 662 100 668 101
rect 662 96 663 100
rect 667 96 668 100
rect 662 95 668 96
rect 750 100 756 101
rect 750 96 751 100
rect 755 96 756 100
rect 750 95 756 96
rect 846 100 852 101
rect 846 96 847 100
rect 851 96 852 100
rect 846 95 852 96
rect 942 100 948 101
rect 942 96 943 100
rect 947 96 948 100
rect 942 95 948 96
rect 1030 100 1036 101
rect 1030 96 1031 100
rect 1035 96 1036 100
rect 1030 95 1036 96
rect 1118 100 1124 101
rect 1118 96 1119 100
rect 1123 96 1124 100
rect 1118 95 1124 96
rect 1214 100 1220 101
rect 1214 96 1215 100
rect 1219 96 1220 100
rect 1214 95 1220 96
rect 1310 100 1316 101
rect 1310 96 1311 100
rect 1315 96 1316 100
rect 1310 95 1316 96
rect 1406 100 1412 101
rect 1406 96 1407 100
rect 1411 96 1412 100
rect 1406 95 1412 96
rect 1494 100 1500 101
rect 1494 96 1495 100
rect 1499 96 1500 100
rect 1494 95 1500 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1670 100 1676 101
rect 1670 96 1671 100
rect 1675 96 1676 100
rect 1766 99 1767 103
rect 1771 99 1772 103
rect 1766 98 1772 99
rect 1670 95 1676 96
<< m3c >>
rect 1807 3496 1811 3500
rect 2007 3495 2011 3499
rect 2239 3495 2243 3499
rect 2455 3495 2459 3499
rect 2655 3495 2659 3499
rect 2855 3495 2859 3499
rect 3047 3495 3051 3499
rect 3247 3495 3251 3499
rect 3463 3496 3467 3500
rect 1807 3479 1811 3483
rect 2007 3476 2011 3480
rect 2239 3476 2243 3480
rect 2455 3476 2459 3480
rect 2655 3476 2659 3480
rect 2855 3476 2859 3480
rect 3047 3476 3051 3480
rect 3247 3476 3251 3480
rect 3463 3479 3467 3483
rect 111 3460 115 3464
rect 455 3459 459 3463
rect 543 3459 547 3463
rect 631 3459 635 3463
rect 719 3459 723 3463
rect 807 3459 811 3463
rect 895 3459 899 3463
rect 983 3459 987 3463
rect 1071 3459 1075 3463
rect 1159 3459 1163 3463
rect 1767 3460 1771 3464
rect 111 3443 115 3447
rect 455 3440 459 3444
rect 543 3440 547 3444
rect 631 3440 635 3444
rect 719 3440 723 3444
rect 807 3440 811 3444
rect 895 3440 899 3444
rect 983 3440 987 3444
rect 1071 3440 1075 3444
rect 1159 3440 1163 3444
rect 1767 3443 1771 3447
rect 1807 3429 1811 3433
rect 1831 3432 1835 3436
rect 1943 3432 1947 3436
rect 2079 3432 2083 3436
rect 2215 3432 2219 3436
rect 2351 3432 2355 3436
rect 2479 3432 2483 3436
rect 2599 3432 2603 3436
rect 2719 3432 2723 3436
rect 2847 3432 2851 3436
rect 2975 3432 2979 3436
rect 3463 3429 3467 3433
rect 1807 3412 1811 3416
rect 1831 3413 1835 3417
rect 1943 3413 1947 3417
rect 2079 3413 2083 3417
rect 2215 3413 2219 3417
rect 2351 3413 2355 3417
rect 2479 3413 2483 3417
rect 2599 3413 2603 3417
rect 2719 3413 2723 3417
rect 2847 3413 2851 3417
rect 2975 3413 2979 3417
rect 3463 3412 3467 3416
rect 111 3393 115 3397
rect 415 3396 419 3400
rect 503 3396 507 3400
rect 591 3396 595 3400
rect 679 3396 683 3400
rect 767 3396 771 3400
rect 855 3396 859 3400
rect 943 3396 947 3400
rect 1031 3396 1035 3400
rect 1119 3396 1123 3400
rect 1207 3396 1211 3400
rect 1303 3396 1307 3400
rect 1767 3393 1771 3397
rect 111 3376 115 3380
rect 415 3377 419 3381
rect 503 3377 507 3381
rect 591 3377 595 3381
rect 679 3377 683 3381
rect 767 3377 771 3381
rect 855 3377 859 3381
rect 943 3377 947 3381
rect 1031 3377 1035 3381
rect 1119 3377 1123 3381
rect 1207 3377 1211 3381
rect 1303 3377 1307 3381
rect 1767 3376 1771 3380
rect 1807 3360 1811 3364
rect 1831 3359 1835 3363
rect 1951 3359 1955 3363
rect 2095 3359 2099 3363
rect 2239 3359 2243 3363
rect 2383 3359 2387 3363
rect 2519 3359 2523 3363
rect 2647 3359 2651 3363
rect 2775 3359 2779 3363
rect 2903 3359 2907 3363
rect 3039 3359 3043 3363
rect 3463 3360 3467 3364
rect 1807 3343 1811 3347
rect 1831 3340 1835 3344
rect 1951 3340 1955 3344
rect 2095 3340 2099 3344
rect 2239 3340 2243 3344
rect 2383 3340 2387 3344
rect 2519 3340 2523 3344
rect 2647 3340 2651 3344
rect 2775 3340 2779 3344
rect 2903 3340 2907 3344
rect 3039 3340 3043 3344
rect 3463 3343 3467 3347
rect 111 3328 115 3332
rect 399 3327 403 3331
rect 495 3327 499 3331
rect 599 3327 603 3331
rect 703 3327 707 3331
rect 807 3327 811 3331
rect 911 3327 915 3331
rect 1015 3327 1019 3331
rect 1119 3327 1123 3331
rect 1223 3327 1227 3331
rect 1327 3327 1331 3331
rect 1767 3328 1771 3332
rect 111 3311 115 3315
rect 399 3308 403 3312
rect 495 3308 499 3312
rect 599 3308 603 3312
rect 703 3308 707 3312
rect 807 3308 811 3312
rect 911 3308 915 3312
rect 1015 3308 1019 3312
rect 1119 3308 1123 3312
rect 1223 3308 1227 3312
rect 1327 3308 1331 3312
rect 1767 3311 1771 3315
rect 1807 3285 1811 3289
rect 1831 3288 1835 3292
rect 1975 3288 1979 3292
rect 2151 3288 2155 3292
rect 2335 3288 2339 3292
rect 2511 3288 2515 3292
rect 2679 3288 2683 3292
rect 2831 3288 2835 3292
rect 2975 3288 2979 3292
rect 3111 3288 3115 3292
rect 3247 3288 3251 3292
rect 3367 3288 3371 3292
rect 3463 3285 3467 3289
rect 1807 3268 1811 3272
rect 1831 3269 1835 3273
rect 1975 3269 1979 3273
rect 2151 3269 2155 3273
rect 2335 3269 2339 3273
rect 2511 3269 2515 3273
rect 2679 3269 2683 3273
rect 2831 3269 2835 3273
rect 2975 3269 2979 3273
rect 3111 3269 3115 3273
rect 3247 3269 3251 3273
rect 3367 3269 3371 3273
rect 3463 3268 3467 3272
rect 111 3257 115 3261
rect 383 3260 387 3264
rect 495 3260 499 3264
rect 607 3260 611 3264
rect 727 3260 731 3264
rect 847 3260 851 3264
rect 967 3260 971 3264
rect 1087 3260 1091 3264
rect 1207 3260 1211 3264
rect 1335 3260 1339 3264
rect 1767 3257 1771 3261
rect 111 3240 115 3244
rect 383 3241 387 3245
rect 495 3241 499 3245
rect 607 3241 611 3245
rect 727 3241 731 3245
rect 847 3241 851 3245
rect 967 3241 971 3245
rect 1087 3241 1091 3245
rect 1207 3241 1211 3245
rect 1335 3241 1339 3245
rect 1767 3240 1771 3244
rect 1807 3216 1811 3220
rect 1831 3215 1835 3219
rect 2031 3215 2035 3219
rect 2247 3215 2251 3219
rect 2455 3215 2459 3219
rect 2655 3215 2659 3219
rect 2839 3215 2843 3219
rect 3023 3215 3027 3219
rect 3207 3215 3211 3219
rect 3367 3215 3371 3219
rect 3463 3216 3467 3220
rect 1807 3199 1811 3203
rect 111 3192 115 3196
rect 303 3191 307 3195
rect 423 3191 427 3195
rect 543 3191 547 3195
rect 671 3191 675 3195
rect 799 3191 803 3195
rect 927 3191 931 3195
rect 1055 3191 1059 3195
rect 1175 3191 1179 3195
rect 1303 3191 1307 3195
rect 1431 3191 1435 3195
rect 1767 3192 1771 3196
rect 1831 3196 1835 3200
rect 2031 3196 2035 3200
rect 2247 3196 2251 3200
rect 2455 3196 2459 3200
rect 2655 3196 2659 3200
rect 2839 3196 2843 3200
rect 3023 3196 3027 3200
rect 3207 3196 3211 3200
rect 3367 3196 3371 3200
rect 3463 3199 3467 3203
rect 111 3175 115 3179
rect 303 3172 307 3176
rect 423 3172 427 3176
rect 543 3172 547 3176
rect 671 3172 675 3176
rect 799 3172 803 3176
rect 927 3172 931 3176
rect 1055 3172 1059 3176
rect 1175 3172 1179 3176
rect 1303 3172 1307 3176
rect 1431 3172 1435 3176
rect 1767 3175 1771 3179
rect 1807 3149 1811 3153
rect 1839 3152 1843 3156
rect 2031 3152 2035 3156
rect 2223 3152 2227 3156
rect 2407 3152 2411 3156
rect 2575 3152 2579 3156
rect 2735 3152 2739 3156
rect 2879 3152 2883 3156
rect 3007 3152 3011 3156
rect 3135 3152 3139 3156
rect 3263 3152 3267 3156
rect 3367 3152 3371 3156
rect 3463 3149 3467 3153
rect 1807 3132 1811 3136
rect 1839 3133 1843 3137
rect 2031 3133 2035 3137
rect 2223 3133 2227 3137
rect 2407 3133 2411 3137
rect 2575 3133 2579 3137
rect 2735 3133 2739 3137
rect 2879 3133 2883 3137
rect 3007 3133 3011 3137
rect 3135 3133 3139 3137
rect 3263 3133 3267 3137
rect 3367 3133 3371 3137
rect 3463 3132 3467 3136
rect 111 3113 115 3117
rect 175 3116 179 3120
rect 319 3116 323 3120
rect 471 3116 475 3120
rect 623 3116 627 3120
rect 775 3116 779 3120
rect 919 3116 923 3120
rect 1063 3116 1067 3120
rect 1199 3116 1203 3120
rect 1343 3116 1347 3120
rect 1487 3116 1491 3120
rect 1767 3113 1771 3117
rect 111 3096 115 3100
rect 175 3097 179 3101
rect 319 3097 323 3101
rect 471 3097 475 3101
rect 623 3097 627 3101
rect 775 3097 779 3101
rect 919 3097 923 3101
rect 1063 3097 1067 3101
rect 1199 3097 1203 3101
rect 1343 3097 1347 3101
rect 1487 3097 1491 3101
rect 1767 3096 1771 3100
rect 1807 3084 1811 3088
rect 1935 3083 1939 3087
rect 2055 3083 2059 3087
rect 2175 3083 2179 3087
rect 2303 3083 2307 3087
rect 2431 3083 2435 3087
rect 2567 3083 2571 3087
rect 2719 3083 2723 3087
rect 2871 3083 2875 3087
rect 3031 3083 3035 3087
rect 3199 3083 3203 3087
rect 3367 3083 3371 3087
rect 3463 3084 3467 3088
rect 1807 3067 1811 3071
rect 1935 3064 1939 3068
rect 2055 3064 2059 3068
rect 2175 3064 2179 3068
rect 2303 3064 2307 3068
rect 2431 3064 2435 3068
rect 2567 3064 2571 3068
rect 2719 3064 2723 3068
rect 2871 3064 2875 3068
rect 3031 3064 3035 3068
rect 3199 3064 3203 3068
rect 3367 3064 3371 3068
rect 3463 3067 3467 3071
rect 111 3044 115 3048
rect 135 3043 139 3047
rect 263 3043 267 3047
rect 431 3043 435 3047
rect 607 3043 611 3047
rect 791 3043 795 3047
rect 967 3043 971 3047
rect 1143 3043 1147 3047
rect 1327 3043 1331 3047
rect 1511 3043 1515 3047
rect 1767 3044 1771 3048
rect 111 3027 115 3031
rect 135 3024 139 3028
rect 263 3024 267 3028
rect 431 3024 435 3028
rect 607 3024 611 3028
rect 791 3024 795 3028
rect 967 3024 971 3028
rect 1143 3024 1147 3028
rect 1327 3024 1331 3028
rect 1511 3024 1515 3028
rect 1767 3027 1771 3031
rect 1807 3009 1811 3013
rect 2023 3012 2027 3016
rect 2127 3012 2131 3016
rect 2231 3012 2235 3016
rect 2335 3012 2339 3016
rect 2439 3012 2443 3016
rect 2543 3012 2547 3016
rect 2647 3012 2651 3016
rect 2759 3012 2763 3016
rect 3463 3009 3467 3013
rect 1807 2992 1811 2996
rect 2023 2993 2027 2997
rect 2127 2993 2131 2997
rect 2231 2993 2235 2997
rect 2335 2993 2339 2997
rect 2439 2993 2443 2997
rect 2543 2993 2547 2997
rect 2647 2993 2651 2997
rect 2759 2993 2763 2997
rect 3463 2992 3467 2996
rect 111 2973 115 2977
rect 135 2976 139 2980
rect 327 2976 331 2980
rect 535 2976 539 2980
rect 735 2976 739 2980
rect 927 2976 931 2980
rect 1103 2976 1107 2980
rect 1279 2976 1283 2980
rect 1447 2976 1451 2980
rect 1623 2976 1627 2980
rect 1767 2973 1771 2977
rect 111 2956 115 2960
rect 135 2957 139 2961
rect 327 2957 331 2961
rect 535 2957 539 2961
rect 735 2957 739 2961
rect 927 2957 931 2961
rect 1103 2957 1107 2961
rect 1279 2957 1283 2961
rect 1447 2957 1451 2961
rect 1623 2957 1627 2961
rect 1767 2956 1771 2960
rect 1807 2948 1811 2952
rect 2055 2947 2059 2951
rect 2143 2947 2147 2951
rect 2231 2947 2235 2951
rect 2319 2947 2323 2951
rect 2407 2947 2411 2951
rect 2495 2947 2499 2951
rect 2583 2947 2587 2951
rect 2671 2947 2675 2951
rect 2759 2947 2763 2951
rect 2847 2947 2851 2951
rect 3463 2948 3467 2952
rect 1807 2931 1811 2935
rect 2055 2928 2059 2932
rect 2143 2928 2147 2932
rect 2231 2928 2235 2932
rect 2319 2928 2323 2932
rect 2407 2928 2411 2932
rect 2495 2928 2499 2932
rect 2583 2928 2587 2932
rect 2671 2928 2675 2932
rect 2759 2928 2763 2932
rect 2847 2928 2851 2932
rect 3463 2931 3467 2935
rect 111 2904 115 2908
rect 135 2903 139 2907
rect 263 2903 267 2907
rect 431 2903 435 2907
rect 607 2903 611 2907
rect 783 2903 787 2907
rect 951 2903 955 2907
rect 1111 2903 1115 2907
rect 1271 2903 1275 2907
rect 1431 2903 1435 2907
rect 1591 2903 1595 2907
rect 1767 2904 1771 2908
rect 111 2887 115 2891
rect 135 2884 139 2888
rect 263 2884 267 2888
rect 431 2884 435 2888
rect 607 2884 611 2888
rect 783 2884 787 2888
rect 951 2884 955 2888
rect 1111 2884 1115 2888
rect 1271 2884 1275 2888
rect 1431 2884 1435 2888
rect 1591 2884 1595 2888
rect 1767 2887 1771 2891
rect 1807 2873 1811 2877
rect 2071 2876 2075 2880
rect 2175 2876 2179 2880
rect 2271 2876 2275 2880
rect 2367 2876 2371 2880
rect 2471 2876 2475 2880
rect 2575 2876 2579 2880
rect 2679 2876 2683 2880
rect 2783 2876 2787 2880
rect 3463 2873 3467 2877
rect 1807 2856 1811 2860
rect 2071 2857 2075 2861
rect 2175 2857 2179 2861
rect 2271 2857 2275 2861
rect 2367 2857 2371 2861
rect 2471 2857 2475 2861
rect 2575 2857 2579 2861
rect 2679 2857 2683 2861
rect 2783 2857 2787 2861
rect 3463 2856 3467 2860
rect 111 2833 115 2837
rect 135 2836 139 2840
rect 255 2836 259 2840
rect 407 2836 411 2840
rect 567 2836 571 2840
rect 727 2836 731 2840
rect 879 2836 883 2840
rect 1023 2836 1027 2840
rect 1167 2836 1171 2840
rect 1311 2836 1315 2840
rect 1463 2836 1467 2840
rect 1767 2833 1771 2837
rect 111 2816 115 2820
rect 135 2817 139 2821
rect 255 2817 259 2821
rect 407 2817 411 2821
rect 567 2817 571 2821
rect 727 2817 731 2821
rect 879 2817 883 2821
rect 1023 2817 1027 2821
rect 1167 2817 1171 2821
rect 1311 2817 1315 2821
rect 1463 2817 1467 2821
rect 1767 2816 1771 2820
rect 1807 2808 1811 2812
rect 1983 2807 1987 2811
rect 2111 2807 2115 2811
rect 2239 2807 2243 2811
rect 2367 2807 2371 2811
rect 2487 2807 2491 2811
rect 2607 2807 2611 2811
rect 2719 2807 2723 2811
rect 2839 2807 2843 2811
rect 2959 2807 2963 2811
rect 3463 2808 3467 2812
rect 1807 2791 1811 2795
rect 1983 2788 1987 2792
rect 2111 2788 2115 2792
rect 2239 2788 2243 2792
rect 2367 2788 2371 2792
rect 2487 2788 2491 2792
rect 2607 2788 2611 2792
rect 2719 2788 2723 2792
rect 2839 2788 2843 2792
rect 2959 2788 2963 2792
rect 3463 2791 3467 2795
rect 111 2764 115 2768
rect 287 2763 291 2767
rect 391 2763 395 2767
rect 503 2763 507 2767
rect 623 2763 627 2767
rect 743 2763 747 2767
rect 855 2763 859 2767
rect 967 2763 971 2767
rect 1079 2763 1083 2767
rect 1199 2763 1203 2767
rect 1319 2763 1323 2767
rect 1767 2764 1771 2768
rect 111 2747 115 2751
rect 287 2744 291 2748
rect 391 2744 395 2748
rect 503 2744 507 2748
rect 623 2744 627 2748
rect 743 2744 747 2748
rect 855 2744 859 2748
rect 967 2744 971 2748
rect 1079 2744 1083 2748
rect 1199 2744 1203 2748
rect 1319 2744 1323 2748
rect 1767 2747 1771 2751
rect 1807 2737 1811 2741
rect 1887 2740 1891 2744
rect 2031 2740 2035 2744
rect 2183 2740 2187 2744
rect 2335 2740 2339 2744
rect 2479 2740 2483 2744
rect 2623 2740 2627 2744
rect 2767 2740 2771 2744
rect 2911 2740 2915 2744
rect 3055 2740 3059 2744
rect 3463 2737 3467 2741
rect 1807 2720 1811 2724
rect 1887 2721 1891 2725
rect 2031 2721 2035 2725
rect 2183 2721 2187 2725
rect 2335 2721 2339 2725
rect 2479 2721 2483 2725
rect 2623 2721 2627 2725
rect 2767 2721 2771 2725
rect 2911 2721 2915 2725
rect 3055 2721 3059 2725
rect 3463 2720 3467 2724
rect 111 2693 115 2697
rect 479 2696 483 2700
rect 567 2696 571 2700
rect 655 2696 659 2700
rect 743 2696 747 2700
rect 831 2696 835 2700
rect 919 2696 923 2700
rect 1007 2696 1011 2700
rect 1095 2696 1099 2700
rect 1183 2696 1187 2700
rect 1767 2693 1771 2697
rect 111 2676 115 2680
rect 479 2677 483 2681
rect 567 2677 571 2681
rect 655 2677 659 2681
rect 743 2677 747 2681
rect 831 2677 835 2681
rect 919 2677 923 2681
rect 1007 2677 1011 2681
rect 1095 2677 1099 2681
rect 1183 2677 1187 2681
rect 1767 2676 1771 2680
rect 1807 2676 1811 2680
rect 1831 2675 1835 2679
rect 2023 2675 2027 2679
rect 2231 2675 2235 2679
rect 2431 2675 2435 2679
rect 2615 2675 2619 2679
rect 2783 2675 2787 2679
rect 2943 2675 2947 2679
rect 3095 2675 3099 2679
rect 3239 2675 3243 2679
rect 3367 2675 3371 2679
rect 3463 2676 3467 2680
rect 1807 2659 1811 2663
rect 1831 2656 1835 2660
rect 2023 2656 2027 2660
rect 2231 2656 2235 2660
rect 2431 2656 2435 2660
rect 2615 2656 2619 2660
rect 2783 2656 2787 2660
rect 2943 2656 2947 2660
rect 3095 2656 3099 2660
rect 3239 2656 3243 2660
rect 3367 2656 3371 2660
rect 3463 2659 3467 2663
rect 111 2624 115 2628
rect 471 2623 475 2627
rect 559 2623 563 2627
rect 647 2623 651 2627
rect 735 2623 739 2627
rect 823 2623 827 2627
rect 911 2623 915 2627
rect 999 2623 1003 2627
rect 1087 2623 1091 2627
rect 1767 2624 1771 2628
rect 111 2607 115 2611
rect 471 2604 475 2608
rect 559 2604 563 2608
rect 647 2604 651 2608
rect 735 2604 739 2608
rect 823 2604 827 2608
rect 911 2604 915 2608
rect 999 2604 1003 2608
rect 1087 2604 1091 2608
rect 1767 2607 1771 2611
rect 1807 2605 1811 2609
rect 1831 2608 1835 2612
rect 1999 2608 2003 2612
rect 2183 2608 2187 2612
rect 2359 2608 2363 2612
rect 2519 2608 2523 2612
rect 2671 2608 2675 2612
rect 2807 2608 2811 2612
rect 2927 2608 2931 2612
rect 3047 2608 3051 2612
rect 3159 2608 3163 2612
rect 3271 2608 3275 2612
rect 3367 2608 3371 2612
rect 3463 2605 3467 2609
rect 1807 2588 1811 2592
rect 1831 2589 1835 2593
rect 1999 2589 2003 2593
rect 2183 2589 2187 2593
rect 2359 2589 2363 2593
rect 2519 2589 2523 2593
rect 2671 2589 2675 2593
rect 2807 2589 2811 2593
rect 2927 2589 2931 2593
rect 3047 2589 3051 2593
rect 3159 2589 3163 2593
rect 3271 2589 3275 2593
rect 3367 2589 3371 2593
rect 3463 2588 3467 2592
rect 111 2545 115 2549
rect 223 2548 227 2552
rect 311 2548 315 2552
rect 407 2548 411 2552
rect 503 2548 507 2552
rect 591 2548 595 2552
rect 679 2548 683 2552
rect 767 2548 771 2552
rect 855 2548 859 2552
rect 943 2548 947 2552
rect 1031 2548 1035 2552
rect 1119 2548 1123 2552
rect 1215 2548 1219 2552
rect 1311 2548 1315 2552
rect 1407 2548 1411 2552
rect 1495 2548 1499 2552
rect 1583 2548 1587 2552
rect 1671 2548 1675 2552
rect 1767 2545 1771 2549
rect 1807 2536 1811 2540
rect 2207 2535 2211 2539
rect 2799 2535 2803 2539
rect 3367 2535 3371 2539
rect 3463 2536 3467 2540
rect 111 2528 115 2532
rect 223 2529 227 2533
rect 311 2529 315 2533
rect 407 2529 411 2533
rect 503 2529 507 2533
rect 591 2529 595 2533
rect 679 2529 683 2533
rect 767 2529 771 2533
rect 855 2529 859 2533
rect 943 2529 947 2533
rect 1031 2529 1035 2533
rect 1119 2529 1123 2533
rect 1215 2529 1219 2533
rect 1311 2529 1315 2533
rect 1407 2529 1411 2533
rect 1495 2529 1499 2533
rect 1583 2529 1587 2533
rect 1671 2529 1675 2533
rect 1767 2528 1771 2532
rect 1807 2519 1811 2523
rect 2207 2516 2211 2520
rect 2799 2516 2803 2520
rect 3367 2516 3371 2520
rect 3463 2519 3467 2523
rect 111 2484 115 2488
rect 135 2483 139 2487
rect 247 2483 251 2487
rect 391 2483 395 2487
rect 543 2483 547 2487
rect 695 2483 699 2487
rect 839 2483 843 2487
rect 975 2483 979 2487
rect 1103 2483 1107 2487
rect 1231 2483 1235 2487
rect 1351 2483 1355 2487
rect 1463 2483 1467 2487
rect 1575 2483 1579 2487
rect 1671 2483 1675 2487
rect 1767 2484 1771 2488
rect 111 2467 115 2471
rect 135 2464 139 2468
rect 247 2464 251 2468
rect 391 2464 395 2468
rect 543 2464 547 2468
rect 695 2464 699 2468
rect 839 2464 843 2468
rect 975 2464 979 2468
rect 1103 2464 1107 2468
rect 1231 2464 1235 2468
rect 1351 2464 1355 2468
rect 1463 2464 1467 2468
rect 1575 2464 1579 2468
rect 1671 2464 1675 2468
rect 1767 2467 1771 2471
rect 1807 2453 1811 2457
rect 2015 2456 2019 2460
rect 2199 2456 2203 2460
rect 2367 2456 2371 2460
rect 2527 2456 2531 2460
rect 2671 2456 2675 2460
rect 2807 2456 2811 2460
rect 2927 2456 2931 2460
rect 3047 2456 3051 2460
rect 3159 2456 3163 2460
rect 3271 2456 3275 2460
rect 3367 2456 3371 2460
rect 3463 2453 3467 2457
rect 1807 2436 1811 2440
rect 2015 2437 2019 2441
rect 2199 2437 2203 2441
rect 2367 2437 2371 2441
rect 2527 2437 2531 2441
rect 2671 2437 2675 2441
rect 2807 2437 2811 2441
rect 2927 2437 2931 2441
rect 3047 2437 3051 2441
rect 3159 2437 3163 2441
rect 3271 2437 3275 2441
rect 3367 2437 3371 2441
rect 3463 2436 3467 2440
rect 111 2401 115 2405
rect 135 2404 139 2408
rect 239 2404 243 2408
rect 391 2404 395 2408
rect 551 2404 555 2408
rect 719 2404 723 2408
rect 895 2404 899 2408
rect 1063 2404 1067 2408
rect 1239 2404 1243 2408
rect 1415 2404 1419 2408
rect 1591 2404 1595 2408
rect 1767 2401 1771 2405
rect 111 2384 115 2388
rect 135 2385 139 2389
rect 239 2385 243 2389
rect 391 2385 395 2389
rect 551 2385 555 2389
rect 719 2385 723 2389
rect 895 2385 899 2389
rect 1063 2385 1067 2389
rect 1239 2385 1243 2389
rect 1415 2385 1419 2389
rect 1591 2385 1595 2389
rect 1767 2384 1771 2388
rect 1807 2388 1811 2392
rect 1839 2387 1843 2391
rect 2007 2387 2011 2391
rect 2183 2387 2187 2391
rect 2367 2387 2371 2391
rect 2559 2387 2563 2391
rect 2759 2387 2763 2391
rect 2967 2387 2971 2391
rect 3175 2387 3179 2391
rect 3367 2387 3371 2391
rect 3463 2388 3467 2392
rect 1807 2371 1811 2375
rect 1839 2368 1843 2372
rect 2007 2368 2011 2372
rect 2183 2368 2187 2372
rect 2367 2368 2371 2372
rect 2559 2368 2563 2372
rect 2759 2368 2763 2372
rect 2967 2368 2971 2372
rect 3175 2368 3179 2372
rect 3367 2368 3371 2372
rect 3463 2371 3467 2375
rect 111 2332 115 2336
rect 375 2331 379 2335
rect 479 2331 483 2335
rect 599 2331 603 2335
rect 719 2331 723 2335
rect 847 2331 851 2335
rect 975 2331 979 2335
rect 1103 2331 1107 2335
rect 1239 2331 1243 2335
rect 1375 2331 1379 2335
rect 1511 2331 1515 2335
rect 1767 2332 1771 2336
rect 1807 2321 1811 2325
rect 1887 2324 1891 2328
rect 2015 2324 2019 2328
rect 2151 2324 2155 2328
rect 2303 2324 2307 2328
rect 2463 2324 2467 2328
rect 2647 2324 2651 2328
rect 2839 2324 2843 2328
rect 3047 2324 3051 2328
rect 3255 2324 3259 2328
rect 3463 2321 3467 2325
rect 111 2315 115 2319
rect 375 2312 379 2316
rect 479 2312 483 2316
rect 599 2312 603 2316
rect 719 2312 723 2316
rect 847 2312 851 2316
rect 975 2312 979 2316
rect 1103 2312 1107 2316
rect 1239 2312 1243 2316
rect 1375 2312 1379 2316
rect 1511 2312 1515 2316
rect 1767 2315 1771 2319
rect 1807 2304 1811 2308
rect 1887 2305 1891 2309
rect 2015 2305 2019 2309
rect 2151 2305 2155 2309
rect 2303 2305 2307 2309
rect 2463 2305 2467 2309
rect 2647 2305 2651 2309
rect 2839 2305 2843 2309
rect 3047 2305 3051 2309
rect 3255 2305 3259 2309
rect 3463 2304 3467 2308
rect 111 2257 115 2261
rect 575 2260 579 2264
rect 663 2260 667 2264
rect 759 2260 763 2264
rect 863 2260 867 2264
rect 967 2260 971 2264
rect 1079 2260 1083 2264
rect 1191 2260 1195 2264
rect 1303 2260 1307 2264
rect 1415 2260 1419 2264
rect 1767 2257 1771 2261
rect 1807 2256 1811 2260
rect 2039 2255 2043 2259
rect 2135 2255 2139 2259
rect 2239 2255 2243 2259
rect 2343 2255 2347 2259
rect 2463 2255 2467 2259
rect 2591 2255 2595 2259
rect 2735 2255 2739 2259
rect 2887 2255 2891 2259
rect 3047 2255 3051 2259
rect 3215 2255 3219 2259
rect 3367 2255 3371 2259
rect 3463 2256 3467 2260
rect 111 2240 115 2244
rect 575 2241 579 2245
rect 663 2241 667 2245
rect 759 2241 763 2245
rect 863 2241 867 2245
rect 967 2241 971 2245
rect 1079 2241 1083 2245
rect 1191 2241 1195 2245
rect 1303 2241 1307 2245
rect 1415 2241 1419 2245
rect 1767 2240 1771 2244
rect 1807 2239 1811 2243
rect 2039 2236 2043 2240
rect 2135 2236 2139 2240
rect 2239 2236 2243 2240
rect 2343 2236 2347 2240
rect 2463 2236 2467 2240
rect 2591 2236 2595 2240
rect 2735 2236 2739 2240
rect 2887 2236 2891 2240
rect 3047 2236 3051 2240
rect 3215 2236 3219 2240
rect 3367 2236 3371 2240
rect 3463 2239 3467 2243
rect 111 2196 115 2200
rect 439 2195 443 2199
rect 527 2195 531 2199
rect 615 2195 619 2199
rect 703 2195 707 2199
rect 791 2195 795 2199
rect 879 2195 883 2199
rect 967 2195 971 2199
rect 1055 2195 1059 2199
rect 1143 2195 1147 2199
rect 1231 2195 1235 2199
rect 1319 2195 1323 2199
rect 1767 2196 1771 2200
rect 111 2179 115 2183
rect 439 2176 443 2180
rect 527 2176 531 2180
rect 615 2176 619 2180
rect 703 2176 707 2180
rect 791 2176 795 2180
rect 879 2176 883 2180
rect 967 2176 971 2180
rect 1055 2176 1059 2180
rect 1143 2176 1147 2180
rect 1231 2176 1235 2180
rect 1319 2176 1323 2180
rect 1767 2179 1771 2183
rect 1807 2177 1811 2181
rect 2183 2180 2187 2184
rect 2279 2180 2283 2184
rect 2383 2180 2387 2184
rect 2495 2180 2499 2184
rect 2607 2180 2611 2184
rect 2719 2180 2723 2184
rect 2839 2180 2843 2184
rect 2967 2180 2971 2184
rect 3103 2180 3107 2184
rect 3247 2180 3251 2184
rect 3367 2180 3371 2184
rect 3463 2177 3467 2181
rect 1807 2160 1811 2164
rect 2183 2161 2187 2165
rect 2279 2161 2283 2165
rect 2383 2161 2387 2165
rect 2495 2161 2499 2165
rect 2607 2161 2611 2165
rect 2719 2161 2723 2165
rect 2839 2161 2843 2165
rect 2967 2161 2971 2165
rect 3103 2161 3107 2165
rect 3247 2161 3251 2165
rect 3367 2161 3371 2165
rect 3463 2160 3467 2164
rect 111 2113 115 2117
rect 303 2116 307 2120
rect 407 2116 411 2120
rect 519 2116 523 2120
rect 631 2116 635 2120
rect 743 2116 747 2120
rect 863 2116 867 2120
rect 983 2116 987 2120
rect 1767 2113 1771 2117
rect 1807 2108 1811 2112
rect 2135 2107 2139 2111
rect 2255 2107 2259 2111
rect 2383 2107 2387 2111
rect 2519 2107 2523 2111
rect 2655 2107 2659 2111
rect 2783 2107 2787 2111
rect 2911 2107 2915 2111
rect 3031 2107 3035 2111
rect 3151 2107 3155 2111
rect 3271 2107 3275 2111
rect 3367 2107 3371 2111
rect 3463 2108 3467 2112
rect 111 2096 115 2100
rect 303 2097 307 2101
rect 407 2097 411 2101
rect 519 2097 523 2101
rect 631 2097 635 2101
rect 743 2097 747 2101
rect 863 2097 867 2101
rect 983 2097 987 2101
rect 1767 2096 1771 2100
rect 1807 2091 1811 2095
rect 2135 2088 2139 2092
rect 2255 2088 2259 2092
rect 2383 2088 2387 2092
rect 2519 2088 2523 2092
rect 2655 2088 2659 2092
rect 2783 2088 2787 2092
rect 2911 2088 2915 2092
rect 3031 2088 3035 2092
rect 3151 2088 3155 2092
rect 3271 2088 3275 2092
rect 3367 2088 3371 2092
rect 3463 2091 3467 2095
rect 111 2052 115 2056
rect 255 2051 259 2055
rect 375 2051 379 2055
rect 495 2051 499 2055
rect 615 2051 619 2055
rect 727 2051 731 2055
rect 831 2051 835 2055
rect 935 2051 939 2055
rect 1039 2051 1043 2055
rect 1143 2051 1147 2055
rect 1255 2051 1259 2055
rect 1767 2052 1771 2056
rect 111 2035 115 2039
rect 255 2032 259 2036
rect 375 2032 379 2036
rect 495 2032 499 2036
rect 615 2032 619 2036
rect 727 2032 731 2036
rect 831 2032 835 2036
rect 935 2032 939 2036
rect 1039 2032 1043 2036
rect 1143 2032 1147 2036
rect 1255 2032 1259 2036
rect 1767 2035 1771 2039
rect 1807 2033 1811 2037
rect 2247 2036 2251 2040
rect 2415 2036 2419 2040
rect 2575 2036 2579 2040
rect 2727 2036 2731 2040
rect 2871 2036 2875 2040
rect 3007 2036 3011 2040
rect 3135 2036 3139 2040
rect 3263 2036 3267 2040
rect 3367 2036 3371 2040
rect 3463 2033 3467 2037
rect 1807 2016 1811 2020
rect 2247 2017 2251 2021
rect 2415 2017 2419 2021
rect 2575 2017 2579 2021
rect 2727 2017 2731 2021
rect 2871 2017 2875 2021
rect 3007 2017 3011 2021
rect 3135 2017 3139 2021
rect 3263 2017 3267 2021
rect 3367 2017 3371 2021
rect 3463 2016 3467 2020
rect 111 1985 115 1989
rect 359 1988 363 1992
rect 487 1988 491 1992
rect 623 1988 627 1992
rect 759 1988 763 1992
rect 895 1988 899 1992
rect 1023 1988 1027 1992
rect 1151 1988 1155 1992
rect 1271 1988 1275 1992
rect 1399 1988 1403 1992
rect 1527 1988 1531 1992
rect 1767 1985 1771 1989
rect 111 1968 115 1972
rect 359 1969 363 1973
rect 487 1969 491 1973
rect 623 1969 627 1973
rect 759 1969 763 1973
rect 895 1969 899 1973
rect 1023 1969 1027 1973
rect 1151 1969 1155 1973
rect 1271 1969 1275 1973
rect 1399 1969 1403 1973
rect 1527 1969 1531 1973
rect 1767 1968 1771 1972
rect 1807 1956 1811 1960
rect 1831 1955 1835 1959
rect 1919 1955 1923 1959
rect 2047 1955 2051 1959
rect 2183 1955 2187 1959
rect 2327 1955 2331 1959
rect 2471 1955 2475 1959
rect 2615 1955 2619 1959
rect 2751 1955 2755 1959
rect 2887 1955 2891 1959
rect 3031 1955 3035 1959
rect 3175 1955 3179 1959
rect 3319 1955 3323 1959
rect 3463 1956 3467 1960
rect 1807 1939 1811 1943
rect 1831 1936 1835 1940
rect 1919 1936 1923 1940
rect 2047 1936 2051 1940
rect 2183 1936 2187 1940
rect 2327 1936 2331 1940
rect 2471 1936 2475 1940
rect 2615 1936 2619 1940
rect 2751 1936 2755 1940
rect 2887 1936 2891 1940
rect 3031 1936 3035 1940
rect 3175 1936 3179 1940
rect 3319 1936 3323 1940
rect 3463 1939 3467 1943
rect 111 1924 115 1928
rect 447 1923 451 1927
rect 575 1923 579 1927
rect 711 1923 715 1927
rect 847 1923 851 1927
rect 983 1923 987 1927
rect 1119 1923 1123 1927
rect 1255 1923 1259 1927
rect 1383 1923 1387 1927
rect 1519 1923 1523 1927
rect 1655 1923 1659 1927
rect 1767 1924 1771 1928
rect 111 1907 115 1911
rect 447 1904 451 1908
rect 575 1904 579 1908
rect 711 1904 715 1908
rect 847 1904 851 1908
rect 983 1904 987 1908
rect 1119 1904 1123 1908
rect 1255 1904 1259 1908
rect 1383 1904 1387 1908
rect 1519 1904 1523 1908
rect 1655 1904 1659 1908
rect 1767 1907 1771 1911
rect 1807 1885 1811 1889
rect 1831 1888 1835 1892
rect 1919 1888 1923 1892
rect 2039 1888 2043 1892
rect 2167 1888 2171 1892
rect 2303 1888 2307 1892
rect 2455 1888 2459 1892
rect 2615 1888 2619 1892
rect 2791 1888 2795 1892
rect 2983 1888 2987 1892
rect 3183 1888 3187 1892
rect 3367 1888 3371 1892
rect 3463 1885 3467 1889
rect 1807 1868 1811 1872
rect 1831 1869 1835 1873
rect 1919 1869 1923 1873
rect 2039 1869 2043 1873
rect 2167 1869 2171 1873
rect 2303 1869 2307 1873
rect 2455 1869 2459 1873
rect 2615 1869 2619 1873
rect 2791 1869 2795 1873
rect 2983 1869 2987 1873
rect 3183 1869 3187 1873
rect 3367 1869 3371 1873
rect 3463 1868 3467 1872
rect 111 1857 115 1861
rect 559 1860 563 1864
rect 695 1860 699 1864
rect 831 1860 835 1864
rect 959 1860 963 1864
rect 1079 1860 1083 1864
rect 1199 1860 1203 1864
rect 1327 1860 1331 1864
rect 1455 1860 1459 1864
rect 1767 1857 1771 1861
rect 111 1840 115 1844
rect 559 1841 563 1845
rect 695 1841 699 1845
rect 831 1841 835 1845
rect 959 1841 963 1845
rect 1079 1841 1083 1845
rect 1199 1841 1203 1845
rect 1327 1841 1331 1845
rect 1455 1841 1459 1845
rect 1767 1840 1771 1844
rect 1807 1820 1811 1824
rect 1831 1819 1835 1823
rect 1959 1819 1963 1823
rect 2111 1819 2115 1823
rect 2255 1819 2259 1823
rect 2407 1819 2411 1823
rect 2567 1819 2571 1823
rect 2743 1819 2747 1823
rect 2935 1819 2939 1823
rect 3135 1819 3139 1823
rect 3343 1819 3347 1823
rect 3463 1820 3467 1824
rect 1807 1803 1811 1807
rect 1831 1800 1835 1804
rect 1959 1800 1963 1804
rect 2111 1800 2115 1804
rect 2255 1800 2259 1804
rect 2407 1800 2411 1804
rect 2567 1800 2571 1804
rect 2743 1800 2747 1804
rect 2935 1800 2939 1804
rect 3135 1800 3139 1804
rect 3343 1800 3347 1804
rect 3463 1803 3467 1807
rect 111 1788 115 1792
rect 135 1787 139 1791
rect 223 1787 227 1791
rect 311 1787 315 1791
rect 407 1787 411 1791
rect 527 1787 531 1791
rect 655 1787 659 1791
rect 799 1787 803 1791
rect 943 1787 947 1791
rect 1087 1787 1091 1791
rect 1239 1787 1243 1791
rect 1391 1787 1395 1791
rect 1543 1787 1547 1791
rect 1671 1787 1675 1791
rect 1767 1788 1771 1792
rect 111 1771 115 1775
rect 135 1768 139 1772
rect 223 1768 227 1772
rect 311 1768 315 1772
rect 407 1768 411 1772
rect 527 1768 531 1772
rect 655 1768 659 1772
rect 799 1768 803 1772
rect 943 1768 947 1772
rect 1087 1768 1091 1772
rect 1239 1768 1243 1772
rect 1391 1768 1395 1772
rect 1543 1768 1547 1772
rect 1671 1768 1675 1772
rect 1767 1771 1771 1775
rect 1807 1741 1811 1745
rect 1879 1744 1883 1748
rect 2015 1744 2019 1748
rect 2151 1744 2155 1748
rect 2303 1744 2307 1748
rect 2479 1744 2483 1748
rect 2687 1744 2691 1748
rect 2911 1744 2915 1748
rect 3151 1744 3155 1748
rect 3367 1744 3371 1748
rect 3463 1741 3467 1745
rect 1807 1724 1811 1728
rect 1879 1725 1883 1729
rect 2015 1725 2019 1729
rect 2151 1725 2155 1729
rect 2303 1725 2307 1729
rect 2479 1725 2483 1729
rect 2687 1725 2691 1729
rect 2911 1725 2915 1729
rect 3151 1725 3155 1729
rect 3367 1725 3371 1729
rect 3463 1724 3467 1728
rect 111 1709 115 1713
rect 135 1712 139 1716
rect 247 1712 251 1716
rect 399 1712 403 1716
rect 567 1712 571 1716
rect 751 1712 755 1716
rect 935 1712 939 1716
rect 1119 1712 1123 1716
rect 1311 1712 1315 1716
rect 1503 1712 1507 1716
rect 1671 1712 1675 1716
rect 1767 1709 1771 1713
rect 111 1692 115 1696
rect 135 1693 139 1697
rect 247 1693 251 1697
rect 399 1693 403 1697
rect 567 1693 571 1697
rect 751 1693 755 1697
rect 935 1693 939 1697
rect 1119 1693 1123 1697
rect 1311 1693 1315 1697
rect 1503 1693 1507 1697
rect 1671 1693 1675 1697
rect 1767 1692 1771 1696
rect 1807 1672 1811 1676
rect 1831 1671 1835 1675
rect 1935 1671 1939 1675
rect 2063 1671 2067 1675
rect 2183 1671 2187 1675
rect 2311 1671 2315 1675
rect 2439 1671 2443 1675
rect 2575 1671 2579 1675
rect 2727 1671 2731 1675
rect 2887 1671 2891 1675
rect 3047 1671 3051 1675
rect 3215 1671 3219 1675
rect 3367 1671 3371 1675
rect 3463 1672 3467 1676
rect 1807 1655 1811 1659
rect 1831 1652 1835 1656
rect 1935 1652 1939 1656
rect 2063 1652 2067 1656
rect 2183 1652 2187 1656
rect 2311 1652 2315 1656
rect 2439 1652 2443 1656
rect 2575 1652 2579 1656
rect 2727 1652 2731 1656
rect 2887 1652 2891 1656
rect 3047 1652 3051 1656
rect 3215 1652 3219 1656
rect 3367 1652 3371 1656
rect 3463 1655 3467 1659
rect 111 1644 115 1648
rect 191 1643 195 1647
rect 295 1643 299 1647
rect 407 1643 411 1647
rect 535 1643 539 1647
rect 687 1643 691 1647
rect 855 1643 859 1647
rect 1039 1643 1043 1647
rect 1231 1643 1235 1647
rect 1431 1643 1435 1647
rect 1639 1643 1643 1647
rect 1767 1644 1771 1648
rect 111 1627 115 1631
rect 191 1624 195 1628
rect 295 1624 299 1628
rect 407 1624 411 1628
rect 535 1624 539 1628
rect 687 1624 691 1628
rect 855 1624 859 1628
rect 1039 1624 1043 1628
rect 1231 1624 1235 1628
rect 1431 1624 1435 1628
rect 1639 1624 1643 1628
rect 1767 1627 1771 1631
rect 1807 1597 1811 1601
rect 1831 1600 1835 1604
rect 1943 1600 1947 1604
rect 2087 1600 2091 1604
rect 2231 1600 2235 1604
rect 2367 1600 2371 1604
rect 2503 1600 2507 1604
rect 2639 1600 2643 1604
rect 2767 1600 2771 1604
rect 2895 1600 2899 1604
rect 3015 1600 3019 1604
rect 3135 1600 3139 1604
rect 3263 1600 3267 1604
rect 3367 1600 3371 1604
rect 3463 1597 3467 1601
rect 111 1573 115 1577
rect 327 1576 331 1580
rect 431 1576 435 1580
rect 543 1576 547 1580
rect 671 1576 675 1580
rect 815 1576 819 1580
rect 967 1576 971 1580
rect 1119 1576 1123 1580
rect 1279 1576 1283 1580
rect 1439 1576 1443 1580
rect 1607 1576 1611 1580
rect 1807 1580 1811 1584
rect 1831 1581 1835 1585
rect 1943 1581 1947 1585
rect 2087 1581 2091 1585
rect 2231 1581 2235 1585
rect 2367 1581 2371 1585
rect 2503 1581 2507 1585
rect 2639 1581 2643 1585
rect 2767 1581 2771 1585
rect 2895 1581 2899 1585
rect 3015 1581 3019 1585
rect 3135 1581 3139 1585
rect 3263 1581 3267 1585
rect 3367 1581 3371 1585
rect 3463 1580 3467 1584
rect 1767 1573 1771 1577
rect 111 1556 115 1560
rect 327 1557 331 1561
rect 431 1557 435 1561
rect 543 1557 547 1561
rect 671 1557 675 1561
rect 815 1557 819 1561
rect 967 1557 971 1561
rect 1119 1557 1123 1561
rect 1279 1557 1283 1561
rect 1439 1557 1443 1561
rect 1607 1557 1611 1561
rect 1767 1556 1771 1560
rect 1807 1528 1811 1532
rect 1839 1527 1843 1531
rect 1991 1527 1995 1531
rect 2151 1527 2155 1531
rect 2303 1527 2307 1531
rect 2455 1527 2459 1531
rect 2599 1527 2603 1531
rect 2735 1527 2739 1531
rect 2871 1527 2875 1531
rect 3007 1527 3011 1531
rect 3143 1527 3147 1531
rect 3463 1528 3467 1532
rect 111 1508 115 1512
rect 223 1507 227 1511
rect 343 1507 347 1511
rect 471 1507 475 1511
rect 607 1507 611 1511
rect 751 1507 755 1511
rect 895 1507 899 1511
rect 1047 1507 1051 1511
rect 1199 1507 1203 1511
rect 1351 1507 1355 1511
rect 1503 1507 1507 1511
rect 1767 1508 1771 1512
rect 1807 1511 1811 1515
rect 1839 1508 1843 1512
rect 1991 1508 1995 1512
rect 2151 1508 2155 1512
rect 2303 1508 2307 1512
rect 2455 1508 2459 1512
rect 2599 1508 2603 1512
rect 2735 1508 2739 1512
rect 2871 1508 2875 1512
rect 3007 1508 3011 1512
rect 3143 1508 3147 1512
rect 3463 1511 3467 1515
rect 111 1491 115 1495
rect 223 1488 227 1492
rect 343 1488 347 1492
rect 471 1488 475 1492
rect 607 1488 611 1492
rect 751 1488 755 1492
rect 895 1488 899 1492
rect 1047 1488 1051 1492
rect 1199 1488 1203 1492
rect 1351 1488 1355 1492
rect 1503 1488 1507 1492
rect 1767 1491 1771 1495
rect 1807 1453 1811 1457
rect 1943 1456 1947 1460
rect 2055 1456 2059 1460
rect 2191 1456 2195 1460
rect 2335 1456 2339 1460
rect 2479 1456 2483 1460
rect 2631 1456 2635 1460
rect 2783 1456 2787 1460
rect 2935 1456 2939 1460
rect 3087 1456 3091 1460
rect 3239 1456 3243 1460
rect 3463 1453 3467 1457
rect 111 1433 115 1437
rect 135 1436 139 1440
rect 303 1436 307 1440
rect 471 1436 475 1440
rect 631 1436 635 1440
rect 783 1436 787 1440
rect 927 1436 931 1440
rect 1063 1436 1067 1440
rect 1199 1436 1203 1440
rect 1335 1436 1339 1440
rect 1471 1436 1475 1440
rect 1767 1433 1771 1437
rect 1807 1436 1811 1440
rect 1943 1437 1947 1441
rect 2055 1437 2059 1441
rect 2191 1437 2195 1441
rect 2335 1437 2339 1441
rect 2479 1437 2483 1441
rect 2631 1437 2635 1441
rect 2783 1437 2787 1441
rect 2935 1437 2939 1441
rect 3087 1437 3091 1441
rect 3239 1437 3243 1441
rect 3463 1436 3467 1440
rect 111 1416 115 1420
rect 135 1417 139 1421
rect 303 1417 307 1421
rect 471 1417 475 1421
rect 631 1417 635 1421
rect 783 1417 787 1421
rect 927 1417 931 1421
rect 1063 1417 1067 1421
rect 1199 1417 1203 1421
rect 1335 1417 1339 1421
rect 1471 1417 1475 1421
rect 1767 1416 1771 1420
rect 1807 1384 1811 1388
rect 2095 1383 2099 1387
rect 2199 1383 2203 1387
rect 2319 1383 2323 1387
rect 2455 1383 2459 1387
rect 2599 1383 2603 1387
rect 2743 1383 2747 1387
rect 2887 1383 2891 1387
rect 3031 1383 3035 1387
rect 3175 1383 3179 1387
rect 3327 1383 3331 1387
rect 3463 1384 3467 1388
rect 111 1368 115 1372
rect 135 1367 139 1371
rect 279 1367 283 1371
rect 447 1367 451 1371
rect 607 1367 611 1371
rect 759 1367 763 1371
rect 903 1367 907 1371
rect 1031 1367 1035 1371
rect 1159 1367 1163 1371
rect 1287 1367 1291 1371
rect 1415 1367 1419 1371
rect 1767 1368 1771 1372
rect 1807 1367 1811 1371
rect 2095 1364 2099 1368
rect 2199 1364 2203 1368
rect 2319 1364 2323 1368
rect 2455 1364 2459 1368
rect 2599 1364 2603 1368
rect 2743 1364 2747 1368
rect 2887 1364 2891 1368
rect 3031 1364 3035 1368
rect 3175 1364 3179 1368
rect 3327 1364 3331 1368
rect 3463 1367 3467 1371
rect 111 1351 115 1355
rect 135 1348 139 1352
rect 279 1348 283 1352
rect 447 1348 451 1352
rect 607 1348 611 1352
rect 759 1348 763 1352
rect 903 1348 907 1352
rect 1031 1348 1035 1352
rect 1159 1348 1163 1352
rect 1287 1348 1291 1352
rect 1415 1348 1419 1352
rect 1767 1351 1771 1355
rect 1807 1313 1811 1317
rect 2103 1316 2107 1320
rect 2239 1316 2243 1320
rect 2383 1316 2387 1320
rect 2535 1316 2539 1320
rect 2687 1316 2691 1320
rect 2839 1316 2843 1320
rect 2991 1316 2995 1320
rect 3143 1316 3147 1320
rect 3303 1316 3307 1320
rect 3463 1313 3467 1317
rect 111 1297 115 1301
rect 135 1300 139 1304
rect 279 1300 283 1304
rect 439 1300 443 1304
rect 583 1300 587 1304
rect 719 1300 723 1304
rect 847 1300 851 1304
rect 967 1300 971 1304
rect 1079 1300 1083 1304
rect 1191 1300 1195 1304
rect 1311 1300 1315 1304
rect 1767 1297 1771 1301
rect 1807 1296 1811 1300
rect 2103 1297 2107 1301
rect 2239 1297 2243 1301
rect 2383 1297 2387 1301
rect 2535 1297 2539 1301
rect 2687 1297 2691 1301
rect 2839 1297 2843 1301
rect 2991 1297 2995 1301
rect 3143 1297 3147 1301
rect 3303 1297 3307 1301
rect 3463 1296 3467 1300
rect 111 1280 115 1284
rect 135 1281 139 1285
rect 279 1281 283 1285
rect 439 1281 443 1285
rect 583 1281 587 1285
rect 719 1281 723 1285
rect 847 1281 851 1285
rect 967 1281 971 1285
rect 1079 1281 1083 1285
rect 1191 1281 1195 1285
rect 1311 1281 1315 1285
rect 1767 1280 1771 1284
rect 1807 1252 1811 1256
rect 1935 1251 1939 1255
rect 2063 1251 2067 1255
rect 2199 1251 2203 1255
rect 2343 1251 2347 1255
rect 2495 1251 2499 1255
rect 2655 1251 2659 1255
rect 2815 1251 2819 1255
rect 2975 1251 2979 1255
rect 3143 1251 3147 1255
rect 3463 1252 3467 1256
rect 111 1232 115 1236
rect 135 1231 139 1235
rect 239 1231 243 1235
rect 367 1231 371 1235
rect 495 1231 499 1235
rect 615 1231 619 1235
rect 735 1231 739 1235
rect 847 1231 851 1235
rect 959 1231 963 1235
rect 1071 1231 1075 1235
rect 1191 1231 1195 1235
rect 1767 1232 1771 1236
rect 1807 1235 1811 1239
rect 1935 1232 1939 1236
rect 2063 1232 2067 1236
rect 2199 1232 2203 1236
rect 2343 1232 2347 1236
rect 2495 1232 2499 1236
rect 2655 1232 2659 1236
rect 2815 1232 2819 1236
rect 2975 1232 2979 1236
rect 3143 1232 3147 1236
rect 3463 1235 3467 1239
rect 111 1215 115 1219
rect 135 1212 139 1216
rect 239 1212 243 1216
rect 367 1212 371 1216
rect 495 1212 499 1216
rect 615 1212 619 1216
rect 735 1212 739 1216
rect 847 1212 851 1216
rect 959 1212 963 1216
rect 1071 1212 1075 1216
rect 1191 1212 1195 1216
rect 1767 1215 1771 1219
rect 1807 1185 1811 1189
rect 1831 1188 1835 1192
rect 1935 1188 1939 1192
rect 2079 1188 2083 1192
rect 2231 1188 2235 1192
rect 2391 1188 2395 1192
rect 2543 1188 2547 1192
rect 2695 1188 2699 1192
rect 2847 1188 2851 1192
rect 2999 1188 3003 1192
rect 3159 1188 3163 1192
rect 3463 1185 3467 1189
rect 111 1161 115 1165
rect 135 1164 139 1168
rect 239 1164 243 1168
rect 375 1164 379 1168
rect 511 1164 515 1168
rect 655 1164 659 1168
rect 791 1164 795 1168
rect 927 1164 931 1168
rect 1063 1164 1067 1168
rect 1199 1164 1203 1168
rect 1335 1164 1339 1168
rect 1807 1168 1811 1172
rect 1831 1169 1835 1173
rect 1935 1169 1939 1173
rect 2079 1169 2083 1173
rect 2231 1169 2235 1173
rect 2391 1169 2395 1173
rect 2543 1169 2547 1173
rect 2695 1169 2699 1173
rect 2847 1169 2851 1173
rect 2999 1169 3003 1173
rect 3159 1169 3163 1173
rect 3463 1168 3467 1172
rect 1767 1161 1771 1165
rect 111 1144 115 1148
rect 135 1145 139 1149
rect 239 1145 243 1149
rect 375 1145 379 1149
rect 511 1145 515 1149
rect 655 1145 659 1149
rect 791 1145 795 1149
rect 927 1145 931 1149
rect 1063 1145 1067 1149
rect 1199 1145 1203 1149
rect 1335 1145 1339 1149
rect 1767 1144 1771 1148
rect 1807 1112 1811 1116
rect 1863 1111 1867 1115
rect 1983 1111 1987 1115
rect 2111 1111 2115 1115
rect 2247 1111 2251 1115
rect 2383 1111 2387 1115
rect 2511 1111 2515 1115
rect 2639 1111 2643 1115
rect 2759 1111 2763 1115
rect 2871 1111 2875 1115
rect 2975 1111 2979 1115
rect 3079 1111 3083 1115
rect 3183 1111 3187 1115
rect 3279 1111 3283 1115
rect 3367 1111 3371 1115
rect 3463 1112 3467 1116
rect 111 1096 115 1100
rect 191 1095 195 1099
rect 335 1095 339 1099
rect 495 1095 499 1099
rect 655 1095 659 1099
rect 815 1095 819 1099
rect 967 1095 971 1099
rect 1119 1095 1123 1099
rect 1263 1095 1267 1099
rect 1407 1095 1411 1099
rect 1559 1095 1563 1099
rect 1767 1096 1771 1100
rect 1807 1095 1811 1099
rect 1863 1092 1867 1096
rect 1983 1092 1987 1096
rect 2111 1092 2115 1096
rect 2247 1092 2251 1096
rect 2383 1092 2387 1096
rect 2511 1092 2515 1096
rect 2639 1092 2643 1096
rect 2759 1092 2763 1096
rect 2871 1092 2875 1096
rect 2975 1092 2979 1096
rect 3079 1092 3083 1096
rect 3183 1092 3187 1096
rect 3279 1092 3283 1096
rect 3367 1092 3371 1096
rect 3463 1095 3467 1099
rect 111 1079 115 1083
rect 191 1076 195 1080
rect 335 1076 339 1080
rect 495 1076 499 1080
rect 655 1076 659 1080
rect 815 1076 819 1080
rect 967 1076 971 1080
rect 1119 1076 1123 1080
rect 1263 1076 1267 1080
rect 1407 1076 1411 1080
rect 1559 1076 1563 1080
rect 1767 1079 1771 1083
rect 1807 1037 1811 1041
rect 2103 1040 2107 1044
rect 2191 1040 2195 1044
rect 2279 1040 2283 1044
rect 2367 1040 2371 1044
rect 2455 1040 2459 1044
rect 2543 1040 2547 1044
rect 2631 1040 2635 1044
rect 2719 1040 2723 1044
rect 2807 1040 2811 1044
rect 3463 1037 3467 1041
rect 111 1021 115 1025
rect 327 1024 331 1028
rect 463 1024 467 1028
rect 607 1024 611 1028
rect 767 1024 771 1028
rect 927 1024 931 1028
rect 1079 1024 1083 1028
rect 1231 1024 1235 1028
rect 1383 1024 1387 1028
rect 1535 1024 1539 1028
rect 1671 1024 1675 1028
rect 1767 1021 1771 1025
rect 1807 1020 1811 1024
rect 2103 1021 2107 1025
rect 2191 1021 2195 1025
rect 2279 1021 2283 1025
rect 2367 1021 2371 1025
rect 2455 1021 2459 1025
rect 2543 1021 2547 1025
rect 2631 1021 2635 1025
rect 2719 1021 2723 1025
rect 2807 1021 2811 1025
rect 3463 1020 3467 1024
rect 111 1004 115 1008
rect 327 1005 331 1009
rect 463 1005 467 1009
rect 607 1005 611 1009
rect 767 1005 771 1009
rect 927 1005 931 1009
rect 1079 1005 1083 1009
rect 1231 1005 1235 1009
rect 1383 1005 1387 1009
rect 1535 1005 1539 1009
rect 1671 1005 1675 1009
rect 1767 1004 1771 1008
rect 1807 976 1811 980
rect 2311 975 2315 979
rect 2407 975 2411 979
rect 2511 975 2515 979
rect 2623 975 2627 979
rect 2751 975 2755 979
rect 2895 975 2899 979
rect 3055 975 3059 979
rect 3223 975 3227 979
rect 3367 975 3371 979
rect 3463 976 3467 980
rect 111 956 115 960
rect 471 955 475 959
rect 567 955 571 959
rect 671 955 675 959
rect 783 955 787 959
rect 887 955 891 959
rect 991 955 995 959
rect 1095 955 1099 959
rect 1199 955 1203 959
rect 1295 955 1299 959
rect 1391 955 1395 959
rect 1487 955 1491 959
rect 1583 955 1587 959
rect 1671 955 1675 959
rect 1767 956 1771 960
rect 1807 959 1811 963
rect 2311 956 2315 960
rect 2407 956 2411 960
rect 2511 956 2515 960
rect 2623 956 2627 960
rect 2751 956 2755 960
rect 2895 956 2899 960
rect 3055 956 3059 960
rect 3223 956 3227 960
rect 3367 956 3371 960
rect 3463 959 3467 963
rect 111 939 115 943
rect 471 936 475 940
rect 567 936 571 940
rect 671 936 675 940
rect 783 936 787 940
rect 887 936 891 940
rect 991 936 995 940
rect 1095 936 1099 940
rect 1199 936 1203 940
rect 1295 936 1299 940
rect 1391 936 1395 940
rect 1487 936 1491 940
rect 1583 936 1587 940
rect 1671 936 1675 940
rect 1767 939 1771 943
rect 1807 897 1811 901
rect 1831 900 1835 904
rect 1983 900 1987 904
rect 2151 900 2155 904
rect 2327 900 2331 904
rect 2519 900 2523 904
rect 2719 900 2723 904
rect 2935 900 2939 904
rect 3159 900 3163 904
rect 3367 900 3371 904
rect 3463 897 3467 901
rect 111 885 115 889
rect 607 888 611 892
rect 695 888 699 892
rect 791 888 795 892
rect 895 888 899 892
rect 999 888 1003 892
rect 1111 888 1115 892
rect 1223 888 1227 892
rect 1343 888 1347 892
rect 1463 888 1467 892
rect 1583 888 1587 892
rect 1767 885 1771 889
rect 1807 880 1811 884
rect 1831 881 1835 885
rect 1983 881 1987 885
rect 2151 881 2155 885
rect 2327 881 2331 885
rect 2519 881 2523 885
rect 2719 881 2723 885
rect 2935 881 2939 885
rect 3159 881 3163 885
rect 3367 881 3371 885
rect 3463 880 3467 884
rect 111 868 115 872
rect 607 869 611 873
rect 695 869 699 873
rect 791 869 795 873
rect 895 869 899 873
rect 999 869 1003 873
rect 1111 869 1115 873
rect 1223 869 1227 873
rect 1343 869 1347 873
rect 1463 869 1467 873
rect 1583 869 1587 873
rect 1767 868 1771 872
rect 1807 832 1811 836
rect 1831 831 1835 835
rect 1959 831 1963 835
rect 2087 831 2091 835
rect 2207 831 2211 835
rect 2327 831 2331 835
rect 2463 831 2467 835
rect 2615 831 2619 835
rect 2791 831 2795 835
rect 2983 831 2987 835
rect 3183 831 3187 835
rect 3367 831 3371 835
rect 3463 832 3467 836
rect 111 820 115 824
rect 519 819 523 823
rect 615 819 619 823
rect 719 819 723 823
rect 831 819 835 823
rect 951 819 955 823
rect 1071 819 1075 823
rect 1191 819 1195 823
rect 1311 819 1315 823
rect 1431 819 1435 823
rect 1559 819 1563 823
rect 1767 820 1771 824
rect 1807 815 1811 819
rect 1831 812 1835 816
rect 1959 812 1963 816
rect 2087 812 2091 816
rect 2207 812 2211 816
rect 2327 812 2331 816
rect 2463 812 2467 816
rect 2615 812 2619 816
rect 2791 812 2795 816
rect 2983 812 2987 816
rect 3183 812 3187 816
rect 3367 812 3371 816
rect 3463 815 3467 819
rect 111 803 115 807
rect 519 800 523 804
rect 615 800 619 804
rect 719 800 723 804
rect 831 800 835 804
rect 951 800 955 804
rect 1071 800 1075 804
rect 1191 800 1195 804
rect 1311 800 1315 804
rect 1431 800 1435 804
rect 1559 800 1563 804
rect 1767 803 1771 807
rect 1807 761 1811 765
rect 1879 764 1883 768
rect 2015 764 2019 768
rect 2151 764 2155 768
rect 2287 764 2291 768
rect 2423 764 2427 768
rect 2559 764 2563 768
rect 2711 764 2715 768
rect 2871 764 2875 768
rect 3039 764 3043 768
rect 3215 764 3219 768
rect 3367 764 3371 768
rect 3463 761 3467 765
rect 111 749 115 753
rect 383 752 387 756
rect 471 752 475 756
rect 575 752 579 756
rect 679 752 683 756
rect 791 752 795 756
rect 911 752 915 756
rect 1031 752 1035 756
rect 1159 752 1163 756
rect 1287 752 1291 756
rect 1415 752 1419 756
rect 1767 749 1771 753
rect 1807 744 1811 748
rect 1879 745 1883 749
rect 2015 745 2019 749
rect 2151 745 2155 749
rect 2287 745 2291 749
rect 2423 745 2427 749
rect 2559 745 2563 749
rect 2711 745 2715 749
rect 2871 745 2875 749
rect 3039 745 3043 749
rect 3215 745 3219 749
rect 3367 745 3371 749
rect 3463 744 3467 748
rect 111 732 115 736
rect 383 733 387 737
rect 471 733 475 737
rect 575 733 579 737
rect 679 733 683 737
rect 791 733 795 737
rect 911 733 915 737
rect 1031 733 1035 737
rect 1159 733 1163 737
rect 1287 733 1291 737
rect 1415 733 1419 737
rect 1767 732 1771 736
rect 1807 696 1811 700
rect 1831 695 1835 699
rect 1951 695 1955 699
rect 2103 695 2107 699
rect 2263 695 2267 699
rect 2415 695 2419 699
rect 2567 695 2571 699
rect 2719 695 2723 699
rect 2879 695 2883 699
rect 3039 695 3043 699
rect 3199 695 3203 699
rect 3463 696 3467 700
rect 111 680 115 684
rect 247 679 251 683
rect 343 679 347 683
rect 455 679 459 683
rect 567 679 571 683
rect 695 679 699 683
rect 831 679 835 683
rect 983 679 987 683
rect 1151 679 1155 683
rect 1327 679 1331 683
rect 1511 679 1515 683
rect 1671 679 1675 683
rect 1767 680 1771 684
rect 1807 679 1811 683
rect 1831 676 1835 680
rect 1951 676 1955 680
rect 2103 676 2107 680
rect 2263 676 2267 680
rect 2415 676 2419 680
rect 2567 676 2571 680
rect 2719 676 2723 680
rect 2879 676 2883 680
rect 3039 676 3043 680
rect 3199 676 3203 680
rect 3463 679 3467 683
rect 111 663 115 667
rect 247 660 251 664
rect 343 660 347 664
rect 455 660 459 664
rect 567 660 571 664
rect 695 660 699 664
rect 831 660 835 664
rect 983 660 987 664
rect 1151 660 1155 664
rect 1327 660 1331 664
rect 1511 660 1515 664
rect 1671 660 1675 664
rect 1767 663 1771 667
rect 1807 629 1811 633
rect 1975 632 1979 636
rect 2239 632 2243 636
rect 2479 632 2483 636
rect 2687 632 2691 636
rect 2879 632 2883 636
rect 3055 632 3059 636
rect 3223 632 3227 636
rect 3367 632 3371 636
rect 3463 629 3467 633
rect 111 609 115 613
rect 135 612 139 616
rect 231 612 235 616
rect 359 612 363 616
rect 487 612 491 616
rect 623 612 627 616
rect 767 612 771 616
rect 911 612 915 616
rect 1055 612 1059 616
rect 1207 612 1211 616
rect 1367 612 1371 616
rect 1527 612 1531 616
rect 1671 612 1675 616
rect 1767 609 1771 613
rect 1807 612 1811 616
rect 1975 613 1979 617
rect 2239 613 2243 617
rect 2479 613 2483 617
rect 2687 613 2691 617
rect 2879 613 2883 617
rect 3055 613 3059 617
rect 3223 613 3227 617
rect 3367 613 3371 617
rect 3463 612 3467 616
rect 111 592 115 596
rect 135 593 139 597
rect 231 593 235 597
rect 359 593 363 597
rect 487 593 491 597
rect 623 593 627 597
rect 767 593 771 597
rect 911 593 915 597
rect 1055 593 1059 597
rect 1207 593 1211 597
rect 1367 593 1371 597
rect 1527 593 1531 597
rect 1671 593 1675 597
rect 1767 592 1771 596
rect 1807 560 1811 564
rect 1895 559 1899 563
rect 2015 559 2019 563
rect 2143 559 2147 563
rect 2279 559 2283 563
rect 2423 559 2427 563
rect 2567 559 2571 563
rect 2719 559 2723 563
rect 2871 559 2875 563
rect 3031 559 3035 563
rect 3199 559 3203 563
rect 3367 559 3371 563
rect 3463 560 3467 564
rect 111 544 115 548
rect 135 543 139 547
rect 247 543 251 547
rect 407 543 411 547
rect 583 543 587 547
rect 767 543 771 547
rect 951 543 955 547
rect 1135 543 1139 547
rect 1319 543 1323 547
rect 1503 543 1507 547
rect 1671 543 1675 547
rect 1767 544 1771 548
rect 1807 543 1811 547
rect 1895 540 1899 544
rect 2015 540 2019 544
rect 2143 540 2147 544
rect 2279 540 2283 544
rect 2423 540 2427 544
rect 2567 540 2571 544
rect 2719 540 2723 544
rect 2871 540 2875 544
rect 3031 540 3035 544
rect 3199 540 3203 544
rect 3367 540 3371 544
rect 3463 543 3467 547
rect 111 527 115 531
rect 135 524 139 528
rect 247 524 251 528
rect 407 524 411 528
rect 583 524 587 528
rect 767 524 771 528
rect 951 524 955 528
rect 1135 524 1139 528
rect 1319 524 1323 528
rect 1503 524 1507 528
rect 1671 524 1675 528
rect 1767 527 1771 531
rect 1807 489 1811 493
rect 2135 492 2139 496
rect 2239 492 2243 496
rect 2359 492 2363 496
rect 2487 492 2491 496
rect 2615 492 2619 496
rect 2751 492 2755 496
rect 2879 492 2883 496
rect 3007 492 3011 496
rect 3135 492 3139 496
rect 3263 492 3267 496
rect 3367 492 3371 496
rect 3463 489 3467 493
rect 111 473 115 477
rect 247 476 251 480
rect 399 476 403 480
rect 567 476 571 480
rect 735 476 739 480
rect 903 476 907 480
rect 1063 476 1067 480
rect 1223 476 1227 480
rect 1375 476 1379 480
rect 1527 476 1531 480
rect 1671 476 1675 480
rect 1767 473 1771 477
rect 1807 472 1811 476
rect 2135 473 2139 477
rect 2239 473 2243 477
rect 2359 473 2363 477
rect 2487 473 2491 477
rect 2615 473 2619 477
rect 2751 473 2755 477
rect 2879 473 2883 477
rect 3007 473 3011 477
rect 3135 473 3139 477
rect 3263 473 3267 477
rect 3367 473 3371 477
rect 3463 472 3467 476
rect 111 456 115 460
rect 247 457 251 461
rect 399 457 403 461
rect 567 457 571 461
rect 735 457 739 461
rect 903 457 907 461
rect 1063 457 1067 461
rect 1223 457 1227 461
rect 1375 457 1379 461
rect 1527 457 1531 461
rect 1671 457 1675 461
rect 1767 456 1771 460
rect 1807 420 1811 424
rect 2239 419 2243 423
rect 2335 419 2339 423
rect 2447 419 2451 423
rect 2559 419 2563 423
rect 2679 419 2683 423
rect 2799 419 2803 423
rect 2911 419 2915 423
rect 3023 419 3027 423
rect 3143 419 3147 423
rect 3263 419 3267 423
rect 3367 419 3371 423
rect 3463 420 3467 424
rect 111 408 115 412
rect 519 407 523 411
rect 615 407 619 411
rect 719 407 723 411
rect 823 407 827 411
rect 927 407 931 411
rect 1023 407 1027 411
rect 1127 407 1131 411
rect 1231 407 1235 411
rect 1335 407 1339 411
rect 1439 407 1443 411
rect 1767 408 1771 412
rect 1807 403 1811 407
rect 2239 400 2243 404
rect 2335 400 2339 404
rect 2447 400 2451 404
rect 2559 400 2563 404
rect 2679 400 2683 404
rect 2799 400 2803 404
rect 2911 400 2915 404
rect 3023 400 3027 404
rect 3143 400 3147 404
rect 3263 400 3267 404
rect 3367 400 3371 404
rect 3463 403 3467 407
rect 111 391 115 395
rect 519 388 523 392
rect 615 388 619 392
rect 719 388 723 392
rect 823 388 827 392
rect 927 388 931 392
rect 1023 388 1027 392
rect 1127 388 1131 392
rect 1231 388 1235 392
rect 1335 388 1339 392
rect 1439 388 1443 392
rect 1767 391 1771 395
rect 1807 349 1811 353
rect 2063 352 2067 356
rect 2151 352 2155 356
rect 2247 352 2251 356
rect 2359 352 2363 356
rect 2479 352 2483 356
rect 2615 352 2619 356
rect 2759 352 2763 356
rect 2911 352 2915 356
rect 3063 352 3067 356
rect 3223 352 3227 356
rect 3367 352 3371 356
rect 3463 349 3467 353
rect 111 337 115 341
rect 471 340 475 344
rect 559 340 563 344
rect 647 340 651 344
rect 735 340 739 344
rect 823 340 827 344
rect 911 340 915 344
rect 999 340 1003 344
rect 1087 340 1091 344
rect 1175 340 1179 344
rect 1263 340 1267 344
rect 1767 337 1771 341
rect 1807 332 1811 336
rect 2063 333 2067 337
rect 2151 333 2155 337
rect 2247 333 2251 337
rect 2359 333 2363 337
rect 2479 333 2483 337
rect 2615 333 2619 337
rect 2759 333 2763 337
rect 2911 333 2915 337
rect 3063 333 3067 337
rect 3223 333 3227 337
rect 3367 333 3371 337
rect 3463 332 3467 336
rect 111 320 115 324
rect 471 321 475 325
rect 559 321 563 325
rect 647 321 651 325
rect 735 321 739 325
rect 823 321 827 325
rect 911 321 915 325
rect 999 321 1003 325
rect 1087 321 1091 325
rect 1175 321 1179 325
rect 1263 321 1267 325
rect 1767 320 1771 324
rect 1807 284 1811 288
rect 1927 283 1931 287
rect 2039 283 2043 287
rect 2167 283 2171 287
rect 2303 283 2307 287
rect 2447 283 2451 287
rect 2599 283 2603 287
rect 2759 283 2763 287
rect 2919 283 2923 287
rect 3087 283 3091 287
rect 3255 283 3259 287
rect 3463 284 3467 288
rect 111 272 115 276
rect 279 271 283 275
rect 367 271 371 275
rect 463 271 467 275
rect 559 271 563 275
rect 655 271 659 275
rect 751 271 755 275
rect 847 271 851 275
rect 943 271 947 275
rect 1047 271 1051 275
rect 1151 271 1155 275
rect 1767 272 1771 276
rect 1807 267 1811 271
rect 1927 264 1931 268
rect 2039 264 2043 268
rect 2167 264 2171 268
rect 2303 264 2307 268
rect 2447 264 2451 268
rect 2599 264 2603 268
rect 2759 264 2763 268
rect 2919 264 2923 268
rect 3087 264 3091 268
rect 3255 264 3259 268
rect 3463 267 3467 271
rect 111 255 115 259
rect 279 252 283 256
rect 367 252 371 256
rect 463 252 467 256
rect 559 252 563 256
rect 655 252 659 256
rect 751 252 755 256
rect 847 252 851 256
rect 943 252 947 256
rect 1047 252 1051 256
rect 1151 252 1155 256
rect 1767 255 1771 259
rect 1807 213 1811 217
rect 1831 216 1835 220
rect 1927 216 1931 220
rect 2055 216 2059 220
rect 2199 216 2203 220
rect 2351 216 2355 220
rect 2511 216 2515 220
rect 2679 216 2683 220
rect 2847 216 2851 220
rect 3023 216 3027 220
rect 3207 216 3211 220
rect 3367 216 3371 220
rect 3463 213 3467 217
rect 111 201 115 205
rect 167 204 171 208
rect 343 204 347 208
rect 511 204 515 208
rect 679 204 683 208
rect 839 204 843 208
rect 991 204 995 208
rect 1135 204 1139 208
rect 1279 204 1283 208
rect 1431 204 1435 208
rect 1767 201 1771 205
rect 1807 196 1811 200
rect 1831 197 1835 201
rect 1927 197 1931 201
rect 2055 197 2059 201
rect 2199 197 2203 201
rect 2351 197 2355 201
rect 2511 197 2515 201
rect 2679 197 2683 201
rect 2847 197 2851 201
rect 3023 197 3027 201
rect 3207 197 3211 201
rect 3367 197 3371 201
rect 3463 196 3467 200
rect 111 184 115 188
rect 167 185 171 189
rect 343 185 347 189
rect 511 185 515 189
rect 679 185 683 189
rect 839 185 843 189
rect 991 185 995 189
rect 1135 185 1139 189
rect 1279 185 1283 189
rect 1431 185 1435 189
rect 1767 184 1771 188
rect 1807 132 1811 136
rect 1831 131 1835 135
rect 1919 131 1923 135
rect 2039 131 2043 135
rect 2159 131 2163 135
rect 2279 131 2283 135
rect 2399 131 2403 135
rect 2511 131 2515 135
rect 2623 131 2627 135
rect 2735 131 2739 135
rect 2839 131 2843 135
rect 2943 131 2947 135
rect 3055 131 3059 135
rect 3167 131 3171 135
rect 3279 131 3283 135
rect 3367 131 3371 135
rect 3463 132 3467 136
rect 111 116 115 120
rect 135 115 139 119
rect 223 115 227 119
rect 311 115 315 119
rect 399 115 403 119
rect 487 115 491 119
rect 575 115 579 119
rect 663 115 667 119
rect 751 115 755 119
rect 847 115 851 119
rect 943 115 947 119
rect 1031 115 1035 119
rect 1119 115 1123 119
rect 1215 115 1219 119
rect 1311 115 1315 119
rect 1407 115 1411 119
rect 1495 115 1499 119
rect 1583 115 1587 119
rect 1671 115 1675 119
rect 1767 116 1771 120
rect 1807 115 1811 119
rect 1831 112 1835 116
rect 1919 112 1923 116
rect 2039 112 2043 116
rect 2159 112 2163 116
rect 2279 112 2283 116
rect 2399 112 2403 116
rect 2511 112 2515 116
rect 2623 112 2627 116
rect 2735 112 2739 116
rect 2839 112 2843 116
rect 2943 112 2947 116
rect 3055 112 3059 116
rect 3167 112 3171 116
rect 3279 112 3283 116
rect 3367 112 3371 116
rect 3463 115 3467 119
rect 111 99 115 103
rect 135 96 139 100
rect 223 96 227 100
rect 311 96 315 100
rect 399 96 403 100
rect 487 96 491 100
rect 575 96 579 100
rect 663 96 667 100
rect 751 96 755 100
rect 847 96 851 100
rect 943 96 947 100
rect 1031 96 1035 100
rect 1119 96 1123 100
rect 1215 96 1219 100
rect 1311 96 1315 100
rect 1407 96 1411 100
rect 1495 96 1499 100
rect 1583 96 1587 100
rect 1671 96 1675 100
rect 1767 99 1771 103
<< m3 >>
rect 1807 3522 1811 3523
rect 1807 3517 1811 3518
rect 2007 3522 2011 3523
rect 2007 3517 2011 3518
rect 2239 3522 2243 3523
rect 2239 3517 2243 3518
rect 2455 3522 2459 3523
rect 2455 3517 2459 3518
rect 2655 3522 2659 3523
rect 2655 3517 2659 3518
rect 2855 3522 2859 3523
rect 2855 3517 2859 3518
rect 3047 3522 3051 3523
rect 3047 3517 3051 3518
rect 3247 3522 3251 3523
rect 3247 3517 3251 3518
rect 3463 3522 3467 3523
rect 3463 3517 3467 3518
rect 1808 3501 1810 3517
rect 1806 3500 1812 3501
rect 2008 3500 2010 3517
rect 2240 3500 2242 3517
rect 2456 3500 2458 3517
rect 2656 3500 2658 3517
rect 2856 3500 2858 3517
rect 3048 3500 3050 3517
rect 3248 3500 3250 3517
rect 3464 3501 3466 3517
rect 3462 3500 3468 3501
rect 1806 3496 1807 3500
rect 1811 3496 1812 3500
rect 1806 3495 1812 3496
rect 2006 3499 2012 3500
rect 2006 3495 2007 3499
rect 2011 3495 2012 3499
rect 2006 3494 2012 3495
rect 2238 3499 2244 3500
rect 2238 3495 2239 3499
rect 2243 3495 2244 3499
rect 2238 3494 2244 3495
rect 2454 3499 2460 3500
rect 2454 3495 2455 3499
rect 2459 3495 2460 3499
rect 2454 3494 2460 3495
rect 2654 3499 2660 3500
rect 2654 3495 2655 3499
rect 2659 3495 2660 3499
rect 2654 3494 2660 3495
rect 2854 3499 2860 3500
rect 2854 3495 2855 3499
rect 2859 3495 2860 3499
rect 2854 3494 2860 3495
rect 3046 3499 3052 3500
rect 3046 3495 3047 3499
rect 3051 3495 3052 3499
rect 3046 3494 3052 3495
rect 3246 3499 3252 3500
rect 3246 3495 3247 3499
rect 3251 3495 3252 3499
rect 3462 3496 3463 3500
rect 3467 3496 3468 3500
rect 3462 3495 3468 3496
rect 3246 3494 3252 3495
rect 111 3486 115 3487
rect 111 3481 115 3482
rect 455 3486 459 3487
rect 455 3481 459 3482
rect 543 3486 547 3487
rect 543 3481 547 3482
rect 631 3486 635 3487
rect 631 3481 635 3482
rect 719 3486 723 3487
rect 719 3481 723 3482
rect 807 3486 811 3487
rect 807 3481 811 3482
rect 895 3486 899 3487
rect 895 3481 899 3482
rect 983 3486 987 3487
rect 983 3481 987 3482
rect 1071 3486 1075 3487
rect 1071 3481 1075 3482
rect 1159 3486 1163 3487
rect 1159 3481 1163 3482
rect 1767 3486 1771 3487
rect 1767 3481 1771 3482
rect 1806 3483 1812 3484
rect 112 3465 114 3481
rect 110 3464 116 3465
rect 456 3464 458 3481
rect 544 3464 546 3481
rect 632 3464 634 3481
rect 720 3464 722 3481
rect 808 3464 810 3481
rect 896 3464 898 3481
rect 984 3464 986 3481
rect 1072 3464 1074 3481
rect 1160 3464 1162 3481
rect 1768 3465 1770 3481
rect 1806 3479 1807 3483
rect 1811 3479 1812 3483
rect 3462 3483 3468 3484
rect 1806 3478 1812 3479
rect 2006 3480 2012 3481
rect 1766 3464 1772 3465
rect 110 3460 111 3464
rect 115 3460 116 3464
rect 110 3459 116 3460
rect 454 3463 460 3464
rect 454 3459 455 3463
rect 459 3459 460 3463
rect 454 3458 460 3459
rect 542 3463 548 3464
rect 542 3459 543 3463
rect 547 3459 548 3463
rect 542 3458 548 3459
rect 630 3463 636 3464
rect 630 3459 631 3463
rect 635 3459 636 3463
rect 630 3458 636 3459
rect 718 3463 724 3464
rect 718 3459 719 3463
rect 723 3459 724 3463
rect 718 3458 724 3459
rect 806 3463 812 3464
rect 806 3459 807 3463
rect 811 3459 812 3463
rect 806 3458 812 3459
rect 894 3463 900 3464
rect 894 3459 895 3463
rect 899 3459 900 3463
rect 894 3458 900 3459
rect 982 3463 988 3464
rect 982 3459 983 3463
rect 987 3459 988 3463
rect 982 3458 988 3459
rect 1070 3463 1076 3464
rect 1070 3459 1071 3463
rect 1075 3459 1076 3463
rect 1070 3458 1076 3459
rect 1158 3463 1164 3464
rect 1158 3459 1159 3463
rect 1163 3459 1164 3463
rect 1766 3460 1767 3464
rect 1771 3460 1772 3464
rect 1766 3459 1772 3460
rect 1808 3459 1810 3478
rect 2006 3476 2007 3480
rect 2011 3476 2012 3480
rect 2006 3475 2012 3476
rect 2238 3480 2244 3481
rect 2238 3476 2239 3480
rect 2243 3476 2244 3480
rect 2238 3475 2244 3476
rect 2454 3480 2460 3481
rect 2454 3476 2455 3480
rect 2459 3476 2460 3480
rect 2454 3475 2460 3476
rect 2654 3480 2660 3481
rect 2654 3476 2655 3480
rect 2659 3476 2660 3480
rect 2654 3475 2660 3476
rect 2854 3480 2860 3481
rect 2854 3476 2855 3480
rect 2859 3476 2860 3480
rect 2854 3475 2860 3476
rect 3046 3480 3052 3481
rect 3046 3476 3047 3480
rect 3051 3476 3052 3480
rect 3046 3475 3052 3476
rect 3246 3480 3252 3481
rect 3246 3476 3247 3480
rect 3251 3476 3252 3480
rect 3462 3479 3463 3483
rect 3467 3479 3468 3483
rect 3462 3478 3468 3479
rect 3246 3475 3252 3476
rect 2008 3459 2010 3475
rect 2240 3459 2242 3475
rect 2456 3459 2458 3475
rect 2656 3459 2658 3475
rect 2856 3459 2858 3475
rect 3048 3459 3050 3475
rect 3248 3459 3250 3475
rect 3464 3459 3466 3478
rect 1158 3458 1164 3459
rect 1807 3458 1811 3459
rect 1807 3453 1811 3454
rect 1831 3458 1835 3459
rect 1831 3453 1835 3454
rect 1943 3458 1947 3459
rect 1943 3453 1947 3454
rect 2007 3458 2011 3459
rect 2007 3453 2011 3454
rect 2079 3458 2083 3459
rect 2079 3453 2083 3454
rect 2215 3458 2219 3459
rect 2215 3453 2219 3454
rect 2239 3458 2243 3459
rect 2239 3453 2243 3454
rect 2351 3458 2355 3459
rect 2351 3453 2355 3454
rect 2455 3458 2459 3459
rect 2455 3453 2459 3454
rect 2479 3458 2483 3459
rect 2479 3453 2483 3454
rect 2599 3458 2603 3459
rect 2599 3453 2603 3454
rect 2655 3458 2659 3459
rect 2655 3453 2659 3454
rect 2719 3458 2723 3459
rect 2719 3453 2723 3454
rect 2847 3458 2851 3459
rect 2847 3453 2851 3454
rect 2855 3458 2859 3459
rect 2855 3453 2859 3454
rect 2975 3458 2979 3459
rect 2975 3453 2979 3454
rect 3047 3458 3051 3459
rect 3047 3453 3051 3454
rect 3247 3458 3251 3459
rect 3247 3453 3251 3454
rect 3463 3458 3467 3459
rect 3463 3453 3467 3454
rect 110 3447 116 3448
rect 110 3443 111 3447
rect 115 3443 116 3447
rect 1766 3447 1772 3448
rect 110 3442 116 3443
rect 454 3444 460 3445
rect 112 3423 114 3442
rect 454 3440 455 3444
rect 459 3440 460 3444
rect 454 3439 460 3440
rect 542 3444 548 3445
rect 542 3440 543 3444
rect 547 3440 548 3444
rect 542 3439 548 3440
rect 630 3444 636 3445
rect 630 3440 631 3444
rect 635 3440 636 3444
rect 630 3439 636 3440
rect 718 3444 724 3445
rect 718 3440 719 3444
rect 723 3440 724 3444
rect 718 3439 724 3440
rect 806 3444 812 3445
rect 806 3440 807 3444
rect 811 3440 812 3444
rect 806 3439 812 3440
rect 894 3444 900 3445
rect 894 3440 895 3444
rect 899 3440 900 3444
rect 894 3439 900 3440
rect 982 3444 988 3445
rect 982 3440 983 3444
rect 987 3440 988 3444
rect 982 3439 988 3440
rect 1070 3444 1076 3445
rect 1070 3440 1071 3444
rect 1075 3440 1076 3444
rect 1070 3439 1076 3440
rect 1158 3444 1164 3445
rect 1158 3440 1159 3444
rect 1163 3440 1164 3444
rect 1766 3443 1767 3447
rect 1771 3443 1772 3447
rect 1766 3442 1772 3443
rect 1158 3439 1164 3440
rect 456 3423 458 3439
rect 544 3423 546 3439
rect 632 3423 634 3439
rect 720 3423 722 3439
rect 808 3423 810 3439
rect 896 3423 898 3439
rect 984 3423 986 3439
rect 1072 3423 1074 3439
rect 1160 3423 1162 3439
rect 1768 3423 1770 3442
rect 1808 3434 1810 3453
rect 1832 3437 1834 3453
rect 1944 3437 1946 3453
rect 2080 3437 2082 3453
rect 2216 3437 2218 3453
rect 2352 3437 2354 3453
rect 2480 3437 2482 3453
rect 2600 3437 2602 3453
rect 2720 3437 2722 3453
rect 2848 3437 2850 3453
rect 2976 3437 2978 3453
rect 1830 3436 1836 3437
rect 1806 3433 1812 3434
rect 1806 3429 1807 3433
rect 1811 3429 1812 3433
rect 1830 3432 1831 3436
rect 1835 3432 1836 3436
rect 1830 3431 1836 3432
rect 1942 3436 1948 3437
rect 1942 3432 1943 3436
rect 1947 3432 1948 3436
rect 1942 3431 1948 3432
rect 2078 3436 2084 3437
rect 2078 3432 2079 3436
rect 2083 3432 2084 3436
rect 2078 3431 2084 3432
rect 2214 3436 2220 3437
rect 2214 3432 2215 3436
rect 2219 3432 2220 3436
rect 2214 3431 2220 3432
rect 2350 3436 2356 3437
rect 2350 3432 2351 3436
rect 2355 3432 2356 3436
rect 2350 3431 2356 3432
rect 2478 3436 2484 3437
rect 2478 3432 2479 3436
rect 2483 3432 2484 3436
rect 2478 3431 2484 3432
rect 2598 3436 2604 3437
rect 2598 3432 2599 3436
rect 2603 3432 2604 3436
rect 2598 3431 2604 3432
rect 2718 3436 2724 3437
rect 2718 3432 2719 3436
rect 2723 3432 2724 3436
rect 2718 3431 2724 3432
rect 2846 3436 2852 3437
rect 2846 3432 2847 3436
rect 2851 3432 2852 3436
rect 2846 3431 2852 3432
rect 2974 3436 2980 3437
rect 2974 3432 2975 3436
rect 2979 3432 2980 3436
rect 3464 3434 3466 3453
rect 2974 3431 2980 3432
rect 3462 3433 3468 3434
rect 1806 3428 1812 3429
rect 3462 3429 3463 3433
rect 3467 3429 3468 3433
rect 3462 3428 3468 3429
rect 111 3422 115 3423
rect 111 3417 115 3418
rect 415 3422 419 3423
rect 415 3417 419 3418
rect 455 3422 459 3423
rect 455 3417 459 3418
rect 503 3422 507 3423
rect 503 3417 507 3418
rect 543 3422 547 3423
rect 543 3417 547 3418
rect 591 3422 595 3423
rect 591 3417 595 3418
rect 631 3422 635 3423
rect 631 3417 635 3418
rect 679 3422 683 3423
rect 679 3417 683 3418
rect 719 3422 723 3423
rect 719 3417 723 3418
rect 767 3422 771 3423
rect 767 3417 771 3418
rect 807 3422 811 3423
rect 807 3417 811 3418
rect 855 3422 859 3423
rect 855 3417 859 3418
rect 895 3422 899 3423
rect 895 3417 899 3418
rect 943 3422 947 3423
rect 943 3417 947 3418
rect 983 3422 987 3423
rect 983 3417 987 3418
rect 1031 3422 1035 3423
rect 1031 3417 1035 3418
rect 1071 3422 1075 3423
rect 1071 3417 1075 3418
rect 1119 3422 1123 3423
rect 1119 3417 1123 3418
rect 1159 3422 1163 3423
rect 1159 3417 1163 3418
rect 1207 3422 1211 3423
rect 1207 3417 1211 3418
rect 1303 3422 1307 3423
rect 1303 3417 1307 3418
rect 1767 3422 1771 3423
rect 1767 3417 1771 3418
rect 1830 3417 1836 3418
rect 112 3398 114 3417
rect 416 3401 418 3417
rect 504 3401 506 3417
rect 592 3401 594 3417
rect 680 3401 682 3417
rect 768 3401 770 3417
rect 856 3401 858 3417
rect 944 3401 946 3417
rect 1032 3401 1034 3417
rect 1120 3401 1122 3417
rect 1208 3401 1210 3417
rect 1304 3401 1306 3417
rect 414 3400 420 3401
rect 110 3397 116 3398
rect 110 3393 111 3397
rect 115 3393 116 3397
rect 414 3396 415 3400
rect 419 3396 420 3400
rect 414 3395 420 3396
rect 502 3400 508 3401
rect 502 3396 503 3400
rect 507 3396 508 3400
rect 502 3395 508 3396
rect 590 3400 596 3401
rect 590 3396 591 3400
rect 595 3396 596 3400
rect 590 3395 596 3396
rect 678 3400 684 3401
rect 678 3396 679 3400
rect 683 3396 684 3400
rect 678 3395 684 3396
rect 766 3400 772 3401
rect 766 3396 767 3400
rect 771 3396 772 3400
rect 766 3395 772 3396
rect 854 3400 860 3401
rect 854 3396 855 3400
rect 859 3396 860 3400
rect 854 3395 860 3396
rect 942 3400 948 3401
rect 942 3396 943 3400
rect 947 3396 948 3400
rect 942 3395 948 3396
rect 1030 3400 1036 3401
rect 1030 3396 1031 3400
rect 1035 3396 1036 3400
rect 1030 3395 1036 3396
rect 1118 3400 1124 3401
rect 1118 3396 1119 3400
rect 1123 3396 1124 3400
rect 1118 3395 1124 3396
rect 1206 3400 1212 3401
rect 1206 3396 1207 3400
rect 1211 3396 1212 3400
rect 1206 3395 1212 3396
rect 1302 3400 1308 3401
rect 1302 3396 1303 3400
rect 1307 3396 1308 3400
rect 1768 3398 1770 3417
rect 1806 3416 1812 3417
rect 1806 3412 1807 3416
rect 1811 3412 1812 3416
rect 1830 3413 1831 3417
rect 1835 3413 1836 3417
rect 1830 3412 1836 3413
rect 1942 3417 1948 3418
rect 1942 3413 1943 3417
rect 1947 3413 1948 3417
rect 1942 3412 1948 3413
rect 2078 3417 2084 3418
rect 2078 3413 2079 3417
rect 2083 3413 2084 3417
rect 2078 3412 2084 3413
rect 2214 3417 2220 3418
rect 2214 3413 2215 3417
rect 2219 3413 2220 3417
rect 2214 3412 2220 3413
rect 2350 3417 2356 3418
rect 2350 3413 2351 3417
rect 2355 3413 2356 3417
rect 2350 3412 2356 3413
rect 2478 3417 2484 3418
rect 2478 3413 2479 3417
rect 2483 3413 2484 3417
rect 2478 3412 2484 3413
rect 2598 3417 2604 3418
rect 2598 3413 2599 3417
rect 2603 3413 2604 3417
rect 2598 3412 2604 3413
rect 2718 3417 2724 3418
rect 2718 3413 2719 3417
rect 2723 3413 2724 3417
rect 2718 3412 2724 3413
rect 2846 3417 2852 3418
rect 2846 3413 2847 3417
rect 2851 3413 2852 3417
rect 2846 3412 2852 3413
rect 2974 3417 2980 3418
rect 2974 3413 2975 3417
rect 2979 3413 2980 3417
rect 2974 3412 2980 3413
rect 3462 3416 3468 3417
rect 3462 3412 3463 3416
rect 3467 3412 3468 3416
rect 1806 3411 1812 3412
rect 1302 3395 1308 3396
rect 1766 3397 1772 3398
rect 110 3392 116 3393
rect 1766 3393 1767 3397
rect 1771 3393 1772 3397
rect 1766 3392 1772 3393
rect 1808 3387 1810 3411
rect 1832 3387 1834 3412
rect 1944 3387 1946 3412
rect 2080 3387 2082 3412
rect 2216 3387 2218 3412
rect 2352 3387 2354 3412
rect 2480 3387 2482 3412
rect 2600 3387 2602 3412
rect 2720 3387 2722 3412
rect 2848 3387 2850 3412
rect 2976 3387 2978 3412
rect 3462 3411 3468 3412
rect 3464 3387 3466 3411
rect 1807 3386 1811 3387
rect 414 3381 420 3382
rect 110 3380 116 3381
rect 110 3376 111 3380
rect 115 3376 116 3380
rect 414 3377 415 3381
rect 419 3377 420 3381
rect 414 3376 420 3377
rect 502 3381 508 3382
rect 502 3377 503 3381
rect 507 3377 508 3381
rect 502 3376 508 3377
rect 590 3381 596 3382
rect 590 3377 591 3381
rect 595 3377 596 3381
rect 590 3376 596 3377
rect 678 3381 684 3382
rect 678 3377 679 3381
rect 683 3377 684 3381
rect 678 3376 684 3377
rect 766 3381 772 3382
rect 766 3377 767 3381
rect 771 3377 772 3381
rect 766 3376 772 3377
rect 854 3381 860 3382
rect 854 3377 855 3381
rect 859 3377 860 3381
rect 854 3376 860 3377
rect 942 3381 948 3382
rect 942 3377 943 3381
rect 947 3377 948 3381
rect 942 3376 948 3377
rect 1030 3381 1036 3382
rect 1030 3377 1031 3381
rect 1035 3377 1036 3381
rect 1030 3376 1036 3377
rect 1118 3381 1124 3382
rect 1118 3377 1119 3381
rect 1123 3377 1124 3381
rect 1118 3376 1124 3377
rect 1206 3381 1212 3382
rect 1206 3377 1207 3381
rect 1211 3377 1212 3381
rect 1206 3376 1212 3377
rect 1302 3381 1308 3382
rect 1807 3381 1811 3382
rect 1831 3386 1835 3387
rect 1831 3381 1835 3382
rect 1943 3386 1947 3387
rect 1943 3381 1947 3382
rect 1951 3386 1955 3387
rect 1951 3381 1955 3382
rect 2079 3386 2083 3387
rect 2079 3381 2083 3382
rect 2095 3386 2099 3387
rect 2095 3381 2099 3382
rect 2215 3386 2219 3387
rect 2215 3381 2219 3382
rect 2239 3386 2243 3387
rect 2239 3381 2243 3382
rect 2351 3386 2355 3387
rect 2351 3381 2355 3382
rect 2383 3386 2387 3387
rect 2383 3381 2387 3382
rect 2479 3386 2483 3387
rect 2479 3381 2483 3382
rect 2519 3386 2523 3387
rect 2519 3381 2523 3382
rect 2599 3386 2603 3387
rect 2599 3381 2603 3382
rect 2647 3386 2651 3387
rect 2647 3381 2651 3382
rect 2719 3386 2723 3387
rect 2719 3381 2723 3382
rect 2775 3386 2779 3387
rect 2775 3381 2779 3382
rect 2847 3386 2851 3387
rect 2847 3381 2851 3382
rect 2903 3386 2907 3387
rect 2903 3381 2907 3382
rect 2975 3386 2979 3387
rect 2975 3381 2979 3382
rect 3039 3386 3043 3387
rect 3039 3381 3043 3382
rect 3463 3386 3467 3387
rect 3463 3381 3467 3382
rect 1302 3377 1303 3381
rect 1307 3377 1308 3381
rect 1302 3376 1308 3377
rect 1766 3380 1772 3381
rect 1766 3376 1767 3380
rect 1771 3376 1772 3380
rect 110 3375 116 3376
rect 112 3355 114 3375
rect 416 3355 418 3376
rect 504 3355 506 3376
rect 592 3355 594 3376
rect 680 3355 682 3376
rect 768 3355 770 3376
rect 856 3355 858 3376
rect 944 3355 946 3376
rect 1032 3355 1034 3376
rect 1120 3355 1122 3376
rect 1208 3355 1210 3376
rect 1304 3355 1306 3376
rect 1766 3375 1772 3376
rect 1768 3355 1770 3375
rect 1808 3365 1810 3381
rect 1806 3364 1812 3365
rect 1832 3364 1834 3381
rect 1952 3364 1954 3381
rect 2096 3364 2098 3381
rect 2240 3364 2242 3381
rect 2384 3364 2386 3381
rect 2520 3364 2522 3381
rect 2648 3364 2650 3381
rect 2776 3364 2778 3381
rect 2904 3364 2906 3381
rect 3040 3364 3042 3381
rect 3464 3365 3466 3381
rect 3462 3364 3468 3365
rect 1806 3360 1807 3364
rect 1811 3360 1812 3364
rect 1806 3359 1812 3360
rect 1830 3363 1836 3364
rect 1830 3359 1831 3363
rect 1835 3359 1836 3363
rect 1830 3358 1836 3359
rect 1950 3363 1956 3364
rect 1950 3359 1951 3363
rect 1955 3359 1956 3363
rect 1950 3358 1956 3359
rect 2094 3363 2100 3364
rect 2094 3359 2095 3363
rect 2099 3359 2100 3363
rect 2094 3358 2100 3359
rect 2238 3363 2244 3364
rect 2238 3359 2239 3363
rect 2243 3359 2244 3363
rect 2238 3358 2244 3359
rect 2382 3363 2388 3364
rect 2382 3359 2383 3363
rect 2387 3359 2388 3363
rect 2382 3358 2388 3359
rect 2518 3363 2524 3364
rect 2518 3359 2519 3363
rect 2523 3359 2524 3363
rect 2518 3358 2524 3359
rect 2646 3363 2652 3364
rect 2646 3359 2647 3363
rect 2651 3359 2652 3363
rect 2646 3358 2652 3359
rect 2774 3363 2780 3364
rect 2774 3359 2775 3363
rect 2779 3359 2780 3363
rect 2774 3358 2780 3359
rect 2902 3363 2908 3364
rect 2902 3359 2903 3363
rect 2907 3359 2908 3363
rect 2902 3358 2908 3359
rect 3038 3363 3044 3364
rect 3038 3359 3039 3363
rect 3043 3359 3044 3363
rect 3462 3360 3463 3364
rect 3467 3360 3468 3364
rect 3462 3359 3468 3360
rect 3038 3358 3044 3359
rect 111 3354 115 3355
rect 111 3349 115 3350
rect 399 3354 403 3355
rect 399 3349 403 3350
rect 415 3354 419 3355
rect 415 3349 419 3350
rect 495 3354 499 3355
rect 495 3349 499 3350
rect 503 3354 507 3355
rect 503 3349 507 3350
rect 591 3354 595 3355
rect 591 3349 595 3350
rect 599 3354 603 3355
rect 599 3349 603 3350
rect 679 3354 683 3355
rect 679 3349 683 3350
rect 703 3354 707 3355
rect 703 3349 707 3350
rect 767 3354 771 3355
rect 767 3349 771 3350
rect 807 3354 811 3355
rect 807 3349 811 3350
rect 855 3354 859 3355
rect 855 3349 859 3350
rect 911 3354 915 3355
rect 911 3349 915 3350
rect 943 3354 947 3355
rect 943 3349 947 3350
rect 1015 3354 1019 3355
rect 1015 3349 1019 3350
rect 1031 3354 1035 3355
rect 1031 3349 1035 3350
rect 1119 3354 1123 3355
rect 1119 3349 1123 3350
rect 1207 3354 1211 3355
rect 1207 3349 1211 3350
rect 1223 3354 1227 3355
rect 1223 3349 1227 3350
rect 1303 3354 1307 3355
rect 1303 3349 1307 3350
rect 1327 3354 1331 3355
rect 1327 3349 1331 3350
rect 1767 3354 1771 3355
rect 1767 3349 1771 3350
rect 112 3333 114 3349
rect 110 3332 116 3333
rect 400 3332 402 3349
rect 496 3332 498 3349
rect 600 3332 602 3349
rect 704 3332 706 3349
rect 808 3332 810 3349
rect 912 3332 914 3349
rect 1016 3332 1018 3349
rect 1120 3332 1122 3349
rect 1224 3332 1226 3349
rect 1328 3332 1330 3349
rect 1768 3333 1770 3349
rect 1806 3347 1812 3348
rect 1806 3343 1807 3347
rect 1811 3343 1812 3347
rect 3462 3347 3468 3348
rect 1806 3342 1812 3343
rect 1830 3344 1836 3345
rect 1766 3332 1772 3333
rect 110 3328 111 3332
rect 115 3328 116 3332
rect 110 3327 116 3328
rect 398 3331 404 3332
rect 398 3327 399 3331
rect 403 3327 404 3331
rect 398 3326 404 3327
rect 494 3331 500 3332
rect 494 3327 495 3331
rect 499 3327 500 3331
rect 494 3326 500 3327
rect 598 3331 604 3332
rect 598 3327 599 3331
rect 603 3327 604 3331
rect 598 3326 604 3327
rect 702 3331 708 3332
rect 702 3327 703 3331
rect 707 3327 708 3331
rect 702 3326 708 3327
rect 806 3331 812 3332
rect 806 3327 807 3331
rect 811 3327 812 3331
rect 806 3326 812 3327
rect 910 3331 916 3332
rect 910 3327 911 3331
rect 915 3327 916 3331
rect 910 3326 916 3327
rect 1014 3331 1020 3332
rect 1014 3327 1015 3331
rect 1019 3327 1020 3331
rect 1014 3326 1020 3327
rect 1118 3331 1124 3332
rect 1118 3327 1119 3331
rect 1123 3327 1124 3331
rect 1118 3326 1124 3327
rect 1222 3331 1228 3332
rect 1222 3327 1223 3331
rect 1227 3327 1228 3331
rect 1222 3326 1228 3327
rect 1326 3331 1332 3332
rect 1326 3327 1327 3331
rect 1331 3327 1332 3331
rect 1766 3328 1767 3332
rect 1771 3328 1772 3332
rect 1766 3327 1772 3328
rect 1326 3326 1332 3327
rect 110 3315 116 3316
rect 110 3311 111 3315
rect 115 3311 116 3315
rect 1766 3315 1772 3316
rect 1808 3315 1810 3342
rect 1830 3340 1831 3344
rect 1835 3340 1836 3344
rect 1830 3339 1836 3340
rect 1950 3344 1956 3345
rect 1950 3340 1951 3344
rect 1955 3340 1956 3344
rect 1950 3339 1956 3340
rect 2094 3344 2100 3345
rect 2094 3340 2095 3344
rect 2099 3340 2100 3344
rect 2094 3339 2100 3340
rect 2238 3344 2244 3345
rect 2238 3340 2239 3344
rect 2243 3340 2244 3344
rect 2238 3339 2244 3340
rect 2382 3344 2388 3345
rect 2382 3340 2383 3344
rect 2387 3340 2388 3344
rect 2382 3339 2388 3340
rect 2518 3344 2524 3345
rect 2518 3340 2519 3344
rect 2523 3340 2524 3344
rect 2518 3339 2524 3340
rect 2646 3344 2652 3345
rect 2646 3340 2647 3344
rect 2651 3340 2652 3344
rect 2646 3339 2652 3340
rect 2774 3344 2780 3345
rect 2774 3340 2775 3344
rect 2779 3340 2780 3344
rect 2774 3339 2780 3340
rect 2902 3344 2908 3345
rect 2902 3340 2903 3344
rect 2907 3340 2908 3344
rect 2902 3339 2908 3340
rect 3038 3344 3044 3345
rect 3038 3340 3039 3344
rect 3043 3340 3044 3344
rect 3462 3343 3463 3347
rect 3467 3343 3468 3347
rect 3462 3342 3468 3343
rect 3038 3339 3044 3340
rect 1832 3315 1834 3339
rect 1952 3315 1954 3339
rect 2096 3315 2098 3339
rect 2240 3315 2242 3339
rect 2384 3315 2386 3339
rect 2520 3315 2522 3339
rect 2648 3315 2650 3339
rect 2776 3315 2778 3339
rect 2904 3315 2906 3339
rect 3040 3315 3042 3339
rect 3464 3315 3466 3342
rect 110 3310 116 3311
rect 398 3312 404 3313
rect 112 3287 114 3310
rect 398 3308 399 3312
rect 403 3308 404 3312
rect 398 3307 404 3308
rect 494 3312 500 3313
rect 494 3308 495 3312
rect 499 3308 500 3312
rect 494 3307 500 3308
rect 598 3312 604 3313
rect 598 3308 599 3312
rect 603 3308 604 3312
rect 598 3307 604 3308
rect 702 3312 708 3313
rect 702 3308 703 3312
rect 707 3308 708 3312
rect 702 3307 708 3308
rect 806 3312 812 3313
rect 806 3308 807 3312
rect 811 3308 812 3312
rect 806 3307 812 3308
rect 910 3312 916 3313
rect 910 3308 911 3312
rect 915 3308 916 3312
rect 910 3307 916 3308
rect 1014 3312 1020 3313
rect 1014 3308 1015 3312
rect 1019 3308 1020 3312
rect 1014 3307 1020 3308
rect 1118 3312 1124 3313
rect 1118 3308 1119 3312
rect 1123 3308 1124 3312
rect 1118 3307 1124 3308
rect 1222 3312 1228 3313
rect 1222 3308 1223 3312
rect 1227 3308 1228 3312
rect 1222 3307 1228 3308
rect 1326 3312 1332 3313
rect 1326 3308 1327 3312
rect 1331 3308 1332 3312
rect 1766 3311 1767 3315
rect 1771 3311 1772 3315
rect 1766 3310 1772 3311
rect 1807 3314 1811 3315
rect 1326 3307 1332 3308
rect 400 3287 402 3307
rect 496 3287 498 3307
rect 600 3287 602 3307
rect 704 3287 706 3307
rect 808 3287 810 3307
rect 912 3287 914 3307
rect 1016 3287 1018 3307
rect 1120 3287 1122 3307
rect 1224 3287 1226 3307
rect 1328 3287 1330 3307
rect 1768 3287 1770 3310
rect 1807 3309 1811 3310
rect 1831 3314 1835 3315
rect 1831 3309 1835 3310
rect 1951 3314 1955 3315
rect 1951 3309 1955 3310
rect 1975 3314 1979 3315
rect 1975 3309 1979 3310
rect 2095 3314 2099 3315
rect 2095 3309 2099 3310
rect 2151 3314 2155 3315
rect 2151 3309 2155 3310
rect 2239 3314 2243 3315
rect 2239 3309 2243 3310
rect 2335 3314 2339 3315
rect 2335 3309 2339 3310
rect 2383 3314 2387 3315
rect 2383 3309 2387 3310
rect 2511 3314 2515 3315
rect 2511 3309 2515 3310
rect 2519 3314 2523 3315
rect 2519 3309 2523 3310
rect 2647 3314 2651 3315
rect 2647 3309 2651 3310
rect 2679 3314 2683 3315
rect 2679 3309 2683 3310
rect 2775 3314 2779 3315
rect 2775 3309 2779 3310
rect 2831 3314 2835 3315
rect 2831 3309 2835 3310
rect 2903 3314 2907 3315
rect 2903 3309 2907 3310
rect 2975 3314 2979 3315
rect 2975 3309 2979 3310
rect 3039 3314 3043 3315
rect 3039 3309 3043 3310
rect 3111 3314 3115 3315
rect 3111 3309 3115 3310
rect 3247 3314 3251 3315
rect 3247 3309 3251 3310
rect 3367 3314 3371 3315
rect 3367 3309 3371 3310
rect 3463 3314 3467 3315
rect 3463 3309 3467 3310
rect 1808 3290 1810 3309
rect 1832 3293 1834 3309
rect 1976 3293 1978 3309
rect 2152 3293 2154 3309
rect 2336 3293 2338 3309
rect 2512 3293 2514 3309
rect 2680 3293 2682 3309
rect 2832 3293 2834 3309
rect 2976 3293 2978 3309
rect 3112 3293 3114 3309
rect 3248 3293 3250 3309
rect 3368 3293 3370 3309
rect 1830 3292 1836 3293
rect 1806 3289 1812 3290
rect 111 3286 115 3287
rect 111 3281 115 3282
rect 383 3286 387 3287
rect 383 3281 387 3282
rect 399 3286 403 3287
rect 399 3281 403 3282
rect 495 3286 499 3287
rect 495 3281 499 3282
rect 599 3286 603 3287
rect 599 3281 603 3282
rect 607 3286 611 3287
rect 607 3281 611 3282
rect 703 3286 707 3287
rect 703 3281 707 3282
rect 727 3286 731 3287
rect 727 3281 731 3282
rect 807 3286 811 3287
rect 807 3281 811 3282
rect 847 3286 851 3287
rect 847 3281 851 3282
rect 911 3286 915 3287
rect 911 3281 915 3282
rect 967 3286 971 3287
rect 967 3281 971 3282
rect 1015 3286 1019 3287
rect 1015 3281 1019 3282
rect 1087 3286 1091 3287
rect 1087 3281 1091 3282
rect 1119 3286 1123 3287
rect 1119 3281 1123 3282
rect 1207 3286 1211 3287
rect 1207 3281 1211 3282
rect 1223 3286 1227 3287
rect 1223 3281 1227 3282
rect 1327 3286 1331 3287
rect 1327 3281 1331 3282
rect 1335 3286 1339 3287
rect 1335 3281 1339 3282
rect 1767 3286 1771 3287
rect 1806 3285 1807 3289
rect 1811 3285 1812 3289
rect 1830 3288 1831 3292
rect 1835 3288 1836 3292
rect 1830 3287 1836 3288
rect 1974 3292 1980 3293
rect 1974 3288 1975 3292
rect 1979 3288 1980 3292
rect 1974 3287 1980 3288
rect 2150 3292 2156 3293
rect 2150 3288 2151 3292
rect 2155 3288 2156 3292
rect 2150 3287 2156 3288
rect 2334 3292 2340 3293
rect 2334 3288 2335 3292
rect 2339 3288 2340 3292
rect 2334 3287 2340 3288
rect 2510 3292 2516 3293
rect 2510 3288 2511 3292
rect 2515 3288 2516 3292
rect 2510 3287 2516 3288
rect 2678 3292 2684 3293
rect 2678 3288 2679 3292
rect 2683 3288 2684 3292
rect 2678 3287 2684 3288
rect 2830 3292 2836 3293
rect 2830 3288 2831 3292
rect 2835 3288 2836 3292
rect 2830 3287 2836 3288
rect 2974 3292 2980 3293
rect 2974 3288 2975 3292
rect 2979 3288 2980 3292
rect 2974 3287 2980 3288
rect 3110 3292 3116 3293
rect 3110 3288 3111 3292
rect 3115 3288 3116 3292
rect 3110 3287 3116 3288
rect 3246 3292 3252 3293
rect 3246 3288 3247 3292
rect 3251 3288 3252 3292
rect 3246 3287 3252 3288
rect 3366 3292 3372 3293
rect 3366 3288 3367 3292
rect 3371 3288 3372 3292
rect 3464 3290 3466 3309
rect 3366 3287 3372 3288
rect 3462 3289 3468 3290
rect 1806 3284 1812 3285
rect 3462 3285 3463 3289
rect 3467 3285 3468 3289
rect 3462 3284 3468 3285
rect 1767 3281 1771 3282
rect 112 3262 114 3281
rect 384 3265 386 3281
rect 496 3265 498 3281
rect 608 3265 610 3281
rect 728 3265 730 3281
rect 848 3265 850 3281
rect 968 3265 970 3281
rect 1088 3265 1090 3281
rect 1208 3265 1210 3281
rect 1336 3265 1338 3281
rect 382 3264 388 3265
rect 110 3261 116 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 382 3260 383 3264
rect 387 3260 388 3264
rect 382 3259 388 3260
rect 494 3264 500 3265
rect 494 3260 495 3264
rect 499 3260 500 3264
rect 494 3259 500 3260
rect 606 3264 612 3265
rect 606 3260 607 3264
rect 611 3260 612 3264
rect 606 3259 612 3260
rect 726 3264 732 3265
rect 726 3260 727 3264
rect 731 3260 732 3264
rect 726 3259 732 3260
rect 846 3264 852 3265
rect 846 3260 847 3264
rect 851 3260 852 3264
rect 846 3259 852 3260
rect 966 3264 972 3265
rect 966 3260 967 3264
rect 971 3260 972 3264
rect 966 3259 972 3260
rect 1086 3264 1092 3265
rect 1086 3260 1087 3264
rect 1091 3260 1092 3264
rect 1086 3259 1092 3260
rect 1206 3264 1212 3265
rect 1206 3260 1207 3264
rect 1211 3260 1212 3264
rect 1206 3259 1212 3260
rect 1334 3264 1340 3265
rect 1334 3260 1335 3264
rect 1339 3260 1340 3264
rect 1768 3262 1770 3281
rect 1830 3273 1836 3274
rect 1806 3272 1812 3273
rect 1806 3268 1807 3272
rect 1811 3268 1812 3272
rect 1830 3269 1831 3273
rect 1835 3269 1836 3273
rect 1830 3268 1836 3269
rect 1974 3273 1980 3274
rect 1974 3269 1975 3273
rect 1979 3269 1980 3273
rect 1974 3268 1980 3269
rect 2150 3273 2156 3274
rect 2150 3269 2151 3273
rect 2155 3269 2156 3273
rect 2150 3268 2156 3269
rect 2334 3273 2340 3274
rect 2334 3269 2335 3273
rect 2339 3269 2340 3273
rect 2334 3268 2340 3269
rect 2510 3273 2516 3274
rect 2510 3269 2511 3273
rect 2515 3269 2516 3273
rect 2510 3268 2516 3269
rect 2678 3273 2684 3274
rect 2678 3269 2679 3273
rect 2683 3269 2684 3273
rect 2678 3268 2684 3269
rect 2830 3273 2836 3274
rect 2830 3269 2831 3273
rect 2835 3269 2836 3273
rect 2830 3268 2836 3269
rect 2974 3273 2980 3274
rect 2974 3269 2975 3273
rect 2979 3269 2980 3273
rect 2974 3268 2980 3269
rect 3110 3273 3116 3274
rect 3110 3269 3111 3273
rect 3115 3269 3116 3273
rect 3110 3268 3116 3269
rect 3246 3273 3252 3274
rect 3246 3269 3247 3273
rect 3251 3269 3252 3273
rect 3246 3268 3252 3269
rect 3366 3273 3372 3274
rect 3366 3269 3367 3273
rect 3371 3269 3372 3273
rect 3366 3268 3372 3269
rect 3462 3272 3468 3273
rect 3462 3268 3463 3272
rect 3467 3268 3468 3272
rect 1806 3267 1812 3268
rect 1334 3259 1340 3260
rect 1766 3261 1772 3262
rect 110 3256 116 3257
rect 1766 3257 1767 3261
rect 1771 3257 1772 3261
rect 1766 3256 1772 3257
rect 382 3245 388 3246
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 382 3241 383 3245
rect 387 3241 388 3245
rect 382 3240 388 3241
rect 494 3245 500 3246
rect 494 3241 495 3245
rect 499 3241 500 3245
rect 494 3240 500 3241
rect 606 3245 612 3246
rect 606 3241 607 3245
rect 611 3241 612 3245
rect 606 3240 612 3241
rect 726 3245 732 3246
rect 726 3241 727 3245
rect 731 3241 732 3245
rect 726 3240 732 3241
rect 846 3245 852 3246
rect 846 3241 847 3245
rect 851 3241 852 3245
rect 846 3240 852 3241
rect 966 3245 972 3246
rect 966 3241 967 3245
rect 971 3241 972 3245
rect 966 3240 972 3241
rect 1086 3245 1092 3246
rect 1086 3241 1087 3245
rect 1091 3241 1092 3245
rect 1086 3240 1092 3241
rect 1206 3245 1212 3246
rect 1206 3241 1207 3245
rect 1211 3241 1212 3245
rect 1206 3240 1212 3241
rect 1334 3245 1340 3246
rect 1334 3241 1335 3245
rect 1339 3241 1340 3245
rect 1334 3240 1340 3241
rect 1766 3244 1772 3245
rect 1766 3240 1767 3244
rect 1771 3240 1772 3244
rect 1808 3243 1810 3267
rect 1832 3243 1834 3268
rect 1976 3243 1978 3268
rect 2152 3243 2154 3268
rect 2336 3243 2338 3268
rect 2512 3243 2514 3268
rect 2680 3243 2682 3268
rect 2832 3243 2834 3268
rect 2976 3243 2978 3268
rect 3112 3243 3114 3268
rect 3248 3243 3250 3268
rect 3368 3243 3370 3268
rect 3462 3267 3468 3268
rect 3464 3243 3466 3267
rect 110 3239 116 3240
rect 112 3219 114 3239
rect 384 3219 386 3240
rect 496 3219 498 3240
rect 608 3219 610 3240
rect 728 3219 730 3240
rect 848 3219 850 3240
rect 968 3219 970 3240
rect 1088 3219 1090 3240
rect 1208 3219 1210 3240
rect 1336 3219 1338 3240
rect 1766 3239 1772 3240
rect 1807 3242 1811 3243
rect 1768 3219 1770 3239
rect 1807 3237 1811 3238
rect 1831 3242 1835 3243
rect 1831 3237 1835 3238
rect 1975 3242 1979 3243
rect 1975 3237 1979 3238
rect 2031 3242 2035 3243
rect 2031 3237 2035 3238
rect 2151 3242 2155 3243
rect 2151 3237 2155 3238
rect 2247 3242 2251 3243
rect 2247 3237 2251 3238
rect 2335 3242 2339 3243
rect 2335 3237 2339 3238
rect 2455 3242 2459 3243
rect 2455 3237 2459 3238
rect 2511 3242 2515 3243
rect 2511 3237 2515 3238
rect 2655 3242 2659 3243
rect 2655 3237 2659 3238
rect 2679 3242 2683 3243
rect 2679 3237 2683 3238
rect 2831 3242 2835 3243
rect 2831 3237 2835 3238
rect 2839 3242 2843 3243
rect 2839 3237 2843 3238
rect 2975 3242 2979 3243
rect 2975 3237 2979 3238
rect 3023 3242 3027 3243
rect 3023 3237 3027 3238
rect 3111 3242 3115 3243
rect 3111 3237 3115 3238
rect 3207 3242 3211 3243
rect 3207 3237 3211 3238
rect 3247 3242 3251 3243
rect 3247 3237 3251 3238
rect 3367 3242 3371 3243
rect 3367 3237 3371 3238
rect 3463 3242 3467 3243
rect 3463 3237 3467 3238
rect 1808 3221 1810 3237
rect 1806 3220 1812 3221
rect 1832 3220 1834 3237
rect 2032 3220 2034 3237
rect 2248 3220 2250 3237
rect 2456 3220 2458 3237
rect 2656 3220 2658 3237
rect 2840 3220 2842 3237
rect 3024 3220 3026 3237
rect 3208 3220 3210 3237
rect 3368 3220 3370 3237
rect 3464 3221 3466 3237
rect 3462 3220 3468 3221
rect 111 3218 115 3219
rect 111 3213 115 3214
rect 303 3218 307 3219
rect 303 3213 307 3214
rect 383 3218 387 3219
rect 383 3213 387 3214
rect 423 3218 427 3219
rect 423 3213 427 3214
rect 495 3218 499 3219
rect 495 3213 499 3214
rect 543 3218 547 3219
rect 543 3213 547 3214
rect 607 3218 611 3219
rect 607 3213 611 3214
rect 671 3218 675 3219
rect 671 3213 675 3214
rect 727 3218 731 3219
rect 727 3213 731 3214
rect 799 3218 803 3219
rect 799 3213 803 3214
rect 847 3218 851 3219
rect 847 3213 851 3214
rect 927 3218 931 3219
rect 927 3213 931 3214
rect 967 3218 971 3219
rect 967 3213 971 3214
rect 1055 3218 1059 3219
rect 1055 3213 1059 3214
rect 1087 3218 1091 3219
rect 1087 3213 1091 3214
rect 1175 3218 1179 3219
rect 1175 3213 1179 3214
rect 1207 3218 1211 3219
rect 1207 3213 1211 3214
rect 1303 3218 1307 3219
rect 1303 3213 1307 3214
rect 1335 3218 1339 3219
rect 1335 3213 1339 3214
rect 1431 3218 1435 3219
rect 1431 3213 1435 3214
rect 1767 3218 1771 3219
rect 1806 3216 1807 3220
rect 1811 3216 1812 3220
rect 1806 3215 1812 3216
rect 1830 3219 1836 3220
rect 1830 3215 1831 3219
rect 1835 3215 1836 3219
rect 1830 3214 1836 3215
rect 2030 3219 2036 3220
rect 2030 3215 2031 3219
rect 2035 3215 2036 3219
rect 2030 3214 2036 3215
rect 2246 3219 2252 3220
rect 2246 3215 2247 3219
rect 2251 3215 2252 3219
rect 2246 3214 2252 3215
rect 2454 3219 2460 3220
rect 2454 3215 2455 3219
rect 2459 3215 2460 3219
rect 2454 3214 2460 3215
rect 2654 3219 2660 3220
rect 2654 3215 2655 3219
rect 2659 3215 2660 3219
rect 2654 3214 2660 3215
rect 2838 3219 2844 3220
rect 2838 3215 2839 3219
rect 2843 3215 2844 3219
rect 2838 3214 2844 3215
rect 3022 3219 3028 3220
rect 3022 3215 3023 3219
rect 3027 3215 3028 3219
rect 3022 3214 3028 3215
rect 3206 3219 3212 3220
rect 3206 3215 3207 3219
rect 3211 3215 3212 3219
rect 3206 3214 3212 3215
rect 3366 3219 3372 3220
rect 3366 3215 3367 3219
rect 3371 3215 3372 3219
rect 3462 3216 3463 3220
rect 3467 3216 3468 3220
rect 3462 3215 3468 3216
rect 3366 3214 3372 3215
rect 1767 3213 1771 3214
rect 112 3197 114 3213
rect 110 3196 116 3197
rect 304 3196 306 3213
rect 424 3196 426 3213
rect 544 3196 546 3213
rect 672 3196 674 3213
rect 800 3196 802 3213
rect 928 3196 930 3213
rect 1056 3196 1058 3213
rect 1176 3196 1178 3213
rect 1304 3196 1306 3213
rect 1432 3196 1434 3213
rect 1768 3197 1770 3213
rect 1806 3203 1812 3204
rect 1806 3199 1807 3203
rect 1811 3199 1812 3203
rect 3462 3203 3468 3204
rect 1806 3198 1812 3199
rect 1830 3200 1836 3201
rect 1766 3196 1772 3197
rect 110 3192 111 3196
rect 115 3192 116 3196
rect 110 3191 116 3192
rect 302 3195 308 3196
rect 302 3191 303 3195
rect 307 3191 308 3195
rect 302 3190 308 3191
rect 422 3195 428 3196
rect 422 3191 423 3195
rect 427 3191 428 3195
rect 422 3190 428 3191
rect 542 3195 548 3196
rect 542 3191 543 3195
rect 547 3191 548 3195
rect 542 3190 548 3191
rect 670 3195 676 3196
rect 670 3191 671 3195
rect 675 3191 676 3195
rect 670 3190 676 3191
rect 798 3195 804 3196
rect 798 3191 799 3195
rect 803 3191 804 3195
rect 798 3190 804 3191
rect 926 3195 932 3196
rect 926 3191 927 3195
rect 931 3191 932 3195
rect 926 3190 932 3191
rect 1054 3195 1060 3196
rect 1054 3191 1055 3195
rect 1059 3191 1060 3195
rect 1054 3190 1060 3191
rect 1174 3195 1180 3196
rect 1174 3191 1175 3195
rect 1179 3191 1180 3195
rect 1174 3190 1180 3191
rect 1302 3195 1308 3196
rect 1302 3191 1303 3195
rect 1307 3191 1308 3195
rect 1302 3190 1308 3191
rect 1430 3195 1436 3196
rect 1430 3191 1431 3195
rect 1435 3191 1436 3195
rect 1766 3192 1767 3196
rect 1771 3192 1772 3196
rect 1766 3191 1772 3192
rect 1430 3190 1436 3191
rect 110 3179 116 3180
rect 110 3175 111 3179
rect 115 3175 116 3179
rect 1766 3179 1772 3180
rect 1808 3179 1810 3198
rect 1830 3196 1831 3200
rect 1835 3196 1836 3200
rect 1830 3195 1836 3196
rect 2030 3200 2036 3201
rect 2030 3196 2031 3200
rect 2035 3196 2036 3200
rect 2030 3195 2036 3196
rect 2246 3200 2252 3201
rect 2246 3196 2247 3200
rect 2251 3196 2252 3200
rect 2246 3195 2252 3196
rect 2454 3200 2460 3201
rect 2454 3196 2455 3200
rect 2459 3196 2460 3200
rect 2454 3195 2460 3196
rect 2654 3200 2660 3201
rect 2654 3196 2655 3200
rect 2659 3196 2660 3200
rect 2654 3195 2660 3196
rect 2838 3200 2844 3201
rect 2838 3196 2839 3200
rect 2843 3196 2844 3200
rect 2838 3195 2844 3196
rect 3022 3200 3028 3201
rect 3022 3196 3023 3200
rect 3027 3196 3028 3200
rect 3022 3195 3028 3196
rect 3206 3200 3212 3201
rect 3206 3196 3207 3200
rect 3211 3196 3212 3200
rect 3206 3195 3212 3196
rect 3366 3200 3372 3201
rect 3366 3196 3367 3200
rect 3371 3196 3372 3200
rect 3462 3199 3463 3203
rect 3467 3199 3468 3203
rect 3462 3198 3468 3199
rect 3366 3195 3372 3196
rect 1832 3179 1834 3195
rect 2032 3179 2034 3195
rect 2248 3179 2250 3195
rect 2456 3179 2458 3195
rect 2656 3179 2658 3195
rect 2840 3179 2842 3195
rect 3024 3179 3026 3195
rect 3208 3179 3210 3195
rect 3368 3179 3370 3195
rect 3464 3179 3466 3198
rect 110 3174 116 3175
rect 302 3176 308 3177
rect 112 3143 114 3174
rect 302 3172 303 3176
rect 307 3172 308 3176
rect 302 3171 308 3172
rect 422 3176 428 3177
rect 422 3172 423 3176
rect 427 3172 428 3176
rect 422 3171 428 3172
rect 542 3176 548 3177
rect 542 3172 543 3176
rect 547 3172 548 3176
rect 542 3171 548 3172
rect 670 3176 676 3177
rect 670 3172 671 3176
rect 675 3172 676 3176
rect 670 3171 676 3172
rect 798 3176 804 3177
rect 798 3172 799 3176
rect 803 3172 804 3176
rect 798 3171 804 3172
rect 926 3176 932 3177
rect 926 3172 927 3176
rect 931 3172 932 3176
rect 926 3171 932 3172
rect 1054 3176 1060 3177
rect 1054 3172 1055 3176
rect 1059 3172 1060 3176
rect 1054 3171 1060 3172
rect 1174 3176 1180 3177
rect 1174 3172 1175 3176
rect 1179 3172 1180 3176
rect 1174 3171 1180 3172
rect 1302 3176 1308 3177
rect 1302 3172 1303 3176
rect 1307 3172 1308 3176
rect 1302 3171 1308 3172
rect 1430 3176 1436 3177
rect 1430 3172 1431 3176
rect 1435 3172 1436 3176
rect 1766 3175 1767 3179
rect 1771 3175 1772 3179
rect 1766 3174 1772 3175
rect 1807 3178 1811 3179
rect 1430 3171 1436 3172
rect 304 3143 306 3171
rect 424 3143 426 3171
rect 544 3143 546 3171
rect 672 3143 674 3171
rect 800 3143 802 3171
rect 928 3143 930 3171
rect 1056 3143 1058 3171
rect 1176 3143 1178 3171
rect 1304 3143 1306 3171
rect 1432 3143 1434 3171
rect 1768 3143 1770 3174
rect 1807 3173 1811 3174
rect 1831 3178 1835 3179
rect 1831 3173 1835 3174
rect 1839 3178 1843 3179
rect 1839 3173 1843 3174
rect 2031 3178 2035 3179
rect 2031 3173 2035 3174
rect 2223 3178 2227 3179
rect 2223 3173 2227 3174
rect 2247 3178 2251 3179
rect 2247 3173 2251 3174
rect 2407 3178 2411 3179
rect 2407 3173 2411 3174
rect 2455 3178 2459 3179
rect 2455 3173 2459 3174
rect 2575 3178 2579 3179
rect 2575 3173 2579 3174
rect 2655 3178 2659 3179
rect 2655 3173 2659 3174
rect 2735 3178 2739 3179
rect 2735 3173 2739 3174
rect 2839 3178 2843 3179
rect 2839 3173 2843 3174
rect 2879 3178 2883 3179
rect 2879 3173 2883 3174
rect 3007 3178 3011 3179
rect 3007 3173 3011 3174
rect 3023 3178 3027 3179
rect 3023 3173 3027 3174
rect 3135 3178 3139 3179
rect 3135 3173 3139 3174
rect 3207 3178 3211 3179
rect 3207 3173 3211 3174
rect 3263 3178 3267 3179
rect 3263 3173 3267 3174
rect 3367 3178 3371 3179
rect 3367 3173 3371 3174
rect 3463 3178 3467 3179
rect 3463 3173 3467 3174
rect 1808 3154 1810 3173
rect 1840 3157 1842 3173
rect 2032 3157 2034 3173
rect 2224 3157 2226 3173
rect 2408 3157 2410 3173
rect 2576 3157 2578 3173
rect 2736 3157 2738 3173
rect 2880 3157 2882 3173
rect 3008 3157 3010 3173
rect 3136 3157 3138 3173
rect 3264 3157 3266 3173
rect 3368 3157 3370 3173
rect 1838 3156 1844 3157
rect 1806 3153 1812 3154
rect 1806 3149 1807 3153
rect 1811 3149 1812 3153
rect 1838 3152 1839 3156
rect 1843 3152 1844 3156
rect 1838 3151 1844 3152
rect 2030 3156 2036 3157
rect 2030 3152 2031 3156
rect 2035 3152 2036 3156
rect 2030 3151 2036 3152
rect 2222 3156 2228 3157
rect 2222 3152 2223 3156
rect 2227 3152 2228 3156
rect 2222 3151 2228 3152
rect 2406 3156 2412 3157
rect 2406 3152 2407 3156
rect 2411 3152 2412 3156
rect 2406 3151 2412 3152
rect 2574 3156 2580 3157
rect 2574 3152 2575 3156
rect 2579 3152 2580 3156
rect 2574 3151 2580 3152
rect 2734 3156 2740 3157
rect 2734 3152 2735 3156
rect 2739 3152 2740 3156
rect 2734 3151 2740 3152
rect 2878 3156 2884 3157
rect 2878 3152 2879 3156
rect 2883 3152 2884 3156
rect 2878 3151 2884 3152
rect 3006 3156 3012 3157
rect 3006 3152 3007 3156
rect 3011 3152 3012 3156
rect 3006 3151 3012 3152
rect 3134 3156 3140 3157
rect 3134 3152 3135 3156
rect 3139 3152 3140 3156
rect 3134 3151 3140 3152
rect 3262 3156 3268 3157
rect 3262 3152 3263 3156
rect 3267 3152 3268 3156
rect 3262 3151 3268 3152
rect 3366 3156 3372 3157
rect 3366 3152 3367 3156
rect 3371 3152 3372 3156
rect 3464 3154 3466 3173
rect 3366 3151 3372 3152
rect 3462 3153 3468 3154
rect 1806 3148 1812 3149
rect 3462 3149 3463 3153
rect 3467 3149 3468 3153
rect 3462 3148 3468 3149
rect 111 3142 115 3143
rect 111 3137 115 3138
rect 175 3142 179 3143
rect 175 3137 179 3138
rect 303 3142 307 3143
rect 303 3137 307 3138
rect 319 3142 323 3143
rect 319 3137 323 3138
rect 423 3142 427 3143
rect 423 3137 427 3138
rect 471 3142 475 3143
rect 471 3137 475 3138
rect 543 3142 547 3143
rect 543 3137 547 3138
rect 623 3142 627 3143
rect 623 3137 627 3138
rect 671 3142 675 3143
rect 671 3137 675 3138
rect 775 3142 779 3143
rect 775 3137 779 3138
rect 799 3142 803 3143
rect 799 3137 803 3138
rect 919 3142 923 3143
rect 919 3137 923 3138
rect 927 3142 931 3143
rect 927 3137 931 3138
rect 1055 3142 1059 3143
rect 1055 3137 1059 3138
rect 1063 3142 1067 3143
rect 1063 3137 1067 3138
rect 1175 3142 1179 3143
rect 1175 3137 1179 3138
rect 1199 3142 1203 3143
rect 1199 3137 1203 3138
rect 1303 3142 1307 3143
rect 1303 3137 1307 3138
rect 1343 3142 1347 3143
rect 1343 3137 1347 3138
rect 1431 3142 1435 3143
rect 1431 3137 1435 3138
rect 1487 3142 1491 3143
rect 1487 3137 1491 3138
rect 1767 3142 1771 3143
rect 1767 3137 1771 3138
rect 1838 3137 1844 3138
rect 112 3118 114 3137
rect 176 3121 178 3137
rect 320 3121 322 3137
rect 472 3121 474 3137
rect 624 3121 626 3137
rect 776 3121 778 3137
rect 920 3121 922 3137
rect 1064 3121 1066 3137
rect 1200 3121 1202 3137
rect 1344 3121 1346 3137
rect 1488 3121 1490 3137
rect 174 3120 180 3121
rect 110 3117 116 3118
rect 110 3113 111 3117
rect 115 3113 116 3117
rect 174 3116 175 3120
rect 179 3116 180 3120
rect 174 3115 180 3116
rect 318 3120 324 3121
rect 318 3116 319 3120
rect 323 3116 324 3120
rect 318 3115 324 3116
rect 470 3120 476 3121
rect 470 3116 471 3120
rect 475 3116 476 3120
rect 470 3115 476 3116
rect 622 3120 628 3121
rect 622 3116 623 3120
rect 627 3116 628 3120
rect 622 3115 628 3116
rect 774 3120 780 3121
rect 774 3116 775 3120
rect 779 3116 780 3120
rect 774 3115 780 3116
rect 918 3120 924 3121
rect 918 3116 919 3120
rect 923 3116 924 3120
rect 918 3115 924 3116
rect 1062 3120 1068 3121
rect 1062 3116 1063 3120
rect 1067 3116 1068 3120
rect 1062 3115 1068 3116
rect 1198 3120 1204 3121
rect 1198 3116 1199 3120
rect 1203 3116 1204 3120
rect 1198 3115 1204 3116
rect 1342 3120 1348 3121
rect 1342 3116 1343 3120
rect 1347 3116 1348 3120
rect 1342 3115 1348 3116
rect 1486 3120 1492 3121
rect 1486 3116 1487 3120
rect 1491 3116 1492 3120
rect 1768 3118 1770 3137
rect 1806 3136 1812 3137
rect 1806 3132 1807 3136
rect 1811 3132 1812 3136
rect 1838 3133 1839 3137
rect 1843 3133 1844 3137
rect 1838 3132 1844 3133
rect 2030 3137 2036 3138
rect 2030 3133 2031 3137
rect 2035 3133 2036 3137
rect 2030 3132 2036 3133
rect 2222 3137 2228 3138
rect 2222 3133 2223 3137
rect 2227 3133 2228 3137
rect 2222 3132 2228 3133
rect 2406 3137 2412 3138
rect 2406 3133 2407 3137
rect 2411 3133 2412 3137
rect 2406 3132 2412 3133
rect 2574 3137 2580 3138
rect 2574 3133 2575 3137
rect 2579 3133 2580 3137
rect 2574 3132 2580 3133
rect 2734 3137 2740 3138
rect 2734 3133 2735 3137
rect 2739 3133 2740 3137
rect 2734 3132 2740 3133
rect 2878 3137 2884 3138
rect 2878 3133 2879 3137
rect 2883 3133 2884 3137
rect 2878 3132 2884 3133
rect 3006 3137 3012 3138
rect 3006 3133 3007 3137
rect 3011 3133 3012 3137
rect 3006 3132 3012 3133
rect 3134 3137 3140 3138
rect 3134 3133 3135 3137
rect 3139 3133 3140 3137
rect 3134 3132 3140 3133
rect 3262 3137 3268 3138
rect 3262 3133 3263 3137
rect 3267 3133 3268 3137
rect 3262 3132 3268 3133
rect 3366 3137 3372 3138
rect 3366 3133 3367 3137
rect 3371 3133 3372 3137
rect 3366 3132 3372 3133
rect 3462 3136 3468 3137
rect 3462 3132 3463 3136
rect 3467 3132 3468 3136
rect 1806 3131 1812 3132
rect 1486 3115 1492 3116
rect 1766 3117 1772 3118
rect 110 3112 116 3113
rect 1766 3113 1767 3117
rect 1771 3113 1772 3117
rect 1766 3112 1772 3113
rect 1808 3111 1810 3131
rect 1840 3111 1842 3132
rect 2032 3111 2034 3132
rect 2224 3111 2226 3132
rect 2408 3111 2410 3132
rect 2576 3111 2578 3132
rect 2736 3111 2738 3132
rect 2880 3111 2882 3132
rect 3008 3111 3010 3132
rect 3136 3111 3138 3132
rect 3264 3111 3266 3132
rect 3368 3111 3370 3132
rect 3462 3131 3468 3132
rect 3464 3111 3466 3131
rect 1807 3110 1811 3111
rect 1807 3105 1811 3106
rect 1839 3110 1843 3111
rect 1839 3105 1843 3106
rect 1935 3110 1939 3111
rect 1935 3105 1939 3106
rect 2031 3110 2035 3111
rect 2031 3105 2035 3106
rect 2055 3110 2059 3111
rect 2055 3105 2059 3106
rect 2175 3110 2179 3111
rect 2175 3105 2179 3106
rect 2223 3110 2227 3111
rect 2223 3105 2227 3106
rect 2303 3110 2307 3111
rect 2303 3105 2307 3106
rect 2407 3110 2411 3111
rect 2407 3105 2411 3106
rect 2431 3110 2435 3111
rect 2431 3105 2435 3106
rect 2567 3110 2571 3111
rect 2567 3105 2571 3106
rect 2575 3110 2579 3111
rect 2575 3105 2579 3106
rect 2719 3110 2723 3111
rect 2719 3105 2723 3106
rect 2735 3110 2739 3111
rect 2735 3105 2739 3106
rect 2871 3110 2875 3111
rect 2871 3105 2875 3106
rect 2879 3110 2883 3111
rect 2879 3105 2883 3106
rect 3007 3110 3011 3111
rect 3007 3105 3011 3106
rect 3031 3110 3035 3111
rect 3031 3105 3035 3106
rect 3135 3110 3139 3111
rect 3135 3105 3139 3106
rect 3199 3110 3203 3111
rect 3199 3105 3203 3106
rect 3263 3110 3267 3111
rect 3263 3105 3267 3106
rect 3367 3110 3371 3111
rect 3367 3105 3371 3106
rect 3463 3110 3467 3111
rect 3463 3105 3467 3106
rect 174 3101 180 3102
rect 110 3100 116 3101
rect 110 3096 111 3100
rect 115 3096 116 3100
rect 174 3097 175 3101
rect 179 3097 180 3101
rect 174 3096 180 3097
rect 318 3101 324 3102
rect 318 3097 319 3101
rect 323 3097 324 3101
rect 318 3096 324 3097
rect 470 3101 476 3102
rect 470 3097 471 3101
rect 475 3097 476 3101
rect 470 3096 476 3097
rect 622 3101 628 3102
rect 622 3097 623 3101
rect 627 3097 628 3101
rect 622 3096 628 3097
rect 774 3101 780 3102
rect 774 3097 775 3101
rect 779 3097 780 3101
rect 774 3096 780 3097
rect 918 3101 924 3102
rect 918 3097 919 3101
rect 923 3097 924 3101
rect 918 3096 924 3097
rect 1062 3101 1068 3102
rect 1062 3097 1063 3101
rect 1067 3097 1068 3101
rect 1062 3096 1068 3097
rect 1198 3101 1204 3102
rect 1198 3097 1199 3101
rect 1203 3097 1204 3101
rect 1198 3096 1204 3097
rect 1342 3101 1348 3102
rect 1342 3097 1343 3101
rect 1347 3097 1348 3101
rect 1342 3096 1348 3097
rect 1486 3101 1492 3102
rect 1486 3097 1487 3101
rect 1491 3097 1492 3101
rect 1486 3096 1492 3097
rect 1766 3100 1772 3101
rect 1766 3096 1767 3100
rect 1771 3096 1772 3100
rect 110 3095 116 3096
rect 112 3071 114 3095
rect 176 3071 178 3096
rect 320 3071 322 3096
rect 472 3071 474 3096
rect 624 3071 626 3096
rect 776 3071 778 3096
rect 920 3071 922 3096
rect 1064 3071 1066 3096
rect 1200 3071 1202 3096
rect 1344 3071 1346 3096
rect 1488 3071 1490 3096
rect 1766 3095 1772 3096
rect 1768 3071 1770 3095
rect 1808 3089 1810 3105
rect 1806 3088 1812 3089
rect 1936 3088 1938 3105
rect 2056 3088 2058 3105
rect 2176 3088 2178 3105
rect 2304 3088 2306 3105
rect 2432 3088 2434 3105
rect 2568 3088 2570 3105
rect 2720 3088 2722 3105
rect 2872 3088 2874 3105
rect 3032 3088 3034 3105
rect 3200 3088 3202 3105
rect 3368 3088 3370 3105
rect 3464 3089 3466 3105
rect 3462 3088 3468 3089
rect 1806 3084 1807 3088
rect 1811 3084 1812 3088
rect 1806 3083 1812 3084
rect 1934 3087 1940 3088
rect 1934 3083 1935 3087
rect 1939 3083 1940 3087
rect 1934 3082 1940 3083
rect 2054 3087 2060 3088
rect 2054 3083 2055 3087
rect 2059 3083 2060 3087
rect 2054 3082 2060 3083
rect 2174 3087 2180 3088
rect 2174 3083 2175 3087
rect 2179 3083 2180 3087
rect 2174 3082 2180 3083
rect 2302 3087 2308 3088
rect 2302 3083 2303 3087
rect 2307 3083 2308 3087
rect 2302 3082 2308 3083
rect 2430 3087 2436 3088
rect 2430 3083 2431 3087
rect 2435 3083 2436 3087
rect 2430 3082 2436 3083
rect 2566 3087 2572 3088
rect 2566 3083 2567 3087
rect 2571 3083 2572 3087
rect 2566 3082 2572 3083
rect 2718 3087 2724 3088
rect 2718 3083 2719 3087
rect 2723 3083 2724 3087
rect 2718 3082 2724 3083
rect 2870 3087 2876 3088
rect 2870 3083 2871 3087
rect 2875 3083 2876 3087
rect 2870 3082 2876 3083
rect 3030 3087 3036 3088
rect 3030 3083 3031 3087
rect 3035 3083 3036 3087
rect 3030 3082 3036 3083
rect 3198 3087 3204 3088
rect 3198 3083 3199 3087
rect 3203 3083 3204 3087
rect 3198 3082 3204 3083
rect 3366 3087 3372 3088
rect 3366 3083 3367 3087
rect 3371 3083 3372 3087
rect 3462 3084 3463 3088
rect 3467 3084 3468 3088
rect 3462 3083 3468 3084
rect 3366 3082 3372 3083
rect 1806 3071 1812 3072
rect 111 3070 115 3071
rect 111 3065 115 3066
rect 135 3070 139 3071
rect 135 3065 139 3066
rect 175 3070 179 3071
rect 175 3065 179 3066
rect 263 3070 267 3071
rect 263 3065 267 3066
rect 319 3070 323 3071
rect 319 3065 323 3066
rect 431 3070 435 3071
rect 431 3065 435 3066
rect 471 3070 475 3071
rect 471 3065 475 3066
rect 607 3070 611 3071
rect 607 3065 611 3066
rect 623 3070 627 3071
rect 623 3065 627 3066
rect 775 3070 779 3071
rect 775 3065 779 3066
rect 791 3070 795 3071
rect 791 3065 795 3066
rect 919 3070 923 3071
rect 919 3065 923 3066
rect 967 3070 971 3071
rect 967 3065 971 3066
rect 1063 3070 1067 3071
rect 1063 3065 1067 3066
rect 1143 3070 1147 3071
rect 1143 3065 1147 3066
rect 1199 3070 1203 3071
rect 1199 3065 1203 3066
rect 1327 3070 1331 3071
rect 1327 3065 1331 3066
rect 1343 3070 1347 3071
rect 1343 3065 1347 3066
rect 1487 3070 1491 3071
rect 1487 3065 1491 3066
rect 1511 3070 1515 3071
rect 1511 3065 1515 3066
rect 1767 3070 1771 3071
rect 1806 3067 1807 3071
rect 1811 3067 1812 3071
rect 3462 3071 3468 3072
rect 1806 3066 1812 3067
rect 1934 3068 1940 3069
rect 1767 3065 1771 3066
rect 112 3049 114 3065
rect 110 3048 116 3049
rect 136 3048 138 3065
rect 264 3048 266 3065
rect 432 3048 434 3065
rect 608 3048 610 3065
rect 792 3048 794 3065
rect 968 3048 970 3065
rect 1144 3048 1146 3065
rect 1328 3048 1330 3065
rect 1512 3048 1514 3065
rect 1768 3049 1770 3065
rect 1766 3048 1772 3049
rect 110 3044 111 3048
rect 115 3044 116 3048
rect 110 3043 116 3044
rect 134 3047 140 3048
rect 134 3043 135 3047
rect 139 3043 140 3047
rect 134 3042 140 3043
rect 262 3047 268 3048
rect 262 3043 263 3047
rect 267 3043 268 3047
rect 262 3042 268 3043
rect 430 3047 436 3048
rect 430 3043 431 3047
rect 435 3043 436 3047
rect 430 3042 436 3043
rect 606 3047 612 3048
rect 606 3043 607 3047
rect 611 3043 612 3047
rect 606 3042 612 3043
rect 790 3047 796 3048
rect 790 3043 791 3047
rect 795 3043 796 3047
rect 790 3042 796 3043
rect 966 3047 972 3048
rect 966 3043 967 3047
rect 971 3043 972 3047
rect 966 3042 972 3043
rect 1142 3047 1148 3048
rect 1142 3043 1143 3047
rect 1147 3043 1148 3047
rect 1142 3042 1148 3043
rect 1326 3047 1332 3048
rect 1326 3043 1327 3047
rect 1331 3043 1332 3047
rect 1326 3042 1332 3043
rect 1510 3047 1516 3048
rect 1510 3043 1511 3047
rect 1515 3043 1516 3047
rect 1766 3044 1767 3048
rect 1771 3044 1772 3048
rect 1766 3043 1772 3044
rect 1510 3042 1516 3043
rect 1808 3039 1810 3066
rect 1934 3064 1935 3068
rect 1939 3064 1940 3068
rect 1934 3063 1940 3064
rect 2054 3068 2060 3069
rect 2054 3064 2055 3068
rect 2059 3064 2060 3068
rect 2054 3063 2060 3064
rect 2174 3068 2180 3069
rect 2174 3064 2175 3068
rect 2179 3064 2180 3068
rect 2174 3063 2180 3064
rect 2302 3068 2308 3069
rect 2302 3064 2303 3068
rect 2307 3064 2308 3068
rect 2302 3063 2308 3064
rect 2430 3068 2436 3069
rect 2430 3064 2431 3068
rect 2435 3064 2436 3068
rect 2430 3063 2436 3064
rect 2566 3068 2572 3069
rect 2566 3064 2567 3068
rect 2571 3064 2572 3068
rect 2566 3063 2572 3064
rect 2718 3068 2724 3069
rect 2718 3064 2719 3068
rect 2723 3064 2724 3068
rect 2718 3063 2724 3064
rect 2870 3068 2876 3069
rect 2870 3064 2871 3068
rect 2875 3064 2876 3068
rect 2870 3063 2876 3064
rect 3030 3068 3036 3069
rect 3030 3064 3031 3068
rect 3035 3064 3036 3068
rect 3030 3063 3036 3064
rect 3198 3068 3204 3069
rect 3198 3064 3199 3068
rect 3203 3064 3204 3068
rect 3198 3063 3204 3064
rect 3366 3068 3372 3069
rect 3366 3064 3367 3068
rect 3371 3064 3372 3068
rect 3462 3067 3463 3071
rect 3467 3067 3468 3071
rect 3462 3066 3468 3067
rect 3366 3063 3372 3064
rect 1936 3039 1938 3063
rect 2056 3039 2058 3063
rect 2176 3039 2178 3063
rect 2304 3039 2306 3063
rect 2432 3039 2434 3063
rect 2568 3039 2570 3063
rect 2720 3039 2722 3063
rect 2872 3039 2874 3063
rect 3032 3039 3034 3063
rect 3200 3039 3202 3063
rect 3368 3039 3370 3063
rect 3464 3039 3466 3066
rect 1807 3038 1811 3039
rect 1807 3033 1811 3034
rect 1935 3038 1939 3039
rect 1935 3033 1939 3034
rect 2023 3038 2027 3039
rect 2023 3033 2027 3034
rect 2055 3038 2059 3039
rect 2055 3033 2059 3034
rect 2127 3038 2131 3039
rect 2127 3033 2131 3034
rect 2175 3038 2179 3039
rect 2175 3033 2179 3034
rect 2231 3038 2235 3039
rect 2231 3033 2235 3034
rect 2303 3038 2307 3039
rect 2303 3033 2307 3034
rect 2335 3038 2339 3039
rect 2335 3033 2339 3034
rect 2431 3038 2435 3039
rect 2431 3033 2435 3034
rect 2439 3038 2443 3039
rect 2439 3033 2443 3034
rect 2543 3038 2547 3039
rect 2543 3033 2547 3034
rect 2567 3038 2571 3039
rect 2567 3033 2571 3034
rect 2647 3038 2651 3039
rect 2647 3033 2651 3034
rect 2719 3038 2723 3039
rect 2719 3033 2723 3034
rect 2759 3038 2763 3039
rect 2759 3033 2763 3034
rect 2871 3038 2875 3039
rect 2871 3033 2875 3034
rect 3031 3038 3035 3039
rect 3031 3033 3035 3034
rect 3199 3038 3203 3039
rect 3199 3033 3203 3034
rect 3367 3038 3371 3039
rect 3367 3033 3371 3034
rect 3463 3038 3467 3039
rect 3463 3033 3467 3034
rect 110 3031 116 3032
rect 110 3027 111 3031
rect 115 3027 116 3031
rect 1766 3031 1772 3032
rect 110 3026 116 3027
rect 134 3028 140 3029
rect 112 3003 114 3026
rect 134 3024 135 3028
rect 139 3024 140 3028
rect 134 3023 140 3024
rect 262 3028 268 3029
rect 262 3024 263 3028
rect 267 3024 268 3028
rect 262 3023 268 3024
rect 430 3028 436 3029
rect 430 3024 431 3028
rect 435 3024 436 3028
rect 430 3023 436 3024
rect 606 3028 612 3029
rect 606 3024 607 3028
rect 611 3024 612 3028
rect 606 3023 612 3024
rect 790 3028 796 3029
rect 790 3024 791 3028
rect 795 3024 796 3028
rect 790 3023 796 3024
rect 966 3028 972 3029
rect 966 3024 967 3028
rect 971 3024 972 3028
rect 966 3023 972 3024
rect 1142 3028 1148 3029
rect 1142 3024 1143 3028
rect 1147 3024 1148 3028
rect 1142 3023 1148 3024
rect 1326 3028 1332 3029
rect 1326 3024 1327 3028
rect 1331 3024 1332 3028
rect 1326 3023 1332 3024
rect 1510 3028 1516 3029
rect 1510 3024 1511 3028
rect 1515 3024 1516 3028
rect 1766 3027 1767 3031
rect 1771 3027 1772 3031
rect 1766 3026 1772 3027
rect 1510 3023 1516 3024
rect 136 3003 138 3023
rect 264 3003 266 3023
rect 432 3003 434 3023
rect 608 3003 610 3023
rect 792 3003 794 3023
rect 968 3003 970 3023
rect 1144 3003 1146 3023
rect 1328 3003 1330 3023
rect 1512 3003 1514 3023
rect 1768 3003 1770 3026
rect 1808 3014 1810 3033
rect 2024 3017 2026 3033
rect 2128 3017 2130 3033
rect 2232 3017 2234 3033
rect 2336 3017 2338 3033
rect 2440 3017 2442 3033
rect 2544 3017 2546 3033
rect 2648 3017 2650 3033
rect 2760 3017 2762 3033
rect 2022 3016 2028 3017
rect 1806 3013 1812 3014
rect 1806 3009 1807 3013
rect 1811 3009 1812 3013
rect 2022 3012 2023 3016
rect 2027 3012 2028 3016
rect 2022 3011 2028 3012
rect 2126 3016 2132 3017
rect 2126 3012 2127 3016
rect 2131 3012 2132 3016
rect 2126 3011 2132 3012
rect 2230 3016 2236 3017
rect 2230 3012 2231 3016
rect 2235 3012 2236 3016
rect 2230 3011 2236 3012
rect 2334 3016 2340 3017
rect 2334 3012 2335 3016
rect 2339 3012 2340 3016
rect 2334 3011 2340 3012
rect 2438 3016 2444 3017
rect 2438 3012 2439 3016
rect 2443 3012 2444 3016
rect 2438 3011 2444 3012
rect 2542 3016 2548 3017
rect 2542 3012 2543 3016
rect 2547 3012 2548 3016
rect 2542 3011 2548 3012
rect 2646 3016 2652 3017
rect 2646 3012 2647 3016
rect 2651 3012 2652 3016
rect 2646 3011 2652 3012
rect 2758 3016 2764 3017
rect 2758 3012 2759 3016
rect 2763 3012 2764 3016
rect 3464 3014 3466 3033
rect 2758 3011 2764 3012
rect 3462 3013 3468 3014
rect 1806 3008 1812 3009
rect 3462 3009 3463 3013
rect 3467 3009 3468 3013
rect 3462 3008 3468 3009
rect 111 3002 115 3003
rect 111 2997 115 2998
rect 135 3002 139 3003
rect 135 2997 139 2998
rect 263 3002 267 3003
rect 263 2997 267 2998
rect 327 3002 331 3003
rect 327 2997 331 2998
rect 431 3002 435 3003
rect 431 2997 435 2998
rect 535 3002 539 3003
rect 535 2997 539 2998
rect 607 3002 611 3003
rect 607 2997 611 2998
rect 735 3002 739 3003
rect 735 2997 739 2998
rect 791 3002 795 3003
rect 791 2997 795 2998
rect 927 3002 931 3003
rect 927 2997 931 2998
rect 967 3002 971 3003
rect 967 2997 971 2998
rect 1103 3002 1107 3003
rect 1103 2997 1107 2998
rect 1143 3002 1147 3003
rect 1143 2997 1147 2998
rect 1279 3002 1283 3003
rect 1279 2997 1283 2998
rect 1327 3002 1331 3003
rect 1327 2997 1331 2998
rect 1447 3002 1451 3003
rect 1447 2997 1451 2998
rect 1511 3002 1515 3003
rect 1511 2997 1515 2998
rect 1623 3002 1627 3003
rect 1623 2997 1627 2998
rect 1767 3002 1771 3003
rect 1767 2997 1771 2998
rect 2022 2997 2028 2998
rect 112 2978 114 2997
rect 136 2981 138 2997
rect 328 2981 330 2997
rect 536 2981 538 2997
rect 736 2981 738 2997
rect 928 2981 930 2997
rect 1104 2981 1106 2997
rect 1280 2981 1282 2997
rect 1448 2981 1450 2997
rect 1624 2981 1626 2997
rect 134 2980 140 2981
rect 110 2977 116 2978
rect 110 2973 111 2977
rect 115 2973 116 2977
rect 134 2976 135 2980
rect 139 2976 140 2980
rect 134 2975 140 2976
rect 326 2980 332 2981
rect 326 2976 327 2980
rect 331 2976 332 2980
rect 326 2975 332 2976
rect 534 2980 540 2981
rect 534 2976 535 2980
rect 539 2976 540 2980
rect 534 2975 540 2976
rect 734 2980 740 2981
rect 734 2976 735 2980
rect 739 2976 740 2980
rect 734 2975 740 2976
rect 926 2980 932 2981
rect 926 2976 927 2980
rect 931 2976 932 2980
rect 926 2975 932 2976
rect 1102 2980 1108 2981
rect 1102 2976 1103 2980
rect 1107 2976 1108 2980
rect 1102 2975 1108 2976
rect 1278 2980 1284 2981
rect 1278 2976 1279 2980
rect 1283 2976 1284 2980
rect 1278 2975 1284 2976
rect 1446 2980 1452 2981
rect 1446 2976 1447 2980
rect 1451 2976 1452 2980
rect 1446 2975 1452 2976
rect 1622 2980 1628 2981
rect 1622 2976 1623 2980
rect 1627 2976 1628 2980
rect 1768 2978 1770 2997
rect 1806 2996 1812 2997
rect 1806 2992 1807 2996
rect 1811 2992 1812 2996
rect 2022 2993 2023 2997
rect 2027 2993 2028 2997
rect 2022 2992 2028 2993
rect 2126 2997 2132 2998
rect 2126 2993 2127 2997
rect 2131 2993 2132 2997
rect 2126 2992 2132 2993
rect 2230 2997 2236 2998
rect 2230 2993 2231 2997
rect 2235 2993 2236 2997
rect 2230 2992 2236 2993
rect 2334 2997 2340 2998
rect 2334 2993 2335 2997
rect 2339 2993 2340 2997
rect 2334 2992 2340 2993
rect 2438 2997 2444 2998
rect 2438 2993 2439 2997
rect 2443 2993 2444 2997
rect 2438 2992 2444 2993
rect 2542 2997 2548 2998
rect 2542 2993 2543 2997
rect 2547 2993 2548 2997
rect 2542 2992 2548 2993
rect 2646 2997 2652 2998
rect 2646 2993 2647 2997
rect 2651 2993 2652 2997
rect 2646 2992 2652 2993
rect 2758 2997 2764 2998
rect 2758 2993 2759 2997
rect 2763 2993 2764 2997
rect 2758 2992 2764 2993
rect 3462 2996 3468 2997
rect 3462 2992 3463 2996
rect 3467 2992 3468 2996
rect 1806 2991 1812 2992
rect 1622 2975 1628 2976
rect 1766 2977 1772 2978
rect 110 2972 116 2973
rect 1766 2973 1767 2977
rect 1771 2973 1772 2977
rect 1808 2975 1810 2991
rect 2024 2975 2026 2992
rect 2128 2975 2130 2992
rect 2232 2975 2234 2992
rect 2336 2975 2338 2992
rect 2440 2975 2442 2992
rect 2544 2975 2546 2992
rect 2648 2975 2650 2992
rect 2760 2975 2762 2992
rect 3462 2991 3468 2992
rect 3464 2975 3466 2991
rect 1766 2972 1772 2973
rect 1807 2974 1811 2975
rect 1807 2969 1811 2970
rect 2023 2974 2027 2975
rect 2023 2969 2027 2970
rect 2055 2974 2059 2975
rect 2055 2969 2059 2970
rect 2127 2974 2131 2975
rect 2127 2969 2131 2970
rect 2143 2974 2147 2975
rect 2143 2969 2147 2970
rect 2231 2974 2235 2975
rect 2231 2969 2235 2970
rect 2319 2974 2323 2975
rect 2319 2969 2323 2970
rect 2335 2974 2339 2975
rect 2335 2969 2339 2970
rect 2407 2974 2411 2975
rect 2407 2969 2411 2970
rect 2439 2974 2443 2975
rect 2439 2969 2443 2970
rect 2495 2974 2499 2975
rect 2495 2969 2499 2970
rect 2543 2974 2547 2975
rect 2543 2969 2547 2970
rect 2583 2974 2587 2975
rect 2583 2969 2587 2970
rect 2647 2974 2651 2975
rect 2647 2969 2651 2970
rect 2671 2974 2675 2975
rect 2671 2969 2675 2970
rect 2759 2974 2763 2975
rect 2759 2969 2763 2970
rect 2847 2974 2851 2975
rect 2847 2969 2851 2970
rect 3463 2974 3467 2975
rect 3463 2969 3467 2970
rect 134 2961 140 2962
rect 110 2960 116 2961
rect 110 2956 111 2960
rect 115 2956 116 2960
rect 134 2957 135 2961
rect 139 2957 140 2961
rect 134 2956 140 2957
rect 326 2961 332 2962
rect 326 2957 327 2961
rect 331 2957 332 2961
rect 326 2956 332 2957
rect 534 2961 540 2962
rect 534 2957 535 2961
rect 539 2957 540 2961
rect 534 2956 540 2957
rect 734 2961 740 2962
rect 734 2957 735 2961
rect 739 2957 740 2961
rect 734 2956 740 2957
rect 926 2961 932 2962
rect 926 2957 927 2961
rect 931 2957 932 2961
rect 926 2956 932 2957
rect 1102 2961 1108 2962
rect 1102 2957 1103 2961
rect 1107 2957 1108 2961
rect 1102 2956 1108 2957
rect 1278 2961 1284 2962
rect 1278 2957 1279 2961
rect 1283 2957 1284 2961
rect 1278 2956 1284 2957
rect 1446 2961 1452 2962
rect 1446 2957 1447 2961
rect 1451 2957 1452 2961
rect 1446 2956 1452 2957
rect 1622 2961 1628 2962
rect 1622 2957 1623 2961
rect 1627 2957 1628 2961
rect 1622 2956 1628 2957
rect 1766 2960 1772 2961
rect 1766 2956 1767 2960
rect 1771 2956 1772 2960
rect 110 2955 116 2956
rect 112 2931 114 2955
rect 136 2931 138 2956
rect 328 2931 330 2956
rect 536 2931 538 2956
rect 736 2931 738 2956
rect 928 2931 930 2956
rect 1104 2931 1106 2956
rect 1280 2931 1282 2956
rect 1448 2931 1450 2956
rect 1624 2931 1626 2956
rect 1766 2955 1772 2956
rect 1768 2931 1770 2955
rect 1808 2953 1810 2969
rect 1806 2952 1812 2953
rect 2056 2952 2058 2969
rect 2144 2952 2146 2969
rect 2232 2952 2234 2969
rect 2320 2952 2322 2969
rect 2408 2952 2410 2969
rect 2496 2952 2498 2969
rect 2584 2952 2586 2969
rect 2672 2952 2674 2969
rect 2760 2952 2762 2969
rect 2848 2952 2850 2969
rect 3464 2953 3466 2969
rect 3462 2952 3468 2953
rect 1806 2948 1807 2952
rect 1811 2948 1812 2952
rect 1806 2947 1812 2948
rect 2054 2951 2060 2952
rect 2054 2947 2055 2951
rect 2059 2947 2060 2951
rect 2054 2946 2060 2947
rect 2142 2951 2148 2952
rect 2142 2947 2143 2951
rect 2147 2947 2148 2951
rect 2142 2946 2148 2947
rect 2230 2951 2236 2952
rect 2230 2947 2231 2951
rect 2235 2947 2236 2951
rect 2230 2946 2236 2947
rect 2318 2951 2324 2952
rect 2318 2947 2319 2951
rect 2323 2947 2324 2951
rect 2318 2946 2324 2947
rect 2406 2951 2412 2952
rect 2406 2947 2407 2951
rect 2411 2947 2412 2951
rect 2406 2946 2412 2947
rect 2494 2951 2500 2952
rect 2494 2947 2495 2951
rect 2499 2947 2500 2951
rect 2494 2946 2500 2947
rect 2582 2951 2588 2952
rect 2582 2947 2583 2951
rect 2587 2947 2588 2951
rect 2582 2946 2588 2947
rect 2670 2951 2676 2952
rect 2670 2947 2671 2951
rect 2675 2947 2676 2951
rect 2670 2946 2676 2947
rect 2758 2951 2764 2952
rect 2758 2947 2759 2951
rect 2763 2947 2764 2951
rect 2758 2946 2764 2947
rect 2846 2951 2852 2952
rect 2846 2947 2847 2951
rect 2851 2947 2852 2951
rect 3462 2948 3463 2952
rect 3467 2948 3468 2952
rect 3462 2947 3468 2948
rect 2846 2946 2852 2947
rect 1806 2935 1812 2936
rect 1806 2931 1807 2935
rect 1811 2931 1812 2935
rect 3462 2935 3468 2936
rect 111 2930 115 2931
rect 111 2925 115 2926
rect 135 2930 139 2931
rect 135 2925 139 2926
rect 263 2930 267 2931
rect 263 2925 267 2926
rect 327 2930 331 2931
rect 327 2925 331 2926
rect 431 2930 435 2931
rect 431 2925 435 2926
rect 535 2930 539 2931
rect 535 2925 539 2926
rect 607 2930 611 2931
rect 607 2925 611 2926
rect 735 2930 739 2931
rect 735 2925 739 2926
rect 783 2930 787 2931
rect 783 2925 787 2926
rect 927 2930 931 2931
rect 927 2925 931 2926
rect 951 2930 955 2931
rect 951 2925 955 2926
rect 1103 2930 1107 2931
rect 1103 2925 1107 2926
rect 1111 2930 1115 2931
rect 1111 2925 1115 2926
rect 1271 2930 1275 2931
rect 1271 2925 1275 2926
rect 1279 2930 1283 2931
rect 1279 2925 1283 2926
rect 1431 2930 1435 2931
rect 1431 2925 1435 2926
rect 1447 2930 1451 2931
rect 1447 2925 1451 2926
rect 1591 2930 1595 2931
rect 1591 2925 1595 2926
rect 1623 2930 1627 2931
rect 1623 2925 1627 2926
rect 1767 2930 1771 2931
rect 1806 2930 1812 2931
rect 2054 2932 2060 2933
rect 1767 2925 1771 2926
rect 112 2909 114 2925
rect 110 2908 116 2909
rect 136 2908 138 2925
rect 264 2908 266 2925
rect 432 2908 434 2925
rect 608 2908 610 2925
rect 784 2908 786 2925
rect 952 2908 954 2925
rect 1112 2908 1114 2925
rect 1272 2908 1274 2925
rect 1432 2908 1434 2925
rect 1592 2908 1594 2925
rect 1768 2909 1770 2925
rect 1766 2908 1772 2909
rect 110 2904 111 2908
rect 115 2904 116 2908
rect 110 2903 116 2904
rect 134 2907 140 2908
rect 134 2903 135 2907
rect 139 2903 140 2907
rect 134 2902 140 2903
rect 262 2907 268 2908
rect 262 2903 263 2907
rect 267 2903 268 2907
rect 262 2902 268 2903
rect 430 2907 436 2908
rect 430 2903 431 2907
rect 435 2903 436 2907
rect 430 2902 436 2903
rect 606 2907 612 2908
rect 606 2903 607 2907
rect 611 2903 612 2907
rect 606 2902 612 2903
rect 782 2907 788 2908
rect 782 2903 783 2907
rect 787 2903 788 2907
rect 782 2902 788 2903
rect 950 2907 956 2908
rect 950 2903 951 2907
rect 955 2903 956 2907
rect 950 2902 956 2903
rect 1110 2907 1116 2908
rect 1110 2903 1111 2907
rect 1115 2903 1116 2907
rect 1110 2902 1116 2903
rect 1270 2907 1276 2908
rect 1270 2903 1271 2907
rect 1275 2903 1276 2907
rect 1270 2902 1276 2903
rect 1430 2907 1436 2908
rect 1430 2903 1431 2907
rect 1435 2903 1436 2907
rect 1430 2902 1436 2903
rect 1590 2907 1596 2908
rect 1590 2903 1591 2907
rect 1595 2903 1596 2907
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1808 2903 1810 2930
rect 2054 2928 2055 2932
rect 2059 2928 2060 2932
rect 2054 2927 2060 2928
rect 2142 2932 2148 2933
rect 2142 2928 2143 2932
rect 2147 2928 2148 2932
rect 2142 2927 2148 2928
rect 2230 2932 2236 2933
rect 2230 2928 2231 2932
rect 2235 2928 2236 2932
rect 2230 2927 2236 2928
rect 2318 2932 2324 2933
rect 2318 2928 2319 2932
rect 2323 2928 2324 2932
rect 2318 2927 2324 2928
rect 2406 2932 2412 2933
rect 2406 2928 2407 2932
rect 2411 2928 2412 2932
rect 2406 2927 2412 2928
rect 2494 2932 2500 2933
rect 2494 2928 2495 2932
rect 2499 2928 2500 2932
rect 2494 2927 2500 2928
rect 2582 2932 2588 2933
rect 2582 2928 2583 2932
rect 2587 2928 2588 2932
rect 2582 2927 2588 2928
rect 2670 2932 2676 2933
rect 2670 2928 2671 2932
rect 2675 2928 2676 2932
rect 2670 2927 2676 2928
rect 2758 2932 2764 2933
rect 2758 2928 2759 2932
rect 2763 2928 2764 2932
rect 2758 2927 2764 2928
rect 2846 2932 2852 2933
rect 2846 2928 2847 2932
rect 2851 2928 2852 2932
rect 3462 2931 3463 2935
rect 3467 2931 3468 2935
rect 3462 2930 3468 2931
rect 2846 2927 2852 2928
rect 2056 2903 2058 2927
rect 2144 2903 2146 2927
rect 2232 2903 2234 2927
rect 2320 2903 2322 2927
rect 2408 2903 2410 2927
rect 2496 2903 2498 2927
rect 2584 2903 2586 2927
rect 2672 2903 2674 2927
rect 2760 2903 2762 2927
rect 2848 2903 2850 2927
rect 3464 2903 3466 2930
rect 1590 2902 1596 2903
rect 1807 2902 1811 2903
rect 1807 2897 1811 2898
rect 2055 2902 2059 2903
rect 2055 2897 2059 2898
rect 2071 2902 2075 2903
rect 2071 2897 2075 2898
rect 2143 2902 2147 2903
rect 2143 2897 2147 2898
rect 2175 2902 2179 2903
rect 2175 2897 2179 2898
rect 2231 2902 2235 2903
rect 2231 2897 2235 2898
rect 2271 2902 2275 2903
rect 2271 2897 2275 2898
rect 2319 2902 2323 2903
rect 2319 2897 2323 2898
rect 2367 2902 2371 2903
rect 2367 2897 2371 2898
rect 2407 2902 2411 2903
rect 2407 2897 2411 2898
rect 2471 2902 2475 2903
rect 2471 2897 2475 2898
rect 2495 2902 2499 2903
rect 2495 2897 2499 2898
rect 2575 2902 2579 2903
rect 2575 2897 2579 2898
rect 2583 2902 2587 2903
rect 2583 2897 2587 2898
rect 2671 2902 2675 2903
rect 2671 2897 2675 2898
rect 2679 2902 2683 2903
rect 2679 2897 2683 2898
rect 2759 2902 2763 2903
rect 2759 2897 2763 2898
rect 2783 2902 2787 2903
rect 2783 2897 2787 2898
rect 2847 2902 2851 2903
rect 2847 2897 2851 2898
rect 3463 2902 3467 2903
rect 3463 2897 3467 2898
rect 110 2891 116 2892
rect 110 2887 111 2891
rect 115 2887 116 2891
rect 1766 2891 1772 2892
rect 110 2886 116 2887
rect 134 2888 140 2889
rect 112 2863 114 2886
rect 134 2884 135 2888
rect 139 2884 140 2888
rect 134 2883 140 2884
rect 262 2888 268 2889
rect 262 2884 263 2888
rect 267 2884 268 2888
rect 262 2883 268 2884
rect 430 2888 436 2889
rect 430 2884 431 2888
rect 435 2884 436 2888
rect 430 2883 436 2884
rect 606 2888 612 2889
rect 606 2884 607 2888
rect 611 2884 612 2888
rect 606 2883 612 2884
rect 782 2888 788 2889
rect 782 2884 783 2888
rect 787 2884 788 2888
rect 782 2883 788 2884
rect 950 2888 956 2889
rect 950 2884 951 2888
rect 955 2884 956 2888
rect 950 2883 956 2884
rect 1110 2888 1116 2889
rect 1110 2884 1111 2888
rect 1115 2884 1116 2888
rect 1110 2883 1116 2884
rect 1270 2888 1276 2889
rect 1270 2884 1271 2888
rect 1275 2884 1276 2888
rect 1270 2883 1276 2884
rect 1430 2888 1436 2889
rect 1430 2884 1431 2888
rect 1435 2884 1436 2888
rect 1430 2883 1436 2884
rect 1590 2888 1596 2889
rect 1590 2884 1591 2888
rect 1595 2884 1596 2888
rect 1766 2887 1767 2891
rect 1771 2887 1772 2891
rect 1766 2886 1772 2887
rect 1590 2883 1596 2884
rect 136 2863 138 2883
rect 264 2863 266 2883
rect 432 2863 434 2883
rect 608 2863 610 2883
rect 784 2863 786 2883
rect 952 2863 954 2883
rect 1112 2863 1114 2883
rect 1272 2863 1274 2883
rect 1432 2863 1434 2883
rect 1592 2863 1594 2883
rect 1768 2863 1770 2886
rect 1808 2878 1810 2897
rect 2072 2881 2074 2897
rect 2176 2881 2178 2897
rect 2272 2881 2274 2897
rect 2368 2881 2370 2897
rect 2472 2881 2474 2897
rect 2576 2881 2578 2897
rect 2680 2881 2682 2897
rect 2784 2881 2786 2897
rect 2070 2880 2076 2881
rect 1806 2877 1812 2878
rect 1806 2873 1807 2877
rect 1811 2873 1812 2877
rect 2070 2876 2071 2880
rect 2075 2876 2076 2880
rect 2070 2875 2076 2876
rect 2174 2880 2180 2881
rect 2174 2876 2175 2880
rect 2179 2876 2180 2880
rect 2174 2875 2180 2876
rect 2270 2880 2276 2881
rect 2270 2876 2271 2880
rect 2275 2876 2276 2880
rect 2270 2875 2276 2876
rect 2366 2880 2372 2881
rect 2366 2876 2367 2880
rect 2371 2876 2372 2880
rect 2366 2875 2372 2876
rect 2470 2880 2476 2881
rect 2470 2876 2471 2880
rect 2475 2876 2476 2880
rect 2470 2875 2476 2876
rect 2574 2880 2580 2881
rect 2574 2876 2575 2880
rect 2579 2876 2580 2880
rect 2574 2875 2580 2876
rect 2678 2880 2684 2881
rect 2678 2876 2679 2880
rect 2683 2876 2684 2880
rect 2678 2875 2684 2876
rect 2782 2880 2788 2881
rect 2782 2876 2783 2880
rect 2787 2876 2788 2880
rect 3464 2878 3466 2897
rect 2782 2875 2788 2876
rect 3462 2877 3468 2878
rect 1806 2872 1812 2873
rect 3462 2873 3463 2877
rect 3467 2873 3468 2877
rect 3462 2872 3468 2873
rect 111 2862 115 2863
rect 111 2857 115 2858
rect 135 2862 139 2863
rect 135 2857 139 2858
rect 255 2862 259 2863
rect 255 2857 259 2858
rect 263 2862 267 2863
rect 263 2857 267 2858
rect 407 2862 411 2863
rect 407 2857 411 2858
rect 431 2862 435 2863
rect 431 2857 435 2858
rect 567 2862 571 2863
rect 567 2857 571 2858
rect 607 2862 611 2863
rect 607 2857 611 2858
rect 727 2862 731 2863
rect 727 2857 731 2858
rect 783 2862 787 2863
rect 783 2857 787 2858
rect 879 2862 883 2863
rect 879 2857 883 2858
rect 951 2862 955 2863
rect 951 2857 955 2858
rect 1023 2862 1027 2863
rect 1023 2857 1027 2858
rect 1111 2862 1115 2863
rect 1111 2857 1115 2858
rect 1167 2862 1171 2863
rect 1167 2857 1171 2858
rect 1271 2862 1275 2863
rect 1271 2857 1275 2858
rect 1311 2862 1315 2863
rect 1311 2857 1315 2858
rect 1431 2862 1435 2863
rect 1431 2857 1435 2858
rect 1463 2862 1467 2863
rect 1463 2857 1467 2858
rect 1591 2862 1595 2863
rect 1591 2857 1595 2858
rect 1767 2862 1771 2863
rect 2070 2861 2076 2862
rect 1767 2857 1771 2858
rect 1806 2860 1812 2861
rect 112 2838 114 2857
rect 136 2841 138 2857
rect 256 2841 258 2857
rect 408 2841 410 2857
rect 568 2841 570 2857
rect 728 2841 730 2857
rect 880 2841 882 2857
rect 1024 2841 1026 2857
rect 1168 2841 1170 2857
rect 1312 2841 1314 2857
rect 1464 2841 1466 2857
rect 134 2840 140 2841
rect 110 2837 116 2838
rect 110 2833 111 2837
rect 115 2833 116 2837
rect 134 2836 135 2840
rect 139 2836 140 2840
rect 134 2835 140 2836
rect 254 2840 260 2841
rect 254 2836 255 2840
rect 259 2836 260 2840
rect 254 2835 260 2836
rect 406 2840 412 2841
rect 406 2836 407 2840
rect 411 2836 412 2840
rect 406 2835 412 2836
rect 566 2840 572 2841
rect 566 2836 567 2840
rect 571 2836 572 2840
rect 566 2835 572 2836
rect 726 2840 732 2841
rect 726 2836 727 2840
rect 731 2836 732 2840
rect 726 2835 732 2836
rect 878 2840 884 2841
rect 878 2836 879 2840
rect 883 2836 884 2840
rect 878 2835 884 2836
rect 1022 2840 1028 2841
rect 1022 2836 1023 2840
rect 1027 2836 1028 2840
rect 1022 2835 1028 2836
rect 1166 2840 1172 2841
rect 1166 2836 1167 2840
rect 1171 2836 1172 2840
rect 1166 2835 1172 2836
rect 1310 2840 1316 2841
rect 1310 2836 1311 2840
rect 1315 2836 1316 2840
rect 1310 2835 1316 2836
rect 1462 2840 1468 2841
rect 1462 2836 1463 2840
rect 1467 2836 1468 2840
rect 1768 2838 1770 2857
rect 1806 2856 1807 2860
rect 1811 2856 1812 2860
rect 2070 2857 2071 2861
rect 2075 2857 2076 2861
rect 2070 2856 2076 2857
rect 2174 2861 2180 2862
rect 2174 2857 2175 2861
rect 2179 2857 2180 2861
rect 2174 2856 2180 2857
rect 2270 2861 2276 2862
rect 2270 2857 2271 2861
rect 2275 2857 2276 2861
rect 2270 2856 2276 2857
rect 2366 2861 2372 2862
rect 2366 2857 2367 2861
rect 2371 2857 2372 2861
rect 2366 2856 2372 2857
rect 2470 2861 2476 2862
rect 2470 2857 2471 2861
rect 2475 2857 2476 2861
rect 2470 2856 2476 2857
rect 2574 2861 2580 2862
rect 2574 2857 2575 2861
rect 2579 2857 2580 2861
rect 2574 2856 2580 2857
rect 2678 2861 2684 2862
rect 2678 2857 2679 2861
rect 2683 2857 2684 2861
rect 2678 2856 2684 2857
rect 2782 2861 2788 2862
rect 2782 2857 2783 2861
rect 2787 2857 2788 2861
rect 2782 2856 2788 2857
rect 3462 2860 3468 2861
rect 3462 2856 3463 2860
rect 3467 2856 3468 2860
rect 1806 2855 1812 2856
rect 1462 2835 1468 2836
rect 1766 2837 1772 2838
rect 110 2832 116 2833
rect 1766 2833 1767 2837
rect 1771 2833 1772 2837
rect 1808 2835 1810 2855
rect 2072 2835 2074 2856
rect 2176 2835 2178 2856
rect 2272 2835 2274 2856
rect 2368 2835 2370 2856
rect 2472 2835 2474 2856
rect 2576 2835 2578 2856
rect 2680 2835 2682 2856
rect 2784 2835 2786 2856
rect 3462 2855 3468 2856
rect 3464 2835 3466 2855
rect 1766 2832 1772 2833
rect 1807 2834 1811 2835
rect 1807 2829 1811 2830
rect 1983 2834 1987 2835
rect 1983 2829 1987 2830
rect 2071 2834 2075 2835
rect 2071 2829 2075 2830
rect 2111 2834 2115 2835
rect 2111 2829 2115 2830
rect 2175 2834 2179 2835
rect 2175 2829 2179 2830
rect 2239 2834 2243 2835
rect 2239 2829 2243 2830
rect 2271 2834 2275 2835
rect 2271 2829 2275 2830
rect 2367 2834 2371 2835
rect 2367 2829 2371 2830
rect 2471 2834 2475 2835
rect 2471 2829 2475 2830
rect 2487 2834 2491 2835
rect 2487 2829 2491 2830
rect 2575 2834 2579 2835
rect 2575 2829 2579 2830
rect 2607 2834 2611 2835
rect 2607 2829 2611 2830
rect 2679 2834 2683 2835
rect 2679 2829 2683 2830
rect 2719 2834 2723 2835
rect 2719 2829 2723 2830
rect 2783 2834 2787 2835
rect 2783 2829 2787 2830
rect 2839 2834 2843 2835
rect 2839 2829 2843 2830
rect 2959 2834 2963 2835
rect 2959 2829 2963 2830
rect 3463 2834 3467 2835
rect 3463 2829 3467 2830
rect 134 2821 140 2822
rect 110 2820 116 2821
rect 110 2816 111 2820
rect 115 2816 116 2820
rect 134 2817 135 2821
rect 139 2817 140 2821
rect 134 2816 140 2817
rect 254 2821 260 2822
rect 254 2817 255 2821
rect 259 2817 260 2821
rect 254 2816 260 2817
rect 406 2821 412 2822
rect 406 2817 407 2821
rect 411 2817 412 2821
rect 406 2816 412 2817
rect 566 2821 572 2822
rect 566 2817 567 2821
rect 571 2817 572 2821
rect 566 2816 572 2817
rect 726 2821 732 2822
rect 726 2817 727 2821
rect 731 2817 732 2821
rect 726 2816 732 2817
rect 878 2821 884 2822
rect 878 2817 879 2821
rect 883 2817 884 2821
rect 878 2816 884 2817
rect 1022 2821 1028 2822
rect 1022 2817 1023 2821
rect 1027 2817 1028 2821
rect 1022 2816 1028 2817
rect 1166 2821 1172 2822
rect 1166 2817 1167 2821
rect 1171 2817 1172 2821
rect 1166 2816 1172 2817
rect 1310 2821 1316 2822
rect 1310 2817 1311 2821
rect 1315 2817 1316 2821
rect 1310 2816 1316 2817
rect 1462 2821 1468 2822
rect 1462 2817 1463 2821
rect 1467 2817 1468 2821
rect 1462 2816 1468 2817
rect 1766 2820 1772 2821
rect 1766 2816 1767 2820
rect 1771 2816 1772 2820
rect 110 2815 116 2816
rect 112 2791 114 2815
rect 136 2791 138 2816
rect 256 2791 258 2816
rect 408 2791 410 2816
rect 568 2791 570 2816
rect 728 2791 730 2816
rect 880 2791 882 2816
rect 1024 2791 1026 2816
rect 1168 2791 1170 2816
rect 1312 2791 1314 2816
rect 1464 2791 1466 2816
rect 1766 2815 1772 2816
rect 1768 2791 1770 2815
rect 1808 2813 1810 2829
rect 1806 2812 1812 2813
rect 1984 2812 1986 2829
rect 2112 2812 2114 2829
rect 2240 2812 2242 2829
rect 2368 2812 2370 2829
rect 2488 2812 2490 2829
rect 2608 2812 2610 2829
rect 2720 2812 2722 2829
rect 2840 2812 2842 2829
rect 2960 2812 2962 2829
rect 3464 2813 3466 2829
rect 3462 2812 3468 2813
rect 1806 2808 1807 2812
rect 1811 2808 1812 2812
rect 1806 2807 1812 2808
rect 1982 2811 1988 2812
rect 1982 2807 1983 2811
rect 1987 2807 1988 2811
rect 1982 2806 1988 2807
rect 2110 2811 2116 2812
rect 2110 2807 2111 2811
rect 2115 2807 2116 2811
rect 2110 2806 2116 2807
rect 2238 2811 2244 2812
rect 2238 2807 2239 2811
rect 2243 2807 2244 2811
rect 2238 2806 2244 2807
rect 2366 2811 2372 2812
rect 2366 2807 2367 2811
rect 2371 2807 2372 2811
rect 2366 2806 2372 2807
rect 2486 2811 2492 2812
rect 2486 2807 2487 2811
rect 2491 2807 2492 2811
rect 2486 2806 2492 2807
rect 2606 2811 2612 2812
rect 2606 2807 2607 2811
rect 2611 2807 2612 2811
rect 2606 2806 2612 2807
rect 2718 2811 2724 2812
rect 2718 2807 2719 2811
rect 2723 2807 2724 2811
rect 2718 2806 2724 2807
rect 2838 2811 2844 2812
rect 2838 2807 2839 2811
rect 2843 2807 2844 2811
rect 2838 2806 2844 2807
rect 2958 2811 2964 2812
rect 2958 2807 2959 2811
rect 2963 2807 2964 2811
rect 3462 2808 3463 2812
rect 3467 2808 3468 2812
rect 3462 2807 3468 2808
rect 2958 2806 2964 2807
rect 1806 2795 1812 2796
rect 1806 2791 1807 2795
rect 1811 2791 1812 2795
rect 3462 2795 3468 2796
rect 111 2790 115 2791
rect 111 2785 115 2786
rect 135 2790 139 2791
rect 135 2785 139 2786
rect 255 2790 259 2791
rect 255 2785 259 2786
rect 287 2790 291 2791
rect 287 2785 291 2786
rect 391 2790 395 2791
rect 391 2785 395 2786
rect 407 2790 411 2791
rect 407 2785 411 2786
rect 503 2790 507 2791
rect 503 2785 507 2786
rect 567 2790 571 2791
rect 567 2785 571 2786
rect 623 2790 627 2791
rect 623 2785 627 2786
rect 727 2790 731 2791
rect 727 2785 731 2786
rect 743 2790 747 2791
rect 743 2785 747 2786
rect 855 2790 859 2791
rect 855 2785 859 2786
rect 879 2790 883 2791
rect 879 2785 883 2786
rect 967 2790 971 2791
rect 967 2785 971 2786
rect 1023 2790 1027 2791
rect 1023 2785 1027 2786
rect 1079 2790 1083 2791
rect 1079 2785 1083 2786
rect 1167 2790 1171 2791
rect 1167 2785 1171 2786
rect 1199 2790 1203 2791
rect 1199 2785 1203 2786
rect 1311 2790 1315 2791
rect 1311 2785 1315 2786
rect 1319 2790 1323 2791
rect 1319 2785 1323 2786
rect 1463 2790 1467 2791
rect 1463 2785 1467 2786
rect 1767 2790 1771 2791
rect 1806 2790 1812 2791
rect 1982 2792 1988 2793
rect 1767 2785 1771 2786
rect 112 2769 114 2785
rect 110 2768 116 2769
rect 288 2768 290 2785
rect 392 2768 394 2785
rect 504 2768 506 2785
rect 624 2768 626 2785
rect 744 2768 746 2785
rect 856 2768 858 2785
rect 968 2768 970 2785
rect 1080 2768 1082 2785
rect 1200 2768 1202 2785
rect 1320 2768 1322 2785
rect 1768 2769 1770 2785
rect 1766 2768 1772 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 286 2767 292 2768
rect 286 2763 287 2767
rect 291 2763 292 2767
rect 286 2762 292 2763
rect 390 2767 396 2768
rect 390 2763 391 2767
rect 395 2763 396 2767
rect 390 2762 396 2763
rect 502 2767 508 2768
rect 502 2763 503 2767
rect 507 2763 508 2767
rect 502 2762 508 2763
rect 622 2767 628 2768
rect 622 2763 623 2767
rect 627 2763 628 2767
rect 622 2762 628 2763
rect 742 2767 748 2768
rect 742 2763 743 2767
rect 747 2763 748 2767
rect 742 2762 748 2763
rect 854 2767 860 2768
rect 854 2763 855 2767
rect 859 2763 860 2767
rect 854 2762 860 2763
rect 966 2767 972 2768
rect 966 2763 967 2767
rect 971 2763 972 2767
rect 966 2762 972 2763
rect 1078 2767 1084 2768
rect 1078 2763 1079 2767
rect 1083 2763 1084 2767
rect 1078 2762 1084 2763
rect 1198 2767 1204 2768
rect 1198 2763 1199 2767
rect 1203 2763 1204 2767
rect 1198 2762 1204 2763
rect 1318 2767 1324 2768
rect 1318 2763 1319 2767
rect 1323 2763 1324 2767
rect 1766 2764 1767 2768
rect 1771 2764 1772 2768
rect 1808 2767 1810 2790
rect 1982 2788 1983 2792
rect 1987 2788 1988 2792
rect 1982 2787 1988 2788
rect 2110 2792 2116 2793
rect 2110 2788 2111 2792
rect 2115 2788 2116 2792
rect 2110 2787 2116 2788
rect 2238 2792 2244 2793
rect 2238 2788 2239 2792
rect 2243 2788 2244 2792
rect 2238 2787 2244 2788
rect 2366 2792 2372 2793
rect 2366 2788 2367 2792
rect 2371 2788 2372 2792
rect 2366 2787 2372 2788
rect 2486 2792 2492 2793
rect 2486 2788 2487 2792
rect 2491 2788 2492 2792
rect 2486 2787 2492 2788
rect 2606 2792 2612 2793
rect 2606 2788 2607 2792
rect 2611 2788 2612 2792
rect 2606 2787 2612 2788
rect 2718 2792 2724 2793
rect 2718 2788 2719 2792
rect 2723 2788 2724 2792
rect 2718 2787 2724 2788
rect 2838 2792 2844 2793
rect 2838 2788 2839 2792
rect 2843 2788 2844 2792
rect 2838 2787 2844 2788
rect 2958 2792 2964 2793
rect 2958 2788 2959 2792
rect 2963 2788 2964 2792
rect 3462 2791 3463 2795
rect 3467 2791 3468 2795
rect 3462 2790 3468 2791
rect 2958 2787 2964 2788
rect 1984 2767 1986 2787
rect 2112 2767 2114 2787
rect 2240 2767 2242 2787
rect 2368 2767 2370 2787
rect 2488 2767 2490 2787
rect 2608 2767 2610 2787
rect 2720 2767 2722 2787
rect 2840 2767 2842 2787
rect 2960 2767 2962 2787
rect 3464 2767 3466 2790
rect 1766 2763 1772 2764
rect 1807 2766 1811 2767
rect 1318 2762 1324 2763
rect 1807 2761 1811 2762
rect 1887 2766 1891 2767
rect 1887 2761 1891 2762
rect 1983 2766 1987 2767
rect 1983 2761 1987 2762
rect 2031 2766 2035 2767
rect 2031 2761 2035 2762
rect 2111 2766 2115 2767
rect 2111 2761 2115 2762
rect 2183 2766 2187 2767
rect 2183 2761 2187 2762
rect 2239 2766 2243 2767
rect 2239 2761 2243 2762
rect 2335 2766 2339 2767
rect 2335 2761 2339 2762
rect 2367 2766 2371 2767
rect 2367 2761 2371 2762
rect 2479 2766 2483 2767
rect 2479 2761 2483 2762
rect 2487 2766 2491 2767
rect 2487 2761 2491 2762
rect 2607 2766 2611 2767
rect 2607 2761 2611 2762
rect 2623 2766 2627 2767
rect 2623 2761 2627 2762
rect 2719 2766 2723 2767
rect 2719 2761 2723 2762
rect 2767 2766 2771 2767
rect 2767 2761 2771 2762
rect 2839 2766 2843 2767
rect 2839 2761 2843 2762
rect 2911 2766 2915 2767
rect 2911 2761 2915 2762
rect 2959 2766 2963 2767
rect 2959 2761 2963 2762
rect 3055 2766 3059 2767
rect 3055 2761 3059 2762
rect 3463 2766 3467 2767
rect 3463 2761 3467 2762
rect 110 2751 116 2752
rect 110 2747 111 2751
rect 115 2747 116 2751
rect 1766 2751 1772 2752
rect 110 2746 116 2747
rect 286 2748 292 2749
rect 112 2723 114 2746
rect 286 2744 287 2748
rect 291 2744 292 2748
rect 286 2743 292 2744
rect 390 2748 396 2749
rect 390 2744 391 2748
rect 395 2744 396 2748
rect 390 2743 396 2744
rect 502 2748 508 2749
rect 502 2744 503 2748
rect 507 2744 508 2748
rect 502 2743 508 2744
rect 622 2748 628 2749
rect 622 2744 623 2748
rect 627 2744 628 2748
rect 622 2743 628 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 854 2748 860 2749
rect 854 2744 855 2748
rect 859 2744 860 2748
rect 854 2743 860 2744
rect 966 2748 972 2749
rect 966 2744 967 2748
rect 971 2744 972 2748
rect 966 2743 972 2744
rect 1078 2748 1084 2749
rect 1078 2744 1079 2748
rect 1083 2744 1084 2748
rect 1078 2743 1084 2744
rect 1198 2748 1204 2749
rect 1198 2744 1199 2748
rect 1203 2744 1204 2748
rect 1198 2743 1204 2744
rect 1318 2748 1324 2749
rect 1318 2744 1319 2748
rect 1323 2744 1324 2748
rect 1766 2747 1767 2751
rect 1771 2747 1772 2751
rect 1766 2746 1772 2747
rect 1318 2743 1324 2744
rect 288 2723 290 2743
rect 392 2723 394 2743
rect 504 2723 506 2743
rect 624 2723 626 2743
rect 744 2723 746 2743
rect 856 2723 858 2743
rect 968 2723 970 2743
rect 1080 2723 1082 2743
rect 1200 2723 1202 2743
rect 1320 2723 1322 2743
rect 1768 2723 1770 2746
rect 1808 2742 1810 2761
rect 1888 2745 1890 2761
rect 2032 2745 2034 2761
rect 2184 2745 2186 2761
rect 2336 2745 2338 2761
rect 2480 2745 2482 2761
rect 2624 2745 2626 2761
rect 2768 2745 2770 2761
rect 2912 2745 2914 2761
rect 3056 2745 3058 2761
rect 1886 2744 1892 2745
rect 1806 2741 1812 2742
rect 1806 2737 1807 2741
rect 1811 2737 1812 2741
rect 1886 2740 1887 2744
rect 1891 2740 1892 2744
rect 1886 2739 1892 2740
rect 2030 2744 2036 2745
rect 2030 2740 2031 2744
rect 2035 2740 2036 2744
rect 2030 2739 2036 2740
rect 2182 2744 2188 2745
rect 2182 2740 2183 2744
rect 2187 2740 2188 2744
rect 2182 2739 2188 2740
rect 2334 2744 2340 2745
rect 2334 2740 2335 2744
rect 2339 2740 2340 2744
rect 2334 2739 2340 2740
rect 2478 2744 2484 2745
rect 2478 2740 2479 2744
rect 2483 2740 2484 2744
rect 2478 2739 2484 2740
rect 2622 2744 2628 2745
rect 2622 2740 2623 2744
rect 2627 2740 2628 2744
rect 2622 2739 2628 2740
rect 2766 2744 2772 2745
rect 2766 2740 2767 2744
rect 2771 2740 2772 2744
rect 2766 2739 2772 2740
rect 2910 2744 2916 2745
rect 2910 2740 2911 2744
rect 2915 2740 2916 2744
rect 2910 2739 2916 2740
rect 3054 2744 3060 2745
rect 3054 2740 3055 2744
rect 3059 2740 3060 2744
rect 3464 2742 3466 2761
rect 3054 2739 3060 2740
rect 3462 2741 3468 2742
rect 1806 2736 1812 2737
rect 3462 2737 3463 2741
rect 3467 2737 3468 2741
rect 3462 2736 3468 2737
rect 1886 2725 1892 2726
rect 1806 2724 1812 2725
rect 111 2722 115 2723
rect 111 2717 115 2718
rect 287 2722 291 2723
rect 287 2717 291 2718
rect 391 2722 395 2723
rect 391 2717 395 2718
rect 479 2722 483 2723
rect 479 2717 483 2718
rect 503 2722 507 2723
rect 503 2717 507 2718
rect 567 2722 571 2723
rect 567 2717 571 2718
rect 623 2722 627 2723
rect 623 2717 627 2718
rect 655 2722 659 2723
rect 655 2717 659 2718
rect 743 2722 747 2723
rect 743 2717 747 2718
rect 831 2722 835 2723
rect 831 2717 835 2718
rect 855 2722 859 2723
rect 855 2717 859 2718
rect 919 2722 923 2723
rect 919 2717 923 2718
rect 967 2722 971 2723
rect 967 2717 971 2718
rect 1007 2722 1011 2723
rect 1007 2717 1011 2718
rect 1079 2722 1083 2723
rect 1079 2717 1083 2718
rect 1095 2722 1099 2723
rect 1095 2717 1099 2718
rect 1183 2722 1187 2723
rect 1183 2717 1187 2718
rect 1199 2722 1203 2723
rect 1199 2717 1203 2718
rect 1319 2722 1323 2723
rect 1319 2717 1323 2718
rect 1767 2722 1771 2723
rect 1806 2720 1807 2724
rect 1811 2720 1812 2724
rect 1886 2721 1887 2725
rect 1891 2721 1892 2725
rect 1886 2720 1892 2721
rect 2030 2725 2036 2726
rect 2030 2721 2031 2725
rect 2035 2721 2036 2725
rect 2030 2720 2036 2721
rect 2182 2725 2188 2726
rect 2182 2721 2183 2725
rect 2187 2721 2188 2725
rect 2182 2720 2188 2721
rect 2334 2725 2340 2726
rect 2334 2721 2335 2725
rect 2339 2721 2340 2725
rect 2334 2720 2340 2721
rect 2478 2725 2484 2726
rect 2478 2721 2479 2725
rect 2483 2721 2484 2725
rect 2478 2720 2484 2721
rect 2622 2725 2628 2726
rect 2622 2721 2623 2725
rect 2627 2721 2628 2725
rect 2622 2720 2628 2721
rect 2766 2725 2772 2726
rect 2766 2721 2767 2725
rect 2771 2721 2772 2725
rect 2766 2720 2772 2721
rect 2910 2725 2916 2726
rect 2910 2721 2911 2725
rect 2915 2721 2916 2725
rect 2910 2720 2916 2721
rect 3054 2725 3060 2726
rect 3054 2721 3055 2725
rect 3059 2721 3060 2725
rect 3054 2720 3060 2721
rect 3462 2724 3468 2725
rect 3462 2720 3463 2724
rect 3467 2720 3468 2724
rect 1806 2719 1812 2720
rect 1767 2717 1771 2718
rect 112 2698 114 2717
rect 480 2701 482 2717
rect 568 2701 570 2717
rect 656 2701 658 2717
rect 744 2701 746 2717
rect 832 2701 834 2717
rect 920 2701 922 2717
rect 1008 2701 1010 2717
rect 1096 2701 1098 2717
rect 1184 2701 1186 2717
rect 478 2700 484 2701
rect 110 2697 116 2698
rect 110 2693 111 2697
rect 115 2693 116 2697
rect 478 2696 479 2700
rect 483 2696 484 2700
rect 478 2695 484 2696
rect 566 2700 572 2701
rect 566 2696 567 2700
rect 571 2696 572 2700
rect 566 2695 572 2696
rect 654 2700 660 2701
rect 654 2696 655 2700
rect 659 2696 660 2700
rect 654 2695 660 2696
rect 742 2700 748 2701
rect 742 2696 743 2700
rect 747 2696 748 2700
rect 742 2695 748 2696
rect 830 2700 836 2701
rect 830 2696 831 2700
rect 835 2696 836 2700
rect 830 2695 836 2696
rect 918 2700 924 2701
rect 918 2696 919 2700
rect 923 2696 924 2700
rect 918 2695 924 2696
rect 1006 2700 1012 2701
rect 1006 2696 1007 2700
rect 1011 2696 1012 2700
rect 1006 2695 1012 2696
rect 1094 2700 1100 2701
rect 1094 2696 1095 2700
rect 1099 2696 1100 2700
rect 1094 2695 1100 2696
rect 1182 2700 1188 2701
rect 1182 2696 1183 2700
rect 1187 2696 1188 2700
rect 1768 2698 1770 2717
rect 1808 2703 1810 2719
rect 1888 2703 1890 2720
rect 2032 2703 2034 2720
rect 2184 2703 2186 2720
rect 2336 2703 2338 2720
rect 2480 2703 2482 2720
rect 2624 2703 2626 2720
rect 2768 2703 2770 2720
rect 2912 2703 2914 2720
rect 3056 2703 3058 2720
rect 3462 2719 3468 2720
rect 3464 2703 3466 2719
rect 1807 2702 1811 2703
rect 1182 2695 1188 2696
rect 1766 2697 1772 2698
rect 1807 2697 1811 2698
rect 1831 2702 1835 2703
rect 1831 2697 1835 2698
rect 1887 2702 1891 2703
rect 1887 2697 1891 2698
rect 2023 2702 2027 2703
rect 2023 2697 2027 2698
rect 2031 2702 2035 2703
rect 2031 2697 2035 2698
rect 2183 2702 2187 2703
rect 2183 2697 2187 2698
rect 2231 2702 2235 2703
rect 2231 2697 2235 2698
rect 2335 2702 2339 2703
rect 2335 2697 2339 2698
rect 2431 2702 2435 2703
rect 2431 2697 2435 2698
rect 2479 2702 2483 2703
rect 2479 2697 2483 2698
rect 2615 2702 2619 2703
rect 2615 2697 2619 2698
rect 2623 2702 2627 2703
rect 2623 2697 2627 2698
rect 2767 2702 2771 2703
rect 2767 2697 2771 2698
rect 2783 2702 2787 2703
rect 2783 2697 2787 2698
rect 2911 2702 2915 2703
rect 2911 2697 2915 2698
rect 2943 2702 2947 2703
rect 2943 2697 2947 2698
rect 3055 2702 3059 2703
rect 3055 2697 3059 2698
rect 3095 2702 3099 2703
rect 3095 2697 3099 2698
rect 3239 2702 3243 2703
rect 3239 2697 3243 2698
rect 3367 2702 3371 2703
rect 3367 2697 3371 2698
rect 3463 2702 3467 2703
rect 3463 2697 3467 2698
rect 110 2692 116 2693
rect 1766 2693 1767 2697
rect 1771 2693 1772 2697
rect 1766 2692 1772 2693
rect 478 2681 484 2682
rect 110 2680 116 2681
rect 110 2676 111 2680
rect 115 2676 116 2680
rect 478 2677 479 2681
rect 483 2677 484 2681
rect 478 2676 484 2677
rect 566 2681 572 2682
rect 566 2677 567 2681
rect 571 2677 572 2681
rect 566 2676 572 2677
rect 654 2681 660 2682
rect 654 2677 655 2681
rect 659 2677 660 2681
rect 654 2676 660 2677
rect 742 2681 748 2682
rect 742 2677 743 2681
rect 747 2677 748 2681
rect 742 2676 748 2677
rect 830 2681 836 2682
rect 830 2677 831 2681
rect 835 2677 836 2681
rect 830 2676 836 2677
rect 918 2681 924 2682
rect 918 2677 919 2681
rect 923 2677 924 2681
rect 918 2676 924 2677
rect 1006 2681 1012 2682
rect 1006 2677 1007 2681
rect 1011 2677 1012 2681
rect 1006 2676 1012 2677
rect 1094 2681 1100 2682
rect 1094 2677 1095 2681
rect 1099 2677 1100 2681
rect 1094 2676 1100 2677
rect 1182 2681 1188 2682
rect 1808 2681 1810 2697
rect 1182 2677 1183 2681
rect 1187 2677 1188 2681
rect 1182 2676 1188 2677
rect 1766 2680 1772 2681
rect 1766 2676 1767 2680
rect 1771 2676 1772 2680
rect 110 2675 116 2676
rect 112 2651 114 2675
rect 480 2651 482 2676
rect 568 2651 570 2676
rect 656 2651 658 2676
rect 744 2651 746 2676
rect 832 2651 834 2676
rect 920 2651 922 2676
rect 1008 2651 1010 2676
rect 1096 2651 1098 2676
rect 1184 2651 1186 2676
rect 1766 2675 1772 2676
rect 1806 2680 1812 2681
rect 1832 2680 1834 2697
rect 2024 2680 2026 2697
rect 2232 2680 2234 2697
rect 2432 2680 2434 2697
rect 2616 2680 2618 2697
rect 2784 2680 2786 2697
rect 2944 2680 2946 2697
rect 3096 2680 3098 2697
rect 3240 2680 3242 2697
rect 3368 2680 3370 2697
rect 3464 2681 3466 2697
rect 3462 2680 3468 2681
rect 1806 2676 1807 2680
rect 1811 2676 1812 2680
rect 1806 2675 1812 2676
rect 1830 2679 1836 2680
rect 1830 2675 1831 2679
rect 1835 2675 1836 2679
rect 1768 2651 1770 2675
rect 1830 2674 1836 2675
rect 2022 2679 2028 2680
rect 2022 2675 2023 2679
rect 2027 2675 2028 2679
rect 2022 2674 2028 2675
rect 2230 2679 2236 2680
rect 2230 2675 2231 2679
rect 2235 2675 2236 2679
rect 2230 2674 2236 2675
rect 2430 2679 2436 2680
rect 2430 2675 2431 2679
rect 2435 2675 2436 2679
rect 2430 2674 2436 2675
rect 2614 2679 2620 2680
rect 2614 2675 2615 2679
rect 2619 2675 2620 2679
rect 2614 2674 2620 2675
rect 2782 2679 2788 2680
rect 2782 2675 2783 2679
rect 2787 2675 2788 2679
rect 2782 2674 2788 2675
rect 2942 2679 2948 2680
rect 2942 2675 2943 2679
rect 2947 2675 2948 2679
rect 2942 2674 2948 2675
rect 3094 2679 3100 2680
rect 3094 2675 3095 2679
rect 3099 2675 3100 2679
rect 3094 2674 3100 2675
rect 3238 2679 3244 2680
rect 3238 2675 3239 2679
rect 3243 2675 3244 2679
rect 3238 2674 3244 2675
rect 3366 2679 3372 2680
rect 3366 2675 3367 2679
rect 3371 2675 3372 2679
rect 3462 2676 3463 2680
rect 3467 2676 3468 2680
rect 3462 2675 3468 2676
rect 3366 2674 3372 2675
rect 1806 2663 1812 2664
rect 1806 2659 1807 2663
rect 1811 2659 1812 2663
rect 3462 2663 3468 2664
rect 1806 2658 1812 2659
rect 1830 2660 1836 2661
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 471 2650 475 2651
rect 471 2645 475 2646
rect 479 2650 483 2651
rect 479 2645 483 2646
rect 559 2650 563 2651
rect 559 2645 563 2646
rect 567 2650 571 2651
rect 567 2645 571 2646
rect 647 2650 651 2651
rect 647 2645 651 2646
rect 655 2650 659 2651
rect 655 2645 659 2646
rect 735 2650 739 2651
rect 735 2645 739 2646
rect 743 2650 747 2651
rect 743 2645 747 2646
rect 823 2650 827 2651
rect 823 2645 827 2646
rect 831 2650 835 2651
rect 831 2645 835 2646
rect 911 2650 915 2651
rect 911 2645 915 2646
rect 919 2650 923 2651
rect 919 2645 923 2646
rect 999 2650 1003 2651
rect 999 2645 1003 2646
rect 1007 2650 1011 2651
rect 1007 2645 1011 2646
rect 1087 2650 1091 2651
rect 1087 2645 1091 2646
rect 1095 2650 1099 2651
rect 1095 2645 1099 2646
rect 1183 2650 1187 2651
rect 1183 2645 1187 2646
rect 1767 2650 1771 2651
rect 1767 2645 1771 2646
rect 112 2629 114 2645
rect 110 2628 116 2629
rect 472 2628 474 2645
rect 560 2628 562 2645
rect 648 2628 650 2645
rect 736 2628 738 2645
rect 824 2628 826 2645
rect 912 2628 914 2645
rect 1000 2628 1002 2645
rect 1088 2628 1090 2645
rect 1768 2629 1770 2645
rect 1808 2635 1810 2658
rect 1830 2656 1831 2660
rect 1835 2656 1836 2660
rect 1830 2655 1836 2656
rect 2022 2660 2028 2661
rect 2022 2656 2023 2660
rect 2027 2656 2028 2660
rect 2022 2655 2028 2656
rect 2230 2660 2236 2661
rect 2230 2656 2231 2660
rect 2235 2656 2236 2660
rect 2230 2655 2236 2656
rect 2430 2660 2436 2661
rect 2430 2656 2431 2660
rect 2435 2656 2436 2660
rect 2430 2655 2436 2656
rect 2614 2660 2620 2661
rect 2614 2656 2615 2660
rect 2619 2656 2620 2660
rect 2614 2655 2620 2656
rect 2782 2660 2788 2661
rect 2782 2656 2783 2660
rect 2787 2656 2788 2660
rect 2782 2655 2788 2656
rect 2942 2660 2948 2661
rect 2942 2656 2943 2660
rect 2947 2656 2948 2660
rect 2942 2655 2948 2656
rect 3094 2660 3100 2661
rect 3094 2656 3095 2660
rect 3099 2656 3100 2660
rect 3094 2655 3100 2656
rect 3238 2660 3244 2661
rect 3238 2656 3239 2660
rect 3243 2656 3244 2660
rect 3238 2655 3244 2656
rect 3366 2660 3372 2661
rect 3366 2656 3367 2660
rect 3371 2656 3372 2660
rect 3462 2659 3463 2663
rect 3467 2659 3468 2663
rect 3462 2658 3468 2659
rect 3366 2655 3372 2656
rect 1832 2635 1834 2655
rect 2024 2635 2026 2655
rect 2232 2635 2234 2655
rect 2432 2635 2434 2655
rect 2616 2635 2618 2655
rect 2784 2635 2786 2655
rect 2944 2635 2946 2655
rect 3096 2635 3098 2655
rect 3240 2635 3242 2655
rect 3368 2635 3370 2655
rect 3464 2635 3466 2658
rect 1807 2634 1811 2635
rect 1807 2629 1811 2630
rect 1831 2634 1835 2635
rect 1831 2629 1835 2630
rect 1999 2634 2003 2635
rect 1999 2629 2003 2630
rect 2023 2634 2027 2635
rect 2023 2629 2027 2630
rect 2183 2634 2187 2635
rect 2183 2629 2187 2630
rect 2231 2634 2235 2635
rect 2231 2629 2235 2630
rect 2359 2634 2363 2635
rect 2359 2629 2363 2630
rect 2431 2634 2435 2635
rect 2431 2629 2435 2630
rect 2519 2634 2523 2635
rect 2519 2629 2523 2630
rect 2615 2634 2619 2635
rect 2615 2629 2619 2630
rect 2671 2634 2675 2635
rect 2671 2629 2675 2630
rect 2783 2634 2787 2635
rect 2783 2629 2787 2630
rect 2807 2634 2811 2635
rect 2807 2629 2811 2630
rect 2927 2634 2931 2635
rect 2927 2629 2931 2630
rect 2943 2634 2947 2635
rect 2943 2629 2947 2630
rect 3047 2634 3051 2635
rect 3047 2629 3051 2630
rect 3095 2634 3099 2635
rect 3095 2629 3099 2630
rect 3159 2634 3163 2635
rect 3159 2629 3163 2630
rect 3239 2634 3243 2635
rect 3239 2629 3243 2630
rect 3271 2634 3275 2635
rect 3271 2629 3275 2630
rect 3367 2634 3371 2635
rect 3367 2629 3371 2630
rect 3463 2634 3467 2635
rect 3463 2629 3467 2630
rect 1766 2628 1772 2629
rect 110 2624 111 2628
rect 115 2624 116 2628
rect 110 2623 116 2624
rect 470 2627 476 2628
rect 470 2623 471 2627
rect 475 2623 476 2627
rect 470 2622 476 2623
rect 558 2627 564 2628
rect 558 2623 559 2627
rect 563 2623 564 2627
rect 558 2622 564 2623
rect 646 2627 652 2628
rect 646 2623 647 2627
rect 651 2623 652 2627
rect 646 2622 652 2623
rect 734 2627 740 2628
rect 734 2623 735 2627
rect 739 2623 740 2627
rect 734 2622 740 2623
rect 822 2627 828 2628
rect 822 2623 823 2627
rect 827 2623 828 2627
rect 822 2622 828 2623
rect 910 2627 916 2628
rect 910 2623 911 2627
rect 915 2623 916 2627
rect 910 2622 916 2623
rect 998 2627 1004 2628
rect 998 2623 999 2627
rect 1003 2623 1004 2627
rect 998 2622 1004 2623
rect 1086 2627 1092 2628
rect 1086 2623 1087 2627
rect 1091 2623 1092 2627
rect 1766 2624 1767 2628
rect 1771 2624 1772 2628
rect 1766 2623 1772 2624
rect 1086 2622 1092 2623
rect 110 2611 116 2612
rect 110 2607 111 2611
rect 115 2607 116 2611
rect 1766 2611 1772 2612
rect 110 2606 116 2607
rect 470 2608 476 2609
rect 112 2575 114 2606
rect 470 2604 471 2608
rect 475 2604 476 2608
rect 470 2603 476 2604
rect 558 2608 564 2609
rect 558 2604 559 2608
rect 563 2604 564 2608
rect 558 2603 564 2604
rect 646 2608 652 2609
rect 646 2604 647 2608
rect 651 2604 652 2608
rect 646 2603 652 2604
rect 734 2608 740 2609
rect 734 2604 735 2608
rect 739 2604 740 2608
rect 734 2603 740 2604
rect 822 2608 828 2609
rect 822 2604 823 2608
rect 827 2604 828 2608
rect 822 2603 828 2604
rect 910 2608 916 2609
rect 910 2604 911 2608
rect 915 2604 916 2608
rect 910 2603 916 2604
rect 998 2608 1004 2609
rect 998 2604 999 2608
rect 1003 2604 1004 2608
rect 998 2603 1004 2604
rect 1086 2608 1092 2609
rect 1086 2604 1087 2608
rect 1091 2604 1092 2608
rect 1766 2607 1767 2611
rect 1771 2607 1772 2611
rect 1808 2610 1810 2629
rect 1832 2613 1834 2629
rect 2000 2613 2002 2629
rect 2184 2613 2186 2629
rect 2360 2613 2362 2629
rect 2520 2613 2522 2629
rect 2672 2613 2674 2629
rect 2808 2613 2810 2629
rect 2928 2613 2930 2629
rect 3048 2613 3050 2629
rect 3160 2613 3162 2629
rect 3272 2613 3274 2629
rect 3368 2613 3370 2629
rect 1830 2612 1836 2613
rect 1766 2606 1772 2607
rect 1806 2609 1812 2610
rect 1086 2603 1092 2604
rect 472 2575 474 2603
rect 560 2575 562 2603
rect 648 2575 650 2603
rect 736 2575 738 2603
rect 824 2575 826 2603
rect 912 2575 914 2603
rect 1000 2575 1002 2603
rect 1088 2575 1090 2603
rect 1768 2575 1770 2606
rect 1806 2605 1807 2609
rect 1811 2605 1812 2609
rect 1830 2608 1831 2612
rect 1835 2608 1836 2612
rect 1830 2607 1836 2608
rect 1998 2612 2004 2613
rect 1998 2608 1999 2612
rect 2003 2608 2004 2612
rect 1998 2607 2004 2608
rect 2182 2612 2188 2613
rect 2182 2608 2183 2612
rect 2187 2608 2188 2612
rect 2182 2607 2188 2608
rect 2358 2612 2364 2613
rect 2358 2608 2359 2612
rect 2363 2608 2364 2612
rect 2358 2607 2364 2608
rect 2518 2612 2524 2613
rect 2518 2608 2519 2612
rect 2523 2608 2524 2612
rect 2518 2607 2524 2608
rect 2670 2612 2676 2613
rect 2670 2608 2671 2612
rect 2675 2608 2676 2612
rect 2670 2607 2676 2608
rect 2806 2612 2812 2613
rect 2806 2608 2807 2612
rect 2811 2608 2812 2612
rect 2806 2607 2812 2608
rect 2926 2612 2932 2613
rect 2926 2608 2927 2612
rect 2931 2608 2932 2612
rect 2926 2607 2932 2608
rect 3046 2612 3052 2613
rect 3046 2608 3047 2612
rect 3051 2608 3052 2612
rect 3046 2607 3052 2608
rect 3158 2612 3164 2613
rect 3158 2608 3159 2612
rect 3163 2608 3164 2612
rect 3158 2607 3164 2608
rect 3270 2612 3276 2613
rect 3270 2608 3271 2612
rect 3275 2608 3276 2612
rect 3270 2607 3276 2608
rect 3366 2612 3372 2613
rect 3366 2608 3367 2612
rect 3371 2608 3372 2612
rect 3464 2610 3466 2629
rect 3366 2607 3372 2608
rect 3462 2609 3468 2610
rect 1806 2604 1812 2605
rect 3462 2605 3463 2609
rect 3467 2605 3468 2609
rect 3462 2604 3468 2605
rect 1830 2593 1836 2594
rect 1806 2592 1812 2593
rect 1806 2588 1807 2592
rect 1811 2588 1812 2592
rect 1830 2589 1831 2593
rect 1835 2589 1836 2593
rect 1830 2588 1836 2589
rect 1998 2593 2004 2594
rect 1998 2589 1999 2593
rect 2003 2589 2004 2593
rect 1998 2588 2004 2589
rect 2182 2593 2188 2594
rect 2182 2589 2183 2593
rect 2187 2589 2188 2593
rect 2182 2588 2188 2589
rect 2358 2593 2364 2594
rect 2358 2589 2359 2593
rect 2363 2589 2364 2593
rect 2358 2588 2364 2589
rect 2518 2593 2524 2594
rect 2518 2589 2519 2593
rect 2523 2589 2524 2593
rect 2518 2588 2524 2589
rect 2670 2593 2676 2594
rect 2670 2589 2671 2593
rect 2675 2589 2676 2593
rect 2670 2588 2676 2589
rect 2806 2593 2812 2594
rect 2806 2589 2807 2593
rect 2811 2589 2812 2593
rect 2806 2588 2812 2589
rect 2926 2593 2932 2594
rect 2926 2589 2927 2593
rect 2931 2589 2932 2593
rect 2926 2588 2932 2589
rect 3046 2593 3052 2594
rect 3046 2589 3047 2593
rect 3051 2589 3052 2593
rect 3046 2588 3052 2589
rect 3158 2593 3164 2594
rect 3158 2589 3159 2593
rect 3163 2589 3164 2593
rect 3158 2588 3164 2589
rect 3270 2593 3276 2594
rect 3270 2589 3271 2593
rect 3275 2589 3276 2593
rect 3270 2588 3276 2589
rect 3366 2593 3372 2594
rect 3366 2589 3367 2593
rect 3371 2589 3372 2593
rect 3366 2588 3372 2589
rect 3462 2592 3468 2593
rect 3462 2588 3463 2592
rect 3467 2588 3468 2592
rect 1806 2587 1812 2588
rect 111 2574 115 2575
rect 111 2569 115 2570
rect 223 2574 227 2575
rect 223 2569 227 2570
rect 311 2574 315 2575
rect 311 2569 315 2570
rect 407 2574 411 2575
rect 407 2569 411 2570
rect 471 2574 475 2575
rect 471 2569 475 2570
rect 503 2574 507 2575
rect 503 2569 507 2570
rect 559 2574 563 2575
rect 559 2569 563 2570
rect 591 2574 595 2575
rect 591 2569 595 2570
rect 647 2574 651 2575
rect 647 2569 651 2570
rect 679 2574 683 2575
rect 679 2569 683 2570
rect 735 2574 739 2575
rect 735 2569 739 2570
rect 767 2574 771 2575
rect 767 2569 771 2570
rect 823 2574 827 2575
rect 823 2569 827 2570
rect 855 2574 859 2575
rect 855 2569 859 2570
rect 911 2574 915 2575
rect 911 2569 915 2570
rect 943 2574 947 2575
rect 943 2569 947 2570
rect 999 2574 1003 2575
rect 999 2569 1003 2570
rect 1031 2574 1035 2575
rect 1031 2569 1035 2570
rect 1087 2574 1091 2575
rect 1087 2569 1091 2570
rect 1119 2574 1123 2575
rect 1119 2569 1123 2570
rect 1215 2574 1219 2575
rect 1215 2569 1219 2570
rect 1311 2574 1315 2575
rect 1311 2569 1315 2570
rect 1407 2574 1411 2575
rect 1407 2569 1411 2570
rect 1495 2574 1499 2575
rect 1495 2569 1499 2570
rect 1583 2574 1587 2575
rect 1583 2569 1587 2570
rect 1671 2574 1675 2575
rect 1671 2569 1675 2570
rect 1767 2574 1771 2575
rect 1767 2569 1771 2570
rect 112 2550 114 2569
rect 224 2553 226 2569
rect 312 2553 314 2569
rect 408 2553 410 2569
rect 504 2553 506 2569
rect 592 2553 594 2569
rect 680 2553 682 2569
rect 768 2553 770 2569
rect 856 2553 858 2569
rect 944 2553 946 2569
rect 1032 2553 1034 2569
rect 1120 2553 1122 2569
rect 1216 2553 1218 2569
rect 1312 2553 1314 2569
rect 1408 2553 1410 2569
rect 1496 2553 1498 2569
rect 1584 2553 1586 2569
rect 1672 2553 1674 2569
rect 222 2552 228 2553
rect 110 2549 116 2550
rect 110 2545 111 2549
rect 115 2545 116 2549
rect 222 2548 223 2552
rect 227 2548 228 2552
rect 222 2547 228 2548
rect 310 2552 316 2553
rect 310 2548 311 2552
rect 315 2548 316 2552
rect 310 2547 316 2548
rect 406 2552 412 2553
rect 406 2548 407 2552
rect 411 2548 412 2552
rect 406 2547 412 2548
rect 502 2552 508 2553
rect 502 2548 503 2552
rect 507 2548 508 2552
rect 502 2547 508 2548
rect 590 2552 596 2553
rect 590 2548 591 2552
rect 595 2548 596 2552
rect 590 2547 596 2548
rect 678 2552 684 2553
rect 678 2548 679 2552
rect 683 2548 684 2552
rect 678 2547 684 2548
rect 766 2552 772 2553
rect 766 2548 767 2552
rect 771 2548 772 2552
rect 766 2547 772 2548
rect 854 2552 860 2553
rect 854 2548 855 2552
rect 859 2548 860 2552
rect 854 2547 860 2548
rect 942 2552 948 2553
rect 942 2548 943 2552
rect 947 2548 948 2552
rect 942 2547 948 2548
rect 1030 2552 1036 2553
rect 1030 2548 1031 2552
rect 1035 2548 1036 2552
rect 1030 2547 1036 2548
rect 1118 2552 1124 2553
rect 1118 2548 1119 2552
rect 1123 2548 1124 2552
rect 1118 2547 1124 2548
rect 1214 2552 1220 2553
rect 1214 2548 1215 2552
rect 1219 2548 1220 2552
rect 1214 2547 1220 2548
rect 1310 2552 1316 2553
rect 1310 2548 1311 2552
rect 1315 2548 1316 2552
rect 1310 2547 1316 2548
rect 1406 2552 1412 2553
rect 1406 2548 1407 2552
rect 1411 2548 1412 2552
rect 1406 2547 1412 2548
rect 1494 2552 1500 2553
rect 1494 2548 1495 2552
rect 1499 2548 1500 2552
rect 1494 2547 1500 2548
rect 1582 2552 1588 2553
rect 1582 2548 1583 2552
rect 1587 2548 1588 2552
rect 1582 2547 1588 2548
rect 1670 2552 1676 2553
rect 1670 2548 1671 2552
rect 1675 2548 1676 2552
rect 1768 2550 1770 2569
rect 1808 2563 1810 2587
rect 1832 2563 1834 2588
rect 2000 2563 2002 2588
rect 2184 2563 2186 2588
rect 2360 2563 2362 2588
rect 2520 2563 2522 2588
rect 2672 2563 2674 2588
rect 2808 2563 2810 2588
rect 2928 2563 2930 2588
rect 3048 2563 3050 2588
rect 3160 2563 3162 2588
rect 3272 2563 3274 2588
rect 3368 2563 3370 2588
rect 3462 2587 3468 2588
rect 3464 2563 3466 2587
rect 1807 2562 1811 2563
rect 1807 2557 1811 2558
rect 1831 2562 1835 2563
rect 1831 2557 1835 2558
rect 1999 2562 2003 2563
rect 1999 2557 2003 2558
rect 2183 2562 2187 2563
rect 2183 2557 2187 2558
rect 2207 2562 2211 2563
rect 2207 2557 2211 2558
rect 2359 2562 2363 2563
rect 2359 2557 2363 2558
rect 2519 2562 2523 2563
rect 2519 2557 2523 2558
rect 2671 2562 2675 2563
rect 2671 2557 2675 2558
rect 2799 2562 2803 2563
rect 2799 2557 2803 2558
rect 2807 2562 2811 2563
rect 2807 2557 2811 2558
rect 2927 2562 2931 2563
rect 2927 2557 2931 2558
rect 3047 2562 3051 2563
rect 3047 2557 3051 2558
rect 3159 2562 3163 2563
rect 3159 2557 3163 2558
rect 3271 2562 3275 2563
rect 3271 2557 3275 2558
rect 3367 2562 3371 2563
rect 3367 2557 3371 2558
rect 3463 2562 3467 2563
rect 3463 2557 3467 2558
rect 1670 2547 1676 2548
rect 1766 2549 1772 2550
rect 110 2544 116 2545
rect 1766 2545 1767 2549
rect 1771 2545 1772 2549
rect 1766 2544 1772 2545
rect 1808 2541 1810 2557
rect 1806 2540 1812 2541
rect 2208 2540 2210 2557
rect 2800 2540 2802 2557
rect 3368 2540 3370 2557
rect 3464 2541 3466 2557
rect 3462 2540 3468 2541
rect 1806 2536 1807 2540
rect 1811 2536 1812 2540
rect 1806 2535 1812 2536
rect 2206 2539 2212 2540
rect 2206 2535 2207 2539
rect 2211 2535 2212 2539
rect 2206 2534 2212 2535
rect 2798 2539 2804 2540
rect 2798 2535 2799 2539
rect 2803 2535 2804 2539
rect 2798 2534 2804 2535
rect 3366 2539 3372 2540
rect 3366 2535 3367 2539
rect 3371 2535 3372 2539
rect 3462 2536 3463 2540
rect 3467 2536 3468 2540
rect 3462 2535 3468 2536
rect 3366 2534 3372 2535
rect 222 2533 228 2534
rect 110 2532 116 2533
rect 110 2528 111 2532
rect 115 2528 116 2532
rect 222 2529 223 2533
rect 227 2529 228 2533
rect 222 2528 228 2529
rect 310 2533 316 2534
rect 310 2529 311 2533
rect 315 2529 316 2533
rect 310 2528 316 2529
rect 406 2533 412 2534
rect 406 2529 407 2533
rect 411 2529 412 2533
rect 406 2528 412 2529
rect 502 2533 508 2534
rect 502 2529 503 2533
rect 507 2529 508 2533
rect 502 2528 508 2529
rect 590 2533 596 2534
rect 590 2529 591 2533
rect 595 2529 596 2533
rect 590 2528 596 2529
rect 678 2533 684 2534
rect 678 2529 679 2533
rect 683 2529 684 2533
rect 678 2528 684 2529
rect 766 2533 772 2534
rect 766 2529 767 2533
rect 771 2529 772 2533
rect 766 2528 772 2529
rect 854 2533 860 2534
rect 854 2529 855 2533
rect 859 2529 860 2533
rect 854 2528 860 2529
rect 942 2533 948 2534
rect 942 2529 943 2533
rect 947 2529 948 2533
rect 942 2528 948 2529
rect 1030 2533 1036 2534
rect 1030 2529 1031 2533
rect 1035 2529 1036 2533
rect 1030 2528 1036 2529
rect 1118 2533 1124 2534
rect 1118 2529 1119 2533
rect 1123 2529 1124 2533
rect 1118 2528 1124 2529
rect 1214 2533 1220 2534
rect 1214 2529 1215 2533
rect 1219 2529 1220 2533
rect 1214 2528 1220 2529
rect 1310 2533 1316 2534
rect 1310 2529 1311 2533
rect 1315 2529 1316 2533
rect 1310 2528 1316 2529
rect 1406 2533 1412 2534
rect 1406 2529 1407 2533
rect 1411 2529 1412 2533
rect 1406 2528 1412 2529
rect 1494 2533 1500 2534
rect 1494 2529 1495 2533
rect 1499 2529 1500 2533
rect 1494 2528 1500 2529
rect 1582 2533 1588 2534
rect 1582 2529 1583 2533
rect 1587 2529 1588 2533
rect 1582 2528 1588 2529
rect 1670 2533 1676 2534
rect 1670 2529 1671 2533
rect 1675 2529 1676 2533
rect 1670 2528 1676 2529
rect 1766 2532 1772 2533
rect 1766 2528 1767 2532
rect 1771 2528 1772 2532
rect 110 2527 116 2528
rect 112 2511 114 2527
rect 224 2511 226 2528
rect 312 2511 314 2528
rect 408 2511 410 2528
rect 504 2511 506 2528
rect 592 2511 594 2528
rect 680 2511 682 2528
rect 768 2511 770 2528
rect 856 2511 858 2528
rect 944 2511 946 2528
rect 1032 2511 1034 2528
rect 1120 2511 1122 2528
rect 1216 2511 1218 2528
rect 1312 2511 1314 2528
rect 1408 2511 1410 2528
rect 1496 2511 1498 2528
rect 1584 2511 1586 2528
rect 1672 2511 1674 2528
rect 1766 2527 1772 2528
rect 1768 2511 1770 2527
rect 1806 2523 1812 2524
rect 1806 2519 1807 2523
rect 1811 2519 1812 2523
rect 3462 2523 3468 2524
rect 1806 2518 1812 2519
rect 2206 2520 2212 2521
rect 111 2510 115 2511
rect 111 2505 115 2506
rect 135 2510 139 2511
rect 135 2505 139 2506
rect 223 2510 227 2511
rect 223 2505 227 2506
rect 247 2510 251 2511
rect 247 2505 251 2506
rect 311 2510 315 2511
rect 311 2505 315 2506
rect 391 2510 395 2511
rect 391 2505 395 2506
rect 407 2510 411 2511
rect 407 2505 411 2506
rect 503 2510 507 2511
rect 503 2505 507 2506
rect 543 2510 547 2511
rect 543 2505 547 2506
rect 591 2510 595 2511
rect 591 2505 595 2506
rect 679 2510 683 2511
rect 679 2505 683 2506
rect 695 2510 699 2511
rect 695 2505 699 2506
rect 767 2510 771 2511
rect 767 2505 771 2506
rect 839 2510 843 2511
rect 839 2505 843 2506
rect 855 2510 859 2511
rect 855 2505 859 2506
rect 943 2510 947 2511
rect 943 2505 947 2506
rect 975 2510 979 2511
rect 975 2505 979 2506
rect 1031 2510 1035 2511
rect 1031 2505 1035 2506
rect 1103 2510 1107 2511
rect 1103 2505 1107 2506
rect 1119 2510 1123 2511
rect 1119 2505 1123 2506
rect 1215 2510 1219 2511
rect 1215 2505 1219 2506
rect 1231 2510 1235 2511
rect 1231 2505 1235 2506
rect 1311 2510 1315 2511
rect 1311 2505 1315 2506
rect 1351 2510 1355 2511
rect 1351 2505 1355 2506
rect 1407 2510 1411 2511
rect 1407 2505 1411 2506
rect 1463 2510 1467 2511
rect 1463 2505 1467 2506
rect 1495 2510 1499 2511
rect 1495 2505 1499 2506
rect 1575 2510 1579 2511
rect 1575 2505 1579 2506
rect 1583 2510 1587 2511
rect 1583 2505 1587 2506
rect 1671 2510 1675 2511
rect 1671 2505 1675 2506
rect 1767 2510 1771 2511
rect 1767 2505 1771 2506
rect 112 2489 114 2505
rect 110 2488 116 2489
rect 136 2488 138 2505
rect 248 2488 250 2505
rect 392 2488 394 2505
rect 544 2488 546 2505
rect 696 2488 698 2505
rect 840 2488 842 2505
rect 976 2488 978 2505
rect 1104 2488 1106 2505
rect 1232 2488 1234 2505
rect 1352 2488 1354 2505
rect 1464 2488 1466 2505
rect 1576 2488 1578 2505
rect 1672 2488 1674 2505
rect 1768 2489 1770 2505
rect 1766 2488 1772 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 134 2487 140 2488
rect 134 2483 135 2487
rect 139 2483 140 2487
rect 134 2482 140 2483
rect 246 2487 252 2488
rect 246 2483 247 2487
rect 251 2483 252 2487
rect 246 2482 252 2483
rect 390 2487 396 2488
rect 390 2483 391 2487
rect 395 2483 396 2487
rect 390 2482 396 2483
rect 542 2487 548 2488
rect 542 2483 543 2487
rect 547 2483 548 2487
rect 542 2482 548 2483
rect 694 2487 700 2488
rect 694 2483 695 2487
rect 699 2483 700 2487
rect 694 2482 700 2483
rect 838 2487 844 2488
rect 838 2483 839 2487
rect 843 2483 844 2487
rect 838 2482 844 2483
rect 974 2487 980 2488
rect 974 2483 975 2487
rect 979 2483 980 2487
rect 974 2482 980 2483
rect 1102 2487 1108 2488
rect 1102 2483 1103 2487
rect 1107 2483 1108 2487
rect 1102 2482 1108 2483
rect 1230 2487 1236 2488
rect 1230 2483 1231 2487
rect 1235 2483 1236 2487
rect 1230 2482 1236 2483
rect 1350 2487 1356 2488
rect 1350 2483 1351 2487
rect 1355 2483 1356 2487
rect 1350 2482 1356 2483
rect 1462 2487 1468 2488
rect 1462 2483 1463 2487
rect 1467 2483 1468 2487
rect 1462 2482 1468 2483
rect 1574 2487 1580 2488
rect 1574 2483 1575 2487
rect 1579 2483 1580 2487
rect 1574 2482 1580 2483
rect 1670 2487 1676 2488
rect 1670 2483 1671 2487
rect 1675 2483 1676 2487
rect 1766 2484 1767 2488
rect 1771 2484 1772 2488
rect 1766 2483 1772 2484
rect 1808 2483 1810 2518
rect 2206 2516 2207 2520
rect 2211 2516 2212 2520
rect 2206 2515 2212 2516
rect 2798 2520 2804 2521
rect 2798 2516 2799 2520
rect 2803 2516 2804 2520
rect 2798 2515 2804 2516
rect 3366 2520 3372 2521
rect 3366 2516 3367 2520
rect 3371 2516 3372 2520
rect 3462 2519 3463 2523
rect 3467 2519 3468 2523
rect 3462 2518 3468 2519
rect 3366 2515 3372 2516
rect 2208 2483 2210 2515
rect 2800 2483 2802 2515
rect 3368 2483 3370 2515
rect 3464 2483 3466 2518
rect 1670 2482 1676 2483
rect 1807 2482 1811 2483
rect 1807 2477 1811 2478
rect 2015 2482 2019 2483
rect 2015 2477 2019 2478
rect 2199 2482 2203 2483
rect 2199 2477 2203 2478
rect 2207 2482 2211 2483
rect 2207 2477 2211 2478
rect 2367 2482 2371 2483
rect 2367 2477 2371 2478
rect 2527 2482 2531 2483
rect 2527 2477 2531 2478
rect 2671 2482 2675 2483
rect 2671 2477 2675 2478
rect 2799 2482 2803 2483
rect 2799 2477 2803 2478
rect 2807 2482 2811 2483
rect 2807 2477 2811 2478
rect 2927 2482 2931 2483
rect 2927 2477 2931 2478
rect 3047 2482 3051 2483
rect 3047 2477 3051 2478
rect 3159 2482 3163 2483
rect 3159 2477 3163 2478
rect 3271 2482 3275 2483
rect 3271 2477 3275 2478
rect 3367 2482 3371 2483
rect 3367 2477 3371 2478
rect 3463 2482 3467 2483
rect 3463 2477 3467 2478
rect 110 2471 116 2472
rect 110 2467 111 2471
rect 115 2467 116 2471
rect 1766 2471 1772 2472
rect 110 2466 116 2467
rect 134 2468 140 2469
rect 112 2431 114 2466
rect 134 2464 135 2468
rect 139 2464 140 2468
rect 134 2463 140 2464
rect 246 2468 252 2469
rect 246 2464 247 2468
rect 251 2464 252 2468
rect 246 2463 252 2464
rect 390 2468 396 2469
rect 390 2464 391 2468
rect 395 2464 396 2468
rect 390 2463 396 2464
rect 542 2468 548 2469
rect 542 2464 543 2468
rect 547 2464 548 2468
rect 542 2463 548 2464
rect 694 2468 700 2469
rect 694 2464 695 2468
rect 699 2464 700 2468
rect 694 2463 700 2464
rect 838 2468 844 2469
rect 838 2464 839 2468
rect 843 2464 844 2468
rect 838 2463 844 2464
rect 974 2468 980 2469
rect 974 2464 975 2468
rect 979 2464 980 2468
rect 974 2463 980 2464
rect 1102 2468 1108 2469
rect 1102 2464 1103 2468
rect 1107 2464 1108 2468
rect 1102 2463 1108 2464
rect 1230 2468 1236 2469
rect 1230 2464 1231 2468
rect 1235 2464 1236 2468
rect 1230 2463 1236 2464
rect 1350 2468 1356 2469
rect 1350 2464 1351 2468
rect 1355 2464 1356 2468
rect 1350 2463 1356 2464
rect 1462 2468 1468 2469
rect 1462 2464 1463 2468
rect 1467 2464 1468 2468
rect 1462 2463 1468 2464
rect 1574 2468 1580 2469
rect 1574 2464 1575 2468
rect 1579 2464 1580 2468
rect 1574 2463 1580 2464
rect 1670 2468 1676 2469
rect 1670 2464 1671 2468
rect 1675 2464 1676 2468
rect 1766 2467 1767 2471
rect 1771 2467 1772 2471
rect 1766 2466 1772 2467
rect 1670 2463 1676 2464
rect 136 2431 138 2463
rect 248 2431 250 2463
rect 392 2431 394 2463
rect 544 2431 546 2463
rect 696 2431 698 2463
rect 840 2431 842 2463
rect 976 2431 978 2463
rect 1104 2431 1106 2463
rect 1232 2431 1234 2463
rect 1352 2431 1354 2463
rect 1464 2431 1466 2463
rect 1576 2431 1578 2463
rect 1672 2431 1674 2463
rect 1768 2431 1770 2466
rect 1808 2458 1810 2477
rect 2016 2461 2018 2477
rect 2200 2461 2202 2477
rect 2368 2461 2370 2477
rect 2528 2461 2530 2477
rect 2672 2461 2674 2477
rect 2808 2461 2810 2477
rect 2928 2461 2930 2477
rect 3048 2461 3050 2477
rect 3160 2461 3162 2477
rect 3272 2461 3274 2477
rect 3368 2461 3370 2477
rect 2014 2460 2020 2461
rect 1806 2457 1812 2458
rect 1806 2453 1807 2457
rect 1811 2453 1812 2457
rect 2014 2456 2015 2460
rect 2019 2456 2020 2460
rect 2014 2455 2020 2456
rect 2198 2460 2204 2461
rect 2198 2456 2199 2460
rect 2203 2456 2204 2460
rect 2198 2455 2204 2456
rect 2366 2460 2372 2461
rect 2366 2456 2367 2460
rect 2371 2456 2372 2460
rect 2366 2455 2372 2456
rect 2526 2460 2532 2461
rect 2526 2456 2527 2460
rect 2531 2456 2532 2460
rect 2526 2455 2532 2456
rect 2670 2460 2676 2461
rect 2670 2456 2671 2460
rect 2675 2456 2676 2460
rect 2670 2455 2676 2456
rect 2806 2460 2812 2461
rect 2806 2456 2807 2460
rect 2811 2456 2812 2460
rect 2806 2455 2812 2456
rect 2926 2460 2932 2461
rect 2926 2456 2927 2460
rect 2931 2456 2932 2460
rect 2926 2455 2932 2456
rect 3046 2460 3052 2461
rect 3046 2456 3047 2460
rect 3051 2456 3052 2460
rect 3046 2455 3052 2456
rect 3158 2460 3164 2461
rect 3158 2456 3159 2460
rect 3163 2456 3164 2460
rect 3158 2455 3164 2456
rect 3270 2460 3276 2461
rect 3270 2456 3271 2460
rect 3275 2456 3276 2460
rect 3270 2455 3276 2456
rect 3366 2460 3372 2461
rect 3366 2456 3367 2460
rect 3371 2456 3372 2460
rect 3464 2458 3466 2477
rect 3366 2455 3372 2456
rect 3462 2457 3468 2458
rect 1806 2452 1812 2453
rect 3462 2453 3463 2457
rect 3467 2453 3468 2457
rect 3462 2452 3468 2453
rect 2014 2441 2020 2442
rect 1806 2440 1812 2441
rect 1806 2436 1807 2440
rect 1811 2436 1812 2440
rect 2014 2437 2015 2441
rect 2019 2437 2020 2441
rect 2014 2436 2020 2437
rect 2198 2441 2204 2442
rect 2198 2437 2199 2441
rect 2203 2437 2204 2441
rect 2198 2436 2204 2437
rect 2366 2441 2372 2442
rect 2366 2437 2367 2441
rect 2371 2437 2372 2441
rect 2366 2436 2372 2437
rect 2526 2441 2532 2442
rect 2526 2437 2527 2441
rect 2531 2437 2532 2441
rect 2526 2436 2532 2437
rect 2670 2441 2676 2442
rect 2670 2437 2671 2441
rect 2675 2437 2676 2441
rect 2670 2436 2676 2437
rect 2806 2441 2812 2442
rect 2806 2437 2807 2441
rect 2811 2437 2812 2441
rect 2806 2436 2812 2437
rect 2926 2441 2932 2442
rect 2926 2437 2927 2441
rect 2931 2437 2932 2441
rect 2926 2436 2932 2437
rect 3046 2441 3052 2442
rect 3046 2437 3047 2441
rect 3051 2437 3052 2441
rect 3046 2436 3052 2437
rect 3158 2441 3164 2442
rect 3158 2437 3159 2441
rect 3163 2437 3164 2441
rect 3158 2436 3164 2437
rect 3270 2441 3276 2442
rect 3270 2437 3271 2441
rect 3275 2437 3276 2441
rect 3270 2436 3276 2437
rect 3366 2441 3372 2442
rect 3366 2437 3367 2441
rect 3371 2437 3372 2441
rect 3366 2436 3372 2437
rect 3462 2440 3468 2441
rect 3462 2436 3463 2440
rect 3467 2436 3468 2440
rect 1806 2435 1812 2436
rect 111 2430 115 2431
rect 111 2425 115 2426
rect 135 2430 139 2431
rect 135 2425 139 2426
rect 239 2430 243 2431
rect 239 2425 243 2426
rect 247 2430 251 2431
rect 247 2425 251 2426
rect 391 2430 395 2431
rect 391 2425 395 2426
rect 543 2430 547 2431
rect 543 2425 547 2426
rect 551 2430 555 2431
rect 551 2425 555 2426
rect 695 2430 699 2431
rect 695 2425 699 2426
rect 719 2430 723 2431
rect 719 2425 723 2426
rect 839 2430 843 2431
rect 839 2425 843 2426
rect 895 2430 899 2431
rect 895 2425 899 2426
rect 975 2430 979 2431
rect 975 2425 979 2426
rect 1063 2430 1067 2431
rect 1063 2425 1067 2426
rect 1103 2430 1107 2431
rect 1103 2425 1107 2426
rect 1231 2430 1235 2431
rect 1231 2425 1235 2426
rect 1239 2430 1243 2431
rect 1239 2425 1243 2426
rect 1351 2430 1355 2431
rect 1351 2425 1355 2426
rect 1415 2430 1419 2431
rect 1415 2425 1419 2426
rect 1463 2430 1467 2431
rect 1463 2425 1467 2426
rect 1575 2430 1579 2431
rect 1575 2425 1579 2426
rect 1591 2430 1595 2431
rect 1591 2425 1595 2426
rect 1671 2430 1675 2431
rect 1671 2425 1675 2426
rect 1767 2430 1771 2431
rect 1767 2425 1771 2426
rect 112 2406 114 2425
rect 136 2409 138 2425
rect 240 2409 242 2425
rect 392 2409 394 2425
rect 552 2409 554 2425
rect 720 2409 722 2425
rect 896 2409 898 2425
rect 1064 2409 1066 2425
rect 1240 2409 1242 2425
rect 1416 2409 1418 2425
rect 1592 2409 1594 2425
rect 134 2408 140 2409
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 134 2404 135 2408
rect 139 2404 140 2408
rect 134 2403 140 2404
rect 238 2408 244 2409
rect 238 2404 239 2408
rect 243 2404 244 2408
rect 238 2403 244 2404
rect 390 2408 396 2409
rect 390 2404 391 2408
rect 395 2404 396 2408
rect 390 2403 396 2404
rect 550 2408 556 2409
rect 550 2404 551 2408
rect 555 2404 556 2408
rect 550 2403 556 2404
rect 718 2408 724 2409
rect 718 2404 719 2408
rect 723 2404 724 2408
rect 718 2403 724 2404
rect 894 2408 900 2409
rect 894 2404 895 2408
rect 899 2404 900 2408
rect 894 2403 900 2404
rect 1062 2408 1068 2409
rect 1062 2404 1063 2408
rect 1067 2404 1068 2408
rect 1062 2403 1068 2404
rect 1238 2408 1244 2409
rect 1238 2404 1239 2408
rect 1243 2404 1244 2408
rect 1238 2403 1244 2404
rect 1414 2408 1420 2409
rect 1414 2404 1415 2408
rect 1419 2404 1420 2408
rect 1414 2403 1420 2404
rect 1590 2408 1596 2409
rect 1590 2404 1591 2408
rect 1595 2404 1596 2408
rect 1768 2406 1770 2425
rect 1808 2415 1810 2435
rect 2016 2415 2018 2436
rect 2200 2415 2202 2436
rect 2368 2415 2370 2436
rect 2528 2415 2530 2436
rect 2672 2415 2674 2436
rect 2808 2415 2810 2436
rect 2928 2415 2930 2436
rect 3048 2415 3050 2436
rect 3160 2415 3162 2436
rect 3272 2415 3274 2436
rect 3368 2415 3370 2436
rect 3462 2435 3468 2436
rect 3464 2415 3466 2435
rect 1807 2414 1811 2415
rect 1807 2409 1811 2410
rect 1839 2414 1843 2415
rect 1839 2409 1843 2410
rect 2007 2414 2011 2415
rect 2007 2409 2011 2410
rect 2015 2414 2019 2415
rect 2015 2409 2019 2410
rect 2183 2414 2187 2415
rect 2183 2409 2187 2410
rect 2199 2414 2203 2415
rect 2199 2409 2203 2410
rect 2367 2414 2371 2415
rect 2367 2409 2371 2410
rect 2527 2414 2531 2415
rect 2527 2409 2531 2410
rect 2559 2414 2563 2415
rect 2559 2409 2563 2410
rect 2671 2414 2675 2415
rect 2671 2409 2675 2410
rect 2759 2414 2763 2415
rect 2759 2409 2763 2410
rect 2807 2414 2811 2415
rect 2807 2409 2811 2410
rect 2927 2414 2931 2415
rect 2927 2409 2931 2410
rect 2967 2414 2971 2415
rect 2967 2409 2971 2410
rect 3047 2414 3051 2415
rect 3047 2409 3051 2410
rect 3159 2414 3163 2415
rect 3159 2409 3163 2410
rect 3175 2414 3179 2415
rect 3175 2409 3179 2410
rect 3271 2414 3275 2415
rect 3271 2409 3275 2410
rect 3367 2414 3371 2415
rect 3367 2409 3371 2410
rect 3463 2414 3467 2415
rect 3463 2409 3467 2410
rect 1590 2403 1596 2404
rect 1766 2405 1772 2406
rect 110 2400 116 2401
rect 1766 2401 1767 2405
rect 1771 2401 1772 2405
rect 1766 2400 1772 2401
rect 1808 2393 1810 2409
rect 1806 2392 1812 2393
rect 1840 2392 1842 2409
rect 2008 2392 2010 2409
rect 2184 2392 2186 2409
rect 2368 2392 2370 2409
rect 2560 2392 2562 2409
rect 2760 2392 2762 2409
rect 2968 2392 2970 2409
rect 3176 2392 3178 2409
rect 3368 2392 3370 2409
rect 3464 2393 3466 2409
rect 3462 2392 3468 2393
rect 134 2389 140 2390
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 134 2385 135 2389
rect 139 2385 140 2389
rect 134 2384 140 2385
rect 238 2389 244 2390
rect 238 2385 239 2389
rect 243 2385 244 2389
rect 238 2384 244 2385
rect 390 2389 396 2390
rect 390 2385 391 2389
rect 395 2385 396 2389
rect 390 2384 396 2385
rect 550 2389 556 2390
rect 550 2385 551 2389
rect 555 2385 556 2389
rect 550 2384 556 2385
rect 718 2389 724 2390
rect 718 2385 719 2389
rect 723 2385 724 2389
rect 718 2384 724 2385
rect 894 2389 900 2390
rect 894 2385 895 2389
rect 899 2385 900 2389
rect 894 2384 900 2385
rect 1062 2389 1068 2390
rect 1062 2385 1063 2389
rect 1067 2385 1068 2389
rect 1062 2384 1068 2385
rect 1238 2389 1244 2390
rect 1238 2385 1239 2389
rect 1243 2385 1244 2389
rect 1238 2384 1244 2385
rect 1414 2389 1420 2390
rect 1414 2385 1415 2389
rect 1419 2385 1420 2389
rect 1414 2384 1420 2385
rect 1590 2389 1596 2390
rect 1590 2385 1591 2389
rect 1595 2385 1596 2389
rect 1590 2384 1596 2385
rect 1766 2388 1772 2389
rect 1766 2384 1767 2388
rect 1771 2384 1772 2388
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1838 2391 1844 2392
rect 1838 2387 1839 2391
rect 1843 2387 1844 2391
rect 1838 2386 1844 2387
rect 2006 2391 2012 2392
rect 2006 2387 2007 2391
rect 2011 2387 2012 2391
rect 2006 2386 2012 2387
rect 2182 2391 2188 2392
rect 2182 2387 2183 2391
rect 2187 2387 2188 2391
rect 2182 2386 2188 2387
rect 2366 2391 2372 2392
rect 2366 2387 2367 2391
rect 2371 2387 2372 2391
rect 2366 2386 2372 2387
rect 2558 2391 2564 2392
rect 2558 2387 2559 2391
rect 2563 2387 2564 2391
rect 2558 2386 2564 2387
rect 2758 2391 2764 2392
rect 2758 2387 2759 2391
rect 2763 2387 2764 2391
rect 2758 2386 2764 2387
rect 2966 2391 2972 2392
rect 2966 2387 2967 2391
rect 2971 2387 2972 2391
rect 2966 2386 2972 2387
rect 3174 2391 3180 2392
rect 3174 2387 3175 2391
rect 3179 2387 3180 2391
rect 3174 2386 3180 2387
rect 3366 2391 3372 2392
rect 3366 2387 3367 2391
rect 3371 2387 3372 2391
rect 3462 2388 3463 2392
rect 3467 2388 3468 2392
rect 3462 2387 3468 2388
rect 3366 2386 3372 2387
rect 110 2383 116 2384
rect 112 2359 114 2383
rect 136 2359 138 2384
rect 240 2359 242 2384
rect 392 2359 394 2384
rect 552 2359 554 2384
rect 720 2359 722 2384
rect 896 2359 898 2384
rect 1064 2359 1066 2384
rect 1240 2359 1242 2384
rect 1416 2359 1418 2384
rect 1592 2359 1594 2384
rect 1766 2383 1772 2384
rect 1768 2359 1770 2383
rect 1806 2375 1812 2376
rect 1806 2371 1807 2375
rect 1811 2371 1812 2375
rect 3462 2375 3468 2376
rect 1806 2370 1812 2371
rect 1838 2372 1844 2373
rect 111 2358 115 2359
rect 111 2353 115 2354
rect 135 2358 139 2359
rect 135 2353 139 2354
rect 239 2358 243 2359
rect 239 2353 243 2354
rect 375 2358 379 2359
rect 375 2353 379 2354
rect 391 2358 395 2359
rect 391 2353 395 2354
rect 479 2358 483 2359
rect 479 2353 483 2354
rect 551 2358 555 2359
rect 551 2353 555 2354
rect 599 2358 603 2359
rect 599 2353 603 2354
rect 719 2358 723 2359
rect 719 2353 723 2354
rect 847 2358 851 2359
rect 847 2353 851 2354
rect 895 2358 899 2359
rect 895 2353 899 2354
rect 975 2358 979 2359
rect 975 2353 979 2354
rect 1063 2358 1067 2359
rect 1063 2353 1067 2354
rect 1103 2358 1107 2359
rect 1103 2353 1107 2354
rect 1239 2358 1243 2359
rect 1239 2353 1243 2354
rect 1375 2358 1379 2359
rect 1375 2353 1379 2354
rect 1415 2358 1419 2359
rect 1415 2353 1419 2354
rect 1511 2358 1515 2359
rect 1511 2353 1515 2354
rect 1591 2358 1595 2359
rect 1591 2353 1595 2354
rect 1767 2358 1771 2359
rect 1767 2353 1771 2354
rect 112 2337 114 2353
rect 110 2336 116 2337
rect 376 2336 378 2353
rect 480 2336 482 2353
rect 600 2336 602 2353
rect 720 2336 722 2353
rect 848 2336 850 2353
rect 976 2336 978 2353
rect 1104 2336 1106 2353
rect 1240 2336 1242 2353
rect 1376 2336 1378 2353
rect 1512 2336 1514 2353
rect 1768 2337 1770 2353
rect 1808 2351 1810 2370
rect 1838 2368 1839 2372
rect 1843 2368 1844 2372
rect 1838 2367 1844 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2182 2372 2188 2373
rect 2182 2368 2183 2372
rect 2187 2368 2188 2372
rect 2182 2367 2188 2368
rect 2366 2372 2372 2373
rect 2366 2368 2367 2372
rect 2371 2368 2372 2372
rect 2366 2367 2372 2368
rect 2558 2372 2564 2373
rect 2558 2368 2559 2372
rect 2563 2368 2564 2372
rect 2558 2367 2564 2368
rect 2758 2372 2764 2373
rect 2758 2368 2759 2372
rect 2763 2368 2764 2372
rect 2758 2367 2764 2368
rect 2966 2372 2972 2373
rect 2966 2368 2967 2372
rect 2971 2368 2972 2372
rect 2966 2367 2972 2368
rect 3174 2372 3180 2373
rect 3174 2368 3175 2372
rect 3179 2368 3180 2372
rect 3174 2367 3180 2368
rect 3366 2372 3372 2373
rect 3366 2368 3367 2372
rect 3371 2368 3372 2372
rect 3462 2371 3463 2375
rect 3467 2371 3468 2375
rect 3462 2370 3468 2371
rect 3366 2367 3372 2368
rect 1840 2351 1842 2367
rect 2008 2351 2010 2367
rect 2184 2351 2186 2367
rect 2368 2351 2370 2367
rect 2560 2351 2562 2367
rect 2760 2351 2762 2367
rect 2968 2351 2970 2367
rect 3176 2351 3178 2367
rect 3368 2351 3370 2367
rect 3464 2351 3466 2370
rect 1807 2350 1811 2351
rect 1807 2345 1811 2346
rect 1839 2350 1843 2351
rect 1839 2345 1843 2346
rect 1887 2350 1891 2351
rect 1887 2345 1891 2346
rect 2007 2350 2011 2351
rect 2007 2345 2011 2346
rect 2015 2350 2019 2351
rect 2015 2345 2019 2346
rect 2151 2350 2155 2351
rect 2151 2345 2155 2346
rect 2183 2350 2187 2351
rect 2183 2345 2187 2346
rect 2303 2350 2307 2351
rect 2303 2345 2307 2346
rect 2367 2350 2371 2351
rect 2367 2345 2371 2346
rect 2463 2350 2467 2351
rect 2463 2345 2467 2346
rect 2559 2350 2563 2351
rect 2559 2345 2563 2346
rect 2647 2350 2651 2351
rect 2647 2345 2651 2346
rect 2759 2350 2763 2351
rect 2759 2345 2763 2346
rect 2839 2350 2843 2351
rect 2839 2345 2843 2346
rect 2967 2350 2971 2351
rect 2967 2345 2971 2346
rect 3047 2350 3051 2351
rect 3047 2345 3051 2346
rect 3175 2350 3179 2351
rect 3175 2345 3179 2346
rect 3255 2350 3259 2351
rect 3255 2345 3259 2346
rect 3367 2350 3371 2351
rect 3367 2345 3371 2346
rect 3463 2350 3467 2351
rect 3463 2345 3467 2346
rect 1766 2336 1772 2337
rect 110 2332 111 2336
rect 115 2332 116 2336
rect 110 2331 116 2332
rect 374 2335 380 2336
rect 374 2331 375 2335
rect 379 2331 380 2335
rect 374 2330 380 2331
rect 478 2335 484 2336
rect 478 2331 479 2335
rect 483 2331 484 2335
rect 478 2330 484 2331
rect 598 2335 604 2336
rect 598 2331 599 2335
rect 603 2331 604 2335
rect 598 2330 604 2331
rect 718 2335 724 2336
rect 718 2331 719 2335
rect 723 2331 724 2335
rect 718 2330 724 2331
rect 846 2335 852 2336
rect 846 2331 847 2335
rect 851 2331 852 2335
rect 846 2330 852 2331
rect 974 2335 980 2336
rect 974 2331 975 2335
rect 979 2331 980 2335
rect 974 2330 980 2331
rect 1102 2335 1108 2336
rect 1102 2331 1103 2335
rect 1107 2331 1108 2335
rect 1102 2330 1108 2331
rect 1238 2335 1244 2336
rect 1238 2331 1239 2335
rect 1243 2331 1244 2335
rect 1238 2330 1244 2331
rect 1374 2335 1380 2336
rect 1374 2331 1375 2335
rect 1379 2331 1380 2335
rect 1374 2330 1380 2331
rect 1510 2335 1516 2336
rect 1510 2331 1511 2335
rect 1515 2331 1516 2335
rect 1766 2332 1767 2336
rect 1771 2332 1772 2336
rect 1766 2331 1772 2332
rect 1510 2330 1516 2331
rect 1808 2326 1810 2345
rect 1888 2329 1890 2345
rect 2016 2329 2018 2345
rect 2152 2329 2154 2345
rect 2304 2329 2306 2345
rect 2464 2329 2466 2345
rect 2648 2329 2650 2345
rect 2840 2329 2842 2345
rect 3048 2329 3050 2345
rect 3256 2329 3258 2345
rect 1886 2328 1892 2329
rect 1806 2325 1812 2326
rect 1806 2321 1807 2325
rect 1811 2321 1812 2325
rect 1886 2324 1887 2328
rect 1891 2324 1892 2328
rect 1886 2323 1892 2324
rect 2014 2328 2020 2329
rect 2014 2324 2015 2328
rect 2019 2324 2020 2328
rect 2014 2323 2020 2324
rect 2150 2328 2156 2329
rect 2150 2324 2151 2328
rect 2155 2324 2156 2328
rect 2150 2323 2156 2324
rect 2302 2328 2308 2329
rect 2302 2324 2303 2328
rect 2307 2324 2308 2328
rect 2302 2323 2308 2324
rect 2462 2328 2468 2329
rect 2462 2324 2463 2328
rect 2467 2324 2468 2328
rect 2462 2323 2468 2324
rect 2646 2328 2652 2329
rect 2646 2324 2647 2328
rect 2651 2324 2652 2328
rect 2646 2323 2652 2324
rect 2838 2328 2844 2329
rect 2838 2324 2839 2328
rect 2843 2324 2844 2328
rect 2838 2323 2844 2324
rect 3046 2328 3052 2329
rect 3046 2324 3047 2328
rect 3051 2324 3052 2328
rect 3046 2323 3052 2324
rect 3254 2328 3260 2329
rect 3254 2324 3255 2328
rect 3259 2324 3260 2328
rect 3464 2326 3466 2345
rect 3254 2323 3260 2324
rect 3462 2325 3468 2326
rect 1806 2320 1812 2321
rect 3462 2321 3463 2325
rect 3467 2321 3468 2325
rect 3462 2320 3468 2321
rect 110 2319 116 2320
rect 110 2315 111 2319
rect 115 2315 116 2319
rect 1766 2319 1772 2320
rect 110 2314 116 2315
rect 374 2316 380 2317
rect 112 2287 114 2314
rect 374 2312 375 2316
rect 379 2312 380 2316
rect 374 2311 380 2312
rect 478 2316 484 2317
rect 478 2312 479 2316
rect 483 2312 484 2316
rect 478 2311 484 2312
rect 598 2316 604 2317
rect 598 2312 599 2316
rect 603 2312 604 2316
rect 598 2311 604 2312
rect 718 2316 724 2317
rect 718 2312 719 2316
rect 723 2312 724 2316
rect 718 2311 724 2312
rect 846 2316 852 2317
rect 846 2312 847 2316
rect 851 2312 852 2316
rect 846 2311 852 2312
rect 974 2316 980 2317
rect 974 2312 975 2316
rect 979 2312 980 2316
rect 974 2311 980 2312
rect 1102 2316 1108 2317
rect 1102 2312 1103 2316
rect 1107 2312 1108 2316
rect 1102 2311 1108 2312
rect 1238 2316 1244 2317
rect 1238 2312 1239 2316
rect 1243 2312 1244 2316
rect 1238 2311 1244 2312
rect 1374 2316 1380 2317
rect 1374 2312 1375 2316
rect 1379 2312 1380 2316
rect 1374 2311 1380 2312
rect 1510 2316 1516 2317
rect 1510 2312 1511 2316
rect 1515 2312 1516 2316
rect 1766 2315 1767 2319
rect 1771 2315 1772 2319
rect 1766 2314 1772 2315
rect 1510 2311 1516 2312
rect 376 2287 378 2311
rect 480 2287 482 2311
rect 600 2287 602 2311
rect 720 2287 722 2311
rect 848 2287 850 2311
rect 976 2287 978 2311
rect 1104 2287 1106 2311
rect 1240 2287 1242 2311
rect 1376 2287 1378 2311
rect 1512 2287 1514 2311
rect 1768 2287 1770 2314
rect 1886 2309 1892 2310
rect 1806 2308 1812 2309
rect 1806 2304 1807 2308
rect 1811 2304 1812 2308
rect 1886 2305 1887 2309
rect 1891 2305 1892 2309
rect 1886 2304 1892 2305
rect 2014 2309 2020 2310
rect 2014 2305 2015 2309
rect 2019 2305 2020 2309
rect 2014 2304 2020 2305
rect 2150 2309 2156 2310
rect 2150 2305 2151 2309
rect 2155 2305 2156 2309
rect 2150 2304 2156 2305
rect 2302 2309 2308 2310
rect 2302 2305 2303 2309
rect 2307 2305 2308 2309
rect 2302 2304 2308 2305
rect 2462 2309 2468 2310
rect 2462 2305 2463 2309
rect 2467 2305 2468 2309
rect 2462 2304 2468 2305
rect 2646 2309 2652 2310
rect 2646 2305 2647 2309
rect 2651 2305 2652 2309
rect 2646 2304 2652 2305
rect 2838 2309 2844 2310
rect 2838 2305 2839 2309
rect 2843 2305 2844 2309
rect 2838 2304 2844 2305
rect 3046 2309 3052 2310
rect 3046 2305 3047 2309
rect 3051 2305 3052 2309
rect 3046 2304 3052 2305
rect 3254 2309 3260 2310
rect 3254 2305 3255 2309
rect 3259 2305 3260 2309
rect 3254 2304 3260 2305
rect 3462 2308 3468 2309
rect 3462 2304 3463 2308
rect 3467 2304 3468 2308
rect 1806 2303 1812 2304
rect 111 2286 115 2287
rect 111 2281 115 2282
rect 375 2286 379 2287
rect 375 2281 379 2282
rect 479 2286 483 2287
rect 479 2281 483 2282
rect 575 2286 579 2287
rect 575 2281 579 2282
rect 599 2286 603 2287
rect 599 2281 603 2282
rect 663 2286 667 2287
rect 663 2281 667 2282
rect 719 2286 723 2287
rect 719 2281 723 2282
rect 759 2286 763 2287
rect 759 2281 763 2282
rect 847 2286 851 2287
rect 847 2281 851 2282
rect 863 2286 867 2287
rect 863 2281 867 2282
rect 967 2286 971 2287
rect 967 2281 971 2282
rect 975 2286 979 2287
rect 975 2281 979 2282
rect 1079 2286 1083 2287
rect 1079 2281 1083 2282
rect 1103 2286 1107 2287
rect 1103 2281 1107 2282
rect 1191 2286 1195 2287
rect 1191 2281 1195 2282
rect 1239 2286 1243 2287
rect 1239 2281 1243 2282
rect 1303 2286 1307 2287
rect 1303 2281 1307 2282
rect 1375 2286 1379 2287
rect 1375 2281 1379 2282
rect 1415 2286 1419 2287
rect 1415 2281 1419 2282
rect 1511 2286 1515 2287
rect 1511 2281 1515 2282
rect 1767 2286 1771 2287
rect 1808 2283 1810 2303
rect 1888 2283 1890 2304
rect 2016 2283 2018 2304
rect 2152 2283 2154 2304
rect 2304 2283 2306 2304
rect 2464 2283 2466 2304
rect 2648 2283 2650 2304
rect 2840 2283 2842 2304
rect 3048 2283 3050 2304
rect 3256 2283 3258 2304
rect 3462 2303 3468 2304
rect 3464 2283 3466 2303
rect 1767 2281 1771 2282
rect 1807 2282 1811 2283
rect 112 2262 114 2281
rect 576 2265 578 2281
rect 664 2265 666 2281
rect 760 2265 762 2281
rect 864 2265 866 2281
rect 968 2265 970 2281
rect 1080 2265 1082 2281
rect 1192 2265 1194 2281
rect 1304 2265 1306 2281
rect 1416 2265 1418 2281
rect 574 2264 580 2265
rect 110 2261 116 2262
rect 110 2257 111 2261
rect 115 2257 116 2261
rect 574 2260 575 2264
rect 579 2260 580 2264
rect 574 2259 580 2260
rect 662 2264 668 2265
rect 662 2260 663 2264
rect 667 2260 668 2264
rect 662 2259 668 2260
rect 758 2264 764 2265
rect 758 2260 759 2264
rect 763 2260 764 2264
rect 758 2259 764 2260
rect 862 2264 868 2265
rect 862 2260 863 2264
rect 867 2260 868 2264
rect 862 2259 868 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1078 2264 1084 2265
rect 1078 2260 1079 2264
rect 1083 2260 1084 2264
rect 1078 2259 1084 2260
rect 1190 2264 1196 2265
rect 1190 2260 1191 2264
rect 1195 2260 1196 2264
rect 1190 2259 1196 2260
rect 1302 2264 1308 2265
rect 1302 2260 1303 2264
rect 1307 2260 1308 2264
rect 1302 2259 1308 2260
rect 1414 2264 1420 2265
rect 1414 2260 1415 2264
rect 1419 2260 1420 2264
rect 1768 2262 1770 2281
rect 1807 2277 1811 2278
rect 1887 2282 1891 2283
rect 1887 2277 1891 2278
rect 2015 2282 2019 2283
rect 2015 2277 2019 2278
rect 2039 2282 2043 2283
rect 2039 2277 2043 2278
rect 2135 2282 2139 2283
rect 2135 2277 2139 2278
rect 2151 2282 2155 2283
rect 2151 2277 2155 2278
rect 2239 2282 2243 2283
rect 2239 2277 2243 2278
rect 2303 2282 2307 2283
rect 2303 2277 2307 2278
rect 2343 2282 2347 2283
rect 2343 2277 2347 2278
rect 2463 2282 2467 2283
rect 2463 2277 2467 2278
rect 2591 2282 2595 2283
rect 2591 2277 2595 2278
rect 2647 2282 2651 2283
rect 2647 2277 2651 2278
rect 2735 2282 2739 2283
rect 2735 2277 2739 2278
rect 2839 2282 2843 2283
rect 2839 2277 2843 2278
rect 2887 2282 2891 2283
rect 2887 2277 2891 2278
rect 3047 2282 3051 2283
rect 3047 2277 3051 2278
rect 3215 2282 3219 2283
rect 3215 2277 3219 2278
rect 3255 2282 3259 2283
rect 3255 2277 3259 2278
rect 3367 2282 3371 2283
rect 3367 2277 3371 2278
rect 3463 2282 3467 2283
rect 3463 2277 3467 2278
rect 1414 2259 1420 2260
rect 1766 2261 1772 2262
rect 1808 2261 1810 2277
rect 110 2256 116 2257
rect 1766 2257 1767 2261
rect 1771 2257 1772 2261
rect 1766 2256 1772 2257
rect 1806 2260 1812 2261
rect 2040 2260 2042 2277
rect 2136 2260 2138 2277
rect 2240 2260 2242 2277
rect 2344 2260 2346 2277
rect 2464 2260 2466 2277
rect 2592 2260 2594 2277
rect 2736 2260 2738 2277
rect 2888 2260 2890 2277
rect 3048 2260 3050 2277
rect 3216 2260 3218 2277
rect 3368 2260 3370 2277
rect 3464 2261 3466 2277
rect 3462 2260 3468 2261
rect 1806 2256 1807 2260
rect 1811 2256 1812 2260
rect 1806 2255 1812 2256
rect 2038 2259 2044 2260
rect 2038 2255 2039 2259
rect 2043 2255 2044 2259
rect 2038 2254 2044 2255
rect 2134 2259 2140 2260
rect 2134 2255 2135 2259
rect 2139 2255 2140 2259
rect 2134 2254 2140 2255
rect 2238 2259 2244 2260
rect 2238 2255 2239 2259
rect 2243 2255 2244 2259
rect 2238 2254 2244 2255
rect 2342 2259 2348 2260
rect 2342 2255 2343 2259
rect 2347 2255 2348 2259
rect 2342 2254 2348 2255
rect 2462 2259 2468 2260
rect 2462 2255 2463 2259
rect 2467 2255 2468 2259
rect 2462 2254 2468 2255
rect 2590 2259 2596 2260
rect 2590 2255 2591 2259
rect 2595 2255 2596 2259
rect 2590 2254 2596 2255
rect 2734 2259 2740 2260
rect 2734 2255 2735 2259
rect 2739 2255 2740 2259
rect 2734 2254 2740 2255
rect 2886 2259 2892 2260
rect 2886 2255 2887 2259
rect 2891 2255 2892 2259
rect 2886 2254 2892 2255
rect 3046 2259 3052 2260
rect 3046 2255 3047 2259
rect 3051 2255 3052 2259
rect 3046 2254 3052 2255
rect 3214 2259 3220 2260
rect 3214 2255 3215 2259
rect 3219 2255 3220 2259
rect 3214 2254 3220 2255
rect 3366 2259 3372 2260
rect 3366 2255 3367 2259
rect 3371 2255 3372 2259
rect 3462 2256 3463 2260
rect 3467 2256 3468 2260
rect 3462 2255 3468 2256
rect 3366 2254 3372 2255
rect 574 2245 580 2246
rect 110 2244 116 2245
rect 110 2240 111 2244
rect 115 2240 116 2244
rect 574 2241 575 2245
rect 579 2241 580 2245
rect 574 2240 580 2241
rect 662 2245 668 2246
rect 662 2241 663 2245
rect 667 2241 668 2245
rect 662 2240 668 2241
rect 758 2245 764 2246
rect 758 2241 759 2245
rect 763 2241 764 2245
rect 758 2240 764 2241
rect 862 2245 868 2246
rect 862 2241 863 2245
rect 867 2241 868 2245
rect 862 2240 868 2241
rect 966 2245 972 2246
rect 966 2241 967 2245
rect 971 2241 972 2245
rect 966 2240 972 2241
rect 1078 2245 1084 2246
rect 1078 2241 1079 2245
rect 1083 2241 1084 2245
rect 1078 2240 1084 2241
rect 1190 2245 1196 2246
rect 1190 2241 1191 2245
rect 1195 2241 1196 2245
rect 1190 2240 1196 2241
rect 1302 2245 1308 2246
rect 1302 2241 1303 2245
rect 1307 2241 1308 2245
rect 1302 2240 1308 2241
rect 1414 2245 1420 2246
rect 1414 2241 1415 2245
rect 1419 2241 1420 2245
rect 1414 2240 1420 2241
rect 1766 2244 1772 2245
rect 1766 2240 1767 2244
rect 1771 2240 1772 2244
rect 110 2239 116 2240
rect 112 2223 114 2239
rect 576 2223 578 2240
rect 664 2223 666 2240
rect 760 2223 762 2240
rect 864 2223 866 2240
rect 968 2223 970 2240
rect 1080 2223 1082 2240
rect 1192 2223 1194 2240
rect 1304 2223 1306 2240
rect 1416 2223 1418 2240
rect 1766 2239 1772 2240
rect 1806 2243 1812 2244
rect 1806 2239 1807 2243
rect 1811 2239 1812 2243
rect 3462 2243 3468 2244
rect 1768 2223 1770 2239
rect 1806 2238 1812 2239
rect 2038 2240 2044 2241
rect 111 2222 115 2223
rect 111 2217 115 2218
rect 439 2222 443 2223
rect 439 2217 443 2218
rect 527 2222 531 2223
rect 527 2217 531 2218
rect 575 2222 579 2223
rect 575 2217 579 2218
rect 615 2222 619 2223
rect 615 2217 619 2218
rect 663 2222 667 2223
rect 663 2217 667 2218
rect 703 2222 707 2223
rect 703 2217 707 2218
rect 759 2222 763 2223
rect 759 2217 763 2218
rect 791 2222 795 2223
rect 791 2217 795 2218
rect 863 2222 867 2223
rect 863 2217 867 2218
rect 879 2222 883 2223
rect 879 2217 883 2218
rect 967 2222 971 2223
rect 967 2217 971 2218
rect 1055 2222 1059 2223
rect 1055 2217 1059 2218
rect 1079 2222 1083 2223
rect 1079 2217 1083 2218
rect 1143 2222 1147 2223
rect 1143 2217 1147 2218
rect 1191 2222 1195 2223
rect 1191 2217 1195 2218
rect 1231 2222 1235 2223
rect 1231 2217 1235 2218
rect 1303 2222 1307 2223
rect 1303 2217 1307 2218
rect 1319 2222 1323 2223
rect 1319 2217 1323 2218
rect 1415 2222 1419 2223
rect 1415 2217 1419 2218
rect 1767 2222 1771 2223
rect 1767 2217 1771 2218
rect 112 2201 114 2217
rect 110 2200 116 2201
rect 440 2200 442 2217
rect 528 2200 530 2217
rect 616 2200 618 2217
rect 704 2200 706 2217
rect 792 2200 794 2217
rect 880 2200 882 2217
rect 968 2200 970 2217
rect 1056 2200 1058 2217
rect 1144 2200 1146 2217
rect 1232 2200 1234 2217
rect 1320 2200 1322 2217
rect 1768 2201 1770 2217
rect 1808 2207 1810 2238
rect 2038 2236 2039 2240
rect 2043 2236 2044 2240
rect 2038 2235 2044 2236
rect 2134 2240 2140 2241
rect 2134 2236 2135 2240
rect 2139 2236 2140 2240
rect 2134 2235 2140 2236
rect 2238 2240 2244 2241
rect 2238 2236 2239 2240
rect 2243 2236 2244 2240
rect 2238 2235 2244 2236
rect 2342 2240 2348 2241
rect 2342 2236 2343 2240
rect 2347 2236 2348 2240
rect 2342 2235 2348 2236
rect 2462 2240 2468 2241
rect 2462 2236 2463 2240
rect 2467 2236 2468 2240
rect 2462 2235 2468 2236
rect 2590 2240 2596 2241
rect 2590 2236 2591 2240
rect 2595 2236 2596 2240
rect 2590 2235 2596 2236
rect 2734 2240 2740 2241
rect 2734 2236 2735 2240
rect 2739 2236 2740 2240
rect 2734 2235 2740 2236
rect 2886 2240 2892 2241
rect 2886 2236 2887 2240
rect 2891 2236 2892 2240
rect 2886 2235 2892 2236
rect 3046 2240 3052 2241
rect 3046 2236 3047 2240
rect 3051 2236 3052 2240
rect 3046 2235 3052 2236
rect 3214 2240 3220 2241
rect 3214 2236 3215 2240
rect 3219 2236 3220 2240
rect 3214 2235 3220 2236
rect 3366 2240 3372 2241
rect 3366 2236 3367 2240
rect 3371 2236 3372 2240
rect 3462 2239 3463 2243
rect 3467 2239 3468 2243
rect 3462 2238 3468 2239
rect 3366 2235 3372 2236
rect 2040 2207 2042 2235
rect 2136 2207 2138 2235
rect 2240 2207 2242 2235
rect 2344 2207 2346 2235
rect 2464 2207 2466 2235
rect 2592 2207 2594 2235
rect 2736 2207 2738 2235
rect 2888 2207 2890 2235
rect 3048 2207 3050 2235
rect 3216 2207 3218 2235
rect 3368 2207 3370 2235
rect 3464 2207 3466 2238
rect 1807 2206 1811 2207
rect 1807 2201 1811 2202
rect 2039 2206 2043 2207
rect 2039 2201 2043 2202
rect 2135 2206 2139 2207
rect 2135 2201 2139 2202
rect 2183 2206 2187 2207
rect 2183 2201 2187 2202
rect 2239 2206 2243 2207
rect 2239 2201 2243 2202
rect 2279 2206 2283 2207
rect 2279 2201 2283 2202
rect 2343 2206 2347 2207
rect 2343 2201 2347 2202
rect 2383 2206 2387 2207
rect 2383 2201 2387 2202
rect 2463 2206 2467 2207
rect 2463 2201 2467 2202
rect 2495 2206 2499 2207
rect 2495 2201 2499 2202
rect 2591 2206 2595 2207
rect 2591 2201 2595 2202
rect 2607 2206 2611 2207
rect 2607 2201 2611 2202
rect 2719 2206 2723 2207
rect 2719 2201 2723 2202
rect 2735 2206 2739 2207
rect 2735 2201 2739 2202
rect 2839 2206 2843 2207
rect 2839 2201 2843 2202
rect 2887 2206 2891 2207
rect 2887 2201 2891 2202
rect 2967 2206 2971 2207
rect 2967 2201 2971 2202
rect 3047 2206 3051 2207
rect 3047 2201 3051 2202
rect 3103 2206 3107 2207
rect 3103 2201 3107 2202
rect 3215 2206 3219 2207
rect 3215 2201 3219 2202
rect 3247 2206 3251 2207
rect 3247 2201 3251 2202
rect 3367 2206 3371 2207
rect 3367 2201 3371 2202
rect 3463 2206 3467 2207
rect 3463 2201 3467 2202
rect 1766 2200 1772 2201
rect 110 2196 111 2200
rect 115 2196 116 2200
rect 110 2195 116 2196
rect 438 2199 444 2200
rect 438 2195 439 2199
rect 443 2195 444 2199
rect 438 2194 444 2195
rect 526 2199 532 2200
rect 526 2195 527 2199
rect 531 2195 532 2199
rect 526 2194 532 2195
rect 614 2199 620 2200
rect 614 2195 615 2199
rect 619 2195 620 2199
rect 614 2194 620 2195
rect 702 2199 708 2200
rect 702 2195 703 2199
rect 707 2195 708 2199
rect 702 2194 708 2195
rect 790 2199 796 2200
rect 790 2195 791 2199
rect 795 2195 796 2199
rect 790 2194 796 2195
rect 878 2199 884 2200
rect 878 2195 879 2199
rect 883 2195 884 2199
rect 878 2194 884 2195
rect 966 2199 972 2200
rect 966 2195 967 2199
rect 971 2195 972 2199
rect 966 2194 972 2195
rect 1054 2199 1060 2200
rect 1054 2195 1055 2199
rect 1059 2195 1060 2199
rect 1054 2194 1060 2195
rect 1142 2199 1148 2200
rect 1142 2195 1143 2199
rect 1147 2195 1148 2199
rect 1142 2194 1148 2195
rect 1230 2199 1236 2200
rect 1230 2195 1231 2199
rect 1235 2195 1236 2199
rect 1230 2194 1236 2195
rect 1318 2199 1324 2200
rect 1318 2195 1319 2199
rect 1323 2195 1324 2199
rect 1766 2196 1767 2200
rect 1771 2196 1772 2200
rect 1766 2195 1772 2196
rect 1318 2194 1324 2195
rect 110 2183 116 2184
rect 110 2179 111 2183
rect 115 2179 116 2183
rect 1766 2183 1772 2184
rect 110 2178 116 2179
rect 438 2180 444 2181
rect 112 2143 114 2178
rect 438 2176 439 2180
rect 443 2176 444 2180
rect 438 2175 444 2176
rect 526 2180 532 2181
rect 526 2176 527 2180
rect 531 2176 532 2180
rect 526 2175 532 2176
rect 614 2180 620 2181
rect 614 2176 615 2180
rect 619 2176 620 2180
rect 614 2175 620 2176
rect 702 2180 708 2181
rect 702 2176 703 2180
rect 707 2176 708 2180
rect 702 2175 708 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 878 2180 884 2181
rect 878 2176 879 2180
rect 883 2176 884 2180
rect 878 2175 884 2176
rect 966 2180 972 2181
rect 966 2176 967 2180
rect 971 2176 972 2180
rect 966 2175 972 2176
rect 1054 2180 1060 2181
rect 1054 2176 1055 2180
rect 1059 2176 1060 2180
rect 1054 2175 1060 2176
rect 1142 2180 1148 2181
rect 1142 2176 1143 2180
rect 1147 2176 1148 2180
rect 1142 2175 1148 2176
rect 1230 2180 1236 2181
rect 1230 2176 1231 2180
rect 1235 2176 1236 2180
rect 1230 2175 1236 2176
rect 1318 2180 1324 2181
rect 1318 2176 1319 2180
rect 1323 2176 1324 2180
rect 1766 2179 1767 2183
rect 1771 2179 1772 2183
rect 1808 2182 1810 2201
rect 2184 2185 2186 2201
rect 2280 2185 2282 2201
rect 2384 2185 2386 2201
rect 2496 2185 2498 2201
rect 2608 2185 2610 2201
rect 2720 2185 2722 2201
rect 2840 2185 2842 2201
rect 2968 2185 2970 2201
rect 3104 2185 3106 2201
rect 3248 2185 3250 2201
rect 3368 2185 3370 2201
rect 2182 2184 2188 2185
rect 1766 2178 1772 2179
rect 1806 2181 1812 2182
rect 1318 2175 1324 2176
rect 440 2143 442 2175
rect 528 2143 530 2175
rect 616 2143 618 2175
rect 704 2143 706 2175
rect 792 2143 794 2175
rect 880 2143 882 2175
rect 968 2143 970 2175
rect 1056 2143 1058 2175
rect 1144 2143 1146 2175
rect 1232 2143 1234 2175
rect 1320 2143 1322 2175
rect 1768 2143 1770 2178
rect 1806 2177 1807 2181
rect 1811 2177 1812 2181
rect 2182 2180 2183 2184
rect 2187 2180 2188 2184
rect 2182 2179 2188 2180
rect 2278 2184 2284 2185
rect 2278 2180 2279 2184
rect 2283 2180 2284 2184
rect 2278 2179 2284 2180
rect 2382 2184 2388 2185
rect 2382 2180 2383 2184
rect 2387 2180 2388 2184
rect 2382 2179 2388 2180
rect 2494 2184 2500 2185
rect 2494 2180 2495 2184
rect 2499 2180 2500 2184
rect 2494 2179 2500 2180
rect 2606 2184 2612 2185
rect 2606 2180 2607 2184
rect 2611 2180 2612 2184
rect 2606 2179 2612 2180
rect 2718 2184 2724 2185
rect 2718 2180 2719 2184
rect 2723 2180 2724 2184
rect 2718 2179 2724 2180
rect 2838 2184 2844 2185
rect 2838 2180 2839 2184
rect 2843 2180 2844 2184
rect 2838 2179 2844 2180
rect 2966 2184 2972 2185
rect 2966 2180 2967 2184
rect 2971 2180 2972 2184
rect 2966 2179 2972 2180
rect 3102 2184 3108 2185
rect 3102 2180 3103 2184
rect 3107 2180 3108 2184
rect 3102 2179 3108 2180
rect 3246 2184 3252 2185
rect 3246 2180 3247 2184
rect 3251 2180 3252 2184
rect 3246 2179 3252 2180
rect 3366 2184 3372 2185
rect 3366 2180 3367 2184
rect 3371 2180 3372 2184
rect 3464 2182 3466 2201
rect 3366 2179 3372 2180
rect 3462 2181 3468 2182
rect 1806 2176 1812 2177
rect 3462 2177 3463 2181
rect 3467 2177 3468 2181
rect 3462 2176 3468 2177
rect 2182 2165 2188 2166
rect 1806 2164 1812 2165
rect 1806 2160 1807 2164
rect 1811 2160 1812 2164
rect 2182 2161 2183 2165
rect 2187 2161 2188 2165
rect 2182 2160 2188 2161
rect 2278 2165 2284 2166
rect 2278 2161 2279 2165
rect 2283 2161 2284 2165
rect 2278 2160 2284 2161
rect 2382 2165 2388 2166
rect 2382 2161 2383 2165
rect 2387 2161 2388 2165
rect 2382 2160 2388 2161
rect 2494 2165 2500 2166
rect 2494 2161 2495 2165
rect 2499 2161 2500 2165
rect 2494 2160 2500 2161
rect 2606 2165 2612 2166
rect 2606 2161 2607 2165
rect 2611 2161 2612 2165
rect 2606 2160 2612 2161
rect 2718 2165 2724 2166
rect 2718 2161 2719 2165
rect 2723 2161 2724 2165
rect 2718 2160 2724 2161
rect 2838 2165 2844 2166
rect 2838 2161 2839 2165
rect 2843 2161 2844 2165
rect 2838 2160 2844 2161
rect 2966 2165 2972 2166
rect 2966 2161 2967 2165
rect 2971 2161 2972 2165
rect 2966 2160 2972 2161
rect 3102 2165 3108 2166
rect 3102 2161 3103 2165
rect 3107 2161 3108 2165
rect 3102 2160 3108 2161
rect 3246 2165 3252 2166
rect 3246 2161 3247 2165
rect 3251 2161 3252 2165
rect 3246 2160 3252 2161
rect 3366 2165 3372 2166
rect 3366 2161 3367 2165
rect 3371 2161 3372 2165
rect 3366 2160 3372 2161
rect 3462 2164 3468 2165
rect 3462 2160 3463 2164
rect 3467 2160 3468 2164
rect 1806 2159 1812 2160
rect 111 2142 115 2143
rect 111 2137 115 2138
rect 303 2142 307 2143
rect 303 2137 307 2138
rect 407 2142 411 2143
rect 407 2137 411 2138
rect 439 2142 443 2143
rect 439 2137 443 2138
rect 519 2142 523 2143
rect 519 2137 523 2138
rect 527 2142 531 2143
rect 527 2137 531 2138
rect 615 2142 619 2143
rect 615 2137 619 2138
rect 631 2142 635 2143
rect 631 2137 635 2138
rect 703 2142 707 2143
rect 703 2137 707 2138
rect 743 2142 747 2143
rect 743 2137 747 2138
rect 791 2142 795 2143
rect 791 2137 795 2138
rect 863 2142 867 2143
rect 863 2137 867 2138
rect 879 2142 883 2143
rect 879 2137 883 2138
rect 967 2142 971 2143
rect 967 2137 971 2138
rect 983 2142 987 2143
rect 983 2137 987 2138
rect 1055 2142 1059 2143
rect 1055 2137 1059 2138
rect 1143 2142 1147 2143
rect 1143 2137 1147 2138
rect 1231 2142 1235 2143
rect 1231 2137 1235 2138
rect 1319 2142 1323 2143
rect 1319 2137 1323 2138
rect 1767 2142 1771 2143
rect 1767 2137 1771 2138
rect 112 2118 114 2137
rect 304 2121 306 2137
rect 408 2121 410 2137
rect 520 2121 522 2137
rect 632 2121 634 2137
rect 744 2121 746 2137
rect 864 2121 866 2137
rect 984 2121 986 2137
rect 302 2120 308 2121
rect 110 2117 116 2118
rect 110 2113 111 2117
rect 115 2113 116 2117
rect 302 2116 303 2120
rect 307 2116 308 2120
rect 302 2115 308 2116
rect 406 2120 412 2121
rect 406 2116 407 2120
rect 411 2116 412 2120
rect 406 2115 412 2116
rect 518 2120 524 2121
rect 518 2116 519 2120
rect 523 2116 524 2120
rect 518 2115 524 2116
rect 630 2120 636 2121
rect 630 2116 631 2120
rect 635 2116 636 2120
rect 630 2115 636 2116
rect 742 2120 748 2121
rect 742 2116 743 2120
rect 747 2116 748 2120
rect 742 2115 748 2116
rect 862 2120 868 2121
rect 862 2116 863 2120
rect 867 2116 868 2120
rect 862 2115 868 2116
rect 982 2120 988 2121
rect 982 2116 983 2120
rect 987 2116 988 2120
rect 1768 2118 1770 2137
rect 1808 2135 1810 2159
rect 2184 2135 2186 2160
rect 2280 2135 2282 2160
rect 2384 2135 2386 2160
rect 2496 2135 2498 2160
rect 2608 2135 2610 2160
rect 2720 2135 2722 2160
rect 2840 2135 2842 2160
rect 2968 2135 2970 2160
rect 3104 2135 3106 2160
rect 3248 2135 3250 2160
rect 3368 2135 3370 2160
rect 3462 2159 3468 2160
rect 3464 2135 3466 2159
rect 1807 2134 1811 2135
rect 1807 2129 1811 2130
rect 2135 2134 2139 2135
rect 2135 2129 2139 2130
rect 2183 2134 2187 2135
rect 2183 2129 2187 2130
rect 2255 2134 2259 2135
rect 2255 2129 2259 2130
rect 2279 2134 2283 2135
rect 2279 2129 2283 2130
rect 2383 2134 2387 2135
rect 2383 2129 2387 2130
rect 2495 2134 2499 2135
rect 2495 2129 2499 2130
rect 2519 2134 2523 2135
rect 2519 2129 2523 2130
rect 2607 2134 2611 2135
rect 2607 2129 2611 2130
rect 2655 2134 2659 2135
rect 2655 2129 2659 2130
rect 2719 2134 2723 2135
rect 2719 2129 2723 2130
rect 2783 2134 2787 2135
rect 2783 2129 2787 2130
rect 2839 2134 2843 2135
rect 2839 2129 2843 2130
rect 2911 2134 2915 2135
rect 2911 2129 2915 2130
rect 2967 2134 2971 2135
rect 2967 2129 2971 2130
rect 3031 2134 3035 2135
rect 3031 2129 3035 2130
rect 3103 2134 3107 2135
rect 3103 2129 3107 2130
rect 3151 2134 3155 2135
rect 3151 2129 3155 2130
rect 3247 2134 3251 2135
rect 3247 2129 3251 2130
rect 3271 2134 3275 2135
rect 3271 2129 3275 2130
rect 3367 2134 3371 2135
rect 3367 2129 3371 2130
rect 3463 2134 3467 2135
rect 3463 2129 3467 2130
rect 982 2115 988 2116
rect 1766 2117 1772 2118
rect 110 2112 116 2113
rect 1766 2113 1767 2117
rect 1771 2113 1772 2117
rect 1808 2113 1810 2129
rect 1766 2112 1772 2113
rect 1806 2112 1812 2113
rect 2136 2112 2138 2129
rect 2256 2112 2258 2129
rect 2384 2112 2386 2129
rect 2520 2112 2522 2129
rect 2656 2112 2658 2129
rect 2784 2112 2786 2129
rect 2912 2112 2914 2129
rect 3032 2112 3034 2129
rect 3152 2112 3154 2129
rect 3272 2112 3274 2129
rect 3368 2112 3370 2129
rect 3464 2113 3466 2129
rect 3462 2112 3468 2113
rect 1806 2108 1807 2112
rect 1811 2108 1812 2112
rect 1806 2107 1812 2108
rect 2134 2111 2140 2112
rect 2134 2107 2135 2111
rect 2139 2107 2140 2111
rect 2134 2106 2140 2107
rect 2254 2111 2260 2112
rect 2254 2107 2255 2111
rect 2259 2107 2260 2111
rect 2254 2106 2260 2107
rect 2382 2111 2388 2112
rect 2382 2107 2383 2111
rect 2387 2107 2388 2111
rect 2382 2106 2388 2107
rect 2518 2111 2524 2112
rect 2518 2107 2519 2111
rect 2523 2107 2524 2111
rect 2518 2106 2524 2107
rect 2654 2111 2660 2112
rect 2654 2107 2655 2111
rect 2659 2107 2660 2111
rect 2654 2106 2660 2107
rect 2782 2111 2788 2112
rect 2782 2107 2783 2111
rect 2787 2107 2788 2111
rect 2782 2106 2788 2107
rect 2910 2111 2916 2112
rect 2910 2107 2911 2111
rect 2915 2107 2916 2111
rect 2910 2106 2916 2107
rect 3030 2111 3036 2112
rect 3030 2107 3031 2111
rect 3035 2107 3036 2111
rect 3030 2106 3036 2107
rect 3150 2111 3156 2112
rect 3150 2107 3151 2111
rect 3155 2107 3156 2111
rect 3150 2106 3156 2107
rect 3270 2111 3276 2112
rect 3270 2107 3271 2111
rect 3275 2107 3276 2111
rect 3270 2106 3276 2107
rect 3366 2111 3372 2112
rect 3366 2107 3367 2111
rect 3371 2107 3372 2111
rect 3462 2108 3463 2112
rect 3467 2108 3468 2112
rect 3462 2107 3468 2108
rect 3366 2106 3372 2107
rect 302 2101 308 2102
rect 110 2100 116 2101
rect 110 2096 111 2100
rect 115 2096 116 2100
rect 302 2097 303 2101
rect 307 2097 308 2101
rect 302 2096 308 2097
rect 406 2101 412 2102
rect 406 2097 407 2101
rect 411 2097 412 2101
rect 406 2096 412 2097
rect 518 2101 524 2102
rect 518 2097 519 2101
rect 523 2097 524 2101
rect 518 2096 524 2097
rect 630 2101 636 2102
rect 630 2097 631 2101
rect 635 2097 636 2101
rect 630 2096 636 2097
rect 742 2101 748 2102
rect 742 2097 743 2101
rect 747 2097 748 2101
rect 742 2096 748 2097
rect 862 2101 868 2102
rect 862 2097 863 2101
rect 867 2097 868 2101
rect 862 2096 868 2097
rect 982 2101 988 2102
rect 982 2097 983 2101
rect 987 2097 988 2101
rect 982 2096 988 2097
rect 1766 2100 1772 2101
rect 1766 2096 1767 2100
rect 1771 2096 1772 2100
rect 110 2095 116 2096
rect 112 2079 114 2095
rect 304 2079 306 2096
rect 408 2079 410 2096
rect 520 2079 522 2096
rect 632 2079 634 2096
rect 744 2079 746 2096
rect 864 2079 866 2096
rect 984 2079 986 2096
rect 1766 2095 1772 2096
rect 1806 2095 1812 2096
rect 1768 2079 1770 2095
rect 1806 2091 1807 2095
rect 1811 2091 1812 2095
rect 3462 2095 3468 2096
rect 1806 2090 1812 2091
rect 2134 2092 2140 2093
rect 111 2078 115 2079
rect 111 2073 115 2074
rect 255 2078 259 2079
rect 255 2073 259 2074
rect 303 2078 307 2079
rect 303 2073 307 2074
rect 375 2078 379 2079
rect 375 2073 379 2074
rect 407 2078 411 2079
rect 407 2073 411 2074
rect 495 2078 499 2079
rect 495 2073 499 2074
rect 519 2078 523 2079
rect 519 2073 523 2074
rect 615 2078 619 2079
rect 615 2073 619 2074
rect 631 2078 635 2079
rect 631 2073 635 2074
rect 727 2078 731 2079
rect 727 2073 731 2074
rect 743 2078 747 2079
rect 743 2073 747 2074
rect 831 2078 835 2079
rect 831 2073 835 2074
rect 863 2078 867 2079
rect 863 2073 867 2074
rect 935 2078 939 2079
rect 935 2073 939 2074
rect 983 2078 987 2079
rect 983 2073 987 2074
rect 1039 2078 1043 2079
rect 1039 2073 1043 2074
rect 1143 2078 1147 2079
rect 1143 2073 1147 2074
rect 1255 2078 1259 2079
rect 1255 2073 1259 2074
rect 1767 2078 1771 2079
rect 1767 2073 1771 2074
rect 112 2057 114 2073
rect 110 2056 116 2057
rect 256 2056 258 2073
rect 376 2056 378 2073
rect 496 2056 498 2073
rect 616 2056 618 2073
rect 728 2056 730 2073
rect 832 2056 834 2073
rect 936 2056 938 2073
rect 1040 2056 1042 2073
rect 1144 2056 1146 2073
rect 1256 2056 1258 2073
rect 1768 2057 1770 2073
rect 1808 2063 1810 2090
rect 2134 2088 2135 2092
rect 2139 2088 2140 2092
rect 2134 2087 2140 2088
rect 2254 2092 2260 2093
rect 2254 2088 2255 2092
rect 2259 2088 2260 2092
rect 2254 2087 2260 2088
rect 2382 2092 2388 2093
rect 2382 2088 2383 2092
rect 2387 2088 2388 2092
rect 2382 2087 2388 2088
rect 2518 2092 2524 2093
rect 2518 2088 2519 2092
rect 2523 2088 2524 2092
rect 2518 2087 2524 2088
rect 2654 2092 2660 2093
rect 2654 2088 2655 2092
rect 2659 2088 2660 2092
rect 2654 2087 2660 2088
rect 2782 2092 2788 2093
rect 2782 2088 2783 2092
rect 2787 2088 2788 2092
rect 2782 2087 2788 2088
rect 2910 2092 2916 2093
rect 2910 2088 2911 2092
rect 2915 2088 2916 2092
rect 2910 2087 2916 2088
rect 3030 2092 3036 2093
rect 3030 2088 3031 2092
rect 3035 2088 3036 2092
rect 3030 2087 3036 2088
rect 3150 2092 3156 2093
rect 3150 2088 3151 2092
rect 3155 2088 3156 2092
rect 3150 2087 3156 2088
rect 3270 2092 3276 2093
rect 3270 2088 3271 2092
rect 3275 2088 3276 2092
rect 3270 2087 3276 2088
rect 3366 2092 3372 2093
rect 3366 2088 3367 2092
rect 3371 2088 3372 2092
rect 3462 2091 3463 2095
rect 3467 2091 3468 2095
rect 3462 2090 3468 2091
rect 3366 2087 3372 2088
rect 2136 2063 2138 2087
rect 2256 2063 2258 2087
rect 2384 2063 2386 2087
rect 2520 2063 2522 2087
rect 2656 2063 2658 2087
rect 2784 2063 2786 2087
rect 2912 2063 2914 2087
rect 3032 2063 3034 2087
rect 3152 2063 3154 2087
rect 3272 2063 3274 2087
rect 3368 2063 3370 2087
rect 3464 2063 3466 2090
rect 1807 2062 1811 2063
rect 1807 2057 1811 2058
rect 2135 2062 2139 2063
rect 2135 2057 2139 2058
rect 2247 2062 2251 2063
rect 2247 2057 2251 2058
rect 2255 2062 2259 2063
rect 2255 2057 2259 2058
rect 2383 2062 2387 2063
rect 2383 2057 2387 2058
rect 2415 2062 2419 2063
rect 2415 2057 2419 2058
rect 2519 2062 2523 2063
rect 2519 2057 2523 2058
rect 2575 2062 2579 2063
rect 2575 2057 2579 2058
rect 2655 2062 2659 2063
rect 2655 2057 2659 2058
rect 2727 2062 2731 2063
rect 2727 2057 2731 2058
rect 2783 2062 2787 2063
rect 2783 2057 2787 2058
rect 2871 2062 2875 2063
rect 2871 2057 2875 2058
rect 2911 2062 2915 2063
rect 2911 2057 2915 2058
rect 3007 2062 3011 2063
rect 3007 2057 3011 2058
rect 3031 2062 3035 2063
rect 3031 2057 3035 2058
rect 3135 2062 3139 2063
rect 3135 2057 3139 2058
rect 3151 2062 3155 2063
rect 3151 2057 3155 2058
rect 3263 2062 3267 2063
rect 3263 2057 3267 2058
rect 3271 2062 3275 2063
rect 3271 2057 3275 2058
rect 3367 2062 3371 2063
rect 3367 2057 3371 2058
rect 3463 2062 3467 2063
rect 3463 2057 3467 2058
rect 1766 2056 1772 2057
rect 110 2052 111 2056
rect 115 2052 116 2056
rect 110 2051 116 2052
rect 254 2055 260 2056
rect 254 2051 255 2055
rect 259 2051 260 2055
rect 254 2050 260 2051
rect 374 2055 380 2056
rect 374 2051 375 2055
rect 379 2051 380 2055
rect 374 2050 380 2051
rect 494 2055 500 2056
rect 494 2051 495 2055
rect 499 2051 500 2055
rect 494 2050 500 2051
rect 614 2055 620 2056
rect 614 2051 615 2055
rect 619 2051 620 2055
rect 614 2050 620 2051
rect 726 2055 732 2056
rect 726 2051 727 2055
rect 731 2051 732 2055
rect 726 2050 732 2051
rect 830 2055 836 2056
rect 830 2051 831 2055
rect 835 2051 836 2055
rect 830 2050 836 2051
rect 934 2055 940 2056
rect 934 2051 935 2055
rect 939 2051 940 2055
rect 934 2050 940 2051
rect 1038 2055 1044 2056
rect 1038 2051 1039 2055
rect 1043 2051 1044 2055
rect 1038 2050 1044 2051
rect 1142 2055 1148 2056
rect 1142 2051 1143 2055
rect 1147 2051 1148 2055
rect 1142 2050 1148 2051
rect 1254 2055 1260 2056
rect 1254 2051 1255 2055
rect 1259 2051 1260 2055
rect 1766 2052 1767 2056
rect 1771 2052 1772 2056
rect 1766 2051 1772 2052
rect 1254 2050 1260 2051
rect 110 2039 116 2040
rect 110 2035 111 2039
rect 115 2035 116 2039
rect 1766 2039 1772 2040
rect 110 2034 116 2035
rect 254 2036 260 2037
rect 112 2015 114 2034
rect 254 2032 255 2036
rect 259 2032 260 2036
rect 254 2031 260 2032
rect 374 2036 380 2037
rect 374 2032 375 2036
rect 379 2032 380 2036
rect 374 2031 380 2032
rect 494 2036 500 2037
rect 494 2032 495 2036
rect 499 2032 500 2036
rect 494 2031 500 2032
rect 614 2036 620 2037
rect 614 2032 615 2036
rect 619 2032 620 2036
rect 614 2031 620 2032
rect 726 2036 732 2037
rect 726 2032 727 2036
rect 731 2032 732 2036
rect 726 2031 732 2032
rect 830 2036 836 2037
rect 830 2032 831 2036
rect 835 2032 836 2036
rect 830 2031 836 2032
rect 934 2036 940 2037
rect 934 2032 935 2036
rect 939 2032 940 2036
rect 934 2031 940 2032
rect 1038 2036 1044 2037
rect 1038 2032 1039 2036
rect 1043 2032 1044 2036
rect 1038 2031 1044 2032
rect 1142 2036 1148 2037
rect 1142 2032 1143 2036
rect 1147 2032 1148 2036
rect 1142 2031 1148 2032
rect 1254 2036 1260 2037
rect 1254 2032 1255 2036
rect 1259 2032 1260 2036
rect 1766 2035 1767 2039
rect 1771 2035 1772 2039
rect 1808 2038 1810 2057
rect 2248 2041 2250 2057
rect 2416 2041 2418 2057
rect 2576 2041 2578 2057
rect 2728 2041 2730 2057
rect 2872 2041 2874 2057
rect 3008 2041 3010 2057
rect 3136 2041 3138 2057
rect 3264 2041 3266 2057
rect 3368 2041 3370 2057
rect 2246 2040 2252 2041
rect 1766 2034 1772 2035
rect 1806 2037 1812 2038
rect 1254 2031 1260 2032
rect 256 2015 258 2031
rect 376 2015 378 2031
rect 496 2015 498 2031
rect 616 2015 618 2031
rect 728 2015 730 2031
rect 832 2015 834 2031
rect 936 2015 938 2031
rect 1040 2015 1042 2031
rect 1144 2015 1146 2031
rect 1256 2015 1258 2031
rect 1768 2015 1770 2034
rect 1806 2033 1807 2037
rect 1811 2033 1812 2037
rect 2246 2036 2247 2040
rect 2251 2036 2252 2040
rect 2246 2035 2252 2036
rect 2414 2040 2420 2041
rect 2414 2036 2415 2040
rect 2419 2036 2420 2040
rect 2414 2035 2420 2036
rect 2574 2040 2580 2041
rect 2574 2036 2575 2040
rect 2579 2036 2580 2040
rect 2574 2035 2580 2036
rect 2726 2040 2732 2041
rect 2726 2036 2727 2040
rect 2731 2036 2732 2040
rect 2726 2035 2732 2036
rect 2870 2040 2876 2041
rect 2870 2036 2871 2040
rect 2875 2036 2876 2040
rect 2870 2035 2876 2036
rect 3006 2040 3012 2041
rect 3006 2036 3007 2040
rect 3011 2036 3012 2040
rect 3006 2035 3012 2036
rect 3134 2040 3140 2041
rect 3134 2036 3135 2040
rect 3139 2036 3140 2040
rect 3134 2035 3140 2036
rect 3262 2040 3268 2041
rect 3262 2036 3263 2040
rect 3267 2036 3268 2040
rect 3262 2035 3268 2036
rect 3366 2040 3372 2041
rect 3366 2036 3367 2040
rect 3371 2036 3372 2040
rect 3464 2038 3466 2057
rect 3366 2035 3372 2036
rect 3462 2037 3468 2038
rect 1806 2032 1812 2033
rect 3462 2033 3463 2037
rect 3467 2033 3468 2037
rect 3462 2032 3468 2033
rect 2246 2021 2252 2022
rect 1806 2020 1812 2021
rect 1806 2016 1807 2020
rect 1811 2016 1812 2020
rect 2246 2017 2247 2021
rect 2251 2017 2252 2021
rect 2246 2016 2252 2017
rect 2414 2021 2420 2022
rect 2414 2017 2415 2021
rect 2419 2017 2420 2021
rect 2414 2016 2420 2017
rect 2574 2021 2580 2022
rect 2574 2017 2575 2021
rect 2579 2017 2580 2021
rect 2574 2016 2580 2017
rect 2726 2021 2732 2022
rect 2726 2017 2727 2021
rect 2731 2017 2732 2021
rect 2726 2016 2732 2017
rect 2870 2021 2876 2022
rect 2870 2017 2871 2021
rect 2875 2017 2876 2021
rect 2870 2016 2876 2017
rect 3006 2021 3012 2022
rect 3006 2017 3007 2021
rect 3011 2017 3012 2021
rect 3006 2016 3012 2017
rect 3134 2021 3140 2022
rect 3134 2017 3135 2021
rect 3139 2017 3140 2021
rect 3134 2016 3140 2017
rect 3262 2021 3268 2022
rect 3262 2017 3263 2021
rect 3267 2017 3268 2021
rect 3262 2016 3268 2017
rect 3366 2021 3372 2022
rect 3366 2017 3367 2021
rect 3371 2017 3372 2021
rect 3366 2016 3372 2017
rect 3462 2020 3468 2021
rect 3462 2016 3463 2020
rect 3467 2016 3468 2020
rect 1806 2015 1812 2016
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 255 2014 259 2015
rect 255 2009 259 2010
rect 359 2014 363 2015
rect 359 2009 363 2010
rect 375 2014 379 2015
rect 375 2009 379 2010
rect 487 2014 491 2015
rect 487 2009 491 2010
rect 495 2014 499 2015
rect 495 2009 499 2010
rect 615 2014 619 2015
rect 615 2009 619 2010
rect 623 2014 627 2015
rect 623 2009 627 2010
rect 727 2014 731 2015
rect 727 2009 731 2010
rect 759 2014 763 2015
rect 759 2009 763 2010
rect 831 2014 835 2015
rect 831 2009 835 2010
rect 895 2014 899 2015
rect 895 2009 899 2010
rect 935 2014 939 2015
rect 935 2009 939 2010
rect 1023 2014 1027 2015
rect 1023 2009 1027 2010
rect 1039 2014 1043 2015
rect 1039 2009 1043 2010
rect 1143 2014 1147 2015
rect 1143 2009 1147 2010
rect 1151 2014 1155 2015
rect 1151 2009 1155 2010
rect 1255 2014 1259 2015
rect 1255 2009 1259 2010
rect 1271 2014 1275 2015
rect 1271 2009 1275 2010
rect 1399 2014 1403 2015
rect 1399 2009 1403 2010
rect 1527 2014 1531 2015
rect 1527 2009 1531 2010
rect 1767 2014 1771 2015
rect 1767 2009 1771 2010
rect 112 1990 114 2009
rect 360 1993 362 2009
rect 488 1993 490 2009
rect 624 1993 626 2009
rect 760 1993 762 2009
rect 896 1993 898 2009
rect 1024 1993 1026 2009
rect 1152 1993 1154 2009
rect 1272 1993 1274 2009
rect 1400 1993 1402 2009
rect 1528 1993 1530 2009
rect 358 1992 364 1993
rect 110 1989 116 1990
rect 110 1985 111 1989
rect 115 1985 116 1989
rect 358 1988 359 1992
rect 363 1988 364 1992
rect 358 1987 364 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 622 1992 628 1993
rect 622 1988 623 1992
rect 627 1988 628 1992
rect 622 1987 628 1988
rect 758 1992 764 1993
rect 758 1988 759 1992
rect 763 1988 764 1992
rect 758 1987 764 1988
rect 894 1992 900 1993
rect 894 1988 895 1992
rect 899 1988 900 1992
rect 894 1987 900 1988
rect 1022 1992 1028 1993
rect 1022 1988 1023 1992
rect 1027 1988 1028 1992
rect 1022 1987 1028 1988
rect 1150 1992 1156 1993
rect 1150 1988 1151 1992
rect 1155 1988 1156 1992
rect 1150 1987 1156 1988
rect 1270 1992 1276 1993
rect 1270 1988 1271 1992
rect 1275 1988 1276 1992
rect 1270 1987 1276 1988
rect 1398 1992 1404 1993
rect 1398 1988 1399 1992
rect 1403 1988 1404 1992
rect 1398 1987 1404 1988
rect 1526 1992 1532 1993
rect 1526 1988 1527 1992
rect 1531 1988 1532 1992
rect 1768 1990 1770 2009
rect 1526 1987 1532 1988
rect 1766 1989 1772 1990
rect 110 1984 116 1985
rect 1766 1985 1767 1989
rect 1771 1985 1772 1989
rect 1766 1984 1772 1985
rect 1808 1983 1810 2015
rect 2248 1983 2250 2016
rect 2416 1983 2418 2016
rect 2576 1983 2578 2016
rect 2728 1983 2730 2016
rect 2872 1983 2874 2016
rect 3008 1983 3010 2016
rect 3136 1983 3138 2016
rect 3264 1983 3266 2016
rect 3368 1983 3370 2016
rect 3462 2015 3468 2016
rect 3464 1983 3466 2015
rect 1807 1982 1811 1983
rect 1807 1977 1811 1978
rect 1831 1982 1835 1983
rect 1831 1977 1835 1978
rect 1919 1982 1923 1983
rect 1919 1977 1923 1978
rect 2047 1982 2051 1983
rect 2047 1977 2051 1978
rect 2183 1982 2187 1983
rect 2183 1977 2187 1978
rect 2247 1982 2251 1983
rect 2247 1977 2251 1978
rect 2327 1982 2331 1983
rect 2327 1977 2331 1978
rect 2415 1982 2419 1983
rect 2415 1977 2419 1978
rect 2471 1982 2475 1983
rect 2471 1977 2475 1978
rect 2575 1982 2579 1983
rect 2575 1977 2579 1978
rect 2615 1982 2619 1983
rect 2615 1977 2619 1978
rect 2727 1982 2731 1983
rect 2727 1977 2731 1978
rect 2751 1982 2755 1983
rect 2751 1977 2755 1978
rect 2871 1982 2875 1983
rect 2871 1977 2875 1978
rect 2887 1982 2891 1983
rect 2887 1977 2891 1978
rect 3007 1982 3011 1983
rect 3007 1977 3011 1978
rect 3031 1982 3035 1983
rect 3031 1977 3035 1978
rect 3135 1982 3139 1983
rect 3135 1977 3139 1978
rect 3175 1982 3179 1983
rect 3175 1977 3179 1978
rect 3263 1982 3267 1983
rect 3263 1977 3267 1978
rect 3319 1982 3323 1983
rect 3319 1977 3323 1978
rect 3367 1982 3371 1983
rect 3367 1977 3371 1978
rect 3463 1982 3467 1983
rect 3463 1977 3467 1978
rect 358 1973 364 1974
rect 110 1972 116 1973
rect 110 1968 111 1972
rect 115 1968 116 1972
rect 358 1969 359 1973
rect 363 1969 364 1973
rect 358 1968 364 1969
rect 486 1973 492 1974
rect 486 1969 487 1973
rect 491 1969 492 1973
rect 486 1968 492 1969
rect 622 1973 628 1974
rect 622 1969 623 1973
rect 627 1969 628 1973
rect 622 1968 628 1969
rect 758 1973 764 1974
rect 758 1969 759 1973
rect 763 1969 764 1973
rect 758 1968 764 1969
rect 894 1973 900 1974
rect 894 1969 895 1973
rect 899 1969 900 1973
rect 894 1968 900 1969
rect 1022 1973 1028 1974
rect 1022 1969 1023 1973
rect 1027 1969 1028 1973
rect 1022 1968 1028 1969
rect 1150 1973 1156 1974
rect 1150 1969 1151 1973
rect 1155 1969 1156 1973
rect 1150 1968 1156 1969
rect 1270 1973 1276 1974
rect 1270 1969 1271 1973
rect 1275 1969 1276 1973
rect 1270 1968 1276 1969
rect 1398 1973 1404 1974
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1398 1968 1404 1969
rect 1526 1973 1532 1974
rect 1526 1969 1527 1973
rect 1531 1969 1532 1973
rect 1526 1968 1532 1969
rect 1766 1972 1772 1973
rect 1766 1968 1767 1972
rect 1771 1968 1772 1972
rect 110 1967 116 1968
rect 112 1951 114 1967
rect 360 1951 362 1968
rect 488 1951 490 1968
rect 624 1951 626 1968
rect 760 1951 762 1968
rect 896 1951 898 1968
rect 1024 1951 1026 1968
rect 1152 1951 1154 1968
rect 1272 1951 1274 1968
rect 1400 1951 1402 1968
rect 1528 1951 1530 1968
rect 1766 1967 1772 1968
rect 1768 1951 1770 1967
rect 1808 1961 1810 1977
rect 1806 1960 1812 1961
rect 1832 1960 1834 1977
rect 1920 1960 1922 1977
rect 2048 1960 2050 1977
rect 2184 1960 2186 1977
rect 2328 1960 2330 1977
rect 2472 1960 2474 1977
rect 2616 1960 2618 1977
rect 2752 1960 2754 1977
rect 2888 1960 2890 1977
rect 3032 1960 3034 1977
rect 3176 1960 3178 1977
rect 3320 1960 3322 1977
rect 3464 1961 3466 1977
rect 3462 1960 3468 1961
rect 1806 1956 1807 1960
rect 1811 1956 1812 1960
rect 1806 1955 1812 1956
rect 1830 1959 1836 1960
rect 1830 1955 1831 1959
rect 1835 1955 1836 1959
rect 1830 1954 1836 1955
rect 1918 1959 1924 1960
rect 1918 1955 1919 1959
rect 1923 1955 1924 1959
rect 1918 1954 1924 1955
rect 2046 1959 2052 1960
rect 2046 1955 2047 1959
rect 2051 1955 2052 1959
rect 2046 1954 2052 1955
rect 2182 1959 2188 1960
rect 2182 1955 2183 1959
rect 2187 1955 2188 1959
rect 2182 1954 2188 1955
rect 2326 1959 2332 1960
rect 2326 1955 2327 1959
rect 2331 1955 2332 1959
rect 2326 1954 2332 1955
rect 2470 1959 2476 1960
rect 2470 1955 2471 1959
rect 2475 1955 2476 1959
rect 2470 1954 2476 1955
rect 2614 1959 2620 1960
rect 2614 1955 2615 1959
rect 2619 1955 2620 1959
rect 2614 1954 2620 1955
rect 2750 1959 2756 1960
rect 2750 1955 2751 1959
rect 2755 1955 2756 1959
rect 2750 1954 2756 1955
rect 2886 1959 2892 1960
rect 2886 1955 2887 1959
rect 2891 1955 2892 1959
rect 2886 1954 2892 1955
rect 3030 1959 3036 1960
rect 3030 1955 3031 1959
rect 3035 1955 3036 1959
rect 3030 1954 3036 1955
rect 3174 1959 3180 1960
rect 3174 1955 3175 1959
rect 3179 1955 3180 1959
rect 3174 1954 3180 1955
rect 3318 1959 3324 1960
rect 3318 1955 3319 1959
rect 3323 1955 3324 1959
rect 3462 1956 3463 1960
rect 3467 1956 3468 1960
rect 3462 1955 3468 1956
rect 3318 1954 3324 1955
rect 111 1950 115 1951
rect 111 1945 115 1946
rect 359 1950 363 1951
rect 359 1945 363 1946
rect 447 1950 451 1951
rect 447 1945 451 1946
rect 487 1950 491 1951
rect 487 1945 491 1946
rect 575 1950 579 1951
rect 575 1945 579 1946
rect 623 1950 627 1951
rect 623 1945 627 1946
rect 711 1950 715 1951
rect 711 1945 715 1946
rect 759 1950 763 1951
rect 759 1945 763 1946
rect 847 1950 851 1951
rect 847 1945 851 1946
rect 895 1950 899 1951
rect 895 1945 899 1946
rect 983 1950 987 1951
rect 983 1945 987 1946
rect 1023 1950 1027 1951
rect 1023 1945 1027 1946
rect 1119 1950 1123 1951
rect 1119 1945 1123 1946
rect 1151 1950 1155 1951
rect 1151 1945 1155 1946
rect 1255 1950 1259 1951
rect 1255 1945 1259 1946
rect 1271 1950 1275 1951
rect 1271 1945 1275 1946
rect 1383 1950 1387 1951
rect 1383 1945 1387 1946
rect 1399 1950 1403 1951
rect 1399 1945 1403 1946
rect 1519 1950 1523 1951
rect 1519 1945 1523 1946
rect 1527 1950 1531 1951
rect 1527 1945 1531 1946
rect 1655 1950 1659 1951
rect 1655 1945 1659 1946
rect 1767 1950 1771 1951
rect 1767 1945 1771 1946
rect 112 1929 114 1945
rect 110 1928 116 1929
rect 448 1928 450 1945
rect 576 1928 578 1945
rect 712 1928 714 1945
rect 848 1928 850 1945
rect 984 1928 986 1945
rect 1120 1928 1122 1945
rect 1256 1928 1258 1945
rect 1384 1928 1386 1945
rect 1520 1928 1522 1945
rect 1656 1928 1658 1945
rect 1768 1929 1770 1945
rect 1806 1943 1812 1944
rect 1806 1939 1807 1943
rect 1811 1939 1812 1943
rect 3462 1943 3468 1944
rect 1806 1938 1812 1939
rect 1830 1940 1836 1941
rect 1766 1928 1772 1929
rect 110 1924 111 1928
rect 115 1924 116 1928
rect 110 1923 116 1924
rect 446 1927 452 1928
rect 446 1923 447 1927
rect 451 1923 452 1927
rect 446 1922 452 1923
rect 574 1927 580 1928
rect 574 1923 575 1927
rect 579 1923 580 1927
rect 574 1922 580 1923
rect 710 1927 716 1928
rect 710 1923 711 1927
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 846 1927 852 1928
rect 846 1923 847 1927
rect 851 1923 852 1927
rect 846 1922 852 1923
rect 982 1927 988 1928
rect 982 1923 983 1927
rect 987 1923 988 1927
rect 982 1922 988 1923
rect 1118 1927 1124 1928
rect 1118 1923 1119 1927
rect 1123 1923 1124 1927
rect 1118 1922 1124 1923
rect 1254 1927 1260 1928
rect 1254 1923 1255 1927
rect 1259 1923 1260 1927
rect 1254 1922 1260 1923
rect 1382 1927 1388 1928
rect 1382 1923 1383 1927
rect 1387 1923 1388 1927
rect 1382 1922 1388 1923
rect 1518 1927 1524 1928
rect 1518 1923 1519 1927
rect 1523 1923 1524 1927
rect 1518 1922 1524 1923
rect 1654 1927 1660 1928
rect 1654 1923 1655 1927
rect 1659 1923 1660 1927
rect 1766 1924 1767 1928
rect 1771 1924 1772 1928
rect 1766 1923 1772 1924
rect 1654 1922 1660 1923
rect 1808 1915 1810 1938
rect 1830 1936 1831 1940
rect 1835 1936 1836 1940
rect 1830 1935 1836 1936
rect 1918 1940 1924 1941
rect 1918 1936 1919 1940
rect 1923 1936 1924 1940
rect 1918 1935 1924 1936
rect 2046 1940 2052 1941
rect 2046 1936 2047 1940
rect 2051 1936 2052 1940
rect 2046 1935 2052 1936
rect 2182 1940 2188 1941
rect 2182 1936 2183 1940
rect 2187 1936 2188 1940
rect 2182 1935 2188 1936
rect 2326 1940 2332 1941
rect 2326 1936 2327 1940
rect 2331 1936 2332 1940
rect 2326 1935 2332 1936
rect 2470 1940 2476 1941
rect 2470 1936 2471 1940
rect 2475 1936 2476 1940
rect 2470 1935 2476 1936
rect 2614 1940 2620 1941
rect 2614 1936 2615 1940
rect 2619 1936 2620 1940
rect 2614 1935 2620 1936
rect 2750 1940 2756 1941
rect 2750 1936 2751 1940
rect 2755 1936 2756 1940
rect 2750 1935 2756 1936
rect 2886 1940 2892 1941
rect 2886 1936 2887 1940
rect 2891 1936 2892 1940
rect 2886 1935 2892 1936
rect 3030 1940 3036 1941
rect 3030 1936 3031 1940
rect 3035 1936 3036 1940
rect 3030 1935 3036 1936
rect 3174 1940 3180 1941
rect 3174 1936 3175 1940
rect 3179 1936 3180 1940
rect 3174 1935 3180 1936
rect 3318 1940 3324 1941
rect 3318 1936 3319 1940
rect 3323 1936 3324 1940
rect 3462 1939 3463 1943
rect 3467 1939 3468 1943
rect 3462 1938 3468 1939
rect 3318 1935 3324 1936
rect 1832 1915 1834 1935
rect 1920 1915 1922 1935
rect 2048 1915 2050 1935
rect 2184 1915 2186 1935
rect 2328 1915 2330 1935
rect 2472 1915 2474 1935
rect 2616 1915 2618 1935
rect 2752 1915 2754 1935
rect 2888 1915 2890 1935
rect 3032 1915 3034 1935
rect 3176 1915 3178 1935
rect 3320 1915 3322 1935
rect 3464 1915 3466 1938
rect 1807 1914 1811 1915
rect 110 1911 116 1912
rect 110 1907 111 1911
rect 115 1907 116 1911
rect 1766 1911 1772 1912
rect 110 1906 116 1907
rect 446 1908 452 1909
rect 112 1887 114 1906
rect 446 1904 447 1908
rect 451 1904 452 1908
rect 446 1903 452 1904
rect 574 1908 580 1909
rect 574 1904 575 1908
rect 579 1904 580 1908
rect 574 1903 580 1904
rect 710 1908 716 1909
rect 710 1904 711 1908
rect 715 1904 716 1908
rect 710 1903 716 1904
rect 846 1908 852 1909
rect 846 1904 847 1908
rect 851 1904 852 1908
rect 846 1903 852 1904
rect 982 1908 988 1909
rect 982 1904 983 1908
rect 987 1904 988 1908
rect 982 1903 988 1904
rect 1118 1908 1124 1909
rect 1118 1904 1119 1908
rect 1123 1904 1124 1908
rect 1118 1903 1124 1904
rect 1254 1908 1260 1909
rect 1254 1904 1255 1908
rect 1259 1904 1260 1908
rect 1254 1903 1260 1904
rect 1382 1908 1388 1909
rect 1382 1904 1383 1908
rect 1387 1904 1388 1908
rect 1382 1903 1388 1904
rect 1518 1908 1524 1909
rect 1518 1904 1519 1908
rect 1523 1904 1524 1908
rect 1518 1903 1524 1904
rect 1654 1908 1660 1909
rect 1654 1904 1655 1908
rect 1659 1904 1660 1908
rect 1766 1907 1767 1911
rect 1771 1907 1772 1911
rect 1807 1909 1811 1910
rect 1831 1914 1835 1915
rect 1831 1909 1835 1910
rect 1919 1914 1923 1915
rect 1919 1909 1923 1910
rect 2039 1914 2043 1915
rect 2039 1909 2043 1910
rect 2047 1914 2051 1915
rect 2047 1909 2051 1910
rect 2167 1914 2171 1915
rect 2167 1909 2171 1910
rect 2183 1914 2187 1915
rect 2183 1909 2187 1910
rect 2303 1914 2307 1915
rect 2303 1909 2307 1910
rect 2327 1914 2331 1915
rect 2327 1909 2331 1910
rect 2455 1914 2459 1915
rect 2455 1909 2459 1910
rect 2471 1914 2475 1915
rect 2471 1909 2475 1910
rect 2615 1914 2619 1915
rect 2615 1909 2619 1910
rect 2751 1914 2755 1915
rect 2751 1909 2755 1910
rect 2791 1914 2795 1915
rect 2791 1909 2795 1910
rect 2887 1914 2891 1915
rect 2887 1909 2891 1910
rect 2983 1914 2987 1915
rect 2983 1909 2987 1910
rect 3031 1914 3035 1915
rect 3031 1909 3035 1910
rect 3175 1914 3179 1915
rect 3175 1909 3179 1910
rect 3183 1914 3187 1915
rect 3183 1909 3187 1910
rect 3319 1914 3323 1915
rect 3319 1909 3323 1910
rect 3367 1914 3371 1915
rect 3367 1909 3371 1910
rect 3463 1914 3467 1915
rect 3463 1909 3467 1910
rect 1766 1906 1772 1907
rect 1654 1903 1660 1904
rect 448 1887 450 1903
rect 576 1887 578 1903
rect 712 1887 714 1903
rect 848 1887 850 1903
rect 984 1887 986 1903
rect 1120 1887 1122 1903
rect 1256 1887 1258 1903
rect 1384 1887 1386 1903
rect 1520 1887 1522 1903
rect 1656 1887 1658 1903
rect 1768 1887 1770 1906
rect 1808 1890 1810 1909
rect 1832 1893 1834 1909
rect 1920 1893 1922 1909
rect 2040 1893 2042 1909
rect 2168 1893 2170 1909
rect 2304 1893 2306 1909
rect 2456 1893 2458 1909
rect 2616 1893 2618 1909
rect 2792 1893 2794 1909
rect 2984 1893 2986 1909
rect 3184 1893 3186 1909
rect 3368 1893 3370 1909
rect 1830 1892 1836 1893
rect 1806 1889 1812 1890
rect 111 1886 115 1887
rect 111 1881 115 1882
rect 447 1886 451 1887
rect 447 1881 451 1882
rect 559 1886 563 1887
rect 559 1881 563 1882
rect 575 1886 579 1887
rect 575 1881 579 1882
rect 695 1886 699 1887
rect 695 1881 699 1882
rect 711 1886 715 1887
rect 711 1881 715 1882
rect 831 1886 835 1887
rect 831 1881 835 1882
rect 847 1886 851 1887
rect 847 1881 851 1882
rect 959 1886 963 1887
rect 959 1881 963 1882
rect 983 1886 987 1887
rect 983 1881 987 1882
rect 1079 1886 1083 1887
rect 1079 1881 1083 1882
rect 1119 1886 1123 1887
rect 1119 1881 1123 1882
rect 1199 1886 1203 1887
rect 1199 1881 1203 1882
rect 1255 1886 1259 1887
rect 1255 1881 1259 1882
rect 1327 1886 1331 1887
rect 1327 1881 1331 1882
rect 1383 1886 1387 1887
rect 1383 1881 1387 1882
rect 1455 1886 1459 1887
rect 1455 1881 1459 1882
rect 1519 1886 1523 1887
rect 1519 1881 1523 1882
rect 1655 1886 1659 1887
rect 1655 1881 1659 1882
rect 1767 1886 1771 1887
rect 1806 1885 1807 1889
rect 1811 1885 1812 1889
rect 1830 1888 1831 1892
rect 1835 1888 1836 1892
rect 1830 1887 1836 1888
rect 1918 1892 1924 1893
rect 1918 1888 1919 1892
rect 1923 1888 1924 1892
rect 1918 1887 1924 1888
rect 2038 1892 2044 1893
rect 2038 1888 2039 1892
rect 2043 1888 2044 1892
rect 2038 1887 2044 1888
rect 2166 1892 2172 1893
rect 2166 1888 2167 1892
rect 2171 1888 2172 1892
rect 2166 1887 2172 1888
rect 2302 1892 2308 1893
rect 2302 1888 2303 1892
rect 2307 1888 2308 1892
rect 2302 1887 2308 1888
rect 2454 1892 2460 1893
rect 2454 1888 2455 1892
rect 2459 1888 2460 1892
rect 2454 1887 2460 1888
rect 2614 1892 2620 1893
rect 2614 1888 2615 1892
rect 2619 1888 2620 1892
rect 2614 1887 2620 1888
rect 2790 1892 2796 1893
rect 2790 1888 2791 1892
rect 2795 1888 2796 1892
rect 2790 1887 2796 1888
rect 2982 1892 2988 1893
rect 2982 1888 2983 1892
rect 2987 1888 2988 1892
rect 2982 1887 2988 1888
rect 3182 1892 3188 1893
rect 3182 1888 3183 1892
rect 3187 1888 3188 1892
rect 3182 1887 3188 1888
rect 3366 1892 3372 1893
rect 3366 1888 3367 1892
rect 3371 1888 3372 1892
rect 3464 1890 3466 1909
rect 3366 1887 3372 1888
rect 3462 1889 3468 1890
rect 1806 1884 1812 1885
rect 3462 1885 3463 1889
rect 3467 1885 3468 1889
rect 3462 1884 3468 1885
rect 1767 1881 1771 1882
rect 112 1862 114 1881
rect 560 1865 562 1881
rect 696 1865 698 1881
rect 832 1865 834 1881
rect 960 1865 962 1881
rect 1080 1865 1082 1881
rect 1200 1865 1202 1881
rect 1328 1865 1330 1881
rect 1456 1865 1458 1881
rect 558 1864 564 1865
rect 110 1861 116 1862
rect 110 1857 111 1861
rect 115 1857 116 1861
rect 558 1860 559 1864
rect 563 1860 564 1864
rect 558 1859 564 1860
rect 694 1864 700 1865
rect 694 1860 695 1864
rect 699 1860 700 1864
rect 694 1859 700 1860
rect 830 1864 836 1865
rect 830 1860 831 1864
rect 835 1860 836 1864
rect 830 1859 836 1860
rect 958 1864 964 1865
rect 958 1860 959 1864
rect 963 1860 964 1864
rect 958 1859 964 1860
rect 1078 1864 1084 1865
rect 1078 1860 1079 1864
rect 1083 1860 1084 1864
rect 1078 1859 1084 1860
rect 1198 1864 1204 1865
rect 1198 1860 1199 1864
rect 1203 1860 1204 1864
rect 1198 1859 1204 1860
rect 1326 1864 1332 1865
rect 1326 1860 1327 1864
rect 1331 1860 1332 1864
rect 1326 1859 1332 1860
rect 1454 1864 1460 1865
rect 1454 1860 1455 1864
rect 1459 1860 1460 1864
rect 1768 1862 1770 1881
rect 1830 1873 1836 1874
rect 1806 1872 1812 1873
rect 1806 1868 1807 1872
rect 1811 1868 1812 1872
rect 1830 1869 1831 1873
rect 1835 1869 1836 1873
rect 1830 1868 1836 1869
rect 1918 1873 1924 1874
rect 1918 1869 1919 1873
rect 1923 1869 1924 1873
rect 1918 1868 1924 1869
rect 2038 1873 2044 1874
rect 2038 1869 2039 1873
rect 2043 1869 2044 1873
rect 2038 1868 2044 1869
rect 2166 1873 2172 1874
rect 2166 1869 2167 1873
rect 2171 1869 2172 1873
rect 2166 1868 2172 1869
rect 2302 1873 2308 1874
rect 2302 1869 2303 1873
rect 2307 1869 2308 1873
rect 2302 1868 2308 1869
rect 2454 1873 2460 1874
rect 2454 1869 2455 1873
rect 2459 1869 2460 1873
rect 2454 1868 2460 1869
rect 2614 1873 2620 1874
rect 2614 1869 2615 1873
rect 2619 1869 2620 1873
rect 2614 1868 2620 1869
rect 2790 1873 2796 1874
rect 2790 1869 2791 1873
rect 2795 1869 2796 1873
rect 2790 1868 2796 1869
rect 2982 1873 2988 1874
rect 2982 1869 2983 1873
rect 2987 1869 2988 1873
rect 2982 1868 2988 1869
rect 3182 1873 3188 1874
rect 3182 1869 3183 1873
rect 3187 1869 3188 1873
rect 3182 1868 3188 1869
rect 3366 1873 3372 1874
rect 3366 1869 3367 1873
rect 3371 1869 3372 1873
rect 3366 1868 3372 1869
rect 3462 1872 3468 1873
rect 3462 1868 3463 1872
rect 3467 1868 3468 1872
rect 1806 1867 1812 1868
rect 1454 1859 1460 1860
rect 1766 1861 1772 1862
rect 110 1856 116 1857
rect 1766 1857 1767 1861
rect 1771 1857 1772 1861
rect 1766 1856 1772 1857
rect 1808 1847 1810 1867
rect 1832 1847 1834 1868
rect 1920 1847 1922 1868
rect 2040 1847 2042 1868
rect 2168 1847 2170 1868
rect 2304 1847 2306 1868
rect 2456 1847 2458 1868
rect 2616 1847 2618 1868
rect 2792 1847 2794 1868
rect 2984 1847 2986 1868
rect 3184 1847 3186 1868
rect 3368 1847 3370 1868
rect 3462 1867 3468 1868
rect 3464 1847 3466 1867
rect 1807 1846 1811 1847
rect 558 1845 564 1846
rect 110 1844 116 1845
rect 110 1840 111 1844
rect 115 1840 116 1844
rect 558 1841 559 1845
rect 563 1841 564 1845
rect 558 1840 564 1841
rect 694 1845 700 1846
rect 694 1841 695 1845
rect 699 1841 700 1845
rect 694 1840 700 1841
rect 830 1845 836 1846
rect 830 1841 831 1845
rect 835 1841 836 1845
rect 830 1840 836 1841
rect 958 1845 964 1846
rect 958 1841 959 1845
rect 963 1841 964 1845
rect 958 1840 964 1841
rect 1078 1845 1084 1846
rect 1078 1841 1079 1845
rect 1083 1841 1084 1845
rect 1078 1840 1084 1841
rect 1198 1845 1204 1846
rect 1198 1841 1199 1845
rect 1203 1841 1204 1845
rect 1198 1840 1204 1841
rect 1326 1845 1332 1846
rect 1326 1841 1327 1845
rect 1331 1841 1332 1845
rect 1326 1840 1332 1841
rect 1454 1845 1460 1846
rect 1454 1841 1455 1845
rect 1459 1841 1460 1845
rect 1454 1840 1460 1841
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1807 1841 1811 1842
rect 1831 1846 1835 1847
rect 1831 1841 1835 1842
rect 1919 1846 1923 1847
rect 1919 1841 1923 1842
rect 1959 1846 1963 1847
rect 1959 1841 1963 1842
rect 2039 1846 2043 1847
rect 2039 1841 2043 1842
rect 2111 1846 2115 1847
rect 2111 1841 2115 1842
rect 2167 1846 2171 1847
rect 2167 1841 2171 1842
rect 2255 1846 2259 1847
rect 2255 1841 2259 1842
rect 2303 1846 2307 1847
rect 2303 1841 2307 1842
rect 2407 1846 2411 1847
rect 2407 1841 2411 1842
rect 2455 1846 2459 1847
rect 2455 1841 2459 1842
rect 2567 1846 2571 1847
rect 2567 1841 2571 1842
rect 2615 1846 2619 1847
rect 2615 1841 2619 1842
rect 2743 1846 2747 1847
rect 2743 1841 2747 1842
rect 2791 1846 2795 1847
rect 2791 1841 2795 1842
rect 2935 1846 2939 1847
rect 2935 1841 2939 1842
rect 2983 1846 2987 1847
rect 2983 1841 2987 1842
rect 3135 1846 3139 1847
rect 3135 1841 3139 1842
rect 3183 1846 3187 1847
rect 3183 1841 3187 1842
rect 3343 1846 3347 1847
rect 3343 1841 3347 1842
rect 3367 1846 3371 1847
rect 3367 1841 3371 1842
rect 3463 1846 3467 1847
rect 3463 1841 3467 1842
rect 110 1839 116 1840
rect 112 1815 114 1839
rect 560 1815 562 1840
rect 696 1815 698 1840
rect 832 1815 834 1840
rect 960 1815 962 1840
rect 1080 1815 1082 1840
rect 1200 1815 1202 1840
rect 1328 1815 1330 1840
rect 1456 1815 1458 1840
rect 1766 1839 1772 1840
rect 1768 1815 1770 1839
rect 1808 1825 1810 1841
rect 1806 1824 1812 1825
rect 1832 1824 1834 1841
rect 1960 1824 1962 1841
rect 2112 1824 2114 1841
rect 2256 1824 2258 1841
rect 2408 1824 2410 1841
rect 2568 1824 2570 1841
rect 2744 1824 2746 1841
rect 2936 1824 2938 1841
rect 3136 1824 3138 1841
rect 3344 1824 3346 1841
rect 3464 1825 3466 1841
rect 3462 1824 3468 1825
rect 1806 1820 1807 1824
rect 1811 1820 1812 1824
rect 1806 1819 1812 1820
rect 1830 1823 1836 1824
rect 1830 1819 1831 1823
rect 1835 1819 1836 1823
rect 1830 1818 1836 1819
rect 1958 1823 1964 1824
rect 1958 1819 1959 1823
rect 1963 1819 1964 1823
rect 1958 1818 1964 1819
rect 2110 1823 2116 1824
rect 2110 1819 2111 1823
rect 2115 1819 2116 1823
rect 2110 1818 2116 1819
rect 2254 1823 2260 1824
rect 2254 1819 2255 1823
rect 2259 1819 2260 1823
rect 2254 1818 2260 1819
rect 2406 1823 2412 1824
rect 2406 1819 2407 1823
rect 2411 1819 2412 1823
rect 2406 1818 2412 1819
rect 2566 1823 2572 1824
rect 2566 1819 2567 1823
rect 2571 1819 2572 1823
rect 2566 1818 2572 1819
rect 2742 1823 2748 1824
rect 2742 1819 2743 1823
rect 2747 1819 2748 1823
rect 2742 1818 2748 1819
rect 2934 1823 2940 1824
rect 2934 1819 2935 1823
rect 2939 1819 2940 1823
rect 2934 1818 2940 1819
rect 3134 1823 3140 1824
rect 3134 1819 3135 1823
rect 3139 1819 3140 1823
rect 3134 1818 3140 1819
rect 3342 1823 3348 1824
rect 3342 1819 3343 1823
rect 3347 1819 3348 1823
rect 3462 1820 3463 1824
rect 3467 1820 3468 1824
rect 3462 1819 3468 1820
rect 3342 1818 3348 1819
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 135 1814 139 1815
rect 135 1809 139 1810
rect 223 1814 227 1815
rect 223 1809 227 1810
rect 311 1814 315 1815
rect 311 1809 315 1810
rect 407 1814 411 1815
rect 407 1809 411 1810
rect 527 1814 531 1815
rect 527 1809 531 1810
rect 559 1814 563 1815
rect 559 1809 563 1810
rect 655 1814 659 1815
rect 655 1809 659 1810
rect 695 1814 699 1815
rect 695 1809 699 1810
rect 799 1814 803 1815
rect 799 1809 803 1810
rect 831 1814 835 1815
rect 831 1809 835 1810
rect 943 1814 947 1815
rect 943 1809 947 1810
rect 959 1814 963 1815
rect 959 1809 963 1810
rect 1079 1814 1083 1815
rect 1079 1809 1083 1810
rect 1087 1814 1091 1815
rect 1087 1809 1091 1810
rect 1199 1814 1203 1815
rect 1199 1809 1203 1810
rect 1239 1814 1243 1815
rect 1239 1809 1243 1810
rect 1327 1814 1331 1815
rect 1327 1809 1331 1810
rect 1391 1814 1395 1815
rect 1391 1809 1395 1810
rect 1455 1814 1459 1815
rect 1455 1809 1459 1810
rect 1543 1814 1547 1815
rect 1543 1809 1547 1810
rect 1671 1814 1675 1815
rect 1671 1809 1675 1810
rect 1767 1814 1771 1815
rect 1767 1809 1771 1810
rect 112 1793 114 1809
rect 110 1792 116 1793
rect 136 1792 138 1809
rect 224 1792 226 1809
rect 312 1792 314 1809
rect 408 1792 410 1809
rect 528 1792 530 1809
rect 656 1792 658 1809
rect 800 1792 802 1809
rect 944 1792 946 1809
rect 1088 1792 1090 1809
rect 1240 1792 1242 1809
rect 1392 1792 1394 1809
rect 1544 1792 1546 1809
rect 1672 1792 1674 1809
rect 1768 1793 1770 1809
rect 1806 1807 1812 1808
rect 1806 1803 1807 1807
rect 1811 1803 1812 1807
rect 3462 1807 3468 1808
rect 1806 1802 1812 1803
rect 1830 1804 1836 1805
rect 1766 1792 1772 1793
rect 110 1788 111 1792
rect 115 1788 116 1792
rect 110 1787 116 1788
rect 134 1791 140 1792
rect 134 1787 135 1791
rect 139 1787 140 1791
rect 134 1786 140 1787
rect 222 1791 228 1792
rect 222 1787 223 1791
rect 227 1787 228 1791
rect 222 1786 228 1787
rect 310 1791 316 1792
rect 310 1787 311 1791
rect 315 1787 316 1791
rect 310 1786 316 1787
rect 406 1791 412 1792
rect 406 1787 407 1791
rect 411 1787 412 1791
rect 406 1786 412 1787
rect 526 1791 532 1792
rect 526 1787 527 1791
rect 531 1787 532 1791
rect 526 1786 532 1787
rect 654 1791 660 1792
rect 654 1787 655 1791
rect 659 1787 660 1791
rect 654 1786 660 1787
rect 798 1791 804 1792
rect 798 1787 799 1791
rect 803 1787 804 1791
rect 798 1786 804 1787
rect 942 1791 948 1792
rect 942 1787 943 1791
rect 947 1787 948 1791
rect 942 1786 948 1787
rect 1086 1791 1092 1792
rect 1086 1787 1087 1791
rect 1091 1787 1092 1791
rect 1086 1786 1092 1787
rect 1238 1791 1244 1792
rect 1238 1787 1239 1791
rect 1243 1787 1244 1791
rect 1238 1786 1244 1787
rect 1390 1791 1396 1792
rect 1390 1787 1391 1791
rect 1395 1787 1396 1791
rect 1390 1786 1396 1787
rect 1542 1791 1548 1792
rect 1542 1787 1543 1791
rect 1547 1787 1548 1791
rect 1542 1786 1548 1787
rect 1670 1791 1676 1792
rect 1670 1787 1671 1791
rect 1675 1787 1676 1791
rect 1766 1788 1767 1792
rect 1771 1788 1772 1792
rect 1766 1787 1772 1788
rect 1670 1786 1676 1787
rect 110 1775 116 1776
rect 110 1771 111 1775
rect 115 1771 116 1775
rect 1766 1775 1772 1776
rect 110 1770 116 1771
rect 134 1772 140 1773
rect 112 1739 114 1770
rect 134 1768 135 1772
rect 139 1768 140 1772
rect 134 1767 140 1768
rect 222 1772 228 1773
rect 222 1768 223 1772
rect 227 1768 228 1772
rect 222 1767 228 1768
rect 310 1772 316 1773
rect 310 1768 311 1772
rect 315 1768 316 1772
rect 310 1767 316 1768
rect 406 1772 412 1773
rect 406 1768 407 1772
rect 411 1768 412 1772
rect 406 1767 412 1768
rect 526 1772 532 1773
rect 526 1768 527 1772
rect 531 1768 532 1772
rect 526 1767 532 1768
rect 654 1772 660 1773
rect 654 1768 655 1772
rect 659 1768 660 1772
rect 654 1767 660 1768
rect 798 1772 804 1773
rect 798 1768 799 1772
rect 803 1768 804 1772
rect 798 1767 804 1768
rect 942 1772 948 1773
rect 942 1768 943 1772
rect 947 1768 948 1772
rect 942 1767 948 1768
rect 1086 1772 1092 1773
rect 1086 1768 1087 1772
rect 1091 1768 1092 1772
rect 1086 1767 1092 1768
rect 1238 1772 1244 1773
rect 1238 1768 1239 1772
rect 1243 1768 1244 1772
rect 1238 1767 1244 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1542 1772 1548 1773
rect 1542 1768 1543 1772
rect 1547 1768 1548 1772
rect 1542 1767 1548 1768
rect 1670 1772 1676 1773
rect 1670 1768 1671 1772
rect 1675 1768 1676 1772
rect 1766 1771 1767 1775
rect 1771 1771 1772 1775
rect 1808 1771 1810 1802
rect 1830 1800 1831 1804
rect 1835 1800 1836 1804
rect 1830 1799 1836 1800
rect 1958 1804 1964 1805
rect 1958 1800 1959 1804
rect 1963 1800 1964 1804
rect 1958 1799 1964 1800
rect 2110 1804 2116 1805
rect 2110 1800 2111 1804
rect 2115 1800 2116 1804
rect 2110 1799 2116 1800
rect 2254 1804 2260 1805
rect 2254 1800 2255 1804
rect 2259 1800 2260 1804
rect 2254 1799 2260 1800
rect 2406 1804 2412 1805
rect 2406 1800 2407 1804
rect 2411 1800 2412 1804
rect 2406 1799 2412 1800
rect 2566 1804 2572 1805
rect 2566 1800 2567 1804
rect 2571 1800 2572 1804
rect 2566 1799 2572 1800
rect 2742 1804 2748 1805
rect 2742 1800 2743 1804
rect 2747 1800 2748 1804
rect 2742 1799 2748 1800
rect 2934 1804 2940 1805
rect 2934 1800 2935 1804
rect 2939 1800 2940 1804
rect 2934 1799 2940 1800
rect 3134 1804 3140 1805
rect 3134 1800 3135 1804
rect 3139 1800 3140 1804
rect 3134 1799 3140 1800
rect 3342 1804 3348 1805
rect 3342 1800 3343 1804
rect 3347 1800 3348 1804
rect 3462 1803 3463 1807
rect 3467 1803 3468 1807
rect 3462 1802 3468 1803
rect 3342 1799 3348 1800
rect 1832 1771 1834 1799
rect 1960 1771 1962 1799
rect 2112 1771 2114 1799
rect 2256 1771 2258 1799
rect 2408 1771 2410 1799
rect 2568 1771 2570 1799
rect 2744 1771 2746 1799
rect 2936 1771 2938 1799
rect 3136 1771 3138 1799
rect 3344 1771 3346 1799
rect 3464 1771 3466 1802
rect 1766 1770 1772 1771
rect 1807 1770 1811 1771
rect 1670 1767 1676 1768
rect 136 1739 138 1767
rect 224 1739 226 1767
rect 312 1739 314 1767
rect 408 1739 410 1767
rect 528 1739 530 1767
rect 656 1739 658 1767
rect 800 1739 802 1767
rect 944 1739 946 1767
rect 1088 1739 1090 1767
rect 1240 1739 1242 1767
rect 1392 1739 1394 1767
rect 1544 1739 1546 1767
rect 1672 1739 1674 1767
rect 1768 1739 1770 1770
rect 1807 1765 1811 1766
rect 1831 1770 1835 1771
rect 1831 1765 1835 1766
rect 1879 1770 1883 1771
rect 1879 1765 1883 1766
rect 1959 1770 1963 1771
rect 1959 1765 1963 1766
rect 2015 1770 2019 1771
rect 2015 1765 2019 1766
rect 2111 1770 2115 1771
rect 2111 1765 2115 1766
rect 2151 1770 2155 1771
rect 2151 1765 2155 1766
rect 2255 1770 2259 1771
rect 2255 1765 2259 1766
rect 2303 1770 2307 1771
rect 2303 1765 2307 1766
rect 2407 1770 2411 1771
rect 2407 1765 2411 1766
rect 2479 1770 2483 1771
rect 2479 1765 2483 1766
rect 2567 1770 2571 1771
rect 2567 1765 2571 1766
rect 2687 1770 2691 1771
rect 2687 1765 2691 1766
rect 2743 1770 2747 1771
rect 2743 1765 2747 1766
rect 2911 1770 2915 1771
rect 2911 1765 2915 1766
rect 2935 1770 2939 1771
rect 2935 1765 2939 1766
rect 3135 1770 3139 1771
rect 3135 1765 3139 1766
rect 3151 1770 3155 1771
rect 3151 1765 3155 1766
rect 3343 1770 3347 1771
rect 3343 1765 3347 1766
rect 3367 1770 3371 1771
rect 3367 1765 3371 1766
rect 3463 1770 3467 1771
rect 3463 1765 3467 1766
rect 1808 1746 1810 1765
rect 1880 1749 1882 1765
rect 2016 1749 2018 1765
rect 2152 1749 2154 1765
rect 2304 1749 2306 1765
rect 2480 1749 2482 1765
rect 2688 1749 2690 1765
rect 2912 1749 2914 1765
rect 3152 1749 3154 1765
rect 3368 1749 3370 1765
rect 1878 1748 1884 1749
rect 1806 1745 1812 1746
rect 1806 1741 1807 1745
rect 1811 1741 1812 1745
rect 1878 1744 1879 1748
rect 1883 1744 1884 1748
rect 1878 1743 1884 1744
rect 2014 1748 2020 1749
rect 2014 1744 2015 1748
rect 2019 1744 2020 1748
rect 2014 1743 2020 1744
rect 2150 1748 2156 1749
rect 2150 1744 2151 1748
rect 2155 1744 2156 1748
rect 2150 1743 2156 1744
rect 2302 1748 2308 1749
rect 2302 1744 2303 1748
rect 2307 1744 2308 1748
rect 2302 1743 2308 1744
rect 2478 1748 2484 1749
rect 2478 1744 2479 1748
rect 2483 1744 2484 1748
rect 2478 1743 2484 1744
rect 2686 1748 2692 1749
rect 2686 1744 2687 1748
rect 2691 1744 2692 1748
rect 2686 1743 2692 1744
rect 2910 1748 2916 1749
rect 2910 1744 2911 1748
rect 2915 1744 2916 1748
rect 2910 1743 2916 1744
rect 3150 1748 3156 1749
rect 3150 1744 3151 1748
rect 3155 1744 3156 1748
rect 3150 1743 3156 1744
rect 3366 1748 3372 1749
rect 3366 1744 3367 1748
rect 3371 1744 3372 1748
rect 3464 1746 3466 1765
rect 3366 1743 3372 1744
rect 3462 1745 3468 1746
rect 1806 1740 1812 1741
rect 3462 1741 3463 1745
rect 3467 1741 3468 1745
rect 3462 1740 3468 1741
rect 111 1738 115 1739
rect 111 1733 115 1734
rect 135 1738 139 1739
rect 135 1733 139 1734
rect 223 1738 227 1739
rect 223 1733 227 1734
rect 247 1738 251 1739
rect 247 1733 251 1734
rect 311 1738 315 1739
rect 311 1733 315 1734
rect 399 1738 403 1739
rect 399 1733 403 1734
rect 407 1738 411 1739
rect 407 1733 411 1734
rect 527 1738 531 1739
rect 527 1733 531 1734
rect 567 1738 571 1739
rect 567 1733 571 1734
rect 655 1738 659 1739
rect 655 1733 659 1734
rect 751 1738 755 1739
rect 751 1733 755 1734
rect 799 1738 803 1739
rect 799 1733 803 1734
rect 935 1738 939 1739
rect 935 1733 939 1734
rect 943 1738 947 1739
rect 943 1733 947 1734
rect 1087 1738 1091 1739
rect 1087 1733 1091 1734
rect 1119 1738 1123 1739
rect 1119 1733 1123 1734
rect 1239 1738 1243 1739
rect 1239 1733 1243 1734
rect 1311 1738 1315 1739
rect 1311 1733 1315 1734
rect 1391 1738 1395 1739
rect 1391 1733 1395 1734
rect 1503 1738 1507 1739
rect 1503 1733 1507 1734
rect 1543 1738 1547 1739
rect 1543 1733 1547 1734
rect 1671 1738 1675 1739
rect 1671 1733 1675 1734
rect 1767 1738 1771 1739
rect 1767 1733 1771 1734
rect 112 1714 114 1733
rect 136 1717 138 1733
rect 248 1717 250 1733
rect 400 1717 402 1733
rect 568 1717 570 1733
rect 752 1717 754 1733
rect 936 1717 938 1733
rect 1120 1717 1122 1733
rect 1312 1717 1314 1733
rect 1504 1717 1506 1733
rect 1672 1717 1674 1733
rect 134 1716 140 1717
rect 110 1713 116 1714
rect 110 1709 111 1713
rect 115 1709 116 1713
rect 134 1712 135 1716
rect 139 1712 140 1716
rect 134 1711 140 1712
rect 246 1716 252 1717
rect 246 1712 247 1716
rect 251 1712 252 1716
rect 246 1711 252 1712
rect 398 1716 404 1717
rect 398 1712 399 1716
rect 403 1712 404 1716
rect 398 1711 404 1712
rect 566 1716 572 1717
rect 566 1712 567 1716
rect 571 1712 572 1716
rect 566 1711 572 1712
rect 750 1716 756 1717
rect 750 1712 751 1716
rect 755 1712 756 1716
rect 750 1711 756 1712
rect 934 1716 940 1717
rect 934 1712 935 1716
rect 939 1712 940 1716
rect 934 1711 940 1712
rect 1118 1716 1124 1717
rect 1118 1712 1119 1716
rect 1123 1712 1124 1716
rect 1118 1711 1124 1712
rect 1310 1716 1316 1717
rect 1310 1712 1311 1716
rect 1315 1712 1316 1716
rect 1310 1711 1316 1712
rect 1502 1716 1508 1717
rect 1502 1712 1503 1716
rect 1507 1712 1508 1716
rect 1502 1711 1508 1712
rect 1670 1716 1676 1717
rect 1670 1712 1671 1716
rect 1675 1712 1676 1716
rect 1768 1714 1770 1733
rect 1878 1729 1884 1730
rect 1806 1728 1812 1729
rect 1806 1724 1807 1728
rect 1811 1724 1812 1728
rect 1878 1725 1879 1729
rect 1883 1725 1884 1729
rect 1878 1724 1884 1725
rect 2014 1729 2020 1730
rect 2014 1725 2015 1729
rect 2019 1725 2020 1729
rect 2014 1724 2020 1725
rect 2150 1729 2156 1730
rect 2150 1725 2151 1729
rect 2155 1725 2156 1729
rect 2150 1724 2156 1725
rect 2302 1729 2308 1730
rect 2302 1725 2303 1729
rect 2307 1725 2308 1729
rect 2302 1724 2308 1725
rect 2478 1729 2484 1730
rect 2478 1725 2479 1729
rect 2483 1725 2484 1729
rect 2478 1724 2484 1725
rect 2686 1729 2692 1730
rect 2686 1725 2687 1729
rect 2691 1725 2692 1729
rect 2686 1724 2692 1725
rect 2910 1729 2916 1730
rect 2910 1725 2911 1729
rect 2915 1725 2916 1729
rect 2910 1724 2916 1725
rect 3150 1729 3156 1730
rect 3150 1725 3151 1729
rect 3155 1725 3156 1729
rect 3150 1724 3156 1725
rect 3366 1729 3372 1730
rect 3366 1725 3367 1729
rect 3371 1725 3372 1729
rect 3366 1724 3372 1725
rect 3462 1728 3468 1729
rect 3462 1724 3463 1728
rect 3467 1724 3468 1728
rect 1806 1723 1812 1724
rect 1670 1711 1676 1712
rect 1766 1713 1772 1714
rect 110 1708 116 1709
rect 1766 1709 1767 1713
rect 1771 1709 1772 1713
rect 1766 1708 1772 1709
rect 1808 1699 1810 1723
rect 1880 1699 1882 1724
rect 2016 1699 2018 1724
rect 2152 1699 2154 1724
rect 2304 1699 2306 1724
rect 2480 1699 2482 1724
rect 2688 1699 2690 1724
rect 2912 1699 2914 1724
rect 3152 1699 3154 1724
rect 3368 1699 3370 1724
rect 3462 1723 3468 1724
rect 3464 1699 3466 1723
rect 1807 1698 1811 1699
rect 134 1697 140 1698
rect 110 1696 116 1697
rect 110 1692 111 1696
rect 115 1692 116 1696
rect 134 1693 135 1697
rect 139 1693 140 1697
rect 134 1692 140 1693
rect 246 1697 252 1698
rect 246 1693 247 1697
rect 251 1693 252 1697
rect 246 1692 252 1693
rect 398 1697 404 1698
rect 398 1693 399 1697
rect 403 1693 404 1697
rect 398 1692 404 1693
rect 566 1697 572 1698
rect 566 1693 567 1697
rect 571 1693 572 1697
rect 566 1692 572 1693
rect 750 1697 756 1698
rect 750 1693 751 1697
rect 755 1693 756 1697
rect 750 1692 756 1693
rect 934 1697 940 1698
rect 934 1693 935 1697
rect 939 1693 940 1697
rect 934 1692 940 1693
rect 1118 1697 1124 1698
rect 1118 1693 1119 1697
rect 1123 1693 1124 1697
rect 1118 1692 1124 1693
rect 1310 1697 1316 1698
rect 1310 1693 1311 1697
rect 1315 1693 1316 1697
rect 1310 1692 1316 1693
rect 1502 1697 1508 1698
rect 1502 1693 1503 1697
rect 1507 1693 1508 1697
rect 1502 1692 1508 1693
rect 1670 1697 1676 1698
rect 1670 1693 1671 1697
rect 1675 1693 1676 1697
rect 1670 1692 1676 1693
rect 1766 1696 1772 1697
rect 1766 1692 1767 1696
rect 1771 1692 1772 1696
rect 1807 1693 1811 1694
rect 1831 1698 1835 1699
rect 1831 1693 1835 1694
rect 1879 1698 1883 1699
rect 1879 1693 1883 1694
rect 1935 1698 1939 1699
rect 1935 1693 1939 1694
rect 2015 1698 2019 1699
rect 2015 1693 2019 1694
rect 2063 1698 2067 1699
rect 2063 1693 2067 1694
rect 2151 1698 2155 1699
rect 2151 1693 2155 1694
rect 2183 1698 2187 1699
rect 2183 1693 2187 1694
rect 2303 1698 2307 1699
rect 2303 1693 2307 1694
rect 2311 1698 2315 1699
rect 2311 1693 2315 1694
rect 2439 1698 2443 1699
rect 2439 1693 2443 1694
rect 2479 1698 2483 1699
rect 2479 1693 2483 1694
rect 2575 1698 2579 1699
rect 2575 1693 2579 1694
rect 2687 1698 2691 1699
rect 2687 1693 2691 1694
rect 2727 1698 2731 1699
rect 2727 1693 2731 1694
rect 2887 1698 2891 1699
rect 2887 1693 2891 1694
rect 2911 1698 2915 1699
rect 2911 1693 2915 1694
rect 3047 1698 3051 1699
rect 3047 1693 3051 1694
rect 3151 1698 3155 1699
rect 3151 1693 3155 1694
rect 3215 1698 3219 1699
rect 3215 1693 3219 1694
rect 3367 1698 3371 1699
rect 3367 1693 3371 1694
rect 3463 1698 3467 1699
rect 3463 1693 3467 1694
rect 110 1691 116 1692
rect 112 1671 114 1691
rect 136 1671 138 1692
rect 248 1671 250 1692
rect 400 1671 402 1692
rect 568 1671 570 1692
rect 752 1671 754 1692
rect 936 1671 938 1692
rect 1120 1671 1122 1692
rect 1312 1671 1314 1692
rect 1504 1671 1506 1692
rect 1672 1671 1674 1692
rect 1766 1691 1772 1692
rect 1768 1671 1770 1691
rect 1808 1677 1810 1693
rect 1806 1676 1812 1677
rect 1832 1676 1834 1693
rect 1936 1676 1938 1693
rect 2064 1676 2066 1693
rect 2184 1676 2186 1693
rect 2312 1676 2314 1693
rect 2440 1676 2442 1693
rect 2576 1676 2578 1693
rect 2728 1676 2730 1693
rect 2888 1676 2890 1693
rect 3048 1676 3050 1693
rect 3216 1676 3218 1693
rect 3368 1676 3370 1693
rect 3464 1677 3466 1693
rect 3462 1676 3468 1677
rect 1806 1672 1807 1676
rect 1811 1672 1812 1676
rect 1806 1671 1812 1672
rect 1830 1675 1836 1676
rect 1830 1671 1831 1675
rect 1835 1671 1836 1675
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 135 1670 139 1671
rect 135 1665 139 1666
rect 191 1670 195 1671
rect 191 1665 195 1666
rect 247 1670 251 1671
rect 247 1665 251 1666
rect 295 1670 299 1671
rect 295 1665 299 1666
rect 399 1670 403 1671
rect 399 1665 403 1666
rect 407 1670 411 1671
rect 407 1665 411 1666
rect 535 1670 539 1671
rect 535 1665 539 1666
rect 567 1670 571 1671
rect 567 1665 571 1666
rect 687 1670 691 1671
rect 687 1665 691 1666
rect 751 1670 755 1671
rect 751 1665 755 1666
rect 855 1670 859 1671
rect 855 1665 859 1666
rect 935 1670 939 1671
rect 935 1665 939 1666
rect 1039 1670 1043 1671
rect 1039 1665 1043 1666
rect 1119 1670 1123 1671
rect 1119 1665 1123 1666
rect 1231 1670 1235 1671
rect 1231 1665 1235 1666
rect 1311 1670 1315 1671
rect 1311 1665 1315 1666
rect 1431 1670 1435 1671
rect 1431 1665 1435 1666
rect 1503 1670 1507 1671
rect 1503 1665 1507 1666
rect 1639 1670 1643 1671
rect 1639 1665 1643 1666
rect 1671 1670 1675 1671
rect 1671 1665 1675 1666
rect 1767 1670 1771 1671
rect 1830 1670 1836 1671
rect 1934 1675 1940 1676
rect 1934 1671 1935 1675
rect 1939 1671 1940 1675
rect 1934 1670 1940 1671
rect 2062 1675 2068 1676
rect 2062 1671 2063 1675
rect 2067 1671 2068 1675
rect 2062 1670 2068 1671
rect 2182 1675 2188 1676
rect 2182 1671 2183 1675
rect 2187 1671 2188 1675
rect 2182 1670 2188 1671
rect 2310 1675 2316 1676
rect 2310 1671 2311 1675
rect 2315 1671 2316 1675
rect 2310 1670 2316 1671
rect 2438 1675 2444 1676
rect 2438 1671 2439 1675
rect 2443 1671 2444 1675
rect 2438 1670 2444 1671
rect 2574 1675 2580 1676
rect 2574 1671 2575 1675
rect 2579 1671 2580 1675
rect 2574 1670 2580 1671
rect 2726 1675 2732 1676
rect 2726 1671 2727 1675
rect 2731 1671 2732 1675
rect 2726 1670 2732 1671
rect 2886 1675 2892 1676
rect 2886 1671 2887 1675
rect 2891 1671 2892 1675
rect 2886 1670 2892 1671
rect 3046 1675 3052 1676
rect 3046 1671 3047 1675
rect 3051 1671 3052 1675
rect 3046 1670 3052 1671
rect 3214 1675 3220 1676
rect 3214 1671 3215 1675
rect 3219 1671 3220 1675
rect 3214 1670 3220 1671
rect 3366 1675 3372 1676
rect 3366 1671 3367 1675
rect 3371 1671 3372 1675
rect 3462 1672 3463 1676
rect 3467 1672 3468 1676
rect 3462 1671 3468 1672
rect 3366 1670 3372 1671
rect 1767 1665 1771 1666
rect 112 1649 114 1665
rect 110 1648 116 1649
rect 192 1648 194 1665
rect 296 1648 298 1665
rect 408 1648 410 1665
rect 536 1648 538 1665
rect 688 1648 690 1665
rect 856 1648 858 1665
rect 1040 1648 1042 1665
rect 1232 1648 1234 1665
rect 1432 1648 1434 1665
rect 1640 1648 1642 1665
rect 1768 1649 1770 1665
rect 1806 1659 1812 1660
rect 1806 1655 1807 1659
rect 1811 1655 1812 1659
rect 3462 1659 3468 1660
rect 1806 1654 1812 1655
rect 1830 1656 1836 1657
rect 1766 1648 1772 1649
rect 110 1644 111 1648
rect 115 1644 116 1648
rect 110 1643 116 1644
rect 190 1647 196 1648
rect 190 1643 191 1647
rect 195 1643 196 1647
rect 190 1642 196 1643
rect 294 1647 300 1648
rect 294 1643 295 1647
rect 299 1643 300 1647
rect 294 1642 300 1643
rect 406 1647 412 1648
rect 406 1643 407 1647
rect 411 1643 412 1647
rect 406 1642 412 1643
rect 534 1647 540 1648
rect 534 1643 535 1647
rect 539 1643 540 1647
rect 534 1642 540 1643
rect 686 1647 692 1648
rect 686 1643 687 1647
rect 691 1643 692 1647
rect 686 1642 692 1643
rect 854 1647 860 1648
rect 854 1643 855 1647
rect 859 1643 860 1647
rect 854 1642 860 1643
rect 1038 1647 1044 1648
rect 1038 1643 1039 1647
rect 1043 1643 1044 1647
rect 1038 1642 1044 1643
rect 1230 1647 1236 1648
rect 1230 1643 1231 1647
rect 1235 1643 1236 1647
rect 1230 1642 1236 1643
rect 1430 1647 1436 1648
rect 1430 1643 1431 1647
rect 1435 1643 1436 1647
rect 1430 1642 1436 1643
rect 1638 1647 1644 1648
rect 1638 1643 1639 1647
rect 1643 1643 1644 1647
rect 1766 1644 1767 1648
rect 1771 1644 1772 1648
rect 1766 1643 1772 1644
rect 1638 1642 1644 1643
rect 110 1631 116 1632
rect 110 1627 111 1631
rect 115 1627 116 1631
rect 1766 1631 1772 1632
rect 110 1626 116 1627
rect 190 1628 196 1629
rect 112 1603 114 1626
rect 190 1624 191 1628
rect 195 1624 196 1628
rect 190 1623 196 1624
rect 294 1628 300 1629
rect 294 1624 295 1628
rect 299 1624 300 1628
rect 294 1623 300 1624
rect 406 1628 412 1629
rect 406 1624 407 1628
rect 411 1624 412 1628
rect 406 1623 412 1624
rect 534 1628 540 1629
rect 534 1624 535 1628
rect 539 1624 540 1628
rect 534 1623 540 1624
rect 686 1628 692 1629
rect 686 1624 687 1628
rect 691 1624 692 1628
rect 686 1623 692 1624
rect 854 1628 860 1629
rect 854 1624 855 1628
rect 859 1624 860 1628
rect 854 1623 860 1624
rect 1038 1628 1044 1629
rect 1038 1624 1039 1628
rect 1043 1624 1044 1628
rect 1038 1623 1044 1624
rect 1230 1628 1236 1629
rect 1230 1624 1231 1628
rect 1235 1624 1236 1628
rect 1230 1623 1236 1624
rect 1430 1628 1436 1629
rect 1430 1624 1431 1628
rect 1435 1624 1436 1628
rect 1430 1623 1436 1624
rect 1638 1628 1644 1629
rect 1638 1624 1639 1628
rect 1643 1624 1644 1628
rect 1766 1627 1767 1631
rect 1771 1627 1772 1631
rect 1808 1627 1810 1654
rect 1830 1652 1831 1656
rect 1835 1652 1836 1656
rect 1830 1651 1836 1652
rect 1934 1656 1940 1657
rect 1934 1652 1935 1656
rect 1939 1652 1940 1656
rect 1934 1651 1940 1652
rect 2062 1656 2068 1657
rect 2062 1652 2063 1656
rect 2067 1652 2068 1656
rect 2062 1651 2068 1652
rect 2182 1656 2188 1657
rect 2182 1652 2183 1656
rect 2187 1652 2188 1656
rect 2182 1651 2188 1652
rect 2310 1656 2316 1657
rect 2310 1652 2311 1656
rect 2315 1652 2316 1656
rect 2310 1651 2316 1652
rect 2438 1656 2444 1657
rect 2438 1652 2439 1656
rect 2443 1652 2444 1656
rect 2438 1651 2444 1652
rect 2574 1656 2580 1657
rect 2574 1652 2575 1656
rect 2579 1652 2580 1656
rect 2574 1651 2580 1652
rect 2726 1656 2732 1657
rect 2726 1652 2727 1656
rect 2731 1652 2732 1656
rect 2726 1651 2732 1652
rect 2886 1656 2892 1657
rect 2886 1652 2887 1656
rect 2891 1652 2892 1656
rect 2886 1651 2892 1652
rect 3046 1656 3052 1657
rect 3046 1652 3047 1656
rect 3051 1652 3052 1656
rect 3046 1651 3052 1652
rect 3214 1656 3220 1657
rect 3214 1652 3215 1656
rect 3219 1652 3220 1656
rect 3214 1651 3220 1652
rect 3366 1656 3372 1657
rect 3366 1652 3367 1656
rect 3371 1652 3372 1656
rect 3462 1655 3463 1659
rect 3467 1655 3468 1659
rect 3462 1654 3468 1655
rect 3366 1651 3372 1652
rect 1832 1627 1834 1651
rect 1936 1627 1938 1651
rect 2064 1627 2066 1651
rect 2184 1627 2186 1651
rect 2312 1627 2314 1651
rect 2440 1627 2442 1651
rect 2576 1627 2578 1651
rect 2728 1627 2730 1651
rect 2888 1627 2890 1651
rect 3048 1627 3050 1651
rect 3216 1627 3218 1651
rect 3368 1627 3370 1651
rect 3464 1627 3466 1654
rect 1766 1626 1772 1627
rect 1807 1626 1811 1627
rect 1638 1623 1644 1624
rect 192 1603 194 1623
rect 296 1603 298 1623
rect 408 1603 410 1623
rect 536 1603 538 1623
rect 688 1603 690 1623
rect 856 1603 858 1623
rect 1040 1603 1042 1623
rect 1232 1603 1234 1623
rect 1432 1603 1434 1623
rect 1640 1603 1642 1623
rect 1768 1603 1770 1626
rect 1807 1621 1811 1622
rect 1831 1626 1835 1627
rect 1831 1621 1835 1622
rect 1935 1626 1939 1627
rect 1935 1621 1939 1622
rect 1943 1626 1947 1627
rect 1943 1621 1947 1622
rect 2063 1626 2067 1627
rect 2063 1621 2067 1622
rect 2087 1626 2091 1627
rect 2087 1621 2091 1622
rect 2183 1626 2187 1627
rect 2183 1621 2187 1622
rect 2231 1626 2235 1627
rect 2231 1621 2235 1622
rect 2311 1626 2315 1627
rect 2311 1621 2315 1622
rect 2367 1626 2371 1627
rect 2367 1621 2371 1622
rect 2439 1626 2443 1627
rect 2439 1621 2443 1622
rect 2503 1626 2507 1627
rect 2503 1621 2507 1622
rect 2575 1626 2579 1627
rect 2575 1621 2579 1622
rect 2639 1626 2643 1627
rect 2639 1621 2643 1622
rect 2727 1626 2731 1627
rect 2727 1621 2731 1622
rect 2767 1626 2771 1627
rect 2767 1621 2771 1622
rect 2887 1626 2891 1627
rect 2887 1621 2891 1622
rect 2895 1626 2899 1627
rect 2895 1621 2899 1622
rect 3015 1626 3019 1627
rect 3015 1621 3019 1622
rect 3047 1626 3051 1627
rect 3047 1621 3051 1622
rect 3135 1626 3139 1627
rect 3135 1621 3139 1622
rect 3215 1626 3219 1627
rect 3215 1621 3219 1622
rect 3263 1626 3267 1627
rect 3263 1621 3267 1622
rect 3367 1626 3371 1627
rect 3367 1621 3371 1622
rect 3463 1626 3467 1627
rect 3463 1621 3467 1622
rect 111 1602 115 1603
rect 111 1597 115 1598
rect 191 1602 195 1603
rect 191 1597 195 1598
rect 295 1602 299 1603
rect 295 1597 299 1598
rect 327 1602 331 1603
rect 327 1597 331 1598
rect 407 1602 411 1603
rect 407 1597 411 1598
rect 431 1602 435 1603
rect 431 1597 435 1598
rect 535 1602 539 1603
rect 535 1597 539 1598
rect 543 1602 547 1603
rect 543 1597 547 1598
rect 671 1602 675 1603
rect 671 1597 675 1598
rect 687 1602 691 1603
rect 687 1597 691 1598
rect 815 1602 819 1603
rect 815 1597 819 1598
rect 855 1602 859 1603
rect 855 1597 859 1598
rect 967 1602 971 1603
rect 967 1597 971 1598
rect 1039 1602 1043 1603
rect 1039 1597 1043 1598
rect 1119 1602 1123 1603
rect 1119 1597 1123 1598
rect 1231 1602 1235 1603
rect 1231 1597 1235 1598
rect 1279 1602 1283 1603
rect 1279 1597 1283 1598
rect 1431 1602 1435 1603
rect 1431 1597 1435 1598
rect 1439 1602 1443 1603
rect 1439 1597 1443 1598
rect 1607 1602 1611 1603
rect 1607 1597 1611 1598
rect 1639 1602 1643 1603
rect 1639 1597 1643 1598
rect 1767 1602 1771 1603
rect 1808 1602 1810 1621
rect 1832 1605 1834 1621
rect 1944 1605 1946 1621
rect 2088 1605 2090 1621
rect 2232 1605 2234 1621
rect 2368 1605 2370 1621
rect 2504 1605 2506 1621
rect 2640 1605 2642 1621
rect 2768 1605 2770 1621
rect 2896 1605 2898 1621
rect 3016 1605 3018 1621
rect 3136 1605 3138 1621
rect 3264 1605 3266 1621
rect 3368 1605 3370 1621
rect 1830 1604 1836 1605
rect 1767 1597 1771 1598
rect 1806 1601 1812 1602
rect 1806 1597 1807 1601
rect 1811 1597 1812 1601
rect 1830 1600 1831 1604
rect 1835 1600 1836 1604
rect 1830 1599 1836 1600
rect 1942 1604 1948 1605
rect 1942 1600 1943 1604
rect 1947 1600 1948 1604
rect 1942 1599 1948 1600
rect 2086 1604 2092 1605
rect 2086 1600 2087 1604
rect 2091 1600 2092 1604
rect 2086 1599 2092 1600
rect 2230 1604 2236 1605
rect 2230 1600 2231 1604
rect 2235 1600 2236 1604
rect 2230 1599 2236 1600
rect 2366 1604 2372 1605
rect 2366 1600 2367 1604
rect 2371 1600 2372 1604
rect 2366 1599 2372 1600
rect 2502 1604 2508 1605
rect 2502 1600 2503 1604
rect 2507 1600 2508 1604
rect 2502 1599 2508 1600
rect 2638 1604 2644 1605
rect 2638 1600 2639 1604
rect 2643 1600 2644 1604
rect 2638 1599 2644 1600
rect 2766 1604 2772 1605
rect 2766 1600 2767 1604
rect 2771 1600 2772 1604
rect 2766 1599 2772 1600
rect 2894 1604 2900 1605
rect 2894 1600 2895 1604
rect 2899 1600 2900 1604
rect 2894 1599 2900 1600
rect 3014 1604 3020 1605
rect 3014 1600 3015 1604
rect 3019 1600 3020 1604
rect 3014 1599 3020 1600
rect 3134 1604 3140 1605
rect 3134 1600 3135 1604
rect 3139 1600 3140 1604
rect 3134 1599 3140 1600
rect 3262 1604 3268 1605
rect 3262 1600 3263 1604
rect 3267 1600 3268 1604
rect 3262 1599 3268 1600
rect 3366 1604 3372 1605
rect 3366 1600 3367 1604
rect 3371 1600 3372 1604
rect 3464 1602 3466 1621
rect 3366 1599 3372 1600
rect 3462 1601 3468 1602
rect 112 1578 114 1597
rect 328 1581 330 1597
rect 432 1581 434 1597
rect 544 1581 546 1597
rect 672 1581 674 1597
rect 816 1581 818 1597
rect 968 1581 970 1597
rect 1120 1581 1122 1597
rect 1280 1581 1282 1597
rect 1440 1581 1442 1597
rect 1608 1581 1610 1597
rect 326 1580 332 1581
rect 110 1577 116 1578
rect 110 1573 111 1577
rect 115 1573 116 1577
rect 326 1576 327 1580
rect 331 1576 332 1580
rect 326 1575 332 1576
rect 430 1580 436 1581
rect 430 1576 431 1580
rect 435 1576 436 1580
rect 430 1575 436 1576
rect 542 1580 548 1581
rect 542 1576 543 1580
rect 547 1576 548 1580
rect 542 1575 548 1576
rect 670 1580 676 1581
rect 670 1576 671 1580
rect 675 1576 676 1580
rect 670 1575 676 1576
rect 814 1580 820 1581
rect 814 1576 815 1580
rect 819 1576 820 1580
rect 814 1575 820 1576
rect 966 1580 972 1581
rect 966 1576 967 1580
rect 971 1576 972 1580
rect 966 1575 972 1576
rect 1118 1580 1124 1581
rect 1118 1576 1119 1580
rect 1123 1576 1124 1580
rect 1118 1575 1124 1576
rect 1278 1580 1284 1581
rect 1278 1576 1279 1580
rect 1283 1576 1284 1580
rect 1278 1575 1284 1576
rect 1438 1580 1444 1581
rect 1438 1576 1439 1580
rect 1443 1576 1444 1580
rect 1438 1575 1444 1576
rect 1606 1580 1612 1581
rect 1606 1576 1607 1580
rect 1611 1576 1612 1580
rect 1768 1578 1770 1597
rect 1806 1596 1812 1597
rect 3462 1597 3463 1601
rect 3467 1597 3468 1601
rect 3462 1596 3468 1597
rect 1830 1585 1836 1586
rect 1806 1584 1812 1585
rect 1806 1580 1807 1584
rect 1811 1580 1812 1584
rect 1830 1581 1831 1585
rect 1835 1581 1836 1585
rect 1830 1580 1836 1581
rect 1942 1585 1948 1586
rect 1942 1581 1943 1585
rect 1947 1581 1948 1585
rect 1942 1580 1948 1581
rect 2086 1585 2092 1586
rect 2086 1581 2087 1585
rect 2091 1581 2092 1585
rect 2086 1580 2092 1581
rect 2230 1585 2236 1586
rect 2230 1581 2231 1585
rect 2235 1581 2236 1585
rect 2230 1580 2236 1581
rect 2366 1585 2372 1586
rect 2366 1581 2367 1585
rect 2371 1581 2372 1585
rect 2366 1580 2372 1581
rect 2502 1585 2508 1586
rect 2502 1581 2503 1585
rect 2507 1581 2508 1585
rect 2502 1580 2508 1581
rect 2638 1585 2644 1586
rect 2638 1581 2639 1585
rect 2643 1581 2644 1585
rect 2638 1580 2644 1581
rect 2766 1585 2772 1586
rect 2766 1581 2767 1585
rect 2771 1581 2772 1585
rect 2766 1580 2772 1581
rect 2894 1585 2900 1586
rect 2894 1581 2895 1585
rect 2899 1581 2900 1585
rect 2894 1580 2900 1581
rect 3014 1585 3020 1586
rect 3014 1581 3015 1585
rect 3019 1581 3020 1585
rect 3014 1580 3020 1581
rect 3134 1585 3140 1586
rect 3134 1581 3135 1585
rect 3139 1581 3140 1585
rect 3134 1580 3140 1581
rect 3262 1585 3268 1586
rect 3262 1581 3263 1585
rect 3267 1581 3268 1585
rect 3262 1580 3268 1581
rect 3366 1585 3372 1586
rect 3366 1581 3367 1585
rect 3371 1581 3372 1585
rect 3366 1580 3372 1581
rect 3462 1584 3468 1585
rect 3462 1580 3463 1584
rect 3467 1580 3468 1584
rect 1806 1579 1812 1580
rect 1606 1575 1612 1576
rect 1766 1577 1772 1578
rect 110 1572 116 1573
rect 1766 1573 1767 1577
rect 1771 1573 1772 1577
rect 1766 1572 1772 1573
rect 326 1561 332 1562
rect 110 1560 116 1561
rect 110 1556 111 1560
rect 115 1556 116 1560
rect 326 1557 327 1561
rect 331 1557 332 1561
rect 326 1556 332 1557
rect 430 1561 436 1562
rect 430 1557 431 1561
rect 435 1557 436 1561
rect 430 1556 436 1557
rect 542 1561 548 1562
rect 542 1557 543 1561
rect 547 1557 548 1561
rect 542 1556 548 1557
rect 670 1561 676 1562
rect 670 1557 671 1561
rect 675 1557 676 1561
rect 670 1556 676 1557
rect 814 1561 820 1562
rect 814 1557 815 1561
rect 819 1557 820 1561
rect 814 1556 820 1557
rect 966 1561 972 1562
rect 966 1557 967 1561
rect 971 1557 972 1561
rect 966 1556 972 1557
rect 1118 1561 1124 1562
rect 1118 1557 1119 1561
rect 1123 1557 1124 1561
rect 1118 1556 1124 1557
rect 1278 1561 1284 1562
rect 1278 1557 1279 1561
rect 1283 1557 1284 1561
rect 1278 1556 1284 1557
rect 1438 1561 1444 1562
rect 1438 1557 1439 1561
rect 1443 1557 1444 1561
rect 1438 1556 1444 1557
rect 1606 1561 1612 1562
rect 1606 1557 1607 1561
rect 1611 1557 1612 1561
rect 1606 1556 1612 1557
rect 1766 1560 1772 1561
rect 1766 1556 1767 1560
rect 1771 1556 1772 1560
rect 110 1555 116 1556
rect 112 1535 114 1555
rect 328 1535 330 1556
rect 432 1535 434 1556
rect 544 1535 546 1556
rect 672 1535 674 1556
rect 816 1535 818 1556
rect 968 1535 970 1556
rect 1120 1535 1122 1556
rect 1280 1535 1282 1556
rect 1440 1535 1442 1556
rect 1608 1535 1610 1556
rect 1766 1555 1772 1556
rect 1808 1555 1810 1579
rect 1832 1555 1834 1580
rect 1944 1555 1946 1580
rect 2088 1555 2090 1580
rect 2232 1555 2234 1580
rect 2368 1555 2370 1580
rect 2504 1555 2506 1580
rect 2640 1555 2642 1580
rect 2768 1555 2770 1580
rect 2896 1555 2898 1580
rect 3016 1555 3018 1580
rect 3136 1555 3138 1580
rect 3264 1555 3266 1580
rect 3368 1555 3370 1580
rect 3462 1579 3468 1580
rect 3464 1555 3466 1579
rect 1768 1535 1770 1555
rect 1807 1554 1811 1555
rect 1807 1549 1811 1550
rect 1831 1554 1835 1555
rect 1831 1549 1835 1550
rect 1839 1554 1843 1555
rect 1839 1549 1843 1550
rect 1943 1554 1947 1555
rect 1943 1549 1947 1550
rect 1991 1554 1995 1555
rect 1991 1549 1995 1550
rect 2087 1554 2091 1555
rect 2087 1549 2091 1550
rect 2151 1554 2155 1555
rect 2151 1549 2155 1550
rect 2231 1554 2235 1555
rect 2231 1549 2235 1550
rect 2303 1554 2307 1555
rect 2303 1549 2307 1550
rect 2367 1554 2371 1555
rect 2367 1549 2371 1550
rect 2455 1554 2459 1555
rect 2455 1549 2459 1550
rect 2503 1554 2507 1555
rect 2503 1549 2507 1550
rect 2599 1554 2603 1555
rect 2599 1549 2603 1550
rect 2639 1554 2643 1555
rect 2639 1549 2643 1550
rect 2735 1554 2739 1555
rect 2735 1549 2739 1550
rect 2767 1554 2771 1555
rect 2767 1549 2771 1550
rect 2871 1554 2875 1555
rect 2871 1549 2875 1550
rect 2895 1554 2899 1555
rect 2895 1549 2899 1550
rect 3007 1554 3011 1555
rect 3007 1549 3011 1550
rect 3015 1554 3019 1555
rect 3015 1549 3019 1550
rect 3135 1554 3139 1555
rect 3135 1549 3139 1550
rect 3143 1554 3147 1555
rect 3143 1549 3147 1550
rect 3263 1554 3267 1555
rect 3263 1549 3267 1550
rect 3367 1554 3371 1555
rect 3367 1549 3371 1550
rect 3463 1554 3467 1555
rect 3463 1549 3467 1550
rect 111 1534 115 1535
rect 111 1529 115 1530
rect 223 1534 227 1535
rect 223 1529 227 1530
rect 327 1534 331 1535
rect 327 1529 331 1530
rect 343 1534 347 1535
rect 343 1529 347 1530
rect 431 1534 435 1535
rect 431 1529 435 1530
rect 471 1534 475 1535
rect 471 1529 475 1530
rect 543 1534 547 1535
rect 543 1529 547 1530
rect 607 1534 611 1535
rect 607 1529 611 1530
rect 671 1534 675 1535
rect 671 1529 675 1530
rect 751 1534 755 1535
rect 751 1529 755 1530
rect 815 1534 819 1535
rect 815 1529 819 1530
rect 895 1534 899 1535
rect 895 1529 899 1530
rect 967 1534 971 1535
rect 967 1529 971 1530
rect 1047 1534 1051 1535
rect 1047 1529 1051 1530
rect 1119 1534 1123 1535
rect 1119 1529 1123 1530
rect 1199 1534 1203 1535
rect 1199 1529 1203 1530
rect 1279 1534 1283 1535
rect 1279 1529 1283 1530
rect 1351 1534 1355 1535
rect 1351 1529 1355 1530
rect 1439 1534 1443 1535
rect 1439 1529 1443 1530
rect 1503 1534 1507 1535
rect 1503 1529 1507 1530
rect 1607 1534 1611 1535
rect 1607 1529 1611 1530
rect 1767 1534 1771 1535
rect 1808 1533 1810 1549
rect 1767 1529 1771 1530
rect 1806 1532 1812 1533
rect 1840 1532 1842 1549
rect 1992 1532 1994 1549
rect 2152 1532 2154 1549
rect 2304 1532 2306 1549
rect 2456 1532 2458 1549
rect 2600 1532 2602 1549
rect 2736 1532 2738 1549
rect 2872 1532 2874 1549
rect 3008 1532 3010 1549
rect 3144 1532 3146 1549
rect 3464 1533 3466 1549
rect 3462 1532 3468 1533
rect 112 1513 114 1529
rect 110 1512 116 1513
rect 224 1512 226 1529
rect 344 1512 346 1529
rect 472 1512 474 1529
rect 608 1512 610 1529
rect 752 1512 754 1529
rect 896 1512 898 1529
rect 1048 1512 1050 1529
rect 1200 1512 1202 1529
rect 1352 1512 1354 1529
rect 1504 1512 1506 1529
rect 1768 1513 1770 1529
rect 1806 1528 1807 1532
rect 1811 1528 1812 1532
rect 1806 1527 1812 1528
rect 1838 1531 1844 1532
rect 1838 1527 1839 1531
rect 1843 1527 1844 1531
rect 1838 1526 1844 1527
rect 1990 1531 1996 1532
rect 1990 1527 1991 1531
rect 1995 1527 1996 1531
rect 1990 1526 1996 1527
rect 2150 1531 2156 1532
rect 2150 1527 2151 1531
rect 2155 1527 2156 1531
rect 2150 1526 2156 1527
rect 2302 1531 2308 1532
rect 2302 1527 2303 1531
rect 2307 1527 2308 1531
rect 2302 1526 2308 1527
rect 2454 1531 2460 1532
rect 2454 1527 2455 1531
rect 2459 1527 2460 1531
rect 2454 1526 2460 1527
rect 2598 1531 2604 1532
rect 2598 1527 2599 1531
rect 2603 1527 2604 1531
rect 2598 1526 2604 1527
rect 2734 1531 2740 1532
rect 2734 1527 2735 1531
rect 2739 1527 2740 1531
rect 2734 1526 2740 1527
rect 2870 1531 2876 1532
rect 2870 1527 2871 1531
rect 2875 1527 2876 1531
rect 2870 1526 2876 1527
rect 3006 1531 3012 1532
rect 3006 1527 3007 1531
rect 3011 1527 3012 1531
rect 3006 1526 3012 1527
rect 3142 1531 3148 1532
rect 3142 1527 3143 1531
rect 3147 1527 3148 1531
rect 3462 1528 3463 1532
rect 3467 1528 3468 1532
rect 3462 1527 3468 1528
rect 3142 1526 3148 1527
rect 1806 1515 1812 1516
rect 1766 1512 1772 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 222 1511 228 1512
rect 222 1507 223 1511
rect 227 1507 228 1511
rect 222 1506 228 1507
rect 342 1511 348 1512
rect 342 1507 343 1511
rect 347 1507 348 1511
rect 342 1506 348 1507
rect 470 1511 476 1512
rect 470 1507 471 1511
rect 475 1507 476 1511
rect 470 1506 476 1507
rect 606 1511 612 1512
rect 606 1507 607 1511
rect 611 1507 612 1511
rect 606 1506 612 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 894 1511 900 1512
rect 894 1507 895 1511
rect 899 1507 900 1511
rect 894 1506 900 1507
rect 1046 1511 1052 1512
rect 1046 1507 1047 1511
rect 1051 1507 1052 1511
rect 1046 1506 1052 1507
rect 1198 1511 1204 1512
rect 1198 1507 1199 1511
rect 1203 1507 1204 1511
rect 1198 1506 1204 1507
rect 1350 1511 1356 1512
rect 1350 1507 1351 1511
rect 1355 1507 1356 1511
rect 1350 1506 1356 1507
rect 1502 1511 1508 1512
rect 1502 1507 1503 1511
rect 1507 1507 1508 1511
rect 1766 1508 1767 1512
rect 1771 1508 1772 1512
rect 1806 1511 1807 1515
rect 1811 1511 1812 1515
rect 3462 1515 3468 1516
rect 1806 1510 1812 1511
rect 1838 1512 1844 1513
rect 1766 1507 1772 1508
rect 1502 1506 1508 1507
rect 110 1495 116 1496
rect 110 1491 111 1495
rect 115 1491 116 1495
rect 1766 1495 1772 1496
rect 110 1490 116 1491
rect 222 1492 228 1493
rect 112 1463 114 1490
rect 222 1488 223 1492
rect 227 1488 228 1492
rect 222 1487 228 1488
rect 342 1492 348 1493
rect 342 1488 343 1492
rect 347 1488 348 1492
rect 342 1487 348 1488
rect 470 1492 476 1493
rect 470 1488 471 1492
rect 475 1488 476 1492
rect 470 1487 476 1488
rect 606 1492 612 1493
rect 606 1488 607 1492
rect 611 1488 612 1492
rect 606 1487 612 1488
rect 750 1492 756 1493
rect 750 1488 751 1492
rect 755 1488 756 1492
rect 750 1487 756 1488
rect 894 1492 900 1493
rect 894 1488 895 1492
rect 899 1488 900 1492
rect 894 1487 900 1488
rect 1046 1492 1052 1493
rect 1046 1488 1047 1492
rect 1051 1488 1052 1492
rect 1046 1487 1052 1488
rect 1198 1492 1204 1493
rect 1198 1488 1199 1492
rect 1203 1488 1204 1492
rect 1198 1487 1204 1488
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1502 1492 1508 1493
rect 1502 1488 1503 1492
rect 1507 1488 1508 1492
rect 1766 1491 1767 1495
rect 1771 1491 1772 1495
rect 1766 1490 1772 1491
rect 1502 1487 1508 1488
rect 224 1463 226 1487
rect 344 1463 346 1487
rect 472 1463 474 1487
rect 608 1463 610 1487
rect 752 1463 754 1487
rect 896 1463 898 1487
rect 1048 1463 1050 1487
rect 1200 1463 1202 1487
rect 1352 1463 1354 1487
rect 1504 1463 1506 1487
rect 1768 1463 1770 1490
rect 1808 1483 1810 1510
rect 1838 1508 1839 1512
rect 1843 1508 1844 1512
rect 1838 1507 1844 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2150 1512 2156 1513
rect 2150 1508 2151 1512
rect 2155 1508 2156 1512
rect 2150 1507 2156 1508
rect 2302 1512 2308 1513
rect 2302 1508 2303 1512
rect 2307 1508 2308 1512
rect 2302 1507 2308 1508
rect 2454 1512 2460 1513
rect 2454 1508 2455 1512
rect 2459 1508 2460 1512
rect 2454 1507 2460 1508
rect 2598 1512 2604 1513
rect 2598 1508 2599 1512
rect 2603 1508 2604 1512
rect 2598 1507 2604 1508
rect 2734 1512 2740 1513
rect 2734 1508 2735 1512
rect 2739 1508 2740 1512
rect 2734 1507 2740 1508
rect 2870 1512 2876 1513
rect 2870 1508 2871 1512
rect 2875 1508 2876 1512
rect 2870 1507 2876 1508
rect 3006 1512 3012 1513
rect 3006 1508 3007 1512
rect 3011 1508 3012 1512
rect 3006 1507 3012 1508
rect 3142 1512 3148 1513
rect 3142 1508 3143 1512
rect 3147 1508 3148 1512
rect 3462 1511 3463 1515
rect 3467 1511 3468 1515
rect 3462 1510 3468 1511
rect 3142 1507 3148 1508
rect 1840 1483 1842 1507
rect 1992 1483 1994 1507
rect 2152 1483 2154 1507
rect 2304 1483 2306 1507
rect 2456 1483 2458 1507
rect 2600 1483 2602 1507
rect 2736 1483 2738 1507
rect 2872 1483 2874 1507
rect 3008 1483 3010 1507
rect 3144 1483 3146 1507
rect 3464 1483 3466 1510
rect 1807 1482 1811 1483
rect 1807 1477 1811 1478
rect 1839 1482 1843 1483
rect 1839 1477 1843 1478
rect 1943 1482 1947 1483
rect 1943 1477 1947 1478
rect 1991 1482 1995 1483
rect 1991 1477 1995 1478
rect 2055 1482 2059 1483
rect 2055 1477 2059 1478
rect 2151 1482 2155 1483
rect 2151 1477 2155 1478
rect 2191 1482 2195 1483
rect 2191 1477 2195 1478
rect 2303 1482 2307 1483
rect 2303 1477 2307 1478
rect 2335 1482 2339 1483
rect 2335 1477 2339 1478
rect 2455 1482 2459 1483
rect 2455 1477 2459 1478
rect 2479 1482 2483 1483
rect 2479 1477 2483 1478
rect 2599 1482 2603 1483
rect 2599 1477 2603 1478
rect 2631 1482 2635 1483
rect 2631 1477 2635 1478
rect 2735 1482 2739 1483
rect 2735 1477 2739 1478
rect 2783 1482 2787 1483
rect 2783 1477 2787 1478
rect 2871 1482 2875 1483
rect 2871 1477 2875 1478
rect 2935 1482 2939 1483
rect 2935 1477 2939 1478
rect 3007 1482 3011 1483
rect 3007 1477 3011 1478
rect 3087 1482 3091 1483
rect 3087 1477 3091 1478
rect 3143 1482 3147 1483
rect 3143 1477 3147 1478
rect 3239 1482 3243 1483
rect 3239 1477 3243 1478
rect 3463 1482 3467 1483
rect 3463 1477 3467 1478
rect 111 1462 115 1463
rect 111 1457 115 1458
rect 135 1462 139 1463
rect 135 1457 139 1458
rect 223 1462 227 1463
rect 223 1457 227 1458
rect 303 1462 307 1463
rect 303 1457 307 1458
rect 343 1462 347 1463
rect 343 1457 347 1458
rect 471 1462 475 1463
rect 471 1457 475 1458
rect 607 1462 611 1463
rect 607 1457 611 1458
rect 631 1462 635 1463
rect 631 1457 635 1458
rect 751 1462 755 1463
rect 751 1457 755 1458
rect 783 1462 787 1463
rect 783 1457 787 1458
rect 895 1462 899 1463
rect 895 1457 899 1458
rect 927 1462 931 1463
rect 927 1457 931 1458
rect 1047 1462 1051 1463
rect 1047 1457 1051 1458
rect 1063 1462 1067 1463
rect 1063 1457 1067 1458
rect 1199 1462 1203 1463
rect 1199 1457 1203 1458
rect 1335 1462 1339 1463
rect 1335 1457 1339 1458
rect 1351 1462 1355 1463
rect 1351 1457 1355 1458
rect 1471 1462 1475 1463
rect 1471 1457 1475 1458
rect 1503 1462 1507 1463
rect 1503 1457 1507 1458
rect 1767 1462 1771 1463
rect 1808 1458 1810 1477
rect 1944 1461 1946 1477
rect 2056 1461 2058 1477
rect 2192 1461 2194 1477
rect 2336 1461 2338 1477
rect 2480 1461 2482 1477
rect 2632 1461 2634 1477
rect 2784 1461 2786 1477
rect 2936 1461 2938 1477
rect 3088 1461 3090 1477
rect 3240 1461 3242 1477
rect 1942 1460 1948 1461
rect 1767 1457 1771 1458
rect 1806 1457 1812 1458
rect 112 1438 114 1457
rect 136 1441 138 1457
rect 304 1441 306 1457
rect 472 1441 474 1457
rect 632 1441 634 1457
rect 784 1441 786 1457
rect 928 1441 930 1457
rect 1064 1441 1066 1457
rect 1200 1441 1202 1457
rect 1336 1441 1338 1457
rect 1472 1441 1474 1457
rect 134 1440 140 1441
rect 110 1437 116 1438
rect 110 1433 111 1437
rect 115 1433 116 1437
rect 134 1436 135 1440
rect 139 1436 140 1440
rect 134 1435 140 1436
rect 302 1440 308 1441
rect 302 1436 303 1440
rect 307 1436 308 1440
rect 302 1435 308 1436
rect 470 1440 476 1441
rect 470 1436 471 1440
rect 475 1436 476 1440
rect 470 1435 476 1436
rect 630 1440 636 1441
rect 630 1436 631 1440
rect 635 1436 636 1440
rect 630 1435 636 1436
rect 782 1440 788 1441
rect 782 1436 783 1440
rect 787 1436 788 1440
rect 782 1435 788 1436
rect 926 1440 932 1441
rect 926 1436 927 1440
rect 931 1436 932 1440
rect 926 1435 932 1436
rect 1062 1440 1068 1441
rect 1062 1436 1063 1440
rect 1067 1436 1068 1440
rect 1062 1435 1068 1436
rect 1198 1440 1204 1441
rect 1198 1436 1199 1440
rect 1203 1436 1204 1440
rect 1198 1435 1204 1436
rect 1334 1440 1340 1441
rect 1334 1436 1335 1440
rect 1339 1436 1340 1440
rect 1334 1435 1340 1436
rect 1470 1440 1476 1441
rect 1470 1436 1471 1440
rect 1475 1436 1476 1440
rect 1768 1438 1770 1457
rect 1806 1453 1807 1457
rect 1811 1453 1812 1457
rect 1942 1456 1943 1460
rect 1947 1456 1948 1460
rect 1942 1455 1948 1456
rect 2054 1460 2060 1461
rect 2054 1456 2055 1460
rect 2059 1456 2060 1460
rect 2054 1455 2060 1456
rect 2190 1460 2196 1461
rect 2190 1456 2191 1460
rect 2195 1456 2196 1460
rect 2190 1455 2196 1456
rect 2334 1460 2340 1461
rect 2334 1456 2335 1460
rect 2339 1456 2340 1460
rect 2334 1455 2340 1456
rect 2478 1460 2484 1461
rect 2478 1456 2479 1460
rect 2483 1456 2484 1460
rect 2478 1455 2484 1456
rect 2630 1460 2636 1461
rect 2630 1456 2631 1460
rect 2635 1456 2636 1460
rect 2630 1455 2636 1456
rect 2782 1460 2788 1461
rect 2782 1456 2783 1460
rect 2787 1456 2788 1460
rect 2782 1455 2788 1456
rect 2934 1460 2940 1461
rect 2934 1456 2935 1460
rect 2939 1456 2940 1460
rect 2934 1455 2940 1456
rect 3086 1460 3092 1461
rect 3086 1456 3087 1460
rect 3091 1456 3092 1460
rect 3086 1455 3092 1456
rect 3238 1460 3244 1461
rect 3238 1456 3239 1460
rect 3243 1456 3244 1460
rect 3464 1458 3466 1477
rect 3238 1455 3244 1456
rect 3462 1457 3468 1458
rect 1806 1452 1812 1453
rect 3462 1453 3463 1457
rect 3467 1453 3468 1457
rect 3462 1452 3468 1453
rect 1942 1441 1948 1442
rect 1806 1440 1812 1441
rect 1470 1435 1476 1436
rect 1766 1437 1772 1438
rect 110 1432 116 1433
rect 1766 1433 1767 1437
rect 1771 1433 1772 1437
rect 1806 1436 1807 1440
rect 1811 1436 1812 1440
rect 1942 1437 1943 1441
rect 1947 1437 1948 1441
rect 1942 1436 1948 1437
rect 2054 1441 2060 1442
rect 2054 1437 2055 1441
rect 2059 1437 2060 1441
rect 2054 1436 2060 1437
rect 2190 1441 2196 1442
rect 2190 1437 2191 1441
rect 2195 1437 2196 1441
rect 2190 1436 2196 1437
rect 2334 1441 2340 1442
rect 2334 1437 2335 1441
rect 2339 1437 2340 1441
rect 2334 1436 2340 1437
rect 2478 1441 2484 1442
rect 2478 1437 2479 1441
rect 2483 1437 2484 1441
rect 2478 1436 2484 1437
rect 2630 1441 2636 1442
rect 2630 1437 2631 1441
rect 2635 1437 2636 1441
rect 2630 1436 2636 1437
rect 2782 1441 2788 1442
rect 2782 1437 2783 1441
rect 2787 1437 2788 1441
rect 2782 1436 2788 1437
rect 2934 1441 2940 1442
rect 2934 1437 2935 1441
rect 2939 1437 2940 1441
rect 2934 1436 2940 1437
rect 3086 1441 3092 1442
rect 3086 1437 3087 1441
rect 3091 1437 3092 1441
rect 3086 1436 3092 1437
rect 3238 1441 3244 1442
rect 3238 1437 3239 1441
rect 3243 1437 3244 1441
rect 3238 1436 3244 1437
rect 3462 1440 3468 1441
rect 3462 1436 3463 1440
rect 3467 1436 3468 1440
rect 1806 1435 1812 1436
rect 1766 1432 1772 1433
rect 134 1421 140 1422
rect 110 1420 116 1421
rect 110 1416 111 1420
rect 115 1416 116 1420
rect 134 1417 135 1421
rect 139 1417 140 1421
rect 134 1416 140 1417
rect 302 1421 308 1422
rect 302 1417 303 1421
rect 307 1417 308 1421
rect 302 1416 308 1417
rect 470 1421 476 1422
rect 470 1417 471 1421
rect 475 1417 476 1421
rect 470 1416 476 1417
rect 630 1421 636 1422
rect 630 1417 631 1421
rect 635 1417 636 1421
rect 630 1416 636 1417
rect 782 1421 788 1422
rect 782 1417 783 1421
rect 787 1417 788 1421
rect 782 1416 788 1417
rect 926 1421 932 1422
rect 926 1417 927 1421
rect 931 1417 932 1421
rect 926 1416 932 1417
rect 1062 1421 1068 1422
rect 1062 1417 1063 1421
rect 1067 1417 1068 1421
rect 1062 1416 1068 1417
rect 1198 1421 1204 1422
rect 1198 1417 1199 1421
rect 1203 1417 1204 1421
rect 1198 1416 1204 1417
rect 1334 1421 1340 1422
rect 1334 1417 1335 1421
rect 1339 1417 1340 1421
rect 1334 1416 1340 1417
rect 1470 1421 1476 1422
rect 1470 1417 1471 1421
rect 1475 1417 1476 1421
rect 1470 1416 1476 1417
rect 1766 1420 1772 1421
rect 1766 1416 1767 1420
rect 1771 1416 1772 1420
rect 110 1415 116 1416
rect 112 1395 114 1415
rect 136 1395 138 1416
rect 304 1395 306 1416
rect 472 1395 474 1416
rect 632 1395 634 1416
rect 784 1395 786 1416
rect 928 1395 930 1416
rect 1064 1395 1066 1416
rect 1200 1395 1202 1416
rect 1336 1395 1338 1416
rect 1472 1395 1474 1416
rect 1766 1415 1772 1416
rect 1768 1395 1770 1415
rect 1808 1411 1810 1435
rect 1944 1411 1946 1436
rect 2056 1411 2058 1436
rect 2192 1411 2194 1436
rect 2336 1411 2338 1436
rect 2480 1411 2482 1436
rect 2632 1411 2634 1436
rect 2784 1411 2786 1436
rect 2936 1411 2938 1436
rect 3088 1411 3090 1436
rect 3240 1411 3242 1436
rect 3462 1435 3468 1436
rect 3464 1411 3466 1435
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1943 1410 1947 1411
rect 1943 1405 1947 1406
rect 2055 1410 2059 1411
rect 2055 1405 2059 1406
rect 2095 1410 2099 1411
rect 2095 1405 2099 1406
rect 2191 1410 2195 1411
rect 2191 1405 2195 1406
rect 2199 1410 2203 1411
rect 2199 1405 2203 1406
rect 2319 1410 2323 1411
rect 2319 1405 2323 1406
rect 2335 1410 2339 1411
rect 2335 1405 2339 1406
rect 2455 1410 2459 1411
rect 2455 1405 2459 1406
rect 2479 1410 2483 1411
rect 2479 1405 2483 1406
rect 2599 1410 2603 1411
rect 2599 1405 2603 1406
rect 2631 1410 2635 1411
rect 2631 1405 2635 1406
rect 2743 1410 2747 1411
rect 2743 1405 2747 1406
rect 2783 1410 2787 1411
rect 2783 1405 2787 1406
rect 2887 1410 2891 1411
rect 2887 1405 2891 1406
rect 2935 1410 2939 1411
rect 2935 1405 2939 1406
rect 3031 1410 3035 1411
rect 3031 1405 3035 1406
rect 3087 1410 3091 1411
rect 3087 1405 3091 1406
rect 3175 1410 3179 1411
rect 3175 1405 3179 1406
rect 3239 1410 3243 1411
rect 3239 1405 3243 1406
rect 3327 1410 3331 1411
rect 3327 1405 3331 1406
rect 3463 1410 3467 1411
rect 3463 1405 3467 1406
rect 111 1394 115 1395
rect 111 1389 115 1390
rect 135 1394 139 1395
rect 135 1389 139 1390
rect 279 1394 283 1395
rect 279 1389 283 1390
rect 303 1394 307 1395
rect 303 1389 307 1390
rect 447 1394 451 1395
rect 447 1389 451 1390
rect 471 1394 475 1395
rect 471 1389 475 1390
rect 607 1394 611 1395
rect 607 1389 611 1390
rect 631 1394 635 1395
rect 631 1389 635 1390
rect 759 1394 763 1395
rect 759 1389 763 1390
rect 783 1394 787 1395
rect 783 1389 787 1390
rect 903 1394 907 1395
rect 903 1389 907 1390
rect 927 1394 931 1395
rect 927 1389 931 1390
rect 1031 1394 1035 1395
rect 1031 1389 1035 1390
rect 1063 1394 1067 1395
rect 1063 1389 1067 1390
rect 1159 1394 1163 1395
rect 1159 1389 1163 1390
rect 1199 1394 1203 1395
rect 1199 1389 1203 1390
rect 1287 1394 1291 1395
rect 1287 1389 1291 1390
rect 1335 1394 1339 1395
rect 1335 1389 1339 1390
rect 1415 1394 1419 1395
rect 1415 1389 1419 1390
rect 1471 1394 1475 1395
rect 1471 1389 1475 1390
rect 1767 1394 1771 1395
rect 1767 1389 1771 1390
rect 1808 1389 1810 1405
rect 112 1373 114 1389
rect 110 1372 116 1373
rect 136 1372 138 1389
rect 280 1372 282 1389
rect 448 1372 450 1389
rect 608 1372 610 1389
rect 760 1372 762 1389
rect 904 1372 906 1389
rect 1032 1372 1034 1389
rect 1160 1372 1162 1389
rect 1288 1372 1290 1389
rect 1416 1372 1418 1389
rect 1768 1373 1770 1389
rect 1806 1388 1812 1389
rect 2096 1388 2098 1405
rect 2200 1388 2202 1405
rect 2320 1388 2322 1405
rect 2456 1388 2458 1405
rect 2600 1388 2602 1405
rect 2744 1388 2746 1405
rect 2888 1388 2890 1405
rect 3032 1388 3034 1405
rect 3176 1388 3178 1405
rect 3328 1388 3330 1405
rect 3464 1389 3466 1405
rect 3462 1388 3468 1389
rect 1806 1384 1807 1388
rect 1811 1384 1812 1388
rect 1806 1383 1812 1384
rect 2094 1387 2100 1388
rect 2094 1383 2095 1387
rect 2099 1383 2100 1387
rect 2094 1382 2100 1383
rect 2198 1387 2204 1388
rect 2198 1383 2199 1387
rect 2203 1383 2204 1387
rect 2198 1382 2204 1383
rect 2318 1387 2324 1388
rect 2318 1383 2319 1387
rect 2323 1383 2324 1387
rect 2318 1382 2324 1383
rect 2454 1387 2460 1388
rect 2454 1383 2455 1387
rect 2459 1383 2460 1387
rect 2454 1382 2460 1383
rect 2598 1387 2604 1388
rect 2598 1383 2599 1387
rect 2603 1383 2604 1387
rect 2598 1382 2604 1383
rect 2742 1387 2748 1388
rect 2742 1383 2743 1387
rect 2747 1383 2748 1387
rect 2742 1382 2748 1383
rect 2886 1387 2892 1388
rect 2886 1383 2887 1387
rect 2891 1383 2892 1387
rect 2886 1382 2892 1383
rect 3030 1387 3036 1388
rect 3030 1383 3031 1387
rect 3035 1383 3036 1387
rect 3030 1382 3036 1383
rect 3174 1387 3180 1388
rect 3174 1383 3175 1387
rect 3179 1383 3180 1387
rect 3174 1382 3180 1383
rect 3326 1387 3332 1388
rect 3326 1383 3327 1387
rect 3331 1383 3332 1387
rect 3462 1384 3463 1388
rect 3467 1384 3468 1388
rect 3462 1383 3468 1384
rect 3326 1382 3332 1383
rect 1766 1372 1772 1373
rect 110 1368 111 1372
rect 115 1368 116 1372
rect 110 1367 116 1368
rect 134 1371 140 1372
rect 134 1367 135 1371
rect 139 1367 140 1371
rect 134 1366 140 1367
rect 278 1371 284 1372
rect 278 1367 279 1371
rect 283 1367 284 1371
rect 278 1366 284 1367
rect 446 1371 452 1372
rect 446 1367 447 1371
rect 451 1367 452 1371
rect 446 1366 452 1367
rect 606 1371 612 1372
rect 606 1367 607 1371
rect 611 1367 612 1371
rect 606 1366 612 1367
rect 758 1371 764 1372
rect 758 1367 759 1371
rect 763 1367 764 1371
rect 758 1366 764 1367
rect 902 1371 908 1372
rect 902 1367 903 1371
rect 907 1367 908 1371
rect 902 1366 908 1367
rect 1030 1371 1036 1372
rect 1030 1367 1031 1371
rect 1035 1367 1036 1371
rect 1030 1366 1036 1367
rect 1158 1371 1164 1372
rect 1158 1367 1159 1371
rect 1163 1367 1164 1371
rect 1158 1366 1164 1367
rect 1286 1371 1292 1372
rect 1286 1367 1287 1371
rect 1291 1367 1292 1371
rect 1286 1366 1292 1367
rect 1414 1371 1420 1372
rect 1414 1367 1415 1371
rect 1419 1367 1420 1371
rect 1766 1368 1767 1372
rect 1771 1368 1772 1372
rect 1766 1367 1772 1368
rect 1806 1371 1812 1372
rect 1806 1367 1807 1371
rect 1811 1367 1812 1371
rect 3462 1371 3468 1372
rect 1414 1366 1420 1367
rect 1806 1366 1812 1367
rect 2094 1368 2100 1369
rect 110 1355 116 1356
rect 110 1351 111 1355
rect 115 1351 116 1355
rect 1766 1355 1772 1356
rect 110 1350 116 1351
rect 134 1352 140 1353
rect 112 1327 114 1350
rect 134 1348 135 1352
rect 139 1348 140 1352
rect 134 1347 140 1348
rect 278 1352 284 1353
rect 278 1348 279 1352
rect 283 1348 284 1352
rect 278 1347 284 1348
rect 446 1352 452 1353
rect 446 1348 447 1352
rect 451 1348 452 1352
rect 446 1347 452 1348
rect 606 1352 612 1353
rect 606 1348 607 1352
rect 611 1348 612 1352
rect 606 1347 612 1348
rect 758 1352 764 1353
rect 758 1348 759 1352
rect 763 1348 764 1352
rect 758 1347 764 1348
rect 902 1352 908 1353
rect 902 1348 903 1352
rect 907 1348 908 1352
rect 902 1347 908 1348
rect 1030 1352 1036 1353
rect 1030 1348 1031 1352
rect 1035 1348 1036 1352
rect 1030 1347 1036 1348
rect 1158 1352 1164 1353
rect 1158 1348 1159 1352
rect 1163 1348 1164 1352
rect 1158 1347 1164 1348
rect 1286 1352 1292 1353
rect 1286 1348 1287 1352
rect 1291 1348 1292 1352
rect 1286 1347 1292 1348
rect 1414 1352 1420 1353
rect 1414 1348 1415 1352
rect 1419 1348 1420 1352
rect 1766 1351 1767 1355
rect 1771 1351 1772 1355
rect 1766 1350 1772 1351
rect 1414 1347 1420 1348
rect 136 1327 138 1347
rect 280 1327 282 1347
rect 448 1327 450 1347
rect 608 1327 610 1347
rect 760 1327 762 1347
rect 904 1327 906 1347
rect 1032 1327 1034 1347
rect 1160 1327 1162 1347
rect 1288 1327 1290 1347
rect 1416 1327 1418 1347
rect 1768 1327 1770 1350
rect 1808 1343 1810 1366
rect 2094 1364 2095 1368
rect 2099 1364 2100 1368
rect 2094 1363 2100 1364
rect 2198 1368 2204 1369
rect 2198 1364 2199 1368
rect 2203 1364 2204 1368
rect 2198 1363 2204 1364
rect 2318 1368 2324 1369
rect 2318 1364 2319 1368
rect 2323 1364 2324 1368
rect 2318 1363 2324 1364
rect 2454 1368 2460 1369
rect 2454 1364 2455 1368
rect 2459 1364 2460 1368
rect 2454 1363 2460 1364
rect 2598 1368 2604 1369
rect 2598 1364 2599 1368
rect 2603 1364 2604 1368
rect 2598 1363 2604 1364
rect 2742 1368 2748 1369
rect 2742 1364 2743 1368
rect 2747 1364 2748 1368
rect 2742 1363 2748 1364
rect 2886 1368 2892 1369
rect 2886 1364 2887 1368
rect 2891 1364 2892 1368
rect 2886 1363 2892 1364
rect 3030 1368 3036 1369
rect 3030 1364 3031 1368
rect 3035 1364 3036 1368
rect 3030 1363 3036 1364
rect 3174 1368 3180 1369
rect 3174 1364 3175 1368
rect 3179 1364 3180 1368
rect 3174 1363 3180 1364
rect 3326 1368 3332 1369
rect 3326 1364 3327 1368
rect 3331 1364 3332 1368
rect 3462 1367 3463 1371
rect 3467 1367 3468 1371
rect 3462 1366 3468 1367
rect 3326 1363 3332 1364
rect 2096 1343 2098 1363
rect 2200 1343 2202 1363
rect 2320 1343 2322 1363
rect 2456 1343 2458 1363
rect 2600 1343 2602 1363
rect 2744 1343 2746 1363
rect 2888 1343 2890 1363
rect 3032 1343 3034 1363
rect 3176 1343 3178 1363
rect 3328 1343 3330 1363
rect 3464 1343 3466 1366
rect 1807 1342 1811 1343
rect 1807 1337 1811 1338
rect 2095 1342 2099 1343
rect 2095 1337 2099 1338
rect 2103 1342 2107 1343
rect 2103 1337 2107 1338
rect 2199 1342 2203 1343
rect 2199 1337 2203 1338
rect 2239 1342 2243 1343
rect 2239 1337 2243 1338
rect 2319 1342 2323 1343
rect 2319 1337 2323 1338
rect 2383 1342 2387 1343
rect 2383 1337 2387 1338
rect 2455 1342 2459 1343
rect 2455 1337 2459 1338
rect 2535 1342 2539 1343
rect 2535 1337 2539 1338
rect 2599 1342 2603 1343
rect 2599 1337 2603 1338
rect 2687 1342 2691 1343
rect 2687 1337 2691 1338
rect 2743 1342 2747 1343
rect 2743 1337 2747 1338
rect 2839 1342 2843 1343
rect 2839 1337 2843 1338
rect 2887 1342 2891 1343
rect 2887 1337 2891 1338
rect 2991 1342 2995 1343
rect 2991 1337 2995 1338
rect 3031 1342 3035 1343
rect 3031 1337 3035 1338
rect 3143 1342 3147 1343
rect 3143 1337 3147 1338
rect 3175 1342 3179 1343
rect 3175 1337 3179 1338
rect 3303 1342 3307 1343
rect 3303 1337 3307 1338
rect 3327 1342 3331 1343
rect 3327 1337 3331 1338
rect 3463 1342 3467 1343
rect 3463 1337 3467 1338
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 135 1326 139 1327
rect 135 1321 139 1322
rect 279 1326 283 1327
rect 279 1321 283 1322
rect 439 1326 443 1327
rect 439 1321 443 1322
rect 447 1326 451 1327
rect 447 1321 451 1322
rect 583 1326 587 1327
rect 583 1321 587 1322
rect 607 1326 611 1327
rect 607 1321 611 1322
rect 719 1326 723 1327
rect 719 1321 723 1322
rect 759 1326 763 1327
rect 759 1321 763 1322
rect 847 1326 851 1327
rect 847 1321 851 1322
rect 903 1326 907 1327
rect 903 1321 907 1322
rect 967 1326 971 1327
rect 967 1321 971 1322
rect 1031 1326 1035 1327
rect 1031 1321 1035 1322
rect 1079 1326 1083 1327
rect 1079 1321 1083 1322
rect 1159 1326 1163 1327
rect 1159 1321 1163 1322
rect 1191 1326 1195 1327
rect 1191 1321 1195 1322
rect 1287 1326 1291 1327
rect 1287 1321 1291 1322
rect 1311 1326 1315 1327
rect 1311 1321 1315 1322
rect 1415 1326 1419 1327
rect 1415 1321 1419 1322
rect 1767 1326 1771 1327
rect 1767 1321 1771 1322
rect 112 1302 114 1321
rect 136 1305 138 1321
rect 280 1305 282 1321
rect 440 1305 442 1321
rect 584 1305 586 1321
rect 720 1305 722 1321
rect 848 1305 850 1321
rect 968 1305 970 1321
rect 1080 1305 1082 1321
rect 1192 1305 1194 1321
rect 1312 1305 1314 1321
rect 134 1304 140 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 134 1300 135 1304
rect 139 1300 140 1304
rect 134 1299 140 1300
rect 278 1304 284 1305
rect 278 1300 279 1304
rect 283 1300 284 1304
rect 278 1299 284 1300
rect 438 1304 444 1305
rect 438 1300 439 1304
rect 443 1300 444 1304
rect 438 1299 444 1300
rect 582 1304 588 1305
rect 582 1300 583 1304
rect 587 1300 588 1304
rect 582 1299 588 1300
rect 718 1304 724 1305
rect 718 1300 719 1304
rect 723 1300 724 1304
rect 718 1299 724 1300
rect 846 1304 852 1305
rect 846 1300 847 1304
rect 851 1300 852 1304
rect 846 1299 852 1300
rect 966 1304 972 1305
rect 966 1300 967 1304
rect 971 1300 972 1304
rect 966 1299 972 1300
rect 1078 1304 1084 1305
rect 1078 1300 1079 1304
rect 1083 1300 1084 1304
rect 1078 1299 1084 1300
rect 1190 1304 1196 1305
rect 1190 1300 1191 1304
rect 1195 1300 1196 1304
rect 1190 1299 1196 1300
rect 1310 1304 1316 1305
rect 1310 1300 1311 1304
rect 1315 1300 1316 1304
rect 1768 1302 1770 1321
rect 1808 1318 1810 1337
rect 2104 1321 2106 1337
rect 2240 1321 2242 1337
rect 2384 1321 2386 1337
rect 2536 1321 2538 1337
rect 2688 1321 2690 1337
rect 2840 1321 2842 1337
rect 2992 1321 2994 1337
rect 3144 1321 3146 1337
rect 3304 1321 3306 1337
rect 2102 1320 2108 1321
rect 1806 1317 1812 1318
rect 1806 1313 1807 1317
rect 1811 1313 1812 1317
rect 2102 1316 2103 1320
rect 2107 1316 2108 1320
rect 2102 1315 2108 1316
rect 2238 1320 2244 1321
rect 2238 1316 2239 1320
rect 2243 1316 2244 1320
rect 2238 1315 2244 1316
rect 2382 1320 2388 1321
rect 2382 1316 2383 1320
rect 2387 1316 2388 1320
rect 2382 1315 2388 1316
rect 2534 1320 2540 1321
rect 2534 1316 2535 1320
rect 2539 1316 2540 1320
rect 2534 1315 2540 1316
rect 2686 1320 2692 1321
rect 2686 1316 2687 1320
rect 2691 1316 2692 1320
rect 2686 1315 2692 1316
rect 2838 1320 2844 1321
rect 2838 1316 2839 1320
rect 2843 1316 2844 1320
rect 2838 1315 2844 1316
rect 2990 1320 2996 1321
rect 2990 1316 2991 1320
rect 2995 1316 2996 1320
rect 2990 1315 2996 1316
rect 3142 1320 3148 1321
rect 3142 1316 3143 1320
rect 3147 1316 3148 1320
rect 3142 1315 3148 1316
rect 3302 1320 3308 1321
rect 3302 1316 3303 1320
rect 3307 1316 3308 1320
rect 3464 1318 3466 1337
rect 3302 1315 3308 1316
rect 3462 1317 3468 1318
rect 1806 1312 1812 1313
rect 3462 1313 3463 1317
rect 3467 1313 3468 1317
rect 3462 1312 3468 1313
rect 1310 1299 1316 1300
rect 1766 1301 1772 1302
rect 2102 1301 2108 1302
rect 110 1296 116 1297
rect 1766 1297 1767 1301
rect 1771 1297 1772 1301
rect 1766 1296 1772 1297
rect 1806 1300 1812 1301
rect 1806 1296 1807 1300
rect 1811 1296 1812 1300
rect 2102 1297 2103 1301
rect 2107 1297 2108 1301
rect 2102 1296 2108 1297
rect 2238 1301 2244 1302
rect 2238 1297 2239 1301
rect 2243 1297 2244 1301
rect 2238 1296 2244 1297
rect 2382 1301 2388 1302
rect 2382 1297 2383 1301
rect 2387 1297 2388 1301
rect 2382 1296 2388 1297
rect 2534 1301 2540 1302
rect 2534 1297 2535 1301
rect 2539 1297 2540 1301
rect 2534 1296 2540 1297
rect 2686 1301 2692 1302
rect 2686 1297 2687 1301
rect 2691 1297 2692 1301
rect 2686 1296 2692 1297
rect 2838 1301 2844 1302
rect 2838 1297 2839 1301
rect 2843 1297 2844 1301
rect 2838 1296 2844 1297
rect 2990 1301 2996 1302
rect 2990 1297 2991 1301
rect 2995 1297 2996 1301
rect 2990 1296 2996 1297
rect 3142 1301 3148 1302
rect 3142 1297 3143 1301
rect 3147 1297 3148 1301
rect 3142 1296 3148 1297
rect 3302 1301 3308 1302
rect 3302 1297 3303 1301
rect 3307 1297 3308 1301
rect 3302 1296 3308 1297
rect 3462 1300 3468 1301
rect 3462 1296 3463 1300
rect 3467 1296 3468 1300
rect 1806 1295 1812 1296
rect 134 1285 140 1286
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 134 1281 135 1285
rect 139 1281 140 1285
rect 134 1280 140 1281
rect 278 1285 284 1286
rect 278 1281 279 1285
rect 283 1281 284 1285
rect 278 1280 284 1281
rect 438 1285 444 1286
rect 438 1281 439 1285
rect 443 1281 444 1285
rect 438 1280 444 1281
rect 582 1285 588 1286
rect 582 1281 583 1285
rect 587 1281 588 1285
rect 582 1280 588 1281
rect 718 1285 724 1286
rect 718 1281 719 1285
rect 723 1281 724 1285
rect 718 1280 724 1281
rect 846 1285 852 1286
rect 846 1281 847 1285
rect 851 1281 852 1285
rect 846 1280 852 1281
rect 966 1285 972 1286
rect 966 1281 967 1285
rect 971 1281 972 1285
rect 966 1280 972 1281
rect 1078 1285 1084 1286
rect 1078 1281 1079 1285
rect 1083 1281 1084 1285
rect 1078 1280 1084 1281
rect 1190 1285 1196 1286
rect 1190 1281 1191 1285
rect 1195 1281 1196 1285
rect 1190 1280 1196 1281
rect 1310 1285 1316 1286
rect 1310 1281 1311 1285
rect 1315 1281 1316 1285
rect 1310 1280 1316 1281
rect 1766 1284 1772 1285
rect 1766 1280 1767 1284
rect 1771 1280 1772 1284
rect 110 1279 116 1280
rect 112 1259 114 1279
rect 136 1259 138 1280
rect 280 1259 282 1280
rect 440 1259 442 1280
rect 584 1259 586 1280
rect 720 1259 722 1280
rect 848 1259 850 1280
rect 968 1259 970 1280
rect 1080 1259 1082 1280
rect 1192 1259 1194 1280
rect 1312 1259 1314 1280
rect 1766 1279 1772 1280
rect 1808 1279 1810 1295
rect 2104 1279 2106 1296
rect 2240 1279 2242 1296
rect 2384 1279 2386 1296
rect 2536 1279 2538 1296
rect 2688 1279 2690 1296
rect 2840 1279 2842 1296
rect 2992 1279 2994 1296
rect 3144 1279 3146 1296
rect 3304 1279 3306 1296
rect 3462 1295 3468 1296
rect 3464 1279 3466 1295
rect 1768 1259 1770 1279
rect 1807 1278 1811 1279
rect 1807 1273 1811 1274
rect 1935 1278 1939 1279
rect 1935 1273 1939 1274
rect 2063 1278 2067 1279
rect 2063 1273 2067 1274
rect 2103 1278 2107 1279
rect 2103 1273 2107 1274
rect 2199 1278 2203 1279
rect 2199 1273 2203 1274
rect 2239 1278 2243 1279
rect 2239 1273 2243 1274
rect 2343 1278 2347 1279
rect 2343 1273 2347 1274
rect 2383 1278 2387 1279
rect 2383 1273 2387 1274
rect 2495 1278 2499 1279
rect 2495 1273 2499 1274
rect 2535 1278 2539 1279
rect 2535 1273 2539 1274
rect 2655 1278 2659 1279
rect 2655 1273 2659 1274
rect 2687 1278 2691 1279
rect 2687 1273 2691 1274
rect 2815 1278 2819 1279
rect 2815 1273 2819 1274
rect 2839 1278 2843 1279
rect 2839 1273 2843 1274
rect 2975 1278 2979 1279
rect 2975 1273 2979 1274
rect 2991 1278 2995 1279
rect 2991 1273 2995 1274
rect 3143 1278 3147 1279
rect 3143 1273 3147 1274
rect 3303 1278 3307 1279
rect 3303 1273 3307 1274
rect 3463 1278 3467 1279
rect 3463 1273 3467 1274
rect 111 1258 115 1259
rect 111 1253 115 1254
rect 135 1258 139 1259
rect 135 1253 139 1254
rect 239 1258 243 1259
rect 239 1253 243 1254
rect 279 1258 283 1259
rect 279 1253 283 1254
rect 367 1258 371 1259
rect 367 1253 371 1254
rect 439 1258 443 1259
rect 439 1253 443 1254
rect 495 1258 499 1259
rect 495 1253 499 1254
rect 583 1258 587 1259
rect 583 1253 587 1254
rect 615 1258 619 1259
rect 615 1253 619 1254
rect 719 1258 723 1259
rect 719 1253 723 1254
rect 735 1258 739 1259
rect 735 1253 739 1254
rect 847 1258 851 1259
rect 847 1253 851 1254
rect 959 1258 963 1259
rect 959 1253 963 1254
rect 967 1258 971 1259
rect 967 1253 971 1254
rect 1071 1258 1075 1259
rect 1071 1253 1075 1254
rect 1079 1258 1083 1259
rect 1079 1253 1083 1254
rect 1191 1258 1195 1259
rect 1191 1253 1195 1254
rect 1311 1258 1315 1259
rect 1311 1253 1315 1254
rect 1767 1258 1771 1259
rect 1808 1257 1810 1273
rect 1767 1253 1771 1254
rect 1806 1256 1812 1257
rect 1936 1256 1938 1273
rect 2064 1256 2066 1273
rect 2200 1256 2202 1273
rect 2344 1256 2346 1273
rect 2496 1256 2498 1273
rect 2656 1256 2658 1273
rect 2816 1256 2818 1273
rect 2976 1256 2978 1273
rect 3144 1256 3146 1273
rect 3464 1257 3466 1273
rect 3462 1256 3468 1257
rect 112 1237 114 1253
rect 110 1236 116 1237
rect 136 1236 138 1253
rect 240 1236 242 1253
rect 368 1236 370 1253
rect 496 1236 498 1253
rect 616 1236 618 1253
rect 736 1236 738 1253
rect 848 1236 850 1253
rect 960 1236 962 1253
rect 1072 1236 1074 1253
rect 1192 1236 1194 1253
rect 1768 1237 1770 1253
rect 1806 1252 1807 1256
rect 1811 1252 1812 1256
rect 1806 1251 1812 1252
rect 1934 1255 1940 1256
rect 1934 1251 1935 1255
rect 1939 1251 1940 1255
rect 1934 1250 1940 1251
rect 2062 1255 2068 1256
rect 2062 1251 2063 1255
rect 2067 1251 2068 1255
rect 2062 1250 2068 1251
rect 2198 1255 2204 1256
rect 2198 1251 2199 1255
rect 2203 1251 2204 1255
rect 2198 1250 2204 1251
rect 2342 1255 2348 1256
rect 2342 1251 2343 1255
rect 2347 1251 2348 1255
rect 2342 1250 2348 1251
rect 2494 1255 2500 1256
rect 2494 1251 2495 1255
rect 2499 1251 2500 1255
rect 2494 1250 2500 1251
rect 2654 1255 2660 1256
rect 2654 1251 2655 1255
rect 2659 1251 2660 1255
rect 2654 1250 2660 1251
rect 2814 1255 2820 1256
rect 2814 1251 2815 1255
rect 2819 1251 2820 1255
rect 2814 1250 2820 1251
rect 2974 1255 2980 1256
rect 2974 1251 2975 1255
rect 2979 1251 2980 1255
rect 2974 1250 2980 1251
rect 3142 1255 3148 1256
rect 3142 1251 3143 1255
rect 3147 1251 3148 1255
rect 3462 1252 3463 1256
rect 3467 1252 3468 1256
rect 3462 1251 3468 1252
rect 3142 1250 3148 1251
rect 1806 1239 1812 1240
rect 1766 1236 1772 1237
rect 110 1232 111 1236
rect 115 1232 116 1236
rect 110 1231 116 1232
rect 134 1235 140 1236
rect 134 1231 135 1235
rect 139 1231 140 1235
rect 134 1230 140 1231
rect 238 1235 244 1236
rect 238 1231 239 1235
rect 243 1231 244 1235
rect 238 1230 244 1231
rect 366 1235 372 1236
rect 366 1231 367 1235
rect 371 1231 372 1235
rect 366 1230 372 1231
rect 494 1235 500 1236
rect 494 1231 495 1235
rect 499 1231 500 1235
rect 494 1230 500 1231
rect 614 1235 620 1236
rect 614 1231 615 1235
rect 619 1231 620 1235
rect 614 1230 620 1231
rect 734 1235 740 1236
rect 734 1231 735 1235
rect 739 1231 740 1235
rect 734 1230 740 1231
rect 846 1235 852 1236
rect 846 1231 847 1235
rect 851 1231 852 1235
rect 846 1230 852 1231
rect 958 1235 964 1236
rect 958 1231 959 1235
rect 963 1231 964 1235
rect 958 1230 964 1231
rect 1070 1235 1076 1236
rect 1070 1231 1071 1235
rect 1075 1231 1076 1235
rect 1070 1230 1076 1231
rect 1190 1235 1196 1236
rect 1190 1231 1191 1235
rect 1195 1231 1196 1235
rect 1766 1232 1767 1236
rect 1771 1232 1772 1236
rect 1806 1235 1807 1239
rect 1811 1235 1812 1239
rect 3462 1239 3468 1240
rect 1806 1234 1812 1235
rect 1934 1236 1940 1237
rect 1766 1231 1772 1232
rect 1190 1230 1196 1231
rect 110 1219 116 1220
rect 110 1215 111 1219
rect 115 1215 116 1219
rect 1766 1219 1772 1220
rect 110 1214 116 1215
rect 134 1216 140 1217
rect 112 1191 114 1214
rect 134 1212 135 1216
rect 139 1212 140 1216
rect 134 1211 140 1212
rect 238 1216 244 1217
rect 238 1212 239 1216
rect 243 1212 244 1216
rect 238 1211 244 1212
rect 366 1216 372 1217
rect 366 1212 367 1216
rect 371 1212 372 1216
rect 366 1211 372 1212
rect 494 1216 500 1217
rect 494 1212 495 1216
rect 499 1212 500 1216
rect 494 1211 500 1212
rect 614 1216 620 1217
rect 614 1212 615 1216
rect 619 1212 620 1216
rect 614 1211 620 1212
rect 734 1216 740 1217
rect 734 1212 735 1216
rect 739 1212 740 1216
rect 734 1211 740 1212
rect 846 1216 852 1217
rect 846 1212 847 1216
rect 851 1212 852 1216
rect 846 1211 852 1212
rect 958 1216 964 1217
rect 958 1212 959 1216
rect 963 1212 964 1216
rect 958 1211 964 1212
rect 1070 1216 1076 1217
rect 1070 1212 1071 1216
rect 1075 1212 1076 1216
rect 1070 1211 1076 1212
rect 1190 1216 1196 1217
rect 1190 1212 1191 1216
rect 1195 1212 1196 1216
rect 1766 1215 1767 1219
rect 1771 1215 1772 1219
rect 1808 1215 1810 1234
rect 1934 1232 1935 1236
rect 1939 1232 1940 1236
rect 1934 1231 1940 1232
rect 2062 1236 2068 1237
rect 2062 1232 2063 1236
rect 2067 1232 2068 1236
rect 2062 1231 2068 1232
rect 2198 1236 2204 1237
rect 2198 1232 2199 1236
rect 2203 1232 2204 1236
rect 2198 1231 2204 1232
rect 2342 1236 2348 1237
rect 2342 1232 2343 1236
rect 2347 1232 2348 1236
rect 2342 1231 2348 1232
rect 2494 1236 2500 1237
rect 2494 1232 2495 1236
rect 2499 1232 2500 1236
rect 2494 1231 2500 1232
rect 2654 1236 2660 1237
rect 2654 1232 2655 1236
rect 2659 1232 2660 1236
rect 2654 1231 2660 1232
rect 2814 1236 2820 1237
rect 2814 1232 2815 1236
rect 2819 1232 2820 1236
rect 2814 1231 2820 1232
rect 2974 1236 2980 1237
rect 2974 1232 2975 1236
rect 2979 1232 2980 1236
rect 2974 1231 2980 1232
rect 3142 1236 3148 1237
rect 3142 1232 3143 1236
rect 3147 1232 3148 1236
rect 3462 1235 3463 1239
rect 3467 1235 3468 1239
rect 3462 1234 3468 1235
rect 3142 1231 3148 1232
rect 1936 1215 1938 1231
rect 2064 1215 2066 1231
rect 2200 1215 2202 1231
rect 2344 1215 2346 1231
rect 2496 1215 2498 1231
rect 2656 1215 2658 1231
rect 2816 1215 2818 1231
rect 2976 1215 2978 1231
rect 3144 1215 3146 1231
rect 3464 1215 3466 1234
rect 1766 1214 1772 1215
rect 1807 1214 1811 1215
rect 1190 1211 1196 1212
rect 136 1191 138 1211
rect 240 1191 242 1211
rect 368 1191 370 1211
rect 496 1191 498 1211
rect 616 1191 618 1211
rect 736 1191 738 1211
rect 848 1191 850 1211
rect 960 1191 962 1211
rect 1072 1191 1074 1211
rect 1192 1191 1194 1211
rect 1768 1191 1770 1214
rect 1807 1209 1811 1210
rect 1831 1214 1835 1215
rect 1831 1209 1835 1210
rect 1935 1214 1939 1215
rect 1935 1209 1939 1210
rect 2063 1214 2067 1215
rect 2063 1209 2067 1210
rect 2079 1214 2083 1215
rect 2079 1209 2083 1210
rect 2199 1214 2203 1215
rect 2199 1209 2203 1210
rect 2231 1214 2235 1215
rect 2231 1209 2235 1210
rect 2343 1214 2347 1215
rect 2343 1209 2347 1210
rect 2391 1214 2395 1215
rect 2391 1209 2395 1210
rect 2495 1214 2499 1215
rect 2495 1209 2499 1210
rect 2543 1214 2547 1215
rect 2543 1209 2547 1210
rect 2655 1214 2659 1215
rect 2655 1209 2659 1210
rect 2695 1214 2699 1215
rect 2695 1209 2699 1210
rect 2815 1214 2819 1215
rect 2815 1209 2819 1210
rect 2847 1214 2851 1215
rect 2847 1209 2851 1210
rect 2975 1214 2979 1215
rect 2975 1209 2979 1210
rect 2999 1214 3003 1215
rect 2999 1209 3003 1210
rect 3143 1214 3147 1215
rect 3143 1209 3147 1210
rect 3159 1214 3163 1215
rect 3159 1209 3163 1210
rect 3463 1214 3467 1215
rect 3463 1209 3467 1210
rect 111 1190 115 1191
rect 111 1185 115 1186
rect 135 1190 139 1191
rect 135 1185 139 1186
rect 239 1190 243 1191
rect 239 1185 243 1186
rect 367 1190 371 1191
rect 367 1185 371 1186
rect 375 1190 379 1191
rect 375 1185 379 1186
rect 495 1190 499 1191
rect 495 1185 499 1186
rect 511 1190 515 1191
rect 511 1185 515 1186
rect 615 1190 619 1191
rect 615 1185 619 1186
rect 655 1190 659 1191
rect 655 1185 659 1186
rect 735 1190 739 1191
rect 735 1185 739 1186
rect 791 1190 795 1191
rect 791 1185 795 1186
rect 847 1190 851 1191
rect 847 1185 851 1186
rect 927 1190 931 1191
rect 927 1185 931 1186
rect 959 1190 963 1191
rect 959 1185 963 1186
rect 1063 1190 1067 1191
rect 1063 1185 1067 1186
rect 1071 1190 1075 1191
rect 1071 1185 1075 1186
rect 1191 1190 1195 1191
rect 1191 1185 1195 1186
rect 1199 1190 1203 1191
rect 1199 1185 1203 1186
rect 1335 1190 1339 1191
rect 1335 1185 1339 1186
rect 1767 1190 1771 1191
rect 1808 1190 1810 1209
rect 1832 1193 1834 1209
rect 1936 1193 1938 1209
rect 2080 1193 2082 1209
rect 2232 1193 2234 1209
rect 2392 1193 2394 1209
rect 2544 1193 2546 1209
rect 2696 1193 2698 1209
rect 2848 1193 2850 1209
rect 3000 1193 3002 1209
rect 3160 1193 3162 1209
rect 1830 1192 1836 1193
rect 1767 1185 1771 1186
rect 1806 1189 1812 1190
rect 1806 1185 1807 1189
rect 1811 1185 1812 1189
rect 1830 1188 1831 1192
rect 1835 1188 1836 1192
rect 1830 1187 1836 1188
rect 1934 1192 1940 1193
rect 1934 1188 1935 1192
rect 1939 1188 1940 1192
rect 1934 1187 1940 1188
rect 2078 1192 2084 1193
rect 2078 1188 2079 1192
rect 2083 1188 2084 1192
rect 2078 1187 2084 1188
rect 2230 1192 2236 1193
rect 2230 1188 2231 1192
rect 2235 1188 2236 1192
rect 2230 1187 2236 1188
rect 2390 1192 2396 1193
rect 2390 1188 2391 1192
rect 2395 1188 2396 1192
rect 2390 1187 2396 1188
rect 2542 1192 2548 1193
rect 2542 1188 2543 1192
rect 2547 1188 2548 1192
rect 2542 1187 2548 1188
rect 2694 1192 2700 1193
rect 2694 1188 2695 1192
rect 2699 1188 2700 1192
rect 2694 1187 2700 1188
rect 2846 1192 2852 1193
rect 2846 1188 2847 1192
rect 2851 1188 2852 1192
rect 2846 1187 2852 1188
rect 2998 1192 3004 1193
rect 2998 1188 2999 1192
rect 3003 1188 3004 1192
rect 2998 1187 3004 1188
rect 3158 1192 3164 1193
rect 3158 1188 3159 1192
rect 3163 1188 3164 1192
rect 3464 1190 3466 1209
rect 3158 1187 3164 1188
rect 3462 1189 3468 1190
rect 112 1166 114 1185
rect 136 1169 138 1185
rect 240 1169 242 1185
rect 376 1169 378 1185
rect 512 1169 514 1185
rect 656 1169 658 1185
rect 792 1169 794 1185
rect 928 1169 930 1185
rect 1064 1169 1066 1185
rect 1200 1169 1202 1185
rect 1336 1169 1338 1185
rect 134 1168 140 1169
rect 110 1165 116 1166
rect 110 1161 111 1165
rect 115 1161 116 1165
rect 134 1164 135 1168
rect 139 1164 140 1168
rect 134 1163 140 1164
rect 238 1168 244 1169
rect 238 1164 239 1168
rect 243 1164 244 1168
rect 238 1163 244 1164
rect 374 1168 380 1169
rect 374 1164 375 1168
rect 379 1164 380 1168
rect 374 1163 380 1164
rect 510 1168 516 1169
rect 510 1164 511 1168
rect 515 1164 516 1168
rect 510 1163 516 1164
rect 654 1168 660 1169
rect 654 1164 655 1168
rect 659 1164 660 1168
rect 654 1163 660 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 926 1168 932 1169
rect 926 1164 927 1168
rect 931 1164 932 1168
rect 926 1163 932 1164
rect 1062 1168 1068 1169
rect 1062 1164 1063 1168
rect 1067 1164 1068 1168
rect 1062 1163 1068 1164
rect 1198 1168 1204 1169
rect 1198 1164 1199 1168
rect 1203 1164 1204 1168
rect 1198 1163 1204 1164
rect 1334 1168 1340 1169
rect 1334 1164 1335 1168
rect 1339 1164 1340 1168
rect 1768 1166 1770 1185
rect 1806 1184 1812 1185
rect 3462 1185 3463 1189
rect 3467 1185 3468 1189
rect 3462 1184 3468 1185
rect 1830 1173 1836 1174
rect 1806 1172 1812 1173
rect 1806 1168 1807 1172
rect 1811 1168 1812 1172
rect 1830 1169 1831 1173
rect 1835 1169 1836 1173
rect 1830 1168 1836 1169
rect 1934 1173 1940 1174
rect 1934 1169 1935 1173
rect 1939 1169 1940 1173
rect 1934 1168 1940 1169
rect 2078 1173 2084 1174
rect 2078 1169 2079 1173
rect 2083 1169 2084 1173
rect 2078 1168 2084 1169
rect 2230 1173 2236 1174
rect 2230 1169 2231 1173
rect 2235 1169 2236 1173
rect 2230 1168 2236 1169
rect 2390 1173 2396 1174
rect 2390 1169 2391 1173
rect 2395 1169 2396 1173
rect 2390 1168 2396 1169
rect 2542 1173 2548 1174
rect 2542 1169 2543 1173
rect 2547 1169 2548 1173
rect 2542 1168 2548 1169
rect 2694 1173 2700 1174
rect 2694 1169 2695 1173
rect 2699 1169 2700 1173
rect 2694 1168 2700 1169
rect 2846 1173 2852 1174
rect 2846 1169 2847 1173
rect 2851 1169 2852 1173
rect 2846 1168 2852 1169
rect 2998 1173 3004 1174
rect 2998 1169 2999 1173
rect 3003 1169 3004 1173
rect 2998 1168 3004 1169
rect 3158 1173 3164 1174
rect 3158 1169 3159 1173
rect 3163 1169 3164 1173
rect 3158 1168 3164 1169
rect 3462 1172 3468 1173
rect 3462 1168 3463 1172
rect 3467 1168 3468 1172
rect 1806 1167 1812 1168
rect 1334 1163 1340 1164
rect 1766 1165 1772 1166
rect 110 1160 116 1161
rect 1766 1161 1767 1165
rect 1771 1161 1772 1165
rect 1766 1160 1772 1161
rect 134 1149 140 1150
rect 110 1148 116 1149
rect 110 1144 111 1148
rect 115 1144 116 1148
rect 134 1145 135 1149
rect 139 1145 140 1149
rect 134 1144 140 1145
rect 238 1149 244 1150
rect 238 1145 239 1149
rect 243 1145 244 1149
rect 238 1144 244 1145
rect 374 1149 380 1150
rect 374 1145 375 1149
rect 379 1145 380 1149
rect 374 1144 380 1145
rect 510 1149 516 1150
rect 510 1145 511 1149
rect 515 1145 516 1149
rect 510 1144 516 1145
rect 654 1149 660 1150
rect 654 1145 655 1149
rect 659 1145 660 1149
rect 654 1144 660 1145
rect 790 1149 796 1150
rect 790 1145 791 1149
rect 795 1145 796 1149
rect 790 1144 796 1145
rect 926 1149 932 1150
rect 926 1145 927 1149
rect 931 1145 932 1149
rect 926 1144 932 1145
rect 1062 1149 1068 1150
rect 1062 1145 1063 1149
rect 1067 1145 1068 1149
rect 1062 1144 1068 1145
rect 1198 1149 1204 1150
rect 1198 1145 1199 1149
rect 1203 1145 1204 1149
rect 1198 1144 1204 1145
rect 1334 1149 1340 1150
rect 1334 1145 1335 1149
rect 1339 1145 1340 1149
rect 1334 1144 1340 1145
rect 1766 1148 1772 1149
rect 1766 1144 1767 1148
rect 1771 1144 1772 1148
rect 110 1143 116 1144
rect 112 1123 114 1143
rect 136 1123 138 1144
rect 240 1123 242 1144
rect 376 1123 378 1144
rect 512 1123 514 1144
rect 656 1123 658 1144
rect 792 1123 794 1144
rect 928 1123 930 1144
rect 1064 1123 1066 1144
rect 1200 1123 1202 1144
rect 1336 1123 1338 1144
rect 1766 1143 1772 1144
rect 1768 1123 1770 1143
rect 1808 1139 1810 1167
rect 1832 1139 1834 1168
rect 1936 1139 1938 1168
rect 2080 1139 2082 1168
rect 2232 1139 2234 1168
rect 2392 1139 2394 1168
rect 2544 1139 2546 1168
rect 2696 1139 2698 1168
rect 2848 1139 2850 1168
rect 3000 1139 3002 1168
rect 3160 1139 3162 1168
rect 3462 1167 3468 1168
rect 3464 1139 3466 1167
rect 1807 1138 1811 1139
rect 1807 1133 1811 1134
rect 1831 1138 1835 1139
rect 1831 1133 1835 1134
rect 1863 1138 1867 1139
rect 1863 1133 1867 1134
rect 1935 1138 1939 1139
rect 1935 1133 1939 1134
rect 1983 1138 1987 1139
rect 1983 1133 1987 1134
rect 2079 1138 2083 1139
rect 2079 1133 2083 1134
rect 2111 1138 2115 1139
rect 2111 1133 2115 1134
rect 2231 1138 2235 1139
rect 2231 1133 2235 1134
rect 2247 1138 2251 1139
rect 2247 1133 2251 1134
rect 2383 1138 2387 1139
rect 2383 1133 2387 1134
rect 2391 1138 2395 1139
rect 2391 1133 2395 1134
rect 2511 1138 2515 1139
rect 2511 1133 2515 1134
rect 2543 1138 2547 1139
rect 2543 1133 2547 1134
rect 2639 1138 2643 1139
rect 2639 1133 2643 1134
rect 2695 1138 2699 1139
rect 2695 1133 2699 1134
rect 2759 1138 2763 1139
rect 2759 1133 2763 1134
rect 2847 1138 2851 1139
rect 2847 1133 2851 1134
rect 2871 1138 2875 1139
rect 2871 1133 2875 1134
rect 2975 1138 2979 1139
rect 2975 1133 2979 1134
rect 2999 1138 3003 1139
rect 2999 1133 3003 1134
rect 3079 1138 3083 1139
rect 3079 1133 3083 1134
rect 3159 1138 3163 1139
rect 3159 1133 3163 1134
rect 3183 1138 3187 1139
rect 3183 1133 3187 1134
rect 3279 1138 3283 1139
rect 3279 1133 3283 1134
rect 3367 1138 3371 1139
rect 3367 1133 3371 1134
rect 3463 1138 3467 1139
rect 3463 1133 3467 1134
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 135 1122 139 1123
rect 135 1117 139 1118
rect 191 1122 195 1123
rect 191 1117 195 1118
rect 239 1122 243 1123
rect 239 1117 243 1118
rect 335 1122 339 1123
rect 335 1117 339 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 495 1122 499 1123
rect 495 1117 499 1118
rect 511 1122 515 1123
rect 511 1117 515 1118
rect 655 1122 659 1123
rect 655 1117 659 1118
rect 791 1122 795 1123
rect 791 1117 795 1118
rect 815 1122 819 1123
rect 815 1117 819 1118
rect 927 1122 931 1123
rect 927 1117 931 1118
rect 967 1122 971 1123
rect 967 1117 971 1118
rect 1063 1122 1067 1123
rect 1063 1117 1067 1118
rect 1119 1122 1123 1123
rect 1119 1117 1123 1118
rect 1199 1122 1203 1123
rect 1199 1117 1203 1118
rect 1263 1122 1267 1123
rect 1263 1117 1267 1118
rect 1335 1122 1339 1123
rect 1335 1117 1339 1118
rect 1407 1122 1411 1123
rect 1407 1117 1411 1118
rect 1559 1122 1563 1123
rect 1559 1117 1563 1118
rect 1767 1122 1771 1123
rect 1767 1117 1771 1118
rect 1808 1117 1810 1133
rect 112 1101 114 1117
rect 110 1100 116 1101
rect 192 1100 194 1117
rect 336 1100 338 1117
rect 496 1100 498 1117
rect 656 1100 658 1117
rect 816 1100 818 1117
rect 968 1100 970 1117
rect 1120 1100 1122 1117
rect 1264 1100 1266 1117
rect 1408 1100 1410 1117
rect 1560 1100 1562 1117
rect 1768 1101 1770 1117
rect 1806 1116 1812 1117
rect 1864 1116 1866 1133
rect 1984 1116 1986 1133
rect 2112 1116 2114 1133
rect 2248 1116 2250 1133
rect 2384 1116 2386 1133
rect 2512 1116 2514 1133
rect 2640 1116 2642 1133
rect 2760 1116 2762 1133
rect 2872 1116 2874 1133
rect 2976 1116 2978 1133
rect 3080 1116 3082 1133
rect 3184 1116 3186 1133
rect 3280 1116 3282 1133
rect 3368 1116 3370 1133
rect 3464 1117 3466 1133
rect 3462 1116 3468 1117
rect 1806 1112 1807 1116
rect 1811 1112 1812 1116
rect 1806 1111 1812 1112
rect 1862 1115 1868 1116
rect 1862 1111 1863 1115
rect 1867 1111 1868 1115
rect 1862 1110 1868 1111
rect 1982 1115 1988 1116
rect 1982 1111 1983 1115
rect 1987 1111 1988 1115
rect 1982 1110 1988 1111
rect 2110 1115 2116 1116
rect 2110 1111 2111 1115
rect 2115 1111 2116 1115
rect 2110 1110 2116 1111
rect 2246 1115 2252 1116
rect 2246 1111 2247 1115
rect 2251 1111 2252 1115
rect 2246 1110 2252 1111
rect 2382 1115 2388 1116
rect 2382 1111 2383 1115
rect 2387 1111 2388 1115
rect 2382 1110 2388 1111
rect 2510 1115 2516 1116
rect 2510 1111 2511 1115
rect 2515 1111 2516 1115
rect 2510 1110 2516 1111
rect 2638 1115 2644 1116
rect 2638 1111 2639 1115
rect 2643 1111 2644 1115
rect 2638 1110 2644 1111
rect 2758 1115 2764 1116
rect 2758 1111 2759 1115
rect 2763 1111 2764 1115
rect 2758 1110 2764 1111
rect 2870 1115 2876 1116
rect 2870 1111 2871 1115
rect 2875 1111 2876 1115
rect 2870 1110 2876 1111
rect 2974 1115 2980 1116
rect 2974 1111 2975 1115
rect 2979 1111 2980 1115
rect 2974 1110 2980 1111
rect 3078 1115 3084 1116
rect 3078 1111 3079 1115
rect 3083 1111 3084 1115
rect 3078 1110 3084 1111
rect 3182 1115 3188 1116
rect 3182 1111 3183 1115
rect 3187 1111 3188 1115
rect 3182 1110 3188 1111
rect 3278 1115 3284 1116
rect 3278 1111 3279 1115
rect 3283 1111 3284 1115
rect 3278 1110 3284 1111
rect 3366 1115 3372 1116
rect 3366 1111 3367 1115
rect 3371 1111 3372 1115
rect 3462 1112 3463 1116
rect 3467 1112 3468 1116
rect 3462 1111 3468 1112
rect 3366 1110 3372 1111
rect 1766 1100 1772 1101
rect 110 1096 111 1100
rect 115 1096 116 1100
rect 110 1095 116 1096
rect 190 1099 196 1100
rect 190 1095 191 1099
rect 195 1095 196 1099
rect 190 1094 196 1095
rect 334 1099 340 1100
rect 334 1095 335 1099
rect 339 1095 340 1099
rect 334 1094 340 1095
rect 494 1099 500 1100
rect 494 1095 495 1099
rect 499 1095 500 1099
rect 494 1094 500 1095
rect 654 1099 660 1100
rect 654 1095 655 1099
rect 659 1095 660 1099
rect 654 1094 660 1095
rect 814 1099 820 1100
rect 814 1095 815 1099
rect 819 1095 820 1099
rect 814 1094 820 1095
rect 966 1099 972 1100
rect 966 1095 967 1099
rect 971 1095 972 1099
rect 966 1094 972 1095
rect 1118 1099 1124 1100
rect 1118 1095 1119 1099
rect 1123 1095 1124 1099
rect 1118 1094 1124 1095
rect 1262 1099 1268 1100
rect 1262 1095 1263 1099
rect 1267 1095 1268 1099
rect 1262 1094 1268 1095
rect 1406 1099 1412 1100
rect 1406 1095 1407 1099
rect 1411 1095 1412 1099
rect 1406 1094 1412 1095
rect 1558 1099 1564 1100
rect 1558 1095 1559 1099
rect 1563 1095 1564 1099
rect 1766 1096 1767 1100
rect 1771 1096 1772 1100
rect 1766 1095 1772 1096
rect 1806 1099 1812 1100
rect 1806 1095 1807 1099
rect 1811 1095 1812 1099
rect 3462 1099 3468 1100
rect 1558 1094 1564 1095
rect 1806 1094 1812 1095
rect 1862 1096 1868 1097
rect 110 1083 116 1084
rect 110 1079 111 1083
rect 115 1079 116 1083
rect 1766 1083 1772 1084
rect 110 1078 116 1079
rect 190 1080 196 1081
rect 112 1051 114 1078
rect 190 1076 191 1080
rect 195 1076 196 1080
rect 190 1075 196 1076
rect 334 1080 340 1081
rect 334 1076 335 1080
rect 339 1076 340 1080
rect 334 1075 340 1076
rect 494 1080 500 1081
rect 494 1076 495 1080
rect 499 1076 500 1080
rect 494 1075 500 1076
rect 654 1080 660 1081
rect 654 1076 655 1080
rect 659 1076 660 1080
rect 654 1075 660 1076
rect 814 1080 820 1081
rect 814 1076 815 1080
rect 819 1076 820 1080
rect 814 1075 820 1076
rect 966 1080 972 1081
rect 966 1076 967 1080
rect 971 1076 972 1080
rect 966 1075 972 1076
rect 1118 1080 1124 1081
rect 1118 1076 1119 1080
rect 1123 1076 1124 1080
rect 1118 1075 1124 1076
rect 1262 1080 1268 1081
rect 1262 1076 1263 1080
rect 1267 1076 1268 1080
rect 1262 1075 1268 1076
rect 1406 1080 1412 1081
rect 1406 1076 1407 1080
rect 1411 1076 1412 1080
rect 1406 1075 1412 1076
rect 1558 1080 1564 1081
rect 1558 1076 1559 1080
rect 1563 1076 1564 1080
rect 1766 1079 1767 1083
rect 1771 1079 1772 1083
rect 1766 1078 1772 1079
rect 1558 1075 1564 1076
rect 192 1051 194 1075
rect 336 1051 338 1075
rect 496 1051 498 1075
rect 656 1051 658 1075
rect 816 1051 818 1075
rect 968 1051 970 1075
rect 1120 1051 1122 1075
rect 1264 1051 1266 1075
rect 1408 1051 1410 1075
rect 1560 1051 1562 1075
rect 1768 1051 1770 1078
rect 1808 1067 1810 1094
rect 1862 1092 1863 1096
rect 1867 1092 1868 1096
rect 1862 1091 1868 1092
rect 1982 1096 1988 1097
rect 1982 1092 1983 1096
rect 1987 1092 1988 1096
rect 1982 1091 1988 1092
rect 2110 1096 2116 1097
rect 2110 1092 2111 1096
rect 2115 1092 2116 1096
rect 2110 1091 2116 1092
rect 2246 1096 2252 1097
rect 2246 1092 2247 1096
rect 2251 1092 2252 1096
rect 2246 1091 2252 1092
rect 2382 1096 2388 1097
rect 2382 1092 2383 1096
rect 2387 1092 2388 1096
rect 2382 1091 2388 1092
rect 2510 1096 2516 1097
rect 2510 1092 2511 1096
rect 2515 1092 2516 1096
rect 2510 1091 2516 1092
rect 2638 1096 2644 1097
rect 2638 1092 2639 1096
rect 2643 1092 2644 1096
rect 2638 1091 2644 1092
rect 2758 1096 2764 1097
rect 2758 1092 2759 1096
rect 2763 1092 2764 1096
rect 2758 1091 2764 1092
rect 2870 1096 2876 1097
rect 2870 1092 2871 1096
rect 2875 1092 2876 1096
rect 2870 1091 2876 1092
rect 2974 1096 2980 1097
rect 2974 1092 2975 1096
rect 2979 1092 2980 1096
rect 2974 1091 2980 1092
rect 3078 1096 3084 1097
rect 3078 1092 3079 1096
rect 3083 1092 3084 1096
rect 3078 1091 3084 1092
rect 3182 1096 3188 1097
rect 3182 1092 3183 1096
rect 3187 1092 3188 1096
rect 3182 1091 3188 1092
rect 3278 1096 3284 1097
rect 3278 1092 3279 1096
rect 3283 1092 3284 1096
rect 3278 1091 3284 1092
rect 3366 1096 3372 1097
rect 3366 1092 3367 1096
rect 3371 1092 3372 1096
rect 3462 1095 3463 1099
rect 3467 1095 3468 1099
rect 3462 1094 3468 1095
rect 3366 1091 3372 1092
rect 1864 1067 1866 1091
rect 1984 1067 1986 1091
rect 2112 1067 2114 1091
rect 2248 1067 2250 1091
rect 2384 1067 2386 1091
rect 2512 1067 2514 1091
rect 2640 1067 2642 1091
rect 2760 1067 2762 1091
rect 2872 1067 2874 1091
rect 2976 1067 2978 1091
rect 3080 1067 3082 1091
rect 3184 1067 3186 1091
rect 3280 1067 3282 1091
rect 3368 1067 3370 1091
rect 3464 1067 3466 1094
rect 1807 1066 1811 1067
rect 1807 1061 1811 1062
rect 1863 1066 1867 1067
rect 1863 1061 1867 1062
rect 1983 1066 1987 1067
rect 1983 1061 1987 1062
rect 2103 1066 2107 1067
rect 2103 1061 2107 1062
rect 2111 1066 2115 1067
rect 2111 1061 2115 1062
rect 2191 1066 2195 1067
rect 2191 1061 2195 1062
rect 2247 1066 2251 1067
rect 2247 1061 2251 1062
rect 2279 1066 2283 1067
rect 2279 1061 2283 1062
rect 2367 1066 2371 1067
rect 2367 1061 2371 1062
rect 2383 1066 2387 1067
rect 2383 1061 2387 1062
rect 2455 1066 2459 1067
rect 2455 1061 2459 1062
rect 2511 1066 2515 1067
rect 2511 1061 2515 1062
rect 2543 1066 2547 1067
rect 2543 1061 2547 1062
rect 2631 1066 2635 1067
rect 2631 1061 2635 1062
rect 2639 1066 2643 1067
rect 2639 1061 2643 1062
rect 2719 1066 2723 1067
rect 2719 1061 2723 1062
rect 2759 1066 2763 1067
rect 2759 1061 2763 1062
rect 2807 1066 2811 1067
rect 2807 1061 2811 1062
rect 2871 1066 2875 1067
rect 2871 1061 2875 1062
rect 2975 1066 2979 1067
rect 2975 1061 2979 1062
rect 3079 1066 3083 1067
rect 3079 1061 3083 1062
rect 3183 1066 3187 1067
rect 3183 1061 3187 1062
rect 3279 1066 3283 1067
rect 3279 1061 3283 1062
rect 3367 1066 3371 1067
rect 3367 1061 3371 1062
rect 3463 1066 3467 1067
rect 3463 1061 3467 1062
rect 111 1050 115 1051
rect 111 1045 115 1046
rect 191 1050 195 1051
rect 191 1045 195 1046
rect 327 1050 331 1051
rect 327 1045 331 1046
rect 335 1050 339 1051
rect 335 1045 339 1046
rect 463 1050 467 1051
rect 463 1045 467 1046
rect 495 1050 499 1051
rect 495 1045 499 1046
rect 607 1050 611 1051
rect 607 1045 611 1046
rect 655 1050 659 1051
rect 655 1045 659 1046
rect 767 1050 771 1051
rect 767 1045 771 1046
rect 815 1050 819 1051
rect 815 1045 819 1046
rect 927 1050 931 1051
rect 927 1045 931 1046
rect 967 1050 971 1051
rect 967 1045 971 1046
rect 1079 1050 1083 1051
rect 1079 1045 1083 1046
rect 1119 1050 1123 1051
rect 1119 1045 1123 1046
rect 1231 1050 1235 1051
rect 1231 1045 1235 1046
rect 1263 1050 1267 1051
rect 1263 1045 1267 1046
rect 1383 1050 1387 1051
rect 1383 1045 1387 1046
rect 1407 1050 1411 1051
rect 1407 1045 1411 1046
rect 1535 1050 1539 1051
rect 1535 1045 1539 1046
rect 1559 1050 1563 1051
rect 1559 1045 1563 1046
rect 1671 1050 1675 1051
rect 1671 1045 1675 1046
rect 1767 1050 1771 1051
rect 1767 1045 1771 1046
rect 112 1026 114 1045
rect 328 1029 330 1045
rect 464 1029 466 1045
rect 608 1029 610 1045
rect 768 1029 770 1045
rect 928 1029 930 1045
rect 1080 1029 1082 1045
rect 1232 1029 1234 1045
rect 1384 1029 1386 1045
rect 1536 1029 1538 1045
rect 1672 1029 1674 1045
rect 326 1028 332 1029
rect 110 1025 116 1026
rect 110 1021 111 1025
rect 115 1021 116 1025
rect 326 1024 327 1028
rect 331 1024 332 1028
rect 326 1023 332 1024
rect 462 1028 468 1029
rect 462 1024 463 1028
rect 467 1024 468 1028
rect 462 1023 468 1024
rect 606 1028 612 1029
rect 606 1024 607 1028
rect 611 1024 612 1028
rect 606 1023 612 1024
rect 766 1028 772 1029
rect 766 1024 767 1028
rect 771 1024 772 1028
rect 766 1023 772 1024
rect 926 1028 932 1029
rect 926 1024 927 1028
rect 931 1024 932 1028
rect 926 1023 932 1024
rect 1078 1028 1084 1029
rect 1078 1024 1079 1028
rect 1083 1024 1084 1028
rect 1078 1023 1084 1024
rect 1230 1028 1236 1029
rect 1230 1024 1231 1028
rect 1235 1024 1236 1028
rect 1230 1023 1236 1024
rect 1382 1028 1388 1029
rect 1382 1024 1383 1028
rect 1387 1024 1388 1028
rect 1382 1023 1388 1024
rect 1534 1028 1540 1029
rect 1534 1024 1535 1028
rect 1539 1024 1540 1028
rect 1534 1023 1540 1024
rect 1670 1028 1676 1029
rect 1670 1024 1671 1028
rect 1675 1024 1676 1028
rect 1768 1026 1770 1045
rect 1808 1042 1810 1061
rect 2104 1045 2106 1061
rect 2192 1045 2194 1061
rect 2280 1045 2282 1061
rect 2368 1045 2370 1061
rect 2456 1045 2458 1061
rect 2544 1045 2546 1061
rect 2632 1045 2634 1061
rect 2720 1045 2722 1061
rect 2808 1045 2810 1061
rect 2102 1044 2108 1045
rect 1806 1041 1812 1042
rect 1806 1037 1807 1041
rect 1811 1037 1812 1041
rect 2102 1040 2103 1044
rect 2107 1040 2108 1044
rect 2102 1039 2108 1040
rect 2190 1044 2196 1045
rect 2190 1040 2191 1044
rect 2195 1040 2196 1044
rect 2190 1039 2196 1040
rect 2278 1044 2284 1045
rect 2278 1040 2279 1044
rect 2283 1040 2284 1044
rect 2278 1039 2284 1040
rect 2366 1044 2372 1045
rect 2366 1040 2367 1044
rect 2371 1040 2372 1044
rect 2366 1039 2372 1040
rect 2454 1044 2460 1045
rect 2454 1040 2455 1044
rect 2459 1040 2460 1044
rect 2454 1039 2460 1040
rect 2542 1044 2548 1045
rect 2542 1040 2543 1044
rect 2547 1040 2548 1044
rect 2542 1039 2548 1040
rect 2630 1044 2636 1045
rect 2630 1040 2631 1044
rect 2635 1040 2636 1044
rect 2630 1039 2636 1040
rect 2718 1044 2724 1045
rect 2718 1040 2719 1044
rect 2723 1040 2724 1044
rect 2718 1039 2724 1040
rect 2806 1044 2812 1045
rect 2806 1040 2807 1044
rect 2811 1040 2812 1044
rect 3464 1042 3466 1061
rect 2806 1039 2812 1040
rect 3462 1041 3468 1042
rect 1806 1036 1812 1037
rect 3462 1037 3463 1041
rect 3467 1037 3468 1041
rect 3462 1036 3468 1037
rect 1670 1023 1676 1024
rect 1766 1025 1772 1026
rect 2102 1025 2108 1026
rect 110 1020 116 1021
rect 1766 1021 1767 1025
rect 1771 1021 1772 1025
rect 1766 1020 1772 1021
rect 1806 1024 1812 1025
rect 1806 1020 1807 1024
rect 1811 1020 1812 1024
rect 2102 1021 2103 1025
rect 2107 1021 2108 1025
rect 2102 1020 2108 1021
rect 2190 1025 2196 1026
rect 2190 1021 2191 1025
rect 2195 1021 2196 1025
rect 2190 1020 2196 1021
rect 2278 1025 2284 1026
rect 2278 1021 2279 1025
rect 2283 1021 2284 1025
rect 2278 1020 2284 1021
rect 2366 1025 2372 1026
rect 2366 1021 2367 1025
rect 2371 1021 2372 1025
rect 2366 1020 2372 1021
rect 2454 1025 2460 1026
rect 2454 1021 2455 1025
rect 2459 1021 2460 1025
rect 2454 1020 2460 1021
rect 2542 1025 2548 1026
rect 2542 1021 2543 1025
rect 2547 1021 2548 1025
rect 2542 1020 2548 1021
rect 2630 1025 2636 1026
rect 2630 1021 2631 1025
rect 2635 1021 2636 1025
rect 2630 1020 2636 1021
rect 2718 1025 2724 1026
rect 2718 1021 2719 1025
rect 2723 1021 2724 1025
rect 2718 1020 2724 1021
rect 2806 1025 2812 1026
rect 2806 1021 2807 1025
rect 2811 1021 2812 1025
rect 2806 1020 2812 1021
rect 3462 1024 3468 1025
rect 3462 1020 3463 1024
rect 3467 1020 3468 1024
rect 1806 1019 1812 1020
rect 326 1009 332 1010
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 326 1005 327 1009
rect 331 1005 332 1009
rect 326 1004 332 1005
rect 462 1009 468 1010
rect 462 1005 463 1009
rect 467 1005 468 1009
rect 462 1004 468 1005
rect 606 1009 612 1010
rect 606 1005 607 1009
rect 611 1005 612 1009
rect 606 1004 612 1005
rect 766 1009 772 1010
rect 766 1005 767 1009
rect 771 1005 772 1009
rect 766 1004 772 1005
rect 926 1009 932 1010
rect 926 1005 927 1009
rect 931 1005 932 1009
rect 926 1004 932 1005
rect 1078 1009 1084 1010
rect 1078 1005 1079 1009
rect 1083 1005 1084 1009
rect 1078 1004 1084 1005
rect 1230 1009 1236 1010
rect 1230 1005 1231 1009
rect 1235 1005 1236 1009
rect 1230 1004 1236 1005
rect 1382 1009 1388 1010
rect 1382 1005 1383 1009
rect 1387 1005 1388 1009
rect 1382 1004 1388 1005
rect 1534 1009 1540 1010
rect 1534 1005 1535 1009
rect 1539 1005 1540 1009
rect 1534 1004 1540 1005
rect 1670 1009 1676 1010
rect 1670 1005 1671 1009
rect 1675 1005 1676 1009
rect 1670 1004 1676 1005
rect 1766 1008 1772 1009
rect 1766 1004 1767 1008
rect 1771 1004 1772 1008
rect 110 1003 116 1004
rect 112 983 114 1003
rect 328 983 330 1004
rect 464 983 466 1004
rect 608 983 610 1004
rect 768 983 770 1004
rect 928 983 930 1004
rect 1080 983 1082 1004
rect 1232 983 1234 1004
rect 1384 983 1386 1004
rect 1536 983 1538 1004
rect 1672 983 1674 1004
rect 1766 1003 1772 1004
rect 1808 1003 1810 1019
rect 2104 1003 2106 1020
rect 2192 1003 2194 1020
rect 2280 1003 2282 1020
rect 2368 1003 2370 1020
rect 2456 1003 2458 1020
rect 2544 1003 2546 1020
rect 2632 1003 2634 1020
rect 2720 1003 2722 1020
rect 2808 1003 2810 1020
rect 3462 1019 3468 1020
rect 3464 1003 3466 1019
rect 1768 983 1770 1003
rect 1807 1002 1811 1003
rect 1807 997 1811 998
rect 2103 1002 2107 1003
rect 2103 997 2107 998
rect 2191 1002 2195 1003
rect 2191 997 2195 998
rect 2279 1002 2283 1003
rect 2279 997 2283 998
rect 2311 1002 2315 1003
rect 2311 997 2315 998
rect 2367 1002 2371 1003
rect 2367 997 2371 998
rect 2407 1002 2411 1003
rect 2407 997 2411 998
rect 2455 1002 2459 1003
rect 2455 997 2459 998
rect 2511 1002 2515 1003
rect 2511 997 2515 998
rect 2543 1002 2547 1003
rect 2543 997 2547 998
rect 2623 1002 2627 1003
rect 2623 997 2627 998
rect 2631 1002 2635 1003
rect 2631 997 2635 998
rect 2719 1002 2723 1003
rect 2719 997 2723 998
rect 2751 1002 2755 1003
rect 2751 997 2755 998
rect 2807 1002 2811 1003
rect 2807 997 2811 998
rect 2895 1002 2899 1003
rect 2895 997 2899 998
rect 3055 1002 3059 1003
rect 3055 997 3059 998
rect 3223 1002 3227 1003
rect 3223 997 3227 998
rect 3367 1002 3371 1003
rect 3367 997 3371 998
rect 3463 1002 3467 1003
rect 3463 997 3467 998
rect 111 982 115 983
rect 111 977 115 978
rect 327 982 331 983
rect 327 977 331 978
rect 463 982 467 983
rect 463 977 467 978
rect 471 982 475 983
rect 471 977 475 978
rect 567 982 571 983
rect 567 977 571 978
rect 607 982 611 983
rect 607 977 611 978
rect 671 982 675 983
rect 671 977 675 978
rect 767 982 771 983
rect 767 977 771 978
rect 783 982 787 983
rect 783 977 787 978
rect 887 982 891 983
rect 887 977 891 978
rect 927 982 931 983
rect 927 977 931 978
rect 991 982 995 983
rect 991 977 995 978
rect 1079 982 1083 983
rect 1079 977 1083 978
rect 1095 982 1099 983
rect 1095 977 1099 978
rect 1199 982 1203 983
rect 1199 977 1203 978
rect 1231 982 1235 983
rect 1231 977 1235 978
rect 1295 982 1299 983
rect 1295 977 1299 978
rect 1383 982 1387 983
rect 1383 977 1387 978
rect 1391 982 1395 983
rect 1391 977 1395 978
rect 1487 982 1491 983
rect 1487 977 1491 978
rect 1535 982 1539 983
rect 1535 977 1539 978
rect 1583 982 1587 983
rect 1583 977 1587 978
rect 1671 982 1675 983
rect 1671 977 1675 978
rect 1767 982 1771 983
rect 1808 981 1810 997
rect 1767 977 1771 978
rect 1806 980 1812 981
rect 2312 980 2314 997
rect 2408 980 2410 997
rect 2512 980 2514 997
rect 2624 980 2626 997
rect 2752 980 2754 997
rect 2896 980 2898 997
rect 3056 980 3058 997
rect 3224 980 3226 997
rect 3368 980 3370 997
rect 3464 981 3466 997
rect 3462 980 3468 981
rect 112 961 114 977
rect 110 960 116 961
rect 472 960 474 977
rect 568 960 570 977
rect 672 960 674 977
rect 784 960 786 977
rect 888 960 890 977
rect 992 960 994 977
rect 1096 960 1098 977
rect 1200 960 1202 977
rect 1296 960 1298 977
rect 1392 960 1394 977
rect 1488 960 1490 977
rect 1584 960 1586 977
rect 1672 960 1674 977
rect 1768 961 1770 977
rect 1806 976 1807 980
rect 1811 976 1812 980
rect 1806 975 1812 976
rect 2310 979 2316 980
rect 2310 975 2311 979
rect 2315 975 2316 979
rect 2310 974 2316 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 2510 979 2516 980
rect 2510 975 2511 979
rect 2515 975 2516 979
rect 2510 974 2516 975
rect 2622 979 2628 980
rect 2622 975 2623 979
rect 2627 975 2628 979
rect 2622 974 2628 975
rect 2750 979 2756 980
rect 2750 975 2751 979
rect 2755 975 2756 979
rect 2750 974 2756 975
rect 2894 979 2900 980
rect 2894 975 2895 979
rect 2899 975 2900 979
rect 2894 974 2900 975
rect 3054 979 3060 980
rect 3054 975 3055 979
rect 3059 975 3060 979
rect 3054 974 3060 975
rect 3222 979 3228 980
rect 3222 975 3223 979
rect 3227 975 3228 979
rect 3222 974 3228 975
rect 3366 979 3372 980
rect 3366 975 3367 979
rect 3371 975 3372 979
rect 3462 976 3463 980
rect 3467 976 3468 980
rect 3462 975 3468 976
rect 3366 974 3372 975
rect 1806 963 1812 964
rect 1766 960 1772 961
rect 110 956 111 960
rect 115 956 116 960
rect 110 955 116 956
rect 470 959 476 960
rect 470 955 471 959
rect 475 955 476 959
rect 470 954 476 955
rect 566 959 572 960
rect 566 955 567 959
rect 571 955 572 959
rect 566 954 572 955
rect 670 959 676 960
rect 670 955 671 959
rect 675 955 676 959
rect 670 954 676 955
rect 782 959 788 960
rect 782 955 783 959
rect 787 955 788 959
rect 782 954 788 955
rect 886 959 892 960
rect 886 955 887 959
rect 891 955 892 959
rect 886 954 892 955
rect 990 959 996 960
rect 990 955 991 959
rect 995 955 996 959
rect 990 954 996 955
rect 1094 959 1100 960
rect 1094 955 1095 959
rect 1099 955 1100 959
rect 1094 954 1100 955
rect 1198 959 1204 960
rect 1198 955 1199 959
rect 1203 955 1204 959
rect 1198 954 1204 955
rect 1294 959 1300 960
rect 1294 955 1295 959
rect 1299 955 1300 959
rect 1294 954 1300 955
rect 1390 959 1396 960
rect 1390 955 1391 959
rect 1395 955 1396 959
rect 1390 954 1396 955
rect 1486 959 1492 960
rect 1486 955 1487 959
rect 1491 955 1492 959
rect 1486 954 1492 955
rect 1582 959 1588 960
rect 1582 955 1583 959
rect 1587 955 1588 959
rect 1582 954 1588 955
rect 1670 959 1676 960
rect 1670 955 1671 959
rect 1675 955 1676 959
rect 1766 956 1767 960
rect 1771 956 1772 960
rect 1806 959 1807 963
rect 1811 959 1812 963
rect 3462 963 3468 964
rect 1806 958 1812 959
rect 2310 960 2316 961
rect 1766 955 1772 956
rect 1670 954 1676 955
rect 110 943 116 944
rect 110 939 111 943
rect 115 939 116 943
rect 1766 943 1772 944
rect 110 938 116 939
rect 470 940 476 941
rect 112 915 114 938
rect 470 936 471 940
rect 475 936 476 940
rect 470 935 476 936
rect 566 940 572 941
rect 566 936 567 940
rect 571 936 572 940
rect 566 935 572 936
rect 670 940 676 941
rect 670 936 671 940
rect 675 936 676 940
rect 670 935 676 936
rect 782 940 788 941
rect 782 936 783 940
rect 787 936 788 940
rect 782 935 788 936
rect 886 940 892 941
rect 886 936 887 940
rect 891 936 892 940
rect 886 935 892 936
rect 990 940 996 941
rect 990 936 991 940
rect 995 936 996 940
rect 990 935 996 936
rect 1094 940 1100 941
rect 1094 936 1095 940
rect 1099 936 1100 940
rect 1094 935 1100 936
rect 1198 940 1204 941
rect 1198 936 1199 940
rect 1203 936 1204 940
rect 1198 935 1204 936
rect 1294 940 1300 941
rect 1294 936 1295 940
rect 1299 936 1300 940
rect 1294 935 1300 936
rect 1390 940 1396 941
rect 1390 936 1391 940
rect 1395 936 1396 940
rect 1390 935 1396 936
rect 1486 940 1492 941
rect 1486 936 1487 940
rect 1491 936 1492 940
rect 1486 935 1492 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1670 940 1676 941
rect 1670 936 1671 940
rect 1675 936 1676 940
rect 1766 939 1767 943
rect 1771 939 1772 943
rect 1766 938 1772 939
rect 1670 935 1676 936
rect 472 915 474 935
rect 568 915 570 935
rect 672 915 674 935
rect 784 915 786 935
rect 888 915 890 935
rect 992 915 994 935
rect 1096 915 1098 935
rect 1200 915 1202 935
rect 1296 915 1298 935
rect 1392 915 1394 935
rect 1488 915 1490 935
rect 1584 915 1586 935
rect 1672 915 1674 935
rect 1768 915 1770 938
rect 1808 927 1810 958
rect 2310 956 2311 960
rect 2315 956 2316 960
rect 2310 955 2316 956
rect 2406 960 2412 961
rect 2406 956 2407 960
rect 2411 956 2412 960
rect 2406 955 2412 956
rect 2510 960 2516 961
rect 2510 956 2511 960
rect 2515 956 2516 960
rect 2510 955 2516 956
rect 2622 960 2628 961
rect 2622 956 2623 960
rect 2627 956 2628 960
rect 2622 955 2628 956
rect 2750 960 2756 961
rect 2750 956 2751 960
rect 2755 956 2756 960
rect 2750 955 2756 956
rect 2894 960 2900 961
rect 2894 956 2895 960
rect 2899 956 2900 960
rect 2894 955 2900 956
rect 3054 960 3060 961
rect 3054 956 3055 960
rect 3059 956 3060 960
rect 3054 955 3060 956
rect 3222 960 3228 961
rect 3222 956 3223 960
rect 3227 956 3228 960
rect 3222 955 3228 956
rect 3366 960 3372 961
rect 3366 956 3367 960
rect 3371 956 3372 960
rect 3462 959 3463 963
rect 3467 959 3468 963
rect 3462 958 3468 959
rect 3366 955 3372 956
rect 2312 927 2314 955
rect 2408 927 2410 955
rect 2512 927 2514 955
rect 2624 927 2626 955
rect 2752 927 2754 955
rect 2896 927 2898 955
rect 3056 927 3058 955
rect 3224 927 3226 955
rect 3368 927 3370 955
rect 3464 927 3466 958
rect 1807 926 1811 927
rect 1807 921 1811 922
rect 1831 926 1835 927
rect 1831 921 1835 922
rect 1983 926 1987 927
rect 1983 921 1987 922
rect 2151 926 2155 927
rect 2151 921 2155 922
rect 2311 926 2315 927
rect 2311 921 2315 922
rect 2327 926 2331 927
rect 2327 921 2331 922
rect 2407 926 2411 927
rect 2407 921 2411 922
rect 2511 926 2515 927
rect 2511 921 2515 922
rect 2519 926 2523 927
rect 2519 921 2523 922
rect 2623 926 2627 927
rect 2623 921 2627 922
rect 2719 926 2723 927
rect 2719 921 2723 922
rect 2751 926 2755 927
rect 2751 921 2755 922
rect 2895 926 2899 927
rect 2895 921 2899 922
rect 2935 926 2939 927
rect 2935 921 2939 922
rect 3055 926 3059 927
rect 3055 921 3059 922
rect 3159 926 3163 927
rect 3159 921 3163 922
rect 3223 926 3227 927
rect 3223 921 3227 922
rect 3367 926 3371 927
rect 3367 921 3371 922
rect 3463 926 3467 927
rect 3463 921 3467 922
rect 111 914 115 915
rect 111 909 115 910
rect 471 914 475 915
rect 471 909 475 910
rect 567 914 571 915
rect 567 909 571 910
rect 607 914 611 915
rect 607 909 611 910
rect 671 914 675 915
rect 671 909 675 910
rect 695 914 699 915
rect 695 909 699 910
rect 783 914 787 915
rect 783 909 787 910
rect 791 914 795 915
rect 791 909 795 910
rect 887 914 891 915
rect 887 909 891 910
rect 895 914 899 915
rect 895 909 899 910
rect 991 914 995 915
rect 991 909 995 910
rect 999 914 1003 915
rect 999 909 1003 910
rect 1095 914 1099 915
rect 1095 909 1099 910
rect 1111 914 1115 915
rect 1111 909 1115 910
rect 1199 914 1203 915
rect 1199 909 1203 910
rect 1223 914 1227 915
rect 1223 909 1227 910
rect 1295 914 1299 915
rect 1295 909 1299 910
rect 1343 914 1347 915
rect 1343 909 1347 910
rect 1391 914 1395 915
rect 1391 909 1395 910
rect 1463 914 1467 915
rect 1463 909 1467 910
rect 1487 914 1491 915
rect 1487 909 1491 910
rect 1583 914 1587 915
rect 1583 909 1587 910
rect 1671 914 1675 915
rect 1671 909 1675 910
rect 1767 914 1771 915
rect 1767 909 1771 910
rect 112 890 114 909
rect 608 893 610 909
rect 696 893 698 909
rect 792 893 794 909
rect 896 893 898 909
rect 1000 893 1002 909
rect 1112 893 1114 909
rect 1224 893 1226 909
rect 1344 893 1346 909
rect 1464 893 1466 909
rect 1584 893 1586 909
rect 606 892 612 893
rect 110 889 116 890
rect 110 885 111 889
rect 115 885 116 889
rect 606 888 607 892
rect 611 888 612 892
rect 606 887 612 888
rect 694 892 700 893
rect 694 888 695 892
rect 699 888 700 892
rect 694 887 700 888
rect 790 892 796 893
rect 790 888 791 892
rect 795 888 796 892
rect 790 887 796 888
rect 894 892 900 893
rect 894 888 895 892
rect 899 888 900 892
rect 894 887 900 888
rect 998 892 1004 893
rect 998 888 999 892
rect 1003 888 1004 892
rect 998 887 1004 888
rect 1110 892 1116 893
rect 1110 888 1111 892
rect 1115 888 1116 892
rect 1110 887 1116 888
rect 1222 892 1228 893
rect 1222 888 1223 892
rect 1227 888 1228 892
rect 1222 887 1228 888
rect 1342 892 1348 893
rect 1342 888 1343 892
rect 1347 888 1348 892
rect 1342 887 1348 888
rect 1462 892 1468 893
rect 1462 888 1463 892
rect 1467 888 1468 892
rect 1462 887 1468 888
rect 1582 892 1588 893
rect 1582 888 1583 892
rect 1587 888 1588 892
rect 1768 890 1770 909
rect 1808 902 1810 921
rect 1832 905 1834 921
rect 1984 905 1986 921
rect 2152 905 2154 921
rect 2328 905 2330 921
rect 2520 905 2522 921
rect 2720 905 2722 921
rect 2936 905 2938 921
rect 3160 905 3162 921
rect 3368 905 3370 921
rect 1830 904 1836 905
rect 1806 901 1812 902
rect 1806 897 1807 901
rect 1811 897 1812 901
rect 1830 900 1831 904
rect 1835 900 1836 904
rect 1830 899 1836 900
rect 1982 904 1988 905
rect 1982 900 1983 904
rect 1987 900 1988 904
rect 1982 899 1988 900
rect 2150 904 2156 905
rect 2150 900 2151 904
rect 2155 900 2156 904
rect 2150 899 2156 900
rect 2326 904 2332 905
rect 2326 900 2327 904
rect 2331 900 2332 904
rect 2326 899 2332 900
rect 2518 904 2524 905
rect 2518 900 2519 904
rect 2523 900 2524 904
rect 2518 899 2524 900
rect 2718 904 2724 905
rect 2718 900 2719 904
rect 2723 900 2724 904
rect 2718 899 2724 900
rect 2934 904 2940 905
rect 2934 900 2935 904
rect 2939 900 2940 904
rect 2934 899 2940 900
rect 3158 904 3164 905
rect 3158 900 3159 904
rect 3163 900 3164 904
rect 3158 899 3164 900
rect 3366 904 3372 905
rect 3366 900 3367 904
rect 3371 900 3372 904
rect 3464 902 3466 921
rect 3366 899 3372 900
rect 3462 901 3468 902
rect 1806 896 1812 897
rect 3462 897 3463 901
rect 3467 897 3468 901
rect 3462 896 3468 897
rect 1582 887 1588 888
rect 1766 889 1772 890
rect 110 884 116 885
rect 1766 885 1767 889
rect 1771 885 1772 889
rect 1830 885 1836 886
rect 1766 884 1772 885
rect 1806 884 1812 885
rect 1806 880 1807 884
rect 1811 880 1812 884
rect 1830 881 1831 885
rect 1835 881 1836 885
rect 1830 880 1836 881
rect 1982 885 1988 886
rect 1982 881 1983 885
rect 1987 881 1988 885
rect 1982 880 1988 881
rect 2150 885 2156 886
rect 2150 881 2151 885
rect 2155 881 2156 885
rect 2150 880 2156 881
rect 2326 885 2332 886
rect 2326 881 2327 885
rect 2331 881 2332 885
rect 2326 880 2332 881
rect 2518 885 2524 886
rect 2518 881 2519 885
rect 2523 881 2524 885
rect 2518 880 2524 881
rect 2718 885 2724 886
rect 2718 881 2719 885
rect 2723 881 2724 885
rect 2718 880 2724 881
rect 2934 885 2940 886
rect 2934 881 2935 885
rect 2939 881 2940 885
rect 2934 880 2940 881
rect 3158 885 3164 886
rect 3158 881 3159 885
rect 3163 881 3164 885
rect 3158 880 3164 881
rect 3366 885 3372 886
rect 3366 881 3367 885
rect 3371 881 3372 885
rect 3366 880 3372 881
rect 3462 884 3468 885
rect 3462 880 3463 884
rect 3467 880 3468 884
rect 1806 879 1812 880
rect 606 873 612 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 606 869 607 873
rect 611 869 612 873
rect 606 868 612 869
rect 694 873 700 874
rect 694 869 695 873
rect 699 869 700 873
rect 694 868 700 869
rect 790 873 796 874
rect 790 869 791 873
rect 795 869 796 873
rect 790 868 796 869
rect 894 873 900 874
rect 894 869 895 873
rect 899 869 900 873
rect 894 868 900 869
rect 998 873 1004 874
rect 998 869 999 873
rect 1003 869 1004 873
rect 998 868 1004 869
rect 1110 873 1116 874
rect 1110 869 1111 873
rect 1115 869 1116 873
rect 1110 868 1116 869
rect 1222 873 1228 874
rect 1222 869 1223 873
rect 1227 869 1228 873
rect 1222 868 1228 869
rect 1342 873 1348 874
rect 1342 869 1343 873
rect 1347 869 1348 873
rect 1342 868 1348 869
rect 1462 873 1468 874
rect 1462 869 1463 873
rect 1467 869 1468 873
rect 1462 868 1468 869
rect 1582 873 1588 874
rect 1582 869 1583 873
rect 1587 869 1588 873
rect 1582 868 1588 869
rect 1766 872 1772 873
rect 1766 868 1767 872
rect 1771 868 1772 872
rect 110 867 116 868
rect 112 847 114 867
rect 608 847 610 868
rect 696 847 698 868
rect 792 847 794 868
rect 896 847 898 868
rect 1000 847 1002 868
rect 1112 847 1114 868
rect 1224 847 1226 868
rect 1344 847 1346 868
rect 1464 847 1466 868
rect 1584 847 1586 868
rect 1766 867 1772 868
rect 1768 847 1770 867
rect 1808 859 1810 879
rect 1832 859 1834 880
rect 1984 859 1986 880
rect 2152 859 2154 880
rect 2328 859 2330 880
rect 2520 859 2522 880
rect 2720 859 2722 880
rect 2936 859 2938 880
rect 3160 859 3162 880
rect 3368 859 3370 880
rect 3462 879 3468 880
rect 3464 859 3466 879
rect 1807 858 1811 859
rect 1807 853 1811 854
rect 1831 858 1835 859
rect 1831 853 1835 854
rect 1959 858 1963 859
rect 1959 853 1963 854
rect 1983 858 1987 859
rect 1983 853 1987 854
rect 2087 858 2091 859
rect 2087 853 2091 854
rect 2151 858 2155 859
rect 2151 853 2155 854
rect 2207 858 2211 859
rect 2207 853 2211 854
rect 2327 858 2331 859
rect 2327 853 2331 854
rect 2463 858 2467 859
rect 2463 853 2467 854
rect 2519 858 2523 859
rect 2519 853 2523 854
rect 2615 858 2619 859
rect 2615 853 2619 854
rect 2719 858 2723 859
rect 2719 853 2723 854
rect 2791 858 2795 859
rect 2791 853 2795 854
rect 2935 858 2939 859
rect 2935 853 2939 854
rect 2983 858 2987 859
rect 2983 853 2987 854
rect 3159 858 3163 859
rect 3159 853 3163 854
rect 3183 858 3187 859
rect 3183 853 3187 854
rect 3367 858 3371 859
rect 3367 853 3371 854
rect 3463 858 3467 859
rect 3463 853 3467 854
rect 111 846 115 847
rect 111 841 115 842
rect 519 846 523 847
rect 519 841 523 842
rect 607 846 611 847
rect 607 841 611 842
rect 615 846 619 847
rect 615 841 619 842
rect 695 846 699 847
rect 695 841 699 842
rect 719 846 723 847
rect 719 841 723 842
rect 791 846 795 847
rect 791 841 795 842
rect 831 846 835 847
rect 831 841 835 842
rect 895 846 899 847
rect 895 841 899 842
rect 951 846 955 847
rect 951 841 955 842
rect 999 846 1003 847
rect 999 841 1003 842
rect 1071 846 1075 847
rect 1071 841 1075 842
rect 1111 846 1115 847
rect 1111 841 1115 842
rect 1191 846 1195 847
rect 1191 841 1195 842
rect 1223 846 1227 847
rect 1223 841 1227 842
rect 1311 846 1315 847
rect 1311 841 1315 842
rect 1343 846 1347 847
rect 1343 841 1347 842
rect 1431 846 1435 847
rect 1431 841 1435 842
rect 1463 846 1467 847
rect 1463 841 1467 842
rect 1559 846 1563 847
rect 1559 841 1563 842
rect 1583 846 1587 847
rect 1583 841 1587 842
rect 1767 846 1771 847
rect 1767 841 1771 842
rect 112 825 114 841
rect 110 824 116 825
rect 520 824 522 841
rect 616 824 618 841
rect 720 824 722 841
rect 832 824 834 841
rect 952 824 954 841
rect 1072 824 1074 841
rect 1192 824 1194 841
rect 1312 824 1314 841
rect 1432 824 1434 841
rect 1560 824 1562 841
rect 1768 825 1770 841
rect 1808 837 1810 853
rect 1806 836 1812 837
rect 1832 836 1834 853
rect 1960 836 1962 853
rect 2088 836 2090 853
rect 2208 836 2210 853
rect 2328 836 2330 853
rect 2464 836 2466 853
rect 2616 836 2618 853
rect 2792 836 2794 853
rect 2984 836 2986 853
rect 3184 836 3186 853
rect 3368 836 3370 853
rect 3464 837 3466 853
rect 3462 836 3468 837
rect 1806 832 1807 836
rect 1811 832 1812 836
rect 1806 831 1812 832
rect 1830 835 1836 836
rect 1830 831 1831 835
rect 1835 831 1836 835
rect 1830 830 1836 831
rect 1958 835 1964 836
rect 1958 831 1959 835
rect 1963 831 1964 835
rect 1958 830 1964 831
rect 2086 835 2092 836
rect 2086 831 2087 835
rect 2091 831 2092 835
rect 2086 830 2092 831
rect 2206 835 2212 836
rect 2206 831 2207 835
rect 2211 831 2212 835
rect 2206 830 2212 831
rect 2326 835 2332 836
rect 2326 831 2327 835
rect 2331 831 2332 835
rect 2326 830 2332 831
rect 2462 835 2468 836
rect 2462 831 2463 835
rect 2467 831 2468 835
rect 2462 830 2468 831
rect 2614 835 2620 836
rect 2614 831 2615 835
rect 2619 831 2620 835
rect 2614 830 2620 831
rect 2790 835 2796 836
rect 2790 831 2791 835
rect 2795 831 2796 835
rect 2790 830 2796 831
rect 2982 835 2988 836
rect 2982 831 2983 835
rect 2987 831 2988 835
rect 2982 830 2988 831
rect 3182 835 3188 836
rect 3182 831 3183 835
rect 3187 831 3188 835
rect 3182 830 3188 831
rect 3366 835 3372 836
rect 3366 831 3367 835
rect 3371 831 3372 835
rect 3462 832 3463 836
rect 3467 832 3468 836
rect 3462 831 3468 832
rect 3366 830 3372 831
rect 1766 824 1772 825
rect 110 820 111 824
rect 115 820 116 824
rect 110 819 116 820
rect 518 823 524 824
rect 518 819 519 823
rect 523 819 524 823
rect 518 818 524 819
rect 614 823 620 824
rect 614 819 615 823
rect 619 819 620 823
rect 614 818 620 819
rect 718 823 724 824
rect 718 819 719 823
rect 723 819 724 823
rect 718 818 724 819
rect 830 823 836 824
rect 830 819 831 823
rect 835 819 836 823
rect 830 818 836 819
rect 950 823 956 824
rect 950 819 951 823
rect 955 819 956 823
rect 950 818 956 819
rect 1070 823 1076 824
rect 1070 819 1071 823
rect 1075 819 1076 823
rect 1070 818 1076 819
rect 1190 823 1196 824
rect 1190 819 1191 823
rect 1195 819 1196 823
rect 1190 818 1196 819
rect 1310 823 1316 824
rect 1310 819 1311 823
rect 1315 819 1316 823
rect 1310 818 1316 819
rect 1430 823 1436 824
rect 1430 819 1431 823
rect 1435 819 1436 823
rect 1430 818 1436 819
rect 1558 823 1564 824
rect 1558 819 1559 823
rect 1563 819 1564 823
rect 1766 820 1767 824
rect 1771 820 1772 824
rect 1766 819 1772 820
rect 1806 819 1812 820
rect 1558 818 1564 819
rect 1806 815 1807 819
rect 1811 815 1812 819
rect 3462 819 3468 820
rect 1806 814 1812 815
rect 1830 816 1836 817
rect 110 807 116 808
rect 110 803 111 807
rect 115 803 116 807
rect 1766 807 1772 808
rect 110 802 116 803
rect 518 804 524 805
rect 112 779 114 802
rect 518 800 519 804
rect 523 800 524 804
rect 518 799 524 800
rect 614 804 620 805
rect 614 800 615 804
rect 619 800 620 804
rect 614 799 620 800
rect 718 804 724 805
rect 718 800 719 804
rect 723 800 724 804
rect 718 799 724 800
rect 830 804 836 805
rect 830 800 831 804
rect 835 800 836 804
rect 830 799 836 800
rect 950 804 956 805
rect 950 800 951 804
rect 955 800 956 804
rect 950 799 956 800
rect 1070 804 1076 805
rect 1070 800 1071 804
rect 1075 800 1076 804
rect 1070 799 1076 800
rect 1190 804 1196 805
rect 1190 800 1191 804
rect 1195 800 1196 804
rect 1190 799 1196 800
rect 1310 804 1316 805
rect 1310 800 1311 804
rect 1315 800 1316 804
rect 1310 799 1316 800
rect 1430 804 1436 805
rect 1430 800 1431 804
rect 1435 800 1436 804
rect 1430 799 1436 800
rect 1558 804 1564 805
rect 1558 800 1559 804
rect 1563 800 1564 804
rect 1766 803 1767 807
rect 1771 803 1772 807
rect 1766 802 1772 803
rect 1558 799 1564 800
rect 520 779 522 799
rect 616 779 618 799
rect 720 779 722 799
rect 832 779 834 799
rect 952 779 954 799
rect 1072 779 1074 799
rect 1192 779 1194 799
rect 1312 779 1314 799
rect 1432 779 1434 799
rect 1560 779 1562 799
rect 1768 779 1770 802
rect 1808 791 1810 814
rect 1830 812 1831 816
rect 1835 812 1836 816
rect 1830 811 1836 812
rect 1958 816 1964 817
rect 1958 812 1959 816
rect 1963 812 1964 816
rect 1958 811 1964 812
rect 2086 816 2092 817
rect 2086 812 2087 816
rect 2091 812 2092 816
rect 2086 811 2092 812
rect 2206 816 2212 817
rect 2206 812 2207 816
rect 2211 812 2212 816
rect 2206 811 2212 812
rect 2326 816 2332 817
rect 2326 812 2327 816
rect 2331 812 2332 816
rect 2326 811 2332 812
rect 2462 816 2468 817
rect 2462 812 2463 816
rect 2467 812 2468 816
rect 2462 811 2468 812
rect 2614 816 2620 817
rect 2614 812 2615 816
rect 2619 812 2620 816
rect 2614 811 2620 812
rect 2790 816 2796 817
rect 2790 812 2791 816
rect 2795 812 2796 816
rect 2790 811 2796 812
rect 2982 816 2988 817
rect 2982 812 2983 816
rect 2987 812 2988 816
rect 2982 811 2988 812
rect 3182 816 3188 817
rect 3182 812 3183 816
rect 3187 812 3188 816
rect 3182 811 3188 812
rect 3366 816 3372 817
rect 3366 812 3367 816
rect 3371 812 3372 816
rect 3462 815 3463 819
rect 3467 815 3468 819
rect 3462 814 3468 815
rect 3366 811 3372 812
rect 1832 791 1834 811
rect 1960 791 1962 811
rect 2088 791 2090 811
rect 2208 791 2210 811
rect 2328 791 2330 811
rect 2464 791 2466 811
rect 2616 791 2618 811
rect 2792 791 2794 811
rect 2984 791 2986 811
rect 3184 791 3186 811
rect 3368 791 3370 811
rect 3464 791 3466 814
rect 1807 790 1811 791
rect 1807 785 1811 786
rect 1831 790 1835 791
rect 1831 785 1835 786
rect 1879 790 1883 791
rect 1879 785 1883 786
rect 1959 790 1963 791
rect 1959 785 1963 786
rect 2015 790 2019 791
rect 2015 785 2019 786
rect 2087 790 2091 791
rect 2087 785 2091 786
rect 2151 790 2155 791
rect 2151 785 2155 786
rect 2207 790 2211 791
rect 2207 785 2211 786
rect 2287 790 2291 791
rect 2287 785 2291 786
rect 2327 790 2331 791
rect 2327 785 2331 786
rect 2423 790 2427 791
rect 2423 785 2427 786
rect 2463 790 2467 791
rect 2463 785 2467 786
rect 2559 790 2563 791
rect 2559 785 2563 786
rect 2615 790 2619 791
rect 2615 785 2619 786
rect 2711 790 2715 791
rect 2711 785 2715 786
rect 2791 790 2795 791
rect 2791 785 2795 786
rect 2871 790 2875 791
rect 2871 785 2875 786
rect 2983 790 2987 791
rect 2983 785 2987 786
rect 3039 790 3043 791
rect 3039 785 3043 786
rect 3183 790 3187 791
rect 3183 785 3187 786
rect 3215 790 3219 791
rect 3215 785 3219 786
rect 3367 790 3371 791
rect 3367 785 3371 786
rect 3463 790 3467 791
rect 3463 785 3467 786
rect 111 778 115 779
rect 111 773 115 774
rect 383 778 387 779
rect 383 773 387 774
rect 471 778 475 779
rect 471 773 475 774
rect 519 778 523 779
rect 519 773 523 774
rect 575 778 579 779
rect 575 773 579 774
rect 615 778 619 779
rect 615 773 619 774
rect 679 778 683 779
rect 679 773 683 774
rect 719 778 723 779
rect 719 773 723 774
rect 791 778 795 779
rect 791 773 795 774
rect 831 778 835 779
rect 831 773 835 774
rect 911 778 915 779
rect 911 773 915 774
rect 951 778 955 779
rect 951 773 955 774
rect 1031 778 1035 779
rect 1031 773 1035 774
rect 1071 778 1075 779
rect 1071 773 1075 774
rect 1159 778 1163 779
rect 1159 773 1163 774
rect 1191 778 1195 779
rect 1191 773 1195 774
rect 1287 778 1291 779
rect 1287 773 1291 774
rect 1311 778 1315 779
rect 1311 773 1315 774
rect 1415 778 1419 779
rect 1415 773 1419 774
rect 1431 778 1435 779
rect 1431 773 1435 774
rect 1559 778 1563 779
rect 1559 773 1563 774
rect 1767 778 1771 779
rect 1767 773 1771 774
rect 112 754 114 773
rect 384 757 386 773
rect 472 757 474 773
rect 576 757 578 773
rect 680 757 682 773
rect 792 757 794 773
rect 912 757 914 773
rect 1032 757 1034 773
rect 1160 757 1162 773
rect 1288 757 1290 773
rect 1416 757 1418 773
rect 382 756 388 757
rect 110 753 116 754
rect 110 749 111 753
rect 115 749 116 753
rect 382 752 383 756
rect 387 752 388 756
rect 382 751 388 752
rect 470 756 476 757
rect 470 752 471 756
rect 475 752 476 756
rect 470 751 476 752
rect 574 756 580 757
rect 574 752 575 756
rect 579 752 580 756
rect 574 751 580 752
rect 678 756 684 757
rect 678 752 679 756
rect 683 752 684 756
rect 678 751 684 752
rect 790 756 796 757
rect 790 752 791 756
rect 795 752 796 756
rect 790 751 796 752
rect 910 756 916 757
rect 910 752 911 756
rect 915 752 916 756
rect 910 751 916 752
rect 1030 756 1036 757
rect 1030 752 1031 756
rect 1035 752 1036 756
rect 1030 751 1036 752
rect 1158 756 1164 757
rect 1158 752 1159 756
rect 1163 752 1164 756
rect 1158 751 1164 752
rect 1286 756 1292 757
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1414 756 1420 757
rect 1414 752 1415 756
rect 1419 752 1420 756
rect 1768 754 1770 773
rect 1808 766 1810 785
rect 1880 769 1882 785
rect 2016 769 2018 785
rect 2152 769 2154 785
rect 2288 769 2290 785
rect 2424 769 2426 785
rect 2560 769 2562 785
rect 2712 769 2714 785
rect 2872 769 2874 785
rect 3040 769 3042 785
rect 3216 769 3218 785
rect 3368 769 3370 785
rect 1878 768 1884 769
rect 1806 765 1812 766
rect 1806 761 1807 765
rect 1811 761 1812 765
rect 1878 764 1879 768
rect 1883 764 1884 768
rect 1878 763 1884 764
rect 2014 768 2020 769
rect 2014 764 2015 768
rect 2019 764 2020 768
rect 2014 763 2020 764
rect 2150 768 2156 769
rect 2150 764 2151 768
rect 2155 764 2156 768
rect 2150 763 2156 764
rect 2286 768 2292 769
rect 2286 764 2287 768
rect 2291 764 2292 768
rect 2286 763 2292 764
rect 2422 768 2428 769
rect 2422 764 2423 768
rect 2427 764 2428 768
rect 2422 763 2428 764
rect 2558 768 2564 769
rect 2558 764 2559 768
rect 2563 764 2564 768
rect 2558 763 2564 764
rect 2710 768 2716 769
rect 2710 764 2711 768
rect 2715 764 2716 768
rect 2710 763 2716 764
rect 2870 768 2876 769
rect 2870 764 2871 768
rect 2875 764 2876 768
rect 2870 763 2876 764
rect 3038 768 3044 769
rect 3038 764 3039 768
rect 3043 764 3044 768
rect 3038 763 3044 764
rect 3214 768 3220 769
rect 3214 764 3215 768
rect 3219 764 3220 768
rect 3214 763 3220 764
rect 3366 768 3372 769
rect 3366 764 3367 768
rect 3371 764 3372 768
rect 3464 766 3466 785
rect 3366 763 3372 764
rect 3462 765 3468 766
rect 1806 760 1812 761
rect 3462 761 3463 765
rect 3467 761 3468 765
rect 3462 760 3468 761
rect 1414 751 1420 752
rect 1766 753 1772 754
rect 110 748 116 749
rect 1766 749 1767 753
rect 1771 749 1772 753
rect 1878 749 1884 750
rect 1766 748 1772 749
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1878 745 1879 749
rect 1883 745 1884 749
rect 1878 744 1884 745
rect 2014 749 2020 750
rect 2014 745 2015 749
rect 2019 745 2020 749
rect 2014 744 2020 745
rect 2150 749 2156 750
rect 2150 745 2151 749
rect 2155 745 2156 749
rect 2150 744 2156 745
rect 2286 749 2292 750
rect 2286 745 2287 749
rect 2291 745 2292 749
rect 2286 744 2292 745
rect 2422 749 2428 750
rect 2422 745 2423 749
rect 2427 745 2428 749
rect 2422 744 2428 745
rect 2558 749 2564 750
rect 2558 745 2559 749
rect 2563 745 2564 749
rect 2558 744 2564 745
rect 2710 749 2716 750
rect 2710 745 2711 749
rect 2715 745 2716 749
rect 2710 744 2716 745
rect 2870 749 2876 750
rect 2870 745 2871 749
rect 2875 745 2876 749
rect 2870 744 2876 745
rect 3038 749 3044 750
rect 3038 745 3039 749
rect 3043 745 3044 749
rect 3038 744 3044 745
rect 3214 749 3220 750
rect 3214 745 3215 749
rect 3219 745 3220 749
rect 3214 744 3220 745
rect 3366 749 3372 750
rect 3366 745 3367 749
rect 3371 745 3372 749
rect 3366 744 3372 745
rect 3462 748 3468 749
rect 3462 744 3463 748
rect 3467 744 3468 748
rect 1806 743 1812 744
rect 382 737 388 738
rect 110 736 116 737
rect 110 732 111 736
rect 115 732 116 736
rect 382 733 383 737
rect 387 733 388 737
rect 382 732 388 733
rect 470 737 476 738
rect 470 733 471 737
rect 475 733 476 737
rect 470 732 476 733
rect 574 737 580 738
rect 574 733 575 737
rect 579 733 580 737
rect 574 732 580 733
rect 678 737 684 738
rect 678 733 679 737
rect 683 733 684 737
rect 678 732 684 733
rect 790 737 796 738
rect 790 733 791 737
rect 795 733 796 737
rect 790 732 796 733
rect 910 737 916 738
rect 910 733 911 737
rect 915 733 916 737
rect 910 732 916 733
rect 1030 737 1036 738
rect 1030 733 1031 737
rect 1035 733 1036 737
rect 1030 732 1036 733
rect 1158 737 1164 738
rect 1158 733 1159 737
rect 1163 733 1164 737
rect 1158 732 1164 733
rect 1286 737 1292 738
rect 1286 733 1287 737
rect 1291 733 1292 737
rect 1286 732 1292 733
rect 1414 737 1420 738
rect 1414 733 1415 737
rect 1419 733 1420 737
rect 1414 732 1420 733
rect 1766 736 1772 737
rect 1766 732 1767 736
rect 1771 732 1772 736
rect 110 731 116 732
rect 112 707 114 731
rect 384 707 386 732
rect 472 707 474 732
rect 576 707 578 732
rect 680 707 682 732
rect 792 707 794 732
rect 912 707 914 732
rect 1032 707 1034 732
rect 1160 707 1162 732
rect 1288 707 1290 732
rect 1416 707 1418 732
rect 1766 731 1772 732
rect 1768 707 1770 731
rect 1808 723 1810 743
rect 1880 723 1882 744
rect 2016 723 2018 744
rect 2152 723 2154 744
rect 2288 723 2290 744
rect 2424 723 2426 744
rect 2560 723 2562 744
rect 2712 723 2714 744
rect 2872 723 2874 744
rect 3040 723 3042 744
rect 3216 723 3218 744
rect 3368 723 3370 744
rect 3462 743 3468 744
rect 3464 723 3466 743
rect 1807 722 1811 723
rect 1807 717 1811 718
rect 1831 722 1835 723
rect 1831 717 1835 718
rect 1879 722 1883 723
rect 1879 717 1883 718
rect 1951 722 1955 723
rect 1951 717 1955 718
rect 2015 722 2019 723
rect 2015 717 2019 718
rect 2103 722 2107 723
rect 2103 717 2107 718
rect 2151 722 2155 723
rect 2151 717 2155 718
rect 2263 722 2267 723
rect 2263 717 2267 718
rect 2287 722 2291 723
rect 2287 717 2291 718
rect 2415 722 2419 723
rect 2415 717 2419 718
rect 2423 722 2427 723
rect 2423 717 2427 718
rect 2559 722 2563 723
rect 2559 717 2563 718
rect 2567 722 2571 723
rect 2567 717 2571 718
rect 2711 722 2715 723
rect 2711 717 2715 718
rect 2719 722 2723 723
rect 2719 717 2723 718
rect 2871 722 2875 723
rect 2871 717 2875 718
rect 2879 722 2883 723
rect 2879 717 2883 718
rect 3039 722 3043 723
rect 3039 717 3043 718
rect 3199 722 3203 723
rect 3199 717 3203 718
rect 3215 722 3219 723
rect 3215 717 3219 718
rect 3367 722 3371 723
rect 3367 717 3371 718
rect 3463 722 3467 723
rect 3463 717 3467 718
rect 111 706 115 707
rect 111 701 115 702
rect 247 706 251 707
rect 247 701 251 702
rect 343 706 347 707
rect 343 701 347 702
rect 383 706 387 707
rect 383 701 387 702
rect 455 706 459 707
rect 455 701 459 702
rect 471 706 475 707
rect 471 701 475 702
rect 567 706 571 707
rect 567 701 571 702
rect 575 706 579 707
rect 575 701 579 702
rect 679 706 683 707
rect 679 701 683 702
rect 695 706 699 707
rect 695 701 699 702
rect 791 706 795 707
rect 791 701 795 702
rect 831 706 835 707
rect 831 701 835 702
rect 911 706 915 707
rect 911 701 915 702
rect 983 706 987 707
rect 983 701 987 702
rect 1031 706 1035 707
rect 1031 701 1035 702
rect 1151 706 1155 707
rect 1151 701 1155 702
rect 1159 706 1163 707
rect 1159 701 1163 702
rect 1287 706 1291 707
rect 1287 701 1291 702
rect 1327 706 1331 707
rect 1327 701 1331 702
rect 1415 706 1419 707
rect 1415 701 1419 702
rect 1511 706 1515 707
rect 1511 701 1515 702
rect 1671 706 1675 707
rect 1671 701 1675 702
rect 1767 706 1771 707
rect 1767 701 1771 702
rect 1808 701 1810 717
rect 112 685 114 701
rect 110 684 116 685
rect 248 684 250 701
rect 344 684 346 701
rect 456 684 458 701
rect 568 684 570 701
rect 696 684 698 701
rect 832 684 834 701
rect 984 684 986 701
rect 1152 684 1154 701
rect 1328 684 1330 701
rect 1512 684 1514 701
rect 1672 684 1674 701
rect 1768 685 1770 701
rect 1806 700 1812 701
rect 1832 700 1834 717
rect 1952 700 1954 717
rect 2104 700 2106 717
rect 2264 700 2266 717
rect 2416 700 2418 717
rect 2568 700 2570 717
rect 2720 700 2722 717
rect 2880 700 2882 717
rect 3040 700 3042 717
rect 3200 700 3202 717
rect 3464 701 3466 717
rect 3462 700 3468 701
rect 1806 696 1807 700
rect 1811 696 1812 700
rect 1806 695 1812 696
rect 1830 699 1836 700
rect 1830 695 1831 699
rect 1835 695 1836 699
rect 1830 694 1836 695
rect 1950 699 1956 700
rect 1950 695 1951 699
rect 1955 695 1956 699
rect 1950 694 1956 695
rect 2102 699 2108 700
rect 2102 695 2103 699
rect 2107 695 2108 699
rect 2102 694 2108 695
rect 2262 699 2268 700
rect 2262 695 2263 699
rect 2267 695 2268 699
rect 2262 694 2268 695
rect 2414 699 2420 700
rect 2414 695 2415 699
rect 2419 695 2420 699
rect 2414 694 2420 695
rect 2566 699 2572 700
rect 2566 695 2567 699
rect 2571 695 2572 699
rect 2566 694 2572 695
rect 2718 699 2724 700
rect 2718 695 2719 699
rect 2723 695 2724 699
rect 2718 694 2724 695
rect 2878 699 2884 700
rect 2878 695 2879 699
rect 2883 695 2884 699
rect 2878 694 2884 695
rect 3038 699 3044 700
rect 3038 695 3039 699
rect 3043 695 3044 699
rect 3038 694 3044 695
rect 3198 699 3204 700
rect 3198 695 3199 699
rect 3203 695 3204 699
rect 3462 696 3463 700
rect 3467 696 3468 700
rect 3462 695 3468 696
rect 3198 694 3204 695
rect 1766 684 1772 685
rect 110 680 111 684
rect 115 680 116 684
rect 110 679 116 680
rect 246 683 252 684
rect 246 679 247 683
rect 251 679 252 683
rect 246 678 252 679
rect 342 683 348 684
rect 342 679 343 683
rect 347 679 348 683
rect 342 678 348 679
rect 454 683 460 684
rect 454 679 455 683
rect 459 679 460 683
rect 454 678 460 679
rect 566 683 572 684
rect 566 679 567 683
rect 571 679 572 683
rect 566 678 572 679
rect 694 683 700 684
rect 694 679 695 683
rect 699 679 700 683
rect 694 678 700 679
rect 830 683 836 684
rect 830 679 831 683
rect 835 679 836 683
rect 830 678 836 679
rect 982 683 988 684
rect 982 679 983 683
rect 987 679 988 683
rect 982 678 988 679
rect 1150 683 1156 684
rect 1150 679 1151 683
rect 1155 679 1156 683
rect 1150 678 1156 679
rect 1326 683 1332 684
rect 1326 679 1327 683
rect 1331 679 1332 683
rect 1326 678 1332 679
rect 1510 683 1516 684
rect 1510 679 1511 683
rect 1515 679 1516 683
rect 1510 678 1516 679
rect 1670 683 1676 684
rect 1670 679 1671 683
rect 1675 679 1676 683
rect 1766 680 1767 684
rect 1771 680 1772 684
rect 1766 679 1772 680
rect 1806 683 1812 684
rect 1806 679 1807 683
rect 1811 679 1812 683
rect 3462 683 3468 684
rect 1670 678 1676 679
rect 1806 678 1812 679
rect 1830 680 1836 681
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 1766 667 1772 668
rect 110 662 116 663
rect 246 664 252 665
rect 112 639 114 662
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 342 664 348 665
rect 342 660 343 664
rect 347 660 348 664
rect 342 659 348 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 566 664 572 665
rect 566 660 567 664
rect 571 660 572 664
rect 566 659 572 660
rect 694 664 700 665
rect 694 660 695 664
rect 699 660 700 664
rect 694 659 700 660
rect 830 664 836 665
rect 830 660 831 664
rect 835 660 836 664
rect 830 659 836 660
rect 982 664 988 665
rect 982 660 983 664
rect 987 660 988 664
rect 982 659 988 660
rect 1150 664 1156 665
rect 1150 660 1151 664
rect 1155 660 1156 664
rect 1150 659 1156 660
rect 1326 664 1332 665
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1510 664 1516 665
rect 1510 660 1511 664
rect 1515 660 1516 664
rect 1510 659 1516 660
rect 1670 664 1676 665
rect 1670 660 1671 664
rect 1675 660 1676 664
rect 1766 663 1767 667
rect 1771 663 1772 667
rect 1766 662 1772 663
rect 1670 659 1676 660
rect 248 639 250 659
rect 344 639 346 659
rect 456 639 458 659
rect 568 639 570 659
rect 696 639 698 659
rect 832 639 834 659
rect 984 639 986 659
rect 1152 639 1154 659
rect 1328 639 1330 659
rect 1512 639 1514 659
rect 1672 639 1674 659
rect 1768 639 1770 662
rect 1808 659 1810 678
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1950 680 1956 681
rect 1950 676 1951 680
rect 1955 676 1956 680
rect 1950 675 1956 676
rect 2102 680 2108 681
rect 2102 676 2103 680
rect 2107 676 2108 680
rect 2102 675 2108 676
rect 2262 680 2268 681
rect 2262 676 2263 680
rect 2267 676 2268 680
rect 2262 675 2268 676
rect 2414 680 2420 681
rect 2414 676 2415 680
rect 2419 676 2420 680
rect 2414 675 2420 676
rect 2566 680 2572 681
rect 2566 676 2567 680
rect 2571 676 2572 680
rect 2566 675 2572 676
rect 2718 680 2724 681
rect 2718 676 2719 680
rect 2723 676 2724 680
rect 2718 675 2724 676
rect 2878 680 2884 681
rect 2878 676 2879 680
rect 2883 676 2884 680
rect 2878 675 2884 676
rect 3038 680 3044 681
rect 3038 676 3039 680
rect 3043 676 3044 680
rect 3038 675 3044 676
rect 3198 680 3204 681
rect 3198 676 3199 680
rect 3203 676 3204 680
rect 3462 679 3463 683
rect 3467 679 3468 683
rect 3462 678 3468 679
rect 3198 675 3204 676
rect 1832 659 1834 675
rect 1952 659 1954 675
rect 2104 659 2106 675
rect 2264 659 2266 675
rect 2416 659 2418 675
rect 2568 659 2570 675
rect 2720 659 2722 675
rect 2880 659 2882 675
rect 3040 659 3042 675
rect 3200 659 3202 675
rect 3464 659 3466 678
rect 1807 658 1811 659
rect 1807 653 1811 654
rect 1831 658 1835 659
rect 1831 653 1835 654
rect 1951 658 1955 659
rect 1951 653 1955 654
rect 1975 658 1979 659
rect 1975 653 1979 654
rect 2103 658 2107 659
rect 2103 653 2107 654
rect 2239 658 2243 659
rect 2239 653 2243 654
rect 2263 658 2267 659
rect 2263 653 2267 654
rect 2415 658 2419 659
rect 2415 653 2419 654
rect 2479 658 2483 659
rect 2479 653 2483 654
rect 2567 658 2571 659
rect 2567 653 2571 654
rect 2687 658 2691 659
rect 2687 653 2691 654
rect 2719 658 2723 659
rect 2719 653 2723 654
rect 2879 658 2883 659
rect 2879 653 2883 654
rect 3039 658 3043 659
rect 3039 653 3043 654
rect 3055 658 3059 659
rect 3055 653 3059 654
rect 3199 658 3203 659
rect 3199 653 3203 654
rect 3223 658 3227 659
rect 3223 653 3227 654
rect 3367 658 3371 659
rect 3367 653 3371 654
rect 3463 658 3467 659
rect 3463 653 3467 654
rect 111 638 115 639
rect 111 633 115 634
rect 135 638 139 639
rect 135 633 139 634
rect 231 638 235 639
rect 231 633 235 634
rect 247 638 251 639
rect 247 633 251 634
rect 343 638 347 639
rect 343 633 347 634
rect 359 638 363 639
rect 359 633 363 634
rect 455 638 459 639
rect 455 633 459 634
rect 487 638 491 639
rect 487 633 491 634
rect 567 638 571 639
rect 567 633 571 634
rect 623 638 627 639
rect 623 633 627 634
rect 695 638 699 639
rect 695 633 699 634
rect 767 638 771 639
rect 767 633 771 634
rect 831 638 835 639
rect 831 633 835 634
rect 911 638 915 639
rect 911 633 915 634
rect 983 638 987 639
rect 983 633 987 634
rect 1055 638 1059 639
rect 1055 633 1059 634
rect 1151 638 1155 639
rect 1151 633 1155 634
rect 1207 638 1211 639
rect 1207 633 1211 634
rect 1327 638 1331 639
rect 1327 633 1331 634
rect 1367 638 1371 639
rect 1367 633 1371 634
rect 1511 638 1515 639
rect 1511 633 1515 634
rect 1527 638 1531 639
rect 1527 633 1531 634
rect 1671 638 1675 639
rect 1671 633 1675 634
rect 1767 638 1771 639
rect 1808 634 1810 653
rect 1976 637 1978 653
rect 2240 637 2242 653
rect 2480 637 2482 653
rect 2688 637 2690 653
rect 2880 637 2882 653
rect 3056 637 3058 653
rect 3224 637 3226 653
rect 3368 637 3370 653
rect 1974 636 1980 637
rect 1767 633 1771 634
rect 1806 633 1812 634
rect 112 614 114 633
rect 136 617 138 633
rect 232 617 234 633
rect 360 617 362 633
rect 488 617 490 633
rect 624 617 626 633
rect 768 617 770 633
rect 912 617 914 633
rect 1056 617 1058 633
rect 1208 617 1210 633
rect 1368 617 1370 633
rect 1528 617 1530 633
rect 1672 617 1674 633
rect 134 616 140 617
rect 110 613 116 614
rect 110 609 111 613
rect 115 609 116 613
rect 134 612 135 616
rect 139 612 140 616
rect 134 611 140 612
rect 230 616 236 617
rect 230 612 231 616
rect 235 612 236 616
rect 230 611 236 612
rect 358 616 364 617
rect 358 612 359 616
rect 363 612 364 616
rect 358 611 364 612
rect 486 616 492 617
rect 486 612 487 616
rect 491 612 492 616
rect 486 611 492 612
rect 622 616 628 617
rect 622 612 623 616
rect 627 612 628 616
rect 622 611 628 612
rect 766 616 772 617
rect 766 612 767 616
rect 771 612 772 616
rect 766 611 772 612
rect 910 616 916 617
rect 910 612 911 616
rect 915 612 916 616
rect 910 611 916 612
rect 1054 616 1060 617
rect 1054 612 1055 616
rect 1059 612 1060 616
rect 1054 611 1060 612
rect 1206 616 1212 617
rect 1206 612 1207 616
rect 1211 612 1212 616
rect 1206 611 1212 612
rect 1366 616 1372 617
rect 1366 612 1367 616
rect 1371 612 1372 616
rect 1366 611 1372 612
rect 1526 616 1532 617
rect 1526 612 1527 616
rect 1531 612 1532 616
rect 1526 611 1532 612
rect 1670 616 1676 617
rect 1670 612 1671 616
rect 1675 612 1676 616
rect 1768 614 1770 633
rect 1806 629 1807 633
rect 1811 629 1812 633
rect 1974 632 1975 636
rect 1979 632 1980 636
rect 1974 631 1980 632
rect 2238 636 2244 637
rect 2238 632 2239 636
rect 2243 632 2244 636
rect 2238 631 2244 632
rect 2478 636 2484 637
rect 2478 632 2479 636
rect 2483 632 2484 636
rect 2478 631 2484 632
rect 2686 636 2692 637
rect 2686 632 2687 636
rect 2691 632 2692 636
rect 2686 631 2692 632
rect 2878 636 2884 637
rect 2878 632 2879 636
rect 2883 632 2884 636
rect 2878 631 2884 632
rect 3054 636 3060 637
rect 3054 632 3055 636
rect 3059 632 3060 636
rect 3054 631 3060 632
rect 3222 636 3228 637
rect 3222 632 3223 636
rect 3227 632 3228 636
rect 3222 631 3228 632
rect 3366 636 3372 637
rect 3366 632 3367 636
rect 3371 632 3372 636
rect 3464 634 3466 653
rect 3366 631 3372 632
rect 3462 633 3468 634
rect 1806 628 1812 629
rect 3462 629 3463 633
rect 3467 629 3468 633
rect 3462 628 3468 629
rect 1974 617 1980 618
rect 1806 616 1812 617
rect 1670 611 1676 612
rect 1766 613 1772 614
rect 110 608 116 609
rect 1766 609 1767 613
rect 1771 609 1772 613
rect 1806 612 1807 616
rect 1811 612 1812 616
rect 1974 613 1975 617
rect 1979 613 1980 617
rect 1974 612 1980 613
rect 2238 617 2244 618
rect 2238 613 2239 617
rect 2243 613 2244 617
rect 2238 612 2244 613
rect 2478 617 2484 618
rect 2478 613 2479 617
rect 2483 613 2484 617
rect 2478 612 2484 613
rect 2686 617 2692 618
rect 2686 613 2687 617
rect 2691 613 2692 617
rect 2686 612 2692 613
rect 2878 617 2884 618
rect 2878 613 2879 617
rect 2883 613 2884 617
rect 2878 612 2884 613
rect 3054 617 3060 618
rect 3054 613 3055 617
rect 3059 613 3060 617
rect 3054 612 3060 613
rect 3222 617 3228 618
rect 3222 613 3223 617
rect 3227 613 3228 617
rect 3222 612 3228 613
rect 3366 617 3372 618
rect 3366 613 3367 617
rect 3371 613 3372 617
rect 3366 612 3372 613
rect 3462 616 3468 617
rect 3462 612 3463 616
rect 3467 612 3468 616
rect 1806 611 1812 612
rect 1766 608 1772 609
rect 134 597 140 598
rect 110 596 116 597
rect 110 592 111 596
rect 115 592 116 596
rect 134 593 135 597
rect 139 593 140 597
rect 134 592 140 593
rect 230 597 236 598
rect 230 593 231 597
rect 235 593 236 597
rect 230 592 236 593
rect 358 597 364 598
rect 358 593 359 597
rect 363 593 364 597
rect 358 592 364 593
rect 486 597 492 598
rect 486 593 487 597
rect 491 593 492 597
rect 486 592 492 593
rect 622 597 628 598
rect 622 593 623 597
rect 627 593 628 597
rect 622 592 628 593
rect 766 597 772 598
rect 766 593 767 597
rect 771 593 772 597
rect 766 592 772 593
rect 910 597 916 598
rect 910 593 911 597
rect 915 593 916 597
rect 910 592 916 593
rect 1054 597 1060 598
rect 1054 593 1055 597
rect 1059 593 1060 597
rect 1054 592 1060 593
rect 1206 597 1212 598
rect 1206 593 1207 597
rect 1211 593 1212 597
rect 1206 592 1212 593
rect 1366 597 1372 598
rect 1366 593 1367 597
rect 1371 593 1372 597
rect 1366 592 1372 593
rect 1526 597 1532 598
rect 1526 593 1527 597
rect 1531 593 1532 597
rect 1526 592 1532 593
rect 1670 597 1676 598
rect 1670 593 1671 597
rect 1675 593 1676 597
rect 1670 592 1676 593
rect 1766 596 1772 597
rect 1766 592 1767 596
rect 1771 592 1772 596
rect 110 591 116 592
rect 112 571 114 591
rect 136 571 138 592
rect 232 571 234 592
rect 360 571 362 592
rect 488 571 490 592
rect 624 571 626 592
rect 768 571 770 592
rect 912 571 914 592
rect 1056 571 1058 592
rect 1208 571 1210 592
rect 1368 571 1370 592
rect 1528 571 1530 592
rect 1672 571 1674 592
rect 1766 591 1772 592
rect 1768 571 1770 591
rect 1808 587 1810 611
rect 1976 587 1978 612
rect 2240 587 2242 612
rect 2480 587 2482 612
rect 2688 587 2690 612
rect 2880 587 2882 612
rect 3056 587 3058 612
rect 3224 587 3226 612
rect 3368 587 3370 612
rect 3462 611 3468 612
rect 3464 587 3466 611
rect 1807 586 1811 587
rect 1807 581 1811 582
rect 1895 586 1899 587
rect 1895 581 1899 582
rect 1975 586 1979 587
rect 1975 581 1979 582
rect 2015 586 2019 587
rect 2015 581 2019 582
rect 2143 586 2147 587
rect 2143 581 2147 582
rect 2239 586 2243 587
rect 2239 581 2243 582
rect 2279 586 2283 587
rect 2279 581 2283 582
rect 2423 586 2427 587
rect 2423 581 2427 582
rect 2479 586 2483 587
rect 2479 581 2483 582
rect 2567 586 2571 587
rect 2567 581 2571 582
rect 2687 586 2691 587
rect 2687 581 2691 582
rect 2719 586 2723 587
rect 2719 581 2723 582
rect 2871 586 2875 587
rect 2871 581 2875 582
rect 2879 586 2883 587
rect 2879 581 2883 582
rect 3031 586 3035 587
rect 3031 581 3035 582
rect 3055 586 3059 587
rect 3055 581 3059 582
rect 3199 586 3203 587
rect 3199 581 3203 582
rect 3223 586 3227 587
rect 3223 581 3227 582
rect 3367 586 3371 587
rect 3367 581 3371 582
rect 3463 586 3467 587
rect 3463 581 3467 582
rect 111 570 115 571
rect 111 565 115 566
rect 135 570 139 571
rect 135 565 139 566
rect 231 570 235 571
rect 231 565 235 566
rect 247 570 251 571
rect 247 565 251 566
rect 359 570 363 571
rect 359 565 363 566
rect 407 570 411 571
rect 407 565 411 566
rect 487 570 491 571
rect 487 565 491 566
rect 583 570 587 571
rect 583 565 587 566
rect 623 570 627 571
rect 623 565 627 566
rect 767 570 771 571
rect 767 565 771 566
rect 911 570 915 571
rect 911 565 915 566
rect 951 570 955 571
rect 951 565 955 566
rect 1055 570 1059 571
rect 1055 565 1059 566
rect 1135 570 1139 571
rect 1135 565 1139 566
rect 1207 570 1211 571
rect 1207 565 1211 566
rect 1319 570 1323 571
rect 1319 565 1323 566
rect 1367 570 1371 571
rect 1367 565 1371 566
rect 1503 570 1507 571
rect 1503 565 1507 566
rect 1527 570 1531 571
rect 1527 565 1531 566
rect 1671 570 1675 571
rect 1671 565 1675 566
rect 1767 570 1771 571
rect 1767 565 1771 566
rect 1808 565 1810 581
rect 112 549 114 565
rect 110 548 116 549
rect 136 548 138 565
rect 248 548 250 565
rect 408 548 410 565
rect 584 548 586 565
rect 768 548 770 565
rect 952 548 954 565
rect 1136 548 1138 565
rect 1320 548 1322 565
rect 1504 548 1506 565
rect 1672 548 1674 565
rect 1768 549 1770 565
rect 1806 564 1812 565
rect 1896 564 1898 581
rect 2016 564 2018 581
rect 2144 564 2146 581
rect 2280 564 2282 581
rect 2424 564 2426 581
rect 2568 564 2570 581
rect 2720 564 2722 581
rect 2872 564 2874 581
rect 3032 564 3034 581
rect 3200 564 3202 581
rect 3368 564 3370 581
rect 3464 565 3466 581
rect 3462 564 3468 565
rect 1806 560 1807 564
rect 1811 560 1812 564
rect 1806 559 1812 560
rect 1894 563 1900 564
rect 1894 559 1895 563
rect 1899 559 1900 563
rect 1894 558 1900 559
rect 2014 563 2020 564
rect 2014 559 2015 563
rect 2019 559 2020 563
rect 2014 558 2020 559
rect 2142 563 2148 564
rect 2142 559 2143 563
rect 2147 559 2148 563
rect 2142 558 2148 559
rect 2278 563 2284 564
rect 2278 559 2279 563
rect 2283 559 2284 563
rect 2278 558 2284 559
rect 2422 563 2428 564
rect 2422 559 2423 563
rect 2427 559 2428 563
rect 2422 558 2428 559
rect 2566 563 2572 564
rect 2566 559 2567 563
rect 2571 559 2572 563
rect 2566 558 2572 559
rect 2718 563 2724 564
rect 2718 559 2719 563
rect 2723 559 2724 563
rect 2718 558 2724 559
rect 2870 563 2876 564
rect 2870 559 2871 563
rect 2875 559 2876 563
rect 2870 558 2876 559
rect 3030 563 3036 564
rect 3030 559 3031 563
rect 3035 559 3036 563
rect 3030 558 3036 559
rect 3198 563 3204 564
rect 3198 559 3199 563
rect 3203 559 3204 563
rect 3198 558 3204 559
rect 3366 563 3372 564
rect 3366 559 3367 563
rect 3371 559 3372 563
rect 3462 560 3463 564
rect 3467 560 3468 564
rect 3462 559 3468 560
rect 3366 558 3372 559
rect 1766 548 1772 549
rect 110 544 111 548
rect 115 544 116 548
rect 110 543 116 544
rect 134 547 140 548
rect 134 543 135 547
rect 139 543 140 547
rect 134 542 140 543
rect 246 547 252 548
rect 246 543 247 547
rect 251 543 252 547
rect 246 542 252 543
rect 406 547 412 548
rect 406 543 407 547
rect 411 543 412 547
rect 406 542 412 543
rect 582 547 588 548
rect 582 543 583 547
rect 587 543 588 547
rect 582 542 588 543
rect 766 547 772 548
rect 766 543 767 547
rect 771 543 772 547
rect 766 542 772 543
rect 950 547 956 548
rect 950 543 951 547
rect 955 543 956 547
rect 950 542 956 543
rect 1134 547 1140 548
rect 1134 543 1135 547
rect 1139 543 1140 547
rect 1134 542 1140 543
rect 1318 547 1324 548
rect 1318 543 1319 547
rect 1323 543 1324 547
rect 1318 542 1324 543
rect 1502 547 1508 548
rect 1502 543 1503 547
rect 1507 543 1508 547
rect 1502 542 1508 543
rect 1670 547 1676 548
rect 1670 543 1671 547
rect 1675 543 1676 547
rect 1766 544 1767 548
rect 1771 544 1772 548
rect 1766 543 1772 544
rect 1806 547 1812 548
rect 1806 543 1807 547
rect 1811 543 1812 547
rect 3462 547 3468 548
rect 1670 542 1676 543
rect 1806 542 1812 543
rect 1894 544 1900 545
rect 110 531 116 532
rect 110 527 111 531
rect 115 527 116 531
rect 1766 531 1772 532
rect 110 526 116 527
rect 134 528 140 529
rect 112 503 114 526
rect 134 524 135 528
rect 139 524 140 528
rect 134 523 140 524
rect 246 528 252 529
rect 246 524 247 528
rect 251 524 252 528
rect 246 523 252 524
rect 406 528 412 529
rect 406 524 407 528
rect 411 524 412 528
rect 406 523 412 524
rect 582 528 588 529
rect 582 524 583 528
rect 587 524 588 528
rect 582 523 588 524
rect 766 528 772 529
rect 766 524 767 528
rect 771 524 772 528
rect 766 523 772 524
rect 950 528 956 529
rect 950 524 951 528
rect 955 524 956 528
rect 950 523 956 524
rect 1134 528 1140 529
rect 1134 524 1135 528
rect 1139 524 1140 528
rect 1134 523 1140 524
rect 1318 528 1324 529
rect 1318 524 1319 528
rect 1323 524 1324 528
rect 1318 523 1324 524
rect 1502 528 1508 529
rect 1502 524 1503 528
rect 1507 524 1508 528
rect 1502 523 1508 524
rect 1670 528 1676 529
rect 1670 524 1671 528
rect 1675 524 1676 528
rect 1766 527 1767 531
rect 1771 527 1772 531
rect 1766 526 1772 527
rect 1670 523 1676 524
rect 136 503 138 523
rect 248 503 250 523
rect 408 503 410 523
rect 584 503 586 523
rect 768 503 770 523
rect 952 503 954 523
rect 1136 503 1138 523
rect 1320 503 1322 523
rect 1504 503 1506 523
rect 1672 503 1674 523
rect 1768 503 1770 526
rect 1808 519 1810 542
rect 1894 540 1895 544
rect 1899 540 1900 544
rect 1894 539 1900 540
rect 2014 544 2020 545
rect 2014 540 2015 544
rect 2019 540 2020 544
rect 2014 539 2020 540
rect 2142 544 2148 545
rect 2142 540 2143 544
rect 2147 540 2148 544
rect 2142 539 2148 540
rect 2278 544 2284 545
rect 2278 540 2279 544
rect 2283 540 2284 544
rect 2278 539 2284 540
rect 2422 544 2428 545
rect 2422 540 2423 544
rect 2427 540 2428 544
rect 2422 539 2428 540
rect 2566 544 2572 545
rect 2566 540 2567 544
rect 2571 540 2572 544
rect 2566 539 2572 540
rect 2718 544 2724 545
rect 2718 540 2719 544
rect 2723 540 2724 544
rect 2718 539 2724 540
rect 2870 544 2876 545
rect 2870 540 2871 544
rect 2875 540 2876 544
rect 2870 539 2876 540
rect 3030 544 3036 545
rect 3030 540 3031 544
rect 3035 540 3036 544
rect 3030 539 3036 540
rect 3198 544 3204 545
rect 3198 540 3199 544
rect 3203 540 3204 544
rect 3198 539 3204 540
rect 3366 544 3372 545
rect 3366 540 3367 544
rect 3371 540 3372 544
rect 3462 543 3463 547
rect 3467 543 3468 547
rect 3462 542 3468 543
rect 3366 539 3372 540
rect 1896 519 1898 539
rect 2016 519 2018 539
rect 2144 519 2146 539
rect 2280 519 2282 539
rect 2424 519 2426 539
rect 2568 519 2570 539
rect 2720 519 2722 539
rect 2872 519 2874 539
rect 3032 519 3034 539
rect 3200 519 3202 539
rect 3368 519 3370 539
rect 3464 519 3466 542
rect 1807 518 1811 519
rect 1807 513 1811 514
rect 1895 518 1899 519
rect 1895 513 1899 514
rect 2015 518 2019 519
rect 2015 513 2019 514
rect 2135 518 2139 519
rect 2135 513 2139 514
rect 2143 518 2147 519
rect 2143 513 2147 514
rect 2239 518 2243 519
rect 2239 513 2243 514
rect 2279 518 2283 519
rect 2279 513 2283 514
rect 2359 518 2363 519
rect 2359 513 2363 514
rect 2423 518 2427 519
rect 2423 513 2427 514
rect 2487 518 2491 519
rect 2487 513 2491 514
rect 2567 518 2571 519
rect 2567 513 2571 514
rect 2615 518 2619 519
rect 2615 513 2619 514
rect 2719 518 2723 519
rect 2719 513 2723 514
rect 2751 518 2755 519
rect 2751 513 2755 514
rect 2871 518 2875 519
rect 2871 513 2875 514
rect 2879 518 2883 519
rect 2879 513 2883 514
rect 3007 518 3011 519
rect 3007 513 3011 514
rect 3031 518 3035 519
rect 3031 513 3035 514
rect 3135 518 3139 519
rect 3135 513 3139 514
rect 3199 518 3203 519
rect 3199 513 3203 514
rect 3263 518 3267 519
rect 3263 513 3267 514
rect 3367 518 3371 519
rect 3367 513 3371 514
rect 3463 518 3467 519
rect 3463 513 3467 514
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 247 502 251 503
rect 247 497 251 498
rect 399 502 403 503
rect 399 497 403 498
rect 407 502 411 503
rect 407 497 411 498
rect 567 502 571 503
rect 567 497 571 498
rect 583 502 587 503
rect 583 497 587 498
rect 735 502 739 503
rect 735 497 739 498
rect 767 502 771 503
rect 767 497 771 498
rect 903 502 907 503
rect 903 497 907 498
rect 951 502 955 503
rect 951 497 955 498
rect 1063 502 1067 503
rect 1063 497 1067 498
rect 1135 502 1139 503
rect 1135 497 1139 498
rect 1223 502 1227 503
rect 1223 497 1227 498
rect 1319 502 1323 503
rect 1319 497 1323 498
rect 1375 502 1379 503
rect 1375 497 1379 498
rect 1503 502 1507 503
rect 1503 497 1507 498
rect 1527 502 1531 503
rect 1527 497 1531 498
rect 1671 502 1675 503
rect 1671 497 1675 498
rect 1767 502 1771 503
rect 1767 497 1771 498
rect 112 478 114 497
rect 248 481 250 497
rect 400 481 402 497
rect 568 481 570 497
rect 736 481 738 497
rect 904 481 906 497
rect 1064 481 1066 497
rect 1224 481 1226 497
rect 1376 481 1378 497
rect 1528 481 1530 497
rect 1672 481 1674 497
rect 246 480 252 481
rect 110 477 116 478
rect 110 473 111 477
rect 115 473 116 477
rect 246 476 247 480
rect 251 476 252 480
rect 246 475 252 476
rect 398 480 404 481
rect 398 476 399 480
rect 403 476 404 480
rect 398 475 404 476
rect 566 480 572 481
rect 566 476 567 480
rect 571 476 572 480
rect 566 475 572 476
rect 734 480 740 481
rect 734 476 735 480
rect 739 476 740 480
rect 734 475 740 476
rect 902 480 908 481
rect 902 476 903 480
rect 907 476 908 480
rect 902 475 908 476
rect 1062 480 1068 481
rect 1062 476 1063 480
rect 1067 476 1068 480
rect 1062 475 1068 476
rect 1222 480 1228 481
rect 1222 476 1223 480
rect 1227 476 1228 480
rect 1222 475 1228 476
rect 1374 480 1380 481
rect 1374 476 1375 480
rect 1379 476 1380 480
rect 1374 475 1380 476
rect 1526 480 1532 481
rect 1526 476 1527 480
rect 1531 476 1532 480
rect 1526 475 1532 476
rect 1670 480 1676 481
rect 1670 476 1671 480
rect 1675 476 1676 480
rect 1768 478 1770 497
rect 1808 494 1810 513
rect 2136 497 2138 513
rect 2240 497 2242 513
rect 2360 497 2362 513
rect 2488 497 2490 513
rect 2616 497 2618 513
rect 2752 497 2754 513
rect 2880 497 2882 513
rect 3008 497 3010 513
rect 3136 497 3138 513
rect 3264 497 3266 513
rect 3368 497 3370 513
rect 2134 496 2140 497
rect 1806 493 1812 494
rect 1806 489 1807 493
rect 1811 489 1812 493
rect 2134 492 2135 496
rect 2139 492 2140 496
rect 2134 491 2140 492
rect 2238 496 2244 497
rect 2238 492 2239 496
rect 2243 492 2244 496
rect 2238 491 2244 492
rect 2358 496 2364 497
rect 2358 492 2359 496
rect 2363 492 2364 496
rect 2358 491 2364 492
rect 2486 496 2492 497
rect 2486 492 2487 496
rect 2491 492 2492 496
rect 2486 491 2492 492
rect 2614 496 2620 497
rect 2614 492 2615 496
rect 2619 492 2620 496
rect 2614 491 2620 492
rect 2750 496 2756 497
rect 2750 492 2751 496
rect 2755 492 2756 496
rect 2750 491 2756 492
rect 2878 496 2884 497
rect 2878 492 2879 496
rect 2883 492 2884 496
rect 2878 491 2884 492
rect 3006 496 3012 497
rect 3006 492 3007 496
rect 3011 492 3012 496
rect 3006 491 3012 492
rect 3134 496 3140 497
rect 3134 492 3135 496
rect 3139 492 3140 496
rect 3134 491 3140 492
rect 3262 496 3268 497
rect 3262 492 3263 496
rect 3267 492 3268 496
rect 3262 491 3268 492
rect 3366 496 3372 497
rect 3366 492 3367 496
rect 3371 492 3372 496
rect 3464 494 3466 513
rect 3366 491 3372 492
rect 3462 493 3468 494
rect 1806 488 1812 489
rect 3462 489 3463 493
rect 3467 489 3468 493
rect 3462 488 3468 489
rect 1670 475 1676 476
rect 1766 477 1772 478
rect 2134 477 2140 478
rect 110 472 116 473
rect 1766 473 1767 477
rect 1771 473 1772 477
rect 1766 472 1772 473
rect 1806 476 1812 477
rect 1806 472 1807 476
rect 1811 472 1812 476
rect 2134 473 2135 477
rect 2139 473 2140 477
rect 2134 472 2140 473
rect 2238 477 2244 478
rect 2238 473 2239 477
rect 2243 473 2244 477
rect 2238 472 2244 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 2486 477 2492 478
rect 2486 473 2487 477
rect 2491 473 2492 477
rect 2486 472 2492 473
rect 2614 477 2620 478
rect 2614 473 2615 477
rect 2619 473 2620 477
rect 2614 472 2620 473
rect 2750 477 2756 478
rect 2750 473 2751 477
rect 2755 473 2756 477
rect 2750 472 2756 473
rect 2878 477 2884 478
rect 2878 473 2879 477
rect 2883 473 2884 477
rect 2878 472 2884 473
rect 3006 477 3012 478
rect 3006 473 3007 477
rect 3011 473 3012 477
rect 3006 472 3012 473
rect 3134 477 3140 478
rect 3134 473 3135 477
rect 3139 473 3140 477
rect 3134 472 3140 473
rect 3262 477 3268 478
rect 3262 473 3263 477
rect 3267 473 3268 477
rect 3262 472 3268 473
rect 3366 477 3372 478
rect 3366 473 3367 477
rect 3371 473 3372 477
rect 3366 472 3372 473
rect 3462 476 3468 477
rect 3462 472 3463 476
rect 3467 472 3468 476
rect 1806 471 1812 472
rect 246 461 252 462
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 246 457 247 461
rect 251 457 252 461
rect 246 456 252 457
rect 398 461 404 462
rect 398 457 399 461
rect 403 457 404 461
rect 398 456 404 457
rect 566 461 572 462
rect 566 457 567 461
rect 571 457 572 461
rect 566 456 572 457
rect 734 461 740 462
rect 734 457 735 461
rect 739 457 740 461
rect 734 456 740 457
rect 902 461 908 462
rect 902 457 903 461
rect 907 457 908 461
rect 902 456 908 457
rect 1062 461 1068 462
rect 1062 457 1063 461
rect 1067 457 1068 461
rect 1062 456 1068 457
rect 1222 461 1228 462
rect 1222 457 1223 461
rect 1227 457 1228 461
rect 1222 456 1228 457
rect 1374 461 1380 462
rect 1374 457 1375 461
rect 1379 457 1380 461
rect 1374 456 1380 457
rect 1526 461 1532 462
rect 1526 457 1527 461
rect 1531 457 1532 461
rect 1526 456 1532 457
rect 1670 461 1676 462
rect 1670 457 1671 461
rect 1675 457 1676 461
rect 1670 456 1676 457
rect 1766 460 1772 461
rect 1766 456 1767 460
rect 1771 456 1772 460
rect 110 455 116 456
rect 112 435 114 455
rect 248 435 250 456
rect 400 435 402 456
rect 568 435 570 456
rect 736 435 738 456
rect 904 435 906 456
rect 1064 435 1066 456
rect 1224 435 1226 456
rect 1376 435 1378 456
rect 1528 435 1530 456
rect 1672 435 1674 456
rect 1766 455 1772 456
rect 1768 435 1770 455
rect 1808 447 1810 471
rect 2136 447 2138 472
rect 2240 447 2242 472
rect 2360 447 2362 472
rect 2488 447 2490 472
rect 2616 447 2618 472
rect 2752 447 2754 472
rect 2880 447 2882 472
rect 3008 447 3010 472
rect 3136 447 3138 472
rect 3264 447 3266 472
rect 3368 447 3370 472
rect 3462 471 3468 472
rect 3464 447 3466 471
rect 1807 446 1811 447
rect 1807 441 1811 442
rect 2135 446 2139 447
rect 2135 441 2139 442
rect 2239 446 2243 447
rect 2239 441 2243 442
rect 2335 446 2339 447
rect 2335 441 2339 442
rect 2359 446 2363 447
rect 2359 441 2363 442
rect 2447 446 2451 447
rect 2447 441 2451 442
rect 2487 446 2491 447
rect 2487 441 2491 442
rect 2559 446 2563 447
rect 2559 441 2563 442
rect 2615 446 2619 447
rect 2615 441 2619 442
rect 2679 446 2683 447
rect 2679 441 2683 442
rect 2751 446 2755 447
rect 2751 441 2755 442
rect 2799 446 2803 447
rect 2799 441 2803 442
rect 2879 446 2883 447
rect 2879 441 2883 442
rect 2911 446 2915 447
rect 2911 441 2915 442
rect 3007 446 3011 447
rect 3007 441 3011 442
rect 3023 446 3027 447
rect 3023 441 3027 442
rect 3135 446 3139 447
rect 3135 441 3139 442
rect 3143 446 3147 447
rect 3143 441 3147 442
rect 3263 446 3267 447
rect 3263 441 3267 442
rect 3367 446 3371 447
rect 3367 441 3371 442
rect 3463 446 3467 447
rect 3463 441 3467 442
rect 111 434 115 435
rect 111 429 115 430
rect 247 434 251 435
rect 247 429 251 430
rect 399 434 403 435
rect 399 429 403 430
rect 519 434 523 435
rect 519 429 523 430
rect 567 434 571 435
rect 567 429 571 430
rect 615 434 619 435
rect 615 429 619 430
rect 719 434 723 435
rect 719 429 723 430
rect 735 434 739 435
rect 735 429 739 430
rect 823 434 827 435
rect 823 429 827 430
rect 903 434 907 435
rect 903 429 907 430
rect 927 434 931 435
rect 927 429 931 430
rect 1023 434 1027 435
rect 1023 429 1027 430
rect 1063 434 1067 435
rect 1063 429 1067 430
rect 1127 434 1131 435
rect 1127 429 1131 430
rect 1223 434 1227 435
rect 1223 429 1227 430
rect 1231 434 1235 435
rect 1231 429 1235 430
rect 1335 434 1339 435
rect 1335 429 1339 430
rect 1375 434 1379 435
rect 1375 429 1379 430
rect 1439 434 1443 435
rect 1439 429 1443 430
rect 1527 434 1531 435
rect 1527 429 1531 430
rect 1671 434 1675 435
rect 1671 429 1675 430
rect 1767 434 1771 435
rect 1767 429 1771 430
rect 112 413 114 429
rect 110 412 116 413
rect 520 412 522 429
rect 616 412 618 429
rect 720 412 722 429
rect 824 412 826 429
rect 928 412 930 429
rect 1024 412 1026 429
rect 1128 412 1130 429
rect 1232 412 1234 429
rect 1336 412 1338 429
rect 1440 412 1442 429
rect 1768 413 1770 429
rect 1808 425 1810 441
rect 1806 424 1812 425
rect 2240 424 2242 441
rect 2336 424 2338 441
rect 2448 424 2450 441
rect 2560 424 2562 441
rect 2680 424 2682 441
rect 2800 424 2802 441
rect 2912 424 2914 441
rect 3024 424 3026 441
rect 3144 424 3146 441
rect 3264 424 3266 441
rect 3368 424 3370 441
rect 3464 425 3466 441
rect 3462 424 3468 425
rect 1806 420 1807 424
rect 1811 420 1812 424
rect 1806 419 1812 420
rect 2238 423 2244 424
rect 2238 419 2239 423
rect 2243 419 2244 423
rect 2238 418 2244 419
rect 2334 423 2340 424
rect 2334 419 2335 423
rect 2339 419 2340 423
rect 2334 418 2340 419
rect 2446 423 2452 424
rect 2446 419 2447 423
rect 2451 419 2452 423
rect 2446 418 2452 419
rect 2558 423 2564 424
rect 2558 419 2559 423
rect 2563 419 2564 423
rect 2558 418 2564 419
rect 2678 423 2684 424
rect 2678 419 2679 423
rect 2683 419 2684 423
rect 2678 418 2684 419
rect 2798 423 2804 424
rect 2798 419 2799 423
rect 2803 419 2804 423
rect 2798 418 2804 419
rect 2910 423 2916 424
rect 2910 419 2911 423
rect 2915 419 2916 423
rect 2910 418 2916 419
rect 3022 423 3028 424
rect 3022 419 3023 423
rect 3027 419 3028 423
rect 3022 418 3028 419
rect 3142 423 3148 424
rect 3142 419 3143 423
rect 3147 419 3148 423
rect 3142 418 3148 419
rect 3262 423 3268 424
rect 3262 419 3263 423
rect 3267 419 3268 423
rect 3262 418 3268 419
rect 3366 423 3372 424
rect 3366 419 3367 423
rect 3371 419 3372 423
rect 3462 420 3463 424
rect 3467 420 3468 424
rect 3462 419 3468 420
rect 3366 418 3372 419
rect 1766 412 1772 413
rect 110 408 111 412
rect 115 408 116 412
rect 110 407 116 408
rect 518 411 524 412
rect 518 407 519 411
rect 523 407 524 411
rect 518 406 524 407
rect 614 411 620 412
rect 614 407 615 411
rect 619 407 620 411
rect 614 406 620 407
rect 718 411 724 412
rect 718 407 719 411
rect 723 407 724 411
rect 718 406 724 407
rect 822 411 828 412
rect 822 407 823 411
rect 827 407 828 411
rect 822 406 828 407
rect 926 411 932 412
rect 926 407 927 411
rect 931 407 932 411
rect 926 406 932 407
rect 1022 411 1028 412
rect 1022 407 1023 411
rect 1027 407 1028 411
rect 1022 406 1028 407
rect 1126 411 1132 412
rect 1126 407 1127 411
rect 1131 407 1132 411
rect 1126 406 1132 407
rect 1230 411 1236 412
rect 1230 407 1231 411
rect 1235 407 1236 411
rect 1230 406 1236 407
rect 1334 411 1340 412
rect 1334 407 1335 411
rect 1339 407 1340 411
rect 1334 406 1340 407
rect 1438 411 1444 412
rect 1438 407 1439 411
rect 1443 407 1444 411
rect 1766 408 1767 412
rect 1771 408 1772 412
rect 1766 407 1772 408
rect 1806 407 1812 408
rect 1438 406 1444 407
rect 1806 403 1807 407
rect 1811 403 1812 407
rect 3462 407 3468 408
rect 1806 402 1812 403
rect 2238 404 2244 405
rect 110 395 116 396
rect 110 391 111 395
rect 115 391 116 395
rect 1766 395 1772 396
rect 110 390 116 391
rect 518 392 524 393
rect 112 367 114 390
rect 518 388 519 392
rect 523 388 524 392
rect 518 387 524 388
rect 614 392 620 393
rect 614 388 615 392
rect 619 388 620 392
rect 614 387 620 388
rect 718 392 724 393
rect 718 388 719 392
rect 723 388 724 392
rect 718 387 724 388
rect 822 392 828 393
rect 822 388 823 392
rect 827 388 828 392
rect 822 387 828 388
rect 926 392 932 393
rect 926 388 927 392
rect 931 388 932 392
rect 926 387 932 388
rect 1022 392 1028 393
rect 1022 388 1023 392
rect 1027 388 1028 392
rect 1022 387 1028 388
rect 1126 392 1132 393
rect 1126 388 1127 392
rect 1131 388 1132 392
rect 1126 387 1132 388
rect 1230 392 1236 393
rect 1230 388 1231 392
rect 1235 388 1236 392
rect 1230 387 1236 388
rect 1334 392 1340 393
rect 1334 388 1335 392
rect 1339 388 1340 392
rect 1334 387 1340 388
rect 1438 392 1444 393
rect 1438 388 1439 392
rect 1443 388 1444 392
rect 1766 391 1767 395
rect 1771 391 1772 395
rect 1766 390 1772 391
rect 1438 387 1444 388
rect 520 367 522 387
rect 616 367 618 387
rect 720 367 722 387
rect 824 367 826 387
rect 928 367 930 387
rect 1024 367 1026 387
rect 1128 367 1130 387
rect 1232 367 1234 387
rect 1336 367 1338 387
rect 1440 367 1442 387
rect 1768 367 1770 390
rect 1808 379 1810 402
rect 2238 400 2239 404
rect 2243 400 2244 404
rect 2238 399 2244 400
rect 2334 404 2340 405
rect 2334 400 2335 404
rect 2339 400 2340 404
rect 2334 399 2340 400
rect 2446 404 2452 405
rect 2446 400 2447 404
rect 2451 400 2452 404
rect 2446 399 2452 400
rect 2558 404 2564 405
rect 2558 400 2559 404
rect 2563 400 2564 404
rect 2558 399 2564 400
rect 2678 404 2684 405
rect 2678 400 2679 404
rect 2683 400 2684 404
rect 2678 399 2684 400
rect 2798 404 2804 405
rect 2798 400 2799 404
rect 2803 400 2804 404
rect 2798 399 2804 400
rect 2910 404 2916 405
rect 2910 400 2911 404
rect 2915 400 2916 404
rect 2910 399 2916 400
rect 3022 404 3028 405
rect 3022 400 3023 404
rect 3027 400 3028 404
rect 3022 399 3028 400
rect 3142 404 3148 405
rect 3142 400 3143 404
rect 3147 400 3148 404
rect 3142 399 3148 400
rect 3262 404 3268 405
rect 3262 400 3263 404
rect 3267 400 3268 404
rect 3262 399 3268 400
rect 3366 404 3372 405
rect 3366 400 3367 404
rect 3371 400 3372 404
rect 3462 403 3463 407
rect 3467 403 3468 407
rect 3462 402 3468 403
rect 3366 399 3372 400
rect 2240 379 2242 399
rect 2336 379 2338 399
rect 2448 379 2450 399
rect 2560 379 2562 399
rect 2680 379 2682 399
rect 2800 379 2802 399
rect 2912 379 2914 399
rect 3024 379 3026 399
rect 3144 379 3146 399
rect 3264 379 3266 399
rect 3368 379 3370 399
rect 3464 379 3466 402
rect 1807 378 1811 379
rect 1807 373 1811 374
rect 2063 378 2067 379
rect 2063 373 2067 374
rect 2151 378 2155 379
rect 2151 373 2155 374
rect 2239 378 2243 379
rect 2239 373 2243 374
rect 2247 378 2251 379
rect 2247 373 2251 374
rect 2335 378 2339 379
rect 2335 373 2339 374
rect 2359 378 2363 379
rect 2359 373 2363 374
rect 2447 378 2451 379
rect 2447 373 2451 374
rect 2479 378 2483 379
rect 2479 373 2483 374
rect 2559 378 2563 379
rect 2559 373 2563 374
rect 2615 378 2619 379
rect 2615 373 2619 374
rect 2679 378 2683 379
rect 2679 373 2683 374
rect 2759 378 2763 379
rect 2759 373 2763 374
rect 2799 378 2803 379
rect 2799 373 2803 374
rect 2911 378 2915 379
rect 2911 373 2915 374
rect 3023 378 3027 379
rect 3023 373 3027 374
rect 3063 378 3067 379
rect 3063 373 3067 374
rect 3143 378 3147 379
rect 3143 373 3147 374
rect 3223 378 3227 379
rect 3223 373 3227 374
rect 3263 378 3267 379
rect 3263 373 3267 374
rect 3367 378 3371 379
rect 3367 373 3371 374
rect 3463 378 3467 379
rect 3463 373 3467 374
rect 111 366 115 367
rect 111 361 115 362
rect 471 366 475 367
rect 471 361 475 362
rect 519 366 523 367
rect 519 361 523 362
rect 559 366 563 367
rect 559 361 563 362
rect 615 366 619 367
rect 615 361 619 362
rect 647 366 651 367
rect 647 361 651 362
rect 719 366 723 367
rect 719 361 723 362
rect 735 366 739 367
rect 735 361 739 362
rect 823 366 827 367
rect 823 361 827 362
rect 911 366 915 367
rect 911 361 915 362
rect 927 366 931 367
rect 927 361 931 362
rect 999 366 1003 367
rect 999 361 1003 362
rect 1023 366 1027 367
rect 1023 361 1027 362
rect 1087 366 1091 367
rect 1087 361 1091 362
rect 1127 366 1131 367
rect 1127 361 1131 362
rect 1175 366 1179 367
rect 1175 361 1179 362
rect 1231 366 1235 367
rect 1231 361 1235 362
rect 1263 366 1267 367
rect 1263 361 1267 362
rect 1335 366 1339 367
rect 1335 361 1339 362
rect 1439 366 1443 367
rect 1439 361 1443 362
rect 1767 366 1771 367
rect 1767 361 1771 362
rect 112 342 114 361
rect 472 345 474 361
rect 560 345 562 361
rect 648 345 650 361
rect 736 345 738 361
rect 824 345 826 361
rect 912 345 914 361
rect 1000 345 1002 361
rect 1088 345 1090 361
rect 1176 345 1178 361
rect 1264 345 1266 361
rect 470 344 476 345
rect 110 341 116 342
rect 110 337 111 341
rect 115 337 116 341
rect 470 340 471 344
rect 475 340 476 344
rect 470 339 476 340
rect 558 344 564 345
rect 558 340 559 344
rect 563 340 564 344
rect 558 339 564 340
rect 646 344 652 345
rect 646 340 647 344
rect 651 340 652 344
rect 646 339 652 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 822 344 828 345
rect 822 340 823 344
rect 827 340 828 344
rect 822 339 828 340
rect 910 344 916 345
rect 910 340 911 344
rect 915 340 916 344
rect 910 339 916 340
rect 998 344 1004 345
rect 998 340 999 344
rect 1003 340 1004 344
rect 998 339 1004 340
rect 1086 344 1092 345
rect 1086 340 1087 344
rect 1091 340 1092 344
rect 1086 339 1092 340
rect 1174 344 1180 345
rect 1174 340 1175 344
rect 1179 340 1180 344
rect 1174 339 1180 340
rect 1262 344 1268 345
rect 1262 340 1263 344
rect 1267 340 1268 344
rect 1768 342 1770 361
rect 1808 354 1810 373
rect 2064 357 2066 373
rect 2152 357 2154 373
rect 2248 357 2250 373
rect 2360 357 2362 373
rect 2480 357 2482 373
rect 2616 357 2618 373
rect 2760 357 2762 373
rect 2912 357 2914 373
rect 3064 357 3066 373
rect 3224 357 3226 373
rect 3368 357 3370 373
rect 2062 356 2068 357
rect 1806 353 1812 354
rect 1806 349 1807 353
rect 1811 349 1812 353
rect 2062 352 2063 356
rect 2067 352 2068 356
rect 2062 351 2068 352
rect 2150 356 2156 357
rect 2150 352 2151 356
rect 2155 352 2156 356
rect 2150 351 2156 352
rect 2246 356 2252 357
rect 2246 352 2247 356
rect 2251 352 2252 356
rect 2246 351 2252 352
rect 2358 356 2364 357
rect 2358 352 2359 356
rect 2363 352 2364 356
rect 2358 351 2364 352
rect 2478 356 2484 357
rect 2478 352 2479 356
rect 2483 352 2484 356
rect 2478 351 2484 352
rect 2614 356 2620 357
rect 2614 352 2615 356
rect 2619 352 2620 356
rect 2614 351 2620 352
rect 2758 356 2764 357
rect 2758 352 2759 356
rect 2763 352 2764 356
rect 2758 351 2764 352
rect 2910 356 2916 357
rect 2910 352 2911 356
rect 2915 352 2916 356
rect 2910 351 2916 352
rect 3062 356 3068 357
rect 3062 352 3063 356
rect 3067 352 3068 356
rect 3062 351 3068 352
rect 3222 356 3228 357
rect 3222 352 3223 356
rect 3227 352 3228 356
rect 3222 351 3228 352
rect 3366 356 3372 357
rect 3366 352 3367 356
rect 3371 352 3372 356
rect 3464 354 3466 373
rect 3366 351 3372 352
rect 3462 353 3468 354
rect 1806 348 1812 349
rect 3462 349 3463 353
rect 3467 349 3468 353
rect 3462 348 3468 349
rect 1262 339 1268 340
rect 1766 341 1772 342
rect 110 336 116 337
rect 1766 337 1767 341
rect 1771 337 1772 341
rect 2062 337 2068 338
rect 1766 336 1772 337
rect 1806 336 1812 337
rect 1806 332 1807 336
rect 1811 332 1812 336
rect 2062 333 2063 337
rect 2067 333 2068 337
rect 2062 332 2068 333
rect 2150 337 2156 338
rect 2150 333 2151 337
rect 2155 333 2156 337
rect 2150 332 2156 333
rect 2246 337 2252 338
rect 2246 333 2247 337
rect 2251 333 2252 337
rect 2246 332 2252 333
rect 2358 337 2364 338
rect 2358 333 2359 337
rect 2363 333 2364 337
rect 2358 332 2364 333
rect 2478 337 2484 338
rect 2478 333 2479 337
rect 2483 333 2484 337
rect 2478 332 2484 333
rect 2614 337 2620 338
rect 2614 333 2615 337
rect 2619 333 2620 337
rect 2614 332 2620 333
rect 2758 337 2764 338
rect 2758 333 2759 337
rect 2763 333 2764 337
rect 2758 332 2764 333
rect 2910 337 2916 338
rect 2910 333 2911 337
rect 2915 333 2916 337
rect 2910 332 2916 333
rect 3062 337 3068 338
rect 3062 333 3063 337
rect 3067 333 3068 337
rect 3062 332 3068 333
rect 3222 337 3228 338
rect 3222 333 3223 337
rect 3227 333 3228 337
rect 3222 332 3228 333
rect 3366 337 3372 338
rect 3366 333 3367 337
rect 3371 333 3372 337
rect 3366 332 3372 333
rect 3462 336 3468 337
rect 3462 332 3463 336
rect 3467 332 3468 336
rect 1806 331 1812 332
rect 470 325 476 326
rect 110 324 116 325
rect 110 320 111 324
rect 115 320 116 324
rect 470 321 471 325
rect 475 321 476 325
rect 470 320 476 321
rect 558 325 564 326
rect 558 321 559 325
rect 563 321 564 325
rect 558 320 564 321
rect 646 325 652 326
rect 646 321 647 325
rect 651 321 652 325
rect 646 320 652 321
rect 734 325 740 326
rect 734 321 735 325
rect 739 321 740 325
rect 734 320 740 321
rect 822 325 828 326
rect 822 321 823 325
rect 827 321 828 325
rect 822 320 828 321
rect 910 325 916 326
rect 910 321 911 325
rect 915 321 916 325
rect 910 320 916 321
rect 998 325 1004 326
rect 998 321 999 325
rect 1003 321 1004 325
rect 998 320 1004 321
rect 1086 325 1092 326
rect 1086 321 1087 325
rect 1091 321 1092 325
rect 1086 320 1092 321
rect 1174 325 1180 326
rect 1174 321 1175 325
rect 1179 321 1180 325
rect 1174 320 1180 321
rect 1262 325 1268 326
rect 1262 321 1263 325
rect 1267 321 1268 325
rect 1262 320 1268 321
rect 1766 324 1772 325
rect 1766 320 1767 324
rect 1771 320 1772 324
rect 110 319 116 320
rect 112 299 114 319
rect 472 299 474 320
rect 560 299 562 320
rect 648 299 650 320
rect 736 299 738 320
rect 824 299 826 320
rect 912 299 914 320
rect 1000 299 1002 320
rect 1088 299 1090 320
rect 1176 299 1178 320
rect 1264 299 1266 320
rect 1766 319 1772 320
rect 1768 299 1770 319
rect 1808 311 1810 331
rect 2064 311 2066 332
rect 2152 311 2154 332
rect 2248 311 2250 332
rect 2360 311 2362 332
rect 2480 311 2482 332
rect 2616 311 2618 332
rect 2760 311 2762 332
rect 2912 311 2914 332
rect 3064 311 3066 332
rect 3224 311 3226 332
rect 3368 311 3370 332
rect 3462 331 3468 332
rect 3464 311 3466 331
rect 1807 310 1811 311
rect 1807 305 1811 306
rect 1927 310 1931 311
rect 1927 305 1931 306
rect 2039 310 2043 311
rect 2039 305 2043 306
rect 2063 310 2067 311
rect 2063 305 2067 306
rect 2151 310 2155 311
rect 2151 305 2155 306
rect 2167 310 2171 311
rect 2167 305 2171 306
rect 2247 310 2251 311
rect 2247 305 2251 306
rect 2303 310 2307 311
rect 2303 305 2307 306
rect 2359 310 2363 311
rect 2359 305 2363 306
rect 2447 310 2451 311
rect 2447 305 2451 306
rect 2479 310 2483 311
rect 2479 305 2483 306
rect 2599 310 2603 311
rect 2599 305 2603 306
rect 2615 310 2619 311
rect 2615 305 2619 306
rect 2759 310 2763 311
rect 2759 305 2763 306
rect 2911 310 2915 311
rect 2911 305 2915 306
rect 2919 310 2923 311
rect 2919 305 2923 306
rect 3063 310 3067 311
rect 3063 305 3067 306
rect 3087 310 3091 311
rect 3087 305 3091 306
rect 3223 310 3227 311
rect 3223 305 3227 306
rect 3255 310 3259 311
rect 3255 305 3259 306
rect 3367 310 3371 311
rect 3367 305 3371 306
rect 3463 310 3467 311
rect 3463 305 3467 306
rect 111 298 115 299
rect 111 293 115 294
rect 279 298 283 299
rect 279 293 283 294
rect 367 298 371 299
rect 367 293 371 294
rect 463 298 467 299
rect 463 293 467 294
rect 471 298 475 299
rect 471 293 475 294
rect 559 298 563 299
rect 559 293 563 294
rect 647 298 651 299
rect 647 293 651 294
rect 655 298 659 299
rect 655 293 659 294
rect 735 298 739 299
rect 735 293 739 294
rect 751 298 755 299
rect 751 293 755 294
rect 823 298 827 299
rect 823 293 827 294
rect 847 298 851 299
rect 847 293 851 294
rect 911 298 915 299
rect 911 293 915 294
rect 943 298 947 299
rect 943 293 947 294
rect 999 298 1003 299
rect 999 293 1003 294
rect 1047 298 1051 299
rect 1047 293 1051 294
rect 1087 298 1091 299
rect 1087 293 1091 294
rect 1151 298 1155 299
rect 1151 293 1155 294
rect 1175 298 1179 299
rect 1175 293 1179 294
rect 1263 298 1267 299
rect 1263 293 1267 294
rect 1767 298 1771 299
rect 1767 293 1771 294
rect 112 277 114 293
rect 110 276 116 277
rect 280 276 282 293
rect 368 276 370 293
rect 464 276 466 293
rect 560 276 562 293
rect 656 276 658 293
rect 752 276 754 293
rect 848 276 850 293
rect 944 276 946 293
rect 1048 276 1050 293
rect 1152 276 1154 293
rect 1768 277 1770 293
rect 1808 289 1810 305
rect 1806 288 1812 289
rect 1928 288 1930 305
rect 2040 288 2042 305
rect 2168 288 2170 305
rect 2304 288 2306 305
rect 2448 288 2450 305
rect 2600 288 2602 305
rect 2760 288 2762 305
rect 2920 288 2922 305
rect 3088 288 3090 305
rect 3256 288 3258 305
rect 3464 289 3466 305
rect 3462 288 3468 289
rect 1806 284 1807 288
rect 1811 284 1812 288
rect 1806 283 1812 284
rect 1926 287 1932 288
rect 1926 283 1927 287
rect 1931 283 1932 287
rect 1926 282 1932 283
rect 2038 287 2044 288
rect 2038 283 2039 287
rect 2043 283 2044 287
rect 2038 282 2044 283
rect 2166 287 2172 288
rect 2166 283 2167 287
rect 2171 283 2172 287
rect 2166 282 2172 283
rect 2302 287 2308 288
rect 2302 283 2303 287
rect 2307 283 2308 287
rect 2302 282 2308 283
rect 2446 287 2452 288
rect 2446 283 2447 287
rect 2451 283 2452 287
rect 2446 282 2452 283
rect 2598 287 2604 288
rect 2598 283 2599 287
rect 2603 283 2604 287
rect 2598 282 2604 283
rect 2758 287 2764 288
rect 2758 283 2759 287
rect 2763 283 2764 287
rect 2758 282 2764 283
rect 2918 287 2924 288
rect 2918 283 2919 287
rect 2923 283 2924 287
rect 2918 282 2924 283
rect 3086 287 3092 288
rect 3086 283 3087 287
rect 3091 283 3092 287
rect 3086 282 3092 283
rect 3254 287 3260 288
rect 3254 283 3255 287
rect 3259 283 3260 287
rect 3462 284 3463 288
rect 3467 284 3468 288
rect 3462 283 3468 284
rect 3254 282 3260 283
rect 1766 276 1772 277
rect 110 272 111 276
rect 115 272 116 276
rect 110 271 116 272
rect 278 275 284 276
rect 278 271 279 275
rect 283 271 284 275
rect 278 270 284 271
rect 366 275 372 276
rect 366 271 367 275
rect 371 271 372 275
rect 366 270 372 271
rect 462 275 468 276
rect 462 271 463 275
rect 467 271 468 275
rect 462 270 468 271
rect 558 275 564 276
rect 558 271 559 275
rect 563 271 564 275
rect 558 270 564 271
rect 654 275 660 276
rect 654 271 655 275
rect 659 271 660 275
rect 654 270 660 271
rect 750 275 756 276
rect 750 271 751 275
rect 755 271 756 275
rect 750 270 756 271
rect 846 275 852 276
rect 846 271 847 275
rect 851 271 852 275
rect 846 270 852 271
rect 942 275 948 276
rect 942 271 943 275
rect 947 271 948 275
rect 942 270 948 271
rect 1046 275 1052 276
rect 1046 271 1047 275
rect 1051 271 1052 275
rect 1046 270 1052 271
rect 1150 275 1156 276
rect 1150 271 1151 275
rect 1155 271 1156 275
rect 1766 272 1767 276
rect 1771 272 1772 276
rect 1766 271 1772 272
rect 1806 271 1812 272
rect 1150 270 1156 271
rect 1806 267 1807 271
rect 1811 267 1812 271
rect 3462 271 3468 272
rect 1806 266 1812 267
rect 1926 268 1932 269
rect 110 259 116 260
rect 110 255 111 259
rect 115 255 116 259
rect 1766 259 1772 260
rect 110 254 116 255
rect 278 256 284 257
rect 112 231 114 254
rect 278 252 279 256
rect 283 252 284 256
rect 278 251 284 252
rect 366 256 372 257
rect 366 252 367 256
rect 371 252 372 256
rect 366 251 372 252
rect 462 256 468 257
rect 462 252 463 256
rect 467 252 468 256
rect 462 251 468 252
rect 558 256 564 257
rect 558 252 559 256
rect 563 252 564 256
rect 558 251 564 252
rect 654 256 660 257
rect 654 252 655 256
rect 659 252 660 256
rect 654 251 660 252
rect 750 256 756 257
rect 750 252 751 256
rect 755 252 756 256
rect 750 251 756 252
rect 846 256 852 257
rect 846 252 847 256
rect 851 252 852 256
rect 846 251 852 252
rect 942 256 948 257
rect 942 252 943 256
rect 947 252 948 256
rect 942 251 948 252
rect 1046 256 1052 257
rect 1046 252 1047 256
rect 1051 252 1052 256
rect 1046 251 1052 252
rect 1150 256 1156 257
rect 1150 252 1151 256
rect 1155 252 1156 256
rect 1766 255 1767 259
rect 1771 255 1772 259
rect 1766 254 1772 255
rect 1150 251 1156 252
rect 280 231 282 251
rect 368 231 370 251
rect 464 231 466 251
rect 560 231 562 251
rect 656 231 658 251
rect 752 231 754 251
rect 848 231 850 251
rect 944 231 946 251
rect 1048 231 1050 251
rect 1152 231 1154 251
rect 1768 231 1770 254
rect 1808 243 1810 266
rect 1926 264 1927 268
rect 1931 264 1932 268
rect 1926 263 1932 264
rect 2038 268 2044 269
rect 2038 264 2039 268
rect 2043 264 2044 268
rect 2038 263 2044 264
rect 2166 268 2172 269
rect 2166 264 2167 268
rect 2171 264 2172 268
rect 2166 263 2172 264
rect 2302 268 2308 269
rect 2302 264 2303 268
rect 2307 264 2308 268
rect 2302 263 2308 264
rect 2446 268 2452 269
rect 2446 264 2447 268
rect 2451 264 2452 268
rect 2446 263 2452 264
rect 2598 268 2604 269
rect 2598 264 2599 268
rect 2603 264 2604 268
rect 2598 263 2604 264
rect 2758 268 2764 269
rect 2758 264 2759 268
rect 2763 264 2764 268
rect 2758 263 2764 264
rect 2918 268 2924 269
rect 2918 264 2919 268
rect 2923 264 2924 268
rect 2918 263 2924 264
rect 3086 268 3092 269
rect 3086 264 3087 268
rect 3091 264 3092 268
rect 3086 263 3092 264
rect 3254 268 3260 269
rect 3254 264 3255 268
rect 3259 264 3260 268
rect 3462 267 3463 271
rect 3467 267 3468 271
rect 3462 266 3468 267
rect 3254 263 3260 264
rect 1928 243 1930 263
rect 2040 243 2042 263
rect 2168 243 2170 263
rect 2304 243 2306 263
rect 2448 243 2450 263
rect 2600 243 2602 263
rect 2760 243 2762 263
rect 2920 243 2922 263
rect 3088 243 3090 263
rect 3256 243 3258 263
rect 3464 243 3466 266
rect 1807 242 1811 243
rect 1807 237 1811 238
rect 1831 242 1835 243
rect 1831 237 1835 238
rect 1927 242 1931 243
rect 1927 237 1931 238
rect 2039 242 2043 243
rect 2039 237 2043 238
rect 2055 242 2059 243
rect 2055 237 2059 238
rect 2167 242 2171 243
rect 2167 237 2171 238
rect 2199 242 2203 243
rect 2199 237 2203 238
rect 2303 242 2307 243
rect 2303 237 2307 238
rect 2351 242 2355 243
rect 2351 237 2355 238
rect 2447 242 2451 243
rect 2447 237 2451 238
rect 2511 242 2515 243
rect 2511 237 2515 238
rect 2599 242 2603 243
rect 2599 237 2603 238
rect 2679 242 2683 243
rect 2679 237 2683 238
rect 2759 242 2763 243
rect 2759 237 2763 238
rect 2847 242 2851 243
rect 2847 237 2851 238
rect 2919 242 2923 243
rect 2919 237 2923 238
rect 3023 242 3027 243
rect 3023 237 3027 238
rect 3087 242 3091 243
rect 3087 237 3091 238
rect 3207 242 3211 243
rect 3207 237 3211 238
rect 3255 242 3259 243
rect 3255 237 3259 238
rect 3367 242 3371 243
rect 3367 237 3371 238
rect 3463 242 3467 243
rect 3463 237 3467 238
rect 111 230 115 231
rect 111 225 115 226
rect 167 230 171 231
rect 167 225 171 226
rect 279 230 283 231
rect 279 225 283 226
rect 343 230 347 231
rect 343 225 347 226
rect 367 230 371 231
rect 367 225 371 226
rect 463 230 467 231
rect 463 225 467 226
rect 511 230 515 231
rect 511 225 515 226
rect 559 230 563 231
rect 559 225 563 226
rect 655 230 659 231
rect 655 225 659 226
rect 679 230 683 231
rect 679 225 683 226
rect 751 230 755 231
rect 751 225 755 226
rect 839 230 843 231
rect 839 225 843 226
rect 847 230 851 231
rect 847 225 851 226
rect 943 230 947 231
rect 943 225 947 226
rect 991 230 995 231
rect 991 225 995 226
rect 1047 230 1051 231
rect 1047 225 1051 226
rect 1135 230 1139 231
rect 1135 225 1139 226
rect 1151 230 1155 231
rect 1151 225 1155 226
rect 1279 230 1283 231
rect 1279 225 1283 226
rect 1431 230 1435 231
rect 1431 225 1435 226
rect 1767 230 1771 231
rect 1767 225 1771 226
rect 112 206 114 225
rect 168 209 170 225
rect 344 209 346 225
rect 512 209 514 225
rect 680 209 682 225
rect 840 209 842 225
rect 992 209 994 225
rect 1136 209 1138 225
rect 1280 209 1282 225
rect 1432 209 1434 225
rect 166 208 172 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 166 204 167 208
rect 171 204 172 208
rect 166 203 172 204
rect 342 208 348 209
rect 342 204 343 208
rect 347 204 348 208
rect 342 203 348 204
rect 510 208 516 209
rect 510 204 511 208
rect 515 204 516 208
rect 510 203 516 204
rect 678 208 684 209
rect 678 204 679 208
rect 683 204 684 208
rect 678 203 684 204
rect 838 208 844 209
rect 838 204 839 208
rect 843 204 844 208
rect 838 203 844 204
rect 990 208 996 209
rect 990 204 991 208
rect 995 204 996 208
rect 990 203 996 204
rect 1134 208 1140 209
rect 1134 204 1135 208
rect 1139 204 1140 208
rect 1134 203 1140 204
rect 1278 208 1284 209
rect 1278 204 1279 208
rect 1283 204 1284 208
rect 1278 203 1284 204
rect 1430 208 1436 209
rect 1430 204 1431 208
rect 1435 204 1436 208
rect 1768 206 1770 225
rect 1808 218 1810 237
rect 1832 221 1834 237
rect 1928 221 1930 237
rect 2056 221 2058 237
rect 2200 221 2202 237
rect 2352 221 2354 237
rect 2512 221 2514 237
rect 2680 221 2682 237
rect 2848 221 2850 237
rect 3024 221 3026 237
rect 3208 221 3210 237
rect 3368 221 3370 237
rect 1830 220 1836 221
rect 1806 217 1812 218
rect 1806 213 1807 217
rect 1811 213 1812 217
rect 1830 216 1831 220
rect 1835 216 1836 220
rect 1830 215 1836 216
rect 1926 220 1932 221
rect 1926 216 1927 220
rect 1931 216 1932 220
rect 1926 215 1932 216
rect 2054 220 2060 221
rect 2054 216 2055 220
rect 2059 216 2060 220
rect 2054 215 2060 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2350 220 2356 221
rect 2350 216 2351 220
rect 2355 216 2356 220
rect 2350 215 2356 216
rect 2510 220 2516 221
rect 2510 216 2511 220
rect 2515 216 2516 220
rect 2510 215 2516 216
rect 2678 220 2684 221
rect 2678 216 2679 220
rect 2683 216 2684 220
rect 2678 215 2684 216
rect 2846 220 2852 221
rect 2846 216 2847 220
rect 2851 216 2852 220
rect 2846 215 2852 216
rect 3022 220 3028 221
rect 3022 216 3023 220
rect 3027 216 3028 220
rect 3022 215 3028 216
rect 3206 220 3212 221
rect 3206 216 3207 220
rect 3211 216 3212 220
rect 3206 215 3212 216
rect 3366 220 3372 221
rect 3366 216 3367 220
rect 3371 216 3372 220
rect 3464 218 3466 237
rect 3366 215 3372 216
rect 3462 217 3468 218
rect 1806 212 1812 213
rect 3462 213 3463 217
rect 3467 213 3468 217
rect 3462 212 3468 213
rect 1430 203 1436 204
rect 1766 205 1772 206
rect 110 200 116 201
rect 1766 201 1767 205
rect 1771 201 1772 205
rect 1830 201 1836 202
rect 1766 200 1772 201
rect 1806 200 1812 201
rect 1806 196 1807 200
rect 1811 196 1812 200
rect 1830 197 1831 201
rect 1835 197 1836 201
rect 1830 196 1836 197
rect 1926 201 1932 202
rect 1926 197 1927 201
rect 1931 197 1932 201
rect 1926 196 1932 197
rect 2054 201 2060 202
rect 2054 197 2055 201
rect 2059 197 2060 201
rect 2054 196 2060 197
rect 2198 201 2204 202
rect 2198 197 2199 201
rect 2203 197 2204 201
rect 2198 196 2204 197
rect 2350 201 2356 202
rect 2350 197 2351 201
rect 2355 197 2356 201
rect 2350 196 2356 197
rect 2510 201 2516 202
rect 2510 197 2511 201
rect 2515 197 2516 201
rect 2510 196 2516 197
rect 2678 201 2684 202
rect 2678 197 2679 201
rect 2683 197 2684 201
rect 2678 196 2684 197
rect 2846 201 2852 202
rect 2846 197 2847 201
rect 2851 197 2852 201
rect 2846 196 2852 197
rect 3022 201 3028 202
rect 3022 197 3023 201
rect 3027 197 3028 201
rect 3022 196 3028 197
rect 3206 201 3212 202
rect 3206 197 3207 201
rect 3211 197 3212 201
rect 3206 196 3212 197
rect 3366 201 3372 202
rect 3366 197 3367 201
rect 3371 197 3372 201
rect 3366 196 3372 197
rect 3462 200 3468 201
rect 3462 196 3463 200
rect 3467 196 3468 200
rect 1806 195 1812 196
rect 166 189 172 190
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 166 185 167 189
rect 171 185 172 189
rect 166 184 172 185
rect 342 189 348 190
rect 342 185 343 189
rect 347 185 348 189
rect 342 184 348 185
rect 510 189 516 190
rect 510 185 511 189
rect 515 185 516 189
rect 510 184 516 185
rect 678 189 684 190
rect 678 185 679 189
rect 683 185 684 189
rect 678 184 684 185
rect 838 189 844 190
rect 838 185 839 189
rect 843 185 844 189
rect 838 184 844 185
rect 990 189 996 190
rect 990 185 991 189
rect 995 185 996 189
rect 990 184 996 185
rect 1134 189 1140 190
rect 1134 185 1135 189
rect 1139 185 1140 189
rect 1134 184 1140 185
rect 1278 189 1284 190
rect 1278 185 1279 189
rect 1283 185 1284 189
rect 1278 184 1284 185
rect 1430 189 1436 190
rect 1430 185 1431 189
rect 1435 185 1436 189
rect 1430 184 1436 185
rect 1766 188 1772 189
rect 1766 184 1767 188
rect 1771 184 1772 188
rect 110 183 116 184
rect 112 143 114 183
rect 168 143 170 184
rect 344 143 346 184
rect 512 143 514 184
rect 680 143 682 184
rect 840 143 842 184
rect 992 143 994 184
rect 1136 143 1138 184
rect 1280 143 1282 184
rect 1432 143 1434 184
rect 1766 183 1772 184
rect 1768 143 1770 183
rect 1808 159 1810 195
rect 1832 159 1834 196
rect 1928 159 1930 196
rect 2056 159 2058 196
rect 2200 159 2202 196
rect 2352 159 2354 196
rect 2512 159 2514 196
rect 2680 159 2682 196
rect 2848 159 2850 196
rect 3024 159 3026 196
rect 3208 159 3210 196
rect 3368 159 3370 196
rect 3462 195 3468 196
rect 3464 159 3466 195
rect 1807 158 1811 159
rect 1807 153 1811 154
rect 1831 158 1835 159
rect 1831 153 1835 154
rect 1919 158 1923 159
rect 1919 153 1923 154
rect 1927 158 1931 159
rect 1927 153 1931 154
rect 2039 158 2043 159
rect 2039 153 2043 154
rect 2055 158 2059 159
rect 2055 153 2059 154
rect 2159 158 2163 159
rect 2159 153 2163 154
rect 2199 158 2203 159
rect 2199 153 2203 154
rect 2279 158 2283 159
rect 2279 153 2283 154
rect 2351 158 2355 159
rect 2351 153 2355 154
rect 2399 158 2403 159
rect 2399 153 2403 154
rect 2511 158 2515 159
rect 2511 153 2515 154
rect 2623 158 2627 159
rect 2623 153 2627 154
rect 2679 158 2683 159
rect 2679 153 2683 154
rect 2735 158 2739 159
rect 2735 153 2739 154
rect 2839 158 2843 159
rect 2839 153 2843 154
rect 2847 158 2851 159
rect 2847 153 2851 154
rect 2943 158 2947 159
rect 2943 153 2947 154
rect 3023 158 3027 159
rect 3023 153 3027 154
rect 3055 158 3059 159
rect 3055 153 3059 154
rect 3167 158 3171 159
rect 3167 153 3171 154
rect 3207 158 3211 159
rect 3207 153 3211 154
rect 3279 158 3283 159
rect 3279 153 3283 154
rect 3367 158 3371 159
rect 3367 153 3371 154
rect 3463 158 3467 159
rect 3463 153 3467 154
rect 111 142 115 143
rect 111 137 115 138
rect 135 142 139 143
rect 135 137 139 138
rect 167 142 171 143
rect 167 137 171 138
rect 223 142 227 143
rect 223 137 227 138
rect 311 142 315 143
rect 311 137 315 138
rect 343 142 347 143
rect 343 137 347 138
rect 399 142 403 143
rect 399 137 403 138
rect 487 142 491 143
rect 487 137 491 138
rect 511 142 515 143
rect 511 137 515 138
rect 575 142 579 143
rect 575 137 579 138
rect 663 142 667 143
rect 663 137 667 138
rect 679 142 683 143
rect 679 137 683 138
rect 751 142 755 143
rect 751 137 755 138
rect 839 142 843 143
rect 839 137 843 138
rect 847 142 851 143
rect 847 137 851 138
rect 943 142 947 143
rect 943 137 947 138
rect 991 142 995 143
rect 991 137 995 138
rect 1031 142 1035 143
rect 1031 137 1035 138
rect 1119 142 1123 143
rect 1119 137 1123 138
rect 1135 142 1139 143
rect 1135 137 1139 138
rect 1215 142 1219 143
rect 1215 137 1219 138
rect 1279 142 1283 143
rect 1279 137 1283 138
rect 1311 142 1315 143
rect 1311 137 1315 138
rect 1407 142 1411 143
rect 1407 137 1411 138
rect 1431 142 1435 143
rect 1431 137 1435 138
rect 1495 142 1499 143
rect 1495 137 1499 138
rect 1583 142 1587 143
rect 1583 137 1587 138
rect 1671 142 1675 143
rect 1671 137 1675 138
rect 1767 142 1771 143
rect 1767 137 1771 138
rect 1808 137 1810 153
rect 112 121 114 137
rect 110 120 116 121
rect 136 120 138 137
rect 224 120 226 137
rect 312 120 314 137
rect 400 120 402 137
rect 488 120 490 137
rect 576 120 578 137
rect 664 120 666 137
rect 752 120 754 137
rect 848 120 850 137
rect 944 120 946 137
rect 1032 120 1034 137
rect 1120 120 1122 137
rect 1216 120 1218 137
rect 1312 120 1314 137
rect 1408 120 1410 137
rect 1496 120 1498 137
rect 1584 120 1586 137
rect 1672 120 1674 137
rect 1768 121 1770 137
rect 1806 136 1812 137
rect 1832 136 1834 153
rect 1920 136 1922 153
rect 2040 136 2042 153
rect 2160 136 2162 153
rect 2280 136 2282 153
rect 2400 136 2402 153
rect 2512 136 2514 153
rect 2624 136 2626 153
rect 2736 136 2738 153
rect 2840 136 2842 153
rect 2944 136 2946 153
rect 3056 136 3058 153
rect 3168 136 3170 153
rect 3280 136 3282 153
rect 3368 136 3370 153
rect 3464 137 3466 153
rect 3462 136 3468 137
rect 1806 132 1807 136
rect 1811 132 1812 136
rect 1806 131 1812 132
rect 1830 135 1836 136
rect 1830 131 1831 135
rect 1835 131 1836 135
rect 1830 130 1836 131
rect 1918 135 1924 136
rect 1918 131 1919 135
rect 1923 131 1924 135
rect 1918 130 1924 131
rect 2038 135 2044 136
rect 2038 131 2039 135
rect 2043 131 2044 135
rect 2038 130 2044 131
rect 2158 135 2164 136
rect 2158 131 2159 135
rect 2163 131 2164 135
rect 2158 130 2164 131
rect 2278 135 2284 136
rect 2278 131 2279 135
rect 2283 131 2284 135
rect 2278 130 2284 131
rect 2398 135 2404 136
rect 2398 131 2399 135
rect 2403 131 2404 135
rect 2398 130 2404 131
rect 2510 135 2516 136
rect 2510 131 2511 135
rect 2515 131 2516 135
rect 2510 130 2516 131
rect 2622 135 2628 136
rect 2622 131 2623 135
rect 2627 131 2628 135
rect 2622 130 2628 131
rect 2734 135 2740 136
rect 2734 131 2735 135
rect 2739 131 2740 135
rect 2734 130 2740 131
rect 2838 135 2844 136
rect 2838 131 2839 135
rect 2843 131 2844 135
rect 2838 130 2844 131
rect 2942 135 2948 136
rect 2942 131 2943 135
rect 2947 131 2948 135
rect 2942 130 2948 131
rect 3054 135 3060 136
rect 3054 131 3055 135
rect 3059 131 3060 135
rect 3054 130 3060 131
rect 3166 135 3172 136
rect 3166 131 3167 135
rect 3171 131 3172 135
rect 3166 130 3172 131
rect 3278 135 3284 136
rect 3278 131 3279 135
rect 3283 131 3284 135
rect 3278 130 3284 131
rect 3366 135 3372 136
rect 3366 131 3367 135
rect 3371 131 3372 135
rect 3462 132 3463 136
rect 3467 132 3468 136
rect 3462 131 3468 132
rect 3366 130 3372 131
rect 1766 120 1772 121
rect 110 116 111 120
rect 115 116 116 120
rect 110 115 116 116
rect 134 119 140 120
rect 134 115 135 119
rect 139 115 140 119
rect 134 114 140 115
rect 222 119 228 120
rect 222 115 223 119
rect 227 115 228 119
rect 222 114 228 115
rect 310 119 316 120
rect 310 115 311 119
rect 315 115 316 119
rect 310 114 316 115
rect 398 119 404 120
rect 398 115 399 119
rect 403 115 404 119
rect 398 114 404 115
rect 486 119 492 120
rect 486 115 487 119
rect 491 115 492 119
rect 486 114 492 115
rect 574 119 580 120
rect 574 115 575 119
rect 579 115 580 119
rect 574 114 580 115
rect 662 119 668 120
rect 662 115 663 119
rect 667 115 668 119
rect 662 114 668 115
rect 750 119 756 120
rect 750 115 751 119
rect 755 115 756 119
rect 750 114 756 115
rect 846 119 852 120
rect 846 115 847 119
rect 851 115 852 119
rect 846 114 852 115
rect 942 119 948 120
rect 942 115 943 119
rect 947 115 948 119
rect 942 114 948 115
rect 1030 119 1036 120
rect 1030 115 1031 119
rect 1035 115 1036 119
rect 1030 114 1036 115
rect 1118 119 1124 120
rect 1118 115 1119 119
rect 1123 115 1124 119
rect 1118 114 1124 115
rect 1214 119 1220 120
rect 1214 115 1215 119
rect 1219 115 1220 119
rect 1214 114 1220 115
rect 1310 119 1316 120
rect 1310 115 1311 119
rect 1315 115 1316 119
rect 1310 114 1316 115
rect 1406 119 1412 120
rect 1406 115 1407 119
rect 1411 115 1412 119
rect 1406 114 1412 115
rect 1494 119 1500 120
rect 1494 115 1495 119
rect 1499 115 1500 119
rect 1494 114 1500 115
rect 1582 119 1588 120
rect 1582 115 1583 119
rect 1587 115 1588 119
rect 1582 114 1588 115
rect 1670 119 1676 120
rect 1670 115 1671 119
rect 1675 115 1676 119
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 119 1812 120
rect 1806 115 1807 119
rect 1811 115 1812 119
rect 3462 119 3468 120
rect 1670 114 1676 115
rect 1806 114 1812 115
rect 1830 116 1836 117
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 1766 103 1772 104
rect 110 98 116 99
rect 134 100 140 101
rect 112 79 114 98
rect 134 96 135 100
rect 139 96 140 100
rect 134 95 140 96
rect 222 100 228 101
rect 222 96 223 100
rect 227 96 228 100
rect 222 95 228 96
rect 310 100 316 101
rect 310 96 311 100
rect 315 96 316 100
rect 310 95 316 96
rect 398 100 404 101
rect 398 96 399 100
rect 403 96 404 100
rect 398 95 404 96
rect 486 100 492 101
rect 486 96 487 100
rect 491 96 492 100
rect 486 95 492 96
rect 574 100 580 101
rect 574 96 575 100
rect 579 96 580 100
rect 574 95 580 96
rect 662 100 668 101
rect 662 96 663 100
rect 667 96 668 100
rect 662 95 668 96
rect 750 100 756 101
rect 750 96 751 100
rect 755 96 756 100
rect 750 95 756 96
rect 846 100 852 101
rect 846 96 847 100
rect 851 96 852 100
rect 846 95 852 96
rect 942 100 948 101
rect 942 96 943 100
rect 947 96 948 100
rect 942 95 948 96
rect 1030 100 1036 101
rect 1030 96 1031 100
rect 1035 96 1036 100
rect 1030 95 1036 96
rect 1118 100 1124 101
rect 1118 96 1119 100
rect 1123 96 1124 100
rect 1118 95 1124 96
rect 1214 100 1220 101
rect 1214 96 1215 100
rect 1219 96 1220 100
rect 1214 95 1220 96
rect 1310 100 1316 101
rect 1310 96 1311 100
rect 1315 96 1316 100
rect 1310 95 1316 96
rect 1406 100 1412 101
rect 1406 96 1407 100
rect 1411 96 1412 100
rect 1406 95 1412 96
rect 1494 100 1500 101
rect 1494 96 1495 100
rect 1499 96 1500 100
rect 1494 95 1500 96
rect 1582 100 1588 101
rect 1582 96 1583 100
rect 1587 96 1588 100
rect 1582 95 1588 96
rect 1670 100 1676 101
rect 1670 96 1671 100
rect 1675 96 1676 100
rect 1766 99 1767 103
rect 1771 99 1772 103
rect 1766 98 1772 99
rect 1670 95 1676 96
rect 136 79 138 95
rect 224 79 226 95
rect 312 79 314 95
rect 400 79 402 95
rect 488 79 490 95
rect 576 79 578 95
rect 664 79 666 95
rect 752 79 754 95
rect 848 79 850 95
rect 944 79 946 95
rect 1032 79 1034 95
rect 1120 79 1122 95
rect 1216 79 1218 95
rect 1312 79 1314 95
rect 1408 79 1410 95
rect 1496 79 1498 95
rect 1584 79 1586 95
rect 1672 79 1674 95
rect 1768 79 1770 98
rect 1808 95 1810 114
rect 1830 112 1831 116
rect 1835 112 1836 116
rect 1830 111 1836 112
rect 1918 116 1924 117
rect 1918 112 1919 116
rect 1923 112 1924 116
rect 1918 111 1924 112
rect 2038 116 2044 117
rect 2038 112 2039 116
rect 2043 112 2044 116
rect 2038 111 2044 112
rect 2158 116 2164 117
rect 2158 112 2159 116
rect 2163 112 2164 116
rect 2158 111 2164 112
rect 2278 116 2284 117
rect 2278 112 2279 116
rect 2283 112 2284 116
rect 2278 111 2284 112
rect 2398 116 2404 117
rect 2398 112 2399 116
rect 2403 112 2404 116
rect 2398 111 2404 112
rect 2510 116 2516 117
rect 2510 112 2511 116
rect 2515 112 2516 116
rect 2510 111 2516 112
rect 2622 116 2628 117
rect 2622 112 2623 116
rect 2627 112 2628 116
rect 2622 111 2628 112
rect 2734 116 2740 117
rect 2734 112 2735 116
rect 2739 112 2740 116
rect 2734 111 2740 112
rect 2838 116 2844 117
rect 2838 112 2839 116
rect 2843 112 2844 116
rect 2838 111 2844 112
rect 2942 116 2948 117
rect 2942 112 2943 116
rect 2947 112 2948 116
rect 2942 111 2948 112
rect 3054 116 3060 117
rect 3054 112 3055 116
rect 3059 112 3060 116
rect 3054 111 3060 112
rect 3166 116 3172 117
rect 3166 112 3167 116
rect 3171 112 3172 116
rect 3166 111 3172 112
rect 3278 116 3284 117
rect 3278 112 3279 116
rect 3283 112 3284 116
rect 3278 111 3284 112
rect 3366 116 3372 117
rect 3366 112 3367 116
rect 3371 112 3372 116
rect 3462 115 3463 119
rect 3467 115 3468 119
rect 3462 114 3468 115
rect 3366 111 3372 112
rect 1832 95 1834 111
rect 1920 95 1922 111
rect 2040 95 2042 111
rect 2160 95 2162 111
rect 2280 95 2282 111
rect 2400 95 2402 111
rect 2512 95 2514 111
rect 2624 95 2626 111
rect 2736 95 2738 111
rect 2840 95 2842 111
rect 2944 95 2946 111
rect 3056 95 3058 111
rect 3168 95 3170 111
rect 3280 95 3282 111
rect 3368 95 3370 111
rect 3464 95 3466 114
rect 1807 94 1811 95
rect 1807 89 1811 90
rect 1831 94 1835 95
rect 1831 89 1835 90
rect 1919 94 1923 95
rect 1919 89 1923 90
rect 2039 94 2043 95
rect 2039 89 2043 90
rect 2159 94 2163 95
rect 2159 89 2163 90
rect 2279 94 2283 95
rect 2279 89 2283 90
rect 2399 94 2403 95
rect 2399 89 2403 90
rect 2511 94 2515 95
rect 2511 89 2515 90
rect 2623 94 2627 95
rect 2623 89 2627 90
rect 2735 94 2739 95
rect 2735 89 2739 90
rect 2839 94 2843 95
rect 2839 89 2843 90
rect 2943 94 2947 95
rect 2943 89 2947 90
rect 3055 94 3059 95
rect 3055 89 3059 90
rect 3167 94 3171 95
rect 3167 89 3171 90
rect 3279 94 3283 95
rect 3279 89 3283 90
rect 3367 94 3371 95
rect 3367 89 3371 90
rect 3463 94 3467 95
rect 3463 89 3467 90
rect 111 78 115 79
rect 111 73 115 74
rect 135 78 139 79
rect 135 73 139 74
rect 223 78 227 79
rect 223 73 227 74
rect 311 78 315 79
rect 311 73 315 74
rect 399 78 403 79
rect 399 73 403 74
rect 487 78 491 79
rect 487 73 491 74
rect 575 78 579 79
rect 575 73 579 74
rect 663 78 667 79
rect 663 73 667 74
rect 751 78 755 79
rect 751 73 755 74
rect 847 78 851 79
rect 847 73 851 74
rect 943 78 947 79
rect 943 73 947 74
rect 1031 78 1035 79
rect 1031 73 1035 74
rect 1119 78 1123 79
rect 1119 73 1123 74
rect 1215 78 1219 79
rect 1215 73 1219 74
rect 1311 78 1315 79
rect 1311 73 1315 74
rect 1407 78 1411 79
rect 1407 73 1411 74
rect 1495 78 1499 79
rect 1495 73 1499 74
rect 1583 78 1587 79
rect 1583 73 1587 74
rect 1671 78 1675 79
rect 1671 73 1675 74
rect 1767 78 1771 79
rect 1767 73 1771 74
<< m4c >>
rect 1807 3518 1811 3522
rect 2007 3518 2011 3522
rect 2239 3518 2243 3522
rect 2455 3518 2459 3522
rect 2655 3518 2659 3522
rect 2855 3518 2859 3522
rect 3047 3518 3051 3522
rect 3247 3518 3251 3522
rect 3463 3518 3467 3522
rect 111 3482 115 3486
rect 455 3482 459 3486
rect 543 3482 547 3486
rect 631 3482 635 3486
rect 719 3482 723 3486
rect 807 3482 811 3486
rect 895 3482 899 3486
rect 983 3482 987 3486
rect 1071 3482 1075 3486
rect 1159 3482 1163 3486
rect 1767 3482 1771 3486
rect 1807 3454 1811 3458
rect 1831 3454 1835 3458
rect 1943 3454 1947 3458
rect 2007 3454 2011 3458
rect 2079 3454 2083 3458
rect 2215 3454 2219 3458
rect 2239 3454 2243 3458
rect 2351 3454 2355 3458
rect 2455 3454 2459 3458
rect 2479 3454 2483 3458
rect 2599 3454 2603 3458
rect 2655 3454 2659 3458
rect 2719 3454 2723 3458
rect 2847 3454 2851 3458
rect 2855 3454 2859 3458
rect 2975 3454 2979 3458
rect 3047 3454 3051 3458
rect 3247 3454 3251 3458
rect 3463 3454 3467 3458
rect 111 3418 115 3422
rect 415 3418 419 3422
rect 455 3418 459 3422
rect 503 3418 507 3422
rect 543 3418 547 3422
rect 591 3418 595 3422
rect 631 3418 635 3422
rect 679 3418 683 3422
rect 719 3418 723 3422
rect 767 3418 771 3422
rect 807 3418 811 3422
rect 855 3418 859 3422
rect 895 3418 899 3422
rect 943 3418 947 3422
rect 983 3418 987 3422
rect 1031 3418 1035 3422
rect 1071 3418 1075 3422
rect 1119 3418 1123 3422
rect 1159 3418 1163 3422
rect 1207 3418 1211 3422
rect 1303 3418 1307 3422
rect 1767 3418 1771 3422
rect 1807 3382 1811 3386
rect 1831 3382 1835 3386
rect 1943 3382 1947 3386
rect 1951 3382 1955 3386
rect 2079 3382 2083 3386
rect 2095 3382 2099 3386
rect 2215 3382 2219 3386
rect 2239 3382 2243 3386
rect 2351 3382 2355 3386
rect 2383 3382 2387 3386
rect 2479 3382 2483 3386
rect 2519 3382 2523 3386
rect 2599 3382 2603 3386
rect 2647 3382 2651 3386
rect 2719 3382 2723 3386
rect 2775 3382 2779 3386
rect 2847 3382 2851 3386
rect 2903 3382 2907 3386
rect 2975 3382 2979 3386
rect 3039 3382 3043 3386
rect 3463 3382 3467 3386
rect 111 3350 115 3354
rect 399 3350 403 3354
rect 415 3350 419 3354
rect 495 3350 499 3354
rect 503 3350 507 3354
rect 591 3350 595 3354
rect 599 3350 603 3354
rect 679 3350 683 3354
rect 703 3350 707 3354
rect 767 3350 771 3354
rect 807 3350 811 3354
rect 855 3350 859 3354
rect 911 3350 915 3354
rect 943 3350 947 3354
rect 1015 3350 1019 3354
rect 1031 3350 1035 3354
rect 1119 3350 1123 3354
rect 1207 3350 1211 3354
rect 1223 3350 1227 3354
rect 1303 3350 1307 3354
rect 1327 3350 1331 3354
rect 1767 3350 1771 3354
rect 1807 3310 1811 3314
rect 1831 3310 1835 3314
rect 1951 3310 1955 3314
rect 1975 3310 1979 3314
rect 2095 3310 2099 3314
rect 2151 3310 2155 3314
rect 2239 3310 2243 3314
rect 2335 3310 2339 3314
rect 2383 3310 2387 3314
rect 2511 3310 2515 3314
rect 2519 3310 2523 3314
rect 2647 3310 2651 3314
rect 2679 3310 2683 3314
rect 2775 3310 2779 3314
rect 2831 3310 2835 3314
rect 2903 3310 2907 3314
rect 2975 3310 2979 3314
rect 3039 3310 3043 3314
rect 3111 3310 3115 3314
rect 3247 3310 3251 3314
rect 3367 3310 3371 3314
rect 3463 3310 3467 3314
rect 111 3282 115 3286
rect 383 3282 387 3286
rect 399 3282 403 3286
rect 495 3282 499 3286
rect 599 3282 603 3286
rect 607 3282 611 3286
rect 703 3282 707 3286
rect 727 3282 731 3286
rect 807 3282 811 3286
rect 847 3282 851 3286
rect 911 3282 915 3286
rect 967 3282 971 3286
rect 1015 3282 1019 3286
rect 1087 3282 1091 3286
rect 1119 3282 1123 3286
rect 1207 3282 1211 3286
rect 1223 3282 1227 3286
rect 1327 3282 1331 3286
rect 1335 3282 1339 3286
rect 1767 3282 1771 3286
rect 1807 3238 1811 3242
rect 1831 3238 1835 3242
rect 1975 3238 1979 3242
rect 2031 3238 2035 3242
rect 2151 3238 2155 3242
rect 2247 3238 2251 3242
rect 2335 3238 2339 3242
rect 2455 3238 2459 3242
rect 2511 3238 2515 3242
rect 2655 3238 2659 3242
rect 2679 3238 2683 3242
rect 2831 3238 2835 3242
rect 2839 3238 2843 3242
rect 2975 3238 2979 3242
rect 3023 3238 3027 3242
rect 3111 3238 3115 3242
rect 3207 3238 3211 3242
rect 3247 3238 3251 3242
rect 3367 3238 3371 3242
rect 3463 3238 3467 3242
rect 111 3214 115 3218
rect 303 3214 307 3218
rect 383 3214 387 3218
rect 423 3214 427 3218
rect 495 3214 499 3218
rect 543 3214 547 3218
rect 607 3214 611 3218
rect 671 3214 675 3218
rect 727 3214 731 3218
rect 799 3214 803 3218
rect 847 3214 851 3218
rect 927 3214 931 3218
rect 967 3214 971 3218
rect 1055 3214 1059 3218
rect 1087 3214 1091 3218
rect 1175 3214 1179 3218
rect 1207 3214 1211 3218
rect 1303 3214 1307 3218
rect 1335 3214 1339 3218
rect 1431 3214 1435 3218
rect 1767 3214 1771 3218
rect 1807 3174 1811 3178
rect 1831 3174 1835 3178
rect 1839 3174 1843 3178
rect 2031 3174 2035 3178
rect 2223 3174 2227 3178
rect 2247 3174 2251 3178
rect 2407 3174 2411 3178
rect 2455 3174 2459 3178
rect 2575 3174 2579 3178
rect 2655 3174 2659 3178
rect 2735 3174 2739 3178
rect 2839 3174 2843 3178
rect 2879 3174 2883 3178
rect 3007 3174 3011 3178
rect 3023 3174 3027 3178
rect 3135 3174 3139 3178
rect 3207 3174 3211 3178
rect 3263 3174 3267 3178
rect 3367 3174 3371 3178
rect 3463 3174 3467 3178
rect 111 3138 115 3142
rect 175 3138 179 3142
rect 303 3138 307 3142
rect 319 3138 323 3142
rect 423 3138 427 3142
rect 471 3138 475 3142
rect 543 3138 547 3142
rect 623 3138 627 3142
rect 671 3138 675 3142
rect 775 3138 779 3142
rect 799 3138 803 3142
rect 919 3138 923 3142
rect 927 3138 931 3142
rect 1055 3138 1059 3142
rect 1063 3138 1067 3142
rect 1175 3138 1179 3142
rect 1199 3138 1203 3142
rect 1303 3138 1307 3142
rect 1343 3138 1347 3142
rect 1431 3138 1435 3142
rect 1487 3138 1491 3142
rect 1767 3138 1771 3142
rect 1807 3106 1811 3110
rect 1839 3106 1843 3110
rect 1935 3106 1939 3110
rect 2031 3106 2035 3110
rect 2055 3106 2059 3110
rect 2175 3106 2179 3110
rect 2223 3106 2227 3110
rect 2303 3106 2307 3110
rect 2407 3106 2411 3110
rect 2431 3106 2435 3110
rect 2567 3106 2571 3110
rect 2575 3106 2579 3110
rect 2719 3106 2723 3110
rect 2735 3106 2739 3110
rect 2871 3106 2875 3110
rect 2879 3106 2883 3110
rect 3007 3106 3011 3110
rect 3031 3106 3035 3110
rect 3135 3106 3139 3110
rect 3199 3106 3203 3110
rect 3263 3106 3267 3110
rect 3367 3106 3371 3110
rect 3463 3106 3467 3110
rect 111 3066 115 3070
rect 135 3066 139 3070
rect 175 3066 179 3070
rect 263 3066 267 3070
rect 319 3066 323 3070
rect 431 3066 435 3070
rect 471 3066 475 3070
rect 607 3066 611 3070
rect 623 3066 627 3070
rect 775 3066 779 3070
rect 791 3066 795 3070
rect 919 3066 923 3070
rect 967 3066 971 3070
rect 1063 3066 1067 3070
rect 1143 3066 1147 3070
rect 1199 3066 1203 3070
rect 1327 3066 1331 3070
rect 1343 3066 1347 3070
rect 1487 3066 1491 3070
rect 1511 3066 1515 3070
rect 1767 3066 1771 3070
rect 1807 3034 1811 3038
rect 1935 3034 1939 3038
rect 2023 3034 2027 3038
rect 2055 3034 2059 3038
rect 2127 3034 2131 3038
rect 2175 3034 2179 3038
rect 2231 3034 2235 3038
rect 2303 3034 2307 3038
rect 2335 3034 2339 3038
rect 2431 3034 2435 3038
rect 2439 3034 2443 3038
rect 2543 3034 2547 3038
rect 2567 3034 2571 3038
rect 2647 3034 2651 3038
rect 2719 3034 2723 3038
rect 2759 3034 2763 3038
rect 2871 3034 2875 3038
rect 3031 3034 3035 3038
rect 3199 3034 3203 3038
rect 3367 3034 3371 3038
rect 3463 3034 3467 3038
rect 111 2998 115 3002
rect 135 2998 139 3002
rect 263 2998 267 3002
rect 327 2998 331 3002
rect 431 2998 435 3002
rect 535 2998 539 3002
rect 607 2998 611 3002
rect 735 2998 739 3002
rect 791 2998 795 3002
rect 927 2998 931 3002
rect 967 2998 971 3002
rect 1103 2998 1107 3002
rect 1143 2998 1147 3002
rect 1279 2998 1283 3002
rect 1327 2998 1331 3002
rect 1447 2998 1451 3002
rect 1511 2998 1515 3002
rect 1623 2998 1627 3002
rect 1767 2998 1771 3002
rect 1807 2970 1811 2974
rect 2023 2970 2027 2974
rect 2055 2970 2059 2974
rect 2127 2970 2131 2974
rect 2143 2970 2147 2974
rect 2231 2970 2235 2974
rect 2319 2970 2323 2974
rect 2335 2970 2339 2974
rect 2407 2970 2411 2974
rect 2439 2970 2443 2974
rect 2495 2970 2499 2974
rect 2543 2970 2547 2974
rect 2583 2970 2587 2974
rect 2647 2970 2651 2974
rect 2671 2970 2675 2974
rect 2759 2970 2763 2974
rect 2847 2970 2851 2974
rect 3463 2970 3467 2974
rect 111 2926 115 2930
rect 135 2926 139 2930
rect 263 2926 267 2930
rect 327 2926 331 2930
rect 431 2926 435 2930
rect 535 2926 539 2930
rect 607 2926 611 2930
rect 735 2926 739 2930
rect 783 2926 787 2930
rect 927 2926 931 2930
rect 951 2926 955 2930
rect 1103 2926 1107 2930
rect 1111 2926 1115 2930
rect 1271 2926 1275 2930
rect 1279 2926 1283 2930
rect 1431 2926 1435 2930
rect 1447 2926 1451 2930
rect 1591 2926 1595 2930
rect 1623 2926 1627 2930
rect 1767 2926 1771 2930
rect 1807 2898 1811 2902
rect 2055 2898 2059 2902
rect 2071 2898 2075 2902
rect 2143 2898 2147 2902
rect 2175 2898 2179 2902
rect 2231 2898 2235 2902
rect 2271 2898 2275 2902
rect 2319 2898 2323 2902
rect 2367 2898 2371 2902
rect 2407 2898 2411 2902
rect 2471 2898 2475 2902
rect 2495 2898 2499 2902
rect 2575 2898 2579 2902
rect 2583 2898 2587 2902
rect 2671 2898 2675 2902
rect 2679 2898 2683 2902
rect 2759 2898 2763 2902
rect 2783 2898 2787 2902
rect 2847 2898 2851 2902
rect 3463 2898 3467 2902
rect 111 2858 115 2862
rect 135 2858 139 2862
rect 255 2858 259 2862
rect 263 2858 267 2862
rect 407 2858 411 2862
rect 431 2858 435 2862
rect 567 2858 571 2862
rect 607 2858 611 2862
rect 727 2858 731 2862
rect 783 2858 787 2862
rect 879 2858 883 2862
rect 951 2858 955 2862
rect 1023 2858 1027 2862
rect 1111 2858 1115 2862
rect 1167 2858 1171 2862
rect 1271 2858 1275 2862
rect 1311 2858 1315 2862
rect 1431 2858 1435 2862
rect 1463 2858 1467 2862
rect 1591 2858 1595 2862
rect 1767 2858 1771 2862
rect 1807 2830 1811 2834
rect 1983 2830 1987 2834
rect 2071 2830 2075 2834
rect 2111 2830 2115 2834
rect 2175 2830 2179 2834
rect 2239 2830 2243 2834
rect 2271 2830 2275 2834
rect 2367 2830 2371 2834
rect 2471 2830 2475 2834
rect 2487 2830 2491 2834
rect 2575 2830 2579 2834
rect 2607 2830 2611 2834
rect 2679 2830 2683 2834
rect 2719 2830 2723 2834
rect 2783 2830 2787 2834
rect 2839 2830 2843 2834
rect 2959 2830 2963 2834
rect 3463 2830 3467 2834
rect 111 2786 115 2790
rect 135 2786 139 2790
rect 255 2786 259 2790
rect 287 2786 291 2790
rect 391 2786 395 2790
rect 407 2786 411 2790
rect 503 2786 507 2790
rect 567 2786 571 2790
rect 623 2786 627 2790
rect 727 2786 731 2790
rect 743 2786 747 2790
rect 855 2786 859 2790
rect 879 2786 883 2790
rect 967 2786 971 2790
rect 1023 2786 1027 2790
rect 1079 2786 1083 2790
rect 1167 2786 1171 2790
rect 1199 2786 1203 2790
rect 1311 2786 1315 2790
rect 1319 2786 1323 2790
rect 1463 2786 1467 2790
rect 1767 2786 1771 2790
rect 1807 2762 1811 2766
rect 1887 2762 1891 2766
rect 1983 2762 1987 2766
rect 2031 2762 2035 2766
rect 2111 2762 2115 2766
rect 2183 2762 2187 2766
rect 2239 2762 2243 2766
rect 2335 2762 2339 2766
rect 2367 2762 2371 2766
rect 2479 2762 2483 2766
rect 2487 2762 2491 2766
rect 2607 2762 2611 2766
rect 2623 2762 2627 2766
rect 2719 2762 2723 2766
rect 2767 2762 2771 2766
rect 2839 2762 2843 2766
rect 2911 2762 2915 2766
rect 2959 2762 2963 2766
rect 3055 2762 3059 2766
rect 3463 2762 3467 2766
rect 111 2718 115 2722
rect 287 2718 291 2722
rect 391 2718 395 2722
rect 479 2718 483 2722
rect 503 2718 507 2722
rect 567 2718 571 2722
rect 623 2718 627 2722
rect 655 2718 659 2722
rect 743 2718 747 2722
rect 831 2718 835 2722
rect 855 2718 859 2722
rect 919 2718 923 2722
rect 967 2718 971 2722
rect 1007 2718 1011 2722
rect 1079 2718 1083 2722
rect 1095 2718 1099 2722
rect 1183 2718 1187 2722
rect 1199 2718 1203 2722
rect 1319 2718 1323 2722
rect 1767 2718 1771 2722
rect 1807 2698 1811 2702
rect 1831 2698 1835 2702
rect 1887 2698 1891 2702
rect 2023 2698 2027 2702
rect 2031 2698 2035 2702
rect 2183 2698 2187 2702
rect 2231 2698 2235 2702
rect 2335 2698 2339 2702
rect 2431 2698 2435 2702
rect 2479 2698 2483 2702
rect 2615 2698 2619 2702
rect 2623 2698 2627 2702
rect 2767 2698 2771 2702
rect 2783 2698 2787 2702
rect 2911 2698 2915 2702
rect 2943 2698 2947 2702
rect 3055 2698 3059 2702
rect 3095 2698 3099 2702
rect 3239 2698 3243 2702
rect 3367 2698 3371 2702
rect 3463 2698 3467 2702
rect 111 2646 115 2650
rect 471 2646 475 2650
rect 479 2646 483 2650
rect 559 2646 563 2650
rect 567 2646 571 2650
rect 647 2646 651 2650
rect 655 2646 659 2650
rect 735 2646 739 2650
rect 743 2646 747 2650
rect 823 2646 827 2650
rect 831 2646 835 2650
rect 911 2646 915 2650
rect 919 2646 923 2650
rect 999 2646 1003 2650
rect 1007 2646 1011 2650
rect 1087 2646 1091 2650
rect 1095 2646 1099 2650
rect 1183 2646 1187 2650
rect 1767 2646 1771 2650
rect 1807 2630 1811 2634
rect 1831 2630 1835 2634
rect 1999 2630 2003 2634
rect 2023 2630 2027 2634
rect 2183 2630 2187 2634
rect 2231 2630 2235 2634
rect 2359 2630 2363 2634
rect 2431 2630 2435 2634
rect 2519 2630 2523 2634
rect 2615 2630 2619 2634
rect 2671 2630 2675 2634
rect 2783 2630 2787 2634
rect 2807 2630 2811 2634
rect 2927 2630 2931 2634
rect 2943 2630 2947 2634
rect 3047 2630 3051 2634
rect 3095 2630 3099 2634
rect 3159 2630 3163 2634
rect 3239 2630 3243 2634
rect 3271 2630 3275 2634
rect 3367 2630 3371 2634
rect 3463 2630 3467 2634
rect 111 2570 115 2574
rect 223 2570 227 2574
rect 311 2570 315 2574
rect 407 2570 411 2574
rect 471 2570 475 2574
rect 503 2570 507 2574
rect 559 2570 563 2574
rect 591 2570 595 2574
rect 647 2570 651 2574
rect 679 2570 683 2574
rect 735 2570 739 2574
rect 767 2570 771 2574
rect 823 2570 827 2574
rect 855 2570 859 2574
rect 911 2570 915 2574
rect 943 2570 947 2574
rect 999 2570 1003 2574
rect 1031 2570 1035 2574
rect 1087 2570 1091 2574
rect 1119 2570 1123 2574
rect 1215 2570 1219 2574
rect 1311 2570 1315 2574
rect 1407 2570 1411 2574
rect 1495 2570 1499 2574
rect 1583 2570 1587 2574
rect 1671 2570 1675 2574
rect 1767 2570 1771 2574
rect 1807 2558 1811 2562
rect 1831 2558 1835 2562
rect 1999 2558 2003 2562
rect 2183 2558 2187 2562
rect 2207 2558 2211 2562
rect 2359 2558 2363 2562
rect 2519 2558 2523 2562
rect 2671 2558 2675 2562
rect 2799 2558 2803 2562
rect 2807 2558 2811 2562
rect 2927 2558 2931 2562
rect 3047 2558 3051 2562
rect 3159 2558 3163 2562
rect 3271 2558 3275 2562
rect 3367 2558 3371 2562
rect 3463 2558 3467 2562
rect 111 2506 115 2510
rect 135 2506 139 2510
rect 223 2506 227 2510
rect 247 2506 251 2510
rect 311 2506 315 2510
rect 391 2506 395 2510
rect 407 2506 411 2510
rect 503 2506 507 2510
rect 543 2506 547 2510
rect 591 2506 595 2510
rect 679 2506 683 2510
rect 695 2506 699 2510
rect 767 2506 771 2510
rect 839 2506 843 2510
rect 855 2506 859 2510
rect 943 2506 947 2510
rect 975 2506 979 2510
rect 1031 2506 1035 2510
rect 1103 2506 1107 2510
rect 1119 2506 1123 2510
rect 1215 2506 1219 2510
rect 1231 2506 1235 2510
rect 1311 2506 1315 2510
rect 1351 2506 1355 2510
rect 1407 2506 1411 2510
rect 1463 2506 1467 2510
rect 1495 2506 1499 2510
rect 1575 2506 1579 2510
rect 1583 2506 1587 2510
rect 1671 2506 1675 2510
rect 1767 2506 1771 2510
rect 1807 2478 1811 2482
rect 2015 2478 2019 2482
rect 2199 2478 2203 2482
rect 2207 2478 2211 2482
rect 2367 2478 2371 2482
rect 2527 2478 2531 2482
rect 2671 2478 2675 2482
rect 2799 2478 2803 2482
rect 2807 2478 2811 2482
rect 2927 2478 2931 2482
rect 3047 2478 3051 2482
rect 3159 2478 3163 2482
rect 3271 2478 3275 2482
rect 3367 2478 3371 2482
rect 3463 2478 3467 2482
rect 111 2426 115 2430
rect 135 2426 139 2430
rect 239 2426 243 2430
rect 247 2426 251 2430
rect 391 2426 395 2430
rect 543 2426 547 2430
rect 551 2426 555 2430
rect 695 2426 699 2430
rect 719 2426 723 2430
rect 839 2426 843 2430
rect 895 2426 899 2430
rect 975 2426 979 2430
rect 1063 2426 1067 2430
rect 1103 2426 1107 2430
rect 1231 2426 1235 2430
rect 1239 2426 1243 2430
rect 1351 2426 1355 2430
rect 1415 2426 1419 2430
rect 1463 2426 1467 2430
rect 1575 2426 1579 2430
rect 1591 2426 1595 2430
rect 1671 2426 1675 2430
rect 1767 2426 1771 2430
rect 1807 2410 1811 2414
rect 1839 2410 1843 2414
rect 2007 2410 2011 2414
rect 2015 2410 2019 2414
rect 2183 2410 2187 2414
rect 2199 2410 2203 2414
rect 2367 2410 2371 2414
rect 2527 2410 2531 2414
rect 2559 2410 2563 2414
rect 2671 2410 2675 2414
rect 2759 2410 2763 2414
rect 2807 2410 2811 2414
rect 2927 2410 2931 2414
rect 2967 2410 2971 2414
rect 3047 2410 3051 2414
rect 3159 2410 3163 2414
rect 3175 2410 3179 2414
rect 3271 2410 3275 2414
rect 3367 2410 3371 2414
rect 3463 2410 3467 2414
rect 111 2354 115 2358
rect 135 2354 139 2358
rect 239 2354 243 2358
rect 375 2354 379 2358
rect 391 2354 395 2358
rect 479 2354 483 2358
rect 551 2354 555 2358
rect 599 2354 603 2358
rect 719 2354 723 2358
rect 847 2354 851 2358
rect 895 2354 899 2358
rect 975 2354 979 2358
rect 1063 2354 1067 2358
rect 1103 2354 1107 2358
rect 1239 2354 1243 2358
rect 1375 2354 1379 2358
rect 1415 2354 1419 2358
rect 1511 2354 1515 2358
rect 1591 2354 1595 2358
rect 1767 2354 1771 2358
rect 1807 2346 1811 2350
rect 1839 2346 1843 2350
rect 1887 2346 1891 2350
rect 2007 2346 2011 2350
rect 2015 2346 2019 2350
rect 2151 2346 2155 2350
rect 2183 2346 2187 2350
rect 2303 2346 2307 2350
rect 2367 2346 2371 2350
rect 2463 2346 2467 2350
rect 2559 2346 2563 2350
rect 2647 2346 2651 2350
rect 2759 2346 2763 2350
rect 2839 2346 2843 2350
rect 2967 2346 2971 2350
rect 3047 2346 3051 2350
rect 3175 2346 3179 2350
rect 3255 2346 3259 2350
rect 3367 2346 3371 2350
rect 3463 2346 3467 2350
rect 111 2282 115 2286
rect 375 2282 379 2286
rect 479 2282 483 2286
rect 575 2282 579 2286
rect 599 2282 603 2286
rect 663 2282 667 2286
rect 719 2282 723 2286
rect 759 2282 763 2286
rect 847 2282 851 2286
rect 863 2282 867 2286
rect 967 2282 971 2286
rect 975 2282 979 2286
rect 1079 2282 1083 2286
rect 1103 2282 1107 2286
rect 1191 2282 1195 2286
rect 1239 2282 1243 2286
rect 1303 2282 1307 2286
rect 1375 2282 1379 2286
rect 1415 2282 1419 2286
rect 1511 2282 1515 2286
rect 1767 2282 1771 2286
rect 1807 2278 1811 2282
rect 1887 2278 1891 2282
rect 2015 2278 2019 2282
rect 2039 2278 2043 2282
rect 2135 2278 2139 2282
rect 2151 2278 2155 2282
rect 2239 2278 2243 2282
rect 2303 2278 2307 2282
rect 2343 2278 2347 2282
rect 2463 2278 2467 2282
rect 2591 2278 2595 2282
rect 2647 2278 2651 2282
rect 2735 2278 2739 2282
rect 2839 2278 2843 2282
rect 2887 2278 2891 2282
rect 3047 2278 3051 2282
rect 3215 2278 3219 2282
rect 3255 2278 3259 2282
rect 3367 2278 3371 2282
rect 3463 2278 3467 2282
rect 111 2218 115 2222
rect 439 2218 443 2222
rect 527 2218 531 2222
rect 575 2218 579 2222
rect 615 2218 619 2222
rect 663 2218 667 2222
rect 703 2218 707 2222
rect 759 2218 763 2222
rect 791 2218 795 2222
rect 863 2218 867 2222
rect 879 2218 883 2222
rect 967 2218 971 2222
rect 1055 2218 1059 2222
rect 1079 2218 1083 2222
rect 1143 2218 1147 2222
rect 1191 2218 1195 2222
rect 1231 2218 1235 2222
rect 1303 2218 1307 2222
rect 1319 2218 1323 2222
rect 1415 2218 1419 2222
rect 1767 2218 1771 2222
rect 1807 2202 1811 2206
rect 2039 2202 2043 2206
rect 2135 2202 2139 2206
rect 2183 2202 2187 2206
rect 2239 2202 2243 2206
rect 2279 2202 2283 2206
rect 2343 2202 2347 2206
rect 2383 2202 2387 2206
rect 2463 2202 2467 2206
rect 2495 2202 2499 2206
rect 2591 2202 2595 2206
rect 2607 2202 2611 2206
rect 2719 2202 2723 2206
rect 2735 2202 2739 2206
rect 2839 2202 2843 2206
rect 2887 2202 2891 2206
rect 2967 2202 2971 2206
rect 3047 2202 3051 2206
rect 3103 2202 3107 2206
rect 3215 2202 3219 2206
rect 3247 2202 3251 2206
rect 3367 2202 3371 2206
rect 3463 2202 3467 2206
rect 111 2138 115 2142
rect 303 2138 307 2142
rect 407 2138 411 2142
rect 439 2138 443 2142
rect 519 2138 523 2142
rect 527 2138 531 2142
rect 615 2138 619 2142
rect 631 2138 635 2142
rect 703 2138 707 2142
rect 743 2138 747 2142
rect 791 2138 795 2142
rect 863 2138 867 2142
rect 879 2138 883 2142
rect 967 2138 971 2142
rect 983 2138 987 2142
rect 1055 2138 1059 2142
rect 1143 2138 1147 2142
rect 1231 2138 1235 2142
rect 1319 2138 1323 2142
rect 1767 2138 1771 2142
rect 1807 2130 1811 2134
rect 2135 2130 2139 2134
rect 2183 2130 2187 2134
rect 2255 2130 2259 2134
rect 2279 2130 2283 2134
rect 2383 2130 2387 2134
rect 2495 2130 2499 2134
rect 2519 2130 2523 2134
rect 2607 2130 2611 2134
rect 2655 2130 2659 2134
rect 2719 2130 2723 2134
rect 2783 2130 2787 2134
rect 2839 2130 2843 2134
rect 2911 2130 2915 2134
rect 2967 2130 2971 2134
rect 3031 2130 3035 2134
rect 3103 2130 3107 2134
rect 3151 2130 3155 2134
rect 3247 2130 3251 2134
rect 3271 2130 3275 2134
rect 3367 2130 3371 2134
rect 3463 2130 3467 2134
rect 111 2074 115 2078
rect 255 2074 259 2078
rect 303 2074 307 2078
rect 375 2074 379 2078
rect 407 2074 411 2078
rect 495 2074 499 2078
rect 519 2074 523 2078
rect 615 2074 619 2078
rect 631 2074 635 2078
rect 727 2074 731 2078
rect 743 2074 747 2078
rect 831 2074 835 2078
rect 863 2074 867 2078
rect 935 2074 939 2078
rect 983 2074 987 2078
rect 1039 2074 1043 2078
rect 1143 2074 1147 2078
rect 1255 2074 1259 2078
rect 1767 2074 1771 2078
rect 1807 2058 1811 2062
rect 2135 2058 2139 2062
rect 2247 2058 2251 2062
rect 2255 2058 2259 2062
rect 2383 2058 2387 2062
rect 2415 2058 2419 2062
rect 2519 2058 2523 2062
rect 2575 2058 2579 2062
rect 2655 2058 2659 2062
rect 2727 2058 2731 2062
rect 2783 2058 2787 2062
rect 2871 2058 2875 2062
rect 2911 2058 2915 2062
rect 3007 2058 3011 2062
rect 3031 2058 3035 2062
rect 3135 2058 3139 2062
rect 3151 2058 3155 2062
rect 3263 2058 3267 2062
rect 3271 2058 3275 2062
rect 3367 2058 3371 2062
rect 3463 2058 3467 2062
rect 111 2010 115 2014
rect 255 2010 259 2014
rect 359 2010 363 2014
rect 375 2010 379 2014
rect 487 2010 491 2014
rect 495 2010 499 2014
rect 615 2010 619 2014
rect 623 2010 627 2014
rect 727 2010 731 2014
rect 759 2010 763 2014
rect 831 2010 835 2014
rect 895 2010 899 2014
rect 935 2010 939 2014
rect 1023 2010 1027 2014
rect 1039 2010 1043 2014
rect 1143 2010 1147 2014
rect 1151 2010 1155 2014
rect 1255 2010 1259 2014
rect 1271 2010 1275 2014
rect 1399 2010 1403 2014
rect 1527 2010 1531 2014
rect 1767 2010 1771 2014
rect 1807 1978 1811 1982
rect 1831 1978 1835 1982
rect 1919 1978 1923 1982
rect 2047 1978 2051 1982
rect 2183 1978 2187 1982
rect 2247 1978 2251 1982
rect 2327 1978 2331 1982
rect 2415 1978 2419 1982
rect 2471 1978 2475 1982
rect 2575 1978 2579 1982
rect 2615 1978 2619 1982
rect 2727 1978 2731 1982
rect 2751 1978 2755 1982
rect 2871 1978 2875 1982
rect 2887 1978 2891 1982
rect 3007 1978 3011 1982
rect 3031 1978 3035 1982
rect 3135 1978 3139 1982
rect 3175 1978 3179 1982
rect 3263 1978 3267 1982
rect 3319 1978 3323 1982
rect 3367 1978 3371 1982
rect 3463 1978 3467 1982
rect 111 1946 115 1950
rect 359 1946 363 1950
rect 447 1946 451 1950
rect 487 1946 491 1950
rect 575 1946 579 1950
rect 623 1946 627 1950
rect 711 1946 715 1950
rect 759 1946 763 1950
rect 847 1946 851 1950
rect 895 1946 899 1950
rect 983 1946 987 1950
rect 1023 1946 1027 1950
rect 1119 1946 1123 1950
rect 1151 1946 1155 1950
rect 1255 1946 1259 1950
rect 1271 1946 1275 1950
rect 1383 1946 1387 1950
rect 1399 1946 1403 1950
rect 1519 1946 1523 1950
rect 1527 1946 1531 1950
rect 1655 1946 1659 1950
rect 1767 1946 1771 1950
rect 1807 1910 1811 1914
rect 1831 1910 1835 1914
rect 1919 1910 1923 1914
rect 2039 1910 2043 1914
rect 2047 1910 2051 1914
rect 2167 1910 2171 1914
rect 2183 1910 2187 1914
rect 2303 1910 2307 1914
rect 2327 1910 2331 1914
rect 2455 1910 2459 1914
rect 2471 1910 2475 1914
rect 2615 1910 2619 1914
rect 2751 1910 2755 1914
rect 2791 1910 2795 1914
rect 2887 1910 2891 1914
rect 2983 1910 2987 1914
rect 3031 1910 3035 1914
rect 3175 1910 3179 1914
rect 3183 1910 3187 1914
rect 3319 1910 3323 1914
rect 3367 1910 3371 1914
rect 3463 1910 3467 1914
rect 111 1882 115 1886
rect 447 1882 451 1886
rect 559 1882 563 1886
rect 575 1882 579 1886
rect 695 1882 699 1886
rect 711 1882 715 1886
rect 831 1882 835 1886
rect 847 1882 851 1886
rect 959 1882 963 1886
rect 983 1882 987 1886
rect 1079 1882 1083 1886
rect 1119 1882 1123 1886
rect 1199 1882 1203 1886
rect 1255 1882 1259 1886
rect 1327 1882 1331 1886
rect 1383 1882 1387 1886
rect 1455 1882 1459 1886
rect 1519 1882 1523 1886
rect 1655 1882 1659 1886
rect 1767 1882 1771 1886
rect 1807 1842 1811 1846
rect 1831 1842 1835 1846
rect 1919 1842 1923 1846
rect 1959 1842 1963 1846
rect 2039 1842 2043 1846
rect 2111 1842 2115 1846
rect 2167 1842 2171 1846
rect 2255 1842 2259 1846
rect 2303 1842 2307 1846
rect 2407 1842 2411 1846
rect 2455 1842 2459 1846
rect 2567 1842 2571 1846
rect 2615 1842 2619 1846
rect 2743 1842 2747 1846
rect 2791 1842 2795 1846
rect 2935 1842 2939 1846
rect 2983 1842 2987 1846
rect 3135 1842 3139 1846
rect 3183 1842 3187 1846
rect 3343 1842 3347 1846
rect 3367 1842 3371 1846
rect 3463 1842 3467 1846
rect 111 1810 115 1814
rect 135 1810 139 1814
rect 223 1810 227 1814
rect 311 1810 315 1814
rect 407 1810 411 1814
rect 527 1810 531 1814
rect 559 1810 563 1814
rect 655 1810 659 1814
rect 695 1810 699 1814
rect 799 1810 803 1814
rect 831 1810 835 1814
rect 943 1810 947 1814
rect 959 1810 963 1814
rect 1079 1810 1083 1814
rect 1087 1810 1091 1814
rect 1199 1810 1203 1814
rect 1239 1810 1243 1814
rect 1327 1810 1331 1814
rect 1391 1810 1395 1814
rect 1455 1810 1459 1814
rect 1543 1810 1547 1814
rect 1671 1810 1675 1814
rect 1767 1810 1771 1814
rect 1807 1766 1811 1770
rect 1831 1766 1835 1770
rect 1879 1766 1883 1770
rect 1959 1766 1963 1770
rect 2015 1766 2019 1770
rect 2111 1766 2115 1770
rect 2151 1766 2155 1770
rect 2255 1766 2259 1770
rect 2303 1766 2307 1770
rect 2407 1766 2411 1770
rect 2479 1766 2483 1770
rect 2567 1766 2571 1770
rect 2687 1766 2691 1770
rect 2743 1766 2747 1770
rect 2911 1766 2915 1770
rect 2935 1766 2939 1770
rect 3135 1766 3139 1770
rect 3151 1766 3155 1770
rect 3343 1766 3347 1770
rect 3367 1766 3371 1770
rect 3463 1766 3467 1770
rect 111 1734 115 1738
rect 135 1734 139 1738
rect 223 1734 227 1738
rect 247 1734 251 1738
rect 311 1734 315 1738
rect 399 1734 403 1738
rect 407 1734 411 1738
rect 527 1734 531 1738
rect 567 1734 571 1738
rect 655 1734 659 1738
rect 751 1734 755 1738
rect 799 1734 803 1738
rect 935 1734 939 1738
rect 943 1734 947 1738
rect 1087 1734 1091 1738
rect 1119 1734 1123 1738
rect 1239 1734 1243 1738
rect 1311 1734 1315 1738
rect 1391 1734 1395 1738
rect 1503 1734 1507 1738
rect 1543 1734 1547 1738
rect 1671 1734 1675 1738
rect 1767 1734 1771 1738
rect 1807 1694 1811 1698
rect 1831 1694 1835 1698
rect 1879 1694 1883 1698
rect 1935 1694 1939 1698
rect 2015 1694 2019 1698
rect 2063 1694 2067 1698
rect 2151 1694 2155 1698
rect 2183 1694 2187 1698
rect 2303 1694 2307 1698
rect 2311 1694 2315 1698
rect 2439 1694 2443 1698
rect 2479 1694 2483 1698
rect 2575 1694 2579 1698
rect 2687 1694 2691 1698
rect 2727 1694 2731 1698
rect 2887 1694 2891 1698
rect 2911 1694 2915 1698
rect 3047 1694 3051 1698
rect 3151 1694 3155 1698
rect 3215 1694 3219 1698
rect 3367 1694 3371 1698
rect 3463 1694 3467 1698
rect 111 1666 115 1670
rect 135 1666 139 1670
rect 191 1666 195 1670
rect 247 1666 251 1670
rect 295 1666 299 1670
rect 399 1666 403 1670
rect 407 1666 411 1670
rect 535 1666 539 1670
rect 567 1666 571 1670
rect 687 1666 691 1670
rect 751 1666 755 1670
rect 855 1666 859 1670
rect 935 1666 939 1670
rect 1039 1666 1043 1670
rect 1119 1666 1123 1670
rect 1231 1666 1235 1670
rect 1311 1666 1315 1670
rect 1431 1666 1435 1670
rect 1503 1666 1507 1670
rect 1639 1666 1643 1670
rect 1671 1666 1675 1670
rect 1767 1666 1771 1670
rect 1807 1622 1811 1626
rect 1831 1622 1835 1626
rect 1935 1622 1939 1626
rect 1943 1622 1947 1626
rect 2063 1622 2067 1626
rect 2087 1622 2091 1626
rect 2183 1622 2187 1626
rect 2231 1622 2235 1626
rect 2311 1622 2315 1626
rect 2367 1622 2371 1626
rect 2439 1622 2443 1626
rect 2503 1622 2507 1626
rect 2575 1622 2579 1626
rect 2639 1622 2643 1626
rect 2727 1622 2731 1626
rect 2767 1622 2771 1626
rect 2887 1622 2891 1626
rect 2895 1622 2899 1626
rect 3015 1622 3019 1626
rect 3047 1622 3051 1626
rect 3135 1622 3139 1626
rect 3215 1622 3219 1626
rect 3263 1622 3267 1626
rect 3367 1622 3371 1626
rect 3463 1622 3467 1626
rect 111 1598 115 1602
rect 191 1598 195 1602
rect 295 1598 299 1602
rect 327 1598 331 1602
rect 407 1598 411 1602
rect 431 1598 435 1602
rect 535 1598 539 1602
rect 543 1598 547 1602
rect 671 1598 675 1602
rect 687 1598 691 1602
rect 815 1598 819 1602
rect 855 1598 859 1602
rect 967 1598 971 1602
rect 1039 1598 1043 1602
rect 1119 1598 1123 1602
rect 1231 1598 1235 1602
rect 1279 1598 1283 1602
rect 1431 1598 1435 1602
rect 1439 1598 1443 1602
rect 1607 1598 1611 1602
rect 1639 1598 1643 1602
rect 1767 1598 1771 1602
rect 1807 1550 1811 1554
rect 1831 1550 1835 1554
rect 1839 1550 1843 1554
rect 1943 1550 1947 1554
rect 1991 1550 1995 1554
rect 2087 1550 2091 1554
rect 2151 1550 2155 1554
rect 2231 1550 2235 1554
rect 2303 1550 2307 1554
rect 2367 1550 2371 1554
rect 2455 1550 2459 1554
rect 2503 1550 2507 1554
rect 2599 1550 2603 1554
rect 2639 1550 2643 1554
rect 2735 1550 2739 1554
rect 2767 1550 2771 1554
rect 2871 1550 2875 1554
rect 2895 1550 2899 1554
rect 3007 1550 3011 1554
rect 3015 1550 3019 1554
rect 3135 1550 3139 1554
rect 3143 1550 3147 1554
rect 3263 1550 3267 1554
rect 3367 1550 3371 1554
rect 3463 1550 3467 1554
rect 111 1530 115 1534
rect 223 1530 227 1534
rect 327 1530 331 1534
rect 343 1530 347 1534
rect 431 1530 435 1534
rect 471 1530 475 1534
rect 543 1530 547 1534
rect 607 1530 611 1534
rect 671 1530 675 1534
rect 751 1530 755 1534
rect 815 1530 819 1534
rect 895 1530 899 1534
rect 967 1530 971 1534
rect 1047 1530 1051 1534
rect 1119 1530 1123 1534
rect 1199 1530 1203 1534
rect 1279 1530 1283 1534
rect 1351 1530 1355 1534
rect 1439 1530 1443 1534
rect 1503 1530 1507 1534
rect 1607 1530 1611 1534
rect 1767 1530 1771 1534
rect 1807 1478 1811 1482
rect 1839 1478 1843 1482
rect 1943 1478 1947 1482
rect 1991 1478 1995 1482
rect 2055 1478 2059 1482
rect 2151 1478 2155 1482
rect 2191 1478 2195 1482
rect 2303 1478 2307 1482
rect 2335 1478 2339 1482
rect 2455 1478 2459 1482
rect 2479 1478 2483 1482
rect 2599 1478 2603 1482
rect 2631 1478 2635 1482
rect 2735 1478 2739 1482
rect 2783 1478 2787 1482
rect 2871 1478 2875 1482
rect 2935 1478 2939 1482
rect 3007 1478 3011 1482
rect 3087 1478 3091 1482
rect 3143 1478 3147 1482
rect 3239 1478 3243 1482
rect 3463 1478 3467 1482
rect 111 1458 115 1462
rect 135 1458 139 1462
rect 223 1458 227 1462
rect 303 1458 307 1462
rect 343 1458 347 1462
rect 471 1458 475 1462
rect 607 1458 611 1462
rect 631 1458 635 1462
rect 751 1458 755 1462
rect 783 1458 787 1462
rect 895 1458 899 1462
rect 927 1458 931 1462
rect 1047 1458 1051 1462
rect 1063 1458 1067 1462
rect 1199 1458 1203 1462
rect 1335 1458 1339 1462
rect 1351 1458 1355 1462
rect 1471 1458 1475 1462
rect 1503 1458 1507 1462
rect 1767 1458 1771 1462
rect 1807 1406 1811 1410
rect 1943 1406 1947 1410
rect 2055 1406 2059 1410
rect 2095 1406 2099 1410
rect 2191 1406 2195 1410
rect 2199 1406 2203 1410
rect 2319 1406 2323 1410
rect 2335 1406 2339 1410
rect 2455 1406 2459 1410
rect 2479 1406 2483 1410
rect 2599 1406 2603 1410
rect 2631 1406 2635 1410
rect 2743 1406 2747 1410
rect 2783 1406 2787 1410
rect 2887 1406 2891 1410
rect 2935 1406 2939 1410
rect 3031 1406 3035 1410
rect 3087 1406 3091 1410
rect 3175 1406 3179 1410
rect 3239 1406 3243 1410
rect 3327 1406 3331 1410
rect 3463 1406 3467 1410
rect 111 1390 115 1394
rect 135 1390 139 1394
rect 279 1390 283 1394
rect 303 1390 307 1394
rect 447 1390 451 1394
rect 471 1390 475 1394
rect 607 1390 611 1394
rect 631 1390 635 1394
rect 759 1390 763 1394
rect 783 1390 787 1394
rect 903 1390 907 1394
rect 927 1390 931 1394
rect 1031 1390 1035 1394
rect 1063 1390 1067 1394
rect 1159 1390 1163 1394
rect 1199 1390 1203 1394
rect 1287 1390 1291 1394
rect 1335 1390 1339 1394
rect 1415 1390 1419 1394
rect 1471 1390 1475 1394
rect 1767 1390 1771 1394
rect 1807 1338 1811 1342
rect 2095 1338 2099 1342
rect 2103 1338 2107 1342
rect 2199 1338 2203 1342
rect 2239 1338 2243 1342
rect 2319 1338 2323 1342
rect 2383 1338 2387 1342
rect 2455 1338 2459 1342
rect 2535 1338 2539 1342
rect 2599 1338 2603 1342
rect 2687 1338 2691 1342
rect 2743 1338 2747 1342
rect 2839 1338 2843 1342
rect 2887 1338 2891 1342
rect 2991 1338 2995 1342
rect 3031 1338 3035 1342
rect 3143 1338 3147 1342
rect 3175 1338 3179 1342
rect 3303 1338 3307 1342
rect 3327 1338 3331 1342
rect 3463 1338 3467 1342
rect 111 1322 115 1326
rect 135 1322 139 1326
rect 279 1322 283 1326
rect 439 1322 443 1326
rect 447 1322 451 1326
rect 583 1322 587 1326
rect 607 1322 611 1326
rect 719 1322 723 1326
rect 759 1322 763 1326
rect 847 1322 851 1326
rect 903 1322 907 1326
rect 967 1322 971 1326
rect 1031 1322 1035 1326
rect 1079 1322 1083 1326
rect 1159 1322 1163 1326
rect 1191 1322 1195 1326
rect 1287 1322 1291 1326
rect 1311 1322 1315 1326
rect 1415 1322 1419 1326
rect 1767 1322 1771 1326
rect 1807 1274 1811 1278
rect 1935 1274 1939 1278
rect 2063 1274 2067 1278
rect 2103 1274 2107 1278
rect 2199 1274 2203 1278
rect 2239 1274 2243 1278
rect 2343 1274 2347 1278
rect 2383 1274 2387 1278
rect 2495 1274 2499 1278
rect 2535 1274 2539 1278
rect 2655 1274 2659 1278
rect 2687 1274 2691 1278
rect 2815 1274 2819 1278
rect 2839 1274 2843 1278
rect 2975 1274 2979 1278
rect 2991 1274 2995 1278
rect 3143 1274 3147 1278
rect 3303 1274 3307 1278
rect 3463 1274 3467 1278
rect 111 1254 115 1258
rect 135 1254 139 1258
rect 239 1254 243 1258
rect 279 1254 283 1258
rect 367 1254 371 1258
rect 439 1254 443 1258
rect 495 1254 499 1258
rect 583 1254 587 1258
rect 615 1254 619 1258
rect 719 1254 723 1258
rect 735 1254 739 1258
rect 847 1254 851 1258
rect 959 1254 963 1258
rect 967 1254 971 1258
rect 1071 1254 1075 1258
rect 1079 1254 1083 1258
rect 1191 1254 1195 1258
rect 1311 1254 1315 1258
rect 1767 1254 1771 1258
rect 1807 1210 1811 1214
rect 1831 1210 1835 1214
rect 1935 1210 1939 1214
rect 2063 1210 2067 1214
rect 2079 1210 2083 1214
rect 2199 1210 2203 1214
rect 2231 1210 2235 1214
rect 2343 1210 2347 1214
rect 2391 1210 2395 1214
rect 2495 1210 2499 1214
rect 2543 1210 2547 1214
rect 2655 1210 2659 1214
rect 2695 1210 2699 1214
rect 2815 1210 2819 1214
rect 2847 1210 2851 1214
rect 2975 1210 2979 1214
rect 2999 1210 3003 1214
rect 3143 1210 3147 1214
rect 3159 1210 3163 1214
rect 3463 1210 3467 1214
rect 111 1186 115 1190
rect 135 1186 139 1190
rect 239 1186 243 1190
rect 367 1186 371 1190
rect 375 1186 379 1190
rect 495 1186 499 1190
rect 511 1186 515 1190
rect 615 1186 619 1190
rect 655 1186 659 1190
rect 735 1186 739 1190
rect 791 1186 795 1190
rect 847 1186 851 1190
rect 927 1186 931 1190
rect 959 1186 963 1190
rect 1063 1186 1067 1190
rect 1071 1186 1075 1190
rect 1191 1186 1195 1190
rect 1199 1186 1203 1190
rect 1335 1186 1339 1190
rect 1767 1186 1771 1190
rect 1807 1134 1811 1138
rect 1831 1134 1835 1138
rect 1863 1134 1867 1138
rect 1935 1134 1939 1138
rect 1983 1134 1987 1138
rect 2079 1134 2083 1138
rect 2111 1134 2115 1138
rect 2231 1134 2235 1138
rect 2247 1134 2251 1138
rect 2383 1134 2387 1138
rect 2391 1134 2395 1138
rect 2511 1134 2515 1138
rect 2543 1134 2547 1138
rect 2639 1134 2643 1138
rect 2695 1134 2699 1138
rect 2759 1134 2763 1138
rect 2847 1134 2851 1138
rect 2871 1134 2875 1138
rect 2975 1134 2979 1138
rect 2999 1134 3003 1138
rect 3079 1134 3083 1138
rect 3159 1134 3163 1138
rect 3183 1134 3187 1138
rect 3279 1134 3283 1138
rect 3367 1134 3371 1138
rect 3463 1134 3467 1138
rect 111 1118 115 1122
rect 135 1118 139 1122
rect 191 1118 195 1122
rect 239 1118 243 1122
rect 335 1118 339 1122
rect 375 1118 379 1122
rect 495 1118 499 1122
rect 511 1118 515 1122
rect 655 1118 659 1122
rect 791 1118 795 1122
rect 815 1118 819 1122
rect 927 1118 931 1122
rect 967 1118 971 1122
rect 1063 1118 1067 1122
rect 1119 1118 1123 1122
rect 1199 1118 1203 1122
rect 1263 1118 1267 1122
rect 1335 1118 1339 1122
rect 1407 1118 1411 1122
rect 1559 1118 1563 1122
rect 1767 1118 1771 1122
rect 1807 1062 1811 1066
rect 1863 1062 1867 1066
rect 1983 1062 1987 1066
rect 2103 1062 2107 1066
rect 2111 1062 2115 1066
rect 2191 1062 2195 1066
rect 2247 1062 2251 1066
rect 2279 1062 2283 1066
rect 2367 1062 2371 1066
rect 2383 1062 2387 1066
rect 2455 1062 2459 1066
rect 2511 1062 2515 1066
rect 2543 1062 2547 1066
rect 2631 1062 2635 1066
rect 2639 1062 2643 1066
rect 2719 1062 2723 1066
rect 2759 1062 2763 1066
rect 2807 1062 2811 1066
rect 2871 1062 2875 1066
rect 2975 1062 2979 1066
rect 3079 1062 3083 1066
rect 3183 1062 3187 1066
rect 3279 1062 3283 1066
rect 3367 1062 3371 1066
rect 3463 1062 3467 1066
rect 111 1046 115 1050
rect 191 1046 195 1050
rect 327 1046 331 1050
rect 335 1046 339 1050
rect 463 1046 467 1050
rect 495 1046 499 1050
rect 607 1046 611 1050
rect 655 1046 659 1050
rect 767 1046 771 1050
rect 815 1046 819 1050
rect 927 1046 931 1050
rect 967 1046 971 1050
rect 1079 1046 1083 1050
rect 1119 1046 1123 1050
rect 1231 1046 1235 1050
rect 1263 1046 1267 1050
rect 1383 1046 1387 1050
rect 1407 1046 1411 1050
rect 1535 1046 1539 1050
rect 1559 1046 1563 1050
rect 1671 1046 1675 1050
rect 1767 1046 1771 1050
rect 1807 998 1811 1002
rect 2103 998 2107 1002
rect 2191 998 2195 1002
rect 2279 998 2283 1002
rect 2311 998 2315 1002
rect 2367 998 2371 1002
rect 2407 998 2411 1002
rect 2455 998 2459 1002
rect 2511 998 2515 1002
rect 2543 998 2547 1002
rect 2623 998 2627 1002
rect 2631 998 2635 1002
rect 2719 998 2723 1002
rect 2751 998 2755 1002
rect 2807 998 2811 1002
rect 2895 998 2899 1002
rect 3055 998 3059 1002
rect 3223 998 3227 1002
rect 3367 998 3371 1002
rect 3463 998 3467 1002
rect 111 978 115 982
rect 327 978 331 982
rect 463 978 467 982
rect 471 978 475 982
rect 567 978 571 982
rect 607 978 611 982
rect 671 978 675 982
rect 767 978 771 982
rect 783 978 787 982
rect 887 978 891 982
rect 927 978 931 982
rect 991 978 995 982
rect 1079 978 1083 982
rect 1095 978 1099 982
rect 1199 978 1203 982
rect 1231 978 1235 982
rect 1295 978 1299 982
rect 1383 978 1387 982
rect 1391 978 1395 982
rect 1487 978 1491 982
rect 1535 978 1539 982
rect 1583 978 1587 982
rect 1671 978 1675 982
rect 1767 978 1771 982
rect 1807 922 1811 926
rect 1831 922 1835 926
rect 1983 922 1987 926
rect 2151 922 2155 926
rect 2311 922 2315 926
rect 2327 922 2331 926
rect 2407 922 2411 926
rect 2511 922 2515 926
rect 2519 922 2523 926
rect 2623 922 2627 926
rect 2719 922 2723 926
rect 2751 922 2755 926
rect 2895 922 2899 926
rect 2935 922 2939 926
rect 3055 922 3059 926
rect 3159 922 3163 926
rect 3223 922 3227 926
rect 3367 922 3371 926
rect 3463 922 3467 926
rect 111 910 115 914
rect 471 910 475 914
rect 567 910 571 914
rect 607 910 611 914
rect 671 910 675 914
rect 695 910 699 914
rect 783 910 787 914
rect 791 910 795 914
rect 887 910 891 914
rect 895 910 899 914
rect 991 910 995 914
rect 999 910 1003 914
rect 1095 910 1099 914
rect 1111 910 1115 914
rect 1199 910 1203 914
rect 1223 910 1227 914
rect 1295 910 1299 914
rect 1343 910 1347 914
rect 1391 910 1395 914
rect 1463 910 1467 914
rect 1487 910 1491 914
rect 1583 910 1587 914
rect 1671 910 1675 914
rect 1767 910 1771 914
rect 1807 854 1811 858
rect 1831 854 1835 858
rect 1959 854 1963 858
rect 1983 854 1987 858
rect 2087 854 2091 858
rect 2151 854 2155 858
rect 2207 854 2211 858
rect 2327 854 2331 858
rect 2463 854 2467 858
rect 2519 854 2523 858
rect 2615 854 2619 858
rect 2719 854 2723 858
rect 2791 854 2795 858
rect 2935 854 2939 858
rect 2983 854 2987 858
rect 3159 854 3163 858
rect 3183 854 3187 858
rect 3367 854 3371 858
rect 3463 854 3467 858
rect 111 842 115 846
rect 519 842 523 846
rect 607 842 611 846
rect 615 842 619 846
rect 695 842 699 846
rect 719 842 723 846
rect 791 842 795 846
rect 831 842 835 846
rect 895 842 899 846
rect 951 842 955 846
rect 999 842 1003 846
rect 1071 842 1075 846
rect 1111 842 1115 846
rect 1191 842 1195 846
rect 1223 842 1227 846
rect 1311 842 1315 846
rect 1343 842 1347 846
rect 1431 842 1435 846
rect 1463 842 1467 846
rect 1559 842 1563 846
rect 1583 842 1587 846
rect 1767 842 1771 846
rect 1807 786 1811 790
rect 1831 786 1835 790
rect 1879 786 1883 790
rect 1959 786 1963 790
rect 2015 786 2019 790
rect 2087 786 2091 790
rect 2151 786 2155 790
rect 2207 786 2211 790
rect 2287 786 2291 790
rect 2327 786 2331 790
rect 2423 786 2427 790
rect 2463 786 2467 790
rect 2559 786 2563 790
rect 2615 786 2619 790
rect 2711 786 2715 790
rect 2791 786 2795 790
rect 2871 786 2875 790
rect 2983 786 2987 790
rect 3039 786 3043 790
rect 3183 786 3187 790
rect 3215 786 3219 790
rect 3367 786 3371 790
rect 3463 786 3467 790
rect 111 774 115 778
rect 383 774 387 778
rect 471 774 475 778
rect 519 774 523 778
rect 575 774 579 778
rect 615 774 619 778
rect 679 774 683 778
rect 719 774 723 778
rect 791 774 795 778
rect 831 774 835 778
rect 911 774 915 778
rect 951 774 955 778
rect 1031 774 1035 778
rect 1071 774 1075 778
rect 1159 774 1163 778
rect 1191 774 1195 778
rect 1287 774 1291 778
rect 1311 774 1315 778
rect 1415 774 1419 778
rect 1431 774 1435 778
rect 1559 774 1563 778
rect 1767 774 1771 778
rect 1807 718 1811 722
rect 1831 718 1835 722
rect 1879 718 1883 722
rect 1951 718 1955 722
rect 2015 718 2019 722
rect 2103 718 2107 722
rect 2151 718 2155 722
rect 2263 718 2267 722
rect 2287 718 2291 722
rect 2415 718 2419 722
rect 2423 718 2427 722
rect 2559 718 2563 722
rect 2567 718 2571 722
rect 2711 718 2715 722
rect 2719 718 2723 722
rect 2871 718 2875 722
rect 2879 718 2883 722
rect 3039 718 3043 722
rect 3199 718 3203 722
rect 3215 718 3219 722
rect 3367 718 3371 722
rect 3463 718 3467 722
rect 111 702 115 706
rect 247 702 251 706
rect 343 702 347 706
rect 383 702 387 706
rect 455 702 459 706
rect 471 702 475 706
rect 567 702 571 706
rect 575 702 579 706
rect 679 702 683 706
rect 695 702 699 706
rect 791 702 795 706
rect 831 702 835 706
rect 911 702 915 706
rect 983 702 987 706
rect 1031 702 1035 706
rect 1151 702 1155 706
rect 1159 702 1163 706
rect 1287 702 1291 706
rect 1327 702 1331 706
rect 1415 702 1419 706
rect 1511 702 1515 706
rect 1671 702 1675 706
rect 1767 702 1771 706
rect 1807 654 1811 658
rect 1831 654 1835 658
rect 1951 654 1955 658
rect 1975 654 1979 658
rect 2103 654 2107 658
rect 2239 654 2243 658
rect 2263 654 2267 658
rect 2415 654 2419 658
rect 2479 654 2483 658
rect 2567 654 2571 658
rect 2687 654 2691 658
rect 2719 654 2723 658
rect 2879 654 2883 658
rect 3039 654 3043 658
rect 3055 654 3059 658
rect 3199 654 3203 658
rect 3223 654 3227 658
rect 3367 654 3371 658
rect 3463 654 3467 658
rect 111 634 115 638
rect 135 634 139 638
rect 231 634 235 638
rect 247 634 251 638
rect 343 634 347 638
rect 359 634 363 638
rect 455 634 459 638
rect 487 634 491 638
rect 567 634 571 638
rect 623 634 627 638
rect 695 634 699 638
rect 767 634 771 638
rect 831 634 835 638
rect 911 634 915 638
rect 983 634 987 638
rect 1055 634 1059 638
rect 1151 634 1155 638
rect 1207 634 1211 638
rect 1327 634 1331 638
rect 1367 634 1371 638
rect 1511 634 1515 638
rect 1527 634 1531 638
rect 1671 634 1675 638
rect 1767 634 1771 638
rect 1807 582 1811 586
rect 1895 582 1899 586
rect 1975 582 1979 586
rect 2015 582 2019 586
rect 2143 582 2147 586
rect 2239 582 2243 586
rect 2279 582 2283 586
rect 2423 582 2427 586
rect 2479 582 2483 586
rect 2567 582 2571 586
rect 2687 582 2691 586
rect 2719 582 2723 586
rect 2871 582 2875 586
rect 2879 582 2883 586
rect 3031 582 3035 586
rect 3055 582 3059 586
rect 3199 582 3203 586
rect 3223 582 3227 586
rect 3367 582 3371 586
rect 3463 582 3467 586
rect 111 566 115 570
rect 135 566 139 570
rect 231 566 235 570
rect 247 566 251 570
rect 359 566 363 570
rect 407 566 411 570
rect 487 566 491 570
rect 583 566 587 570
rect 623 566 627 570
rect 767 566 771 570
rect 911 566 915 570
rect 951 566 955 570
rect 1055 566 1059 570
rect 1135 566 1139 570
rect 1207 566 1211 570
rect 1319 566 1323 570
rect 1367 566 1371 570
rect 1503 566 1507 570
rect 1527 566 1531 570
rect 1671 566 1675 570
rect 1767 566 1771 570
rect 1807 514 1811 518
rect 1895 514 1899 518
rect 2015 514 2019 518
rect 2135 514 2139 518
rect 2143 514 2147 518
rect 2239 514 2243 518
rect 2279 514 2283 518
rect 2359 514 2363 518
rect 2423 514 2427 518
rect 2487 514 2491 518
rect 2567 514 2571 518
rect 2615 514 2619 518
rect 2719 514 2723 518
rect 2751 514 2755 518
rect 2871 514 2875 518
rect 2879 514 2883 518
rect 3007 514 3011 518
rect 3031 514 3035 518
rect 3135 514 3139 518
rect 3199 514 3203 518
rect 3263 514 3267 518
rect 3367 514 3371 518
rect 3463 514 3467 518
rect 111 498 115 502
rect 135 498 139 502
rect 247 498 251 502
rect 399 498 403 502
rect 407 498 411 502
rect 567 498 571 502
rect 583 498 587 502
rect 735 498 739 502
rect 767 498 771 502
rect 903 498 907 502
rect 951 498 955 502
rect 1063 498 1067 502
rect 1135 498 1139 502
rect 1223 498 1227 502
rect 1319 498 1323 502
rect 1375 498 1379 502
rect 1503 498 1507 502
rect 1527 498 1531 502
rect 1671 498 1675 502
rect 1767 498 1771 502
rect 1807 442 1811 446
rect 2135 442 2139 446
rect 2239 442 2243 446
rect 2335 442 2339 446
rect 2359 442 2363 446
rect 2447 442 2451 446
rect 2487 442 2491 446
rect 2559 442 2563 446
rect 2615 442 2619 446
rect 2679 442 2683 446
rect 2751 442 2755 446
rect 2799 442 2803 446
rect 2879 442 2883 446
rect 2911 442 2915 446
rect 3007 442 3011 446
rect 3023 442 3027 446
rect 3135 442 3139 446
rect 3143 442 3147 446
rect 3263 442 3267 446
rect 3367 442 3371 446
rect 3463 442 3467 446
rect 111 430 115 434
rect 247 430 251 434
rect 399 430 403 434
rect 519 430 523 434
rect 567 430 571 434
rect 615 430 619 434
rect 719 430 723 434
rect 735 430 739 434
rect 823 430 827 434
rect 903 430 907 434
rect 927 430 931 434
rect 1023 430 1027 434
rect 1063 430 1067 434
rect 1127 430 1131 434
rect 1223 430 1227 434
rect 1231 430 1235 434
rect 1335 430 1339 434
rect 1375 430 1379 434
rect 1439 430 1443 434
rect 1527 430 1531 434
rect 1671 430 1675 434
rect 1767 430 1771 434
rect 1807 374 1811 378
rect 2063 374 2067 378
rect 2151 374 2155 378
rect 2239 374 2243 378
rect 2247 374 2251 378
rect 2335 374 2339 378
rect 2359 374 2363 378
rect 2447 374 2451 378
rect 2479 374 2483 378
rect 2559 374 2563 378
rect 2615 374 2619 378
rect 2679 374 2683 378
rect 2759 374 2763 378
rect 2799 374 2803 378
rect 2911 374 2915 378
rect 3023 374 3027 378
rect 3063 374 3067 378
rect 3143 374 3147 378
rect 3223 374 3227 378
rect 3263 374 3267 378
rect 3367 374 3371 378
rect 3463 374 3467 378
rect 111 362 115 366
rect 471 362 475 366
rect 519 362 523 366
rect 559 362 563 366
rect 615 362 619 366
rect 647 362 651 366
rect 719 362 723 366
rect 735 362 739 366
rect 823 362 827 366
rect 911 362 915 366
rect 927 362 931 366
rect 999 362 1003 366
rect 1023 362 1027 366
rect 1087 362 1091 366
rect 1127 362 1131 366
rect 1175 362 1179 366
rect 1231 362 1235 366
rect 1263 362 1267 366
rect 1335 362 1339 366
rect 1439 362 1443 366
rect 1767 362 1771 366
rect 1807 306 1811 310
rect 1927 306 1931 310
rect 2039 306 2043 310
rect 2063 306 2067 310
rect 2151 306 2155 310
rect 2167 306 2171 310
rect 2247 306 2251 310
rect 2303 306 2307 310
rect 2359 306 2363 310
rect 2447 306 2451 310
rect 2479 306 2483 310
rect 2599 306 2603 310
rect 2615 306 2619 310
rect 2759 306 2763 310
rect 2911 306 2915 310
rect 2919 306 2923 310
rect 3063 306 3067 310
rect 3087 306 3091 310
rect 3223 306 3227 310
rect 3255 306 3259 310
rect 3367 306 3371 310
rect 3463 306 3467 310
rect 111 294 115 298
rect 279 294 283 298
rect 367 294 371 298
rect 463 294 467 298
rect 471 294 475 298
rect 559 294 563 298
rect 647 294 651 298
rect 655 294 659 298
rect 735 294 739 298
rect 751 294 755 298
rect 823 294 827 298
rect 847 294 851 298
rect 911 294 915 298
rect 943 294 947 298
rect 999 294 1003 298
rect 1047 294 1051 298
rect 1087 294 1091 298
rect 1151 294 1155 298
rect 1175 294 1179 298
rect 1263 294 1267 298
rect 1767 294 1771 298
rect 1807 238 1811 242
rect 1831 238 1835 242
rect 1927 238 1931 242
rect 2039 238 2043 242
rect 2055 238 2059 242
rect 2167 238 2171 242
rect 2199 238 2203 242
rect 2303 238 2307 242
rect 2351 238 2355 242
rect 2447 238 2451 242
rect 2511 238 2515 242
rect 2599 238 2603 242
rect 2679 238 2683 242
rect 2759 238 2763 242
rect 2847 238 2851 242
rect 2919 238 2923 242
rect 3023 238 3027 242
rect 3087 238 3091 242
rect 3207 238 3211 242
rect 3255 238 3259 242
rect 3367 238 3371 242
rect 3463 238 3467 242
rect 111 226 115 230
rect 167 226 171 230
rect 279 226 283 230
rect 343 226 347 230
rect 367 226 371 230
rect 463 226 467 230
rect 511 226 515 230
rect 559 226 563 230
rect 655 226 659 230
rect 679 226 683 230
rect 751 226 755 230
rect 839 226 843 230
rect 847 226 851 230
rect 943 226 947 230
rect 991 226 995 230
rect 1047 226 1051 230
rect 1135 226 1139 230
rect 1151 226 1155 230
rect 1279 226 1283 230
rect 1431 226 1435 230
rect 1767 226 1771 230
rect 1807 154 1811 158
rect 1831 154 1835 158
rect 1919 154 1923 158
rect 1927 154 1931 158
rect 2039 154 2043 158
rect 2055 154 2059 158
rect 2159 154 2163 158
rect 2199 154 2203 158
rect 2279 154 2283 158
rect 2351 154 2355 158
rect 2399 154 2403 158
rect 2511 154 2515 158
rect 2623 154 2627 158
rect 2679 154 2683 158
rect 2735 154 2739 158
rect 2839 154 2843 158
rect 2847 154 2851 158
rect 2943 154 2947 158
rect 3023 154 3027 158
rect 3055 154 3059 158
rect 3167 154 3171 158
rect 3207 154 3211 158
rect 3279 154 3283 158
rect 3367 154 3371 158
rect 3463 154 3467 158
rect 111 138 115 142
rect 135 138 139 142
rect 167 138 171 142
rect 223 138 227 142
rect 311 138 315 142
rect 343 138 347 142
rect 399 138 403 142
rect 487 138 491 142
rect 511 138 515 142
rect 575 138 579 142
rect 663 138 667 142
rect 679 138 683 142
rect 751 138 755 142
rect 839 138 843 142
rect 847 138 851 142
rect 943 138 947 142
rect 991 138 995 142
rect 1031 138 1035 142
rect 1119 138 1123 142
rect 1135 138 1139 142
rect 1215 138 1219 142
rect 1279 138 1283 142
rect 1311 138 1315 142
rect 1407 138 1411 142
rect 1431 138 1435 142
rect 1495 138 1499 142
rect 1583 138 1587 142
rect 1671 138 1675 142
rect 1767 138 1771 142
rect 1807 90 1811 94
rect 1831 90 1835 94
rect 1919 90 1923 94
rect 2039 90 2043 94
rect 2159 90 2163 94
rect 2279 90 2283 94
rect 2399 90 2403 94
rect 2511 90 2515 94
rect 2623 90 2627 94
rect 2735 90 2739 94
rect 2839 90 2843 94
rect 2943 90 2947 94
rect 3055 90 3059 94
rect 3167 90 3171 94
rect 3279 90 3283 94
rect 3367 90 3371 94
rect 3463 90 3467 94
rect 111 74 115 78
rect 135 74 139 78
rect 223 74 227 78
rect 311 74 315 78
rect 399 74 403 78
rect 487 74 491 78
rect 575 74 579 78
rect 663 74 667 78
rect 751 74 755 78
rect 847 74 851 78
rect 943 74 947 78
rect 1031 74 1035 78
rect 1119 74 1123 78
rect 1215 74 1219 78
rect 1311 74 1315 78
rect 1407 74 1411 78
rect 1495 74 1499 78
rect 1583 74 1587 78
rect 1671 74 1675 78
rect 1767 74 1771 78
<< m4 >>
rect 1790 3517 1791 3523
rect 1797 3522 3499 3523
rect 1797 3518 1807 3522
rect 1811 3518 2007 3522
rect 2011 3518 2239 3522
rect 2243 3518 2455 3522
rect 2459 3518 2655 3522
rect 2659 3518 2855 3522
rect 2859 3518 3047 3522
rect 3051 3518 3247 3522
rect 3251 3518 3463 3522
rect 3467 3518 3499 3522
rect 1797 3517 3499 3518
rect 3505 3517 3506 3523
rect 96 3481 97 3487
rect 103 3486 1791 3487
rect 103 3482 111 3486
rect 115 3482 455 3486
rect 459 3482 543 3486
rect 547 3482 631 3486
rect 635 3482 719 3486
rect 723 3482 807 3486
rect 811 3482 895 3486
rect 899 3482 983 3486
rect 987 3482 1071 3486
rect 1075 3482 1159 3486
rect 1163 3482 1767 3486
rect 1771 3482 1791 3486
rect 103 3481 1791 3482
rect 1797 3481 1798 3487
rect 1778 3453 1779 3459
rect 1785 3458 3487 3459
rect 1785 3454 1807 3458
rect 1811 3454 1831 3458
rect 1835 3454 1943 3458
rect 1947 3454 2007 3458
rect 2011 3454 2079 3458
rect 2083 3454 2215 3458
rect 2219 3454 2239 3458
rect 2243 3454 2351 3458
rect 2355 3454 2455 3458
rect 2459 3454 2479 3458
rect 2483 3454 2599 3458
rect 2603 3454 2655 3458
rect 2659 3454 2719 3458
rect 2723 3454 2847 3458
rect 2851 3454 2855 3458
rect 2859 3454 2975 3458
rect 2979 3454 3047 3458
rect 3051 3454 3247 3458
rect 3251 3454 3463 3458
rect 3467 3454 3487 3458
rect 1785 3453 3487 3454
rect 3493 3453 3494 3459
rect 84 3417 85 3423
rect 91 3422 1779 3423
rect 91 3418 111 3422
rect 115 3418 415 3422
rect 419 3418 455 3422
rect 459 3418 503 3422
rect 507 3418 543 3422
rect 547 3418 591 3422
rect 595 3418 631 3422
rect 635 3418 679 3422
rect 683 3418 719 3422
rect 723 3418 767 3422
rect 771 3418 807 3422
rect 811 3418 855 3422
rect 859 3418 895 3422
rect 899 3418 943 3422
rect 947 3418 983 3422
rect 987 3418 1031 3422
rect 1035 3418 1071 3422
rect 1075 3418 1119 3422
rect 1123 3418 1159 3422
rect 1163 3418 1207 3422
rect 1211 3418 1303 3422
rect 1307 3418 1767 3422
rect 1771 3418 1779 3422
rect 91 3417 1779 3418
rect 1785 3417 1786 3423
rect 1790 3381 1791 3387
rect 1797 3386 3499 3387
rect 1797 3382 1807 3386
rect 1811 3382 1831 3386
rect 1835 3382 1943 3386
rect 1947 3382 1951 3386
rect 1955 3382 2079 3386
rect 2083 3382 2095 3386
rect 2099 3382 2215 3386
rect 2219 3382 2239 3386
rect 2243 3382 2351 3386
rect 2355 3382 2383 3386
rect 2387 3382 2479 3386
rect 2483 3382 2519 3386
rect 2523 3382 2599 3386
rect 2603 3382 2647 3386
rect 2651 3382 2719 3386
rect 2723 3382 2775 3386
rect 2779 3382 2847 3386
rect 2851 3382 2903 3386
rect 2907 3382 2975 3386
rect 2979 3382 3039 3386
rect 3043 3382 3463 3386
rect 3467 3382 3499 3386
rect 1797 3381 3499 3382
rect 3505 3381 3506 3387
rect 96 3349 97 3355
rect 103 3354 1791 3355
rect 103 3350 111 3354
rect 115 3350 399 3354
rect 403 3350 415 3354
rect 419 3350 495 3354
rect 499 3350 503 3354
rect 507 3350 591 3354
rect 595 3350 599 3354
rect 603 3350 679 3354
rect 683 3350 703 3354
rect 707 3350 767 3354
rect 771 3350 807 3354
rect 811 3350 855 3354
rect 859 3350 911 3354
rect 915 3350 943 3354
rect 947 3350 1015 3354
rect 1019 3350 1031 3354
rect 1035 3350 1119 3354
rect 1123 3350 1207 3354
rect 1211 3350 1223 3354
rect 1227 3350 1303 3354
rect 1307 3350 1327 3354
rect 1331 3350 1767 3354
rect 1771 3350 1791 3354
rect 103 3349 1791 3350
rect 1797 3349 1798 3355
rect 1778 3309 1779 3315
rect 1785 3314 3487 3315
rect 1785 3310 1807 3314
rect 1811 3310 1831 3314
rect 1835 3310 1951 3314
rect 1955 3310 1975 3314
rect 1979 3310 2095 3314
rect 2099 3310 2151 3314
rect 2155 3310 2239 3314
rect 2243 3310 2335 3314
rect 2339 3310 2383 3314
rect 2387 3310 2511 3314
rect 2515 3310 2519 3314
rect 2523 3310 2647 3314
rect 2651 3310 2679 3314
rect 2683 3310 2775 3314
rect 2779 3310 2831 3314
rect 2835 3310 2903 3314
rect 2907 3310 2975 3314
rect 2979 3310 3039 3314
rect 3043 3310 3111 3314
rect 3115 3310 3247 3314
rect 3251 3310 3367 3314
rect 3371 3310 3463 3314
rect 3467 3310 3487 3314
rect 1785 3309 3487 3310
rect 3493 3309 3494 3315
rect 84 3281 85 3287
rect 91 3286 1779 3287
rect 91 3282 111 3286
rect 115 3282 383 3286
rect 387 3282 399 3286
rect 403 3282 495 3286
rect 499 3282 599 3286
rect 603 3282 607 3286
rect 611 3282 703 3286
rect 707 3282 727 3286
rect 731 3282 807 3286
rect 811 3282 847 3286
rect 851 3282 911 3286
rect 915 3282 967 3286
rect 971 3282 1015 3286
rect 1019 3282 1087 3286
rect 1091 3282 1119 3286
rect 1123 3282 1207 3286
rect 1211 3282 1223 3286
rect 1227 3282 1327 3286
rect 1331 3282 1335 3286
rect 1339 3282 1767 3286
rect 1771 3282 1779 3286
rect 91 3281 1779 3282
rect 1785 3281 1786 3287
rect 1790 3237 1791 3243
rect 1797 3242 3499 3243
rect 1797 3238 1807 3242
rect 1811 3238 1831 3242
rect 1835 3238 1975 3242
rect 1979 3238 2031 3242
rect 2035 3238 2151 3242
rect 2155 3238 2247 3242
rect 2251 3238 2335 3242
rect 2339 3238 2455 3242
rect 2459 3238 2511 3242
rect 2515 3238 2655 3242
rect 2659 3238 2679 3242
rect 2683 3238 2831 3242
rect 2835 3238 2839 3242
rect 2843 3238 2975 3242
rect 2979 3238 3023 3242
rect 3027 3238 3111 3242
rect 3115 3238 3207 3242
rect 3211 3238 3247 3242
rect 3251 3238 3367 3242
rect 3371 3238 3463 3242
rect 3467 3238 3499 3242
rect 1797 3237 3499 3238
rect 3505 3237 3506 3243
rect 96 3213 97 3219
rect 103 3218 1791 3219
rect 103 3214 111 3218
rect 115 3214 303 3218
rect 307 3214 383 3218
rect 387 3214 423 3218
rect 427 3214 495 3218
rect 499 3214 543 3218
rect 547 3214 607 3218
rect 611 3214 671 3218
rect 675 3214 727 3218
rect 731 3214 799 3218
rect 803 3214 847 3218
rect 851 3214 927 3218
rect 931 3214 967 3218
rect 971 3214 1055 3218
rect 1059 3214 1087 3218
rect 1091 3214 1175 3218
rect 1179 3214 1207 3218
rect 1211 3214 1303 3218
rect 1307 3214 1335 3218
rect 1339 3214 1431 3218
rect 1435 3214 1767 3218
rect 1771 3214 1791 3218
rect 103 3213 1791 3214
rect 1797 3213 1798 3219
rect 1778 3173 1779 3179
rect 1785 3178 3487 3179
rect 1785 3174 1807 3178
rect 1811 3174 1831 3178
rect 1835 3174 1839 3178
rect 1843 3174 2031 3178
rect 2035 3174 2223 3178
rect 2227 3174 2247 3178
rect 2251 3174 2407 3178
rect 2411 3174 2455 3178
rect 2459 3174 2575 3178
rect 2579 3174 2655 3178
rect 2659 3174 2735 3178
rect 2739 3174 2839 3178
rect 2843 3174 2879 3178
rect 2883 3174 3007 3178
rect 3011 3174 3023 3178
rect 3027 3174 3135 3178
rect 3139 3174 3207 3178
rect 3211 3174 3263 3178
rect 3267 3174 3367 3178
rect 3371 3174 3463 3178
rect 3467 3174 3487 3178
rect 1785 3173 3487 3174
rect 3493 3173 3494 3179
rect 84 3137 85 3143
rect 91 3142 1779 3143
rect 91 3138 111 3142
rect 115 3138 175 3142
rect 179 3138 303 3142
rect 307 3138 319 3142
rect 323 3138 423 3142
rect 427 3138 471 3142
rect 475 3138 543 3142
rect 547 3138 623 3142
rect 627 3138 671 3142
rect 675 3138 775 3142
rect 779 3138 799 3142
rect 803 3138 919 3142
rect 923 3138 927 3142
rect 931 3138 1055 3142
rect 1059 3138 1063 3142
rect 1067 3138 1175 3142
rect 1179 3138 1199 3142
rect 1203 3138 1303 3142
rect 1307 3138 1343 3142
rect 1347 3138 1431 3142
rect 1435 3138 1487 3142
rect 1491 3138 1767 3142
rect 1771 3138 1779 3142
rect 91 3137 1779 3138
rect 1785 3137 1786 3143
rect 1790 3105 1791 3111
rect 1797 3110 3499 3111
rect 1797 3106 1807 3110
rect 1811 3106 1839 3110
rect 1843 3106 1935 3110
rect 1939 3106 2031 3110
rect 2035 3106 2055 3110
rect 2059 3106 2175 3110
rect 2179 3106 2223 3110
rect 2227 3106 2303 3110
rect 2307 3106 2407 3110
rect 2411 3106 2431 3110
rect 2435 3106 2567 3110
rect 2571 3106 2575 3110
rect 2579 3106 2719 3110
rect 2723 3106 2735 3110
rect 2739 3106 2871 3110
rect 2875 3106 2879 3110
rect 2883 3106 3007 3110
rect 3011 3106 3031 3110
rect 3035 3106 3135 3110
rect 3139 3106 3199 3110
rect 3203 3106 3263 3110
rect 3267 3106 3367 3110
rect 3371 3106 3463 3110
rect 3467 3106 3499 3110
rect 1797 3105 3499 3106
rect 3505 3105 3506 3111
rect 96 3065 97 3071
rect 103 3070 1791 3071
rect 103 3066 111 3070
rect 115 3066 135 3070
rect 139 3066 175 3070
rect 179 3066 263 3070
rect 267 3066 319 3070
rect 323 3066 431 3070
rect 435 3066 471 3070
rect 475 3066 607 3070
rect 611 3066 623 3070
rect 627 3066 775 3070
rect 779 3066 791 3070
rect 795 3066 919 3070
rect 923 3066 967 3070
rect 971 3066 1063 3070
rect 1067 3066 1143 3070
rect 1147 3066 1199 3070
rect 1203 3066 1327 3070
rect 1331 3066 1343 3070
rect 1347 3066 1487 3070
rect 1491 3066 1511 3070
rect 1515 3066 1767 3070
rect 1771 3066 1791 3070
rect 103 3065 1791 3066
rect 1797 3065 1798 3071
rect 1778 3033 1779 3039
rect 1785 3038 3487 3039
rect 1785 3034 1807 3038
rect 1811 3034 1935 3038
rect 1939 3034 2023 3038
rect 2027 3034 2055 3038
rect 2059 3034 2127 3038
rect 2131 3034 2175 3038
rect 2179 3034 2231 3038
rect 2235 3034 2303 3038
rect 2307 3034 2335 3038
rect 2339 3034 2431 3038
rect 2435 3034 2439 3038
rect 2443 3034 2543 3038
rect 2547 3034 2567 3038
rect 2571 3034 2647 3038
rect 2651 3034 2719 3038
rect 2723 3034 2759 3038
rect 2763 3034 2871 3038
rect 2875 3034 3031 3038
rect 3035 3034 3199 3038
rect 3203 3034 3367 3038
rect 3371 3034 3463 3038
rect 3467 3034 3487 3038
rect 1785 3033 3487 3034
rect 3493 3033 3494 3039
rect 84 2997 85 3003
rect 91 3002 1779 3003
rect 91 2998 111 3002
rect 115 2998 135 3002
rect 139 2998 263 3002
rect 267 2998 327 3002
rect 331 2998 431 3002
rect 435 2998 535 3002
rect 539 2998 607 3002
rect 611 2998 735 3002
rect 739 2998 791 3002
rect 795 2998 927 3002
rect 931 2998 967 3002
rect 971 2998 1103 3002
rect 1107 2998 1143 3002
rect 1147 2998 1279 3002
rect 1283 2998 1327 3002
rect 1331 2998 1447 3002
rect 1451 2998 1511 3002
rect 1515 2998 1623 3002
rect 1627 2998 1767 3002
rect 1771 2998 1779 3002
rect 91 2997 1779 2998
rect 1785 2997 1786 3003
rect 1790 2969 1791 2975
rect 1797 2974 3499 2975
rect 1797 2970 1807 2974
rect 1811 2970 2023 2974
rect 2027 2970 2055 2974
rect 2059 2970 2127 2974
rect 2131 2970 2143 2974
rect 2147 2970 2231 2974
rect 2235 2970 2319 2974
rect 2323 2970 2335 2974
rect 2339 2970 2407 2974
rect 2411 2970 2439 2974
rect 2443 2970 2495 2974
rect 2499 2970 2543 2974
rect 2547 2970 2583 2974
rect 2587 2970 2647 2974
rect 2651 2970 2671 2974
rect 2675 2970 2759 2974
rect 2763 2970 2847 2974
rect 2851 2970 3463 2974
rect 3467 2970 3499 2974
rect 1797 2969 3499 2970
rect 3505 2969 3506 2975
rect 96 2925 97 2931
rect 103 2930 1791 2931
rect 103 2926 111 2930
rect 115 2926 135 2930
rect 139 2926 263 2930
rect 267 2926 327 2930
rect 331 2926 431 2930
rect 435 2926 535 2930
rect 539 2926 607 2930
rect 611 2926 735 2930
rect 739 2926 783 2930
rect 787 2926 927 2930
rect 931 2926 951 2930
rect 955 2926 1103 2930
rect 1107 2926 1111 2930
rect 1115 2926 1271 2930
rect 1275 2926 1279 2930
rect 1283 2926 1431 2930
rect 1435 2926 1447 2930
rect 1451 2926 1591 2930
rect 1595 2926 1623 2930
rect 1627 2926 1767 2930
rect 1771 2926 1791 2930
rect 103 2925 1791 2926
rect 1797 2925 1798 2931
rect 1778 2897 1779 2903
rect 1785 2902 3487 2903
rect 1785 2898 1807 2902
rect 1811 2898 2055 2902
rect 2059 2898 2071 2902
rect 2075 2898 2143 2902
rect 2147 2898 2175 2902
rect 2179 2898 2231 2902
rect 2235 2898 2271 2902
rect 2275 2898 2319 2902
rect 2323 2898 2367 2902
rect 2371 2898 2407 2902
rect 2411 2898 2471 2902
rect 2475 2898 2495 2902
rect 2499 2898 2575 2902
rect 2579 2898 2583 2902
rect 2587 2898 2671 2902
rect 2675 2898 2679 2902
rect 2683 2898 2759 2902
rect 2763 2898 2783 2902
rect 2787 2898 2847 2902
rect 2851 2898 3463 2902
rect 3467 2898 3487 2902
rect 1785 2897 3487 2898
rect 3493 2897 3494 2903
rect 84 2857 85 2863
rect 91 2862 1779 2863
rect 91 2858 111 2862
rect 115 2858 135 2862
rect 139 2858 255 2862
rect 259 2858 263 2862
rect 267 2858 407 2862
rect 411 2858 431 2862
rect 435 2858 567 2862
rect 571 2858 607 2862
rect 611 2858 727 2862
rect 731 2858 783 2862
rect 787 2858 879 2862
rect 883 2858 951 2862
rect 955 2858 1023 2862
rect 1027 2858 1111 2862
rect 1115 2858 1167 2862
rect 1171 2858 1271 2862
rect 1275 2858 1311 2862
rect 1315 2858 1431 2862
rect 1435 2858 1463 2862
rect 1467 2858 1591 2862
rect 1595 2858 1767 2862
rect 1771 2858 1779 2862
rect 91 2857 1779 2858
rect 1785 2857 1786 2863
rect 1790 2829 1791 2835
rect 1797 2834 3499 2835
rect 1797 2830 1807 2834
rect 1811 2830 1983 2834
rect 1987 2830 2071 2834
rect 2075 2830 2111 2834
rect 2115 2830 2175 2834
rect 2179 2830 2239 2834
rect 2243 2830 2271 2834
rect 2275 2830 2367 2834
rect 2371 2830 2471 2834
rect 2475 2830 2487 2834
rect 2491 2830 2575 2834
rect 2579 2830 2607 2834
rect 2611 2830 2679 2834
rect 2683 2830 2719 2834
rect 2723 2830 2783 2834
rect 2787 2830 2839 2834
rect 2843 2830 2959 2834
rect 2963 2830 3463 2834
rect 3467 2830 3499 2834
rect 1797 2829 3499 2830
rect 3505 2829 3506 2835
rect 96 2785 97 2791
rect 103 2790 1791 2791
rect 103 2786 111 2790
rect 115 2786 135 2790
rect 139 2786 255 2790
rect 259 2786 287 2790
rect 291 2786 391 2790
rect 395 2786 407 2790
rect 411 2786 503 2790
rect 507 2786 567 2790
rect 571 2786 623 2790
rect 627 2786 727 2790
rect 731 2786 743 2790
rect 747 2786 855 2790
rect 859 2786 879 2790
rect 883 2786 967 2790
rect 971 2786 1023 2790
rect 1027 2786 1079 2790
rect 1083 2786 1167 2790
rect 1171 2786 1199 2790
rect 1203 2786 1311 2790
rect 1315 2786 1319 2790
rect 1323 2786 1463 2790
rect 1467 2786 1767 2790
rect 1771 2786 1791 2790
rect 103 2785 1791 2786
rect 1797 2785 1798 2791
rect 1778 2761 1779 2767
rect 1785 2766 3487 2767
rect 1785 2762 1807 2766
rect 1811 2762 1887 2766
rect 1891 2762 1983 2766
rect 1987 2762 2031 2766
rect 2035 2762 2111 2766
rect 2115 2762 2183 2766
rect 2187 2762 2239 2766
rect 2243 2762 2335 2766
rect 2339 2762 2367 2766
rect 2371 2762 2479 2766
rect 2483 2762 2487 2766
rect 2491 2762 2607 2766
rect 2611 2762 2623 2766
rect 2627 2762 2719 2766
rect 2723 2762 2767 2766
rect 2771 2762 2839 2766
rect 2843 2762 2911 2766
rect 2915 2762 2959 2766
rect 2963 2762 3055 2766
rect 3059 2762 3463 2766
rect 3467 2762 3487 2766
rect 1785 2761 3487 2762
rect 3493 2761 3494 2767
rect 84 2717 85 2723
rect 91 2722 1779 2723
rect 91 2718 111 2722
rect 115 2718 287 2722
rect 291 2718 391 2722
rect 395 2718 479 2722
rect 483 2718 503 2722
rect 507 2718 567 2722
rect 571 2718 623 2722
rect 627 2718 655 2722
rect 659 2718 743 2722
rect 747 2718 831 2722
rect 835 2718 855 2722
rect 859 2718 919 2722
rect 923 2718 967 2722
rect 971 2718 1007 2722
rect 1011 2718 1079 2722
rect 1083 2718 1095 2722
rect 1099 2718 1183 2722
rect 1187 2718 1199 2722
rect 1203 2718 1319 2722
rect 1323 2718 1767 2722
rect 1771 2718 1779 2722
rect 91 2717 1779 2718
rect 1785 2717 1786 2723
rect 1790 2697 1791 2703
rect 1797 2702 3499 2703
rect 1797 2698 1807 2702
rect 1811 2698 1831 2702
rect 1835 2698 1887 2702
rect 1891 2698 2023 2702
rect 2027 2698 2031 2702
rect 2035 2698 2183 2702
rect 2187 2698 2231 2702
rect 2235 2698 2335 2702
rect 2339 2698 2431 2702
rect 2435 2698 2479 2702
rect 2483 2698 2615 2702
rect 2619 2698 2623 2702
rect 2627 2698 2767 2702
rect 2771 2698 2783 2702
rect 2787 2698 2911 2702
rect 2915 2698 2943 2702
rect 2947 2698 3055 2702
rect 3059 2698 3095 2702
rect 3099 2698 3239 2702
rect 3243 2698 3367 2702
rect 3371 2698 3463 2702
rect 3467 2698 3499 2702
rect 1797 2697 3499 2698
rect 3505 2697 3506 2703
rect 96 2645 97 2651
rect 103 2650 1791 2651
rect 103 2646 111 2650
rect 115 2646 471 2650
rect 475 2646 479 2650
rect 483 2646 559 2650
rect 563 2646 567 2650
rect 571 2646 647 2650
rect 651 2646 655 2650
rect 659 2646 735 2650
rect 739 2646 743 2650
rect 747 2646 823 2650
rect 827 2646 831 2650
rect 835 2646 911 2650
rect 915 2646 919 2650
rect 923 2646 999 2650
rect 1003 2646 1007 2650
rect 1011 2646 1087 2650
rect 1091 2646 1095 2650
rect 1099 2646 1183 2650
rect 1187 2646 1767 2650
rect 1771 2646 1791 2650
rect 103 2645 1791 2646
rect 1797 2645 1798 2651
rect 1778 2629 1779 2635
rect 1785 2634 3487 2635
rect 1785 2630 1807 2634
rect 1811 2630 1831 2634
rect 1835 2630 1999 2634
rect 2003 2630 2023 2634
rect 2027 2630 2183 2634
rect 2187 2630 2231 2634
rect 2235 2630 2359 2634
rect 2363 2630 2431 2634
rect 2435 2630 2519 2634
rect 2523 2630 2615 2634
rect 2619 2630 2671 2634
rect 2675 2630 2783 2634
rect 2787 2630 2807 2634
rect 2811 2630 2927 2634
rect 2931 2630 2943 2634
rect 2947 2630 3047 2634
rect 3051 2630 3095 2634
rect 3099 2630 3159 2634
rect 3163 2630 3239 2634
rect 3243 2630 3271 2634
rect 3275 2630 3367 2634
rect 3371 2630 3463 2634
rect 3467 2630 3487 2634
rect 1785 2629 3487 2630
rect 3493 2629 3494 2635
rect 84 2569 85 2575
rect 91 2574 1779 2575
rect 91 2570 111 2574
rect 115 2570 223 2574
rect 227 2570 311 2574
rect 315 2570 407 2574
rect 411 2570 471 2574
rect 475 2570 503 2574
rect 507 2570 559 2574
rect 563 2570 591 2574
rect 595 2570 647 2574
rect 651 2570 679 2574
rect 683 2570 735 2574
rect 739 2570 767 2574
rect 771 2570 823 2574
rect 827 2570 855 2574
rect 859 2570 911 2574
rect 915 2570 943 2574
rect 947 2570 999 2574
rect 1003 2570 1031 2574
rect 1035 2570 1087 2574
rect 1091 2570 1119 2574
rect 1123 2570 1215 2574
rect 1219 2570 1311 2574
rect 1315 2570 1407 2574
rect 1411 2570 1495 2574
rect 1499 2570 1583 2574
rect 1587 2570 1671 2574
rect 1675 2570 1767 2574
rect 1771 2570 1779 2574
rect 91 2569 1779 2570
rect 1785 2569 1786 2575
rect 1790 2557 1791 2563
rect 1797 2562 3499 2563
rect 1797 2558 1807 2562
rect 1811 2558 1831 2562
rect 1835 2558 1999 2562
rect 2003 2558 2183 2562
rect 2187 2558 2207 2562
rect 2211 2558 2359 2562
rect 2363 2558 2519 2562
rect 2523 2558 2671 2562
rect 2675 2558 2799 2562
rect 2803 2558 2807 2562
rect 2811 2558 2927 2562
rect 2931 2558 3047 2562
rect 3051 2558 3159 2562
rect 3163 2558 3271 2562
rect 3275 2558 3367 2562
rect 3371 2558 3463 2562
rect 3467 2558 3499 2562
rect 1797 2557 3499 2558
rect 3505 2557 3506 2563
rect 96 2505 97 2511
rect 103 2510 1791 2511
rect 103 2506 111 2510
rect 115 2506 135 2510
rect 139 2506 223 2510
rect 227 2506 247 2510
rect 251 2506 311 2510
rect 315 2506 391 2510
rect 395 2506 407 2510
rect 411 2506 503 2510
rect 507 2506 543 2510
rect 547 2506 591 2510
rect 595 2506 679 2510
rect 683 2506 695 2510
rect 699 2506 767 2510
rect 771 2506 839 2510
rect 843 2506 855 2510
rect 859 2506 943 2510
rect 947 2506 975 2510
rect 979 2506 1031 2510
rect 1035 2506 1103 2510
rect 1107 2506 1119 2510
rect 1123 2506 1215 2510
rect 1219 2506 1231 2510
rect 1235 2506 1311 2510
rect 1315 2506 1351 2510
rect 1355 2506 1407 2510
rect 1411 2506 1463 2510
rect 1467 2506 1495 2510
rect 1499 2506 1575 2510
rect 1579 2506 1583 2510
rect 1587 2506 1671 2510
rect 1675 2506 1767 2510
rect 1771 2506 1791 2510
rect 103 2505 1791 2506
rect 1797 2505 1798 2511
rect 1778 2477 1779 2483
rect 1785 2482 3487 2483
rect 1785 2478 1807 2482
rect 1811 2478 2015 2482
rect 2019 2478 2199 2482
rect 2203 2478 2207 2482
rect 2211 2478 2367 2482
rect 2371 2478 2527 2482
rect 2531 2478 2671 2482
rect 2675 2478 2799 2482
rect 2803 2478 2807 2482
rect 2811 2478 2927 2482
rect 2931 2478 3047 2482
rect 3051 2478 3159 2482
rect 3163 2478 3271 2482
rect 3275 2478 3367 2482
rect 3371 2478 3463 2482
rect 3467 2478 3487 2482
rect 1785 2477 3487 2478
rect 3493 2477 3494 2483
rect 84 2425 85 2431
rect 91 2430 1779 2431
rect 91 2426 111 2430
rect 115 2426 135 2430
rect 139 2426 239 2430
rect 243 2426 247 2430
rect 251 2426 391 2430
rect 395 2426 543 2430
rect 547 2426 551 2430
rect 555 2426 695 2430
rect 699 2426 719 2430
rect 723 2426 839 2430
rect 843 2426 895 2430
rect 899 2426 975 2430
rect 979 2426 1063 2430
rect 1067 2426 1103 2430
rect 1107 2426 1231 2430
rect 1235 2426 1239 2430
rect 1243 2426 1351 2430
rect 1355 2426 1415 2430
rect 1419 2426 1463 2430
rect 1467 2426 1575 2430
rect 1579 2426 1591 2430
rect 1595 2426 1671 2430
rect 1675 2426 1767 2430
rect 1771 2426 1779 2430
rect 91 2425 1779 2426
rect 1785 2425 1786 2431
rect 1790 2409 1791 2415
rect 1797 2414 3499 2415
rect 1797 2410 1807 2414
rect 1811 2410 1839 2414
rect 1843 2410 2007 2414
rect 2011 2410 2015 2414
rect 2019 2410 2183 2414
rect 2187 2410 2199 2414
rect 2203 2410 2367 2414
rect 2371 2410 2527 2414
rect 2531 2410 2559 2414
rect 2563 2410 2671 2414
rect 2675 2410 2759 2414
rect 2763 2410 2807 2414
rect 2811 2410 2927 2414
rect 2931 2410 2967 2414
rect 2971 2410 3047 2414
rect 3051 2410 3159 2414
rect 3163 2410 3175 2414
rect 3179 2410 3271 2414
rect 3275 2410 3367 2414
rect 3371 2410 3463 2414
rect 3467 2410 3499 2414
rect 1797 2409 3499 2410
rect 3505 2409 3506 2415
rect 1778 2363 1779 2369
rect 1785 2363 1810 2369
rect 96 2353 97 2359
rect 103 2358 1791 2359
rect 103 2354 111 2358
rect 115 2354 135 2358
rect 139 2354 239 2358
rect 243 2354 375 2358
rect 379 2354 391 2358
rect 395 2354 479 2358
rect 483 2354 551 2358
rect 555 2354 599 2358
rect 603 2354 719 2358
rect 723 2354 847 2358
rect 851 2354 895 2358
rect 899 2354 975 2358
rect 979 2354 1063 2358
rect 1067 2354 1103 2358
rect 1107 2354 1239 2358
rect 1243 2354 1375 2358
rect 1379 2354 1415 2358
rect 1419 2354 1511 2358
rect 1515 2354 1591 2358
rect 1595 2354 1767 2358
rect 1771 2354 1791 2358
rect 103 2353 1791 2354
rect 1797 2353 1798 2359
rect 1804 2351 1810 2363
rect 1804 2350 3487 2351
rect 1804 2346 1807 2350
rect 1811 2346 1839 2350
rect 1843 2346 1887 2350
rect 1891 2346 2007 2350
rect 2011 2346 2015 2350
rect 2019 2346 2151 2350
rect 2155 2346 2183 2350
rect 2187 2346 2303 2350
rect 2307 2346 2367 2350
rect 2371 2346 2463 2350
rect 2467 2346 2559 2350
rect 2563 2346 2647 2350
rect 2651 2346 2759 2350
rect 2763 2346 2839 2350
rect 2843 2346 2967 2350
rect 2971 2346 3047 2350
rect 3051 2346 3175 2350
rect 3179 2346 3255 2350
rect 3259 2346 3367 2350
rect 3371 2346 3463 2350
rect 3467 2346 3487 2350
rect 1804 2345 3487 2346
rect 3493 2345 3494 2351
rect 84 2281 85 2287
rect 91 2286 1779 2287
rect 91 2282 111 2286
rect 115 2282 375 2286
rect 379 2282 479 2286
rect 483 2282 575 2286
rect 579 2282 599 2286
rect 603 2282 663 2286
rect 667 2282 719 2286
rect 723 2282 759 2286
rect 763 2282 847 2286
rect 851 2282 863 2286
rect 867 2282 967 2286
rect 971 2282 975 2286
rect 979 2282 1079 2286
rect 1083 2282 1103 2286
rect 1107 2282 1191 2286
rect 1195 2282 1239 2286
rect 1243 2282 1303 2286
rect 1307 2282 1375 2286
rect 1379 2282 1415 2286
rect 1419 2282 1511 2286
rect 1515 2282 1767 2286
rect 1771 2282 1779 2286
rect 91 2281 1779 2282
rect 1785 2281 1786 2287
rect 1790 2277 1791 2283
rect 1797 2282 3499 2283
rect 1797 2278 1807 2282
rect 1811 2278 1887 2282
rect 1891 2278 2015 2282
rect 2019 2278 2039 2282
rect 2043 2278 2135 2282
rect 2139 2278 2151 2282
rect 2155 2278 2239 2282
rect 2243 2278 2303 2282
rect 2307 2278 2343 2282
rect 2347 2278 2463 2282
rect 2467 2278 2591 2282
rect 2595 2278 2647 2282
rect 2651 2278 2735 2282
rect 2739 2278 2839 2282
rect 2843 2278 2887 2282
rect 2891 2278 3047 2282
rect 3051 2278 3215 2282
rect 3219 2278 3255 2282
rect 3259 2278 3367 2282
rect 3371 2278 3463 2282
rect 3467 2278 3499 2282
rect 1797 2277 3499 2278
rect 3505 2277 3506 2283
rect 96 2217 97 2223
rect 103 2222 1791 2223
rect 103 2218 111 2222
rect 115 2218 439 2222
rect 443 2218 527 2222
rect 531 2218 575 2222
rect 579 2218 615 2222
rect 619 2218 663 2222
rect 667 2218 703 2222
rect 707 2218 759 2222
rect 763 2218 791 2222
rect 795 2218 863 2222
rect 867 2218 879 2222
rect 883 2218 967 2222
rect 971 2218 1055 2222
rect 1059 2218 1079 2222
rect 1083 2218 1143 2222
rect 1147 2218 1191 2222
rect 1195 2218 1231 2222
rect 1235 2218 1303 2222
rect 1307 2218 1319 2222
rect 1323 2218 1415 2222
rect 1419 2218 1767 2222
rect 1771 2218 1791 2222
rect 103 2217 1791 2218
rect 1797 2217 1798 2223
rect 1778 2201 1779 2207
rect 1785 2206 3487 2207
rect 1785 2202 1807 2206
rect 1811 2202 2039 2206
rect 2043 2202 2135 2206
rect 2139 2202 2183 2206
rect 2187 2202 2239 2206
rect 2243 2202 2279 2206
rect 2283 2202 2343 2206
rect 2347 2202 2383 2206
rect 2387 2202 2463 2206
rect 2467 2202 2495 2206
rect 2499 2202 2591 2206
rect 2595 2202 2607 2206
rect 2611 2202 2719 2206
rect 2723 2202 2735 2206
rect 2739 2202 2839 2206
rect 2843 2202 2887 2206
rect 2891 2202 2967 2206
rect 2971 2202 3047 2206
rect 3051 2202 3103 2206
rect 3107 2202 3215 2206
rect 3219 2202 3247 2206
rect 3251 2202 3367 2206
rect 3371 2202 3463 2206
rect 3467 2202 3487 2206
rect 1785 2201 3487 2202
rect 3493 2201 3494 2207
rect 84 2137 85 2143
rect 91 2142 1779 2143
rect 91 2138 111 2142
rect 115 2138 303 2142
rect 307 2138 407 2142
rect 411 2138 439 2142
rect 443 2138 519 2142
rect 523 2138 527 2142
rect 531 2138 615 2142
rect 619 2138 631 2142
rect 635 2138 703 2142
rect 707 2138 743 2142
rect 747 2138 791 2142
rect 795 2138 863 2142
rect 867 2138 879 2142
rect 883 2138 967 2142
rect 971 2138 983 2142
rect 987 2138 1055 2142
rect 1059 2138 1143 2142
rect 1147 2138 1231 2142
rect 1235 2138 1319 2142
rect 1323 2138 1767 2142
rect 1771 2138 1779 2142
rect 91 2137 1779 2138
rect 1785 2137 1786 2143
rect 1790 2129 1791 2135
rect 1797 2134 3499 2135
rect 1797 2130 1807 2134
rect 1811 2130 2135 2134
rect 2139 2130 2183 2134
rect 2187 2130 2255 2134
rect 2259 2130 2279 2134
rect 2283 2130 2383 2134
rect 2387 2130 2495 2134
rect 2499 2130 2519 2134
rect 2523 2130 2607 2134
rect 2611 2130 2655 2134
rect 2659 2130 2719 2134
rect 2723 2130 2783 2134
rect 2787 2130 2839 2134
rect 2843 2130 2911 2134
rect 2915 2130 2967 2134
rect 2971 2130 3031 2134
rect 3035 2130 3103 2134
rect 3107 2130 3151 2134
rect 3155 2130 3247 2134
rect 3251 2130 3271 2134
rect 3275 2130 3367 2134
rect 3371 2130 3463 2134
rect 3467 2130 3499 2134
rect 1797 2129 3499 2130
rect 3505 2129 3506 2135
rect 96 2073 97 2079
rect 103 2078 1791 2079
rect 103 2074 111 2078
rect 115 2074 255 2078
rect 259 2074 303 2078
rect 307 2074 375 2078
rect 379 2074 407 2078
rect 411 2074 495 2078
rect 499 2074 519 2078
rect 523 2074 615 2078
rect 619 2074 631 2078
rect 635 2074 727 2078
rect 731 2074 743 2078
rect 747 2074 831 2078
rect 835 2074 863 2078
rect 867 2074 935 2078
rect 939 2074 983 2078
rect 987 2074 1039 2078
rect 1043 2074 1143 2078
rect 1147 2074 1255 2078
rect 1259 2074 1767 2078
rect 1771 2074 1791 2078
rect 103 2073 1791 2074
rect 1797 2073 1798 2079
rect 1778 2057 1779 2063
rect 1785 2062 3487 2063
rect 1785 2058 1807 2062
rect 1811 2058 2135 2062
rect 2139 2058 2247 2062
rect 2251 2058 2255 2062
rect 2259 2058 2383 2062
rect 2387 2058 2415 2062
rect 2419 2058 2519 2062
rect 2523 2058 2575 2062
rect 2579 2058 2655 2062
rect 2659 2058 2727 2062
rect 2731 2058 2783 2062
rect 2787 2058 2871 2062
rect 2875 2058 2911 2062
rect 2915 2058 3007 2062
rect 3011 2058 3031 2062
rect 3035 2058 3135 2062
rect 3139 2058 3151 2062
rect 3155 2058 3263 2062
rect 3267 2058 3271 2062
rect 3275 2058 3367 2062
rect 3371 2058 3463 2062
rect 3467 2058 3487 2062
rect 1785 2057 3487 2058
rect 3493 2057 3494 2063
rect 84 2009 85 2015
rect 91 2014 1779 2015
rect 91 2010 111 2014
rect 115 2010 255 2014
rect 259 2010 359 2014
rect 363 2010 375 2014
rect 379 2010 487 2014
rect 491 2010 495 2014
rect 499 2010 615 2014
rect 619 2010 623 2014
rect 627 2010 727 2014
rect 731 2010 759 2014
rect 763 2010 831 2014
rect 835 2010 895 2014
rect 899 2010 935 2014
rect 939 2010 1023 2014
rect 1027 2010 1039 2014
rect 1043 2010 1143 2014
rect 1147 2010 1151 2014
rect 1155 2010 1255 2014
rect 1259 2010 1271 2014
rect 1275 2010 1399 2014
rect 1403 2010 1527 2014
rect 1531 2010 1767 2014
rect 1771 2010 1779 2014
rect 91 2009 1779 2010
rect 1785 2009 1786 2015
rect 1790 1977 1791 1983
rect 1797 1982 3499 1983
rect 1797 1978 1807 1982
rect 1811 1978 1831 1982
rect 1835 1978 1919 1982
rect 1923 1978 2047 1982
rect 2051 1978 2183 1982
rect 2187 1978 2247 1982
rect 2251 1978 2327 1982
rect 2331 1978 2415 1982
rect 2419 1978 2471 1982
rect 2475 1978 2575 1982
rect 2579 1978 2615 1982
rect 2619 1978 2727 1982
rect 2731 1978 2751 1982
rect 2755 1978 2871 1982
rect 2875 1978 2887 1982
rect 2891 1978 3007 1982
rect 3011 1978 3031 1982
rect 3035 1978 3135 1982
rect 3139 1978 3175 1982
rect 3179 1978 3263 1982
rect 3267 1978 3319 1982
rect 3323 1978 3367 1982
rect 3371 1978 3463 1982
rect 3467 1978 3499 1982
rect 1797 1977 3499 1978
rect 3505 1977 3506 1983
rect 96 1945 97 1951
rect 103 1950 1791 1951
rect 103 1946 111 1950
rect 115 1946 359 1950
rect 363 1946 447 1950
rect 451 1946 487 1950
rect 491 1946 575 1950
rect 579 1946 623 1950
rect 627 1946 711 1950
rect 715 1946 759 1950
rect 763 1946 847 1950
rect 851 1946 895 1950
rect 899 1946 983 1950
rect 987 1946 1023 1950
rect 1027 1946 1119 1950
rect 1123 1946 1151 1950
rect 1155 1946 1255 1950
rect 1259 1946 1271 1950
rect 1275 1946 1383 1950
rect 1387 1946 1399 1950
rect 1403 1946 1519 1950
rect 1523 1946 1527 1950
rect 1531 1946 1655 1950
rect 1659 1946 1767 1950
rect 1771 1946 1791 1950
rect 103 1945 1791 1946
rect 1797 1945 1798 1951
rect 1778 1909 1779 1915
rect 1785 1914 3487 1915
rect 1785 1910 1807 1914
rect 1811 1910 1831 1914
rect 1835 1910 1919 1914
rect 1923 1910 2039 1914
rect 2043 1910 2047 1914
rect 2051 1910 2167 1914
rect 2171 1910 2183 1914
rect 2187 1910 2303 1914
rect 2307 1910 2327 1914
rect 2331 1910 2455 1914
rect 2459 1910 2471 1914
rect 2475 1910 2615 1914
rect 2619 1910 2751 1914
rect 2755 1910 2791 1914
rect 2795 1910 2887 1914
rect 2891 1910 2983 1914
rect 2987 1910 3031 1914
rect 3035 1910 3175 1914
rect 3179 1910 3183 1914
rect 3187 1910 3319 1914
rect 3323 1910 3367 1914
rect 3371 1910 3463 1914
rect 3467 1910 3487 1914
rect 1785 1909 3487 1910
rect 3493 1909 3494 1915
rect 84 1881 85 1887
rect 91 1886 1779 1887
rect 91 1882 111 1886
rect 115 1882 447 1886
rect 451 1882 559 1886
rect 563 1882 575 1886
rect 579 1882 695 1886
rect 699 1882 711 1886
rect 715 1882 831 1886
rect 835 1882 847 1886
rect 851 1882 959 1886
rect 963 1882 983 1886
rect 987 1882 1079 1886
rect 1083 1882 1119 1886
rect 1123 1882 1199 1886
rect 1203 1882 1255 1886
rect 1259 1882 1327 1886
rect 1331 1882 1383 1886
rect 1387 1882 1455 1886
rect 1459 1882 1519 1886
rect 1523 1882 1655 1886
rect 1659 1882 1767 1886
rect 1771 1882 1779 1886
rect 91 1881 1779 1882
rect 1785 1881 1786 1887
rect 1790 1841 1791 1847
rect 1797 1846 3499 1847
rect 1797 1842 1807 1846
rect 1811 1842 1831 1846
rect 1835 1842 1919 1846
rect 1923 1842 1959 1846
rect 1963 1842 2039 1846
rect 2043 1842 2111 1846
rect 2115 1842 2167 1846
rect 2171 1842 2255 1846
rect 2259 1842 2303 1846
rect 2307 1842 2407 1846
rect 2411 1842 2455 1846
rect 2459 1842 2567 1846
rect 2571 1842 2615 1846
rect 2619 1842 2743 1846
rect 2747 1842 2791 1846
rect 2795 1842 2935 1846
rect 2939 1842 2983 1846
rect 2987 1842 3135 1846
rect 3139 1842 3183 1846
rect 3187 1842 3343 1846
rect 3347 1842 3367 1846
rect 3371 1842 3463 1846
rect 3467 1842 3499 1846
rect 1797 1841 3499 1842
rect 3505 1841 3506 1847
rect 96 1809 97 1815
rect 103 1814 1791 1815
rect 103 1810 111 1814
rect 115 1810 135 1814
rect 139 1810 223 1814
rect 227 1810 311 1814
rect 315 1810 407 1814
rect 411 1810 527 1814
rect 531 1810 559 1814
rect 563 1810 655 1814
rect 659 1810 695 1814
rect 699 1810 799 1814
rect 803 1810 831 1814
rect 835 1810 943 1814
rect 947 1810 959 1814
rect 963 1810 1079 1814
rect 1083 1810 1087 1814
rect 1091 1810 1199 1814
rect 1203 1810 1239 1814
rect 1243 1810 1327 1814
rect 1331 1810 1391 1814
rect 1395 1810 1455 1814
rect 1459 1810 1543 1814
rect 1547 1810 1671 1814
rect 1675 1810 1767 1814
rect 1771 1810 1791 1814
rect 103 1809 1791 1810
rect 1797 1809 1798 1815
rect 1778 1765 1779 1771
rect 1785 1770 3487 1771
rect 1785 1766 1807 1770
rect 1811 1766 1831 1770
rect 1835 1766 1879 1770
rect 1883 1766 1959 1770
rect 1963 1766 2015 1770
rect 2019 1766 2111 1770
rect 2115 1766 2151 1770
rect 2155 1766 2255 1770
rect 2259 1766 2303 1770
rect 2307 1766 2407 1770
rect 2411 1766 2479 1770
rect 2483 1766 2567 1770
rect 2571 1766 2687 1770
rect 2691 1766 2743 1770
rect 2747 1766 2911 1770
rect 2915 1766 2935 1770
rect 2939 1766 3135 1770
rect 3139 1766 3151 1770
rect 3155 1766 3343 1770
rect 3347 1766 3367 1770
rect 3371 1766 3463 1770
rect 3467 1766 3487 1770
rect 1785 1765 3487 1766
rect 3493 1765 3494 1771
rect 84 1733 85 1739
rect 91 1738 1779 1739
rect 91 1734 111 1738
rect 115 1734 135 1738
rect 139 1734 223 1738
rect 227 1734 247 1738
rect 251 1734 311 1738
rect 315 1734 399 1738
rect 403 1734 407 1738
rect 411 1734 527 1738
rect 531 1734 567 1738
rect 571 1734 655 1738
rect 659 1734 751 1738
rect 755 1734 799 1738
rect 803 1734 935 1738
rect 939 1734 943 1738
rect 947 1734 1087 1738
rect 1091 1734 1119 1738
rect 1123 1734 1239 1738
rect 1243 1734 1311 1738
rect 1315 1734 1391 1738
rect 1395 1734 1503 1738
rect 1507 1734 1543 1738
rect 1547 1734 1671 1738
rect 1675 1734 1767 1738
rect 1771 1734 1779 1738
rect 91 1733 1779 1734
rect 1785 1733 1786 1739
rect 1790 1693 1791 1699
rect 1797 1698 3499 1699
rect 1797 1694 1807 1698
rect 1811 1694 1831 1698
rect 1835 1694 1879 1698
rect 1883 1694 1935 1698
rect 1939 1694 2015 1698
rect 2019 1694 2063 1698
rect 2067 1694 2151 1698
rect 2155 1694 2183 1698
rect 2187 1694 2303 1698
rect 2307 1694 2311 1698
rect 2315 1694 2439 1698
rect 2443 1694 2479 1698
rect 2483 1694 2575 1698
rect 2579 1694 2687 1698
rect 2691 1694 2727 1698
rect 2731 1694 2887 1698
rect 2891 1694 2911 1698
rect 2915 1694 3047 1698
rect 3051 1694 3151 1698
rect 3155 1694 3215 1698
rect 3219 1694 3367 1698
rect 3371 1694 3463 1698
rect 3467 1694 3499 1698
rect 1797 1693 3499 1694
rect 3505 1693 3506 1699
rect 96 1665 97 1671
rect 103 1670 1791 1671
rect 103 1666 111 1670
rect 115 1666 135 1670
rect 139 1666 191 1670
rect 195 1666 247 1670
rect 251 1666 295 1670
rect 299 1666 399 1670
rect 403 1666 407 1670
rect 411 1666 535 1670
rect 539 1666 567 1670
rect 571 1666 687 1670
rect 691 1666 751 1670
rect 755 1666 855 1670
rect 859 1666 935 1670
rect 939 1666 1039 1670
rect 1043 1666 1119 1670
rect 1123 1666 1231 1670
rect 1235 1666 1311 1670
rect 1315 1666 1431 1670
rect 1435 1666 1503 1670
rect 1507 1666 1639 1670
rect 1643 1666 1671 1670
rect 1675 1666 1767 1670
rect 1771 1666 1791 1670
rect 103 1665 1791 1666
rect 1797 1665 1798 1671
rect 1778 1621 1779 1627
rect 1785 1626 3487 1627
rect 1785 1622 1807 1626
rect 1811 1622 1831 1626
rect 1835 1622 1935 1626
rect 1939 1622 1943 1626
rect 1947 1622 2063 1626
rect 2067 1622 2087 1626
rect 2091 1622 2183 1626
rect 2187 1622 2231 1626
rect 2235 1622 2311 1626
rect 2315 1622 2367 1626
rect 2371 1622 2439 1626
rect 2443 1622 2503 1626
rect 2507 1622 2575 1626
rect 2579 1622 2639 1626
rect 2643 1622 2727 1626
rect 2731 1622 2767 1626
rect 2771 1622 2887 1626
rect 2891 1622 2895 1626
rect 2899 1622 3015 1626
rect 3019 1622 3047 1626
rect 3051 1622 3135 1626
rect 3139 1622 3215 1626
rect 3219 1622 3263 1626
rect 3267 1622 3367 1626
rect 3371 1622 3463 1626
rect 3467 1622 3487 1626
rect 1785 1621 3487 1622
rect 3493 1621 3494 1627
rect 84 1597 85 1603
rect 91 1602 1779 1603
rect 91 1598 111 1602
rect 115 1598 191 1602
rect 195 1598 295 1602
rect 299 1598 327 1602
rect 331 1598 407 1602
rect 411 1598 431 1602
rect 435 1598 535 1602
rect 539 1598 543 1602
rect 547 1598 671 1602
rect 675 1598 687 1602
rect 691 1598 815 1602
rect 819 1598 855 1602
rect 859 1598 967 1602
rect 971 1598 1039 1602
rect 1043 1598 1119 1602
rect 1123 1598 1231 1602
rect 1235 1598 1279 1602
rect 1283 1598 1431 1602
rect 1435 1598 1439 1602
rect 1443 1598 1607 1602
rect 1611 1598 1639 1602
rect 1643 1598 1767 1602
rect 1771 1598 1779 1602
rect 91 1597 1779 1598
rect 1785 1597 1786 1603
rect 1790 1549 1791 1555
rect 1797 1554 3499 1555
rect 1797 1550 1807 1554
rect 1811 1550 1831 1554
rect 1835 1550 1839 1554
rect 1843 1550 1943 1554
rect 1947 1550 1991 1554
rect 1995 1550 2087 1554
rect 2091 1550 2151 1554
rect 2155 1550 2231 1554
rect 2235 1550 2303 1554
rect 2307 1550 2367 1554
rect 2371 1550 2455 1554
rect 2459 1550 2503 1554
rect 2507 1550 2599 1554
rect 2603 1550 2639 1554
rect 2643 1550 2735 1554
rect 2739 1550 2767 1554
rect 2771 1550 2871 1554
rect 2875 1550 2895 1554
rect 2899 1550 3007 1554
rect 3011 1550 3015 1554
rect 3019 1550 3135 1554
rect 3139 1550 3143 1554
rect 3147 1550 3263 1554
rect 3267 1550 3367 1554
rect 3371 1550 3463 1554
rect 3467 1550 3499 1554
rect 1797 1549 3499 1550
rect 3505 1549 3506 1555
rect 96 1529 97 1535
rect 103 1534 1791 1535
rect 103 1530 111 1534
rect 115 1530 223 1534
rect 227 1530 327 1534
rect 331 1530 343 1534
rect 347 1530 431 1534
rect 435 1530 471 1534
rect 475 1530 543 1534
rect 547 1530 607 1534
rect 611 1530 671 1534
rect 675 1530 751 1534
rect 755 1530 815 1534
rect 819 1530 895 1534
rect 899 1530 967 1534
rect 971 1530 1047 1534
rect 1051 1530 1119 1534
rect 1123 1530 1199 1534
rect 1203 1530 1279 1534
rect 1283 1530 1351 1534
rect 1355 1530 1439 1534
rect 1443 1530 1503 1534
rect 1507 1530 1607 1534
rect 1611 1530 1767 1534
rect 1771 1530 1791 1534
rect 103 1529 1791 1530
rect 1797 1529 1798 1535
rect 1778 1477 1779 1483
rect 1785 1482 3487 1483
rect 1785 1478 1807 1482
rect 1811 1478 1839 1482
rect 1843 1478 1943 1482
rect 1947 1478 1991 1482
rect 1995 1478 2055 1482
rect 2059 1478 2151 1482
rect 2155 1478 2191 1482
rect 2195 1478 2303 1482
rect 2307 1478 2335 1482
rect 2339 1478 2455 1482
rect 2459 1478 2479 1482
rect 2483 1478 2599 1482
rect 2603 1478 2631 1482
rect 2635 1478 2735 1482
rect 2739 1478 2783 1482
rect 2787 1478 2871 1482
rect 2875 1478 2935 1482
rect 2939 1478 3007 1482
rect 3011 1478 3087 1482
rect 3091 1478 3143 1482
rect 3147 1478 3239 1482
rect 3243 1478 3463 1482
rect 3467 1478 3487 1482
rect 1785 1477 3487 1478
rect 3493 1477 3494 1483
rect 84 1457 85 1463
rect 91 1462 1779 1463
rect 91 1458 111 1462
rect 115 1458 135 1462
rect 139 1458 223 1462
rect 227 1458 303 1462
rect 307 1458 343 1462
rect 347 1458 471 1462
rect 475 1458 607 1462
rect 611 1458 631 1462
rect 635 1458 751 1462
rect 755 1458 783 1462
rect 787 1458 895 1462
rect 899 1458 927 1462
rect 931 1458 1047 1462
rect 1051 1458 1063 1462
rect 1067 1458 1199 1462
rect 1203 1458 1335 1462
rect 1339 1458 1351 1462
rect 1355 1458 1471 1462
rect 1475 1458 1503 1462
rect 1507 1458 1767 1462
rect 1771 1458 1779 1462
rect 91 1457 1779 1458
rect 1785 1457 1786 1463
rect 1790 1405 1791 1411
rect 1797 1410 3499 1411
rect 1797 1406 1807 1410
rect 1811 1406 1943 1410
rect 1947 1406 2055 1410
rect 2059 1406 2095 1410
rect 2099 1406 2191 1410
rect 2195 1406 2199 1410
rect 2203 1406 2319 1410
rect 2323 1406 2335 1410
rect 2339 1406 2455 1410
rect 2459 1406 2479 1410
rect 2483 1406 2599 1410
rect 2603 1406 2631 1410
rect 2635 1406 2743 1410
rect 2747 1406 2783 1410
rect 2787 1406 2887 1410
rect 2891 1406 2935 1410
rect 2939 1406 3031 1410
rect 3035 1406 3087 1410
rect 3091 1406 3175 1410
rect 3179 1406 3239 1410
rect 3243 1406 3327 1410
rect 3331 1406 3463 1410
rect 3467 1406 3499 1410
rect 1797 1405 3499 1406
rect 3505 1405 3506 1411
rect 96 1389 97 1395
rect 103 1394 1791 1395
rect 103 1390 111 1394
rect 115 1390 135 1394
rect 139 1390 279 1394
rect 283 1390 303 1394
rect 307 1390 447 1394
rect 451 1390 471 1394
rect 475 1390 607 1394
rect 611 1390 631 1394
rect 635 1390 759 1394
rect 763 1390 783 1394
rect 787 1390 903 1394
rect 907 1390 927 1394
rect 931 1390 1031 1394
rect 1035 1390 1063 1394
rect 1067 1390 1159 1394
rect 1163 1390 1199 1394
rect 1203 1390 1287 1394
rect 1291 1390 1335 1394
rect 1339 1390 1415 1394
rect 1419 1390 1471 1394
rect 1475 1390 1767 1394
rect 1771 1390 1791 1394
rect 103 1389 1791 1390
rect 1797 1389 1798 1395
rect 1778 1337 1779 1343
rect 1785 1342 3487 1343
rect 1785 1338 1807 1342
rect 1811 1338 2095 1342
rect 2099 1338 2103 1342
rect 2107 1338 2199 1342
rect 2203 1338 2239 1342
rect 2243 1338 2319 1342
rect 2323 1338 2383 1342
rect 2387 1338 2455 1342
rect 2459 1338 2535 1342
rect 2539 1338 2599 1342
rect 2603 1338 2687 1342
rect 2691 1338 2743 1342
rect 2747 1338 2839 1342
rect 2843 1338 2887 1342
rect 2891 1338 2991 1342
rect 2995 1338 3031 1342
rect 3035 1338 3143 1342
rect 3147 1338 3175 1342
rect 3179 1338 3303 1342
rect 3307 1338 3327 1342
rect 3331 1338 3463 1342
rect 3467 1338 3487 1342
rect 1785 1337 3487 1338
rect 3493 1337 3494 1343
rect 84 1321 85 1327
rect 91 1326 1779 1327
rect 91 1322 111 1326
rect 115 1322 135 1326
rect 139 1322 279 1326
rect 283 1322 439 1326
rect 443 1322 447 1326
rect 451 1322 583 1326
rect 587 1322 607 1326
rect 611 1322 719 1326
rect 723 1322 759 1326
rect 763 1322 847 1326
rect 851 1322 903 1326
rect 907 1322 967 1326
rect 971 1322 1031 1326
rect 1035 1322 1079 1326
rect 1083 1322 1159 1326
rect 1163 1322 1191 1326
rect 1195 1322 1287 1326
rect 1291 1322 1311 1326
rect 1315 1322 1415 1326
rect 1419 1322 1767 1326
rect 1771 1322 1779 1326
rect 91 1321 1779 1322
rect 1785 1321 1786 1327
rect 1790 1273 1791 1279
rect 1797 1278 3499 1279
rect 1797 1274 1807 1278
rect 1811 1274 1935 1278
rect 1939 1274 2063 1278
rect 2067 1274 2103 1278
rect 2107 1274 2199 1278
rect 2203 1274 2239 1278
rect 2243 1274 2343 1278
rect 2347 1274 2383 1278
rect 2387 1274 2495 1278
rect 2499 1274 2535 1278
rect 2539 1274 2655 1278
rect 2659 1274 2687 1278
rect 2691 1274 2815 1278
rect 2819 1274 2839 1278
rect 2843 1274 2975 1278
rect 2979 1274 2991 1278
rect 2995 1274 3143 1278
rect 3147 1274 3303 1278
rect 3307 1274 3463 1278
rect 3467 1274 3499 1278
rect 1797 1273 3499 1274
rect 3505 1273 3506 1279
rect 96 1253 97 1259
rect 103 1258 1791 1259
rect 103 1254 111 1258
rect 115 1254 135 1258
rect 139 1254 239 1258
rect 243 1254 279 1258
rect 283 1254 367 1258
rect 371 1254 439 1258
rect 443 1254 495 1258
rect 499 1254 583 1258
rect 587 1254 615 1258
rect 619 1254 719 1258
rect 723 1254 735 1258
rect 739 1254 847 1258
rect 851 1254 959 1258
rect 963 1254 967 1258
rect 971 1254 1071 1258
rect 1075 1254 1079 1258
rect 1083 1254 1191 1258
rect 1195 1254 1311 1258
rect 1315 1254 1767 1258
rect 1771 1254 1791 1258
rect 103 1253 1791 1254
rect 1797 1253 1798 1259
rect 1778 1209 1779 1215
rect 1785 1214 3487 1215
rect 1785 1210 1807 1214
rect 1811 1210 1831 1214
rect 1835 1210 1935 1214
rect 1939 1210 2063 1214
rect 2067 1210 2079 1214
rect 2083 1210 2199 1214
rect 2203 1210 2231 1214
rect 2235 1210 2343 1214
rect 2347 1210 2391 1214
rect 2395 1210 2495 1214
rect 2499 1210 2543 1214
rect 2547 1210 2655 1214
rect 2659 1210 2695 1214
rect 2699 1210 2815 1214
rect 2819 1210 2847 1214
rect 2851 1210 2975 1214
rect 2979 1210 2999 1214
rect 3003 1210 3143 1214
rect 3147 1210 3159 1214
rect 3163 1210 3463 1214
rect 3467 1210 3487 1214
rect 1785 1209 3487 1210
rect 3493 1209 3494 1215
rect 84 1185 85 1191
rect 91 1190 1779 1191
rect 91 1186 111 1190
rect 115 1186 135 1190
rect 139 1186 239 1190
rect 243 1186 367 1190
rect 371 1186 375 1190
rect 379 1186 495 1190
rect 499 1186 511 1190
rect 515 1186 615 1190
rect 619 1186 655 1190
rect 659 1186 735 1190
rect 739 1186 791 1190
rect 795 1186 847 1190
rect 851 1186 927 1190
rect 931 1186 959 1190
rect 963 1186 1063 1190
rect 1067 1186 1071 1190
rect 1075 1186 1191 1190
rect 1195 1186 1199 1190
rect 1203 1186 1335 1190
rect 1339 1186 1767 1190
rect 1771 1186 1779 1190
rect 91 1185 1779 1186
rect 1785 1185 1786 1191
rect 1790 1133 1791 1139
rect 1797 1138 3499 1139
rect 1797 1134 1807 1138
rect 1811 1134 1831 1138
rect 1835 1134 1863 1138
rect 1867 1134 1935 1138
rect 1939 1134 1983 1138
rect 1987 1134 2079 1138
rect 2083 1134 2111 1138
rect 2115 1134 2231 1138
rect 2235 1134 2247 1138
rect 2251 1134 2383 1138
rect 2387 1134 2391 1138
rect 2395 1134 2511 1138
rect 2515 1134 2543 1138
rect 2547 1134 2639 1138
rect 2643 1134 2695 1138
rect 2699 1134 2759 1138
rect 2763 1134 2847 1138
rect 2851 1134 2871 1138
rect 2875 1134 2975 1138
rect 2979 1134 2999 1138
rect 3003 1134 3079 1138
rect 3083 1134 3159 1138
rect 3163 1134 3183 1138
rect 3187 1134 3279 1138
rect 3283 1134 3367 1138
rect 3371 1134 3463 1138
rect 3467 1134 3499 1138
rect 1797 1133 3499 1134
rect 3505 1133 3506 1139
rect 96 1117 97 1123
rect 103 1122 1791 1123
rect 103 1118 111 1122
rect 115 1118 135 1122
rect 139 1118 191 1122
rect 195 1118 239 1122
rect 243 1118 335 1122
rect 339 1118 375 1122
rect 379 1118 495 1122
rect 499 1118 511 1122
rect 515 1118 655 1122
rect 659 1118 791 1122
rect 795 1118 815 1122
rect 819 1118 927 1122
rect 931 1118 967 1122
rect 971 1118 1063 1122
rect 1067 1118 1119 1122
rect 1123 1118 1199 1122
rect 1203 1118 1263 1122
rect 1267 1118 1335 1122
rect 1339 1118 1407 1122
rect 1411 1118 1559 1122
rect 1563 1118 1767 1122
rect 1771 1118 1791 1122
rect 103 1117 1791 1118
rect 1797 1117 1798 1123
rect 1778 1061 1779 1067
rect 1785 1066 3487 1067
rect 1785 1062 1807 1066
rect 1811 1062 1863 1066
rect 1867 1062 1983 1066
rect 1987 1062 2103 1066
rect 2107 1062 2111 1066
rect 2115 1062 2191 1066
rect 2195 1062 2247 1066
rect 2251 1062 2279 1066
rect 2283 1062 2367 1066
rect 2371 1062 2383 1066
rect 2387 1062 2455 1066
rect 2459 1062 2511 1066
rect 2515 1062 2543 1066
rect 2547 1062 2631 1066
rect 2635 1062 2639 1066
rect 2643 1062 2719 1066
rect 2723 1062 2759 1066
rect 2763 1062 2807 1066
rect 2811 1062 2871 1066
rect 2875 1062 2975 1066
rect 2979 1062 3079 1066
rect 3083 1062 3183 1066
rect 3187 1062 3279 1066
rect 3283 1062 3367 1066
rect 3371 1062 3463 1066
rect 3467 1062 3487 1066
rect 1785 1061 3487 1062
rect 3493 1061 3494 1067
rect 84 1045 85 1051
rect 91 1050 1779 1051
rect 91 1046 111 1050
rect 115 1046 191 1050
rect 195 1046 327 1050
rect 331 1046 335 1050
rect 339 1046 463 1050
rect 467 1046 495 1050
rect 499 1046 607 1050
rect 611 1046 655 1050
rect 659 1046 767 1050
rect 771 1046 815 1050
rect 819 1046 927 1050
rect 931 1046 967 1050
rect 971 1046 1079 1050
rect 1083 1046 1119 1050
rect 1123 1046 1231 1050
rect 1235 1046 1263 1050
rect 1267 1046 1383 1050
rect 1387 1046 1407 1050
rect 1411 1046 1535 1050
rect 1539 1046 1559 1050
rect 1563 1046 1671 1050
rect 1675 1046 1767 1050
rect 1771 1046 1779 1050
rect 91 1045 1779 1046
rect 1785 1045 1786 1051
rect 1790 997 1791 1003
rect 1797 1002 3499 1003
rect 1797 998 1807 1002
rect 1811 998 2103 1002
rect 2107 998 2191 1002
rect 2195 998 2279 1002
rect 2283 998 2311 1002
rect 2315 998 2367 1002
rect 2371 998 2407 1002
rect 2411 998 2455 1002
rect 2459 998 2511 1002
rect 2515 998 2543 1002
rect 2547 998 2623 1002
rect 2627 998 2631 1002
rect 2635 998 2719 1002
rect 2723 998 2751 1002
rect 2755 998 2807 1002
rect 2811 998 2895 1002
rect 2899 998 3055 1002
rect 3059 998 3223 1002
rect 3227 998 3367 1002
rect 3371 998 3463 1002
rect 3467 998 3499 1002
rect 1797 997 3499 998
rect 3505 997 3506 1003
rect 96 977 97 983
rect 103 982 1791 983
rect 103 978 111 982
rect 115 978 327 982
rect 331 978 463 982
rect 467 978 471 982
rect 475 978 567 982
rect 571 978 607 982
rect 611 978 671 982
rect 675 978 767 982
rect 771 978 783 982
rect 787 978 887 982
rect 891 978 927 982
rect 931 978 991 982
rect 995 978 1079 982
rect 1083 978 1095 982
rect 1099 978 1199 982
rect 1203 978 1231 982
rect 1235 978 1295 982
rect 1299 978 1383 982
rect 1387 978 1391 982
rect 1395 978 1487 982
rect 1491 978 1535 982
rect 1539 978 1583 982
rect 1587 978 1671 982
rect 1675 978 1767 982
rect 1771 978 1791 982
rect 103 977 1791 978
rect 1797 977 1798 983
rect 1778 921 1779 927
rect 1785 926 3487 927
rect 1785 922 1807 926
rect 1811 922 1831 926
rect 1835 922 1983 926
rect 1987 922 2151 926
rect 2155 922 2311 926
rect 2315 922 2327 926
rect 2331 922 2407 926
rect 2411 922 2511 926
rect 2515 922 2519 926
rect 2523 922 2623 926
rect 2627 922 2719 926
rect 2723 922 2751 926
rect 2755 922 2895 926
rect 2899 922 2935 926
rect 2939 922 3055 926
rect 3059 922 3159 926
rect 3163 922 3223 926
rect 3227 922 3367 926
rect 3371 922 3463 926
rect 3467 922 3487 926
rect 1785 921 3487 922
rect 3493 921 3494 927
rect 84 909 85 915
rect 91 914 1779 915
rect 91 910 111 914
rect 115 910 471 914
rect 475 910 567 914
rect 571 910 607 914
rect 611 910 671 914
rect 675 910 695 914
rect 699 910 783 914
rect 787 910 791 914
rect 795 910 887 914
rect 891 910 895 914
rect 899 910 991 914
rect 995 910 999 914
rect 1003 910 1095 914
rect 1099 910 1111 914
rect 1115 910 1199 914
rect 1203 910 1223 914
rect 1227 910 1295 914
rect 1299 910 1343 914
rect 1347 910 1391 914
rect 1395 910 1463 914
rect 1467 910 1487 914
rect 1491 910 1583 914
rect 1587 910 1671 914
rect 1675 910 1767 914
rect 1771 910 1779 914
rect 91 909 1779 910
rect 1785 909 1786 915
rect 1790 853 1791 859
rect 1797 858 3499 859
rect 1797 854 1807 858
rect 1811 854 1831 858
rect 1835 854 1959 858
rect 1963 854 1983 858
rect 1987 854 2087 858
rect 2091 854 2151 858
rect 2155 854 2207 858
rect 2211 854 2327 858
rect 2331 854 2463 858
rect 2467 854 2519 858
rect 2523 854 2615 858
rect 2619 854 2719 858
rect 2723 854 2791 858
rect 2795 854 2935 858
rect 2939 854 2983 858
rect 2987 854 3159 858
rect 3163 854 3183 858
rect 3187 854 3367 858
rect 3371 854 3463 858
rect 3467 854 3499 858
rect 1797 853 3499 854
rect 3505 853 3506 859
rect 96 841 97 847
rect 103 846 1791 847
rect 103 842 111 846
rect 115 842 519 846
rect 523 842 607 846
rect 611 842 615 846
rect 619 842 695 846
rect 699 842 719 846
rect 723 842 791 846
rect 795 842 831 846
rect 835 842 895 846
rect 899 842 951 846
rect 955 842 999 846
rect 1003 842 1071 846
rect 1075 842 1111 846
rect 1115 842 1191 846
rect 1195 842 1223 846
rect 1227 842 1311 846
rect 1315 842 1343 846
rect 1347 842 1431 846
rect 1435 842 1463 846
rect 1467 842 1559 846
rect 1563 842 1583 846
rect 1587 842 1767 846
rect 1771 842 1791 846
rect 103 841 1791 842
rect 1797 841 1798 847
rect 1778 785 1779 791
rect 1785 790 3487 791
rect 1785 786 1807 790
rect 1811 786 1831 790
rect 1835 786 1879 790
rect 1883 786 1959 790
rect 1963 786 2015 790
rect 2019 786 2087 790
rect 2091 786 2151 790
rect 2155 786 2207 790
rect 2211 786 2287 790
rect 2291 786 2327 790
rect 2331 786 2423 790
rect 2427 786 2463 790
rect 2467 786 2559 790
rect 2563 786 2615 790
rect 2619 786 2711 790
rect 2715 786 2791 790
rect 2795 786 2871 790
rect 2875 786 2983 790
rect 2987 786 3039 790
rect 3043 786 3183 790
rect 3187 786 3215 790
rect 3219 786 3367 790
rect 3371 786 3463 790
rect 3467 786 3487 790
rect 1785 785 3487 786
rect 3493 785 3494 791
rect 84 773 85 779
rect 91 778 1779 779
rect 91 774 111 778
rect 115 774 383 778
rect 387 774 471 778
rect 475 774 519 778
rect 523 774 575 778
rect 579 774 615 778
rect 619 774 679 778
rect 683 774 719 778
rect 723 774 791 778
rect 795 774 831 778
rect 835 774 911 778
rect 915 774 951 778
rect 955 774 1031 778
rect 1035 774 1071 778
rect 1075 774 1159 778
rect 1163 774 1191 778
rect 1195 774 1287 778
rect 1291 774 1311 778
rect 1315 774 1415 778
rect 1419 774 1431 778
rect 1435 774 1559 778
rect 1563 774 1767 778
rect 1771 774 1779 778
rect 91 773 1779 774
rect 1785 773 1786 779
rect 1790 717 1791 723
rect 1797 722 3499 723
rect 1797 718 1807 722
rect 1811 718 1831 722
rect 1835 718 1879 722
rect 1883 718 1951 722
rect 1955 718 2015 722
rect 2019 718 2103 722
rect 2107 718 2151 722
rect 2155 718 2263 722
rect 2267 718 2287 722
rect 2291 718 2415 722
rect 2419 718 2423 722
rect 2427 718 2559 722
rect 2563 718 2567 722
rect 2571 718 2711 722
rect 2715 718 2719 722
rect 2723 718 2871 722
rect 2875 718 2879 722
rect 2883 718 3039 722
rect 3043 718 3199 722
rect 3203 718 3215 722
rect 3219 718 3367 722
rect 3371 718 3463 722
rect 3467 718 3499 722
rect 1797 717 3499 718
rect 3505 717 3506 723
rect 96 701 97 707
rect 103 706 1791 707
rect 103 702 111 706
rect 115 702 247 706
rect 251 702 343 706
rect 347 702 383 706
rect 387 702 455 706
rect 459 702 471 706
rect 475 702 567 706
rect 571 702 575 706
rect 579 702 679 706
rect 683 702 695 706
rect 699 702 791 706
rect 795 702 831 706
rect 835 702 911 706
rect 915 702 983 706
rect 987 702 1031 706
rect 1035 702 1151 706
rect 1155 702 1159 706
rect 1163 702 1287 706
rect 1291 702 1327 706
rect 1331 702 1415 706
rect 1419 702 1511 706
rect 1515 702 1671 706
rect 1675 702 1767 706
rect 1771 702 1791 706
rect 103 701 1791 702
rect 1797 701 1798 707
rect 1778 653 1779 659
rect 1785 658 3487 659
rect 1785 654 1807 658
rect 1811 654 1831 658
rect 1835 654 1951 658
rect 1955 654 1975 658
rect 1979 654 2103 658
rect 2107 654 2239 658
rect 2243 654 2263 658
rect 2267 654 2415 658
rect 2419 654 2479 658
rect 2483 654 2567 658
rect 2571 654 2687 658
rect 2691 654 2719 658
rect 2723 654 2879 658
rect 2883 654 3039 658
rect 3043 654 3055 658
rect 3059 654 3199 658
rect 3203 654 3223 658
rect 3227 654 3367 658
rect 3371 654 3463 658
rect 3467 654 3487 658
rect 1785 653 3487 654
rect 3493 653 3494 659
rect 84 633 85 639
rect 91 638 1779 639
rect 91 634 111 638
rect 115 634 135 638
rect 139 634 231 638
rect 235 634 247 638
rect 251 634 343 638
rect 347 634 359 638
rect 363 634 455 638
rect 459 634 487 638
rect 491 634 567 638
rect 571 634 623 638
rect 627 634 695 638
rect 699 634 767 638
rect 771 634 831 638
rect 835 634 911 638
rect 915 634 983 638
rect 987 634 1055 638
rect 1059 634 1151 638
rect 1155 634 1207 638
rect 1211 634 1327 638
rect 1331 634 1367 638
rect 1371 634 1511 638
rect 1515 634 1527 638
rect 1531 634 1671 638
rect 1675 634 1767 638
rect 1771 634 1779 638
rect 91 633 1779 634
rect 1785 633 1786 639
rect 1790 581 1791 587
rect 1797 586 3499 587
rect 1797 582 1807 586
rect 1811 582 1895 586
rect 1899 582 1975 586
rect 1979 582 2015 586
rect 2019 582 2143 586
rect 2147 582 2239 586
rect 2243 582 2279 586
rect 2283 582 2423 586
rect 2427 582 2479 586
rect 2483 582 2567 586
rect 2571 582 2687 586
rect 2691 582 2719 586
rect 2723 582 2871 586
rect 2875 582 2879 586
rect 2883 582 3031 586
rect 3035 582 3055 586
rect 3059 582 3199 586
rect 3203 582 3223 586
rect 3227 582 3367 586
rect 3371 582 3463 586
rect 3467 582 3499 586
rect 1797 581 3499 582
rect 3505 581 3506 587
rect 96 565 97 571
rect 103 570 1791 571
rect 103 566 111 570
rect 115 566 135 570
rect 139 566 231 570
rect 235 566 247 570
rect 251 566 359 570
rect 363 566 407 570
rect 411 566 487 570
rect 491 566 583 570
rect 587 566 623 570
rect 627 566 767 570
rect 771 566 911 570
rect 915 566 951 570
rect 955 566 1055 570
rect 1059 566 1135 570
rect 1139 566 1207 570
rect 1211 566 1319 570
rect 1323 566 1367 570
rect 1371 566 1503 570
rect 1507 566 1527 570
rect 1531 566 1671 570
rect 1675 566 1767 570
rect 1771 566 1791 570
rect 103 565 1791 566
rect 1797 565 1798 571
rect 1778 513 1779 519
rect 1785 518 3487 519
rect 1785 514 1807 518
rect 1811 514 1895 518
rect 1899 514 2015 518
rect 2019 514 2135 518
rect 2139 514 2143 518
rect 2147 514 2239 518
rect 2243 514 2279 518
rect 2283 514 2359 518
rect 2363 514 2423 518
rect 2427 514 2487 518
rect 2491 514 2567 518
rect 2571 514 2615 518
rect 2619 514 2719 518
rect 2723 514 2751 518
rect 2755 514 2871 518
rect 2875 514 2879 518
rect 2883 514 3007 518
rect 3011 514 3031 518
rect 3035 514 3135 518
rect 3139 514 3199 518
rect 3203 514 3263 518
rect 3267 514 3367 518
rect 3371 514 3463 518
rect 3467 514 3487 518
rect 1785 513 3487 514
rect 3493 513 3494 519
rect 84 497 85 503
rect 91 502 1779 503
rect 91 498 111 502
rect 115 498 135 502
rect 139 498 247 502
rect 251 498 399 502
rect 403 498 407 502
rect 411 498 567 502
rect 571 498 583 502
rect 587 498 735 502
rect 739 498 767 502
rect 771 498 903 502
rect 907 498 951 502
rect 955 498 1063 502
rect 1067 498 1135 502
rect 1139 498 1223 502
rect 1227 498 1319 502
rect 1323 498 1375 502
rect 1379 498 1503 502
rect 1507 498 1527 502
rect 1531 498 1671 502
rect 1675 498 1767 502
rect 1771 498 1779 502
rect 91 497 1779 498
rect 1785 497 1786 503
rect 1790 441 1791 447
rect 1797 446 3499 447
rect 1797 442 1807 446
rect 1811 442 2135 446
rect 2139 442 2239 446
rect 2243 442 2335 446
rect 2339 442 2359 446
rect 2363 442 2447 446
rect 2451 442 2487 446
rect 2491 442 2559 446
rect 2563 442 2615 446
rect 2619 442 2679 446
rect 2683 442 2751 446
rect 2755 442 2799 446
rect 2803 442 2879 446
rect 2883 442 2911 446
rect 2915 442 3007 446
rect 3011 442 3023 446
rect 3027 442 3135 446
rect 3139 442 3143 446
rect 3147 442 3263 446
rect 3267 442 3367 446
rect 3371 442 3463 446
rect 3467 442 3499 446
rect 1797 441 3499 442
rect 3505 441 3506 447
rect 96 429 97 435
rect 103 434 1791 435
rect 103 430 111 434
rect 115 430 247 434
rect 251 430 399 434
rect 403 430 519 434
rect 523 430 567 434
rect 571 430 615 434
rect 619 430 719 434
rect 723 430 735 434
rect 739 430 823 434
rect 827 430 903 434
rect 907 430 927 434
rect 931 430 1023 434
rect 1027 430 1063 434
rect 1067 430 1127 434
rect 1131 430 1223 434
rect 1227 430 1231 434
rect 1235 430 1335 434
rect 1339 430 1375 434
rect 1379 430 1439 434
rect 1443 430 1527 434
rect 1531 430 1671 434
rect 1675 430 1767 434
rect 1771 430 1791 434
rect 103 429 1791 430
rect 1797 429 1798 435
rect 1778 373 1779 379
rect 1785 378 3487 379
rect 1785 374 1807 378
rect 1811 374 2063 378
rect 2067 374 2151 378
rect 2155 374 2239 378
rect 2243 374 2247 378
rect 2251 374 2335 378
rect 2339 374 2359 378
rect 2363 374 2447 378
rect 2451 374 2479 378
rect 2483 374 2559 378
rect 2563 374 2615 378
rect 2619 374 2679 378
rect 2683 374 2759 378
rect 2763 374 2799 378
rect 2803 374 2911 378
rect 2915 374 3023 378
rect 3027 374 3063 378
rect 3067 374 3143 378
rect 3147 374 3223 378
rect 3227 374 3263 378
rect 3267 374 3367 378
rect 3371 374 3463 378
rect 3467 374 3487 378
rect 1785 373 3487 374
rect 3493 373 3494 379
rect 84 361 85 367
rect 91 366 1779 367
rect 91 362 111 366
rect 115 362 471 366
rect 475 362 519 366
rect 523 362 559 366
rect 563 362 615 366
rect 619 362 647 366
rect 651 362 719 366
rect 723 362 735 366
rect 739 362 823 366
rect 827 362 911 366
rect 915 362 927 366
rect 931 362 999 366
rect 1003 362 1023 366
rect 1027 362 1087 366
rect 1091 362 1127 366
rect 1131 362 1175 366
rect 1179 362 1231 366
rect 1235 362 1263 366
rect 1267 362 1335 366
rect 1339 362 1439 366
rect 1443 362 1767 366
rect 1771 362 1779 366
rect 91 361 1779 362
rect 1785 361 1786 367
rect 1790 305 1791 311
rect 1797 310 3499 311
rect 1797 306 1807 310
rect 1811 306 1927 310
rect 1931 306 2039 310
rect 2043 306 2063 310
rect 2067 306 2151 310
rect 2155 306 2167 310
rect 2171 306 2247 310
rect 2251 306 2303 310
rect 2307 306 2359 310
rect 2363 306 2447 310
rect 2451 306 2479 310
rect 2483 306 2599 310
rect 2603 306 2615 310
rect 2619 306 2759 310
rect 2763 306 2911 310
rect 2915 306 2919 310
rect 2923 306 3063 310
rect 3067 306 3087 310
rect 3091 306 3223 310
rect 3227 306 3255 310
rect 3259 306 3367 310
rect 3371 306 3463 310
rect 3467 306 3499 310
rect 1797 305 3499 306
rect 3505 305 3506 311
rect 96 293 97 299
rect 103 298 1791 299
rect 103 294 111 298
rect 115 294 279 298
rect 283 294 367 298
rect 371 294 463 298
rect 467 294 471 298
rect 475 294 559 298
rect 563 294 647 298
rect 651 294 655 298
rect 659 294 735 298
rect 739 294 751 298
rect 755 294 823 298
rect 827 294 847 298
rect 851 294 911 298
rect 915 294 943 298
rect 947 294 999 298
rect 1003 294 1047 298
rect 1051 294 1087 298
rect 1091 294 1151 298
rect 1155 294 1175 298
rect 1179 294 1263 298
rect 1267 294 1767 298
rect 1771 294 1791 298
rect 103 293 1791 294
rect 1797 293 1798 299
rect 1778 237 1779 243
rect 1785 242 3487 243
rect 1785 238 1807 242
rect 1811 238 1831 242
rect 1835 238 1927 242
rect 1931 238 2039 242
rect 2043 238 2055 242
rect 2059 238 2167 242
rect 2171 238 2199 242
rect 2203 238 2303 242
rect 2307 238 2351 242
rect 2355 238 2447 242
rect 2451 238 2511 242
rect 2515 238 2599 242
rect 2603 238 2679 242
rect 2683 238 2759 242
rect 2763 238 2847 242
rect 2851 238 2919 242
rect 2923 238 3023 242
rect 3027 238 3087 242
rect 3091 238 3207 242
rect 3211 238 3255 242
rect 3259 238 3367 242
rect 3371 238 3463 242
rect 3467 238 3487 242
rect 1785 237 3487 238
rect 3493 237 3494 243
rect 84 225 85 231
rect 91 230 1779 231
rect 91 226 111 230
rect 115 226 167 230
rect 171 226 279 230
rect 283 226 343 230
rect 347 226 367 230
rect 371 226 463 230
rect 467 226 511 230
rect 515 226 559 230
rect 563 226 655 230
rect 659 226 679 230
rect 683 226 751 230
rect 755 226 839 230
rect 843 226 847 230
rect 851 226 943 230
rect 947 226 991 230
rect 995 226 1047 230
rect 1051 226 1135 230
rect 1139 226 1151 230
rect 1155 226 1279 230
rect 1283 226 1431 230
rect 1435 226 1767 230
rect 1771 226 1779 230
rect 91 225 1779 226
rect 1785 225 1786 231
rect 1790 153 1791 159
rect 1797 158 3499 159
rect 1797 154 1807 158
rect 1811 154 1831 158
rect 1835 154 1919 158
rect 1923 154 1927 158
rect 1931 154 2039 158
rect 2043 154 2055 158
rect 2059 154 2159 158
rect 2163 154 2199 158
rect 2203 154 2279 158
rect 2283 154 2351 158
rect 2355 154 2399 158
rect 2403 154 2511 158
rect 2515 154 2623 158
rect 2627 154 2679 158
rect 2683 154 2735 158
rect 2739 154 2839 158
rect 2843 154 2847 158
rect 2851 154 2943 158
rect 2947 154 3023 158
rect 3027 154 3055 158
rect 3059 154 3167 158
rect 3171 154 3207 158
rect 3211 154 3279 158
rect 3283 154 3367 158
rect 3371 154 3463 158
rect 3467 154 3499 158
rect 1797 153 3499 154
rect 3505 153 3506 159
rect 96 137 97 143
rect 103 142 1791 143
rect 103 138 111 142
rect 115 138 135 142
rect 139 138 167 142
rect 171 138 223 142
rect 227 138 311 142
rect 315 138 343 142
rect 347 138 399 142
rect 403 138 487 142
rect 491 138 511 142
rect 515 138 575 142
rect 579 138 663 142
rect 667 138 679 142
rect 683 138 751 142
rect 755 138 839 142
rect 843 138 847 142
rect 851 138 943 142
rect 947 138 991 142
rect 995 138 1031 142
rect 1035 138 1119 142
rect 1123 138 1135 142
rect 1139 138 1215 142
rect 1219 138 1279 142
rect 1283 138 1311 142
rect 1315 138 1407 142
rect 1411 138 1431 142
rect 1435 138 1495 142
rect 1499 138 1583 142
rect 1587 138 1671 142
rect 1675 138 1767 142
rect 1771 138 1791 142
rect 103 137 1791 138
rect 1797 137 1798 143
rect 1778 89 1779 95
rect 1785 94 3487 95
rect 1785 90 1807 94
rect 1811 90 1831 94
rect 1835 90 1919 94
rect 1923 90 2039 94
rect 2043 90 2159 94
rect 2163 90 2279 94
rect 2283 90 2399 94
rect 2403 90 2511 94
rect 2515 90 2623 94
rect 2627 90 2735 94
rect 2739 90 2839 94
rect 2843 90 2943 94
rect 2947 90 3055 94
rect 3059 90 3167 94
rect 3171 90 3279 94
rect 3283 90 3367 94
rect 3371 90 3463 94
rect 3467 90 3487 94
rect 1785 89 3487 90
rect 3493 89 3494 95
rect 84 73 85 79
rect 91 78 1779 79
rect 91 74 111 78
rect 115 74 135 78
rect 139 74 223 78
rect 227 74 311 78
rect 315 74 399 78
rect 403 74 487 78
rect 491 74 575 78
rect 579 74 663 78
rect 667 74 751 78
rect 755 74 847 78
rect 851 74 943 78
rect 947 74 1031 78
rect 1035 74 1119 78
rect 1123 74 1215 78
rect 1219 74 1311 78
rect 1315 74 1407 78
rect 1411 74 1495 78
rect 1499 74 1583 78
rect 1587 74 1671 78
rect 1675 74 1767 78
rect 1771 74 1779 78
rect 91 73 1779 74
rect 1785 73 1786 79
<< m5c >>
rect 1791 3517 1797 3523
rect 3499 3517 3505 3523
rect 97 3481 103 3487
rect 1791 3481 1797 3487
rect 1779 3453 1785 3459
rect 3487 3453 3493 3459
rect 85 3417 91 3423
rect 1779 3417 1785 3423
rect 1791 3381 1797 3387
rect 3499 3381 3505 3387
rect 97 3349 103 3355
rect 1791 3349 1797 3355
rect 1779 3309 1785 3315
rect 3487 3309 3493 3315
rect 85 3281 91 3287
rect 1779 3281 1785 3287
rect 1791 3237 1797 3243
rect 3499 3237 3505 3243
rect 97 3213 103 3219
rect 1791 3213 1797 3219
rect 1779 3173 1785 3179
rect 3487 3173 3493 3179
rect 85 3137 91 3143
rect 1779 3137 1785 3143
rect 1791 3105 1797 3111
rect 3499 3105 3505 3111
rect 97 3065 103 3071
rect 1791 3065 1797 3071
rect 1779 3033 1785 3039
rect 3487 3033 3493 3039
rect 85 2997 91 3003
rect 1779 2997 1785 3003
rect 1791 2969 1797 2975
rect 3499 2969 3505 2975
rect 97 2925 103 2931
rect 1791 2925 1797 2931
rect 1779 2897 1785 2903
rect 3487 2897 3493 2903
rect 85 2857 91 2863
rect 1779 2857 1785 2863
rect 1791 2829 1797 2835
rect 3499 2829 3505 2835
rect 97 2785 103 2791
rect 1791 2785 1797 2791
rect 1779 2761 1785 2767
rect 3487 2761 3493 2767
rect 85 2717 91 2723
rect 1779 2717 1785 2723
rect 1791 2697 1797 2703
rect 3499 2697 3505 2703
rect 97 2645 103 2651
rect 1791 2645 1797 2651
rect 1779 2629 1785 2635
rect 3487 2629 3493 2635
rect 85 2569 91 2575
rect 1779 2569 1785 2575
rect 1791 2557 1797 2563
rect 3499 2557 3505 2563
rect 97 2505 103 2511
rect 1791 2505 1797 2511
rect 1779 2477 1785 2483
rect 3487 2477 3493 2483
rect 85 2425 91 2431
rect 1779 2425 1785 2431
rect 1791 2409 1797 2415
rect 3499 2409 3505 2415
rect 1779 2363 1785 2369
rect 97 2353 103 2359
rect 1791 2353 1797 2359
rect 3487 2345 3493 2351
rect 85 2281 91 2287
rect 1779 2281 1785 2287
rect 1791 2277 1797 2283
rect 3499 2277 3505 2283
rect 97 2217 103 2223
rect 1791 2217 1797 2223
rect 1779 2201 1785 2207
rect 3487 2201 3493 2207
rect 85 2137 91 2143
rect 1779 2137 1785 2143
rect 1791 2129 1797 2135
rect 3499 2129 3505 2135
rect 97 2073 103 2079
rect 1791 2073 1797 2079
rect 1779 2057 1785 2063
rect 3487 2057 3493 2063
rect 85 2009 91 2015
rect 1779 2009 1785 2015
rect 1791 1977 1797 1983
rect 3499 1977 3505 1983
rect 97 1945 103 1951
rect 1791 1945 1797 1951
rect 1779 1909 1785 1915
rect 3487 1909 3493 1915
rect 85 1881 91 1887
rect 1779 1881 1785 1887
rect 1791 1841 1797 1847
rect 3499 1841 3505 1847
rect 97 1809 103 1815
rect 1791 1809 1797 1815
rect 1779 1765 1785 1771
rect 3487 1765 3493 1771
rect 85 1733 91 1739
rect 1779 1733 1785 1739
rect 1791 1693 1797 1699
rect 3499 1693 3505 1699
rect 97 1665 103 1671
rect 1791 1665 1797 1671
rect 1779 1621 1785 1627
rect 3487 1621 3493 1627
rect 85 1597 91 1603
rect 1779 1597 1785 1603
rect 1791 1549 1797 1555
rect 3499 1549 3505 1555
rect 97 1529 103 1535
rect 1791 1529 1797 1535
rect 1779 1477 1785 1483
rect 3487 1477 3493 1483
rect 85 1457 91 1463
rect 1779 1457 1785 1463
rect 1791 1405 1797 1411
rect 3499 1405 3505 1411
rect 97 1389 103 1395
rect 1791 1389 1797 1395
rect 1779 1337 1785 1343
rect 3487 1337 3493 1343
rect 85 1321 91 1327
rect 1779 1321 1785 1327
rect 1791 1273 1797 1279
rect 3499 1273 3505 1279
rect 97 1253 103 1259
rect 1791 1253 1797 1259
rect 1779 1209 1785 1215
rect 3487 1209 3493 1215
rect 85 1185 91 1191
rect 1779 1185 1785 1191
rect 1791 1133 1797 1139
rect 3499 1133 3505 1139
rect 97 1117 103 1123
rect 1791 1117 1797 1123
rect 1779 1061 1785 1067
rect 3487 1061 3493 1067
rect 85 1045 91 1051
rect 1779 1045 1785 1051
rect 1791 997 1797 1003
rect 3499 997 3505 1003
rect 97 977 103 983
rect 1791 977 1797 983
rect 1779 921 1785 927
rect 3487 921 3493 927
rect 85 909 91 915
rect 1779 909 1785 915
rect 1791 853 1797 859
rect 3499 853 3505 859
rect 97 841 103 847
rect 1791 841 1797 847
rect 1779 785 1785 791
rect 3487 785 3493 791
rect 85 773 91 779
rect 1779 773 1785 779
rect 1791 717 1797 723
rect 3499 717 3505 723
rect 97 701 103 707
rect 1791 701 1797 707
rect 1779 653 1785 659
rect 3487 653 3493 659
rect 85 633 91 639
rect 1779 633 1785 639
rect 1791 581 1797 587
rect 3499 581 3505 587
rect 97 565 103 571
rect 1791 565 1797 571
rect 1779 513 1785 519
rect 3487 513 3493 519
rect 85 497 91 503
rect 1779 497 1785 503
rect 1791 441 1797 447
rect 3499 441 3505 447
rect 97 429 103 435
rect 1791 429 1797 435
rect 1779 373 1785 379
rect 3487 373 3493 379
rect 85 361 91 367
rect 1779 361 1785 367
rect 1791 305 1797 311
rect 3499 305 3505 311
rect 97 293 103 299
rect 1791 293 1797 299
rect 1779 237 1785 243
rect 3487 237 3493 243
rect 85 225 91 231
rect 1779 225 1785 231
rect 1791 153 1797 159
rect 3499 153 3505 159
rect 97 137 103 143
rect 1791 137 1797 143
rect 1779 89 1785 95
rect 3487 89 3493 95
rect 85 73 91 79
rect 1779 73 1785 79
<< m5 >>
rect 84 3423 92 3528
rect 84 3417 85 3423
rect 91 3417 92 3423
rect 84 3287 92 3417
rect 84 3281 85 3287
rect 91 3281 92 3287
rect 84 3143 92 3281
rect 84 3137 85 3143
rect 91 3137 92 3143
rect 84 3003 92 3137
rect 84 2997 85 3003
rect 91 2997 92 3003
rect 84 2863 92 2997
rect 84 2857 85 2863
rect 91 2857 92 2863
rect 84 2723 92 2857
rect 84 2717 85 2723
rect 91 2717 92 2723
rect 84 2575 92 2717
rect 84 2569 85 2575
rect 91 2569 92 2575
rect 84 2431 92 2569
rect 84 2425 85 2431
rect 91 2425 92 2431
rect 84 2287 92 2425
rect 84 2281 85 2287
rect 91 2281 92 2287
rect 84 2143 92 2281
rect 84 2137 85 2143
rect 91 2137 92 2143
rect 84 2015 92 2137
rect 84 2009 85 2015
rect 91 2009 92 2015
rect 84 1887 92 2009
rect 84 1881 85 1887
rect 91 1881 92 1887
rect 84 1739 92 1881
rect 84 1733 85 1739
rect 91 1733 92 1739
rect 84 1603 92 1733
rect 84 1597 85 1603
rect 91 1597 92 1603
rect 84 1463 92 1597
rect 84 1457 85 1463
rect 91 1457 92 1463
rect 84 1327 92 1457
rect 84 1321 85 1327
rect 91 1321 92 1327
rect 84 1191 92 1321
rect 84 1185 85 1191
rect 91 1185 92 1191
rect 84 1051 92 1185
rect 84 1045 85 1051
rect 91 1045 92 1051
rect 84 915 92 1045
rect 84 909 85 915
rect 91 909 92 915
rect 84 779 92 909
rect 84 773 85 779
rect 91 773 92 779
rect 84 639 92 773
rect 84 633 85 639
rect 91 633 92 639
rect 84 503 92 633
rect 84 497 85 503
rect 91 497 92 503
rect 84 367 92 497
rect 84 361 85 367
rect 91 361 92 367
rect 84 231 92 361
rect 84 225 85 231
rect 91 225 92 231
rect 84 79 92 225
rect 84 73 85 79
rect 91 73 92 79
rect 84 72 92 73
rect 96 3487 104 3528
rect 96 3481 97 3487
rect 103 3481 104 3487
rect 96 3355 104 3481
rect 96 3349 97 3355
rect 103 3349 104 3355
rect 96 3219 104 3349
rect 96 3213 97 3219
rect 103 3213 104 3219
rect 96 3071 104 3213
rect 96 3065 97 3071
rect 103 3065 104 3071
rect 96 2931 104 3065
rect 96 2925 97 2931
rect 103 2925 104 2931
rect 96 2791 104 2925
rect 96 2785 97 2791
rect 103 2785 104 2791
rect 96 2651 104 2785
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2511 104 2645
rect 96 2505 97 2511
rect 103 2505 104 2511
rect 96 2359 104 2505
rect 96 2353 97 2359
rect 103 2353 104 2359
rect 96 2223 104 2353
rect 96 2217 97 2223
rect 103 2217 104 2223
rect 96 2079 104 2217
rect 96 2073 97 2079
rect 103 2073 104 2079
rect 96 1951 104 2073
rect 96 1945 97 1951
rect 103 1945 104 1951
rect 96 1815 104 1945
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1671 104 1809
rect 96 1665 97 1671
rect 103 1665 104 1671
rect 96 1535 104 1665
rect 96 1529 97 1535
rect 103 1529 104 1535
rect 96 1395 104 1529
rect 96 1389 97 1395
rect 103 1389 104 1395
rect 96 1259 104 1389
rect 96 1253 97 1259
rect 103 1253 104 1259
rect 96 1123 104 1253
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 983 104 1117
rect 96 977 97 983
rect 103 977 104 983
rect 96 847 104 977
rect 96 841 97 847
rect 103 841 104 847
rect 96 707 104 841
rect 96 701 97 707
rect 103 701 104 707
rect 96 571 104 701
rect 96 565 97 571
rect 103 565 104 571
rect 96 435 104 565
rect 96 429 97 435
rect 103 429 104 435
rect 96 299 104 429
rect 96 293 97 299
rect 103 293 104 299
rect 96 143 104 293
rect 96 137 97 143
rect 103 137 104 143
rect 96 72 104 137
rect 1778 3459 1786 3528
rect 1778 3453 1779 3459
rect 1785 3453 1786 3459
rect 1778 3423 1786 3453
rect 1778 3417 1779 3423
rect 1785 3417 1786 3423
rect 1778 3315 1786 3417
rect 1778 3309 1779 3315
rect 1785 3309 1786 3315
rect 1778 3287 1786 3309
rect 1778 3281 1779 3287
rect 1785 3281 1786 3287
rect 1778 3179 1786 3281
rect 1778 3173 1779 3179
rect 1785 3173 1786 3179
rect 1778 3143 1786 3173
rect 1778 3137 1779 3143
rect 1785 3137 1786 3143
rect 1778 3039 1786 3137
rect 1778 3033 1779 3039
rect 1785 3033 1786 3039
rect 1778 3003 1786 3033
rect 1778 2997 1779 3003
rect 1785 2997 1786 3003
rect 1778 2903 1786 2997
rect 1778 2897 1779 2903
rect 1785 2897 1786 2903
rect 1778 2863 1786 2897
rect 1778 2857 1779 2863
rect 1785 2857 1786 2863
rect 1778 2767 1786 2857
rect 1778 2761 1779 2767
rect 1785 2761 1786 2767
rect 1778 2723 1786 2761
rect 1778 2717 1779 2723
rect 1785 2717 1786 2723
rect 1778 2635 1786 2717
rect 1778 2629 1779 2635
rect 1785 2629 1786 2635
rect 1778 2575 1786 2629
rect 1778 2569 1779 2575
rect 1785 2569 1786 2575
rect 1778 2483 1786 2569
rect 1778 2477 1779 2483
rect 1785 2477 1786 2483
rect 1778 2431 1786 2477
rect 1778 2425 1779 2431
rect 1785 2425 1786 2431
rect 1778 2369 1786 2425
rect 1778 2363 1779 2369
rect 1785 2363 1786 2369
rect 1778 2287 1786 2363
rect 1778 2281 1779 2287
rect 1785 2281 1786 2287
rect 1778 2207 1786 2281
rect 1778 2201 1779 2207
rect 1785 2201 1786 2207
rect 1778 2143 1786 2201
rect 1778 2137 1779 2143
rect 1785 2137 1786 2143
rect 1778 2063 1786 2137
rect 1778 2057 1779 2063
rect 1785 2057 1786 2063
rect 1778 2015 1786 2057
rect 1778 2009 1779 2015
rect 1785 2009 1786 2015
rect 1778 1915 1786 2009
rect 1778 1909 1779 1915
rect 1785 1909 1786 1915
rect 1778 1887 1786 1909
rect 1778 1881 1779 1887
rect 1785 1881 1786 1887
rect 1778 1771 1786 1881
rect 1778 1765 1779 1771
rect 1785 1765 1786 1771
rect 1778 1739 1786 1765
rect 1778 1733 1779 1739
rect 1785 1733 1786 1739
rect 1778 1627 1786 1733
rect 1778 1621 1779 1627
rect 1785 1621 1786 1627
rect 1778 1603 1786 1621
rect 1778 1597 1779 1603
rect 1785 1597 1786 1603
rect 1778 1483 1786 1597
rect 1778 1477 1779 1483
rect 1785 1477 1786 1483
rect 1778 1463 1786 1477
rect 1778 1457 1779 1463
rect 1785 1457 1786 1463
rect 1778 1343 1786 1457
rect 1778 1337 1779 1343
rect 1785 1337 1786 1343
rect 1778 1327 1786 1337
rect 1778 1321 1779 1327
rect 1785 1321 1786 1327
rect 1778 1215 1786 1321
rect 1778 1209 1779 1215
rect 1785 1209 1786 1215
rect 1778 1191 1786 1209
rect 1778 1185 1779 1191
rect 1785 1185 1786 1191
rect 1778 1067 1786 1185
rect 1778 1061 1779 1067
rect 1785 1061 1786 1067
rect 1778 1051 1786 1061
rect 1778 1045 1779 1051
rect 1785 1045 1786 1051
rect 1778 927 1786 1045
rect 1778 921 1779 927
rect 1785 921 1786 927
rect 1778 915 1786 921
rect 1778 909 1779 915
rect 1785 909 1786 915
rect 1778 791 1786 909
rect 1778 785 1779 791
rect 1785 785 1786 791
rect 1778 779 1786 785
rect 1778 773 1779 779
rect 1785 773 1786 779
rect 1778 659 1786 773
rect 1778 653 1779 659
rect 1785 653 1786 659
rect 1778 639 1786 653
rect 1778 633 1779 639
rect 1785 633 1786 639
rect 1778 519 1786 633
rect 1778 513 1779 519
rect 1785 513 1786 519
rect 1778 503 1786 513
rect 1778 497 1779 503
rect 1785 497 1786 503
rect 1778 379 1786 497
rect 1778 373 1779 379
rect 1785 373 1786 379
rect 1778 367 1786 373
rect 1778 361 1779 367
rect 1785 361 1786 367
rect 1778 243 1786 361
rect 1778 237 1779 243
rect 1785 237 1786 243
rect 1778 231 1786 237
rect 1778 225 1779 231
rect 1785 225 1786 231
rect 1778 95 1786 225
rect 1778 89 1779 95
rect 1785 89 1786 95
rect 1778 79 1786 89
rect 1778 73 1779 79
rect 1785 73 1786 79
rect 1778 72 1786 73
rect 1790 3523 1798 3528
rect 1790 3517 1791 3523
rect 1797 3517 1798 3523
rect 1790 3487 1798 3517
rect 1790 3481 1791 3487
rect 1797 3481 1798 3487
rect 1790 3387 1798 3481
rect 1790 3381 1791 3387
rect 1797 3381 1798 3387
rect 1790 3355 1798 3381
rect 1790 3349 1791 3355
rect 1797 3349 1798 3355
rect 1790 3243 1798 3349
rect 1790 3237 1791 3243
rect 1797 3237 1798 3243
rect 1790 3219 1798 3237
rect 1790 3213 1791 3219
rect 1797 3213 1798 3219
rect 1790 3111 1798 3213
rect 1790 3105 1791 3111
rect 1797 3105 1798 3111
rect 1790 3071 1798 3105
rect 1790 3065 1791 3071
rect 1797 3065 1798 3071
rect 1790 2975 1798 3065
rect 1790 2969 1791 2975
rect 1797 2969 1798 2975
rect 1790 2931 1798 2969
rect 1790 2925 1791 2931
rect 1797 2925 1798 2931
rect 1790 2835 1798 2925
rect 1790 2829 1791 2835
rect 1797 2829 1798 2835
rect 1790 2791 1798 2829
rect 1790 2785 1791 2791
rect 1797 2785 1798 2791
rect 1790 2703 1798 2785
rect 1790 2697 1791 2703
rect 1797 2697 1798 2703
rect 1790 2651 1798 2697
rect 1790 2645 1791 2651
rect 1797 2645 1798 2651
rect 1790 2563 1798 2645
rect 1790 2557 1791 2563
rect 1797 2557 1798 2563
rect 1790 2511 1798 2557
rect 1790 2505 1791 2511
rect 1797 2505 1798 2511
rect 1790 2415 1798 2505
rect 1790 2409 1791 2415
rect 1797 2409 1798 2415
rect 1790 2359 1798 2409
rect 1790 2353 1791 2359
rect 1797 2353 1798 2359
rect 1790 2283 1798 2353
rect 1790 2277 1791 2283
rect 1797 2277 1798 2283
rect 1790 2223 1798 2277
rect 1790 2217 1791 2223
rect 1797 2217 1798 2223
rect 1790 2135 1798 2217
rect 1790 2129 1791 2135
rect 1797 2129 1798 2135
rect 1790 2079 1798 2129
rect 1790 2073 1791 2079
rect 1797 2073 1798 2079
rect 1790 1983 1798 2073
rect 1790 1977 1791 1983
rect 1797 1977 1798 1983
rect 1790 1951 1798 1977
rect 1790 1945 1791 1951
rect 1797 1945 1798 1951
rect 1790 1847 1798 1945
rect 1790 1841 1791 1847
rect 1797 1841 1798 1847
rect 1790 1815 1798 1841
rect 1790 1809 1791 1815
rect 1797 1809 1798 1815
rect 1790 1699 1798 1809
rect 1790 1693 1791 1699
rect 1797 1693 1798 1699
rect 1790 1671 1798 1693
rect 1790 1665 1791 1671
rect 1797 1665 1798 1671
rect 1790 1555 1798 1665
rect 1790 1549 1791 1555
rect 1797 1549 1798 1555
rect 1790 1535 1798 1549
rect 1790 1529 1791 1535
rect 1797 1529 1798 1535
rect 1790 1411 1798 1529
rect 1790 1405 1791 1411
rect 1797 1405 1798 1411
rect 1790 1395 1798 1405
rect 1790 1389 1791 1395
rect 1797 1389 1798 1395
rect 1790 1279 1798 1389
rect 1790 1273 1791 1279
rect 1797 1273 1798 1279
rect 1790 1259 1798 1273
rect 1790 1253 1791 1259
rect 1797 1253 1798 1259
rect 1790 1139 1798 1253
rect 1790 1133 1791 1139
rect 1797 1133 1798 1139
rect 1790 1123 1798 1133
rect 1790 1117 1791 1123
rect 1797 1117 1798 1123
rect 1790 1003 1798 1117
rect 1790 997 1791 1003
rect 1797 997 1798 1003
rect 1790 983 1798 997
rect 1790 977 1791 983
rect 1797 977 1798 983
rect 1790 859 1798 977
rect 1790 853 1791 859
rect 1797 853 1798 859
rect 1790 847 1798 853
rect 1790 841 1791 847
rect 1797 841 1798 847
rect 1790 723 1798 841
rect 1790 717 1791 723
rect 1797 717 1798 723
rect 1790 707 1798 717
rect 1790 701 1791 707
rect 1797 701 1798 707
rect 1790 587 1798 701
rect 1790 581 1791 587
rect 1797 581 1798 587
rect 1790 571 1798 581
rect 1790 565 1791 571
rect 1797 565 1798 571
rect 1790 447 1798 565
rect 1790 441 1791 447
rect 1797 441 1798 447
rect 1790 435 1798 441
rect 1790 429 1791 435
rect 1797 429 1798 435
rect 1790 311 1798 429
rect 1790 305 1791 311
rect 1797 305 1798 311
rect 1790 299 1798 305
rect 1790 293 1791 299
rect 1797 293 1798 299
rect 1790 159 1798 293
rect 1790 153 1791 159
rect 1797 153 1798 159
rect 1790 143 1798 153
rect 1790 137 1791 143
rect 1797 137 1798 143
rect 1790 72 1798 137
rect 3486 3459 3494 3528
rect 3486 3453 3487 3459
rect 3493 3453 3494 3459
rect 3486 3315 3494 3453
rect 3486 3309 3487 3315
rect 3493 3309 3494 3315
rect 3486 3179 3494 3309
rect 3486 3173 3487 3179
rect 3493 3173 3494 3179
rect 3486 3039 3494 3173
rect 3486 3033 3487 3039
rect 3493 3033 3494 3039
rect 3486 2903 3494 3033
rect 3486 2897 3487 2903
rect 3493 2897 3494 2903
rect 3486 2767 3494 2897
rect 3486 2761 3487 2767
rect 3493 2761 3494 2767
rect 3486 2635 3494 2761
rect 3486 2629 3487 2635
rect 3493 2629 3494 2635
rect 3486 2483 3494 2629
rect 3486 2477 3487 2483
rect 3493 2477 3494 2483
rect 3486 2351 3494 2477
rect 3486 2345 3487 2351
rect 3493 2345 3494 2351
rect 3486 2207 3494 2345
rect 3486 2201 3487 2207
rect 3493 2201 3494 2207
rect 3486 2063 3494 2201
rect 3486 2057 3487 2063
rect 3493 2057 3494 2063
rect 3486 1915 3494 2057
rect 3486 1909 3487 1915
rect 3493 1909 3494 1915
rect 3486 1771 3494 1909
rect 3486 1765 3487 1771
rect 3493 1765 3494 1771
rect 3486 1627 3494 1765
rect 3486 1621 3487 1627
rect 3493 1621 3494 1627
rect 3486 1483 3494 1621
rect 3486 1477 3487 1483
rect 3493 1477 3494 1483
rect 3486 1343 3494 1477
rect 3486 1337 3487 1343
rect 3493 1337 3494 1343
rect 3486 1215 3494 1337
rect 3486 1209 3487 1215
rect 3493 1209 3494 1215
rect 3486 1067 3494 1209
rect 3486 1061 3487 1067
rect 3493 1061 3494 1067
rect 3486 927 3494 1061
rect 3486 921 3487 927
rect 3493 921 3494 927
rect 3486 791 3494 921
rect 3486 785 3487 791
rect 3493 785 3494 791
rect 3486 659 3494 785
rect 3486 653 3487 659
rect 3493 653 3494 659
rect 3486 519 3494 653
rect 3486 513 3487 519
rect 3493 513 3494 519
rect 3486 379 3494 513
rect 3486 373 3487 379
rect 3493 373 3494 379
rect 3486 243 3494 373
rect 3486 237 3487 243
rect 3493 237 3494 243
rect 3486 95 3494 237
rect 3486 89 3487 95
rect 3493 89 3494 95
rect 3486 72 3494 89
rect 3498 3523 3506 3528
rect 3498 3517 3499 3523
rect 3505 3517 3506 3523
rect 3498 3387 3506 3517
rect 3498 3381 3499 3387
rect 3505 3381 3506 3387
rect 3498 3243 3506 3381
rect 3498 3237 3499 3243
rect 3505 3237 3506 3243
rect 3498 3111 3506 3237
rect 3498 3105 3499 3111
rect 3505 3105 3506 3111
rect 3498 2975 3506 3105
rect 3498 2969 3499 2975
rect 3505 2969 3506 2975
rect 3498 2835 3506 2969
rect 3498 2829 3499 2835
rect 3505 2829 3506 2835
rect 3498 2703 3506 2829
rect 3498 2697 3499 2703
rect 3505 2697 3506 2703
rect 3498 2563 3506 2697
rect 3498 2557 3499 2563
rect 3505 2557 3506 2563
rect 3498 2415 3506 2557
rect 3498 2409 3499 2415
rect 3505 2409 3506 2415
rect 3498 2283 3506 2409
rect 3498 2277 3499 2283
rect 3505 2277 3506 2283
rect 3498 2135 3506 2277
rect 3498 2129 3499 2135
rect 3505 2129 3506 2135
rect 3498 1983 3506 2129
rect 3498 1977 3499 1983
rect 3505 1977 3506 1983
rect 3498 1847 3506 1977
rect 3498 1841 3499 1847
rect 3505 1841 3506 1847
rect 3498 1699 3506 1841
rect 3498 1693 3499 1699
rect 3505 1693 3506 1699
rect 3498 1555 3506 1693
rect 3498 1549 3499 1555
rect 3505 1549 3506 1555
rect 3498 1411 3506 1549
rect 3498 1405 3499 1411
rect 3505 1405 3506 1411
rect 3498 1279 3506 1405
rect 3498 1273 3499 1279
rect 3505 1273 3506 1279
rect 3498 1139 3506 1273
rect 3498 1133 3499 1139
rect 3505 1133 3506 1139
rect 3498 1003 3506 1133
rect 3498 997 3499 1003
rect 3505 997 3506 1003
rect 3498 859 3506 997
rect 3498 853 3499 859
rect 3505 853 3506 859
rect 3498 723 3506 853
rect 3498 717 3499 723
rect 3505 717 3506 723
rect 3498 587 3506 717
rect 3498 581 3499 587
rect 3505 581 3506 587
rect 3498 447 3506 581
rect 3498 441 3499 447
rect 3505 441 3506 447
rect 3498 311 3506 441
rect 3498 305 3499 311
rect 3505 305 3506 311
rect 3498 159 3506 305
rect 3498 153 3499 159
rect 3505 153 3506 159
rect 3498 72 3506 153
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220321
transform 1 0 3456 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220321
transform 1 0 1800 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220321
transform 1 0 3456 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220321
transform 1 0 1800 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220321
transform 1 0 3456 0 1 3340
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220321
transform 1 0 1800 0 1 3340
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220321
transform 1 0 3456 0 -1 3292
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220321
transform 1 0 1800 0 -1 3292
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220321
transform 1 0 3456 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220321
transform 1 0 1800 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220321
transform 1 0 3456 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220321
transform 1 0 1800 0 -1 3156
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220321
transform 1 0 3456 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220321
transform 1 0 1800 0 1 3064
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220321
transform 1 0 3456 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220321
transform 1 0 1800 0 -1 3016
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220321
transform 1 0 3456 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220321
transform 1 0 1800 0 1 2928
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220321
transform 1 0 3456 0 -1 2880
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220321
transform 1 0 1800 0 -1 2880
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220321
transform 1 0 3456 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220321
transform 1 0 1800 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220321
transform 1 0 3456 0 -1 2744
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220321
transform 1 0 1800 0 -1 2744
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220321
transform 1 0 3456 0 1 2656
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220321
transform 1 0 1800 0 1 2656
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220321
transform 1 0 3456 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220321
transform 1 0 1800 0 -1 2612
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220321
transform 1 0 3456 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220321
transform 1 0 1800 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220321
transform 1 0 3456 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220321
transform 1 0 1800 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220321
transform 1 0 3456 0 1 2368
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220321
transform 1 0 1800 0 1 2368
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220321
transform 1 0 3456 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220321
transform 1 0 1800 0 -1 2328
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220321
transform 1 0 3456 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220321
transform 1 0 1800 0 1 2236
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220321
transform 1 0 3456 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220321
transform 1 0 1800 0 -1 2184
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220321
transform 1 0 3456 0 1 2088
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220321
transform 1 0 1800 0 1 2088
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220321
transform 1 0 3456 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220321
transform 1 0 1800 0 -1 2040
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220321
transform 1 0 3456 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220321
transform 1 0 1800 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220321
transform 1 0 3456 0 -1 1892
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220321
transform 1 0 1800 0 -1 1892
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220321
transform 1 0 3456 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220321
transform 1 0 1800 0 1 1800
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220321
transform 1 0 3456 0 -1 1748
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220321
transform 1 0 1800 0 -1 1748
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220321
transform 1 0 3456 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220321
transform 1 0 1800 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220321
transform 1 0 3456 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220321
transform 1 0 1800 0 -1 1604
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220321
transform 1 0 3456 0 1 1508
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220321
transform 1 0 1800 0 1 1508
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220321
transform 1 0 3456 0 -1 1460
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220321
transform 1 0 1800 0 -1 1460
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220321
transform 1 0 3456 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220321
transform 1 0 1800 0 1 1364
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220321
transform 1 0 3456 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220321
transform 1 0 1800 0 -1 1320
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220321
transform 1 0 3456 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220321
transform 1 0 1800 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220321
transform 1 0 3456 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220321
transform 1 0 1800 0 -1 1192
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220321
transform 1 0 3456 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220321
transform 1 0 1800 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220321
transform 1 0 3456 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220321
transform 1 0 1800 0 -1 1044
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220321
transform 1 0 3456 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220321
transform 1 0 1800 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220321
transform 1 0 3456 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220321
transform 1 0 1800 0 -1 904
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220321
transform 1 0 3456 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220321
transform 1 0 1800 0 1 812
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220321
transform 1 0 3456 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220321
transform 1 0 1800 0 -1 768
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220321
transform 1 0 3456 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220321
transform 1 0 1800 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220321
transform 1 0 3456 0 -1 636
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220321
transform 1 0 1800 0 -1 636
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220321
transform 1 0 3456 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220321
transform 1 0 1800 0 1 540
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220321
transform 1 0 3456 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220321
transform 1 0 1800 0 -1 496
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220321
transform 1 0 3456 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220321
transform 1 0 1800 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220321
transform 1 0 3456 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220321
transform 1 0 1800 0 -1 356
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220321
transform 1 0 3456 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220321
transform 1 0 1800 0 1 264
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220321
transform 1 0 3456 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220321
transform 1 0 1800 0 -1 220
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220321
transform 1 0 3456 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220321
transform 1 0 1800 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220321
transform 1 0 1760 0 1 3440
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220321
transform 1 0 104 0 1 3440
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220321
transform 1 0 1760 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220321
transform 1 0 104 0 -1 3400
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220321
transform 1 0 1760 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220321
transform 1 0 104 0 1 3308
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220321
transform 1 0 1760 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220321
transform 1 0 104 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220321
transform 1 0 1760 0 1 3172
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220321
transform 1 0 104 0 1 3172
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220321
transform 1 0 1760 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220321
transform 1 0 104 0 -1 3120
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220321
transform 1 0 1760 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220321
transform 1 0 104 0 1 3024
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220321
transform 1 0 1760 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220321
transform 1 0 104 0 -1 2980
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220321
transform 1 0 1760 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220321
transform 1 0 104 0 1 2884
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220321
transform 1 0 1760 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220321
transform 1 0 104 0 -1 2840
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220321
transform 1 0 1760 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220321
transform 1 0 104 0 1 2744
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220321
transform 1 0 1760 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220321
transform 1 0 104 0 -1 2700
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220321
transform 1 0 1760 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220321
transform 1 0 104 0 1 2604
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220321
transform 1 0 1760 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220321
transform 1 0 104 0 -1 2552
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220321
transform 1 0 1760 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220321
transform 1 0 104 0 1 2464
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220321
transform 1 0 1760 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220321
transform 1 0 104 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220321
transform 1 0 1760 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220321
transform 1 0 104 0 1 2312
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220321
transform 1 0 1760 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220321
transform 1 0 104 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220321
transform 1 0 1760 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220321
transform 1 0 104 0 1 2176
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220321
transform 1 0 1760 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220321
transform 1 0 104 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220321
transform 1 0 1760 0 1 2032
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220321
transform 1 0 104 0 1 2032
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220321
transform 1 0 1760 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220321
transform 1 0 104 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220321
transform 1 0 1760 0 1 1904
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220321
transform 1 0 104 0 1 1904
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220321
transform 1 0 1760 0 -1 1864
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220321
transform 1 0 104 0 -1 1864
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220321
transform 1 0 1760 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220321
transform 1 0 104 0 1 1768
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220321
transform 1 0 1760 0 -1 1716
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220321
transform 1 0 104 0 -1 1716
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220321
transform 1 0 1760 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220321
transform 1 0 104 0 1 1624
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220321
transform 1 0 1760 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220321
transform 1 0 104 0 -1 1580
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220321
transform 1 0 1760 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220321
transform 1 0 104 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220321
transform 1 0 1760 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220321
transform 1 0 104 0 -1 1440
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220321
transform 1 0 1760 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220321
transform 1 0 104 0 1 1348
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220321
transform 1 0 1760 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220321
transform 1 0 104 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220321
transform 1 0 1760 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220321
transform 1 0 104 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220321
transform 1 0 1760 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220321
transform 1 0 104 0 -1 1168
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220321
transform 1 0 1760 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220321
transform 1 0 104 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220321
transform 1 0 1760 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220321
transform 1 0 104 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220321
transform 1 0 1760 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220321
transform 1 0 104 0 1 936
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220321
transform 1 0 1760 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220321
transform 1 0 104 0 -1 892
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220321
transform 1 0 1760 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220321
transform 1 0 104 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220321
transform 1 0 1760 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220321
transform 1 0 104 0 -1 756
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220321
transform 1 0 1760 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220321
transform 1 0 104 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220321
transform 1 0 1760 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220321
transform 1 0 104 0 -1 616
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220321
transform 1 0 1760 0 1 524
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220321
transform 1 0 104 0 1 524
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220321
transform 1 0 1760 0 -1 480
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220321
transform 1 0 104 0 -1 480
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220321
transform 1 0 1760 0 1 388
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220321
transform 1 0 104 0 1 388
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220321
transform 1 0 1760 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220321
transform 1 0 104 0 -1 344
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220321
transform 1 0 1760 0 1 252
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220321
transform 1 0 104 0 1 252
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220321
transform 1 0 1760 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220321
transform 1 0 104 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220321
transform 1 0 1760 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220321
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0cell_0_0gcelem2x0  tst_5999_6
timestamp 1731220321
transform 1 0 3240 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5998_6
timestamp 1731220321
transform 1 0 3040 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5997_6
timestamp 1731220321
transform 1 0 2848 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5996_6
timestamp 1731220321
transform 1 0 2648 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5995_6
timestamp 1731220321
transform 1 0 2968 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5994_6
timestamp 1731220321
transform 1 0 2840 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5993_6
timestamp 1731220321
transform 1 0 2712 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5992_6
timestamp 1731220321
transform 1 0 2592 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5991_6
timestamp 1731220321
transform 1 0 2472 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5990_6
timestamp 1731220321
transform 1 0 2512 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5989_6
timestamp 1731220321
transform 1 0 2640 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5988_6
timestamp 1731220321
transform 1 0 2768 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5987_6
timestamp 1731220321
transform 1 0 3032 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5986_6
timestamp 1731220321
transform 1 0 2896 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5985_6
timestamp 1731220321
transform 1 0 2824 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5984_6
timestamp 1731220321
transform 1 0 2672 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5983_6
timestamp 1731220321
transform 1 0 2968 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5982_6
timestamp 1731220321
transform 1 0 3104 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5981_6
timestamp 1731220321
transform 1 0 3240 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5980_6
timestamp 1731220321
transform 1 0 3360 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5979_6
timestamp 1731220321
transform 1 0 3360 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5978_6
timestamp 1731220321
transform 1 0 3360 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5977_6
timestamp 1731220321
transform 1 0 3256 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5976_6
timestamp 1731220321
transform 1 0 3360 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5975_6
timestamp 1731220321
transform 1 0 3192 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5974_6
timestamp 1731220321
transform 1 0 3128 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5973_6
timestamp 1731220321
transform 1 0 3000 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5972_6
timestamp 1731220321
transform 1 0 3200 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5971_6
timestamp 1731220321
transform 1 0 3016 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5970_6
timestamp 1731220321
transform 1 0 2832 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5969_6
timestamp 1731220321
transform 1 0 2648 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5968_6
timestamp 1731220321
transform 1 0 2568 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5967_6
timestamp 1731220321
transform 1 0 2728 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5966_6
timestamp 1731220321
transform 1 0 2872 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5965_6
timestamp 1731220321
transform 1 0 3024 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5964_6
timestamp 1731220321
transform 1 0 2864 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5963_6
timestamp 1731220321
transform 1 0 2712 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5962_6
timestamp 1731220321
transform 1 0 2560 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5961_6
timestamp 1731220321
transform 1 0 2752 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5960_6
timestamp 1731220321
transform 1 0 2640 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5959_6
timestamp 1731220321
transform 1 0 2536 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5958_6
timestamp 1731220321
transform 1 0 2432 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5957_6
timestamp 1731220321
transform 1 0 2664 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5956_6
timestamp 1731220321
transform 1 0 2576 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5955_6
timestamp 1731220321
transform 1 0 2488 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5954_6
timestamp 1731220321
transform 1 0 2400 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5953_6
timestamp 1731220321
transform 1 0 2224 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5952_6
timestamp 1731220321
transform 1 0 2752 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5951_6
timestamp 1731220321
transform 1 0 2840 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5950_6
timestamp 1731220321
transform 1 0 2776 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5949_6
timestamp 1731220321
transform 1 0 2672 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5948_6
timestamp 1731220321
transform 1 0 2568 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5947_6
timestamp 1731220321
transform 1 0 2464 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5946_6
timestamp 1731220321
transform 1 0 2480 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5945_6
timestamp 1731220321
transform 1 0 2600 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5944_6
timestamp 1731220321
transform 1 0 2712 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5943_6
timestamp 1731220321
transform 1 0 2952 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5942_6
timestamp 1731220321
transform 1 0 2832 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5941_6
timestamp 1731220321
transform 1 0 2760 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5940_6
timestamp 1731220321
transform 1 0 2616 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5939_6
timestamp 1731220321
transform 1 0 2904 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5938_6
timestamp 1731220321
transform 1 0 3048 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5937_6
timestamp 1731220321
transform 1 0 3088 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5936_6
timestamp 1731220321
transform 1 0 2936 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5935_6
timestamp 1731220321
transform 1 0 2776 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5934_6
timestamp 1731220321
transform 1 0 2608 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5933_6
timestamp 1731220321
transform 1 0 2512 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5932_6
timestamp 1731220321
transform 1 0 2664 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5931_6
timestamp 1731220321
transform 1 0 2800 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5930_6
timestamp 1731220321
transform 1 0 2920 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5929_6
timestamp 1731220321
transform 1 0 3040 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5928_6
timestamp 1731220321
transform 1 0 3152 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5927_6
timestamp 1731220321
transform 1 0 3264 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5926_6
timestamp 1731220321
transform 1 0 3232 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5925_6
timestamp 1731220321
transform 1 0 3360 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5924_6
timestamp 1731220321
transform 1 0 3360 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5923_6
timestamp 1731220321
transform 1 0 2792 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5922_6
timestamp 1731220321
transform 1 0 3360 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5921_6
timestamp 1731220321
transform 1 0 3360 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5920_6
timestamp 1731220321
transform 1 0 3360 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5919_6
timestamp 1731220321
transform 1 0 3360 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5918_6
timestamp 1731220321
transform 1 0 3360 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5917_6
timestamp 1731220321
transform 1 0 3360 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5916_6
timestamp 1731220321
transform 1 0 3360 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5915_6
timestamp 1731220321
transform 1 0 3360 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5914_6
timestamp 1731220321
transform 1 0 3360 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5913_6
timestamp 1731220321
transform 1 0 3360 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5912_6
timestamp 1731220321
transform 1 0 3256 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5911_6
timestamp 1731220321
transform 1 0 3128 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5910_6
timestamp 1731220321
transform 1 0 3208 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5909_6
timestamp 1731220321
transform 1 0 3336 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5908_6
timestamp 1731220321
transform 1 0 3312 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5907_6
timestamp 1731220321
transform 1 0 3360 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5906_6
timestamp 1731220321
transform 1 0 3208 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5905_6
timestamp 1731220321
transform 1 0 3248 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5904_6
timestamp 1731220321
transform 1 0 3168 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5903_6
timestamp 1731220321
transform 1 0 3264 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5902_6
timestamp 1731220321
transform 1 0 3152 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5901_6
timestamp 1731220321
transform 1 0 3040 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5900_6
timestamp 1731220321
transform 1 0 2920 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5899_6
timestamp 1731220321
transform 1 0 2800 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5898_6
timestamp 1731220321
transform 1 0 2664 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5897_6
timestamp 1731220321
transform 1 0 2520 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5896_6
timestamp 1731220321
transform 1 0 2552 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5895_6
timestamp 1731220321
transform 1 0 2752 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5894_6
timestamp 1731220321
transform 1 0 2960 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5893_6
timestamp 1731220321
transform 1 0 3040 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5892_6
timestamp 1731220321
transform 1 0 2832 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5891_6
timestamp 1731220321
transform 1 0 2640 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5890_6
timestamp 1731220321
transform 1 0 2456 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5889_6
timestamp 1731220321
transform 1 0 2584 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5888_6
timestamp 1731220321
transform 1 0 2728 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5887_6
timestamp 1731220321
transform 1 0 2880 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5886_6
timestamp 1731220321
transform 1 0 3040 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5885_6
timestamp 1731220321
transform 1 0 2960 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5884_6
timestamp 1731220321
transform 1 0 2832 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5883_6
timestamp 1731220321
transform 1 0 2712 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5882_6
timestamp 1731220321
transform 1 0 3240 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5881_6
timestamp 1731220321
transform 1 0 3096 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5880_6
timestamp 1731220321
transform 1 0 3024 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5879_6
timestamp 1731220321
transform 1 0 2904 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5878_6
timestamp 1731220321
transform 1 0 2776 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5877_6
timestamp 1731220321
transform 1 0 3144 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5876_6
timestamp 1731220321
transform 1 0 3264 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5875_6
timestamp 1731220321
transform 1 0 3256 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5874_6
timestamp 1731220321
transform 1 0 3128 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5873_6
timestamp 1731220321
transform 1 0 3000 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5872_6
timestamp 1731220321
transform 1 0 2864 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5871_6
timestamp 1731220321
transform 1 0 2720 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5870_6
timestamp 1731220321
transform 1 0 3168 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5869_6
timestamp 1731220321
transform 1 0 3024 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5868_6
timestamp 1731220321
transform 1 0 2880 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5867_6
timestamp 1731220321
transform 1 0 2744 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5866_6
timestamp 1731220321
transform 1 0 2608 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5865_6
timestamp 1731220321
transform 1 0 3176 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5864_6
timestamp 1731220321
transform 1 0 2976 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5863_6
timestamp 1731220321
transform 1 0 2784 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5862_6
timestamp 1731220321
transform 1 0 2608 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5861_6
timestamp 1731220321
transform 1 0 3128 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5860_6
timestamp 1731220321
transform 1 0 2928 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5859_6
timestamp 1731220321
transform 1 0 2736 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5858_6
timestamp 1731220321
transform 1 0 2560 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5857_6
timestamp 1731220321
transform 1 0 2400 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5856_6
timestamp 1731220321
transform 1 0 2472 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5855_6
timestamp 1731220321
transform 1 0 2680 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5854_6
timestamp 1731220321
transform 1 0 3144 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5853_6
timestamp 1731220321
transform 1 0 2904 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5852_6
timestamp 1731220321
transform 1 0 2720 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5851_6
timestamp 1731220321
transform 1 0 2568 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5850_6
timestamp 1731220321
transform 1 0 2432 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5849_6
timestamp 1731220321
transform 1 0 2880 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5848_6
timestamp 1731220321
transform 1 0 3040 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5847_6
timestamp 1731220321
transform 1 0 3008 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5846_6
timestamp 1731220321
transform 1 0 2888 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5845_6
timestamp 1731220321
transform 1 0 2760 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5844_6
timestamp 1731220321
transform 1 0 2632 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5843_6
timestamp 1731220321
transform 1 0 2496 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5842_6
timestamp 1731220321
transform 1 0 2592 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5841_6
timestamp 1731220321
transform 1 0 2728 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5840_6
timestamp 1731220321
transform 1 0 2864 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5839_6
timestamp 1731220321
transform 1 0 3000 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5838_6
timestamp 1731220321
transform 1 0 3136 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5837_6
timestamp 1731220321
transform 1 0 3232 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5836_6
timestamp 1731220321
transform 1 0 3080 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5835_6
timestamp 1731220321
transform 1 0 2928 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5834_6
timestamp 1731220321
transform 1 0 2776 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5833_6
timestamp 1731220321
transform 1 0 2880 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5832_6
timestamp 1731220321
transform 1 0 3024 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5831_6
timestamp 1731220321
transform 1 0 3168 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5830_6
timestamp 1731220321
transform 1 0 3320 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5829_6
timestamp 1731220321
transform 1 0 3296 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5828_6
timestamp 1731220321
transform 1 0 3136 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5827_6
timestamp 1731220321
transform 1 0 2984 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5826_6
timestamp 1731220321
transform 1 0 2832 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5825_6
timestamp 1731220321
transform 1 0 3136 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5824_6
timestamp 1731220321
transform 1 0 2968 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5823_6
timestamp 1731220321
transform 1 0 2808 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5822_6
timestamp 1731220321
transform 1 0 2688 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5821_6
timestamp 1731220321
transform 1 0 2840 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5820_6
timestamp 1731220321
transform 1 0 3152 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5819_6
timestamp 1731220321
transform 1 0 2992 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5818_6
timestamp 1731220321
transform 1 0 2864 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5817_6
timestamp 1731220321
transform 1 0 2752 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5816_6
timestamp 1731220321
transform 1 0 2632 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5815_6
timestamp 1731220321
transform 1 0 2968 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5814_6
timestamp 1731220321
transform 1 0 3072 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5813_6
timestamp 1731220321
transform 1 0 3176 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5812_6
timestamp 1731220321
transform 1 0 3272 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5811_6
timestamp 1731220321
transform 1 0 3360 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5810_6
timestamp 1731220321
transform 1 0 3360 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5809_6
timestamp 1731220321
transform 1 0 3360 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5808_6
timestamp 1731220321
transform 1 0 3360 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5807_6
timestamp 1731220321
transform 1 0 3360 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5806_6
timestamp 1731220321
transform 1 0 3360 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5805_6
timestamp 1731220321
transform 1 0 3360 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5804_6
timestamp 1731220321
transform 1 0 3360 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5803_6
timestamp 1731220321
transform 1 0 3360 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5802_6
timestamp 1731220321
transform 1 0 3360 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5801_6
timestamp 1731220321
transform 1 0 3360 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5800_6
timestamp 1731220321
transform 1 0 3360 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5799_6
timestamp 1731220321
transform 1 0 3272 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5798_6
timestamp 1731220321
transform 1 0 3160 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5797_6
timestamp 1731220321
transform 1 0 3200 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5796_6
timestamp 1731220321
transform 1 0 3248 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5795_6
timestamp 1731220321
transform 1 0 3256 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5794_6
timestamp 1731220321
transform 1 0 3256 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5793_6
timestamp 1731220321
transform 1 0 3128 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5792_6
timestamp 1731220321
transform 1 0 3216 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5791_6
timestamp 1731220321
transform 1 0 3048 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5790_6
timestamp 1731220321
transform 1 0 3032 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5789_6
timestamp 1731220321
transform 1 0 2872 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5788_6
timestamp 1731220321
transform 1 0 2680 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5787_6
timestamp 1731220321
transform 1 0 2472 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5786_6
timestamp 1731220321
transform 1 0 2864 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5785_6
timestamp 1731220321
transform 1 0 3192 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5784_6
timestamp 1731220321
transform 1 0 3024 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5783_6
timestamp 1731220321
transform 1 0 3000 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5782_6
timestamp 1731220321
transform 1 0 2872 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5781_6
timestamp 1731220321
transform 1 0 3136 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5780_6
timestamp 1731220321
transform 1 0 3016 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5779_6
timestamp 1731220321
transform 1 0 2904 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5778_6
timestamp 1731220321
transform 1 0 2904 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5777_6
timestamp 1731220321
transform 1 0 3056 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5776_6
timestamp 1731220321
transform 1 0 3216 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5775_6
timestamp 1731220321
transform 1 0 3080 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5774_6
timestamp 1731220321
transform 1 0 2912 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5773_6
timestamp 1731220321
transform 1 0 2752 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5772_6
timestamp 1731220321
transform 1 0 2840 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5771_6
timestamp 1731220321
transform 1 0 3016 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5770_6
timestamp 1731220321
transform 1 0 3048 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5769_6
timestamp 1731220321
transform 1 0 2936 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5768_6
timestamp 1731220321
transform 1 0 2832 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5767_6
timestamp 1731220321
transform 1 0 2728 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5766_6
timestamp 1731220321
transform 1 0 2616 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5765_6
timestamp 1731220321
transform 1 0 2504 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5764_6
timestamp 1731220321
transform 1 0 2392 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5763_6
timestamp 1731220321
transform 1 0 2504 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5762_6
timestamp 1731220321
transform 1 0 2672 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5761_6
timestamp 1731220321
transform 1 0 2592 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5760_6
timestamp 1731220321
transform 1 0 2608 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5759_6
timestamp 1731220321
transform 1 0 2752 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5758_6
timestamp 1731220321
transform 1 0 2792 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5757_6
timestamp 1731220321
transform 1 0 2744 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5756_6
timestamp 1731220321
transform 1 0 2712 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5755_6
timestamp 1731220321
transform 1 0 2560 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5754_6
timestamp 1731220321
transform 1 0 2560 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5753_6
timestamp 1731220321
transform 1 0 2712 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5752_6
timestamp 1731220321
transform 1 0 2872 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5751_6
timestamp 1731220321
transform 1 0 3192 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5750_6
timestamp 1731220321
transform 1 0 3208 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5749_6
timestamp 1731220321
transform 1 0 3032 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5748_6
timestamp 1731220321
transform 1 0 2864 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5747_6
timestamp 1731220321
transform 1 0 2704 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5746_6
timestamp 1731220321
transform 1 0 2552 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5745_6
timestamp 1731220321
transform 1 0 3176 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5744_6
timestamp 1731220321
transform 1 0 2976 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5743_6
timestamp 1731220321
transform 1 0 2784 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5742_6
timestamp 1731220321
transform 1 0 2608 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5741_6
timestamp 1731220321
transform 1 0 2456 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5740_6
timestamp 1731220321
transform 1 0 2320 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5739_6
timestamp 1731220321
transform 1 0 2512 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5738_6
timestamp 1731220321
transform 1 0 2712 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5737_6
timestamp 1731220321
transform 1 0 3152 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5736_6
timestamp 1731220321
transform 1 0 2928 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5735_6
timestamp 1731220321
transform 1 0 2744 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5734_6
timestamp 1731220321
transform 1 0 2616 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5733_6
timestamp 1731220321
transform 1 0 3216 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5732_6
timestamp 1731220321
transform 1 0 3048 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5731_6
timestamp 1731220321
transform 1 0 2888 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5730_6
timestamp 1731220321
transform 1 0 2800 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5729_6
timestamp 1731220321
transform 1 0 2712 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5728_6
timestamp 1731220321
transform 1 0 2624 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5727_6
timestamp 1731220321
transform 1 0 2536 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5726_6
timestamp 1731220321
transform 1 0 2504 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5725_6
timestamp 1731220321
transform 1 0 2536 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5724_6
timestamp 1731220321
transform 1 0 2488 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5723_6
timestamp 1731220321
transform 1 0 2648 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5722_6
timestamp 1731220321
transform 1 0 2680 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5721_6
timestamp 1731220321
transform 1 0 2736 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5720_6
timestamp 1731220321
transform 1 0 2624 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5719_6
timestamp 1731220321
transform 1 0 2448 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5718_6
timestamp 1731220321
transform 1 0 2360 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5717_6
timestamp 1731220321
transform 1 0 2304 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5716_6
timestamp 1731220321
transform 1 0 2296 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5715_6
timestamp 1731220321
transform 1 0 2248 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5714_6
timestamp 1731220321
transform 1 0 2448 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5713_6
timestamp 1731220321
transform 1 0 2464 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5712_6
timestamp 1731220321
transform 1 0 2568 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5711_6
timestamp 1731220321
transform 1 0 2408 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5710_6
timestamp 1731220321
transform 1 0 2240 0 -1 2060
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5709_6
timestamp 1731220321
transform 1 0 2128 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5708_6
timestamp 1731220321
transform 1 0 2248 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5707_6
timestamp 1731220321
transform 1 0 2376 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5706_6
timestamp 1731220321
transform 1 0 2512 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5705_6
timestamp 1731220321
transform 1 0 2648 0 1 2068
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5704_6
timestamp 1731220321
transform 1 0 2600 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5703_6
timestamp 1731220321
transform 1 0 2488 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5702_6
timestamp 1731220321
transform 1 0 2376 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5701_6
timestamp 1731220321
transform 1 0 2272 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5700_6
timestamp 1731220321
transform 1 0 2176 0 -1 2204
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5699_6
timestamp 1731220321
transform 1 0 2456 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5698_6
timestamp 1731220321
transform 1 0 2336 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5697_6
timestamp 1731220321
transform 1 0 2232 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5696_6
timestamp 1731220321
transform 1 0 2128 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5695_6
timestamp 1731220321
transform 1 0 2032 0 1 2216
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5694_6
timestamp 1731220321
transform 1 0 2296 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5693_6
timestamp 1731220321
transform 1 0 2144 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5692_6
timestamp 1731220321
transform 1 0 2008 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5691_6
timestamp 1731220321
transform 1 0 1880 0 -1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5690_6
timestamp 1731220321
transform 1 0 1832 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5689_6
timestamp 1731220321
transform 1 0 2000 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5688_6
timestamp 1731220321
transform 1 0 2176 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5687_6
timestamp 1731220321
transform 1 0 2360 0 1 2348
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5686_6
timestamp 1731220321
transform 1 0 2360 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5685_6
timestamp 1731220321
transform 1 0 2192 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5684_6
timestamp 1731220321
transform 1 0 2008 0 -1 2480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5683_6
timestamp 1731220321
transform 1 0 2200 0 1 2496
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5682_6
timestamp 1731220321
transform 1 0 2352 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5681_6
timestamp 1731220321
transform 1 0 2424 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5680_6
timestamp 1731220321
transform 1 0 2472 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5679_6
timestamp 1731220321
transform 1 0 2328 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5678_6
timestamp 1731220321
transform 1 0 2360 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5677_6
timestamp 1731220321
transform 1 0 2360 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5676_6
timestamp 1731220321
transform 1 0 2312 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5675_6
timestamp 1731220321
transform 1 0 2328 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5674_6
timestamp 1731220321
transform 1 0 2296 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5673_6
timestamp 1731220321
transform 1 0 2424 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5672_6
timestamp 1731220321
transform 1 0 2400 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5671_6
timestamp 1731220321
transform 1 0 2448 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5670_6
timestamp 1731220321
transform 1 0 2240 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5669_6
timestamp 1731220321
transform 1 0 2328 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5668_6
timestamp 1731220321
transform 1 0 2504 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5667_6
timestamp 1731220321
transform 1 0 2376 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5666_6
timestamp 1731220321
transform 1 0 2232 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5665_6
timestamp 1731220321
transform 1 0 2208 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5664_6
timestamp 1731220321
transform 1 0 2344 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5663_6
timestamp 1731220321
transform 1 0 2448 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5662_6
timestamp 1731220321
transform 1 0 2232 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5661_6
timestamp 1731220321
transform 1 0 2000 0 1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5660_6
timestamp 1731220321
transform 1 0 1936 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5659_6
timestamp 1731220321
transform 1 0 1824 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5658_6
timestamp 1731220321
transform 1 0 2072 0 -1 3456
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5657_6
timestamp 1731220321
transform 1 0 2088 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5656_6
timestamp 1731220321
transform 1 0 1944 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5655_6
timestamp 1731220321
transform 1 0 1824 0 1 3320
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5654_6
timestamp 1731220321
transform 1 0 1824 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5653_6
timestamp 1731220321
transform 1 0 1968 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5652_6
timestamp 1731220321
transform 1 0 2144 0 -1 3312
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5651_6
timestamp 1731220321
transform 1 0 2024 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5650_6
timestamp 1731220321
transform 1 0 1824 0 1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5649_6
timestamp 1731220321
transform 1 0 1832 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5648_6
timestamp 1731220321
transform 1 0 2024 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5647_6
timestamp 1731220321
transform 1 0 2216 0 -1 3176
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5646_6
timestamp 1731220321
transform 1 0 2168 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5645_6
timestamp 1731220321
transform 1 0 2048 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5644_6
timestamp 1731220321
transform 1 0 1928 0 1 3044
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5643_6
timestamp 1731220321
transform 1 0 2016 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5642_6
timestamp 1731220321
transform 1 0 2224 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5641_6
timestamp 1731220321
transform 1 0 2120 0 -1 3036
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5640_6
timestamp 1731220321
transform 1 0 2048 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5639_6
timestamp 1731220321
transform 1 0 2136 0 1 2908
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5638_6
timestamp 1731220321
transform 1 0 2264 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5637_6
timestamp 1731220321
transform 1 0 2168 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5636_6
timestamp 1731220321
transform 1 0 2064 0 -1 2900
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5635_6
timestamp 1731220321
transform 1 0 1976 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5634_6
timestamp 1731220321
transform 1 0 2104 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5633_6
timestamp 1731220321
transform 1 0 2232 0 1 2768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5632_6
timestamp 1731220321
transform 1 0 2176 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5631_6
timestamp 1731220321
transform 1 0 2024 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5630_6
timestamp 1731220321
transform 1 0 1880 0 -1 2764
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5629_6
timestamp 1731220321
transform 1 0 1824 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5628_6
timestamp 1731220321
transform 1 0 2016 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5627_6
timestamp 1731220321
transform 1 0 2224 0 1 2636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5626_6
timestamp 1731220321
transform 1 0 2176 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5625_6
timestamp 1731220321
transform 1 0 1992 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5624_6
timestamp 1731220321
transform 1 0 1824 0 -1 2632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5623_6
timestamp 1731220321
transform 1 0 1664 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5622_6
timestamp 1731220321
transform 1 0 1576 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5621_6
timestamp 1731220321
transform 1 0 1488 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5620_6
timestamp 1731220321
transform 1 0 1400 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5619_6
timestamp 1731220321
transform 1 0 1664 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5618_6
timestamp 1731220321
transform 1 0 1568 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5617_6
timestamp 1731220321
transform 1 0 1456 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5616_6
timestamp 1731220321
transform 1 0 1304 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5615_6
timestamp 1731220321
transform 1 0 1208 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5614_6
timestamp 1731220321
transform 1 0 1112 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5613_6
timestamp 1731220321
transform 1 0 1024 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5612_6
timestamp 1731220321
transform 1 0 936 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5611_6
timestamp 1731220321
transform 1 0 848 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5610_6
timestamp 1731220321
transform 1 0 1096 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5609_6
timestamp 1731220321
transform 1 0 1224 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5608_6
timestamp 1731220321
transform 1 0 1344 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5607_6
timestamp 1731220321
transform 1 0 1232 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5606_6
timestamp 1731220321
transform 1 0 1408 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5605_6
timestamp 1731220321
transform 1 0 1584 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5604_6
timestamp 1731220321
transform 1 0 1504 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5603_6
timestamp 1731220321
transform 1 0 1368 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5602_6
timestamp 1731220321
transform 1 0 1232 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5601_6
timestamp 1731220321
transform 1 0 1184 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5600_6
timestamp 1731220321
transform 1 0 1296 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5599_6
timestamp 1731220321
transform 1 0 1408 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5598_6
timestamp 1731220321
transform 1 0 1312 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5597_6
timestamp 1731220321
transform 1 0 1224 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5596_6
timestamp 1731220321
transform 1 0 1136 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5595_6
timestamp 1731220321
transform 1 0 1048 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5594_6
timestamp 1731220321
transform 1 0 960 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5593_6
timestamp 1731220321
transform 1 0 872 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5592_6
timestamp 1731220321
transform 1 0 656 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5591_6
timestamp 1731220321
transform 1 0 568 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5590_6
timestamp 1731220321
transform 1 0 712 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5589_6
timestamp 1731220321
transform 1 0 592 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5588_6
timestamp 1731220321
transform 1 0 472 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5587_6
timestamp 1731220321
transform 1 0 368 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5586_6
timestamp 1731220321
transform 1 0 712 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5585_6
timestamp 1731220321
transform 1 0 544 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5584_6
timestamp 1731220321
transform 1 0 384 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5583_6
timestamp 1731220321
transform 1 0 232 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5582_6
timestamp 1731220321
transform 1 0 128 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5581_6
timestamp 1731220321
transform 1 0 128 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5580_6
timestamp 1731220321
transform 1 0 240 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5579_6
timestamp 1731220321
transform 1 0 688 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5578_6
timestamp 1731220321
transform 1 0 536 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5577_6
timestamp 1731220321
transform 1 0 384 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5576_6
timestamp 1731220321
transform 1 0 304 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5575_6
timestamp 1731220321
transform 1 0 216 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5574_6
timestamp 1731220321
transform 1 0 400 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5573_6
timestamp 1731220321
transform 1 0 584 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5572_6
timestamp 1731220321
transform 1 0 496 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5571_6
timestamp 1731220321
transform 1 0 464 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5570_6
timestamp 1731220321
transform 1 0 552 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5569_6
timestamp 1731220321
transform 1 0 640 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5568_6
timestamp 1731220321
transform 1 0 728 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5567_6
timestamp 1731220321
transform 1 0 816 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5566_6
timestamp 1731220321
transform 1 0 824 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5565_6
timestamp 1731220321
transform 1 0 736 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5564_6
timestamp 1731220321
transform 1 0 648 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5563_6
timestamp 1731220321
transform 1 0 560 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5562_6
timestamp 1731220321
transform 1 0 472 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5561_6
timestamp 1731220321
transform 1 0 736 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5560_6
timestamp 1731220321
transform 1 0 616 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5559_6
timestamp 1731220321
transform 1 0 496 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5558_6
timestamp 1731220321
transform 1 0 384 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5557_6
timestamp 1731220321
transform 1 0 280 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5556_6
timestamp 1731220321
transform 1 0 720 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5555_6
timestamp 1731220321
transform 1 0 560 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5554_6
timestamp 1731220321
transform 1 0 400 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5553_6
timestamp 1731220321
transform 1 0 248 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5552_6
timestamp 1731220321
transform 1 0 128 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5551_6
timestamp 1731220321
transform 1 0 776 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5550_6
timestamp 1731220321
transform 1 0 600 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5549_6
timestamp 1731220321
transform 1 0 424 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5548_6
timestamp 1731220321
transform 1 0 256 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5547_6
timestamp 1731220321
transform 1 0 128 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5546_6
timestamp 1731220321
transform 1 0 128 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5545_6
timestamp 1731220321
transform 1 0 728 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5544_6
timestamp 1731220321
transform 1 0 528 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5543_6
timestamp 1731220321
transform 1 0 320 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5542_6
timestamp 1731220321
transform 1 0 256 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5541_6
timestamp 1731220321
transform 1 0 128 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5540_6
timestamp 1731220321
transform 1 0 784 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5539_6
timestamp 1731220321
transform 1 0 600 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5538_6
timestamp 1731220321
transform 1 0 424 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5537_6
timestamp 1731220321
transform 1 0 312 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5536_6
timestamp 1731220321
transform 1 0 168 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5535_6
timestamp 1731220321
transform 1 0 768 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5534_6
timestamp 1731220321
transform 1 0 616 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5533_6
timestamp 1731220321
transform 1 0 464 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5532_6
timestamp 1731220321
transform 1 0 416 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5531_6
timestamp 1731220321
transform 1 0 296 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5530_6
timestamp 1731220321
transform 1 0 792 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5529_6
timestamp 1731220321
transform 1 0 664 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5528_6
timestamp 1731220321
transform 1 0 536 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5527_6
timestamp 1731220321
transform 1 0 488 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5526_6
timestamp 1731220321
transform 1 0 376 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5525_6
timestamp 1731220321
transform 1 0 600 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5524_6
timestamp 1731220321
transform 1 0 720 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5523_6
timestamp 1731220321
transform 1 0 840 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5522_6
timestamp 1731220321
transform 1 0 800 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5521_6
timestamp 1731220321
transform 1 0 696 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5520_6
timestamp 1731220321
transform 1 0 592 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5519_6
timestamp 1731220321
transform 1 0 488 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5518_6
timestamp 1731220321
transform 1 0 392 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5517_6
timestamp 1731220321
transform 1 0 408 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5516_6
timestamp 1731220321
transform 1 0 496 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5515_6
timestamp 1731220321
transform 1 0 760 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5514_6
timestamp 1731220321
transform 1 0 672 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5513_6
timestamp 1731220321
transform 1 0 584 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5512_6
timestamp 1731220321
transform 1 0 536 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5511_6
timestamp 1731220321
transform 1 0 448 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5510_6
timestamp 1731220321
transform 1 0 624 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5509_6
timestamp 1731220321
transform 1 0 712 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5508_6
timestamp 1731220321
transform 1 0 800 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5507_6
timestamp 1731220321
transform 1 0 888 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5506_6
timestamp 1731220321
transform 1 0 976 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5505_6
timestamp 1731220321
transform 1 0 1152 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5504_6
timestamp 1731220321
transform 1 0 1064 0 1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5503_6
timestamp 1731220321
transform 1 0 1024 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5502_6
timestamp 1731220321
transform 1 0 936 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5501_6
timestamp 1731220321
transform 1 0 848 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5500_6
timestamp 1731220321
transform 1 0 1112 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5499_6
timestamp 1731220321
transform 1 0 1296 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5498_6
timestamp 1731220321
transform 1 0 1200 0 -1 3420
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5497_6
timestamp 1731220321
transform 1 0 1112 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5496_6
timestamp 1731220321
transform 1 0 1008 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5495_6
timestamp 1731220321
transform 1 0 904 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5494_6
timestamp 1731220321
transform 1 0 1216 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5493_6
timestamp 1731220321
transform 1 0 1320 0 1 3288
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5492_6
timestamp 1731220321
transform 1 0 1328 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5491_6
timestamp 1731220321
transform 1 0 1200 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5490_6
timestamp 1731220321
transform 1 0 1080 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5489_6
timestamp 1731220321
transform 1 0 960 0 -1 3284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5488_6
timestamp 1731220321
transform 1 0 920 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5487_6
timestamp 1731220321
transform 1 0 1048 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5486_6
timestamp 1731220321
transform 1 0 1168 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5485_6
timestamp 1731220321
transform 1 0 1424 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5484_6
timestamp 1731220321
transform 1 0 1296 0 1 3152
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5483_6
timestamp 1731220321
transform 1 0 1192 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5482_6
timestamp 1731220321
transform 1 0 1056 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5481_6
timestamp 1731220321
transform 1 0 912 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5480_6
timestamp 1731220321
transform 1 0 1336 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5479_6
timestamp 1731220321
transform 1 0 1480 0 -1 3140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5478_6
timestamp 1731220321
transform 1 0 1504 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5477_6
timestamp 1731220321
transform 1 0 1320 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5476_6
timestamp 1731220321
transform 1 0 1136 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5475_6
timestamp 1731220321
transform 1 0 960 0 1 3004
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5474_6
timestamp 1731220321
transform 1 0 920 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5473_6
timestamp 1731220321
transform 1 0 1096 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5472_6
timestamp 1731220321
transform 1 0 1272 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5471_6
timestamp 1731220321
transform 1 0 1440 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5470_6
timestamp 1731220321
transform 1 0 1616 0 -1 3000
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5469_6
timestamp 1731220321
transform 1 0 1584 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5468_6
timestamp 1731220321
transform 1 0 1424 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5467_6
timestamp 1731220321
transform 1 0 1264 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5466_6
timestamp 1731220321
transform 1 0 1104 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5465_6
timestamp 1731220321
transform 1 0 944 0 1 2864
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5464_6
timestamp 1731220321
transform 1 0 1456 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5463_6
timestamp 1731220321
transform 1 0 1304 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5462_6
timestamp 1731220321
transform 1 0 1160 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5461_6
timestamp 1731220321
transform 1 0 1016 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5460_6
timestamp 1731220321
transform 1 0 872 0 -1 2860
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5459_6
timestamp 1731220321
transform 1 0 1312 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5458_6
timestamp 1731220321
transform 1 0 1192 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5457_6
timestamp 1731220321
transform 1 0 1072 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5456_6
timestamp 1731220321
transform 1 0 960 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5455_6
timestamp 1731220321
transform 1 0 848 0 1 2724
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5454_6
timestamp 1731220321
transform 1 0 1176 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5453_6
timestamp 1731220321
transform 1 0 1088 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5452_6
timestamp 1731220321
transform 1 0 1000 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5451_6
timestamp 1731220321
transform 1 0 912 0 -1 2720
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5450_6
timestamp 1731220321
transform 1 0 1080 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5449_6
timestamp 1731220321
transform 1 0 992 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5448_6
timestamp 1731220321
transform 1 0 904 0 1 2584
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5447_6
timestamp 1731220321
transform 1 0 760 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5446_6
timestamp 1731220321
transform 1 0 672 0 -1 2572
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5445_6
timestamp 1731220321
transform 1 0 832 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5444_6
timestamp 1731220321
transform 1 0 968 0 1 2444
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5443_6
timestamp 1731220321
transform 1 0 1056 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5442_6
timestamp 1731220321
transform 1 0 888 0 -1 2428
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5441_6
timestamp 1731220321
transform 1 0 840 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5440_6
timestamp 1731220321
transform 1 0 968 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5439_6
timestamp 1731220321
transform 1 0 1096 0 1 2292
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5438_6
timestamp 1731220321
transform 1 0 1072 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5437_6
timestamp 1731220321
transform 1 0 960 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5436_6
timestamp 1731220321
transform 1 0 856 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5435_6
timestamp 1731220321
transform 1 0 752 0 -1 2284
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5434_6
timestamp 1731220321
transform 1 0 784 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5433_6
timestamp 1731220321
transform 1 0 696 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5432_6
timestamp 1731220321
transform 1 0 608 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5431_6
timestamp 1731220321
transform 1 0 520 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5430_6
timestamp 1731220321
transform 1 0 432 0 1 2156
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5429_6
timestamp 1731220321
transform 1 0 624 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5428_6
timestamp 1731220321
transform 1 0 512 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5427_6
timestamp 1731220321
transform 1 0 400 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5426_6
timestamp 1731220321
transform 1 0 296 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5425_6
timestamp 1731220321
transform 1 0 248 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5424_6
timestamp 1731220321
transform 1 0 368 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5423_6
timestamp 1731220321
transform 1 0 488 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5422_6
timestamp 1731220321
transform 1 0 480 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5421_6
timestamp 1731220321
transform 1 0 352 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5420_6
timestamp 1731220321
transform 1 0 616 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5419_6
timestamp 1731220321
transform 1 0 704 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5418_6
timestamp 1731220321
transform 1 0 568 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5417_6
timestamp 1731220321
transform 1 0 440 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5416_6
timestamp 1731220321
transform 1 0 552 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5415_6
timestamp 1731220321
transform 1 0 688 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5414_6
timestamp 1731220321
transform 1 0 824 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5413_6
timestamp 1731220321
transform 1 0 840 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5412_6
timestamp 1731220321
transform 1 0 976 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5411_6
timestamp 1731220321
transform 1 0 888 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5410_6
timestamp 1731220321
transform 1 0 752 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5409_6
timestamp 1731220321
transform 1 0 720 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5408_6
timestamp 1731220321
transform 1 0 608 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5407_6
timestamp 1731220321
transform 1 0 736 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5406_6
timestamp 1731220321
transform 1 0 856 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5405_6
timestamp 1731220321
transform 1 0 976 0 -1 2140
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5404_6
timestamp 1731220321
transform 1 0 928 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5403_6
timestamp 1731220321
transform 1 0 824 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5402_6
timestamp 1731220321
transform 1 0 1032 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5401_6
timestamp 1731220321
transform 1 0 1136 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5400_6
timestamp 1731220321
transform 1 0 1248 0 1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5399_6
timestamp 1731220321
transform 1 0 1144 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5398_6
timestamp 1731220321
transform 1 0 1016 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5397_6
timestamp 1731220321
transform 1 0 1264 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5396_6
timestamp 1731220321
transform 1 0 1392 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5395_6
timestamp 1731220321
transform 1 0 1520 0 -1 2012
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5394_6
timestamp 1731220321
transform 1 0 1648 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5393_6
timestamp 1731220321
transform 1 0 1512 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5392_6
timestamp 1731220321
transform 1 0 1376 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5391_6
timestamp 1731220321
transform 1 0 1248 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5390_6
timestamp 1731220321
transform 1 0 1112 0 1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5389_6
timestamp 1731220321
transform 1 0 1448 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5388_6
timestamp 1731220321
transform 1 0 1320 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5387_6
timestamp 1731220321
transform 1 0 1192 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5386_6
timestamp 1731220321
transform 1 0 1072 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5385_6
timestamp 1731220321
transform 1 0 952 0 -1 1884
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5384_6
timestamp 1731220321
transform 1 0 1232 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5383_6
timestamp 1731220321
transform 1 0 1080 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5382_6
timestamp 1731220321
transform 1 0 936 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5381_6
timestamp 1731220321
transform 1 0 928 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5380_6
timestamp 1731220321
transform 1 0 1112 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5379_6
timestamp 1731220321
transform 1 0 1224 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5378_6
timestamp 1731220321
transform 1 0 1032 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5377_6
timestamp 1731220321
transform 1 0 848 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5376_6
timestamp 1731220321
transform 1 0 960 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5375_6
timestamp 1731220321
transform 1 0 1112 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5374_6
timestamp 1731220321
transform 1 0 1192 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5373_6
timestamp 1731220321
transform 1 0 1040 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5372_6
timestamp 1731220321
transform 1 0 888 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5371_6
timestamp 1731220321
transform 1 0 1056 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5370_6
timestamp 1731220321
transform 1 0 920 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5369_6
timestamp 1731220321
transform 1 0 896 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5368_6
timestamp 1731220321
transform 1 0 1024 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5367_6
timestamp 1731220321
transform 1 0 1152 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5366_6
timestamp 1731220321
transform 1 0 1184 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5365_6
timestamp 1731220321
transform 1 0 1304 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5364_6
timestamp 1731220321
transform 1 0 1408 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5363_6
timestamp 1731220321
transform 1 0 1280 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5362_6
timestamp 1731220321
transform 1 0 1192 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5361_6
timestamp 1731220321
transform 1 0 1328 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5360_6
timestamp 1731220321
transform 1 0 1464 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5359_6
timestamp 1731220321
transform 1 0 1496 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5358_6
timestamp 1731220321
transform 1 0 1344 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5357_6
timestamp 1731220321
transform 1 0 1272 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5356_6
timestamp 1731220321
transform 1 0 1600 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5355_6
timestamp 1731220321
transform 1 0 1432 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5354_6
timestamp 1731220321
transform 1 0 1424 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5353_6
timestamp 1731220321
transform 1 0 1632 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5352_6
timestamp 1731220321
transform 1 0 1664 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5351_6
timestamp 1731220321
transform 1 0 1496 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5350_6
timestamp 1731220321
transform 1 0 1304 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5349_6
timestamp 1731220321
transform 1 0 1384 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5348_6
timestamp 1731220321
transform 1 0 1536 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5347_6
timestamp 1731220321
transform 1 0 1664 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5346_6
timestamp 1731220321
transform 1 0 1824 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5345_6
timestamp 1731220321
transform 1 0 1824 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5344_6
timestamp 1731220321
transform 1 0 1912 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5343_6
timestamp 1731220321
transform 1 0 1824 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5342_6
timestamp 1731220321
transform 1 0 1912 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5341_6
timestamp 1731220321
transform 1 0 2040 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5340_6
timestamp 1731220321
transform 1 0 2176 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5339_6
timestamp 1731220321
transform 1 0 2320 0 1 1916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5338_6
timestamp 1731220321
transform 1 0 2296 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5337_6
timestamp 1731220321
transform 1 0 2160 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5336_6
timestamp 1731220321
transform 1 0 2032 0 -1 1912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5335_6
timestamp 1731220321
transform 1 0 2104 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5334_6
timestamp 1731220321
transform 1 0 1952 0 1 1780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5333_6
timestamp 1731220321
transform 1 0 1872 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5332_6
timestamp 1731220321
transform 1 0 2008 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5331_6
timestamp 1731220321
transform 1 0 2144 0 -1 1768
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5330_6
timestamp 1731220321
transform 1 0 2176 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5329_6
timestamp 1731220321
transform 1 0 2056 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5328_6
timestamp 1731220321
transform 1 0 1928 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5327_6
timestamp 1731220321
transform 1 0 1824 0 1 1632
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5326_6
timestamp 1731220321
transform 1 0 1824 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5325_6
timestamp 1731220321
transform 1 0 1936 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5324_6
timestamp 1731220321
transform 1 0 2080 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5323_6
timestamp 1731220321
transform 1 0 2224 0 -1 1624
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5322_6
timestamp 1731220321
transform 1 0 2296 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5321_6
timestamp 1731220321
transform 1 0 2144 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5320_6
timestamp 1731220321
transform 1 0 1984 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5319_6
timestamp 1731220321
transform 1 0 1832 0 1 1488
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5318_6
timestamp 1731220321
transform 1 0 1936 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5317_6
timestamp 1731220321
transform 1 0 2048 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5316_6
timestamp 1731220321
transform 1 0 2184 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5315_6
timestamp 1731220321
transform 1 0 2472 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5314_6
timestamp 1731220321
transform 1 0 2328 0 -1 1480
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5313_6
timestamp 1731220321
transform 1 0 2312 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5312_6
timestamp 1731220321
transform 1 0 2192 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5311_6
timestamp 1731220321
transform 1 0 2088 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5310_6
timestamp 1731220321
transform 1 0 2448 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5309_6
timestamp 1731220321
transform 1 0 2592 0 1 1344
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5308_6
timestamp 1731220321
transform 1 0 2528 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5307_6
timestamp 1731220321
transform 1 0 2376 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5306_6
timestamp 1731220321
transform 1 0 2232 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5305_6
timestamp 1731220321
transform 1 0 2096 0 -1 1340
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5304_6
timestamp 1731220321
transform 1 0 2336 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5303_6
timestamp 1731220321
transform 1 0 2192 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5302_6
timestamp 1731220321
transform 1 0 2056 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5301_6
timestamp 1731220321
transform 1 0 1928 0 1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5300_6
timestamp 1731220321
transform 1 0 2384 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5299_6
timestamp 1731220321
transform 1 0 2224 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5298_6
timestamp 1731220321
transform 1 0 2072 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5297_6
timestamp 1731220321
transform 1 0 1928 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5296_6
timestamp 1731220321
transform 1 0 1824 0 -1 1212
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5295_6
timestamp 1731220321
transform 1 0 1856 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5294_6
timestamp 1731220321
transform 1 0 1976 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5293_6
timestamp 1731220321
transform 1 0 2104 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5292_6
timestamp 1731220321
transform 1 0 2240 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5291_6
timestamp 1731220321
transform 1 0 2376 0 1 1072
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5290_6
timestamp 1731220321
transform 1 0 2272 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5289_6
timestamp 1731220321
transform 1 0 2184 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5288_6
timestamp 1731220321
transform 1 0 2096 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5287_6
timestamp 1731220321
transform 1 0 2360 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5286_6
timestamp 1731220321
transform 1 0 2448 0 -1 1064
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5285_6
timestamp 1731220321
transform 1 0 2504 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5284_6
timestamp 1731220321
transform 1 0 2400 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5283_6
timestamp 1731220321
transform 1 0 2304 0 1 936
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5282_6
timestamp 1731220321
transform 1 0 2144 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5281_6
timestamp 1731220321
transform 1 0 1976 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5280_6
timestamp 1731220321
transform 1 0 2080 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5279_6
timestamp 1731220321
transform 1 0 2320 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5278_6
timestamp 1731220321
transform 1 0 2200 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5277_6
timestamp 1731220321
transform 1 0 2144 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5276_6
timestamp 1731220321
transform 1 0 2280 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5275_6
timestamp 1731220321
transform 1 0 2416 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5274_6
timestamp 1731220321
transform 1 0 2408 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5273_6
timestamp 1731220321
transform 1 0 2256 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5272_6
timestamp 1731220321
transform 1 0 2096 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5271_6
timestamp 1731220321
transform 1 0 2232 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5270_6
timestamp 1731220321
transform 1 0 1968 0 -1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5269_6
timestamp 1731220321
transform 1 0 1888 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5268_6
timestamp 1731220321
transform 1 0 2008 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5267_6
timestamp 1731220321
transform 1 0 2136 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5266_6
timestamp 1731220321
transform 1 0 2272 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5265_6
timestamp 1731220321
transform 1 0 2416 0 1 520
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5264_6
timestamp 1731220321
transform 1 0 2352 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5263_6
timestamp 1731220321
transform 1 0 2232 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5262_6
timestamp 1731220321
transform 1 0 2128 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5261_6
timestamp 1731220321
transform 1 0 2480 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5260_6
timestamp 1731220321
transform 1 0 2608 0 -1 516
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5259_6
timestamp 1731220321
transform 1 0 2672 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5258_6
timestamp 1731220321
transform 1 0 2552 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5257_6
timestamp 1731220321
transform 1 0 2440 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5256_6
timestamp 1731220321
transform 1 0 2328 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5255_6
timestamp 1731220321
transform 1 0 2232 0 1 380
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5254_6
timestamp 1731220321
transform 1 0 2472 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5253_6
timestamp 1731220321
transform 1 0 2352 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5252_6
timestamp 1731220321
transform 1 0 2240 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5251_6
timestamp 1731220321
transform 1 0 2144 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5250_6
timestamp 1731220321
transform 1 0 2056 0 -1 376
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5249_6
timestamp 1731220321
transform 1 0 2440 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5248_6
timestamp 1731220321
transform 1 0 2296 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5247_6
timestamp 1731220321
transform 1 0 2160 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5246_6
timestamp 1731220321
transform 1 0 2032 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5245_6
timestamp 1731220321
transform 1 0 1920 0 1 244
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5244_6
timestamp 1731220321
transform 1 0 2344 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5243_6
timestamp 1731220321
transform 1 0 2192 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5242_6
timestamp 1731220321
transform 1 0 2048 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5241_6
timestamp 1731220321
transform 1 0 1920 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5240_6
timestamp 1731220321
transform 1 0 1824 0 -1 240
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5239_6
timestamp 1731220321
transform 1 0 2272 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5238_6
timestamp 1731220321
transform 1 0 2152 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5237_6
timestamp 1731220321
transform 1 0 2032 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5236_6
timestamp 1731220321
transform 1 0 1912 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5235_6
timestamp 1731220321
transform 1 0 1824 0 1 92
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5234_6
timestamp 1731220321
transform 1 0 1664 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5233_6
timestamp 1731220321
transform 1 0 1576 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5232_6
timestamp 1731220321
transform 1 0 1488 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5231_6
timestamp 1731220321
transform 1 0 1400 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5230_6
timestamp 1731220321
transform 1 0 1304 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5229_6
timestamp 1731220321
transform 1 0 1208 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5228_6
timestamp 1731220321
transform 1 0 1112 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5227_6
timestamp 1731220321
transform 1 0 1024 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5226_6
timestamp 1731220321
transform 1 0 936 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5225_6
timestamp 1731220321
transform 1 0 840 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5224_6
timestamp 1731220321
transform 1 0 1424 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5223_6
timestamp 1731220321
transform 1 0 1272 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5222_6
timestamp 1731220321
transform 1 0 1128 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5221_6
timestamp 1731220321
transform 1 0 984 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5220_6
timestamp 1731220321
transform 1 0 832 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5219_6
timestamp 1731220321
transform 1 0 1144 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5218_6
timestamp 1731220321
transform 1 0 1040 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5217_6
timestamp 1731220321
transform 1 0 936 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5216_6
timestamp 1731220321
transform 1 0 840 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5215_6
timestamp 1731220321
transform 1 0 744 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5214_6
timestamp 1731220321
transform 1 0 904 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5213_6
timestamp 1731220321
transform 1 0 992 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5212_6
timestamp 1731220321
transform 1 0 1080 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5211_6
timestamp 1731220321
transform 1 0 1256 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5210_6
timestamp 1731220321
transform 1 0 1168 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5209_6
timestamp 1731220321
transform 1 0 1120 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5208_6
timestamp 1731220321
transform 1 0 1016 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5207_6
timestamp 1731220321
transform 1 0 1224 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5206_6
timestamp 1731220321
transform 1 0 1432 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5205_6
timestamp 1731220321
transform 1 0 1328 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5204_6
timestamp 1731220321
transform 1 0 1216 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5203_6
timestamp 1731220321
transform 1 0 1056 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5202_6
timestamp 1731220321
transform 1 0 1368 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5201_6
timestamp 1731220321
transform 1 0 1520 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5200_6
timestamp 1731220321
transform 1 0 1664 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5199_6
timestamp 1731220321
transform 1 0 1664 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5198_6
timestamp 1731220321
transform 1 0 1496 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5197_6
timestamp 1731220321
transform 1 0 1312 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5196_6
timestamp 1731220321
transform 1 0 1520 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5195_6
timestamp 1731220321
transform 1 0 1664 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5194_6
timestamp 1731220321
transform 1 0 1664 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5193_6
timestamp 1731220321
transform 1 0 1824 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5192_6
timestamp 1731220321
transform 1 0 1944 0 1 656
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5191_6
timestamp 1731220321
transform 1 0 1872 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5190_6
timestamp 1731220321
transform 1 0 2008 0 -1 788
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5189_6
timestamp 1731220321
transform 1 0 1952 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5188_6
timestamp 1731220321
transform 1 0 1824 0 1 792
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5187_6
timestamp 1731220321
transform 1 0 1824 0 -1 924
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5186_6
timestamp 1731220321
transform 1 0 1664 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5185_6
timestamp 1731220321
transform 1 0 1576 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5184_6
timestamp 1731220321
transform 1 0 1480 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5183_6
timestamp 1731220321
transform 1 0 1664 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5182_6
timestamp 1731220321
transform 1 0 1528 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5181_6
timestamp 1731220321
transform 1 0 1376 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5180_6
timestamp 1731220321
transform 1 0 1384 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5179_6
timestamp 1731220321
transform 1 0 1288 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5178_6
timestamp 1731220321
transform 1 0 1192 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5177_6
timestamp 1731220321
transform 1 0 1088 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5176_6
timestamp 1731220321
transform 1 0 1336 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5175_6
timestamp 1731220321
transform 1 0 1456 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5174_6
timestamp 1731220321
transform 1 0 1576 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5173_6
timestamp 1731220321
transform 1 0 1552 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5172_6
timestamp 1731220321
transform 1 0 1424 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5171_6
timestamp 1731220321
transform 1 0 1304 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5170_6
timestamp 1731220321
transform 1 0 1184 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5169_6
timestamp 1731220321
transform 1 0 1152 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5168_6
timestamp 1731220321
transform 1 0 1280 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5167_6
timestamp 1731220321
transform 1 0 1408 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5166_6
timestamp 1731220321
transform 1 0 1504 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5165_6
timestamp 1731220321
transform 1 0 1320 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5164_6
timestamp 1731220321
transform 1 0 1144 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5163_6
timestamp 1731220321
transform 1 0 1360 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5162_6
timestamp 1731220321
transform 1 0 1200 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5161_6
timestamp 1731220321
transform 1 0 1048 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5160_6
timestamp 1731220321
transform 1 0 1128 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5159_6
timestamp 1731220321
transform 1 0 944 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5158_6
timestamp 1731220321
transform 1 0 904 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5157_6
timestamp 1731220321
transform 1 0 760 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5156_6
timestamp 1731220321
transform 1 0 824 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5155_6
timestamp 1731220321
transform 1 0 976 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5154_6
timestamp 1731220321
transform 1 0 904 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5153_6
timestamp 1731220321
transform 1 0 1024 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5152_6
timestamp 1731220321
transform 1 0 1064 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5151_6
timestamp 1731220321
transform 1 0 1216 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5150_6
timestamp 1731220321
transform 1 0 1104 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5149_6
timestamp 1731220321
transform 1 0 984 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5148_6
timestamp 1731220321
transform 1 0 1072 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5147_6
timestamp 1731220321
transform 1 0 1224 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5146_6
timestamp 1731220321
transform 1 0 1552 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5145_6
timestamp 1731220321
transform 1 0 1400 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5144_6
timestamp 1731220321
transform 1 0 1256 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5143_6
timestamp 1731220321
transform 1 0 1112 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5142_6
timestamp 1731220321
transform 1 0 960 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5141_6
timestamp 1731220321
transform 1 0 1328 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5140_6
timestamp 1731220321
transform 1 0 1192 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5139_6
timestamp 1731220321
transform 1 0 1056 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5138_6
timestamp 1731220321
transform 1 0 920 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5137_6
timestamp 1731220321
transform 1 0 784 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5136_6
timestamp 1731220321
transform 1 0 1184 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5135_6
timestamp 1731220321
transform 1 0 1064 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5134_6
timestamp 1731220321
transform 1 0 952 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5133_6
timestamp 1731220321
transform 1 0 840 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5132_6
timestamp 1731220321
transform 1 0 728 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5131_6
timestamp 1731220321
transform 1 0 1072 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5130_6
timestamp 1731220321
transform 1 0 960 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5129_6
timestamp 1731220321
transform 1 0 840 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5128_6
timestamp 1731220321
transform 1 0 712 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5127_6
timestamp 1731220321
transform 1 0 608 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5126_6
timestamp 1731220321
transform 1 0 576 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5125_6
timestamp 1731220321
transform 1 0 432 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5124_6
timestamp 1731220321
transform 1 0 272 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5123_6
timestamp 1731220321
transform 1 0 600 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5122_6
timestamp 1731220321
transform 1 0 752 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5121_6
timestamp 1731220321
transform 1 0 776 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5120_6
timestamp 1731220321
transform 1 0 624 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5119_6
timestamp 1731220321
transform 1 0 464 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5118_6
timestamp 1731220321
transform 1 0 600 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5117_6
timestamp 1731220321
transform 1 0 744 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5116_6
timestamp 1731220321
transform 1 0 808 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5115_6
timestamp 1731220321
transform 1 0 664 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5114_6
timestamp 1731220321
transform 1 0 536 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5113_6
timestamp 1731220321
transform 1 0 528 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5112_6
timestamp 1731220321
transform 1 0 680 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5111_6
timestamp 1731220321
transform 1 0 560 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5110_6
timestamp 1731220321
transform 1 0 744 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5109_6
timestamp 1731220321
transform 1 0 792 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5108_6
timestamp 1731220321
transform 1 0 648 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5107_6
timestamp 1731220321
transform 1 0 520 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5106_6
timestamp 1731220321
transform 1 0 400 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5105_6
timestamp 1731220321
transform 1 0 304 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5104_6
timestamp 1731220321
transform 1 0 216 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5103_6
timestamp 1731220321
transform 1 0 128 0 1 1748
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5102_6
timestamp 1731220321
transform 1 0 128 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5101_6
timestamp 1731220321
transform 1 0 240 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_5100_6
timestamp 1731220321
transform 1 0 392 0 -1 1736
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_599_6
timestamp 1731220321
transform 1 0 400 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_598_6
timestamp 1731220321
transform 1 0 288 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_597_6
timestamp 1731220321
transform 1 0 184 0 1 1604
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_596_6
timestamp 1731220321
transform 1 0 320 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_595_6
timestamp 1731220321
transform 1 0 424 0 -1 1600
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_594_6
timestamp 1731220321
transform 1 0 464 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_593_6
timestamp 1731220321
transform 1 0 336 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_592_6
timestamp 1731220321
transform 1 0 216 0 1 1468
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_591_6
timestamp 1731220321
transform 1 0 128 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_590_6
timestamp 1731220321
transform 1 0 296 0 -1 1460
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_589_6
timestamp 1731220321
transform 1 0 440 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_588_6
timestamp 1731220321
transform 1 0 272 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_587_6
timestamp 1731220321
transform 1 0 128 0 1 1328
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_586_6
timestamp 1731220321
transform 1 0 128 0 -1 1324
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_585_6
timestamp 1731220321
transform 1 0 128 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_584_6
timestamp 1731220321
transform 1 0 232 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_583_6
timestamp 1731220321
transform 1 0 360 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_582_6
timestamp 1731220321
transform 1 0 488 0 1 1192
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_581_6
timestamp 1731220321
transform 1 0 648 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_580_6
timestamp 1731220321
transform 1 0 504 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_579_6
timestamp 1731220321
transform 1 0 368 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_578_6
timestamp 1731220321
transform 1 0 232 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_577_6
timestamp 1731220321
transform 1 0 128 0 -1 1188
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_576_6
timestamp 1731220321
transform 1 0 184 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_575_6
timestamp 1731220321
transform 1 0 328 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_574_6
timestamp 1731220321
transform 1 0 488 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_573_6
timestamp 1731220321
transform 1 0 808 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_572_6
timestamp 1731220321
transform 1 0 648 0 1 1056
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_571_6
timestamp 1731220321
transform 1 0 600 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_570_6
timestamp 1731220321
transform 1 0 456 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_569_6
timestamp 1731220321
transform 1 0 320 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_568_6
timestamp 1731220321
transform 1 0 760 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_567_6
timestamp 1731220321
transform 1 0 920 0 -1 1048
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_566_6
timestamp 1731220321
transform 1 0 880 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_565_6
timestamp 1731220321
transform 1 0 776 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_564_6
timestamp 1731220321
transform 1 0 664 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_563_6
timestamp 1731220321
transform 1 0 560 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_562_6
timestamp 1731220321
transform 1 0 464 0 1 916
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_561_6
timestamp 1731220321
transform 1 0 600 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_560_6
timestamp 1731220321
transform 1 0 688 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_559_6
timestamp 1731220321
transform 1 0 784 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_558_6
timestamp 1731220321
transform 1 0 888 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_557_6
timestamp 1731220321
transform 1 0 992 0 -1 912
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_556_6
timestamp 1731220321
transform 1 0 944 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_555_6
timestamp 1731220321
transform 1 0 824 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_554_6
timestamp 1731220321
transform 1 0 712 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_553_6
timestamp 1731220321
transform 1 0 608 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_552_6
timestamp 1731220321
transform 1 0 512 0 1 780
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_551_6
timestamp 1731220321
transform 1 0 784 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_550_6
timestamp 1731220321
transform 1 0 672 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_549_6
timestamp 1731220321
transform 1 0 568 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_548_6
timestamp 1731220321
transform 1 0 464 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_547_6
timestamp 1731220321
transform 1 0 376 0 -1 776
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_546_6
timestamp 1731220321
transform 1 0 688 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_545_6
timestamp 1731220321
transform 1 0 560 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_544_6
timestamp 1731220321
transform 1 0 448 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_543_6
timestamp 1731220321
transform 1 0 336 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_542_6
timestamp 1731220321
transform 1 0 240 0 1 640
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_541_6
timestamp 1731220321
transform 1 0 616 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_540_6
timestamp 1731220321
transform 1 0 480 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_539_6
timestamp 1731220321
transform 1 0 352 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_538_6
timestamp 1731220321
transform 1 0 224 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_537_6
timestamp 1731220321
transform 1 0 128 0 -1 636
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_536_6
timestamp 1731220321
transform 1 0 128 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_535_6
timestamp 1731220321
transform 1 0 240 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_534_6
timestamp 1731220321
transform 1 0 400 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_533_6
timestamp 1731220321
transform 1 0 760 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_532_6
timestamp 1731220321
transform 1 0 576 0 1 504
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_531_6
timestamp 1731220321
transform 1 0 560 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_530_6
timestamp 1731220321
transform 1 0 392 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_529_6
timestamp 1731220321
transform 1 0 240 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_528_6
timestamp 1731220321
transform 1 0 728 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_527_6
timestamp 1731220321
transform 1 0 896 0 -1 500
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_526_6
timestamp 1731220321
transform 1 0 920 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_525_6
timestamp 1731220321
transform 1 0 712 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_524_6
timestamp 1731220321
transform 1 0 608 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_523_6
timestamp 1731220321
transform 1 0 512 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_522_6
timestamp 1731220321
transform 1 0 816 0 1 368
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_521_6
timestamp 1731220321
transform 1 0 816 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_520_6
timestamp 1731220321
transform 1 0 728 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_519_6
timestamp 1731220321
transform 1 0 640 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_518_6
timestamp 1731220321
transform 1 0 552 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_517_6
timestamp 1731220321
transform 1 0 464 0 -1 364
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_516_6
timestamp 1731220321
transform 1 0 648 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_515_6
timestamp 1731220321
transform 1 0 552 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_514_6
timestamp 1731220321
transform 1 0 456 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_513_6
timestamp 1731220321
transform 1 0 360 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_512_6
timestamp 1731220321
transform 1 0 272 0 1 232
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_511_6
timestamp 1731220321
transform 1 0 672 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_510_6
timestamp 1731220321
transform 1 0 504 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_59_6
timestamp 1731220321
transform 1 0 336 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_58_6
timestamp 1731220321
transform 1 0 160 0 -1 228
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_57_6
timestamp 1731220321
transform 1 0 744 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_56_6
timestamp 1731220321
transform 1 0 656 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_55_6
timestamp 1731220321
transform 1 0 568 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_54_6
timestamp 1731220321
transform 1 0 480 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_53_6
timestamp 1731220321
transform 1 0 392 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_52_6
timestamp 1731220321
transform 1 0 304 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_51_6
timestamp 1731220321
transform 1 0 216 0 1 76
box 8 4 84 60
use _0_0cell_0_0gcelem2x0  tst_50_6
timestamp 1731220321
transform 1 0 128 0 1 76
box 8 4 84 60
<< end >>
