magic
tech sky130l
timestamp 1730768378
<< m1 >>
rect 1424 1501 1428 1535
rect 1568 1347 1572 1499
rect 1000 631 1004 663
rect 296 471 300 503
<< m2c >>
rect 241 1725 245 1729
rect 377 1725 381 1729
rect 513 1725 517 1729
rect 649 1725 653 1729
rect 784 1725 788 1729
rect 111 1721 115 1725
rect 1719 1721 1723 1725
rect 111 1703 115 1707
rect 1719 1703 1723 1707
rect 111 1629 115 1633
rect 1719 1629 1723 1633
rect 111 1611 115 1615
rect 1719 1611 1723 1615
rect 328 1607 332 1611
rect 464 1607 468 1611
rect 600 1607 604 1611
rect 736 1607 740 1611
rect 872 1607 876 1611
rect 1424 1535 1428 1539
rect 593 1497 597 1501
rect 729 1497 733 1501
rect 865 1497 869 1501
rect 1001 1497 1005 1501
rect 1136 1497 1140 1501
rect 1273 1497 1277 1501
rect 1409 1497 1413 1501
rect 1424 1497 1428 1501
rect 1545 1497 1549 1501
rect 1568 1499 1572 1503
rect 111 1493 115 1497
rect 111 1475 115 1479
rect 111 1401 115 1405
rect 111 1383 115 1387
rect 824 1379 828 1383
rect 968 1379 972 1383
rect 1112 1379 1116 1383
rect 1256 1379 1260 1383
rect 1400 1379 1404 1383
rect 1544 1379 1548 1383
rect 1680 1497 1684 1501
rect 1719 1493 1723 1497
rect 1719 1475 1723 1479
rect 1719 1401 1723 1405
rect 1719 1383 1723 1387
rect 1680 1379 1684 1383
rect 1568 1343 1572 1347
rect 288 1273 292 1277
rect 520 1273 524 1277
rect 784 1273 788 1277
rect 1080 1273 1084 1277
rect 1392 1273 1396 1277
rect 1680 1273 1684 1277
rect 111 1269 115 1273
rect 1719 1269 1723 1273
rect 111 1251 115 1255
rect 1719 1251 1723 1255
rect 111 1189 115 1193
rect 1719 1189 1723 1193
rect 111 1171 115 1175
rect 1719 1171 1723 1175
rect 240 1167 244 1171
rect 416 1167 420 1171
rect 640 1167 644 1171
rect 880 1167 884 1171
rect 1144 1167 1148 1171
rect 1416 1167 1420 1171
rect 1680 1167 1684 1171
rect 329 1053 333 1057
rect 569 1053 573 1057
rect 825 1053 829 1057
rect 1096 1053 1100 1057
rect 1376 1053 1380 1057
rect 1664 1053 1668 1057
rect 111 1049 115 1053
rect 1719 1049 1723 1053
rect 111 1031 115 1035
rect 1719 1031 1723 1035
rect 111 973 115 977
rect 1719 973 1723 977
rect 111 955 115 959
rect 1719 955 1723 959
rect 544 951 548 955
rect 728 951 732 955
rect 936 951 940 955
rect 1160 951 1164 955
rect 1392 951 1396 955
rect 1624 951 1628 955
rect 793 845 797 849
rect 929 845 933 849
rect 1065 845 1069 849
rect 1201 845 1205 849
rect 1336 845 1340 849
rect 1472 845 1476 849
rect 1608 845 1612 849
rect 111 841 115 845
rect 1719 841 1723 845
rect 111 823 115 827
rect 1719 823 1723 827
rect 111 753 115 757
rect 1719 753 1723 757
rect 111 735 115 739
rect 1719 735 1723 739
rect 896 731 900 735
rect 1032 731 1036 735
rect 1168 731 1172 735
rect 1304 731 1308 735
rect 1440 731 1444 735
rect 1576 731 1580 735
rect 1000 663 1004 667
rect 617 625 621 629
rect 784 625 788 629
rect 960 625 964 629
rect 1000 627 1004 631
rect 1136 625 1140 629
rect 1321 625 1325 629
rect 1512 625 1516 629
rect 111 621 115 625
rect 1719 621 1723 625
rect 111 603 115 607
rect 1719 603 1723 607
rect 111 525 115 529
rect 1719 525 1723 529
rect 111 507 115 511
rect 1719 507 1723 511
rect 248 503 252 507
rect 296 503 300 507
rect 440 503 444 507
rect 632 503 636 507
rect 824 503 828 507
rect 1016 503 1020 507
rect 1208 503 1212 507
rect 1408 503 1412 507
rect 1608 503 1612 507
rect 296 467 300 471
rect 241 381 245 385
rect 457 381 461 385
rect 721 381 725 385
rect 1000 381 1004 385
rect 1288 381 1292 385
rect 1576 381 1580 385
rect 111 377 115 381
rect 1719 377 1723 381
rect 111 359 115 363
rect 1719 359 1723 363
rect 111 293 115 297
rect 1719 293 1723 297
rect 111 275 115 279
rect 1719 275 1723 279
rect 304 271 308 275
rect 536 271 540 275
rect 768 271 772 275
rect 1000 271 1004 275
rect 1232 271 1236 275
rect 1464 271 1468 275
rect 1680 271 1684 275
rect 417 153 421 157
rect 553 153 557 157
rect 697 153 701 157
rect 849 153 853 157
rect 1009 153 1013 157
rect 1177 153 1181 157
rect 1344 153 1348 157
rect 1680 153 1684 157
rect 111 149 115 153
rect 1719 149 1723 153
rect 111 131 115 135
rect 1719 131 1723 135
<< m2 >>
rect 242 1767 248 1768
rect 242 1763 243 1767
rect 247 1766 248 1767
rect 378 1767 384 1768
rect 247 1764 285 1766
rect 247 1763 248 1764
rect 242 1762 248 1763
rect 378 1763 379 1767
rect 383 1766 384 1767
rect 514 1767 520 1768
rect 383 1764 421 1766
rect 383 1763 384 1764
rect 378 1762 384 1763
rect 514 1763 515 1767
rect 519 1766 520 1767
rect 650 1767 656 1768
rect 519 1764 557 1766
rect 519 1763 520 1764
rect 514 1762 520 1763
rect 650 1763 651 1767
rect 655 1766 656 1767
rect 655 1764 693 1766
rect 655 1763 656 1764
rect 650 1762 656 1763
rect 240 1729 248 1730
rect 110 1725 116 1726
rect 110 1721 111 1725
rect 115 1721 116 1725
rect 240 1725 241 1729
rect 247 1725 248 1729
rect 240 1724 248 1725
rect 376 1729 384 1730
rect 376 1725 377 1729
rect 383 1725 384 1729
rect 376 1724 384 1725
rect 512 1729 520 1730
rect 512 1725 513 1729
rect 519 1725 520 1729
rect 512 1724 520 1725
rect 648 1729 656 1730
rect 648 1725 649 1729
rect 655 1725 656 1729
rect 648 1724 656 1725
rect 766 1729 772 1730
rect 766 1725 767 1729
rect 771 1728 772 1729
rect 783 1729 789 1730
rect 783 1728 784 1729
rect 771 1726 784 1728
rect 771 1725 772 1726
rect 766 1724 772 1725
rect 783 1725 784 1726
rect 788 1725 789 1729
rect 783 1724 789 1725
rect 1718 1725 1724 1726
rect 110 1720 116 1721
rect 134 1723 140 1724
rect 134 1719 135 1723
rect 139 1719 140 1723
rect 134 1718 140 1719
rect 270 1723 276 1724
rect 270 1719 271 1723
rect 275 1719 276 1723
rect 270 1718 276 1719
rect 406 1723 412 1724
rect 406 1719 407 1723
rect 411 1719 412 1723
rect 406 1718 412 1719
rect 542 1723 548 1724
rect 542 1719 543 1723
rect 547 1719 548 1723
rect 542 1718 548 1719
rect 678 1723 684 1724
rect 678 1719 679 1723
rect 683 1719 684 1723
rect 1718 1721 1719 1725
rect 1723 1721 1724 1725
rect 1718 1720 1724 1721
rect 678 1718 684 1719
rect 158 1708 164 1709
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 158 1704 159 1708
rect 163 1704 164 1708
rect 158 1703 164 1704
rect 294 1708 300 1709
rect 294 1704 295 1708
rect 299 1704 300 1708
rect 294 1703 300 1704
rect 430 1708 436 1709
rect 430 1704 431 1708
rect 435 1704 436 1708
rect 430 1703 436 1704
rect 566 1708 572 1709
rect 566 1704 567 1708
rect 571 1704 572 1708
rect 566 1703 572 1704
rect 702 1708 708 1709
rect 702 1704 703 1708
rect 707 1704 708 1708
rect 702 1703 708 1704
rect 1718 1707 1724 1708
rect 1718 1703 1719 1707
rect 1723 1703 1724 1707
rect 110 1702 116 1703
rect 1718 1702 1724 1703
rect 110 1633 116 1634
rect 1718 1633 1724 1634
rect 110 1629 111 1633
rect 115 1629 116 1633
rect 110 1628 116 1629
rect 246 1632 252 1633
rect 246 1628 247 1632
rect 251 1628 252 1632
rect 246 1627 252 1628
rect 382 1632 388 1633
rect 382 1628 383 1632
rect 387 1628 388 1632
rect 382 1627 388 1628
rect 518 1632 524 1633
rect 518 1628 519 1632
rect 523 1628 524 1632
rect 518 1627 524 1628
rect 654 1632 660 1633
rect 654 1628 655 1632
rect 659 1628 660 1632
rect 654 1627 660 1628
rect 790 1632 796 1633
rect 790 1628 791 1632
rect 795 1628 796 1632
rect 1718 1629 1719 1633
rect 1723 1629 1724 1633
rect 1718 1628 1724 1629
rect 790 1627 796 1628
rect 222 1617 228 1618
rect 110 1615 116 1616
rect 110 1611 111 1615
rect 115 1611 116 1615
rect 222 1613 223 1617
rect 227 1613 228 1617
rect 222 1612 228 1613
rect 358 1617 364 1618
rect 358 1613 359 1617
rect 363 1613 364 1617
rect 358 1612 364 1613
rect 494 1617 500 1618
rect 494 1613 495 1617
rect 499 1613 500 1617
rect 494 1612 500 1613
rect 630 1617 636 1618
rect 630 1613 631 1617
rect 635 1613 636 1617
rect 630 1612 636 1613
rect 766 1617 772 1618
rect 766 1613 767 1617
rect 771 1613 772 1617
rect 766 1612 772 1613
rect 1718 1615 1724 1616
rect 110 1610 116 1611
rect 327 1611 333 1612
rect 327 1607 328 1611
rect 332 1610 333 1611
rect 370 1611 376 1612
rect 370 1610 371 1611
rect 332 1608 371 1610
rect 332 1607 333 1608
rect 327 1606 333 1607
rect 370 1607 371 1608
rect 375 1607 376 1611
rect 370 1606 376 1607
rect 463 1611 469 1612
rect 463 1607 464 1611
rect 468 1610 469 1611
rect 506 1611 512 1612
rect 506 1610 507 1611
rect 468 1608 507 1610
rect 468 1607 469 1608
rect 463 1606 469 1607
rect 506 1607 507 1608
rect 511 1607 512 1611
rect 506 1606 512 1607
rect 599 1611 605 1612
rect 599 1607 600 1611
rect 604 1610 605 1611
rect 642 1611 648 1612
rect 642 1610 643 1611
rect 604 1608 643 1610
rect 604 1607 605 1608
rect 599 1606 605 1607
rect 642 1607 643 1608
rect 647 1607 648 1611
rect 642 1606 648 1607
rect 735 1611 741 1612
rect 735 1607 736 1611
rect 740 1610 741 1611
rect 778 1611 784 1612
rect 778 1610 779 1611
rect 740 1608 779 1610
rect 740 1607 741 1608
rect 735 1606 741 1607
rect 778 1607 779 1608
rect 783 1607 784 1611
rect 871 1611 877 1612
rect 871 1610 872 1611
rect 778 1606 784 1607
rect 788 1608 872 1610
rect 586 1603 592 1604
rect 586 1599 587 1603
rect 591 1602 592 1603
rect 788 1602 790 1608
rect 871 1607 872 1608
rect 876 1607 877 1611
rect 1718 1611 1719 1615
rect 1723 1611 1724 1615
rect 1718 1610 1724 1611
rect 871 1606 877 1607
rect 591 1600 790 1602
rect 591 1599 592 1600
rect 586 1598 592 1599
rect 306 1575 312 1576
rect 306 1571 307 1575
rect 311 1571 312 1575
rect 306 1570 312 1571
rect 370 1575 376 1576
rect 370 1571 371 1575
rect 375 1571 376 1575
rect 370 1570 376 1571
rect 506 1575 512 1576
rect 506 1571 507 1575
rect 511 1571 512 1575
rect 506 1570 512 1571
rect 642 1575 648 1576
rect 642 1571 643 1575
rect 647 1571 648 1575
rect 642 1570 648 1571
rect 778 1575 784 1576
rect 778 1571 779 1575
rect 783 1571 784 1575
rect 778 1570 784 1571
rect 586 1539 592 1540
rect 586 1538 587 1539
rect 573 1536 587 1538
rect 586 1535 587 1536
rect 591 1535 592 1539
rect 586 1534 592 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1538 604 1539
rect 730 1539 736 1540
rect 603 1536 637 1538
rect 603 1535 604 1536
rect 598 1534 604 1535
rect 730 1535 731 1539
rect 735 1538 736 1539
rect 874 1539 880 1540
rect 735 1536 773 1538
rect 735 1535 736 1536
rect 730 1534 736 1535
rect 874 1535 875 1539
rect 879 1538 880 1539
rect 1002 1539 1008 1540
rect 879 1536 909 1538
rect 879 1535 880 1536
rect 874 1534 880 1535
rect 1002 1535 1003 1539
rect 1007 1538 1008 1539
rect 1274 1539 1280 1540
rect 1007 1536 1045 1538
rect 1007 1535 1008 1536
rect 1002 1534 1008 1535
rect 1274 1535 1275 1539
rect 1279 1538 1280 1539
rect 1423 1539 1429 1540
rect 1279 1536 1317 1538
rect 1279 1535 1280 1536
rect 1274 1534 1280 1535
rect 1423 1535 1424 1539
rect 1428 1538 1429 1539
rect 1546 1539 1552 1540
rect 1428 1536 1453 1538
rect 1428 1535 1429 1536
rect 1423 1534 1429 1535
rect 1546 1535 1547 1539
rect 1551 1538 1552 1539
rect 1551 1536 1589 1538
rect 1551 1535 1552 1536
rect 1546 1534 1552 1535
rect 1248 1530 1250 1533
rect 1286 1531 1292 1532
rect 1286 1530 1287 1531
rect 1248 1528 1287 1530
rect 1286 1527 1287 1528
rect 1291 1527 1292 1531
rect 1286 1526 1292 1527
rect 1567 1503 1573 1504
rect 592 1501 604 1502
rect 110 1497 116 1498
rect 110 1493 111 1497
rect 115 1493 116 1497
rect 592 1497 593 1501
rect 597 1497 599 1501
rect 603 1497 604 1501
rect 592 1496 604 1497
rect 728 1501 736 1502
rect 728 1497 729 1501
rect 735 1497 736 1501
rect 728 1496 736 1497
rect 864 1501 870 1502
rect 864 1497 865 1501
rect 869 1500 870 1501
rect 874 1501 880 1502
rect 874 1500 875 1501
rect 869 1498 875 1500
rect 869 1497 870 1498
rect 864 1496 870 1497
rect 874 1497 875 1498
rect 879 1497 880 1501
rect 874 1496 880 1497
rect 1000 1501 1008 1502
rect 1000 1497 1001 1501
rect 1007 1497 1008 1501
rect 1000 1496 1008 1497
rect 1118 1501 1124 1502
rect 1118 1497 1119 1501
rect 1123 1500 1124 1501
rect 1135 1501 1141 1502
rect 1135 1500 1136 1501
rect 1123 1498 1136 1500
rect 1123 1497 1124 1498
rect 1118 1496 1124 1497
rect 1135 1497 1136 1498
rect 1140 1497 1141 1501
rect 1135 1496 1141 1497
rect 1272 1501 1280 1502
rect 1272 1497 1273 1501
rect 1279 1497 1280 1501
rect 1272 1496 1280 1497
rect 1408 1501 1414 1502
rect 1408 1497 1409 1501
rect 1413 1500 1414 1501
rect 1423 1501 1429 1502
rect 1423 1500 1424 1501
rect 1413 1498 1424 1500
rect 1413 1497 1414 1498
rect 1408 1496 1414 1497
rect 1423 1497 1424 1498
rect 1428 1497 1429 1501
rect 1423 1496 1429 1497
rect 1544 1501 1552 1502
rect 1544 1497 1545 1501
rect 1551 1497 1552 1501
rect 1567 1499 1568 1503
rect 1572 1502 1573 1503
rect 1572 1500 1662 1502
rect 1679 1501 1685 1502
rect 1679 1500 1680 1501
rect 1572 1499 1573 1500
rect 1567 1498 1573 1499
rect 1660 1498 1680 1500
rect 1544 1496 1552 1497
rect 1679 1497 1680 1498
rect 1684 1497 1685 1501
rect 1679 1496 1685 1497
rect 1718 1497 1724 1498
rect 110 1492 116 1493
rect 486 1495 492 1496
rect 486 1491 487 1495
rect 491 1491 492 1495
rect 486 1490 492 1491
rect 622 1495 628 1496
rect 622 1491 623 1495
rect 627 1491 628 1495
rect 622 1490 628 1491
rect 758 1495 764 1496
rect 758 1491 759 1495
rect 763 1491 764 1495
rect 758 1490 764 1491
rect 894 1495 900 1496
rect 894 1491 895 1495
rect 899 1491 900 1495
rect 894 1490 900 1491
rect 1030 1495 1036 1496
rect 1030 1491 1031 1495
rect 1035 1491 1036 1495
rect 1030 1490 1036 1491
rect 1166 1495 1172 1496
rect 1166 1491 1167 1495
rect 1171 1491 1172 1495
rect 1166 1490 1172 1491
rect 1302 1495 1308 1496
rect 1302 1491 1303 1495
rect 1307 1491 1308 1495
rect 1302 1490 1308 1491
rect 1438 1495 1444 1496
rect 1438 1491 1439 1495
rect 1443 1491 1444 1495
rect 1438 1490 1444 1491
rect 1574 1495 1580 1496
rect 1574 1491 1575 1495
rect 1579 1491 1580 1495
rect 1718 1493 1719 1497
rect 1723 1493 1724 1497
rect 1718 1492 1724 1493
rect 1574 1490 1580 1491
rect 510 1480 516 1481
rect 110 1479 116 1480
rect 110 1475 111 1479
rect 115 1475 116 1479
rect 510 1476 511 1480
rect 515 1476 516 1480
rect 510 1475 516 1476
rect 646 1480 652 1481
rect 646 1476 647 1480
rect 651 1476 652 1480
rect 646 1475 652 1476
rect 782 1480 788 1481
rect 782 1476 783 1480
rect 787 1476 788 1480
rect 782 1475 788 1476
rect 918 1480 924 1481
rect 918 1476 919 1480
rect 923 1476 924 1480
rect 918 1475 924 1476
rect 1054 1480 1060 1481
rect 1054 1476 1055 1480
rect 1059 1476 1060 1480
rect 1054 1475 1060 1476
rect 1190 1480 1196 1481
rect 1190 1476 1191 1480
rect 1195 1476 1196 1480
rect 1190 1475 1196 1476
rect 1326 1480 1332 1481
rect 1326 1476 1327 1480
rect 1331 1476 1332 1480
rect 1326 1475 1332 1476
rect 1462 1480 1468 1481
rect 1462 1476 1463 1480
rect 1467 1476 1468 1480
rect 1462 1475 1468 1476
rect 1598 1480 1604 1481
rect 1598 1476 1599 1480
rect 1603 1476 1604 1480
rect 1598 1475 1604 1476
rect 1718 1479 1724 1480
rect 1718 1475 1719 1479
rect 1723 1475 1724 1479
rect 110 1474 116 1475
rect 1718 1474 1724 1475
rect 110 1405 116 1406
rect 1718 1405 1724 1406
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 110 1400 116 1401
rect 742 1404 748 1405
rect 742 1400 743 1404
rect 747 1400 748 1404
rect 742 1399 748 1400
rect 886 1404 892 1405
rect 886 1400 887 1404
rect 891 1400 892 1404
rect 886 1399 892 1400
rect 1030 1404 1036 1405
rect 1030 1400 1031 1404
rect 1035 1400 1036 1404
rect 1030 1399 1036 1400
rect 1174 1404 1180 1405
rect 1174 1400 1175 1404
rect 1179 1400 1180 1404
rect 1174 1399 1180 1400
rect 1318 1404 1324 1405
rect 1318 1400 1319 1404
rect 1323 1400 1324 1404
rect 1318 1399 1324 1400
rect 1462 1404 1468 1405
rect 1462 1400 1463 1404
rect 1467 1400 1468 1404
rect 1462 1399 1468 1400
rect 1598 1404 1604 1405
rect 1598 1400 1599 1404
rect 1603 1400 1604 1404
rect 1718 1401 1719 1405
rect 1723 1401 1724 1405
rect 1718 1400 1724 1401
rect 1598 1399 1604 1400
rect 718 1389 724 1390
rect 110 1387 116 1388
rect 110 1383 111 1387
rect 115 1383 116 1387
rect 718 1385 719 1389
rect 723 1385 724 1389
rect 718 1384 724 1385
rect 862 1389 868 1390
rect 862 1385 863 1389
rect 867 1385 868 1389
rect 862 1384 868 1385
rect 1006 1389 1012 1390
rect 1006 1385 1007 1389
rect 1011 1385 1012 1389
rect 1006 1384 1012 1385
rect 1150 1389 1156 1390
rect 1150 1385 1151 1389
rect 1155 1385 1156 1389
rect 1150 1384 1156 1385
rect 1294 1389 1300 1390
rect 1294 1385 1295 1389
rect 1299 1385 1300 1389
rect 1294 1384 1300 1385
rect 1438 1389 1444 1390
rect 1438 1385 1439 1389
rect 1443 1385 1444 1389
rect 1438 1384 1444 1385
rect 1574 1389 1580 1390
rect 1574 1385 1575 1389
rect 1579 1385 1580 1389
rect 1574 1384 1580 1385
rect 1718 1387 1724 1388
rect 110 1382 116 1383
rect 823 1383 829 1384
rect 823 1379 824 1383
rect 828 1382 829 1383
rect 874 1383 880 1384
rect 874 1382 875 1383
rect 828 1380 875 1382
rect 828 1379 829 1380
rect 823 1378 829 1379
rect 874 1379 875 1380
rect 879 1379 880 1383
rect 874 1378 880 1379
rect 967 1383 973 1384
rect 967 1379 968 1383
rect 972 1382 973 1383
rect 1018 1383 1024 1384
rect 1018 1382 1019 1383
rect 972 1380 1019 1382
rect 972 1379 973 1380
rect 967 1378 973 1379
rect 1018 1379 1019 1380
rect 1023 1379 1024 1383
rect 1018 1378 1024 1379
rect 1111 1383 1117 1384
rect 1111 1379 1112 1383
rect 1116 1382 1117 1383
rect 1162 1383 1168 1384
rect 1162 1382 1163 1383
rect 1116 1380 1163 1382
rect 1116 1379 1117 1380
rect 1111 1378 1117 1379
rect 1162 1379 1163 1380
rect 1167 1379 1168 1383
rect 1162 1378 1168 1379
rect 1255 1383 1264 1384
rect 1255 1379 1256 1383
rect 1263 1379 1264 1383
rect 1255 1378 1264 1379
rect 1286 1383 1292 1384
rect 1286 1379 1287 1383
rect 1291 1382 1292 1383
rect 1399 1383 1405 1384
rect 1399 1382 1400 1383
rect 1291 1380 1400 1382
rect 1291 1379 1292 1380
rect 1286 1378 1292 1379
rect 1399 1379 1400 1380
rect 1404 1379 1405 1383
rect 1399 1378 1405 1379
rect 1543 1383 1549 1384
rect 1543 1379 1544 1383
rect 1548 1382 1549 1383
rect 1586 1383 1592 1384
rect 1586 1382 1587 1383
rect 1548 1380 1587 1382
rect 1548 1379 1549 1380
rect 1543 1378 1549 1379
rect 1586 1379 1587 1380
rect 1591 1379 1592 1383
rect 1586 1378 1592 1379
rect 1674 1383 1685 1384
rect 1674 1379 1675 1383
rect 1679 1379 1680 1383
rect 1684 1379 1685 1383
rect 1718 1383 1719 1387
rect 1723 1383 1724 1387
rect 1718 1382 1724 1383
rect 1674 1378 1685 1379
rect 1118 1363 1124 1364
rect 1118 1362 1119 1363
rect 864 1360 1119 1362
rect 864 1346 866 1360
rect 1118 1359 1119 1360
rect 1123 1359 1124 1363
rect 1118 1358 1124 1359
rect 805 1344 866 1346
rect 874 1347 880 1348
rect 874 1343 875 1347
rect 879 1343 880 1347
rect 874 1342 880 1343
rect 1018 1347 1024 1348
rect 1018 1343 1019 1347
rect 1023 1343 1024 1347
rect 1018 1342 1024 1343
rect 1162 1347 1168 1348
rect 1162 1343 1163 1347
rect 1167 1343 1168 1347
rect 1162 1342 1168 1343
rect 1378 1347 1384 1348
rect 1378 1343 1379 1347
rect 1383 1343 1384 1347
rect 1567 1347 1573 1348
rect 1567 1346 1568 1347
rect 1525 1344 1568 1346
rect 1378 1342 1384 1343
rect 1567 1343 1568 1344
rect 1572 1343 1573 1347
rect 1567 1342 1573 1343
rect 1586 1347 1592 1348
rect 1586 1343 1587 1347
rect 1591 1343 1592 1347
rect 1586 1342 1592 1343
rect 358 1315 364 1316
rect 358 1314 359 1315
rect 269 1312 359 1314
rect 358 1311 359 1312
rect 363 1311 364 1315
rect 530 1315 536 1316
rect 530 1314 531 1315
rect 501 1312 531 1314
rect 358 1310 364 1311
rect 530 1311 531 1312
rect 535 1311 536 1315
rect 886 1315 892 1316
rect 886 1314 887 1315
rect 765 1312 887 1314
rect 530 1310 536 1311
rect 886 1311 887 1312
rect 891 1311 892 1315
rect 1190 1315 1196 1316
rect 1190 1314 1191 1315
rect 1061 1312 1191 1314
rect 886 1310 892 1311
rect 1190 1311 1191 1312
rect 1195 1311 1196 1315
rect 1190 1310 1196 1311
rect 1258 1315 1264 1316
rect 1258 1311 1259 1315
rect 1263 1314 1264 1315
rect 1674 1315 1680 1316
rect 1674 1314 1675 1315
rect 1263 1312 1301 1314
rect 1661 1312 1675 1314
rect 1263 1311 1264 1312
rect 1258 1310 1264 1311
rect 1674 1311 1675 1312
rect 1679 1311 1680 1315
rect 1674 1310 1680 1311
rect 358 1279 364 1280
rect 270 1277 276 1278
rect 110 1273 116 1274
rect 110 1269 111 1273
rect 115 1269 116 1273
rect 270 1273 271 1277
rect 275 1276 276 1277
rect 287 1277 293 1278
rect 287 1276 288 1277
rect 275 1274 288 1276
rect 275 1273 276 1274
rect 270 1272 276 1273
rect 287 1273 288 1274
rect 292 1273 293 1277
rect 358 1275 359 1279
rect 363 1278 364 1279
rect 530 1279 536 1280
rect 363 1276 502 1278
rect 519 1277 525 1278
rect 519 1276 520 1277
rect 363 1275 364 1276
rect 358 1274 364 1275
rect 500 1274 520 1276
rect 287 1272 293 1273
rect 519 1273 520 1274
rect 524 1273 525 1277
rect 530 1275 531 1279
rect 535 1278 536 1279
rect 886 1279 892 1280
rect 535 1276 766 1278
rect 783 1277 789 1278
rect 783 1276 784 1277
rect 535 1275 536 1276
rect 530 1274 536 1275
rect 764 1274 784 1276
rect 519 1272 525 1273
rect 783 1273 784 1274
rect 788 1273 789 1277
rect 886 1275 887 1279
rect 891 1278 892 1279
rect 1190 1279 1196 1280
rect 891 1276 1062 1278
rect 1079 1277 1085 1278
rect 1079 1276 1080 1277
rect 891 1275 892 1276
rect 886 1274 892 1275
rect 1060 1274 1080 1276
rect 783 1272 789 1273
rect 1079 1273 1080 1274
rect 1084 1273 1085 1277
rect 1190 1275 1191 1279
rect 1195 1278 1196 1279
rect 1195 1276 1374 1278
rect 1391 1277 1397 1278
rect 1391 1276 1392 1277
rect 1195 1275 1196 1276
rect 1190 1274 1196 1275
rect 1372 1274 1392 1276
rect 1079 1272 1085 1273
rect 1391 1273 1392 1274
rect 1396 1273 1397 1277
rect 1391 1272 1397 1273
rect 1666 1277 1672 1278
rect 1666 1273 1667 1277
rect 1671 1276 1672 1277
rect 1679 1277 1685 1278
rect 1679 1276 1680 1277
rect 1671 1274 1680 1276
rect 1671 1273 1672 1274
rect 1666 1272 1672 1273
rect 1679 1273 1680 1274
rect 1684 1273 1685 1277
rect 1679 1272 1685 1273
rect 1718 1273 1724 1274
rect 110 1268 116 1269
rect 182 1271 188 1272
rect 182 1267 183 1271
rect 187 1267 188 1271
rect 182 1266 188 1267
rect 414 1271 420 1272
rect 414 1267 415 1271
rect 419 1267 420 1271
rect 414 1266 420 1267
rect 678 1271 684 1272
rect 678 1267 679 1271
rect 683 1267 684 1271
rect 678 1266 684 1267
rect 974 1271 980 1272
rect 974 1267 975 1271
rect 979 1267 980 1271
rect 974 1266 980 1267
rect 1286 1271 1292 1272
rect 1286 1267 1287 1271
rect 1291 1267 1292 1271
rect 1286 1266 1292 1267
rect 1574 1271 1580 1272
rect 1574 1267 1575 1271
rect 1579 1267 1580 1271
rect 1718 1269 1719 1273
rect 1723 1269 1724 1273
rect 1718 1268 1724 1269
rect 1574 1266 1580 1267
rect 206 1256 212 1257
rect 110 1255 116 1256
rect 110 1251 111 1255
rect 115 1251 116 1255
rect 206 1252 207 1256
rect 211 1252 212 1256
rect 206 1251 212 1252
rect 438 1256 444 1257
rect 438 1252 439 1256
rect 443 1252 444 1256
rect 438 1251 444 1252
rect 702 1256 708 1257
rect 702 1252 703 1256
rect 707 1252 708 1256
rect 702 1251 708 1252
rect 998 1256 1004 1257
rect 998 1252 999 1256
rect 1003 1252 1004 1256
rect 998 1251 1004 1252
rect 1310 1256 1316 1257
rect 1310 1252 1311 1256
rect 1315 1252 1316 1256
rect 1310 1251 1316 1252
rect 1598 1256 1604 1257
rect 1598 1252 1599 1256
rect 1603 1252 1604 1256
rect 1598 1251 1604 1252
rect 1718 1255 1724 1256
rect 1718 1251 1719 1255
rect 1723 1251 1724 1255
rect 110 1250 116 1251
rect 1718 1250 1724 1251
rect 110 1193 116 1194
rect 1718 1193 1724 1194
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 110 1188 116 1189
rect 158 1192 164 1193
rect 158 1188 159 1192
rect 163 1188 164 1192
rect 158 1187 164 1188
rect 334 1192 340 1193
rect 334 1188 335 1192
rect 339 1188 340 1192
rect 334 1187 340 1188
rect 558 1192 564 1193
rect 558 1188 559 1192
rect 563 1188 564 1192
rect 558 1187 564 1188
rect 798 1192 804 1193
rect 798 1188 799 1192
rect 803 1188 804 1192
rect 798 1187 804 1188
rect 1062 1192 1068 1193
rect 1062 1188 1063 1192
rect 1067 1188 1068 1192
rect 1062 1187 1068 1188
rect 1334 1192 1340 1193
rect 1334 1188 1335 1192
rect 1339 1188 1340 1192
rect 1334 1187 1340 1188
rect 1598 1192 1604 1193
rect 1598 1188 1599 1192
rect 1603 1188 1604 1192
rect 1718 1189 1719 1193
rect 1723 1189 1724 1193
rect 1718 1188 1724 1189
rect 1598 1187 1604 1188
rect 134 1177 140 1178
rect 110 1175 116 1176
rect 110 1171 111 1175
rect 115 1171 116 1175
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 310 1177 316 1178
rect 310 1173 311 1177
rect 315 1173 316 1177
rect 310 1172 316 1173
rect 534 1177 540 1178
rect 534 1173 535 1177
rect 539 1173 540 1177
rect 534 1172 540 1173
rect 774 1177 780 1178
rect 774 1173 775 1177
rect 779 1173 780 1177
rect 774 1172 780 1173
rect 1038 1177 1044 1178
rect 1038 1173 1039 1177
rect 1043 1173 1044 1177
rect 1038 1172 1044 1173
rect 1310 1177 1316 1178
rect 1310 1173 1311 1177
rect 1315 1173 1316 1177
rect 1310 1172 1316 1173
rect 1574 1177 1580 1178
rect 1574 1173 1575 1177
rect 1579 1173 1580 1177
rect 1574 1172 1580 1173
rect 1718 1175 1724 1176
rect 110 1170 116 1171
rect 239 1171 245 1172
rect 239 1167 240 1171
rect 244 1170 245 1171
rect 322 1171 328 1172
rect 322 1170 323 1171
rect 244 1168 323 1170
rect 244 1167 245 1168
rect 239 1166 245 1167
rect 322 1167 323 1168
rect 327 1167 328 1171
rect 322 1166 328 1167
rect 415 1171 421 1172
rect 415 1167 416 1171
rect 420 1170 421 1171
rect 546 1171 552 1172
rect 546 1170 547 1171
rect 420 1168 547 1170
rect 420 1167 421 1168
rect 415 1166 421 1167
rect 546 1167 547 1168
rect 551 1167 552 1171
rect 546 1166 552 1167
rect 639 1171 645 1172
rect 639 1167 640 1171
rect 644 1170 645 1171
rect 786 1171 792 1172
rect 786 1170 787 1171
rect 644 1168 787 1170
rect 644 1167 645 1168
rect 639 1166 645 1167
rect 786 1167 787 1168
rect 791 1167 792 1171
rect 786 1166 792 1167
rect 879 1171 885 1172
rect 879 1167 880 1171
rect 884 1170 885 1171
rect 1050 1171 1056 1172
rect 1050 1170 1051 1171
rect 884 1168 1051 1170
rect 884 1167 885 1168
rect 879 1166 885 1167
rect 1050 1167 1051 1168
rect 1055 1167 1056 1171
rect 1050 1166 1056 1167
rect 1090 1171 1096 1172
rect 1090 1167 1091 1171
rect 1095 1170 1096 1171
rect 1143 1171 1149 1172
rect 1143 1170 1144 1171
rect 1095 1168 1144 1170
rect 1095 1167 1096 1168
rect 1090 1166 1096 1167
rect 1143 1167 1144 1168
rect 1148 1167 1149 1171
rect 1143 1166 1149 1167
rect 1378 1171 1384 1172
rect 1378 1167 1379 1171
rect 1383 1170 1384 1171
rect 1415 1171 1421 1172
rect 1415 1170 1416 1171
rect 1383 1168 1416 1170
rect 1383 1167 1384 1168
rect 1378 1166 1384 1167
rect 1415 1167 1416 1168
rect 1420 1167 1421 1171
rect 1415 1166 1421 1167
rect 1658 1171 1664 1172
rect 1658 1167 1659 1171
rect 1663 1170 1664 1171
rect 1679 1171 1685 1172
rect 1679 1170 1680 1171
rect 1663 1168 1680 1170
rect 1663 1167 1664 1168
rect 1658 1166 1664 1167
rect 1679 1167 1680 1168
rect 1684 1167 1685 1171
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1718 1170 1724 1171
rect 1679 1166 1685 1167
rect 270 1135 276 1136
rect 270 1134 271 1135
rect 221 1132 271 1134
rect 270 1131 271 1132
rect 275 1131 276 1135
rect 270 1130 276 1131
rect 322 1135 328 1136
rect 322 1131 323 1135
rect 327 1131 328 1135
rect 322 1130 328 1131
rect 546 1135 552 1136
rect 546 1131 547 1135
rect 551 1131 552 1135
rect 546 1130 552 1131
rect 786 1135 792 1136
rect 786 1131 787 1135
rect 791 1131 792 1135
rect 786 1130 792 1131
rect 1050 1135 1056 1136
rect 1050 1131 1051 1135
rect 1055 1131 1056 1135
rect 1050 1130 1056 1131
rect 1374 1135 1380 1136
rect 1374 1131 1375 1135
rect 1379 1131 1380 1135
rect 1666 1135 1672 1136
rect 1666 1134 1667 1135
rect 1661 1132 1667 1134
rect 1374 1130 1380 1131
rect 1666 1131 1667 1132
rect 1671 1131 1672 1135
rect 1666 1130 1672 1131
rect 1090 1107 1096 1108
rect 1090 1106 1091 1107
rect 324 1104 1091 1106
rect 324 1094 326 1104
rect 1090 1103 1091 1104
rect 1095 1103 1096 1107
rect 1090 1102 1096 1103
rect 309 1092 326 1094
rect 330 1095 336 1096
rect 330 1091 331 1095
rect 335 1094 336 1095
rect 586 1095 592 1096
rect 335 1092 477 1094
rect 335 1091 336 1092
rect 330 1090 336 1091
rect 586 1091 587 1095
rect 591 1094 592 1095
rect 842 1095 848 1096
rect 591 1092 733 1094
rect 591 1091 592 1092
rect 586 1090 592 1091
rect 842 1091 843 1095
rect 847 1094 848 1095
rect 1454 1095 1460 1096
rect 1454 1094 1455 1095
rect 847 1092 1005 1094
rect 1357 1092 1455 1094
rect 847 1091 848 1092
rect 842 1090 848 1091
rect 1454 1091 1455 1092
rect 1459 1091 1460 1095
rect 1658 1095 1664 1096
rect 1658 1094 1659 1095
rect 1645 1092 1659 1094
rect 1454 1090 1460 1091
rect 1658 1091 1659 1092
rect 1663 1091 1664 1095
rect 1658 1090 1664 1091
rect 328 1057 336 1058
rect 110 1053 116 1054
rect 110 1049 111 1053
rect 115 1049 116 1053
rect 328 1053 329 1057
rect 335 1053 336 1057
rect 328 1052 336 1053
rect 568 1057 574 1058
rect 568 1053 569 1057
rect 573 1056 574 1057
rect 586 1057 592 1058
rect 586 1056 587 1057
rect 573 1054 587 1056
rect 573 1053 574 1054
rect 568 1052 574 1053
rect 586 1053 587 1054
rect 591 1053 592 1057
rect 586 1052 592 1053
rect 824 1057 830 1058
rect 824 1053 825 1057
rect 829 1056 830 1057
rect 842 1057 848 1058
rect 842 1056 843 1057
rect 829 1054 843 1056
rect 829 1053 830 1054
rect 824 1052 830 1053
rect 842 1053 843 1054
rect 847 1053 848 1057
rect 842 1052 848 1053
rect 1094 1057 1101 1058
rect 1094 1053 1095 1057
rect 1100 1053 1101 1057
rect 1094 1052 1101 1053
rect 1374 1057 1381 1058
rect 1374 1053 1375 1057
rect 1380 1053 1381 1057
rect 1374 1052 1381 1053
rect 1646 1057 1652 1058
rect 1646 1053 1647 1057
rect 1651 1056 1652 1057
rect 1663 1057 1669 1058
rect 1663 1056 1664 1057
rect 1651 1054 1664 1056
rect 1651 1053 1652 1054
rect 1646 1052 1652 1053
rect 1663 1053 1664 1054
rect 1668 1053 1669 1057
rect 1663 1052 1669 1053
rect 1718 1053 1724 1054
rect 110 1048 116 1049
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 462 1051 468 1052
rect 462 1047 463 1051
rect 467 1047 468 1051
rect 462 1046 468 1047
rect 718 1051 724 1052
rect 718 1047 719 1051
rect 723 1047 724 1051
rect 718 1046 724 1047
rect 990 1051 996 1052
rect 990 1047 991 1051
rect 995 1047 996 1051
rect 990 1046 996 1047
rect 1270 1051 1276 1052
rect 1270 1047 1271 1051
rect 1275 1047 1276 1051
rect 1270 1046 1276 1047
rect 1558 1051 1564 1052
rect 1558 1047 1559 1051
rect 1563 1047 1564 1051
rect 1718 1049 1719 1053
rect 1723 1049 1724 1053
rect 1718 1048 1724 1049
rect 1558 1046 1564 1047
rect 246 1036 252 1037
rect 110 1035 116 1036
rect 110 1031 111 1035
rect 115 1031 116 1035
rect 246 1032 247 1036
rect 251 1032 252 1036
rect 246 1031 252 1032
rect 486 1036 492 1037
rect 486 1032 487 1036
rect 491 1032 492 1036
rect 486 1031 492 1032
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 1014 1036 1020 1037
rect 1014 1032 1015 1036
rect 1019 1032 1020 1036
rect 1014 1031 1020 1032
rect 1294 1036 1300 1037
rect 1294 1032 1295 1036
rect 1299 1032 1300 1036
rect 1294 1031 1300 1032
rect 1582 1036 1588 1037
rect 1582 1032 1583 1036
rect 1587 1032 1588 1036
rect 1582 1031 1588 1032
rect 1718 1035 1724 1036
rect 1718 1031 1719 1035
rect 1723 1031 1724 1035
rect 110 1030 116 1031
rect 1718 1030 1724 1031
rect 558 991 564 992
rect 558 987 559 991
rect 563 990 564 991
rect 1094 991 1100 992
rect 1094 990 1095 991
rect 563 988 1095 990
rect 563 987 564 988
rect 558 986 564 987
rect 1094 987 1095 988
rect 1099 987 1100 991
rect 1094 986 1100 987
rect 110 977 116 978
rect 1718 977 1724 978
rect 110 973 111 977
rect 115 973 116 977
rect 110 972 116 973
rect 462 976 468 977
rect 462 972 463 976
rect 467 972 468 976
rect 462 971 468 972
rect 646 976 652 977
rect 646 972 647 976
rect 651 972 652 976
rect 646 971 652 972
rect 854 976 860 977
rect 854 972 855 976
rect 859 972 860 976
rect 854 971 860 972
rect 1078 976 1084 977
rect 1078 972 1079 976
rect 1083 972 1084 976
rect 1078 971 1084 972
rect 1310 976 1316 977
rect 1310 972 1311 976
rect 1315 972 1316 976
rect 1310 971 1316 972
rect 1542 976 1548 977
rect 1542 972 1543 976
rect 1547 972 1548 976
rect 1718 973 1719 977
rect 1723 973 1724 977
rect 1718 972 1724 973
rect 1542 971 1548 972
rect 438 961 444 962
rect 110 959 116 960
rect 110 955 111 959
rect 115 955 116 959
rect 438 957 439 961
rect 443 957 444 961
rect 438 956 444 957
rect 622 961 628 962
rect 622 957 623 961
rect 627 957 628 961
rect 622 956 628 957
rect 830 961 836 962
rect 830 957 831 961
rect 835 957 836 961
rect 830 956 836 957
rect 1054 961 1060 962
rect 1054 957 1055 961
rect 1059 957 1060 961
rect 1054 956 1060 957
rect 1286 961 1292 962
rect 1286 957 1287 961
rect 1291 957 1292 961
rect 1286 956 1292 957
rect 1518 961 1524 962
rect 1518 957 1519 961
rect 1523 957 1524 961
rect 1518 956 1524 957
rect 1718 959 1724 960
rect 110 954 116 955
rect 543 955 549 956
rect 543 951 544 955
rect 548 954 549 955
rect 634 955 640 956
rect 634 954 635 955
rect 548 952 635 954
rect 548 951 549 952
rect 543 950 549 951
rect 634 951 635 952
rect 639 951 640 955
rect 634 950 640 951
rect 727 955 733 956
rect 727 951 728 955
rect 732 954 733 955
rect 842 955 848 956
rect 842 954 843 955
rect 732 952 843 954
rect 732 951 733 952
rect 727 950 733 951
rect 842 951 843 952
rect 847 951 848 955
rect 842 950 848 951
rect 935 955 941 956
rect 935 951 936 955
rect 940 954 941 955
rect 1066 955 1072 956
rect 1066 954 1067 955
rect 940 952 1067 954
rect 940 951 941 952
rect 935 950 941 951
rect 1066 951 1067 952
rect 1071 951 1072 955
rect 1066 950 1072 951
rect 1159 955 1165 956
rect 1159 951 1160 955
rect 1164 954 1165 955
rect 1298 955 1304 956
rect 1298 954 1299 955
rect 1164 952 1299 954
rect 1164 951 1165 952
rect 1159 950 1165 951
rect 1298 951 1299 952
rect 1303 951 1304 955
rect 1391 955 1397 956
rect 1391 954 1392 955
rect 1298 950 1304 951
rect 1308 952 1392 954
rect 786 947 792 948
rect 786 943 787 947
rect 791 946 792 947
rect 1308 946 1310 952
rect 1391 951 1392 952
rect 1396 951 1397 955
rect 1391 950 1397 951
rect 1602 955 1608 956
rect 1602 951 1603 955
rect 1607 954 1608 955
rect 1623 955 1629 956
rect 1623 954 1624 955
rect 1607 952 1624 954
rect 1607 951 1608 952
rect 1602 950 1608 951
rect 1623 951 1624 952
rect 1628 951 1629 955
rect 1718 955 1719 959
rect 1723 955 1724 959
rect 1718 954 1724 955
rect 1623 950 1629 951
rect 791 944 1310 946
rect 791 943 792 944
rect 786 942 792 943
rect 558 919 564 920
rect 558 918 559 919
rect 525 916 559 918
rect 558 915 559 916
rect 563 915 564 919
rect 558 914 564 915
rect 634 919 640 920
rect 634 915 635 919
rect 639 915 640 919
rect 634 914 640 915
rect 842 919 848 920
rect 842 915 843 919
rect 847 915 848 919
rect 842 914 848 915
rect 1066 919 1072 920
rect 1066 915 1067 919
rect 1071 915 1072 919
rect 1066 914 1072 915
rect 1298 919 1304 920
rect 1298 915 1299 919
rect 1303 915 1304 919
rect 1646 919 1652 920
rect 1646 918 1647 919
rect 1605 916 1647 918
rect 1298 914 1304 915
rect 1646 915 1647 916
rect 1651 915 1652 919
rect 1646 914 1652 915
rect 786 887 792 888
rect 786 886 787 887
rect 773 884 787 886
rect 786 883 787 884
rect 791 883 792 887
rect 786 882 792 883
rect 794 887 800 888
rect 794 883 795 887
rect 799 886 800 887
rect 930 887 936 888
rect 799 884 837 886
rect 799 883 800 884
rect 794 882 800 883
rect 930 883 931 887
rect 935 886 936 887
rect 1066 887 1072 888
rect 935 884 973 886
rect 935 883 936 884
rect 930 882 936 883
rect 1066 883 1067 887
rect 1071 886 1072 887
rect 1202 887 1208 888
rect 1071 884 1109 886
rect 1071 883 1072 884
rect 1066 882 1072 883
rect 1202 883 1203 887
rect 1207 886 1208 887
rect 1602 887 1608 888
rect 1602 886 1603 887
rect 1207 884 1245 886
rect 1589 884 1603 886
rect 1207 883 1208 884
rect 1202 882 1208 883
rect 1450 883 1456 884
rect 1450 879 1451 883
rect 1455 879 1456 883
rect 1602 883 1603 884
rect 1607 883 1608 887
rect 1602 882 1608 883
rect 1450 878 1456 879
rect 792 849 800 850
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 792 845 793 849
rect 799 845 800 849
rect 792 844 800 845
rect 928 849 936 850
rect 928 845 929 849
rect 935 845 936 849
rect 928 844 936 845
rect 1064 849 1072 850
rect 1064 845 1065 849
rect 1071 845 1072 849
rect 1064 844 1072 845
rect 1200 849 1208 850
rect 1200 845 1201 849
rect 1207 845 1208 849
rect 1200 844 1208 845
rect 1318 849 1324 850
rect 1318 845 1319 849
rect 1323 848 1324 849
rect 1335 849 1341 850
rect 1335 848 1336 849
rect 1323 846 1336 848
rect 1323 845 1324 846
rect 1318 844 1324 845
rect 1335 845 1336 846
rect 1340 845 1341 849
rect 1335 844 1341 845
rect 1458 849 1464 850
rect 1458 845 1459 849
rect 1463 848 1464 849
rect 1471 849 1477 850
rect 1471 848 1472 849
rect 1463 846 1472 848
rect 1463 845 1464 846
rect 1458 844 1464 845
rect 1471 845 1472 846
rect 1476 845 1477 849
rect 1471 844 1477 845
rect 1590 849 1596 850
rect 1590 845 1591 849
rect 1595 848 1596 849
rect 1607 849 1613 850
rect 1607 848 1608 849
rect 1595 846 1608 848
rect 1595 845 1596 846
rect 1590 844 1596 845
rect 1607 845 1608 846
rect 1612 845 1613 849
rect 1607 844 1613 845
rect 1718 845 1724 846
rect 110 840 116 841
rect 686 843 692 844
rect 686 839 687 843
rect 691 839 692 843
rect 686 838 692 839
rect 822 843 828 844
rect 822 839 823 843
rect 827 839 828 843
rect 822 838 828 839
rect 958 843 964 844
rect 958 839 959 843
rect 963 839 964 843
rect 958 838 964 839
rect 1094 843 1100 844
rect 1094 839 1095 843
rect 1099 839 1100 843
rect 1094 838 1100 839
rect 1230 843 1236 844
rect 1230 839 1231 843
rect 1235 839 1236 843
rect 1230 838 1236 839
rect 1366 843 1372 844
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 1502 843 1508 844
rect 1502 839 1503 843
rect 1507 839 1508 843
rect 1718 841 1719 845
rect 1723 841 1724 845
rect 1718 840 1724 841
rect 1502 838 1508 839
rect 710 828 716 829
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 710 824 711 828
rect 715 824 716 828
rect 710 823 716 824
rect 846 828 852 829
rect 846 824 847 828
rect 851 824 852 828
rect 846 823 852 824
rect 982 828 988 829
rect 982 824 983 828
rect 987 824 988 828
rect 982 823 988 824
rect 1118 828 1124 829
rect 1118 824 1119 828
rect 1123 824 1124 828
rect 1118 823 1124 824
rect 1254 828 1260 829
rect 1254 824 1255 828
rect 1259 824 1260 828
rect 1254 823 1260 824
rect 1390 828 1396 829
rect 1390 824 1391 828
rect 1395 824 1396 828
rect 1390 823 1396 824
rect 1526 828 1532 829
rect 1526 824 1527 828
rect 1531 824 1532 828
rect 1526 823 1532 824
rect 1718 827 1724 828
rect 1718 823 1719 827
rect 1723 823 1724 827
rect 110 822 116 823
rect 1718 822 1724 823
rect 110 757 116 758
rect 1718 757 1724 758
rect 110 753 111 757
rect 115 753 116 757
rect 110 752 116 753
rect 814 756 820 757
rect 814 752 815 756
rect 819 752 820 756
rect 814 751 820 752
rect 950 756 956 757
rect 950 752 951 756
rect 955 752 956 756
rect 950 751 956 752
rect 1086 756 1092 757
rect 1086 752 1087 756
rect 1091 752 1092 756
rect 1086 751 1092 752
rect 1222 756 1228 757
rect 1222 752 1223 756
rect 1227 752 1228 756
rect 1222 751 1228 752
rect 1358 756 1364 757
rect 1358 752 1359 756
rect 1363 752 1364 756
rect 1358 751 1364 752
rect 1494 756 1500 757
rect 1494 752 1495 756
rect 1499 752 1500 756
rect 1718 753 1719 757
rect 1723 753 1724 757
rect 1718 752 1724 753
rect 1494 751 1500 752
rect 790 741 796 742
rect 110 739 116 740
rect 110 735 111 739
rect 115 735 116 739
rect 790 737 791 741
rect 795 737 796 741
rect 790 736 796 737
rect 926 741 932 742
rect 926 737 927 741
rect 931 737 932 741
rect 926 736 932 737
rect 1062 741 1068 742
rect 1062 737 1063 741
rect 1067 737 1068 741
rect 1062 736 1068 737
rect 1198 741 1204 742
rect 1198 737 1199 741
rect 1203 737 1204 741
rect 1198 736 1204 737
rect 1334 741 1340 742
rect 1334 737 1335 741
rect 1339 737 1340 741
rect 1334 736 1340 737
rect 1470 741 1476 742
rect 1470 737 1471 741
rect 1475 737 1476 741
rect 1470 736 1476 737
rect 1718 739 1724 740
rect 110 734 116 735
rect 895 735 901 736
rect 895 731 896 735
rect 900 734 901 735
rect 938 735 944 736
rect 938 734 939 735
rect 900 732 939 734
rect 900 731 901 732
rect 895 730 901 731
rect 938 731 939 732
rect 943 731 944 735
rect 938 730 944 731
rect 1022 735 1028 736
rect 1022 731 1023 735
rect 1027 734 1028 735
rect 1031 735 1037 736
rect 1031 734 1032 735
rect 1027 732 1032 734
rect 1027 731 1028 732
rect 1022 730 1028 731
rect 1031 731 1032 732
rect 1036 731 1037 735
rect 1031 730 1037 731
rect 1098 735 1104 736
rect 1098 731 1099 735
rect 1103 734 1104 735
rect 1167 735 1173 736
rect 1167 734 1168 735
rect 1103 732 1168 734
rect 1103 731 1104 732
rect 1098 730 1104 731
rect 1167 731 1168 732
rect 1172 731 1173 735
rect 1167 730 1173 731
rect 1178 735 1184 736
rect 1178 731 1179 735
rect 1183 734 1184 735
rect 1303 735 1309 736
rect 1303 734 1304 735
rect 1183 732 1304 734
rect 1183 731 1184 732
rect 1178 730 1184 731
rect 1303 731 1304 732
rect 1308 731 1309 735
rect 1303 730 1309 731
rect 1439 735 1445 736
rect 1439 731 1440 735
rect 1444 734 1445 735
rect 1450 735 1456 736
rect 1450 734 1451 735
rect 1444 732 1451 734
rect 1444 731 1445 732
rect 1439 730 1445 731
rect 1450 731 1451 732
rect 1455 731 1456 735
rect 1450 730 1456 731
rect 1506 735 1512 736
rect 1506 731 1507 735
rect 1511 734 1512 735
rect 1575 735 1581 736
rect 1575 734 1576 735
rect 1511 732 1576 734
rect 1511 731 1512 732
rect 1506 730 1512 731
rect 1575 731 1576 732
rect 1580 731 1581 735
rect 1718 735 1719 739
rect 1723 735 1724 739
rect 1718 734 1724 735
rect 1575 730 1581 731
rect 874 699 880 700
rect 874 695 875 699
rect 879 695 880 699
rect 874 694 880 695
rect 938 699 944 700
rect 938 695 939 699
rect 943 695 944 699
rect 1178 699 1184 700
rect 1178 698 1179 699
rect 1149 696 1179 698
rect 938 694 944 695
rect 1178 695 1179 696
rect 1183 695 1184 699
rect 1318 699 1324 700
rect 1318 698 1319 699
rect 1285 696 1319 698
rect 1178 694 1184 695
rect 1318 695 1319 696
rect 1323 695 1324 699
rect 1318 694 1324 695
rect 1326 699 1332 700
rect 1326 695 1327 699
rect 1331 698 1332 699
rect 1590 699 1596 700
rect 1590 698 1591 699
rect 1331 696 1349 698
rect 1557 696 1591 698
rect 1331 695 1332 696
rect 1326 694 1332 695
rect 1590 695 1591 696
rect 1595 695 1596 699
rect 1590 694 1596 695
rect 638 667 644 668
rect 594 663 600 664
rect 594 659 595 663
rect 599 659 600 663
rect 638 663 639 667
rect 643 666 644 667
rect 999 667 1005 668
rect 999 666 1000 667
rect 643 664 693 666
rect 941 664 1000 666
rect 643 663 644 664
rect 638 662 644 663
rect 999 663 1000 664
rect 1004 663 1005 667
rect 999 662 1005 663
rect 1022 667 1028 668
rect 1022 663 1023 667
rect 1027 666 1028 667
rect 1206 667 1212 668
rect 1027 664 1045 666
rect 1027 663 1028 664
rect 1022 662 1028 663
rect 1206 663 1207 667
rect 1211 666 1212 667
rect 1506 667 1512 668
rect 1506 666 1507 667
rect 1211 664 1229 666
rect 1493 664 1507 666
rect 1211 663 1212 664
rect 1206 662 1212 663
rect 1506 663 1507 664
rect 1511 663 1512 667
rect 1506 662 1512 663
rect 594 658 600 659
rect 619 636 942 638
rect 594 635 600 636
rect 594 631 595 635
rect 599 634 600 635
rect 619 634 621 636
rect 599 632 621 634
rect 599 631 600 632
rect 594 630 600 631
rect 638 631 644 632
rect 638 630 639 631
rect 616 629 639 630
rect 110 625 116 626
rect 110 621 111 625
rect 115 621 116 625
rect 616 625 617 629
rect 621 628 639 629
rect 621 625 622 628
rect 638 627 639 628
rect 643 627 644 631
rect 638 626 644 627
rect 782 629 789 630
rect 616 624 622 625
rect 782 625 783 629
rect 788 625 789 629
rect 940 628 942 636
rect 999 631 1005 632
rect 959 629 965 630
rect 959 628 960 629
rect 940 626 960 628
rect 782 624 789 625
rect 959 625 960 626
rect 964 625 965 629
rect 999 627 1000 631
rect 1004 630 1005 631
rect 1004 628 1118 630
rect 1135 629 1141 630
rect 1135 628 1136 629
rect 1004 627 1005 628
rect 999 626 1005 627
rect 1116 626 1136 628
rect 959 624 965 625
rect 1135 625 1136 626
rect 1140 625 1141 629
rect 1135 624 1141 625
rect 1320 629 1332 630
rect 1320 625 1321 629
rect 1325 625 1327 629
rect 1331 625 1332 629
rect 1320 624 1332 625
rect 1494 629 1500 630
rect 1494 625 1495 629
rect 1499 628 1500 629
rect 1511 629 1517 630
rect 1511 628 1512 629
rect 1499 626 1512 628
rect 1499 625 1500 626
rect 1494 624 1500 625
rect 1511 625 1512 626
rect 1516 625 1517 629
rect 1511 624 1517 625
rect 1718 625 1724 626
rect 110 620 116 621
rect 510 623 516 624
rect 510 619 511 623
rect 515 619 516 623
rect 510 618 516 619
rect 678 623 684 624
rect 678 619 679 623
rect 683 619 684 623
rect 678 618 684 619
rect 854 623 860 624
rect 854 619 855 623
rect 859 619 860 623
rect 854 618 860 619
rect 1030 623 1036 624
rect 1030 619 1031 623
rect 1035 619 1036 623
rect 1030 618 1036 619
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1406 623 1412 624
rect 1406 619 1407 623
rect 1411 619 1412 623
rect 1718 621 1719 625
rect 1723 621 1724 625
rect 1718 620 1724 621
rect 1406 618 1412 619
rect 534 608 540 609
rect 110 607 116 608
rect 110 603 111 607
rect 115 603 116 607
rect 534 604 535 608
rect 539 604 540 608
rect 534 603 540 604
rect 702 608 708 609
rect 702 604 703 608
rect 707 604 708 608
rect 702 603 708 604
rect 878 608 884 609
rect 878 604 879 608
rect 883 604 884 608
rect 878 603 884 604
rect 1054 608 1060 609
rect 1054 604 1055 608
rect 1059 604 1060 608
rect 1054 603 1060 604
rect 1238 608 1244 609
rect 1238 604 1239 608
rect 1243 604 1244 608
rect 1238 603 1244 604
rect 1430 608 1436 609
rect 1430 604 1431 608
rect 1435 604 1436 608
rect 1430 603 1436 604
rect 1718 607 1724 608
rect 1718 603 1719 607
rect 1723 603 1724 607
rect 110 602 116 603
rect 1718 602 1724 603
rect 110 529 116 530
rect 1718 529 1724 530
rect 110 525 111 529
rect 115 525 116 529
rect 110 524 116 525
rect 166 528 172 529
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 550 528 556 529
rect 550 524 551 528
rect 555 524 556 528
rect 550 523 556 524
rect 742 528 748 529
rect 742 524 743 528
rect 747 524 748 528
rect 742 523 748 524
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 1126 528 1132 529
rect 1126 524 1127 528
rect 1131 524 1132 528
rect 1126 523 1132 524
rect 1326 528 1332 529
rect 1326 524 1327 528
rect 1331 524 1332 528
rect 1326 523 1332 524
rect 1526 528 1532 529
rect 1526 524 1527 528
rect 1531 524 1532 528
rect 1718 525 1719 529
rect 1723 525 1724 529
rect 1718 524 1724 525
rect 1526 523 1532 524
rect 142 513 148 514
rect 110 511 116 512
rect 110 507 111 511
rect 115 507 116 511
rect 142 509 143 513
rect 147 509 148 513
rect 142 508 148 509
rect 334 513 340 514
rect 334 509 335 513
rect 339 509 340 513
rect 334 508 340 509
rect 526 513 532 514
rect 526 509 527 513
rect 531 509 532 513
rect 526 508 532 509
rect 718 513 724 514
rect 718 509 719 513
rect 723 509 724 513
rect 718 508 724 509
rect 910 513 916 514
rect 910 509 911 513
rect 915 509 916 513
rect 910 508 916 509
rect 1102 513 1108 514
rect 1102 509 1103 513
rect 1107 509 1108 513
rect 1102 508 1108 509
rect 1302 513 1308 514
rect 1302 509 1303 513
rect 1307 509 1308 513
rect 1302 508 1308 509
rect 1502 513 1508 514
rect 1502 509 1503 513
rect 1507 509 1508 513
rect 1502 508 1508 509
rect 1718 511 1724 512
rect 110 506 116 507
rect 234 507 240 508
rect 234 503 235 507
rect 239 506 240 507
rect 247 507 253 508
rect 247 506 248 507
rect 239 504 248 506
rect 239 503 240 504
rect 234 502 240 503
rect 247 503 248 504
rect 252 503 253 507
rect 247 502 253 503
rect 295 507 301 508
rect 295 503 296 507
rect 300 506 301 507
rect 439 507 445 508
rect 439 506 440 507
rect 300 504 440 506
rect 300 503 301 504
rect 295 502 301 503
rect 439 503 440 504
rect 444 503 445 507
rect 439 502 445 503
rect 474 507 480 508
rect 474 503 475 507
rect 479 506 480 507
rect 631 507 637 508
rect 631 506 632 507
rect 479 504 632 506
rect 479 503 480 504
rect 474 502 480 503
rect 631 503 632 504
rect 636 503 637 507
rect 631 502 637 503
rect 710 507 716 508
rect 710 503 711 507
rect 715 506 716 507
rect 823 507 829 508
rect 823 506 824 507
rect 715 504 824 506
rect 715 503 716 504
rect 710 502 716 503
rect 823 503 824 504
rect 828 503 829 507
rect 823 502 829 503
rect 1015 507 1021 508
rect 1015 503 1016 507
rect 1020 506 1021 507
rect 1114 507 1120 508
rect 1114 506 1115 507
rect 1020 504 1115 506
rect 1020 503 1021 504
rect 1015 502 1021 503
rect 1114 503 1115 504
rect 1119 503 1120 507
rect 1114 502 1120 503
rect 1206 507 1213 508
rect 1206 503 1207 507
rect 1212 503 1213 507
rect 1206 502 1213 503
rect 1407 507 1413 508
rect 1407 503 1408 507
rect 1412 506 1413 507
rect 1514 507 1520 508
rect 1514 506 1515 507
rect 1412 504 1515 506
rect 1412 503 1413 504
rect 1407 502 1413 503
rect 1514 503 1515 504
rect 1519 503 1520 507
rect 1514 502 1520 503
rect 1570 507 1576 508
rect 1570 503 1571 507
rect 1575 506 1576 507
rect 1607 507 1613 508
rect 1607 506 1608 507
rect 1575 504 1608 506
rect 1575 503 1576 504
rect 1570 502 1576 503
rect 1607 503 1608 504
rect 1612 503 1613 507
rect 1718 507 1719 511
rect 1723 507 1724 511
rect 1718 506 1724 507
rect 1607 502 1613 503
rect 295 471 301 472
rect 295 470 296 471
rect 229 468 296 470
rect 295 467 296 468
rect 300 467 301 471
rect 474 471 480 472
rect 474 470 475 471
rect 421 468 475 470
rect 295 466 301 467
rect 474 467 475 468
rect 479 467 480 471
rect 710 471 716 472
rect 710 470 711 471
rect 613 468 711 470
rect 474 466 480 467
rect 710 467 711 468
rect 715 467 716 471
rect 710 466 716 467
rect 782 471 788 472
rect 782 467 783 471
rect 787 467 788 471
rect 1114 471 1120 472
rect 997 468 1102 470
rect 782 466 788 467
rect 1100 454 1102 468
rect 1114 467 1115 471
rect 1119 467 1120 471
rect 1494 471 1500 472
rect 1494 470 1495 471
rect 1389 468 1495 470
rect 1114 466 1120 467
rect 1494 467 1495 468
rect 1499 467 1500 471
rect 1494 466 1500 467
rect 1514 471 1520 472
rect 1514 467 1515 471
rect 1519 467 1520 471
rect 1514 466 1520 467
rect 1274 455 1280 456
rect 1274 454 1275 455
rect 1100 452 1275 454
rect 1274 451 1275 452
rect 1279 451 1280 455
rect 1274 450 1280 451
rect 234 423 240 424
rect 234 422 235 423
rect 221 420 235 422
rect 234 419 235 420
rect 239 419 240 423
rect 234 418 240 419
rect 242 423 248 424
rect 242 419 243 423
rect 247 422 248 423
rect 474 423 480 424
rect 247 420 365 422
rect 247 419 248 420
rect 242 418 248 419
rect 474 419 475 423
rect 479 422 480 423
rect 738 423 744 424
rect 479 420 629 422
rect 479 419 480 420
rect 474 418 480 419
rect 738 419 739 423
rect 743 422 744 423
rect 1570 423 1576 424
rect 1570 422 1571 423
rect 743 420 909 422
rect 1557 420 1571 422
rect 743 419 744 420
rect 738 418 744 419
rect 1266 419 1272 420
rect 1266 415 1267 419
rect 1271 415 1272 419
rect 1570 419 1571 420
rect 1575 419 1576 423
rect 1570 418 1576 419
rect 1266 414 1272 415
rect 240 385 248 386
rect 110 381 116 382
rect 110 377 111 381
rect 115 377 116 381
rect 240 381 241 385
rect 247 381 248 385
rect 240 380 248 381
rect 456 385 462 386
rect 456 381 457 385
rect 461 384 462 385
rect 474 385 480 386
rect 474 384 475 385
rect 461 382 475 384
rect 461 381 462 382
rect 456 380 462 381
rect 474 381 475 382
rect 479 381 480 385
rect 474 380 480 381
rect 720 385 726 386
rect 720 381 721 385
rect 725 384 726 385
rect 738 385 744 386
rect 738 384 739 385
rect 725 382 739 384
rect 725 381 726 382
rect 720 380 726 381
rect 738 381 739 382
rect 743 381 744 385
rect 738 380 744 381
rect 982 385 988 386
rect 982 381 983 385
rect 987 384 988 385
rect 999 385 1005 386
rect 999 384 1000 385
rect 987 382 1000 384
rect 987 381 988 382
rect 982 380 988 381
rect 999 381 1000 382
rect 1004 381 1005 385
rect 999 380 1005 381
rect 1274 385 1280 386
rect 1274 381 1275 385
rect 1279 384 1280 385
rect 1287 385 1293 386
rect 1287 384 1288 385
rect 1279 382 1288 384
rect 1279 381 1280 382
rect 1274 380 1280 381
rect 1287 381 1288 382
rect 1292 381 1293 385
rect 1287 380 1293 381
rect 1558 385 1564 386
rect 1558 381 1559 385
rect 1563 384 1564 385
rect 1575 385 1581 386
rect 1575 384 1576 385
rect 1563 382 1576 384
rect 1563 381 1564 382
rect 1558 380 1564 381
rect 1575 381 1576 382
rect 1580 381 1581 385
rect 1575 380 1581 381
rect 1718 381 1724 382
rect 110 376 116 377
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 350 379 356 380
rect 350 375 351 379
rect 355 375 356 379
rect 350 374 356 375
rect 614 379 620 380
rect 614 375 615 379
rect 619 375 620 379
rect 614 374 620 375
rect 894 379 900 380
rect 894 375 895 379
rect 899 375 900 379
rect 894 374 900 375
rect 1182 379 1188 380
rect 1182 375 1183 379
rect 1187 375 1188 379
rect 1182 374 1188 375
rect 1470 379 1476 380
rect 1470 375 1471 379
rect 1475 375 1476 379
rect 1718 377 1719 381
rect 1723 377 1724 381
rect 1718 376 1724 377
rect 1470 374 1476 375
rect 158 364 164 365
rect 110 363 116 364
rect 110 359 111 363
rect 115 359 116 363
rect 158 360 159 364
rect 163 360 164 364
rect 158 359 164 360
rect 374 364 380 365
rect 374 360 375 364
rect 379 360 380 364
rect 374 359 380 360
rect 638 364 644 365
rect 638 360 639 364
rect 643 360 644 364
rect 638 359 644 360
rect 918 364 924 365
rect 918 360 919 364
rect 923 360 924 364
rect 918 359 924 360
rect 1206 364 1212 365
rect 1206 360 1207 364
rect 1211 360 1212 364
rect 1206 359 1212 360
rect 1494 364 1500 365
rect 1494 360 1495 364
rect 1499 360 1500 364
rect 1494 359 1500 360
rect 1718 363 1724 364
rect 1718 359 1719 363
rect 1723 359 1724 363
rect 110 358 116 359
rect 1718 358 1724 359
rect 110 297 116 298
rect 1718 297 1724 298
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 222 296 228 297
rect 222 292 223 296
rect 227 292 228 296
rect 222 291 228 292
rect 454 296 460 297
rect 454 292 455 296
rect 459 292 460 296
rect 454 291 460 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 918 296 924 297
rect 918 292 919 296
rect 923 292 924 296
rect 918 291 924 292
rect 1150 296 1156 297
rect 1150 292 1151 296
rect 1155 292 1156 296
rect 1150 291 1156 292
rect 1382 296 1388 297
rect 1382 292 1383 296
rect 1387 292 1388 296
rect 1382 291 1388 292
rect 1598 296 1604 297
rect 1598 292 1599 296
rect 1603 292 1604 296
rect 1718 293 1719 297
rect 1723 293 1724 297
rect 1718 292 1724 293
rect 1598 291 1604 292
rect 198 281 204 282
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 198 277 199 281
rect 203 277 204 281
rect 198 276 204 277
rect 430 281 436 282
rect 430 277 431 281
rect 435 277 436 281
rect 430 276 436 277
rect 662 281 668 282
rect 662 277 663 281
rect 667 277 668 281
rect 662 276 668 277
rect 894 281 900 282
rect 894 277 895 281
rect 899 277 900 281
rect 894 276 900 277
rect 1126 281 1132 282
rect 1126 277 1127 281
rect 1131 277 1132 281
rect 1126 276 1132 277
rect 1358 281 1364 282
rect 1358 277 1359 281
rect 1363 277 1364 281
rect 1358 276 1364 277
rect 1574 281 1580 282
rect 1574 277 1575 281
rect 1579 277 1580 281
rect 1574 276 1580 277
rect 1718 279 1724 280
rect 110 274 116 275
rect 302 275 309 276
rect 302 271 303 275
rect 308 271 309 275
rect 302 270 309 271
rect 374 275 380 276
rect 374 271 375 275
rect 379 274 380 275
rect 535 275 541 276
rect 535 274 536 275
rect 379 272 536 274
rect 379 271 380 272
rect 374 270 380 271
rect 535 271 536 272
rect 540 271 541 275
rect 535 270 541 271
rect 546 275 552 276
rect 546 271 547 275
rect 551 274 552 275
rect 767 275 773 276
rect 767 274 768 275
rect 551 272 768 274
rect 551 271 552 272
rect 546 270 552 271
rect 767 271 768 272
rect 772 271 773 275
rect 767 270 773 271
rect 999 275 1005 276
rect 999 271 1000 275
rect 1004 274 1005 275
rect 1138 275 1144 276
rect 1138 274 1139 275
rect 1004 272 1139 274
rect 1004 271 1005 272
rect 999 270 1005 271
rect 1138 271 1139 272
rect 1143 271 1144 275
rect 1138 270 1144 271
rect 1231 275 1237 276
rect 1231 271 1232 275
rect 1236 274 1237 275
rect 1266 275 1272 276
rect 1266 274 1267 275
rect 1236 272 1267 274
rect 1236 271 1237 272
rect 1231 270 1237 271
rect 1266 271 1267 272
rect 1271 271 1272 275
rect 1266 270 1272 271
rect 1463 275 1469 276
rect 1463 271 1464 275
rect 1468 274 1469 275
rect 1586 275 1592 276
rect 1586 274 1587 275
rect 1468 272 1587 274
rect 1468 271 1469 272
rect 1463 270 1469 271
rect 1586 271 1587 272
rect 1591 271 1592 275
rect 1586 270 1592 271
rect 1674 275 1685 276
rect 1674 271 1675 275
rect 1679 271 1680 275
rect 1684 271 1685 275
rect 1718 275 1719 279
rect 1723 275 1724 279
rect 1718 274 1724 275
rect 1674 270 1685 271
rect 982 255 988 256
rect 982 254 983 255
rect 840 252 983 254
rect 374 239 380 240
rect 374 238 375 239
rect 285 236 375 238
rect 374 235 375 236
rect 379 235 380 239
rect 546 239 552 240
rect 546 238 547 239
rect 517 236 547 238
rect 374 234 380 235
rect 546 235 547 236
rect 551 235 552 239
rect 840 238 842 252
rect 982 251 983 252
rect 987 251 988 255
rect 982 250 988 251
rect 1138 239 1144 240
rect 749 236 842 238
rect 981 236 1126 238
rect 546 234 552 235
rect 1124 222 1126 236
rect 1138 235 1139 239
rect 1143 235 1144 239
rect 1558 239 1564 240
rect 1558 238 1559 239
rect 1445 236 1559 238
rect 1138 234 1144 235
rect 1558 235 1559 236
rect 1563 235 1564 239
rect 1558 234 1564 235
rect 1586 239 1592 240
rect 1586 235 1587 239
rect 1591 235 1592 239
rect 1586 234 1592 235
rect 1326 223 1332 224
rect 1326 222 1327 223
rect 1124 220 1327 222
rect 1326 219 1327 220
rect 1331 219 1332 223
rect 1326 218 1332 219
rect 302 195 308 196
rect 302 191 303 195
rect 307 194 308 195
rect 422 195 428 196
rect 307 192 325 194
rect 307 191 308 192
rect 302 190 308 191
rect 422 191 423 195
rect 427 194 428 195
rect 554 195 560 196
rect 427 192 461 194
rect 427 191 428 192
rect 422 190 428 191
rect 554 191 555 195
rect 559 194 560 195
rect 714 195 720 196
rect 559 192 605 194
rect 559 191 560 192
rect 554 190 560 191
rect 714 191 715 195
rect 719 194 720 195
rect 866 195 872 196
rect 719 192 757 194
rect 719 191 720 192
rect 714 190 720 191
rect 866 191 867 195
rect 871 194 872 195
rect 1010 195 1016 196
rect 871 192 917 194
rect 871 191 872 192
rect 866 190 872 191
rect 1010 191 1011 195
rect 1015 194 1016 195
rect 1178 195 1184 196
rect 1015 192 1085 194
rect 1015 191 1016 192
rect 1010 190 1016 191
rect 1178 191 1179 195
rect 1183 194 1184 195
rect 1674 195 1680 196
rect 1674 194 1675 195
rect 1183 192 1253 194
rect 1661 192 1675 194
rect 1183 191 1184 192
rect 1178 190 1184 191
rect 1498 191 1504 192
rect 1498 187 1499 191
rect 1503 187 1504 191
rect 1674 191 1675 192
rect 1679 191 1680 195
rect 1674 190 1680 191
rect 1498 186 1504 187
rect 1498 159 1504 160
rect 416 157 428 158
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 416 153 417 157
rect 421 153 423 157
rect 427 153 428 157
rect 416 152 428 153
rect 552 157 560 158
rect 552 153 553 157
rect 559 153 560 157
rect 552 152 560 153
rect 696 157 702 158
rect 696 153 697 157
rect 701 156 702 157
rect 714 157 720 158
rect 714 156 715 157
rect 701 154 715 156
rect 701 153 702 154
rect 696 152 702 153
rect 714 153 715 154
rect 719 153 720 157
rect 714 152 720 153
rect 848 157 854 158
rect 848 153 849 157
rect 853 156 854 157
rect 866 157 872 158
rect 866 156 867 157
rect 853 154 867 156
rect 853 153 854 154
rect 848 152 854 153
rect 866 153 867 154
rect 871 153 872 157
rect 866 152 872 153
rect 1008 157 1016 158
rect 1008 153 1009 157
rect 1015 153 1016 157
rect 1008 152 1016 153
rect 1176 157 1184 158
rect 1176 153 1177 157
rect 1183 153 1184 157
rect 1176 152 1184 153
rect 1326 157 1332 158
rect 1326 153 1327 157
rect 1331 156 1332 157
rect 1343 157 1349 158
rect 1343 156 1344 157
rect 1331 154 1344 156
rect 1331 153 1332 154
rect 1326 152 1332 153
rect 1343 153 1344 154
rect 1348 153 1349 157
rect 1498 155 1499 159
rect 1503 158 1504 159
rect 1503 156 1662 158
rect 1679 157 1685 158
rect 1679 156 1680 157
rect 1503 155 1504 156
rect 1498 154 1504 155
rect 1660 154 1680 156
rect 1343 152 1349 153
rect 1679 153 1680 154
rect 1684 153 1685 157
rect 1679 152 1685 153
rect 1718 153 1724 154
rect 110 148 116 149
rect 310 151 316 152
rect 310 147 311 151
rect 315 147 316 151
rect 310 146 316 147
rect 446 151 452 152
rect 446 147 447 151
rect 451 147 452 151
rect 446 146 452 147
rect 590 151 596 152
rect 590 147 591 151
rect 595 147 596 151
rect 590 146 596 147
rect 742 151 748 152
rect 742 147 743 151
rect 747 147 748 151
rect 742 146 748 147
rect 902 151 908 152
rect 902 147 903 151
rect 907 147 908 151
rect 902 146 908 147
rect 1070 151 1076 152
rect 1070 147 1071 151
rect 1075 147 1076 151
rect 1070 146 1076 147
rect 1238 151 1244 152
rect 1238 147 1239 151
rect 1243 147 1244 151
rect 1238 146 1244 147
rect 1414 151 1420 152
rect 1414 147 1415 151
rect 1419 147 1420 151
rect 1414 146 1420 147
rect 1574 151 1580 152
rect 1574 147 1575 151
rect 1579 147 1580 151
rect 1718 149 1719 153
rect 1723 149 1724 153
rect 1718 148 1724 149
rect 1574 146 1580 147
rect 334 136 340 137
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 334 132 335 136
rect 339 132 340 136
rect 334 131 340 132
rect 470 136 476 137
rect 470 132 471 136
rect 475 132 476 136
rect 470 131 476 132
rect 614 136 620 137
rect 614 132 615 136
rect 619 132 620 136
rect 614 131 620 132
rect 766 136 772 137
rect 766 132 767 136
rect 771 132 772 136
rect 766 131 772 132
rect 926 136 932 137
rect 926 132 927 136
rect 931 132 932 136
rect 926 131 932 132
rect 1094 136 1100 137
rect 1094 132 1095 136
rect 1099 132 1100 136
rect 1094 131 1100 132
rect 1262 136 1268 137
rect 1262 132 1263 136
rect 1267 132 1268 136
rect 1262 131 1268 132
rect 1438 136 1444 137
rect 1438 132 1439 136
rect 1443 132 1444 136
rect 1438 131 1444 132
rect 1598 136 1604 137
rect 1598 132 1599 136
rect 1603 132 1604 136
rect 1598 131 1604 132
rect 1718 135 1724 136
rect 1718 131 1719 135
rect 1723 131 1724 135
rect 110 130 116 131
rect 1718 130 1724 131
<< m3c >>
rect 243 1763 247 1767
rect 379 1763 383 1767
rect 515 1763 519 1767
rect 651 1763 655 1767
rect 111 1721 115 1725
rect 243 1725 245 1729
rect 245 1725 247 1729
rect 379 1725 381 1729
rect 381 1725 383 1729
rect 515 1725 517 1729
rect 517 1725 519 1729
rect 651 1725 653 1729
rect 653 1725 655 1729
rect 767 1725 771 1729
rect 135 1719 139 1723
rect 271 1719 275 1723
rect 407 1719 411 1723
rect 543 1719 547 1723
rect 679 1719 683 1723
rect 1719 1721 1723 1725
rect 111 1703 115 1707
rect 159 1704 163 1708
rect 295 1704 299 1708
rect 431 1704 435 1708
rect 567 1704 571 1708
rect 703 1704 707 1708
rect 1719 1703 1723 1707
rect 111 1629 115 1633
rect 247 1628 251 1632
rect 383 1628 387 1632
rect 519 1628 523 1632
rect 655 1628 659 1632
rect 791 1628 795 1632
rect 1719 1629 1723 1633
rect 111 1611 115 1615
rect 223 1613 227 1617
rect 359 1613 363 1617
rect 495 1613 499 1617
rect 631 1613 635 1617
rect 767 1613 771 1617
rect 371 1607 375 1611
rect 507 1607 511 1611
rect 643 1607 647 1611
rect 779 1607 783 1611
rect 587 1599 591 1603
rect 1719 1611 1723 1615
rect 307 1571 311 1575
rect 371 1571 375 1575
rect 507 1571 511 1575
rect 643 1571 647 1575
rect 779 1571 783 1575
rect 587 1535 591 1539
rect 599 1535 603 1539
rect 731 1535 735 1539
rect 875 1535 879 1539
rect 1003 1535 1007 1539
rect 1275 1535 1279 1539
rect 1547 1535 1551 1539
rect 1287 1527 1291 1531
rect 111 1493 115 1497
rect 599 1497 603 1501
rect 731 1497 733 1501
rect 733 1497 735 1501
rect 875 1497 879 1501
rect 1003 1497 1005 1501
rect 1005 1497 1007 1501
rect 1119 1497 1123 1501
rect 1275 1497 1277 1501
rect 1277 1497 1279 1501
rect 1547 1497 1549 1501
rect 1549 1497 1551 1501
rect 487 1491 491 1495
rect 623 1491 627 1495
rect 759 1491 763 1495
rect 895 1491 899 1495
rect 1031 1491 1035 1495
rect 1167 1491 1171 1495
rect 1303 1491 1307 1495
rect 1439 1491 1443 1495
rect 1575 1491 1579 1495
rect 1719 1493 1723 1497
rect 111 1475 115 1479
rect 511 1476 515 1480
rect 647 1476 651 1480
rect 783 1476 787 1480
rect 919 1476 923 1480
rect 1055 1476 1059 1480
rect 1191 1476 1195 1480
rect 1327 1476 1331 1480
rect 1463 1476 1467 1480
rect 1599 1476 1603 1480
rect 1719 1475 1723 1479
rect 111 1401 115 1405
rect 743 1400 747 1404
rect 887 1400 891 1404
rect 1031 1400 1035 1404
rect 1175 1400 1179 1404
rect 1319 1400 1323 1404
rect 1463 1400 1467 1404
rect 1599 1400 1603 1404
rect 1719 1401 1723 1405
rect 111 1383 115 1387
rect 719 1385 723 1389
rect 863 1385 867 1389
rect 1007 1385 1011 1389
rect 1151 1385 1155 1389
rect 1295 1385 1299 1389
rect 1439 1385 1443 1389
rect 1575 1385 1579 1389
rect 875 1379 879 1383
rect 1019 1379 1023 1383
rect 1163 1379 1167 1383
rect 1259 1379 1260 1383
rect 1260 1379 1263 1383
rect 1287 1379 1291 1383
rect 1587 1379 1591 1383
rect 1675 1379 1679 1383
rect 1719 1383 1723 1387
rect 1119 1359 1123 1363
rect 875 1343 879 1347
rect 1019 1343 1023 1347
rect 1163 1343 1167 1347
rect 1379 1343 1383 1347
rect 1587 1343 1591 1347
rect 359 1311 363 1315
rect 531 1311 535 1315
rect 887 1311 891 1315
rect 1191 1311 1195 1315
rect 1259 1311 1263 1315
rect 1675 1311 1679 1315
rect 111 1269 115 1273
rect 271 1273 275 1277
rect 359 1275 363 1279
rect 531 1275 535 1279
rect 887 1275 891 1279
rect 1191 1275 1195 1279
rect 1667 1273 1671 1277
rect 183 1267 187 1271
rect 415 1267 419 1271
rect 679 1267 683 1271
rect 975 1267 979 1271
rect 1287 1267 1291 1271
rect 1575 1267 1579 1271
rect 1719 1269 1723 1273
rect 111 1251 115 1255
rect 207 1252 211 1256
rect 439 1252 443 1256
rect 703 1252 707 1256
rect 999 1252 1003 1256
rect 1311 1252 1315 1256
rect 1599 1252 1603 1256
rect 1719 1251 1723 1255
rect 111 1189 115 1193
rect 159 1188 163 1192
rect 335 1188 339 1192
rect 559 1188 563 1192
rect 799 1188 803 1192
rect 1063 1188 1067 1192
rect 1335 1188 1339 1192
rect 1599 1188 1603 1192
rect 1719 1189 1723 1193
rect 111 1171 115 1175
rect 135 1173 139 1177
rect 311 1173 315 1177
rect 535 1173 539 1177
rect 775 1173 779 1177
rect 1039 1173 1043 1177
rect 1311 1173 1315 1177
rect 1575 1173 1579 1177
rect 323 1167 327 1171
rect 547 1167 551 1171
rect 787 1167 791 1171
rect 1051 1167 1055 1171
rect 1091 1167 1095 1171
rect 1379 1167 1383 1171
rect 1659 1167 1663 1171
rect 1719 1171 1723 1175
rect 271 1131 275 1135
rect 323 1131 327 1135
rect 547 1131 551 1135
rect 787 1131 791 1135
rect 1051 1131 1055 1135
rect 1375 1131 1379 1135
rect 1667 1131 1671 1135
rect 1091 1103 1095 1107
rect 331 1091 335 1095
rect 587 1091 591 1095
rect 843 1091 847 1095
rect 1455 1091 1459 1095
rect 1659 1091 1663 1095
rect 111 1049 115 1053
rect 331 1053 333 1057
rect 333 1053 335 1057
rect 587 1053 591 1057
rect 843 1053 847 1057
rect 1095 1053 1096 1057
rect 1096 1053 1099 1057
rect 1375 1053 1376 1057
rect 1376 1053 1379 1057
rect 1647 1053 1651 1057
rect 223 1047 227 1051
rect 463 1047 467 1051
rect 719 1047 723 1051
rect 991 1047 995 1051
rect 1271 1047 1275 1051
rect 1559 1047 1563 1051
rect 1719 1049 1723 1053
rect 111 1031 115 1035
rect 247 1032 251 1036
rect 487 1032 491 1036
rect 743 1032 747 1036
rect 1015 1032 1019 1036
rect 1295 1032 1299 1036
rect 1583 1032 1587 1036
rect 1719 1031 1723 1035
rect 559 987 563 991
rect 1095 987 1099 991
rect 111 973 115 977
rect 463 972 467 976
rect 647 972 651 976
rect 855 972 859 976
rect 1079 972 1083 976
rect 1311 972 1315 976
rect 1543 972 1547 976
rect 1719 973 1723 977
rect 111 955 115 959
rect 439 957 443 961
rect 623 957 627 961
rect 831 957 835 961
rect 1055 957 1059 961
rect 1287 957 1291 961
rect 1519 957 1523 961
rect 635 951 639 955
rect 843 951 847 955
rect 1067 951 1071 955
rect 1299 951 1303 955
rect 787 943 791 947
rect 1603 951 1607 955
rect 1719 955 1723 959
rect 559 915 563 919
rect 635 915 639 919
rect 843 915 847 919
rect 1067 915 1071 919
rect 1299 915 1303 919
rect 1647 915 1651 919
rect 787 883 791 887
rect 795 883 799 887
rect 931 883 935 887
rect 1067 883 1071 887
rect 1203 883 1207 887
rect 1451 879 1455 883
rect 1603 883 1607 887
rect 111 841 115 845
rect 795 845 797 849
rect 797 845 799 849
rect 931 845 933 849
rect 933 845 935 849
rect 1067 845 1069 849
rect 1069 845 1071 849
rect 1203 845 1205 849
rect 1205 845 1207 849
rect 1319 845 1323 849
rect 1459 845 1463 849
rect 1591 845 1595 849
rect 687 839 691 843
rect 823 839 827 843
rect 959 839 963 843
rect 1095 839 1099 843
rect 1231 839 1235 843
rect 1367 839 1371 843
rect 1503 839 1507 843
rect 1719 841 1723 845
rect 111 823 115 827
rect 711 824 715 828
rect 847 824 851 828
rect 983 824 987 828
rect 1119 824 1123 828
rect 1255 824 1259 828
rect 1391 824 1395 828
rect 1527 824 1531 828
rect 1719 823 1723 827
rect 111 753 115 757
rect 815 752 819 756
rect 951 752 955 756
rect 1087 752 1091 756
rect 1223 752 1227 756
rect 1359 752 1363 756
rect 1495 752 1499 756
rect 1719 753 1723 757
rect 111 735 115 739
rect 791 737 795 741
rect 927 737 931 741
rect 1063 737 1067 741
rect 1199 737 1203 741
rect 1335 737 1339 741
rect 1471 737 1475 741
rect 939 731 943 735
rect 1023 731 1027 735
rect 1099 731 1103 735
rect 1179 731 1183 735
rect 1451 731 1455 735
rect 1507 731 1511 735
rect 1719 735 1723 739
rect 875 695 879 699
rect 939 695 943 699
rect 1179 695 1183 699
rect 1319 695 1323 699
rect 1327 695 1331 699
rect 1591 695 1595 699
rect 595 659 599 663
rect 639 663 643 667
rect 1023 663 1027 667
rect 1207 663 1211 667
rect 1507 663 1511 667
rect 595 631 599 635
rect 111 621 115 625
rect 639 627 643 631
rect 783 625 784 629
rect 784 625 787 629
rect 1327 625 1331 629
rect 1495 625 1499 629
rect 511 619 515 623
rect 679 619 683 623
rect 855 619 859 623
rect 1031 619 1035 623
rect 1215 619 1219 623
rect 1407 619 1411 623
rect 1719 621 1723 625
rect 111 603 115 607
rect 535 604 539 608
rect 703 604 707 608
rect 879 604 883 608
rect 1055 604 1059 608
rect 1239 604 1243 608
rect 1431 604 1435 608
rect 1719 603 1723 607
rect 111 525 115 529
rect 167 524 171 528
rect 359 524 363 528
rect 551 524 555 528
rect 743 524 747 528
rect 935 524 939 528
rect 1127 524 1131 528
rect 1327 524 1331 528
rect 1527 524 1531 528
rect 1719 525 1723 529
rect 111 507 115 511
rect 143 509 147 513
rect 335 509 339 513
rect 527 509 531 513
rect 719 509 723 513
rect 911 509 915 513
rect 1103 509 1107 513
rect 1303 509 1307 513
rect 1503 509 1507 513
rect 235 503 239 507
rect 475 503 479 507
rect 711 503 715 507
rect 1115 503 1119 507
rect 1207 503 1208 507
rect 1208 503 1211 507
rect 1515 503 1519 507
rect 1571 503 1575 507
rect 1719 507 1723 511
rect 475 467 479 471
rect 711 467 715 471
rect 783 467 787 471
rect 1115 467 1119 471
rect 1495 467 1499 471
rect 1515 467 1519 471
rect 1275 451 1279 455
rect 235 419 239 423
rect 243 419 247 423
rect 475 419 479 423
rect 739 419 743 423
rect 1267 415 1271 419
rect 1571 419 1575 423
rect 111 377 115 381
rect 243 381 245 385
rect 245 381 247 385
rect 475 381 479 385
rect 739 381 743 385
rect 983 381 987 385
rect 1275 381 1279 385
rect 1559 381 1563 385
rect 135 375 139 379
rect 351 375 355 379
rect 615 375 619 379
rect 895 375 899 379
rect 1183 375 1187 379
rect 1471 375 1475 379
rect 1719 377 1723 381
rect 111 359 115 363
rect 159 360 163 364
rect 375 360 379 364
rect 639 360 643 364
rect 919 360 923 364
rect 1207 360 1211 364
rect 1495 360 1499 364
rect 1719 359 1723 363
rect 111 293 115 297
rect 223 292 227 296
rect 455 292 459 296
rect 687 292 691 296
rect 919 292 923 296
rect 1151 292 1155 296
rect 1383 292 1387 296
rect 1599 292 1603 296
rect 1719 293 1723 297
rect 111 275 115 279
rect 199 277 203 281
rect 431 277 435 281
rect 663 277 667 281
rect 895 277 899 281
rect 1127 277 1131 281
rect 1359 277 1363 281
rect 1575 277 1579 281
rect 303 271 304 275
rect 304 271 307 275
rect 375 271 379 275
rect 547 271 551 275
rect 1139 271 1143 275
rect 1267 271 1271 275
rect 1587 271 1591 275
rect 1675 271 1679 275
rect 1719 275 1723 279
rect 375 235 379 239
rect 547 235 551 239
rect 983 251 987 255
rect 1139 235 1143 239
rect 1559 235 1563 239
rect 1587 235 1591 239
rect 1327 219 1331 223
rect 303 191 307 195
rect 423 191 427 195
rect 555 191 559 195
rect 715 191 719 195
rect 867 191 871 195
rect 1011 191 1015 195
rect 1179 191 1183 195
rect 1499 187 1503 191
rect 1675 191 1679 195
rect 111 149 115 153
rect 423 153 427 157
rect 555 153 557 157
rect 557 153 559 157
rect 715 153 719 157
rect 867 153 871 157
rect 1011 153 1013 157
rect 1013 153 1015 157
rect 1179 153 1181 157
rect 1181 153 1183 157
rect 1327 153 1331 157
rect 1499 155 1503 159
rect 311 147 315 151
rect 447 147 451 151
rect 591 147 595 151
rect 743 147 747 151
rect 903 147 907 151
rect 1071 147 1075 151
rect 1239 147 1243 151
rect 1415 147 1419 151
rect 1575 147 1579 151
rect 1719 149 1723 153
rect 111 131 115 135
rect 335 132 339 136
rect 471 132 475 136
rect 615 132 619 136
rect 767 132 771 136
rect 927 132 931 136
rect 1095 132 1099 136
rect 1263 132 1267 136
rect 1439 132 1443 136
rect 1599 132 1603 136
rect 1719 131 1723 135
<< m3 >>
rect 111 1778 115 1779
rect 111 1773 115 1774
rect 135 1778 139 1779
rect 135 1773 139 1774
rect 271 1778 275 1779
rect 271 1773 275 1774
rect 407 1778 411 1779
rect 407 1773 411 1774
rect 543 1778 547 1779
rect 543 1773 547 1774
rect 679 1778 683 1779
rect 679 1773 683 1774
rect 1719 1778 1723 1779
rect 1719 1773 1723 1774
rect 112 1726 114 1773
rect 110 1725 116 1726
rect 110 1721 111 1725
rect 115 1721 116 1725
rect 136 1724 138 1773
rect 242 1767 248 1768
rect 242 1763 243 1767
rect 247 1763 248 1767
rect 242 1762 248 1763
rect 244 1730 246 1762
rect 242 1729 248 1730
rect 242 1725 243 1729
rect 247 1725 248 1729
rect 242 1724 248 1725
rect 272 1724 274 1773
rect 378 1767 384 1768
rect 378 1763 379 1767
rect 383 1763 384 1767
rect 378 1762 384 1763
rect 380 1730 382 1762
rect 378 1729 384 1730
rect 378 1725 379 1729
rect 383 1725 384 1729
rect 378 1724 384 1725
rect 408 1724 410 1773
rect 514 1767 520 1768
rect 514 1763 515 1767
rect 519 1763 520 1767
rect 514 1762 520 1763
rect 516 1730 518 1762
rect 514 1729 520 1730
rect 514 1725 515 1729
rect 519 1725 520 1729
rect 514 1724 520 1725
rect 544 1724 546 1773
rect 650 1767 656 1768
rect 650 1763 651 1767
rect 655 1763 656 1767
rect 650 1762 656 1763
rect 652 1730 654 1762
rect 650 1729 656 1730
rect 650 1725 651 1729
rect 655 1725 656 1729
rect 650 1724 656 1725
rect 680 1724 682 1773
rect 766 1729 772 1730
rect 766 1725 767 1729
rect 771 1725 772 1729
rect 1720 1726 1722 1773
rect 766 1724 772 1725
rect 1718 1725 1724 1726
rect 110 1720 116 1721
rect 134 1723 140 1724
rect 134 1719 135 1723
rect 139 1719 140 1723
rect 134 1718 140 1719
rect 270 1723 276 1724
rect 270 1719 271 1723
rect 275 1719 276 1723
rect 270 1718 276 1719
rect 406 1723 412 1724
rect 406 1719 407 1723
rect 411 1719 412 1723
rect 406 1718 412 1719
rect 542 1723 548 1724
rect 542 1719 543 1723
rect 547 1719 548 1723
rect 542 1718 548 1719
rect 678 1723 684 1724
rect 678 1719 679 1723
rect 683 1719 684 1723
rect 678 1718 684 1719
rect 158 1708 164 1709
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 158 1704 159 1708
rect 163 1704 164 1708
rect 158 1703 164 1704
rect 294 1708 300 1709
rect 294 1704 295 1708
rect 299 1704 300 1708
rect 294 1703 300 1704
rect 430 1708 436 1709
rect 430 1704 431 1708
rect 435 1704 436 1708
rect 430 1703 436 1704
rect 566 1708 572 1709
rect 566 1704 567 1708
rect 571 1704 572 1708
rect 566 1703 572 1704
rect 702 1708 708 1709
rect 702 1704 703 1708
rect 707 1704 708 1708
rect 702 1703 708 1704
rect 110 1702 116 1703
rect 112 1663 114 1702
rect 160 1663 162 1703
rect 296 1663 298 1703
rect 432 1663 434 1703
rect 568 1663 570 1703
rect 704 1663 706 1703
rect 111 1662 115 1663
rect 111 1657 115 1658
rect 159 1662 163 1663
rect 159 1657 163 1658
rect 247 1662 251 1663
rect 247 1657 251 1658
rect 295 1662 299 1663
rect 295 1657 299 1658
rect 383 1662 387 1663
rect 383 1657 387 1658
rect 431 1662 435 1663
rect 431 1657 435 1658
rect 519 1662 523 1663
rect 519 1657 523 1658
rect 567 1662 571 1663
rect 567 1657 571 1658
rect 655 1662 659 1663
rect 655 1657 659 1658
rect 703 1662 707 1663
rect 703 1657 707 1658
rect 112 1634 114 1657
rect 110 1633 116 1634
rect 248 1633 250 1657
rect 384 1633 386 1657
rect 520 1633 522 1657
rect 656 1633 658 1657
rect 110 1629 111 1633
rect 115 1629 116 1633
rect 110 1628 116 1629
rect 246 1632 252 1633
rect 246 1628 247 1632
rect 251 1628 252 1632
rect 382 1632 388 1633
rect 246 1627 252 1628
rect 307 1628 311 1629
rect 382 1628 383 1632
rect 387 1628 388 1632
rect 382 1627 388 1628
rect 518 1632 524 1633
rect 518 1628 519 1632
rect 523 1628 524 1632
rect 518 1627 524 1628
rect 654 1632 660 1633
rect 654 1628 655 1632
rect 659 1628 660 1632
rect 768 1629 770 1724
rect 1718 1721 1719 1725
rect 1723 1721 1724 1725
rect 1718 1720 1724 1721
rect 1718 1707 1724 1708
rect 1718 1703 1719 1707
rect 1723 1703 1724 1707
rect 1718 1702 1724 1703
rect 1720 1663 1722 1702
rect 791 1662 795 1663
rect 791 1657 795 1658
rect 1719 1662 1723 1663
rect 1719 1657 1723 1658
rect 792 1633 794 1657
rect 1720 1634 1722 1657
rect 1718 1633 1724 1634
rect 790 1632 796 1633
rect 654 1627 660 1628
rect 767 1628 771 1629
rect 307 1623 311 1624
rect 790 1628 791 1632
rect 795 1628 796 1632
rect 1718 1629 1719 1633
rect 1723 1629 1724 1633
rect 1718 1628 1724 1629
rect 790 1627 796 1628
rect 767 1623 771 1624
rect 222 1617 228 1618
rect 110 1615 116 1616
rect 110 1611 111 1615
rect 115 1611 116 1615
rect 222 1613 223 1617
rect 227 1613 228 1617
rect 222 1612 228 1613
rect 110 1610 116 1611
rect 112 1551 114 1610
rect 224 1551 226 1612
rect 308 1576 310 1623
rect 358 1617 364 1618
rect 358 1613 359 1617
rect 363 1613 364 1617
rect 358 1612 364 1613
rect 494 1617 500 1618
rect 494 1613 495 1617
rect 499 1613 500 1617
rect 494 1612 500 1613
rect 630 1617 636 1618
rect 630 1613 631 1617
rect 635 1613 636 1617
rect 630 1612 636 1613
rect 766 1617 772 1618
rect 766 1613 767 1617
rect 771 1613 772 1617
rect 766 1612 772 1613
rect 1718 1615 1724 1616
rect 306 1575 312 1576
rect 306 1571 307 1575
rect 311 1571 312 1575
rect 306 1570 312 1571
rect 360 1551 362 1612
rect 370 1611 376 1612
rect 370 1607 371 1611
rect 375 1607 376 1611
rect 370 1606 376 1607
rect 372 1576 374 1606
rect 370 1575 376 1576
rect 370 1571 371 1575
rect 375 1571 376 1575
rect 370 1570 376 1571
rect 496 1551 498 1612
rect 506 1611 512 1612
rect 506 1607 507 1611
rect 511 1607 512 1611
rect 506 1606 512 1607
rect 508 1576 510 1606
rect 586 1603 592 1604
rect 586 1599 587 1603
rect 591 1599 592 1603
rect 586 1598 592 1599
rect 506 1575 512 1576
rect 506 1571 507 1575
rect 511 1571 512 1575
rect 506 1570 512 1571
rect 111 1550 115 1551
rect 111 1545 115 1546
rect 223 1550 227 1551
rect 223 1545 227 1546
rect 359 1550 363 1551
rect 359 1545 363 1546
rect 487 1550 491 1551
rect 487 1545 491 1546
rect 495 1550 499 1551
rect 495 1545 499 1546
rect 112 1498 114 1545
rect 110 1497 116 1498
rect 110 1493 111 1497
rect 115 1493 116 1497
rect 488 1496 490 1545
rect 588 1540 590 1598
rect 632 1551 634 1612
rect 642 1611 648 1612
rect 642 1607 643 1611
rect 647 1607 648 1611
rect 642 1606 648 1607
rect 644 1576 646 1606
rect 642 1575 648 1576
rect 642 1571 643 1575
rect 647 1571 648 1575
rect 642 1570 648 1571
rect 768 1551 770 1612
rect 778 1611 784 1612
rect 778 1607 779 1611
rect 783 1607 784 1611
rect 1718 1611 1719 1615
rect 1723 1611 1724 1615
rect 1718 1610 1724 1611
rect 778 1606 784 1607
rect 780 1576 782 1606
rect 778 1575 784 1576
rect 778 1571 779 1575
rect 783 1571 784 1575
rect 778 1570 784 1571
rect 1720 1551 1722 1610
rect 623 1550 627 1551
rect 623 1545 627 1546
rect 631 1550 635 1551
rect 631 1545 635 1546
rect 759 1550 763 1551
rect 759 1545 763 1546
rect 767 1550 771 1551
rect 767 1545 771 1546
rect 895 1550 899 1551
rect 895 1545 899 1546
rect 1031 1550 1035 1551
rect 1031 1545 1035 1546
rect 1167 1550 1171 1551
rect 1167 1545 1171 1546
rect 1303 1550 1307 1551
rect 1303 1545 1307 1546
rect 1439 1550 1443 1551
rect 1439 1545 1443 1546
rect 1575 1550 1579 1551
rect 1575 1545 1579 1546
rect 1719 1550 1723 1551
rect 1719 1545 1723 1546
rect 586 1539 592 1540
rect 586 1535 587 1539
rect 591 1535 592 1539
rect 586 1534 592 1535
rect 598 1539 604 1540
rect 598 1535 599 1539
rect 603 1535 604 1539
rect 598 1534 604 1535
rect 600 1502 602 1534
rect 598 1501 604 1502
rect 598 1497 599 1501
rect 603 1497 604 1501
rect 598 1496 604 1497
rect 624 1496 626 1545
rect 730 1539 736 1540
rect 730 1535 731 1539
rect 735 1535 736 1539
rect 730 1534 736 1535
rect 732 1502 734 1534
rect 730 1501 736 1502
rect 730 1497 731 1501
rect 735 1497 736 1501
rect 730 1496 736 1497
rect 760 1496 762 1545
rect 874 1539 880 1540
rect 874 1535 875 1539
rect 879 1535 880 1539
rect 874 1534 880 1535
rect 876 1502 878 1534
rect 874 1501 880 1502
rect 874 1497 875 1501
rect 879 1497 880 1501
rect 874 1496 880 1497
rect 896 1496 898 1545
rect 1002 1539 1008 1540
rect 1002 1535 1003 1539
rect 1007 1535 1008 1539
rect 1002 1534 1008 1535
rect 1004 1502 1006 1534
rect 1002 1501 1008 1502
rect 1002 1497 1003 1501
rect 1007 1497 1008 1501
rect 1002 1496 1008 1497
rect 1032 1496 1034 1545
rect 1118 1501 1124 1502
rect 1118 1497 1119 1501
rect 1123 1497 1124 1501
rect 1118 1496 1124 1497
rect 1168 1496 1170 1545
rect 1274 1539 1280 1540
rect 1274 1535 1275 1539
rect 1279 1535 1280 1539
rect 1274 1534 1280 1535
rect 1276 1502 1278 1534
rect 1286 1531 1292 1532
rect 1286 1527 1287 1531
rect 1291 1527 1292 1531
rect 1286 1526 1292 1527
rect 1274 1501 1280 1502
rect 1274 1497 1275 1501
rect 1279 1497 1280 1501
rect 1274 1496 1280 1497
rect 110 1492 116 1493
rect 486 1495 492 1496
rect 486 1491 487 1495
rect 491 1491 492 1495
rect 486 1490 492 1491
rect 622 1495 628 1496
rect 622 1491 623 1495
rect 627 1491 628 1495
rect 622 1490 628 1491
rect 758 1495 764 1496
rect 758 1491 759 1495
rect 763 1491 764 1495
rect 758 1490 764 1491
rect 894 1495 900 1496
rect 894 1491 895 1495
rect 899 1491 900 1495
rect 894 1490 900 1491
rect 1030 1495 1036 1496
rect 1030 1491 1031 1495
rect 1035 1491 1036 1495
rect 1030 1490 1036 1491
rect 510 1480 516 1481
rect 110 1479 116 1480
rect 110 1475 111 1479
rect 115 1475 116 1479
rect 510 1476 511 1480
rect 515 1476 516 1480
rect 510 1475 516 1476
rect 646 1480 652 1481
rect 646 1476 647 1480
rect 651 1476 652 1480
rect 646 1475 652 1476
rect 782 1480 788 1481
rect 782 1476 783 1480
rect 787 1476 788 1480
rect 782 1475 788 1476
rect 918 1480 924 1481
rect 918 1476 919 1480
rect 923 1476 924 1480
rect 918 1475 924 1476
rect 1054 1480 1060 1481
rect 1054 1476 1055 1480
rect 1059 1476 1060 1480
rect 1054 1475 1060 1476
rect 110 1474 116 1475
rect 112 1435 114 1474
rect 512 1435 514 1475
rect 648 1435 650 1475
rect 784 1435 786 1475
rect 920 1435 922 1475
rect 1056 1435 1058 1475
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 511 1434 515 1435
rect 511 1429 515 1430
rect 647 1434 651 1435
rect 647 1429 651 1430
rect 743 1434 747 1435
rect 743 1429 747 1430
rect 783 1434 787 1435
rect 783 1429 787 1430
rect 887 1434 891 1435
rect 887 1429 891 1430
rect 919 1434 923 1435
rect 919 1429 923 1430
rect 1031 1434 1035 1435
rect 1031 1429 1035 1430
rect 1055 1434 1059 1435
rect 1055 1429 1059 1430
rect 112 1406 114 1429
rect 110 1405 116 1406
rect 744 1405 746 1429
rect 888 1405 890 1429
rect 1032 1405 1034 1429
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 110 1400 116 1401
rect 742 1404 748 1405
rect 742 1400 743 1404
rect 747 1400 748 1404
rect 742 1399 748 1400
rect 886 1404 892 1405
rect 886 1400 887 1404
rect 891 1400 892 1404
rect 886 1399 892 1400
rect 1030 1404 1036 1405
rect 1030 1400 1031 1404
rect 1035 1400 1036 1404
rect 1030 1399 1036 1400
rect 718 1389 724 1390
rect 110 1387 116 1388
rect 110 1383 111 1387
rect 115 1383 116 1387
rect 718 1385 719 1389
rect 723 1385 724 1389
rect 718 1384 724 1385
rect 862 1389 868 1390
rect 862 1385 863 1389
rect 867 1385 868 1389
rect 862 1384 868 1385
rect 1006 1389 1012 1390
rect 1006 1385 1007 1389
rect 1011 1385 1012 1389
rect 1006 1384 1012 1385
rect 110 1382 116 1383
rect 112 1327 114 1382
rect 720 1327 722 1384
rect 864 1327 866 1384
rect 874 1383 880 1384
rect 874 1379 875 1383
rect 879 1379 880 1383
rect 874 1378 880 1379
rect 876 1348 878 1378
rect 874 1347 880 1348
rect 874 1343 875 1347
rect 879 1343 880 1347
rect 874 1342 880 1343
rect 1008 1327 1010 1384
rect 1018 1383 1024 1384
rect 1018 1379 1019 1383
rect 1023 1379 1024 1383
rect 1018 1378 1024 1379
rect 1020 1348 1022 1378
rect 1120 1364 1122 1496
rect 1166 1495 1172 1496
rect 1166 1491 1167 1495
rect 1171 1491 1172 1495
rect 1166 1490 1172 1491
rect 1190 1480 1196 1481
rect 1190 1476 1191 1480
rect 1195 1476 1196 1480
rect 1190 1475 1196 1476
rect 1192 1435 1194 1475
rect 1175 1434 1179 1435
rect 1175 1429 1179 1430
rect 1191 1434 1195 1435
rect 1191 1429 1195 1430
rect 1176 1405 1178 1429
rect 1174 1404 1180 1405
rect 1174 1400 1175 1404
rect 1179 1400 1180 1404
rect 1174 1399 1180 1400
rect 1150 1389 1156 1390
rect 1150 1385 1151 1389
rect 1155 1385 1156 1389
rect 1150 1384 1156 1385
rect 1288 1384 1290 1526
rect 1304 1496 1306 1545
rect 1440 1496 1442 1545
rect 1546 1539 1552 1540
rect 1546 1535 1547 1539
rect 1551 1535 1552 1539
rect 1546 1534 1552 1535
rect 1548 1502 1550 1534
rect 1546 1501 1552 1502
rect 1546 1497 1547 1501
rect 1551 1497 1552 1501
rect 1546 1496 1552 1497
rect 1576 1496 1578 1545
rect 1720 1498 1722 1545
rect 1718 1497 1724 1498
rect 1302 1495 1308 1496
rect 1302 1491 1303 1495
rect 1307 1491 1308 1495
rect 1302 1490 1308 1491
rect 1438 1495 1444 1496
rect 1438 1491 1439 1495
rect 1443 1491 1444 1495
rect 1438 1490 1444 1491
rect 1574 1495 1580 1496
rect 1574 1491 1575 1495
rect 1579 1491 1580 1495
rect 1718 1493 1719 1497
rect 1723 1493 1724 1497
rect 1718 1492 1724 1493
rect 1574 1490 1580 1491
rect 1326 1480 1332 1481
rect 1326 1476 1327 1480
rect 1331 1476 1332 1480
rect 1326 1475 1332 1476
rect 1462 1480 1468 1481
rect 1462 1476 1463 1480
rect 1467 1476 1468 1480
rect 1462 1475 1468 1476
rect 1598 1480 1604 1481
rect 1598 1476 1599 1480
rect 1603 1476 1604 1480
rect 1598 1475 1604 1476
rect 1718 1479 1724 1480
rect 1718 1475 1719 1479
rect 1723 1475 1724 1479
rect 1328 1435 1330 1475
rect 1464 1435 1466 1475
rect 1600 1435 1602 1475
rect 1718 1474 1724 1475
rect 1720 1435 1722 1474
rect 1319 1434 1323 1435
rect 1319 1429 1323 1430
rect 1327 1434 1331 1435
rect 1327 1429 1331 1430
rect 1463 1434 1467 1435
rect 1463 1429 1467 1430
rect 1599 1434 1603 1435
rect 1599 1429 1603 1430
rect 1719 1434 1723 1435
rect 1719 1429 1723 1430
rect 1320 1405 1322 1429
rect 1464 1405 1466 1429
rect 1600 1405 1602 1429
rect 1720 1406 1722 1429
rect 1718 1405 1724 1406
rect 1318 1404 1324 1405
rect 1318 1400 1319 1404
rect 1323 1400 1324 1404
rect 1318 1399 1324 1400
rect 1462 1404 1468 1405
rect 1462 1400 1463 1404
rect 1467 1400 1468 1404
rect 1462 1399 1468 1400
rect 1598 1404 1604 1405
rect 1598 1400 1599 1404
rect 1603 1400 1604 1404
rect 1718 1401 1719 1405
rect 1723 1401 1724 1405
rect 1718 1400 1724 1401
rect 1598 1399 1604 1400
rect 1294 1389 1300 1390
rect 1294 1385 1295 1389
rect 1299 1385 1300 1389
rect 1294 1384 1300 1385
rect 1438 1389 1444 1390
rect 1438 1385 1439 1389
rect 1443 1385 1444 1389
rect 1438 1384 1444 1385
rect 1574 1389 1580 1390
rect 1574 1385 1575 1389
rect 1579 1385 1580 1389
rect 1574 1384 1580 1385
rect 1718 1387 1724 1388
rect 1118 1363 1124 1364
rect 1118 1359 1119 1363
rect 1123 1359 1124 1363
rect 1118 1358 1124 1359
rect 1018 1347 1024 1348
rect 1018 1343 1019 1347
rect 1023 1343 1024 1347
rect 1018 1342 1024 1343
rect 1152 1327 1154 1384
rect 1162 1383 1168 1384
rect 1162 1379 1163 1383
rect 1167 1379 1168 1383
rect 1162 1378 1168 1379
rect 1258 1383 1264 1384
rect 1258 1379 1259 1383
rect 1263 1379 1264 1383
rect 1258 1378 1264 1379
rect 1286 1383 1292 1384
rect 1286 1379 1287 1383
rect 1291 1379 1292 1383
rect 1286 1378 1292 1379
rect 1164 1348 1166 1378
rect 1162 1347 1168 1348
rect 1162 1343 1163 1347
rect 1167 1343 1168 1347
rect 1162 1342 1168 1343
rect 111 1326 115 1327
rect 111 1321 115 1322
rect 183 1326 187 1327
rect 183 1321 187 1322
rect 415 1326 419 1327
rect 415 1321 419 1322
rect 679 1326 683 1327
rect 679 1321 683 1322
rect 719 1326 723 1327
rect 719 1321 723 1322
rect 863 1326 867 1327
rect 863 1321 867 1322
rect 975 1326 979 1327
rect 975 1321 979 1322
rect 1007 1326 1011 1327
rect 1007 1321 1011 1322
rect 1151 1326 1155 1327
rect 1151 1321 1155 1322
rect 112 1274 114 1321
rect 110 1273 116 1274
rect 110 1269 111 1273
rect 115 1269 116 1273
rect 184 1272 186 1321
rect 358 1315 364 1316
rect 358 1311 359 1315
rect 363 1311 364 1315
rect 358 1310 364 1311
rect 360 1280 362 1310
rect 358 1279 364 1280
rect 270 1277 276 1278
rect 270 1273 271 1277
rect 275 1273 276 1277
rect 358 1275 359 1279
rect 363 1275 364 1279
rect 358 1274 364 1275
rect 270 1272 276 1273
rect 416 1272 418 1321
rect 530 1315 536 1316
rect 530 1311 531 1315
rect 535 1311 536 1315
rect 530 1310 536 1311
rect 532 1280 534 1310
rect 530 1279 536 1280
rect 530 1275 531 1279
rect 535 1275 536 1279
rect 530 1274 536 1275
rect 680 1272 682 1321
rect 886 1315 892 1316
rect 886 1311 887 1315
rect 891 1311 892 1315
rect 886 1310 892 1311
rect 888 1280 890 1310
rect 886 1279 892 1280
rect 886 1275 887 1279
rect 891 1275 892 1279
rect 886 1274 892 1275
rect 976 1272 978 1321
rect 1260 1316 1262 1378
rect 1296 1327 1298 1384
rect 1378 1347 1384 1348
rect 1378 1343 1379 1347
rect 1383 1343 1384 1347
rect 1378 1342 1384 1343
rect 1287 1326 1291 1327
rect 1287 1321 1291 1322
rect 1295 1326 1299 1327
rect 1295 1321 1299 1322
rect 1190 1315 1196 1316
rect 1190 1311 1191 1315
rect 1195 1311 1196 1315
rect 1190 1310 1196 1311
rect 1258 1315 1264 1316
rect 1258 1311 1259 1315
rect 1263 1311 1264 1315
rect 1258 1310 1264 1311
rect 1192 1280 1194 1310
rect 1190 1279 1196 1280
rect 1190 1275 1191 1279
rect 1195 1275 1196 1279
rect 1190 1274 1196 1275
rect 1288 1272 1290 1321
rect 110 1268 116 1269
rect 182 1271 188 1272
rect 182 1267 183 1271
rect 187 1267 188 1271
rect 182 1266 188 1267
rect 206 1256 212 1257
rect 110 1255 116 1256
rect 110 1251 111 1255
rect 115 1251 116 1255
rect 206 1252 207 1256
rect 211 1252 212 1256
rect 206 1251 212 1252
rect 110 1250 116 1251
rect 112 1223 114 1250
rect 208 1223 210 1251
rect 111 1222 115 1223
rect 111 1217 115 1218
rect 159 1222 163 1223
rect 159 1217 163 1218
rect 207 1222 211 1223
rect 207 1217 211 1218
rect 112 1194 114 1217
rect 110 1193 116 1194
rect 160 1193 162 1217
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 110 1188 116 1189
rect 158 1192 164 1193
rect 158 1188 159 1192
rect 163 1188 164 1192
rect 158 1187 164 1188
rect 134 1177 140 1178
rect 110 1175 116 1176
rect 110 1171 111 1175
rect 115 1171 116 1175
rect 134 1173 135 1177
rect 139 1173 140 1177
rect 134 1172 140 1173
rect 110 1170 116 1171
rect 112 1107 114 1170
rect 136 1107 138 1172
rect 272 1136 274 1272
rect 414 1271 420 1272
rect 414 1267 415 1271
rect 419 1267 420 1271
rect 414 1266 420 1267
rect 678 1271 684 1272
rect 678 1267 679 1271
rect 683 1267 684 1271
rect 678 1266 684 1267
rect 974 1271 980 1272
rect 974 1267 975 1271
rect 979 1267 980 1271
rect 974 1266 980 1267
rect 1286 1271 1292 1272
rect 1286 1267 1287 1271
rect 1291 1267 1292 1271
rect 1286 1266 1292 1267
rect 438 1256 444 1257
rect 438 1252 439 1256
rect 443 1252 444 1256
rect 438 1251 444 1252
rect 702 1256 708 1257
rect 702 1252 703 1256
rect 707 1252 708 1256
rect 702 1251 708 1252
rect 998 1256 1004 1257
rect 998 1252 999 1256
rect 1003 1252 1004 1256
rect 998 1251 1004 1252
rect 1310 1256 1316 1257
rect 1310 1252 1311 1256
rect 1315 1252 1316 1256
rect 1310 1251 1316 1252
rect 440 1223 442 1251
rect 704 1223 706 1251
rect 1000 1223 1002 1251
rect 1312 1223 1314 1251
rect 335 1222 339 1223
rect 335 1217 339 1218
rect 439 1222 443 1223
rect 439 1217 443 1218
rect 559 1222 563 1223
rect 559 1217 563 1218
rect 703 1222 707 1223
rect 703 1217 707 1218
rect 799 1222 803 1223
rect 799 1217 803 1218
rect 999 1222 1003 1223
rect 999 1217 1003 1218
rect 1063 1222 1067 1223
rect 1063 1217 1067 1218
rect 1311 1222 1315 1223
rect 1311 1217 1315 1218
rect 1335 1222 1339 1223
rect 1335 1217 1339 1218
rect 336 1193 338 1217
rect 560 1193 562 1217
rect 800 1193 802 1217
rect 1064 1193 1066 1217
rect 1336 1193 1338 1217
rect 334 1192 340 1193
rect 334 1188 335 1192
rect 339 1188 340 1192
rect 334 1187 340 1188
rect 558 1192 564 1193
rect 558 1188 559 1192
rect 563 1188 564 1192
rect 558 1187 564 1188
rect 798 1192 804 1193
rect 798 1188 799 1192
rect 803 1188 804 1192
rect 798 1187 804 1188
rect 1062 1192 1068 1193
rect 1062 1188 1063 1192
rect 1067 1188 1068 1192
rect 1062 1187 1068 1188
rect 1334 1192 1340 1193
rect 1334 1188 1335 1192
rect 1339 1188 1340 1192
rect 1334 1187 1340 1188
rect 310 1177 316 1178
rect 310 1173 311 1177
rect 315 1173 316 1177
rect 310 1172 316 1173
rect 534 1177 540 1178
rect 534 1173 535 1177
rect 539 1173 540 1177
rect 534 1172 540 1173
rect 774 1177 780 1178
rect 774 1173 775 1177
rect 779 1173 780 1177
rect 774 1172 780 1173
rect 1038 1177 1044 1178
rect 1038 1173 1039 1177
rect 1043 1173 1044 1177
rect 1038 1172 1044 1173
rect 1310 1177 1316 1178
rect 1310 1173 1311 1177
rect 1315 1173 1316 1177
rect 1310 1172 1316 1173
rect 1380 1172 1382 1342
rect 1440 1327 1442 1384
rect 1576 1327 1578 1384
rect 1586 1383 1592 1384
rect 1586 1379 1587 1383
rect 1591 1379 1592 1383
rect 1586 1378 1592 1379
rect 1674 1383 1680 1384
rect 1674 1379 1675 1383
rect 1679 1379 1680 1383
rect 1718 1383 1719 1387
rect 1723 1383 1724 1387
rect 1718 1382 1724 1383
rect 1674 1378 1680 1379
rect 1588 1348 1590 1378
rect 1586 1347 1592 1348
rect 1586 1343 1587 1347
rect 1591 1343 1592 1347
rect 1586 1342 1592 1343
rect 1439 1326 1443 1327
rect 1439 1321 1443 1322
rect 1575 1326 1579 1327
rect 1575 1321 1579 1322
rect 1576 1272 1578 1321
rect 1676 1316 1678 1378
rect 1720 1327 1722 1382
rect 1719 1326 1723 1327
rect 1719 1321 1723 1322
rect 1674 1315 1680 1316
rect 1674 1311 1675 1315
rect 1679 1311 1680 1315
rect 1674 1310 1680 1311
rect 1666 1277 1672 1278
rect 1666 1273 1667 1277
rect 1671 1273 1672 1277
rect 1720 1274 1722 1321
rect 1666 1272 1672 1273
rect 1718 1273 1724 1274
rect 1574 1271 1580 1272
rect 1574 1267 1575 1271
rect 1579 1267 1580 1271
rect 1574 1266 1580 1267
rect 1598 1256 1604 1257
rect 1598 1252 1599 1256
rect 1603 1252 1604 1256
rect 1598 1251 1604 1252
rect 1600 1223 1602 1251
rect 1599 1222 1603 1223
rect 1599 1217 1603 1218
rect 1600 1193 1602 1217
rect 1598 1192 1604 1193
rect 1598 1188 1599 1192
rect 1603 1188 1604 1192
rect 1598 1187 1604 1188
rect 1574 1177 1580 1178
rect 1574 1173 1575 1177
rect 1579 1173 1580 1177
rect 1574 1172 1580 1173
rect 270 1135 276 1136
rect 270 1131 271 1135
rect 275 1131 276 1135
rect 270 1130 276 1131
rect 312 1107 314 1172
rect 322 1171 328 1172
rect 322 1167 323 1171
rect 327 1167 328 1171
rect 322 1166 328 1167
rect 324 1136 326 1166
rect 322 1135 328 1136
rect 322 1131 323 1135
rect 327 1131 328 1135
rect 322 1130 328 1131
rect 536 1107 538 1172
rect 546 1171 552 1172
rect 546 1167 547 1171
rect 551 1167 552 1171
rect 546 1166 552 1167
rect 548 1136 550 1166
rect 546 1135 552 1136
rect 546 1131 547 1135
rect 551 1131 552 1135
rect 546 1130 552 1131
rect 776 1107 778 1172
rect 786 1171 792 1172
rect 786 1167 787 1171
rect 791 1167 792 1171
rect 786 1166 792 1167
rect 788 1136 790 1166
rect 786 1135 792 1136
rect 786 1131 787 1135
rect 791 1131 792 1135
rect 786 1130 792 1131
rect 1040 1107 1042 1172
rect 1050 1171 1056 1172
rect 1050 1167 1051 1171
rect 1055 1167 1056 1171
rect 1050 1166 1056 1167
rect 1090 1171 1096 1172
rect 1090 1167 1091 1171
rect 1095 1167 1096 1171
rect 1090 1166 1096 1167
rect 1052 1136 1054 1166
rect 1050 1135 1056 1136
rect 1050 1131 1051 1135
rect 1055 1131 1056 1135
rect 1050 1130 1056 1131
rect 1092 1108 1094 1166
rect 1090 1107 1096 1108
rect 1312 1107 1314 1172
rect 1378 1171 1384 1172
rect 1378 1167 1379 1171
rect 1383 1167 1384 1171
rect 1378 1166 1384 1167
rect 1374 1135 1380 1136
rect 1374 1131 1375 1135
rect 1379 1131 1380 1135
rect 1374 1130 1380 1131
rect 111 1106 115 1107
rect 111 1101 115 1102
rect 135 1106 139 1107
rect 135 1101 139 1102
rect 223 1106 227 1107
rect 223 1101 227 1102
rect 311 1106 315 1107
rect 311 1101 315 1102
rect 463 1106 467 1107
rect 463 1101 467 1102
rect 535 1106 539 1107
rect 535 1101 539 1102
rect 719 1106 723 1107
rect 719 1101 723 1102
rect 775 1106 779 1107
rect 775 1101 779 1102
rect 991 1106 995 1107
rect 991 1101 995 1102
rect 1039 1106 1043 1107
rect 1090 1103 1091 1107
rect 1095 1103 1096 1107
rect 1090 1102 1096 1103
rect 1271 1106 1275 1107
rect 1039 1101 1043 1102
rect 1271 1101 1275 1102
rect 1311 1106 1315 1107
rect 1311 1101 1315 1102
rect 112 1054 114 1101
rect 110 1053 116 1054
rect 110 1049 111 1053
rect 115 1049 116 1053
rect 224 1052 226 1101
rect 330 1095 336 1096
rect 330 1091 331 1095
rect 335 1091 336 1095
rect 330 1090 336 1091
rect 332 1058 334 1090
rect 330 1057 336 1058
rect 330 1053 331 1057
rect 335 1053 336 1057
rect 330 1052 336 1053
rect 464 1052 466 1101
rect 586 1095 592 1096
rect 586 1091 587 1095
rect 591 1091 592 1095
rect 586 1090 592 1091
rect 588 1058 590 1090
rect 586 1057 592 1058
rect 586 1053 587 1057
rect 591 1053 592 1057
rect 586 1052 592 1053
rect 720 1052 722 1101
rect 842 1095 848 1096
rect 842 1091 843 1095
rect 847 1091 848 1095
rect 842 1090 848 1091
rect 844 1058 846 1090
rect 842 1057 848 1058
rect 842 1053 843 1057
rect 847 1053 848 1057
rect 842 1052 848 1053
rect 992 1052 994 1101
rect 1094 1057 1100 1058
rect 1094 1053 1095 1057
rect 1099 1053 1100 1057
rect 1094 1052 1100 1053
rect 1272 1052 1274 1101
rect 1376 1058 1378 1130
rect 1576 1107 1578 1172
rect 1658 1171 1664 1172
rect 1658 1167 1659 1171
rect 1663 1167 1664 1171
rect 1658 1166 1664 1167
rect 1559 1106 1563 1107
rect 1559 1101 1563 1102
rect 1575 1106 1579 1107
rect 1575 1101 1579 1102
rect 1454 1095 1460 1096
rect 1454 1091 1455 1095
rect 1459 1091 1460 1095
rect 1454 1090 1460 1091
rect 1374 1057 1380 1058
rect 1374 1053 1375 1057
rect 1379 1053 1380 1057
rect 1374 1052 1380 1053
rect 110 1048 116 1049
rect 222 1051 228 1052
rect 222 1047 223 1051
rect 227 1047 228 1051
rect 222 1046 228 1047
rect 462 1051 468 1052
rect 462 1047 463 1051
rect 467 1047 468 1051
rect 462 1046 468 1047
rect 718 1051 724 1052
rect 718 1047 719 1051
rect 723 1047 724 1051
rect 718 1046 724 1047
rect 990 1051 996 1052
rect 990 1047 991 1051
rect 995 1047 996 1051
rect 990 1046 996 1047
rect 246 1036 252 1037
rect 110 1035 116 1036
rect 110 1031 111 1035
rect 115 1031 116 1035
rect 246 1032 247 1036
rect 251 1032 252 1036
rect 246 1031 252 1032
rect 486 1036 492 1037
rect 486 1032 487 1036
rect 491 1032 492 1036
rect 486 1031 492 1032
rect 742 1036 748 1037
rect 742 1032 743 1036
rect 747 1032 748 1036
rect 742 1031 748 1032
rect 1014 1036 1020 1037
rect 1014 1032 1015 1036
rect 1019 1032 1020 1036
rect 1014 1031 1020 1032
rect 110 1030 116 1031
rect 112 1007 114 1030
rect 248 1007 250 1031
rect 488 1007 490 1031
rect 744 1007 746 1031
rect 1016 1007 1018 1031
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 247 1006 251 1007
rect 247 1001 251 1002
rect 463 1006 467 1007
rect 463 1001 467 1002
rect 487 1006 491 1007
rect 487 1001 491 1002
rect 647 1006 651 1007
rect 647 1001 651 1002
rect 743 1006 747 1007
rect 743 1001 747 1002
rect 855 1006 859 1007
rect 855 1001 859 1002
rect 1015 1006 1019 1007
rect 1015 1001 1019 1002
rect 1079 1006 1083 1007
rect 1079 1001 1083 1002
rect 112 978 114 1001
rect 110 977 116 978
rect 464 977 466 1001
rect 558 991 564 992
rect 558 987 559 991
rect 563 987 564 991
rect 558 986 564 987
rect 110 973 111 977
rect 115 973 116 977
rect 110 972 116 973
rect 462 976 468 977
rect 462 972 463 976
rect 467 972 468 976
rect 462 971 468 972
rect 438 961 444 962
rect 110 959 116 960
rect 110 955 111 959
rect 115 955 116 959
rect 438 957 439 961
rect 443 957 444 961
rect 438 956 444 957
rect 110 954 116 955
rect 112 899 114 954
rect 440 899 442 956
rect 560 920 562 986
rect 648 977 650 1001
rect 856 977 858 1001
rect 1080 977 1082 1001
rect 1096 992 1098 1052
rect 1270 1051 1276 1052
rect 1270 1047 1271 1051
rect 1275 1047 1276 1051
rect 1270 1046 1276 1047
rect 1294 1036 1300 1037
rect 1294 1032 1295 1036
rect 1299 1032 1300 1036
rect 1294 1031 1300 1032
rect 1296 1007 1298 1031
rect 1295 1006 1299 1007
rect 1295 1001 1299 1002
rect 1311 1006 1315 1007
rect 1311 1001 1315 1002
rect 1094 991 1100 992
rect 1094 987 1095 991
rect 1099 987 1100 991
rect 1094 986 1100 987
rect 1312 977 1314 1001
rect 646 976 652 977
rect 646 972 647 976
rect 651 972 652 976
rect 646 971 652 972
rect 854 976 860 977
rect 854 972 855 976
rect 859 972 860 976
rect 854 971 860 972
rect 1078 976 1084 977
rect 1078 972 1079 976
rect 1083 972 1084 976
rect 1078 971 1084 972
rect 1310 976 1316 977
rect 1310 972 1311 976
rect 1315 972 1316 976
rect 1310 971 1316 972
rect 622 961 628 962
rect 622 957 623 961
rect 627 957 628 961
rect 622 956 628 957
rect 830 961 836 962
rect 830 957 831 961
rect 835 957 836 961
rect 830 956 836 957
rect 1054 961 1060 962
rect 1054 957 1055 961
rect 1059 957 1060 961
rect 1054 956 1060 957
rect 1286 961 1292 962
rect 1286 957 1287 961
rect 1291 957 1292 961
rect 1286 956 1292 957
rect 558 919 564 920
rect 558 915 559 919
rect 563 915 564 919
rect 558 914 564 915
rect 624 899 626 956
rect 634 955 640 956
rect 634 951 635 955
rect 639 951 640 955
rect 634 950 640 951
rect 636 920 638 950
rect 786 947 792 948
rect 786 943 787 947
rect 791 943 792 947
rect 786 942 792 943
rect 634 919 640 920
rect 634 915 635 919
rect 639 915 640 919
rect 634 914 640 915
rect 111 898 115 899
rect 111 893 115 894
rect 439 898 443 899
rect 439 893 443 894
rect 623 898 627 899
rect 623 893 627 894
rect 687 898 691 899
rect 687 893 691 894
rect 112 846 114 893
rect 110 845 116 846
rect 110 841 111 845
rect 115 841 116 845
rect 688 844 690 893
rect 788 888 790 942
rect 832 899 834 956
rect 842 955 848 956
rect 842 951 843 955
rect 847 951 848 955
rect 842 950 848 951
rect 844 920 846 950
rect 842 919 848 920
rect 842 915 843 919
rect 847 915 848 919
rect 842 914 848 915
rect 1056 899 1058 956
rect 1066 955 1072 956
rect 1066 951 1067 955
rect 1071 951 1072 955
rect 1066 950 1072 951
rect 1068 920 1070 950
rect 1066 919 1072 920
rect 1066 915 1067 919
rect 1071 915 1072 919
rect 1066 914 1072 915
rect 1288 899 1290 956
rect 1298 955 1304 956
rect 1298 951 1299 955
rect 1303 951 1304 955
rect 1298 950 1304 951
rect 1300 920 1302 950
rect 1298 919 1304 920
rect 1298 915 1299 919
rect 1303 915 1304 919
rect 1298 914 1304 915
rect 823 898 827 899
rect 823 893 827 894
rect 831 898 835 899
rect 831 893 835 894
rect 959 898 963 899
rect 959 893 963 894
rect 1055 898 1059 899
rect 1055 893 1059 894
rect 1095 898 1099 899
rect 1095 893 1099 894
rect 1231 898 1235 899
rect 1231 893 1235 894
rect 1287 898 1291 899
rect 1287 893 1291 894
rect 1367 898 1371 899
rect 1367 893 1371 894
rect 786 887 792 888
rect 786 883 787 887
rect 791 883 792 887
rect 786 882 792 883
rect 794 887 800 888
rect 794 883 795 887
rect 799 883 800 887
rect 794 882 800 883
rect 796 850 798 882
rect 794 849 800 850
rect 794 845 795 849
rect 799 845 800 849
rect 794 844 800 845
rect 824 844 826 893
rect 930 887 936 888
rect 930 883 931 887
rect 935 883 936 887
rect 930 882 936 883
rect 932 850 934 882
rect 930 849 936 850
rect 930 845 931 849
rect 935 845 936 849
rect 930 844 936 845
rect 960 844 962 893
rect 1066 887 1072 888
rect 1066 883 1067 887
rect 1071 883 1072 887
rect 1066 882 1072 883
rect 1068 850 1070 882
rect 1066 849 1072 850
rect 1066 845 1067 849
rect 1071 845 1072 849
rect 1066 844 1072 845
rect 1096 844 1098 893
rect 1202 887 1208 888
rect 1202 883 1203 887
rect 1207 883 1208 887
rect 1202 882 1208 883
rect 1204 850 1206 882
rect 1202 849 1208 850
rect 1202 845 1203 849
rect 1207 845 1208 849
rect 1202 844 1208 845
rect 1232 844 1234 893
rect 1318 849 1324 850
rect 1318 845 1319 849
rect 1323 845 1324 849
rect 1318 844 1324 845
rect 1368 844 1370 893
rect 1456 891 1458 1090
rect 1560 1052 1562 1101
rect 1660 1096 1662 1166
rect 1668 1136 1670 1272
rect 1718 1269 1719 1273
rect 1723 1269 1724 1273
rect 1718 1268 1724 1269
rect 1718 1255 1724 1256
rect 1718 1251 1719 1255
rect 1723 1251 1724 1255
rect 1718 1250 1724 1251
rect 1720 1223 1722 1250
rect 1719 1222 1723 1223
rect 1719 1217 1723 1218
rect 1720 1194 1722 1217
rect 1718 1193 1724 1194
rect 1718 1189 1719 1193
rect 1723 1189 1724 1193
rect 1718 1188 1724 1189
rect 1718 1175 1724 1176
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1718 1170 1724 1171
rect 1666 1135 1672 1136
rect 1666 1131 1667 1135
rect 1671 1131 1672 1135
rect 1666 1130 1672 1131
rect 1720 1107 1722 1170
rect 1719 1106 1723 1107
rect 1719 1101 1723 1102
rect 1658 1095 1664 1096
rect 1658 1091 1659 1095
rect 1663 1091 1664 1095
rect 1658 1090 1664 1091
rect 1646 1057 1652 1058
rect 1646 1053 1647 1057
rect 1651 1053 1652 1057
rect 1720 1054 1722 1101
rect 1646 1052 1652 1053
rect 1718 1053 1724 1054
rect 1558 1051 1564 1052
rect 1558 1047 1559 1051
rect 1563 1047 1564 1051
rect 1558 1046 1564 1047
rect 1582 1036 1588 1037
rect 1582 1032 1583 1036
rect 1587 1032 1588 1036
rect 1582 1031 1588 1032
rect 1584 1007 1586 1031
rect 1543 1006 1547 1007
rect 1543 1001 1547 1002
rect 1583 1006 1587 1007
rect 1583 1001 1587 1002
rect 1544 977 1546 1001
rect 1542 976 1548 977
rect 1542 972 1543 976
rect 1547 972 1548 976
rect 1542 971 1548 972
rect 1518 961 1524 962
rect 1518 957 1519 961
rect 1523 957 1524 961
rect 1518 956 1524 957
rect 1520 899 1522 956
rect 1602 955 1608 956
rect 1602 951 1603 955
rect 1607 951 1608 955
rect 1602 950 1608 951
rect 1503 898 1507 899
rect 1503 893 1507 894
rect 1519 898 1523 899
rect 1519 893 1523 894
rect 1456 889 1462 891
rect 1450 883 1456 884
rect 1450 879 1451 883
rect 1455 879 1456 883
rect 1450 878 1456 879
rect 110 840 116 841
rect 686 843 692 844
rect 686 839 687 843
rect 691 839 692 843
rect 686 838 692 839
rect 822 843 828 844
rect 822 839 823 843
rect 827 839 828 843
rect 822 838 828 839
rect 958 843 964 844
rect 958 839 959 843
rect 963 839 964 843
rect 958 838 964 839
rect 1094 843 1100 844
rect 1094 839 1095 843
rect 1099 839 1100 843
rect 1094 838 1100 839
rect 1230 843 1236 844
rect 1230 839 1231 843
rect 1235 839 1236 843
rect 1230 838 1236 839
rect 710 828 716 829
rect 110 827 116 828
rect 110 823 111 827
rect 115 823 116 827
rect 710 824 711 828
rect 715 824 716 828
rect 710 823 716 824
rect 846 828 852 829
rect 846 824 847 828
rect 851 824 852 828
rect 846 823 852 824
rect 982 828 988 829
rect 982 824 983 828
rect 987 824 988 828
rect 982 823 988 824
rect 1118 828 1124 829
rect 1118 824 1119 828
rect 1123 824 1124 828
rect 1118 823 1124 824
rect 1254 828 1260 829
rect 1254 824 1255 828
rect 1259 824 1260 828
rect 1254 823 1260 824
rect 110 822 116 823
rect 112 787 114 822
rect 712 787 714 823
rect 848 787 850 823
rect 984 787 986 823
rect 1120 787 1122 823
rect 1256 787 1258 823
rect 111 786 115 787
rect 111 781 115 782
rect 711 786 715 787
rect 711 781 715 782
rect 815 786 819 787
rect 815 781 819 782
rect 847 786 851 787
rect 847 781 851 782
rect 951 786 955 787
rect 951 781 955 782
rect 983 786 987 787
rect 983 781 987 782
rect 1087 786 1091 787
rect 1087 781 1091 782
rect 1119 786 1123 787
rect 1119 781 1123 782
rect 1223 786 1227 787
rect 1223 781 1227 782
rect 1255 786 1259 787
rect 1255 781 1259 782
rect 112 758 114 781
rect 110 757 116 758
rect 816 757 818 781
rect 952 757 954 781
rect 1088 757 1090 781
rect 1224 757 1226 781
rect 110 753 111 757
rect 115 753 116 757
rect 110 752 116 753
rect 814 756 820 757
rect 814 752 815 756
rect 819 752 820 756
rect 814 751 820 752
rect 950 756 956 757
rect 950 752 951 756
rect 955 752 956 756
rect 950 751 956 752
rect 1086 756 1092 757
rect 1086 752 1087 756
rect 1091 752 1092 756
rect 1086 751 1092 752
rect 1222 756 1228 757
rect 1222 752 1223 756
rect 1227 752 1228 756
rect 1222 751 1228 752
rect 790 741 796 742
rect 110 739 116 740
rect 110 735 111 739
rect 115 735 116 739
rect 790 737 791 741
rect 795 737 796 741
rect 790 736 796 737
rect 926 741 932 742
rect 926 737 927 741
rect 931 737 932 741
rect 926 736 932 737
rect 1062 741 1068 742
rect 1062 737 1063 741
rect 1067 737 1068 741
rect 1062 736 1068 737
rect 1198 741 1204 742
rect 1198 737 1199 741
rect 1203 737 1204 741
rect 1198 736 1204 737
rect 110 734 116 735
rect 112 679 114 734
rect 792 679 794 736
rect 875 700 879 701
rect 874 695 875 700
rect 879 695 880 700
rect 874 694 880 695
rect 928 679 930 736
rect 938 735 944 736
rect 938 731 939 735
rect 943 731 944 735
rect 938 730 944 731
rect 1022 735 1028 736
rect 1022 731 1023 735
rect 1027 731 1028 735
rect 1022 730 1028 731
rect 940 700 942 730
rect 938 699 944 700
rect 938 695 939 699
rect 943 695 944 699
rect 938 694 944 695
rect 111 678 115 679
rect 111 673 115 674
rect 511 678 515 679
rect 511 673 515 674
rect 679 678 683 679
rect 679 673 683 674
rect 791 678 795 679
rect 791 673 795 674
rect 855 678 859 679
rect 855 673 859 674
rect 927 678 931 679
rect 927 673 931 674
rect 112 626 114 673
rect 110 625 116 626
rect 110 621 111 625
rect 115 621 116 625
rect 512 624 514 673
rect 638 667 644 668
rect 594 663 600 664
rect 594 659 595 663
rect 599 659 600 663
rect 638 663 639 667
rect 643 663 644 667
rect 638 662 644 663
rect 594 658 600 659
rect 596 636 598 658
rect 594 635 600 636
rect 594 631 595 635
rect 599 631 600 635
rect 640 632 642 662
rect 594 630 600 631
rect 638 631 644 632
rect 638 627 639 631
rect 643 627 644 631
rect 638 626 644 627
rect 680 624 682 673
rect 782 629 788 630
rect 782 625 783 629
rect 787 625 788 629
rect 782 624 788 625
rect 856 624 858 673
rect 1024 668 1026 730
rect 1064 679 1066 736
rect 1098 735 1104 736
rect 1098 731 1099 735
rect 1103 731 1104 735
rect 1098 730 1104 731
rect 1178 735 1184 736
rect 1178 731 1179 735
rect 1183 731 1184 735
rect 1178 730 1184 731
rect 1100 701 1102 730
rect 1099 700 1103 701
rect 1180 700 1182 730
rect 1099 695 1103 696
rect 1178 699 1184 700
rect 1178 695 1179 699
rect 1183 695 1184 699
rect 1178 694 1184 695
rect 1200 679 1202 736
rect 1320 700 1322 844
rect 1366 843 1372 844
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 1390 828 1396 829
rect 1390 824 1391 828
rect 1395 824 1396 828
rect 1390 823 1396 824
rect 1392 787 1394 823
rect 1359 786 1363 787
rect 1359 781 1363 782
rect 1391 786 1395 787
rect 1391 781 1395 782
rect 1360 757 1362 781
rect 1358 756 1364 757
rect 1358 752 1359 756
rect 1363 752 1364 756
rect 1358 751 1364 752
rect 1334 741 1340 742
rect 1334 737 1335 741
rect 1339 737 1340 741
rect 1334 736 1340 737
rect 1452 736 1454 878
rect 1460 850 1462 889
rect 1458 849 1464 850
rect 1458 845 1459 849
rect 1463 845 1464 849
rect 1458 844 1464 845
rect 1504 844 1506 893
rect 1604 888 1606 950
rect 1648 920 1650 1052
rect 1718 1049 1719 1053
rect 1723 1049 1724 1053
rect 1718 1048 1724 1049
rect 1718 1035 1724 1036
rect 1718 1031 1719 1035
rect 1723 1031 1724 1035
rect 1718 1030 1724 1031
rect 1720 1007 1722 1030
rect 1719 1006 1723 1007
rect 1719 1001 1723 1002
rect 1720 978 1722 1001
rect 1718 977 1724 978
rect 1718 973 1719 977
rect 1723 973 1724 977
rect 1718 972 1724 973
rect 1718 959 1724 960
rect 1718 955 1719 959
rect 1723 955 1724 959
rect 1718 954 1724 955
rect 1646 919 1652 920
rect 1646 915 1647 919
rect 1651 915 1652 919
rect 1646 914 1652 915
rect 1720 899 1722 954
rect 1719 898 1723 899
rect 1719 893 1723 894
rect 1602 887 1608 888
rect 1602 883 1603 887
rect 1607 883 1608 887
rect 1602 882 1608 883
rect 1590 849 1596 850
rect 1590 845 1591 849
rect 1595 845 1596 849
rect 1720 846 1722 893
rect 1590 844 1596 845
rect 1718 845 1724 846
rect 1502 843 1508 844
rect 1502 839 1503 843
rect 1507 839 1508 843
rect 1502 838 1508 839
rect 1526 828 1532 829
rect 1526 824 1527 828
rect 1531 824 1532 828
rect 1526 823 1532 824
rect 1528 787 1530 823
rect 1495 786 1499 787
rect 1495 781 1499 782
rect 1527 786 1531 787
rect 1527 781 1531 782
rect 1496 757 1498 781
rect 1494 756 1500 757
rect 1494 752 1495 756
rect 1499 752 1500 756
rect 1494 751 1500 752
rect 1470 741 1476 742
rect 1470 737 1471 741
rect 1475 737 1476 741
rect 1470 736 1476 737
rect 1318 699 1324 700
rect 1318 695 1319 699
rect 1323 695 1324 699
rect 1318 694 1324 695
rect 1326 699 1332 700
rect 1326 695 1327 699
rect 1331 695 1332 699
rect 1326 694 1332 695
rect 1031 678 1035 679
rect 1031 673 1035 674
rect 1063 678 1067 679
rect 1063 673 1067 674
rect 1199 678 1203 679
rect 1199 673 1203 674
rect 1215 678 1219 679
rect 1215 673 1219 674
rect 1022 667 1028 668
rect 1022 663 1023 667
rect 1027 663 1028 667
rect 1022 662 1028 663
rect 1032 624 1034 673
rect 1206 667 1212 668
rect 1206 663 1207 667
rect 1211 663 1212 667
rect 1206 662 1212 663
rect 110 620 116 621
rect 510 623 516 624
rect 510 619 511 623
rect 515 619 516 623
rect 510 618 516 619
rect 678 623 684 624
rect 678 619 679 623
rect 683 619 684 623
rect 678 618 684 619
rect 534 608 540 609
rect 110 607 116 608
rect 110 603 111 607
rect 115 603 116 607
rect 534 604 535 608
rect 539 604 540 608
rect 534 603 540 604
rect 702 608 708 609
rect 702 604 703 608
rect 707 604 708 608
rect 702 603 708 604
rect 110 602 116 603
rect 112 559 114 602
rect 536 559 538 603
rect 704 559 706 603
rect 111 558 115 559
rect 111 553 115 554
rect 167 558 171 559
rect 167 553 171 554
rect 359 558 363 559
rect 359 553 363 554
rect 535 558 539 559
rect 535 553 539 554
rect 551 558 555 559
rect 551 553 555 554
rect 703 558 707 559
rect 703 553 707 554
rect 743 558 747 559
rect 743 553 747 554
rect 112 530 114 553
rect 110 529 116 530
rect 168 529 170 553
rect 360 529 362 553
rect 552 529 554 553
rect 744 529 746 553
rect 110 525 111 529
rect 115 525 116 529
rect 110 524 116 525
rect 166 528 172 529
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 550 528 556 529
rect 550 524 551 528
rect 555 524 556 528
rect 550 523 556 524
rect 742 528 748 529
rect 742 524 743 528
rect 747 524 748 528
rect 742 523 748 524
rect 142 513 148 514
rect 110 511 116 512
rect 110 507 111 511
rect 115 507 116 511
rect 142 509 143 513
rect 147 509 148 513
rect 142 508 148 509
rect 334 513 340 514
rect 334 509 335 513
rect 339 509 340 513
rect 334 508 340 509
rect 526 513 532 514
rect 526 509 527 513
rect 531 509 532 513
rect 526 508 532 509
rect 718 513 724 514
rect 718 509 719 513
rect 723 509 724 513
rect 718 508 724 509
rect 110 506 116 507
rect 112 435 114 506
rect 144 435 146 508
rect 234 507 240 508
rect 234 503 235 507
rect 239 503 240 507
rect 234 502 240 503
rect 111 434 115 435
rect 111 429 115 430
rect 135 434 139 435
rect 135 429 139 430
rect 143 434 147 435
rect 143 429 147 430
rect 112 382 114 429
rect 110 381 116 382
rect 110 377 111 381
rect 115 377 116 381
rect 136 380 138 429
rect 236 424 238 502
rect 336 435 338 508
rect 474 507 480 508
rect 474 503 475 507
rect 479 503 480 507
rect 474 502 480 503
rect 476 472 478 502
rect 474 471 480 472
rect 474 467 475 471
rect 479 467 480 471
rect 474 466 480 467
rect 528 435 530 508
rect 710 507 716 508
rect 710 503 711 507
rect 715 503 716 507
rect 710 502 716 503
rect 712 472 714 502
rect 710 471 716 472
rect 710 467 711 471
rect 715 467 716 471
rect 710 466 716 467
rect 720 435 722 508
rect 784 472 786 624
rect 854 623 860 624
rect 854 619 855 623
rect 859 619 860 623
rect 854 618 860 619
rect 1030 623 1036 624
rect 1030 619 1031 623
rect 1035 619 1036 623
rect 1030 618 1036 619
rect 878 608 884 609
rect 878 604 879 608
rect 883 604 884 608
rect 878 603 884 604
rect 1054 608 1060 609
rect 1054 604 1055 608
rect 1059 604 1060 608
rect 1054 603 1060 604
rect 880 559 882 603
rect 1056 559 1058 603
rect 879 558 883 559
rect 879 553 883 554
rect 935 558 939 559
rect 935 553 939 554
rect 1055 558 1059 559
rect 1055 553 1059 554
rect 1127 558 1131 559
rect 1127 553 1131 554
rect 936 529 938 553
rect 1128 529 1130 553
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 1126 528 1132 529
rect 1126 524 1127 528
rect 1131 524 1132 528
rect 1126 523 1132 524
rect 910 513 916 514
rect 910 509 911 513
rect 915 509 916 513
rect 910 508 916 509
rect 1102 513 1108 514
rect 1102 509 1103 513
rect 1107 509 1108 513
rect 1102 508 1108 509
rect 1208 508 1210 662
rect 1216 624 1218 673
rect 1328 630 1330 694
rect 1336 679 1338 736
rect 1450 735 1456 736
rect 1450 731 1451 735
rect 1455 731 1456 735
rect 1450 730 1456 731
rect 1472 679 1474 736
rect 1506 735 1512 736
rect 1506 731 1507 735
rect 1511 731 1512 735
rect 1506 730 1512 731
rect 1335 678 1339 679
rect 1335 673 1339 674
rect 1407 678 1411 679
rect 1407 673 1411 674
rect 1471 678 1475 679
rect 1471 673 1475 674
rect 1326 629 1332 630
rect 1326 625 1327 629
rect 1331 625 1332 629
rect 1326 624 1332 625
rect 1408 624 1410 673
rect 1508 668 1510 730
rect 1592 700 1594 844
rect 1718 841 1719 845
rect 1723 841 1724 845
rect 1718 840 1724 841
rect 1718 827 1724 828
rect 1718 823 1719 827
rect 1723 823 1724 827
rect 1718 822 1724 823
rect 1720 787 1722 822
rect 1719 786 1723 787
rect 1719 781 1723 782
rect 1720 758 1722 781
rect 1718 757 1724 758
rect 1718 753 1719 757
rect 1723 753 1724 757
rect 1718 752 1724 753
rect 1718 739 1724 740
rect 1718 735 1719 739
rect 1723 735 1724 739
rect 1718 734 1724 735
rect 1590 699 1596 700
rect 1590 695 1591 699
rect 1595 695 1596 699
rect 1590 694 1596 695
rect 1720 679 1722 734
rect 1719 678 1723 679
rect 1719 673 1723 674
rect 1506 667 1512 668
rect 1506 663 1507 667
rect 1511 663 1512 667
rect 1506 662 1512 663
rect 1494 629 1500 630
rect 1494 625 1495 629
rect 1499 625 1500 629
rect 1720 626 1722 673
rect 1494 624 1500 625
rect 1718 625 1724 626
rect 1214 623 1220 624
rect 1214 619 1215 623
rect 1219 619 1220 623
rect 1214 618 1220 619
rect 1406 623 1412 624
rect 1406 619 1407 623
rect 1411 619 1412 623
rect 1406 618 1412 619
rect 1238 608 1244 609
rect 1238 604 1239 608
rect 1243 604 1244 608
rect 1238 603 1244 604
rect 1430 608 1436 609
rect 1430 604 1431 608
rect 1435 604 1436 608
rect 1430 603 1436 604
rect 1240 559 1242 603
rect 1432 559 1434 603
rect 1239 558 1243 559
rect 1239 553 1243 554
rect 1327 558 1331 559
rect 1327 553 1331 554
rect 1431 558 1435 559
rect 1431 553 1435 554
rect 1328 529 1330 553
rect 1326 528 1332 529
rect 1326 524 1327 528
rect 1331 524 1332 528
rect 1326 523 1332 524
rect 1302 513 1308 514
rect 1302 509 1303 513
rect 1307 509 1308 513
rect 1302 508 1308 509
rect 782 471 788 472
rect 782 467 783 471
rect 787 467 788 471
rect 782 466 788 467
rect 912 435 914 508
rect 1104 435 1106 508
rect 1114 507 1120 508
rect 1114 503 1115 507
rect 1119 503 1120 507
rect 1114 502 1120 503
rect 1206 507 1212 508
rect 1206 503 1207 507
rect 1211 503 1212 507
rect 1206 502 1212 503
rect 1116 472 1118 502
rect 1114 471 1120 472
rect 1114 467 1115 471
rect 1119 467 1120 471
rect 1114 466 1120 467
rect 1274 455 1280 456
rect 1274 451 1275 455
rect 1279 451 1280 455
rect 1274 450 1280 451
rect 335 434 339 435
rect 335 429 339 430
rect 351 434 355 435
rect 351 429 355 430
rect 527 434 531 435
rect 527 429 531 430
rect 615 434 619 435
rect 615 429 619 430
rect 719 434 723 435
rect 719 429 723 430
rect 895 434 899 435
rect 895 429 899 430
rect 911 434 915 435
rect 911 429 915 430
rect 1103 434 1107 435
rect 1103 429 1107 430
rect 1183 434 1187 435
rect 1183 429 1187 430
rect 234 423 240 424
rect 234 419 235 423
rect 239 419 240 423
rect 234 418 240 419
rect 242 423 248 424
rect 242 419 243 423
rect 247 419 248 423
rect 242 418 248 419
rect 244 386 246 418
rect 242 385 248 386
rect 242 381 243 385
rect 247 381 248 385
rect 242 380 248 381
rect 352 380 354 429
rect 474 423 480 424
rect 474 419 475 423
rect 479 419 480 423
rect 474 418 480 419
rect 476 386 478 418
rect 474 385 480 386
rect 474 381 475 385
rect 479 381 480 385
rect 474 380 480 381
rect 616 380 618 429
rect 738 423 744 424
rect 738 419 739 423
rect 743 419 744 423
rect 738 418 744 419
rect 740 386 742 418
rect 738 385 744 386
rect 738 381 739 385
rect 743 381 744 385
rect 738 380 744 381
rect 896 380 898 429
rect 982 385 988 386
rect 982 381 983 385
rect 987 381 988 385
rect 982 380 988 381
rect 1184 380 1186 429
rect 1266 419 1272 420
rect 1266 415 1267 419
rect 1271 415 1272 419
rect 1266 414 1272 415
rect 110 376 116 377
rect 134 379 140 380
rect 134 375 135 379
rect 139 375 140 379
rect 134 374 140 375
rect 350 379 356 380
rect 350 375 351 379
rect 355 375 356 379
rect 350 374 356 375
rect 614 379 620 380
rect 614 375 615 379
rect 619 375 620 379
rect 614 374 620 375
rect 894 379 900 380
rect 894 375 895 379
rect 899 375 900 379
rect 894 374 900 375
rect 158 364 164 365
rect 110 363 116 364
rect 110 359 111 363
rect 115 359 116 363
rect 158 360 159 364
rect 163 360 164 364
rect 158 359 164 360
rect 374 364 380 365
rect 374 360 375 364
rect 379 360 380 364
rect 374 359 380 360
rect 638 364 644 365
rect 638 360 639 364
rect 643 360 644 364
rect 638 359 644 360
rect 918 364 924 365
rect 918 360 919 364
rect 923 360 924 364
rect 918 359 924 360
rect 110 358 116 359
rect 112 327 114 358
rect 160 327 162 359
rect 376 327 378 359
rect 640 327 642 359
rect 920 327 922 359
rect 111 326 115 327
rect 111 321 115 322
rect 159 326 163 327
rect 159 321 163 322
rect 223 326 227 327
rect 223 321 227 322
rect 375 326 379 327
rect 375 321 379 322
rect 455 326 459 327
rect 455 321 459 322
rect 639 326 643 327
rect 639 321 643 322
rect 687 326 691 327
rect 687 321 691 322
rect 919 326 923 327
rect 919 321 923 322
rect 112 298 114 321
rect 110 297 116 298
rect 224 297 226 321
rect 456 297 458 321
rect 688 297 690 321
rect 920 297 922 321
rect 110 293 111 297
rect 115 293 116 297
rect 110 292 116 293
rect 222 296 228 297
rect 222 292 223 296
rect 227 292 228 296
rect 222 291 228 292
rect 454 296 460 297
rect 454 292 455 296
rect 459 292 460 296
rect 454 291 460 292
rect 686 296 692 297
rect 686 292 687 296
rect 691 292 692 296
rect 686 291 692 292
rect 918 296 924 297
rect 918 292 919 296
rect 923 292 924 296
rect 918 291 924 292
rect 198 281 204 282
rect 110 279 116 280
rect 110 275 111 279
rect 115 275 116 279
rect 198 277 199 281
rect 203 277 204 281
rect 198 276 204 277
rect 430 281 436 282
rect 430 277 431 281
rect 435 277 436 281
rect 430 276 436 277
rect 662 281 668 282
rect 662 277 663 281
rect 667 277 668 281
rect 662 276 668 277
rect 894 281 900 282
rect 894 277 895 281
rect 899 277 900 281
rect 894 276 900 277
rect 110 274 116 275
rect 112 207 114 274
rect 200 207 202 276
rect 302 275 308 276
rect 302 271 303 275
rect 307 271 308 275
rect 302 270 308 271
rect 374 275 380 276
rect 374 271 375 275
rect 379 271 380 275
rect 374 270 380 271
rect 111 206 115 207
rect 111 201 115 202
rect 199 206 203 207
rect 199 201 203 202
rect 112 154 114 201
rect 304 196 306 270
rect 376 240 378 270
rect 374 239 380 240
rect 374 235 375 239
rect 379 235 380 239
rect 374 234 380 235
rect 432 207 434 276
rect 546 275 552 276
rect 546 271 547 275
rect 551 271 552 275
rect 546 270 552 271
rect 548 240 550 270
rect 546 239 552 240
rect 546 235 547 239
rect 551 235 552 239
rect 546 234 552 235
rect 664 207 666 276
rect 896 207 898 276
rect 984 256 986 380
rect 1182 379 1188 380
rect 1182 375 1183 379
rect 1187 375 1188 379
rect 1182 374 1188 375
rect 1206 364 1212 365
rect 1206 360 1207 364
rect 1211 360 1212 364
rect 1206 359 1212 360
rect 1208 327 1210 359
rect 1151 326 1155 327
rect 1151 321 1155 322
rect 1207 326 1211 327
rect 1207 321 1211 322
rect 1152 297 1154 321
rect 1150 296 1156 297
rect 1150 292 1151 296
rect 1155 292 1156 296
rect 1150 291 1156 292
rect 1126 281 1132 282
rect 1126 277 1127 281
rect 1131 277 1132 281
rect 1126 276 1132 277
rect 1268 276 1270 414
rect 1276 386 1278 450
rect 1304 435 1306 508
rect 1496 472 1498 624
rect 1718 621 1719 625
rect 1723 621 1724 625
rect 1718 620 1724 621
rect 1718 607 1724 608
rect 1718 603 1719 607
rect 1723 603 1724 607
rect 1718 602 1724 603
rect 1720 559 1722 602
rect 1527 558 1531 559
rect 1527 553 1531 554
rect 1719 558 1723 559
rect 1719 553 1723 554
rect 1528 529 1530 553
rect 1720 530 1722 553
rect 1718 529 1724 530
rect 1526 528 1532 529
rect 1526 524 1527 528
rect 1531 524 1532 528
rect 1718 525 1719 529
rect 1723 525 1724 529
rect 1718 524 1724 525
rect 1526 523 1532 524
rect 1502 513 1508 514
rect 1502 509 1503 513
rect 1507 509 1508 513
rect 1502 508 1508 509
rect 1718 511 1724 512
rect 1494 471 1500 472
rect 1494 467 1495 471
rect 1499 467 1500 471
rect 1494 466 1500 467
rect 1504 435 1506 508
rect 1514 507 1520 508
rect 1514 503 1515 507
rect 1519 503 1520 507
rect 1514 502 1520 503
rect 1570 507 1576 508
rect 1570 503 1571 507
rect 1575 503 1576 507
rect 1718 507 1719 511
rect 1723 507 1724 511
rect 1718 506 1724 507
rect 1570 502 1576 503
rect 1516 472 1518 502
rect 1514 471 1520 472
rect 1514 467 1515 471
rect 1519 467 1520 471
rect 1514 466 1520 467
rect 1303 434 1307 435
rect 1303 429 1307 430
rect 1471 434 1475 435
rect 1471 429 1475 430
rect 1503 434 1507 435
rect 1503 429 1507 430
rect 1274 385 1280 386
rect 1274 381 1275 385
rect 1279 381 1280 385
rect 1274 380 1280 381
rect 1472 380 1474 429
rect 1572 424 1574 502
rect 1720 435 1722 506
rect 1719 434 1723 435
rect 1719 429 1723 430
rect 1570 423 1576 424
rect 1570 419 1571 423
rect 1575 419 1576 423
rect 1570 418 1576 419
rect 1558 385 1564 386
rect 1558 381 1559 385
rect 1563 381 1564 385
rect 1720 382 1722 429
rect 1558 380 1564 381
rect 1718 381 1724 382
rect 1470 379 1476 380
rect 1470 375 1471 379
rect 1475 375 1476 379
rect 1470 374 1476 375
rect 1494 364 1500 365
rect 1494 360 1495 364
rect 1499 360 1500 364
rect 1494 359 1500 360
rect 1496 327 1498 359
rect 1383 326 1387 327
rect 1383 321 1387 322
rect 1495 326 1499 327
rect 1495 321 1499 322
rect 1384 297 1386 321
rect 1382 296 1388 297
rect 1382 292 1383 296
rect 1387 292 1388 296
rect 1382 291 1388 292
rect 1358 281 1364 282
rect 1358 277 1359 281
rect 1363 277 1364 281
rect 1358 276 1364 277
rect 982 255 988 256
rect 982 251 983 255
rect 987 251 988 255
rect 982 250 988 251
rect 1128 207 1130 276
rect 1138 275 1144 276
rect 1138 271 1139 275
rect 1143 271 1144 275
rect 1138 270 1144 271
rect 1266 275 1272 276
rect 1266 271 1267 275
rect 1271 271 1272 275
rect 1266 270 1272 271
rect 1140 240 1142 270
rect 1138 239 1144 240
rect 1138 235 1139 239
rect 1143 235 1144 239
rect 1138 234 1144 235
rect 1326 223 1332 224
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 1326 218 1332 219
rect 311 206 315 207
rect 311 201 315 202
rect 431 206 435 207
rect 431 201 435 202
rect 447 206 451 207
rect 447 201 451 202
rect 591 206 595 207
rect 591 201 595 202
rect 663 206 667 207
rect 663 201 667 202
rect 743 206 747 207
rect 743 201 747 202
rect 895 206 899 207
rect 895 201 899 202
rect 903 206 907 207
rect 903 201 907 202
rect 1071 206 1075 207
rect 1071 201 1075 202
rect 1127 206 1131 207
rect 1127 201 1131 202
rect 1239 206 1243 207
rect 1239 201 1243 202
rect 302 195 308 196
rect 302 191 303 195
rect 307 191 308 195
rect 302 190 308 191
rect 110 153 116 154
rect 110 149 111 153
rect 115 149 116 153
rect 312 152 314 201
rect 422 195 428 196
rect 422 191 423 195
rect 427 191 428 195
rect 422 190 428 191
rect 424 158 426 190
rect 422 157 428 158
rect 422 153 423 157
rect 427 153 428 157
rect 422 152 428 153
rect 448 152 450 201
rect 554 195 560 196
rect 554 191 555 195
rect 559 191 560 195
rect 554 190 560 191
rect 556 158 558 190
rect 554 157 560 158
rect 554 153 555 157
rect 559 153 560 157
rect 554 152 560 153
rect 592 152 594 201
rect 714 195 720 196
rect 714 191 715 195
rect 719 191 720 195
rect 714 190 720 191
rect 716 158 718 190
rect 714 157 720 158
rect 714 153 715 157
rect 719 153 720 157
rect 714 152 720 153
rect 744 152 746 201
rect 866 195 872 196
rect 866 191 867 195
rect 871 191 872 195
rect 866 190 872 191
rect 868 158 870 190
rect 866 157 872 158
rect 866 153 867 157
rect 871 153 872 157
rect 866 152 872 153
rect 904 152 906 201
rect 1010 195 1016 196
rect 1010 191 1011 195
rect 1015 191 1016 195
rect 1010 190 1016 191
rect 1012 158 1014 190
rect 1010 157 1016 158
rect 1010 153 1011 157
rect 1015 153 1016 157
rect 1010 152 1016 153
rect 1072 152 1074 201
rect 1178 195 1184 196
rect 1178 191 1179 195
rect 1183 191 1184 195
rect 1178 190 1184 191
rect 1180 158 1182 190
rect 1178 157 1184 158
rect 1178 153 1179 157
rect 1183 153 1184 157
rect 1178 152 1184 153
rect 1240 152 1242 201
rect 1328 158 1330 218
rect 1360 207 1362 276
rect 1560 240 1562 380
rect 1718 377 1719 381
rect 1723 377 1724 381
rect 1718 376 1724 377
rect 1718 363 1724 364
rect 1718 359 1719 363
rect 1723 359 1724 363
rect 1718 358 1724 359
rect 1720 327 1722 358
rect 1599 326 1603 327
rect 1599 321 1603 322
rect 1719 326 1723 327
rect 1719 321 1723 322
rect 1600 297 1602 321
rect 1720 298 1722 321
rect 1718 297 1724 298
rect 1598 296 1604 297
rect 1598 292 1599 296
rect 1603 292 1604 296
rect 1718 293 1719 297
rect 1723 293 1724 297
rect 1718 292 1724 293
rect 1598 291 1604 292
rect 1574 281 1580 282
rect 1574 277 1575 281
rect 1579 277 1580 281
rect 1574 276 1580 277
rect 1718 279 1724 280
rect 1558 239 1564 240
rect 1558 235 1559 239
rect 1563 235 1564 239
rect 1558 234 1564 235
rect 1576 207 1578 276
rect 1586 275 1592 276
rect 1586 271 1587 275
rect 1591 271 1592 275
rect 1586 270 1592 271
rect 1674 275 1680 276
rect 1674 271 1675 275
rect 1679 271 1680 275
rect 1718 275 1719 279
rect 1723 275 1724 279
rect 1718 274 1724 275
rect 1674 270 1680 271
rect 1588 240 1590 270
rect 1586 239 1592 240
rect 1586 235 1587 239
rect 1591 235 1592 239
rect 1586 234 1592 235
rect 1359 206 1363 207
rect 1359 201 1363 202
rect 1415 206 1419 207
rect 1415 201 1419 202
rect 1575 206 1579 207
rect 1575 201 1579 202
rect 1326 157 1332 158
rect 1326 153 1327 157
rect 1331 153 1332 157
rect 1326 152 1332 153
rect 1416 152 1418 201
rect 1498 191 1504 192
rect 1498 187 1499 191
rect 1503 187 1504 191
rect 1498 186 1504 187
rect 1500 160 1502 186
rect 1498 159 1504 160
rect 1498 155 1499 159
rect 1503 155 1504 159
rect 1498 154 1504 155
rect 1576 152 1578 201
rect 1676 196 1678 270
rect 1720 207 1722 274
rect 1719 206 1723 207
rect 1719 201 1723 202
rect 1674 195 1680 196
rect 1674 191 1675 195
rect 1679 191 1680 195
rect 1674 190 1680 191
rect 1720 154 1722 201
rect 1718 153 1724 154
rect 110 148 116 149
rect 310 151 316 152
rect 310 147 311 151
rect 315 147 316 151
rect 310 146 316 147
rect 446 151 452 152
rect 446 147 447 151
rect 451 147 452 151
rect 446 146 452 147
rect 590 151 596 152
rect 590 147 591 151
rect 595 147 596 151
rect 590 146 596 147
rect 742 151 748 152
rect 742 147 743 151
rect 747 147 748 151
rect 742 146 748 147
rect 902 151 908 152
rect 902 147 903 151
rect 907 147 908 151
rect 902 146 908 147
rect 1070 151 1076 152
rect 1070 147 1071 151
rect 1075 147 1076 151
rect 1070 146 1076 147
rect 1238 151 1244 152
rect 1238 147 1239 151
rect 1243 147 1244 151
rect 1238 146 1244 147
rect 1414 151 1420 152
rect 1414 147 1415 151
rect 1419 147 1420 151
rect 1414 146 1420 147
rect 1574 151 1580 152
rect 1574 147 1575 151
rect 1579 147 1580 151
rect 1718 149 1719 153
rect 1723 149 1724 153
rect 1718 148 1724 149
rect 1574 146 1580 147
rect 334 136 340 137
rect 110 135 116 136
rect 110 131 111 135
rect 115 131 116 135
rect 334 132 335 136
rect 339 132 340 136
rect 334 131 340 132
rect 470 136 476 137
rect 470 132 471 136
rect 475 132 476 136
rect 470 131 476 132
rect 614 136 620 137
rect 614 132 615 136
rect 619 132 620 136
rect 614 131 620 132
rect 766 136 772 137
rect 766 132 767 136
rect 771 132 772 136
rect 766 131 772 132
rect 926 136 932 137
rect 926 132 927 136
rect 931 132 932 136
rect 926 131 932 132
rect 1094 136 1100 137
rect 1094 132 1095 136
rect 1099 132 1100 136
rect 1094 131 1100 132
rect 1262 136 1268 137
rect 1262 132 1263 136
rect 1267 132 1268 136
rect 1262 131 1268 132
rect 1438 136 1444 137
rect 1438 132 1439 136
rect 1443 132 1444 136
rect 1438 131 1444 132
rect 1598 136 1604 137
rect 1598 132 1599 136
rect 1603 132 1604 136
rect 1598 131 1604 132
rect 1718 135 1724 136
rect 1718 131 1719 135
rect 1723 131 1724 135
rect 110 130 116 131
rect 112 107 114 130
rect 336 107 338 131
rect 472 107 474 131
rect 616 107 618 131
rect 768 107 770 131
rect 928 107 930 131
rect 1096 107 1098 131
rect 1264 107 1266 131
rect 1440 107 1442 131
rect 1600 107 1602 131
rect 1718 130 1724 131
rect 1720 107 1722 130
rect 111 106 115 107
rect 111 101 115 102
rect 335 106 339 107
rect 335 101 339 102
rect 471 106 475 107
rect 471 101 475 102
rect 615 106 619 107
rect 615 101 619 102
rect 767 106 771 107
rect 767 101 771 102
rect 927 106 931 107
rect 927 101 931 102
rect 1095 106 1099 107
rect 1095 101 1099 102
rect 1263 106 1267 107
rect 1263 101 1267 102
rect 1439 106 1443 107
rect 1439 101 1443 102
rect 1599 106 1603 107
rect 1599 101 1603 102
rect 1719 106 1723 107
rect 1719 101 1723 102
<< m4c >>
rect 111 1774 115 1778
rect 135 1774 139 1778
rect 271 1774 275 1778
rect 407 1774 411 1778
rect 543 1774 547 1778
rect 679 1774 683 1778
rect 1719 1774 1723 1778
rect 111 1658 115 1662
rect 159 1658 163 1662
rect 247 1658 251 1662
rect 295 1658 299 1662
rect 383 1658 387 1662
rect 431 1658 435 1662
rect 519 1658 523 1662
rect 567 1658 571 1662
rect 655 1658 659 1662
rect 703 1658 707 1662
rect 307 1624 311 1628
rect 791 1658 795 1662
rect 1719 1658 1723 1662
rect 767 1624 771 1628
rect 111 1546 115 1550
rect 223 1546 227 1550
rect 359 1546 363 1550
rect 487 1546 491 1550
rect 495 1546 499 1550
rect 623 1546 627 1550
rect 631 1546 635 1550
rect 759 1546 763 1550
rect 767 1546 771 1550
rect 895 1546 899 1550
rect 1031 1546 1035 1550
rect 1167 1546 1171 1550
rect 1303 1546 1307 1550
rect 1439 1546 1443 1550
rect 1575 1546 1579 1550
rect 1719 1546 1723 1550
rect 111 1430 115 1434
rect 511 1430 515 1434
rect 647 1430 651 1434
rect 743 1430 747 1434
rect 783 1430 787 1434
rect 887 1430 891 1434
rect 919 1430 923 1434
rect 1031 1430 1035 1434
rect 1055 1430 1059 1434
rect 1175 1430 1179 1434
rect 1191 1430 1195 1434
rect 1319 1430 1323 1434
rect 1327 1430 1331 1434
rect 1463 1430 1467 1434
rect 1599 1430 1603 1434
rect 1719 1430 1723 1434
rect 111 1322 115 1326
rect 183 1322 187 1326
rect 415 1322 419 1326
rect 679 1322 683 1326
rect 719 1322 723 1326
rect 863 1322 867 1326
rect 975 1322 979 1326
rect 1007 1322 1011 1326
rect 1151 1322 1155 1326
rect 1287 1322 1291 1326
rect 1295 1322 1299 1326
rect 111 1218 115 1222
rect 159 1218 163 1222
rect 207 1218 211 1222
rect 335 1218 339 1222
rect 439 1218 443 1222
rect 559 1218 563 1222
rect 703 1218 707 1222
rect 799 1218 803 1222
rect 999 1218 1003 1222
rect 1063 1218 1067 1222
rect 1311 1218 1315 1222
rect 1335 1218 1339 1222
rect 1439 1322 1443 1326
rect 1575 1322 1579 1326
rect 1719 1322 1723 1326
rect 1599 1218 1603 1222
rect 111 1102 115 1106
rect 135 1102 139 1106
rect 223 1102 227 1106
rect 311 1102 315 1106
rect 463 1102 467 1106
rect 535 1102 539 1106
rect 719 1102 723 1106
rect 775 1102 779 1106
rect 991 1102 995 1106
rect 1039 1102 1043 1106
rect 1271 1102 1275 1106
rect 1311 1102 1315 1106
rect 1559 1102 1563 1106
rect 1575 1102 1579 1106
rect 111 1002 115 1006
rect 247 1002 251 1006
rect 463 1002 467 1006
rect 487 1002 491 1006
rect 647 1002 651 1006
rect 743 1002 747 1006
rect 855 1002 859 1006
rect 1015 1002 1019 1006
rect 1079 1002 1083 1006
rect 1295 1002 1299 1006
rect 1311 1002 1315 1006
rect 111 894 115 898
rect 439 894 443 898
rect 623 894 627 898
rect 687 894 691 898
rect 823 894 827 898
rect 831 894 835 898
rect 959 894 963 898
rect 1055 894 1059 898
rect 1095 894 1099 898
rect 1231 894 1235 898
rect 1287 894 1291 898
rect 1367 894 1371 898
rect 1719 1218 1723 1222
rect 1719 1102 1723 1106
rect 1543 1002 1547 1006
rect 1583 1002 1587 1006
rect 1503 894 1507 898
rect 1519 894 1523 898
rect 111 782 115 786
rect 711 782 715 786
rect 815 782 819 786
rect 847 782 851 786
rect 951 782 955 786
rect 983 782 987 786
rect 1087 782 1091 786
rect 1119 782 1123 786
rect 1223 782 1227 786
rect 1255 782 1259 786
rect 875 699 879 700
rect 875 696 879 699
rect 111 674 115 678
rect 511 674 515 678
rect 679 674 683 678
rect 791 674 795 678
rect 855 674 859 678
rect 927 674 931 678
rect 1099 696 1103 700
rect 1359 782 1363 786
rect 1391 782 1395 786
rect 1719 1002 1723 1006
rect 1719 894 1723 898
rect 1495 782 1499 786
rect 1527 782 1531 786
rect 1031 674 1035 678
rect 1063 674 1067 678
rect 1199 674 1203 678
rect 1215 674 1219 678
rect 111 554 115 558
rect 167 554 171 558
rect 359 554 363 558
rect 535 554 539 558
rect 551 554 555 558
rect 703 554 707 558
rect 743 554 747 558
rect 111 430 115 434
rect 135 430 139 434
rect 143 430 147 434
rect 879 554 883 558
rect 935 554 939 558
rect 1055 554 1059 558
rect 1127 554 1131 558
rect 1335 674 1339 678
rect 1407 674 1411 678
rect 1471 674 1475 678
rect 1719 782 1723 786
rect 1719 674 1723 678
rect 1239 554 1243 558
rect 1327 554 1331 558
rect 1431 554 1435 558
rect 335 430 339 434
rect 351 430 355 434
rect 527 430 531 434
rect 615 430 619 434
rect 719 430 723 434
rect 895 430 899 434
rect 911 430 915 434
rect 1103 430 1107 434
rect 1183 430 1187 434
rect 111 322 115 326
rect 159 322 163 326
rect 223 322 227 326
rect 375 322 379 326
rect 455 322 459 326
rect 639 322 643 326
rect 687 322 691 326
rect 919 322 923 326
rect 111 202 115 206
rect 199 202 203 206
rect 1151 322 1155 326
rect 1207 322 1211 326
rect 1527 554 1531 558
rect 1719 554 1723 558
rect 1303 430 1307 434
rect 1471 430 1475 434
rect 1503 430 1507 434
rect 1719 430 1723 434
rect 1383 322 1387 326
rect 1495 322 1499 326
rect 311 202 315 206
rect 431 202 435 206
rect 447 202 451 206
rect 591 202 595 206
rect 663 202 667 206
rect 743 202 747 206
rect 895 202 899 206
rect 903 202 907 206
rect 1071 202 1075 206
rect 1127 202 1131 206
rect 1239 202 1243 206
rect 1599 322 1603 326
rect 1719 322 1723 326
rect 1359 202 1363 206
rect 1415 202 1419 206
rect 1575 202 1579 206
rect 1719 202 1723 206
rect 111 102 115 106
rect 335 102 339 106
rect 471 102 475 106
rect 615 102 619 106
rect 767 102 771 106
rect 927 102 931 106
rect 1095 102 1099 106
rect 1263 102 1267 106
rect 1439 102 1443 106
rect 1599 102 1603 106
rect 1719 102 1723 106
<< m4 >>
rect 96 1773 97 1779
rect 103 1778 1755 1779
rect 103 1774 111 1778
rect 115 1774 135 1778
rect 139 1774 271 1778
rect 275 1774 407 1778
rect 411 1774 543 1778
rect 547 1774 679 1778
rect 683 1774 1719 1778
rect 1723 1774 1755 1778
rect 103 1773 1755 1774
rect 1761 1773 1762 1779
rect 84 1657 85 1663
rect 91 1662 1743 1663
rect 91 1658 111 1662
rect 115 1658 159 1662
rect 163 1658 247 1662
rect 251 1658 295 1662
rect 299 1658 383 1662
rect 387 1658 431 1662
rect 435 1658 519 1662
rect 523 1658 567 1662
rect 571 1658 655 1662
rect 659 1658 703 1662
rect 707 1658 791 1662
rect 795 1658 1719 1662
rect 1723 1658 1743 1662
rect 91 1657 1743 1658
rect 1749 1657 1750 1663
rect 306 1628 312 1629
rect 766 1628 772 1629
rect 306 1624 307 1628
rect 311 1624 767 1628
rect 771 1624 772 1628
rect 306 1623 312 1624
rect 766 1623 772 1624
rect 96 1545 97 1551
rect 103 1550 1755 1551
rect 103 1546 111 1550
rect 115 1546 223 1550
rect 227 1546 359 1550
rect 363 1546 487 1550
rect 491 1546 495 1550
rect 499 1546 623 1550
rect 627 1546 631 1550
rect 635 1546 759 1550
rect 763 1546 767 1550
rect 771 1546 895 1550
rect 899 1546 1031 1550
rect 1035 1546 1167 1550
rect 1171 1546 1303 1550
rect 1307 1546 1439 1550
rect 1443 1546 1575 1550
rect 1579 1546 1719 1550
rect 1723 1546 1755 1550
rect 103 1545 1755 1546
rect 1761 1545 1762 1551
rect 84 1429 85 1435
rect 91 1434 1743 1435
rect 91 1430 111 1434
rect 115 1430 511 1434
rect 515 1430 647 1434
rect 651 1430 743 1434
rect 747 1430 783 1434
rect 787 1430 887 1434
rect 891 1430 919 1434
rect 923 1430 1031 1434
rect 1035 1430 1055 1434
rect 1059 1430 1175 1434
rect 1179 1430 1191 1434
rect 1195 1430 1319 1434
rect 1323 1430 1327 1434
rect 1331 1430 1463 1434
rect 1467 1430 1599 1434
rect 1603 1430 1719 1434
rect 1723 1430 1743 1434
rect 91 1429 1743 1430
rect 1749 1429 1750 1435
rect 96 1321 97 1327
rect 103 1326 1755 1327
rect 103 1322 111 1326
rect 115 1322 183 1326
rect 187 1322 415 1326
rect 419 1322 679 1326
rect 683 1322 719 1326
rect 723 1322 863 1326
rect 867 1322 975 1326
rect 979 1322 1007 1326
rect 1011 1322 1151 1326
rect 1155 1322 1287 1326
rect 1291 1322 1295 1326
rect 1299 1322 1439 1326
rect 1443 1322 1575 1326
rect 1579 1322 1719 1326
rect 1723 1322 1755 1326
rect 103 1321 1755 1322
rect 1761 1321 1762 1327
rect 84 1217 85 1223
rect 91 1222 1743 1223
rect 91 1218 111 1222
rect 115 1218 159 1222
rect 163 1218 207 1222
rect 211 1218 335 1222
rect 339 1218 439 1222
rect 443 1218 559 1222
rect 563 1218 703 1222
rect 707 1218 799 1222
rect 803 1218 999 1222
rect 1003 1218 1063 1222
rect 1067 1218 1311 1222
rect 1315 1218 1335 1222
rect 1339 1218 1599 1222
rect 1603 1218 1719 1222
rect 1723 1218 1743 1222
rect 91 1217 1743 1218
rect 1749 1217 1750 1223
rect 96 1101 97 1107
rect 103 1106 1755 1107
rect 103 1102 111 1106
rect 115 1102 135 1106
rect 139 1102 223 1106
rect 227 1102 311 1106
rect 315 1102 463 1106
rect 467 1102 535 1106
rect 539 1102 719 1106
rect 723 1102 775 1106
rect 779 1102 991 1106
rect 995 1102 1039 1106
rect 1043 1102 1271 1106
rect 1275 1102 1311 1106
rect 1315 1102 1559 1106
rect 1563 1102 1575 1106
rect 1579 1102 1719 1106
rect 1723 1102 1755 1106
rect 103 1101 1755 1102
rect 1761 1101 1762 1107
rect 84 1001 85 1007
rect 91 1006 1743 1007
rect 91 1002 111 1006
rect 115 1002 247 1006
rect 251 1002 463 1006
rect 467 1002 487 1006
rect 491 1002 647 1006
rect 651 1002 743 1006
rect 747 1002 855 1006
rect 859 1002 1015 1006
rect 1019 1002 1079 1006
rect 1083 1002 1295 1006
rect 1299 1002 1311 1006
rect 1315 1002 1543 1006
rect 1547 1002 1583 1006
rect 1587 1002 1719 1006
rect 1723 1002 1743 1006
rect 91 1001 1743 1002
rect 1749 1001 1750 1007
rect 96 893 97 899
rect 103 898 1755 899
rect 103 894 111 898
rect 115 894 439 898
rect 443 894 623 898
rect 627 894 687 898
rect 691 894 823 898
rect 827 894 831 898
rect 835 894 959 898
rect 963 894 1055 898
rect 1059 894 1095 898
rect 1099 894 1231 898
rect 1235 894 1287 898
rect 1291 894 1367 898
rect 1371 894 1503 898
rect 1507 894 1519 898
rect 1523 894 1719 898
rect 1723 894 1755 898
rect 103 893 1755 894
rect 1761 893 1762 899
rect 84 781 85 787
rect 91 786 1743 787
rect 91 782 111 786
rect 115 782 711 786
rect 715 782 815 786
rect 819 782 847 786
rect 851 782 951 786
rect 955 782 983 786
rect 987 782 1087 786
rect 1091 782 1119 786
rect 1123 782 1223 786
rect 1227 782 1255 786
rect 1259 782 1359 786
rect 1363 782 1391 786
rect 1395 782 1495 786
rect 1499 782 1527 786
rect 1531 782 1719 786
rect 1723 782 1743 786
rect 91 781 1743 782
rect 1749 781 1750 787
rect 874 700 880 701
rect 1098 700 1104 701
rect 874 696 875 700
rect 879 696 1099 700
rect 1103 696 1104 700
rect 874 695 880 696
rect 1098 695 1104 696
rect 96 673 97 679
rect 103 678 1755 679
rect 103 674 111 678
rect 115 674 511 678
rect 515 674 679 678
rect 683 674 791 678
rect 795 674 855 678
rect 859 674 927 678
rect 931 674 1031 678
rect 1035 674 1063 678
rect 1067 674 1199 678
rect 1203 674 1215 678
rect 1219 674 1335 678
rect 1339 674 1407 678
rect 1411 674 1471 678
rect 1475 674 1719 678
rect 1723 674 1755 678
rect 103 673 1755 674
rect 1761 673 1762 679
rect 84 553 85 559
rect 91 558 1743 559
rect 91 554 111 558
rect 115 554 167 558
rect 171 554 359 558
rect 363 554 535 558
rect 539 554 551 558
rect 555 554 703 558
rect 707 554 743 558
rect 747 554 879 558
rect 883 554 935 558
rect 939 554 1055 558
rect 1059 554 1127 558
rect 1131 554 1239 558
rect 1243 554 1327 558
rect 1331 554 1431 558
rect 1435 554 1527 558
rect 1531 554 1719 558
rect 1723 554 1743 558
rect 91 553 1743 554
rect 1749 553 1750 559
rect 96 429 97 435
rect 103 434 1755 435
rect 103 430 111 434
rect 115 430 135 434
rect 139 430 143 434
rect 147 430 335 434
rect 339 430 351 434
rect 355 430 527 434
rect 531 430 615 434
rect 619 430 719 434
rect 723 430 895 434
rect 899 430 911 434
rect 915 430 1103 434
rect 1107 430 1183 434
rect 1187 430 1303 434
rect 1307 430 1471 434
rect 1475 430 1503 434
rect 1507 430 1719 434
rect 1723 430 1755 434
rect 103 429 1755 430
rect 1761 429 1762 435
rect 84 321 85 327
rect 91 326 1743 327
rect 91 322 111 326
rect 115 322 159 326
rect 163 322 223 326
rect 227 322 375 326
rect 379 322 455 326
rect 459 322 639 326
rect 643 322 687 326
rect 691 322 919 326
rect 923 322 1151 326
rect 1155 322 1207 326
rect 1211 322 1383 326
rect 1387 322 1495 326
rect 1499 322 1599 326
rect 1603 322 1719 326
rect 1723 322 1743 326
rect 91 321 1743 322
rect 1749 321 1750 327
rect 96 201 97 207
rect 103 206 1755 207
rect 103 202 111 206
rect 115 202 199 206
rect 203 202 311 206
rect 315 202 431 206
rect 435 202 447 206
rect 451 202 591 206
rect 595 202 663 206
rect 667 202 743 206
rect 747 202 895 206
rect 899 202 903 206
rect 907 202 1071 206
rect 1075 202 1127 206
rect 1131 202 1239 206
rect 1243 202 1359 206
rect 1363 202 1415 206
rect 1419 202 1575 206
rect 1579 202 1719 206
rect 1723 202 1755 206
rect 103 201 1755 202
rect 1761 201 1762 207
rect 84 101 85 107
rect 91 106 1743 107
rect 91 102 111 106
rect 115 102 335 106
rect 339 102 471 106
rect 475 102 615 106
rect 619 102 767 106
rect 771 102 927 106
rect 931 102 1095 106
rect 1099 102 1263 106
rect 1267 102 1439 106
rect 1443 102 1599 106
rect 1603 102 1719 106
rect 1723 102 1743 106
rect 91 101 1743 102
rect 1749 101 1750 107
<< m5c >>
rect 97 1773 103 1779
rect 1755 1773 1761 1779
rect 85 1657 91 1663
rect 1743 1657 1749 1663
rect 97 1545 103 1551
rect 1755 1545 1761 1551
rect 85 1429 91 1435
rect 1743 1429 1749 1435
rect 97 1321 103 1327
rect 1755 1321 1761 1327
rect 85 1217 91 1223
rect 1743 1217 1749 1223
rect 97 1101 103 1107
rect 1755 1101 1761 1107
rect 85 1001 91 1007
rect 1743 1001 1749 1007
rect 97 893 103 899
rect 1755 893 1761 899
rect 85 781 91 787
rect 1743 781 1749 787
rect 97 673 103 679
rect 1755 673 1761 679
rect 85 553 91 559
rect 1743 553 1749 559
rect 97 429 103 435
rect 1755 429 1761 435
rect 85 321 91 327
rect 1743 321 1749 327
rect 97 201 103 207
rect 1755 201 1761 207
rect 85 101 91 107
rect 1743 101 1749 107
<< m5 >>
rect 84 1663 92 1800
rect 84 1657 85 1663
rect 91 1657 92 1663
rect 84 1435 92 1657
rect 84 1429 85 1435
rect 91 1429 92 1435
rect 84 1223 92 1429
rect 84 1217 85 1223
rect 91 1217 92 1223
rect 84 1007 92 1217
rect 84 1001 85 1007
rect 91 1001 92 1007
rect 84 787 92 1001
rect 84 781 85 787
rect 91 781 92 787
rect 84 559 92 781
rect 84 553 85 559
rect 91 553 92 559
rect 84 327 92 553
rect 84 321 85 327
rect 91 321 92 327
rect 84 107 92 321
rect 84 101 85 107
rect 91 101 92 107
rect 84 72 92 101
rect 96 1779 104 1800
rect 96 1773 97 1779
rect 103 1773 104 1779
rect 96 1551 104 1773
rect 96 1545 97 1551
rect 103 1545 104 1551
rect 96 1327 104 1545
rect 96 1321 97 1327
rect 103 1321 104 1327
rect 96 1107 104 1321
rect 96 1101 97 1107
rect 103 1101 104 1107
rect 96 899 104 1101
rect 96 893 97 899
rect 103 893 104 899
rect 96 679 104 893
rect 96 673 97 679
rect 103 673 104 679
rect 96 435 104 673
rect 96 429 97 435
rect 103 429 104 435
rect 96 207 104 429
rect 96 201 97 207
rect 103 201 104 207
rect 96 72 104 201
rect 1742 1663 1750 1800
rect 1742 1657 1743 1663
rect 1749 1657 1750 1663
rect 1742 1435 1750 1657
rect 1742 1429 1743 1435
rect 1749 1429 1750 1435
rect 1742 1223 1750 1429
rect 1742 1217 1743 1223
rect 1749 1217 1750 1223
rect 1742 1007 1750 1217
rect 1742 1001 1743 1007
rect 1749 1001 1750 1007
rect 1742 787 1750 1001
rect 1742 781 1743 787
rect 1749 781 1750 787
rect 1742 559 1750 781
rect 1742 553 1743 559
rect 1749 553 1750 559
rect 1742 327 1750 553
rect 1742 321 1743 327
rect 1749 321 1750 327
rect 1742 107 1750 321
rect 1742 101 1743 107
rect 1749 101 1750 107
rect 1742 72 1750 101
rect 1754 1779 1762 1800
rect 1754 1773 1755 1779
rect 1761 1773 1762 1779
rect 1754 1551 1762 1773
rect 1754 1545 1755 1551
rect 1761 1545 1762 1551
rect 1754 1327 1762 1545
rect 1754 1321 1755 1327
rect 1761 1321 1762 1327
rect 1754 1107 1762 1321
rect 1754 1101 1755 1107
rect 1761 1101 1762 1107
rect 1754 899 1762 1101
rect 1754 893 1755 899
rect 1761 893 1762 899
rect 1754 679 1762 893
rect 1754 673 1755 679
rect 1761 673 1762 679
rect 1754 435 1762 673
rect 1754 429 1755 435
rect 1761 429 1762 435
rect 1754 207 1762 429
rect 1754 201 1755 207
rect 1761 201 1762 207
rect 1754 72 1762 201
use welltap_svt  __well_tap__0
timestamp 1730768378
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__0
timestamp 1730768378
transform 1 0 104 0 1 128
box 8 4 12 24
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768378
transform 1 0 304 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_562_6
timestamp 1730768378
transform 1 0 304 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768378
transform 1 0 440 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_563_6
timestamp 1730768378
transform 1 0 440 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768378
transform 1 0 584 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_564_6
timestamp 1730768378
transform 1 0 584 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768378
transform 1 0 736 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_565_6
timestamp 1730768378
transform 1 0 736 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768378
transform 1 0 896 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_566_6
timestamp 1730768378
transform 1 0 896 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768378
transform 1 0 1064 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_567_6
timestamp 1730768378
transform 1 0 1064 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768378
transform 1 0 1232 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_568_6
timestamp 1730768378
transform 1 0 1232 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768378
transform 1 0 1408 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_599_6
timestamp 1730768378
transform 1 0 1408 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768378
transform 1 0 1568 0 1 104
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_598_6
timestamp 1730768378
transform 1 0 1568 0 1 104
box 8 5 126 98
use welltap_svt  __well_tap__1
timestamp 1730768378
transform 1 0 1712 0 1 128
box 8 4 12 24
use welltap_svt  __well_tap__1
timestamp 1730768378
transform 1 0 1712 0 1 128
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768378
transform 1 0 192 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_561_6
timestamp 1730768378
transform 1 0 192 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768378
transform 1 0 424 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_560_6
timestamp 1730768378
transform 1 0 424 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768378
transform 1 0 656 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_559_6
timestamp 1730768378
transform 1 0 656 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768378
transform 1 0 888 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_569_6
timestamp 1730768378
transform 1 0 888 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768378
transform 1 0 1120 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_570_6
timestamp 1730768378
transform 1 0 1120 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768378
transform 1 0 1352 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_596_6
timestamp 1730768378
transform 1 0 1352 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768378
transform 1 0 1568 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_597_6
timestamp 1730768378
transform 1 0 1568 0 -1 324
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768378
transform 1 0 128 0 1 332
box 8 5 126 98
use welltap_svt  __well_tap__2
timestamp 1730768378
transform 1 0 104 0 -1 300
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_555_6
timestamp 1730768378
transform 1 0 128 0 1 332
box 8 5 126 98
use welltap_svt  __well_tap__2
timestamp 1730768378
transform 1 0 104 0 -1 300
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768378
transform 1 0 344 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_556_6
timestamp 1730768378
transform 1 0 344 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768378
transform 1 0 608 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_557_6
timestamp 1730768378
transform 1 0 608 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768378
transform 1 0 888 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_558_6
timestamp 1730768378
transform 1 0 888 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768378
transform 1 0 1176 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_571_6
timestamp 1730768378
transform 1 0 1176 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768378
transform 1 0 1464 0 1 332
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_595_6
timestamp 1730768378
transform 1 0 1464 0 1 332
box 8 5 126 98
use welltap_svt  __well_tap__3
timestamp 1730768378
transform 1 0 1712 0 -1 300
box 8 4 12 24
use welltap_svt  __well_tap__3
timestamp 1730768378
transform 1 0 1712 0 -1 300
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768378
transform 1 0 104 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__4
timestamp 1730768378
transform 1 0 104 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768378
transform 1 0 1712 0 1 356
box 8 4 12 24
use welltap_svt  __well_tap__5
timestamp 1730768378
transform 1 0 1712 0 1 356
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768378
transform 1 0 136 0 -1 556
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768378
transform 1 0 104 0 -1 532
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_554_6
timestamp 1730768378
transform 1 0 136 0 -1 556
box 8 5 126 98
use welltap_svt  __well_tap__6
timestamp 1730768378
transform 1 0 104 0 -1 532
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768378
transform 1 0 328 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_553_6
timestamp 1730768378
transform 1 0 328 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768378
transform 1 0 520 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_552_6
timestamp 1730768378
transform 1 0 520 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768378
transform 1 0 712 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_551_6
timestamp 1730768378
transform 1 0 712 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768378
transform 1 0 904 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_572_6
timestamp 1730768378
transform 1 0 904 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768378
transform 1 0 1096 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_573_6
timestamp 1730768378
transform 1 0 1096 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768378
transform 1 0 1296 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_593_6
timestamp 1730768378
transform 1 0 1296 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768378
transform 1 0 1496 0 -1 556
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_594_6
timestamp 1730768378
transform 1 0 1496 0 -1 556
box 8 5 126 98
use welltap_svt  __well_tap__7
timestamp 1730768378
transform 1 0 1712 0 -1 532
box 8 4 12 24
use welltap_svt  __well_tap__7
timestamp 1730768378
transform 1 0 1712 0 -1 532
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768378
transform 1 0 104 0 1 600
box 8 4 12 24
use welltap_svt  __well_tap__8
timestamp 1730768378
transform 1 0 104 0 1 600
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768378
transform 1 0 504 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_549_6
timestamp 1730768378
transform 1 0 504 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768378
transform 1 0 672 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_550_6
timestamp 1730768378
transform 1 0 672 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768378
transform 1 0 848 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_548_6
timestamp 1730768378
transform 1 0 848 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768378
transform 1 0 1024 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_547_6
timestamp 1730768378
transform 1 0 1024 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768378
transform 1 0 1208 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_574_6
timestamp 1730768378
transform 1 0 1208 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768378
transform 1 0 1400 0 1 576
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_592_6
timestamp 1730768378
transform 1 0 1400 0 1 576
box 8 5 126 98
use welltap_svt  __well_tap__9
timestamp 1730768378
transform 1 0 1712 0 1 600
box 8 4 12 24
use welltap_svt  __well_tap__9
timestamp 1730768378
transform 1 0 1712 0 1 600
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768378
transform 1 0 784 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_545_6
timestamp 1730768378
transform 1 0 784 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768378
transform 1 0 920 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_546_6
timestamp 1730768378
transform 1 0 920 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768378
transform 1 0 1056 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_544_6
timestamp 1730768378
transform 1 0 1056 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768378
transform 1 0 1192 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_543_6
timestamp 1730768378
transform 1 0 1192 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768378
transform 1 0 1328 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_575_6
timestamp 1730768378
transform 1 0 1328 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768378
transform 1 0 1464 0 -1 784
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_591_6
timestamp 1730768378
transform 1 0 1464 0 -1 784
box 8 5 126 98
use welltap_svt  __well_tap__10
timestamp 1730768378
transform 1 0 104 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__10
timestamp 1730768378
transform 1 0 104 0 -1 760
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768378
transform 1 0 680 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_538_6
timestamp 1730768378
transform 1 0 680 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768378
transform 1 0 816 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_539_6
timestamp 1730768378
transform 1 0 816 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768378
transform 1 0 952 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_540_6
timestamp 1730768378
transform 1 0 952 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768378
transform 1 0 1088 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_541_6
timestamp 1730768378
transform 1 0 1088 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768378
transform 1 0 1224 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_542_6
timestamp 1730768378
transform 1 0 1224 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768378
transform 1 0 1360 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_576_6
timestamp 1730768378
transform 1 0 1360 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768378
transform 1 0 1496 0 1 796
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_590_6
timestamp 1730768378
transform 1 0 1496 0 1 796
box 8 5 126 98
use welltap_svt  __well_tap__11
timestamp 1730768378
transform 1 0 1712 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__11
timestamp 1730768378
transform 1 0 1712 0 -1 760
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768378
transform 1 0 104 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__12
timestamp 1730768378
transform 1 0 104 0 1 820
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768378
transform 1 0 432 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_533_6
timestamp 1730768378
transform 1 0 432 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768378
transform 1 0 616 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_534_6
timestamp 1730768378
transform 1 0 616 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768378
transform 1 0 824 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_535_6
timestamp 1730768378
transform 1 0 824 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768378
transform 1 0 1048 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_536_6
timestamp 1730768378
transform 1 0 1048 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768378
transform 1 0 1280 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_537_6
timestamp 1730768378
transform 1 0 1280 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768378
transform 1 0 1512 0 -1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_589_6
timestamp 1730768378
transform 1 0 1512 0 -1 1004
box 8 5 126 98
use welltap_svt  __well_tap__13
timestamp 1730768378
transform 1 0 1712 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__13
timestamp 1730768378
transform 1 0 1712 0 1 820
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730768378
transform 1 0 104 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__14
timestamp 1730768378
transform 1 0 104 0 -1 980
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768378
transform 1 0 216 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_529_6
timestamp 1730768378
transform 1 0 216 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768378
transform 1 0 456 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_530_6
timestamp 1730768378
transform 1 0 456 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768378
transform 1 0 712 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_531_6
timestamp 1730768378
transform 1 0 712 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768378
transform 1 0 984 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_532_6
timestamp 1730768378
transform 1 0 984 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768378
transform 1 0 1264 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_577_6
timestamp 1730768378
transform 1 0 1264 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768378
transform 1 0 1552 0 1 1004
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_588_6
timestamp 1730768378
transform 1 0 1552 0 1 1004
box 8 5 126 98
use welltap_svt  __well_tap__15
timestamp 1730768378
transform 1 0 1712 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__15
timestamp 1730768378
transform 1 0 1712 0 -1 980
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730768378
transform 1 0 104 0 1 1028
box 8 4 12 24
use welltap_svt  __well_tap__16
timestamp 1730768378
transform 1 0 104 0 1 1028
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730768378
transform 1 0 1712 0 1 1028
box 8 4 12 24
use welltap_svt  __well_tap__17
timestamp 1730768378
transform 1 0 1712 0 1 1028
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768378
transform 1 0 128 0 -1 1220
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768378
transform 1 0 104 0 -1 1196
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_524_6
timestamp 1730768378
transform 1 0 128 0 -1 1220
box 8 5 126 98
use welltap_svt  __well_tap__18
timestamp 1730768378
transform 1 0 104 0 -1 1196
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768378
transform 1 0 304 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_525_6
timestamp 1730768378
transform 1 0 304 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768378
transform 1 0 528 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_526_6
timestamp 1730768378
transform 1 0 528 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768378
transform 1 0 768 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_527_6
timestamp 1730768378
transform 1 0 768 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768378
transform 1 0 1032 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_528_6
timestamp 1730768378
transform 1 0 1032 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768378
transform 1 0 1304 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_578_6
timestamp 1730768378
transform 1 0 1304 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768378
transform 1 0 1568 0 -1 1220
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_587_6
timestamp 1730768378
transform 1 0 1568 0 -1 1220
box 8 5 126 98
use welltap_svt  __well_tap__19
timestamp 1730768378
transform 1 0 1712 0 -1 1196
box 8 4 12 24
use welltap_svt  __well_tap__19
timestamp 1730768378
transform 1 0 1712 0 -1 1196
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768378
transform 1 0 176 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768378
transform 1 0 104 0 1 1248
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_523_6
timestamp 1730768378
transform 1 0 176 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__20
timestamp 1730768378
transform 1 0 104 0 1 1248
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768378
transform 1 0 408 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_522_6
timestamp 1730768378
transform 1 0 408 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768378
transform 1 0 672 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_521_6
timestamp 1730768378
transform 1 0 672 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768378
transform 1 0 968 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_520_6
timestamp 1730768378
transform 1 0 968 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768378
transform 1 0 1280 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_519_6
timestamp 1730768378
transform 1 0 1280 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768378
transform 1 0 1568 0 1 1224
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_586_6
timestamp 1730768378
transform 1 0 1568 0 1 1224
box 8 5 126 98
use welltap_svt  __well_tap__21
timestamp 1730768378
transform 1 0 1712 0 1 1248
box 8 4 12 24
use welltap_svt  __well_tap__21
timestamp 1730768378
transform 1 0 1712 0 1 1248
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730768378
transform 1 0 104 0 -1 1408
box 8 4 12 24
use welltap_svt  __well_tap__22
timestamp 1730768378
transform 1 0 104 0 -1 1408
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768378
transform 1 0 712 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_515_6
timestamp 1730768378
transform 1 0 712 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768378
transform 1 0 856 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_516_6
timestamp 1730768378
transform 1 0 856 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768378
transform 1 0 1000 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_517_6
timestamp 1730768378
transform 1 0 1000 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768378
transform 1 0 1144 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_518_6
timestamp 1730768378
transform 1 0 1144 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768378
transform 1 0 1288 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_579_6
timestamp 1730768378
transform 1 0 1288 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768378
transform 1 0 1432 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_584_6
timestamp 1730768378
transform 1 0 1432 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768378
transform 1 0 1568 0 -1 1432
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_585_6
timestamp 1730768378
transform 1 0 1568 0 -1 1432
box 8 5 126 98
use welltap_svt  __well_tap__23
timestamp 1730768378
transform 1 0 1712 0 -1 1408
box 8 4 12 24
use welltap_svt  __well_tap__23
timestamp 1730768378
transform 1 0 1712 0 -1 1408
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768378
transform 1 0 104 0 1 1472
box 8 4 12 24
use welltap_svt  __well_tap__24
timestamp 1730768378
transform 1 0 104 0 1 1472
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768378
transform 1 0 480 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_510_6
timestamp 1730768378
transform 1 0 480 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768378
transform 1 0 616 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_511_6
timestamp 1730768378
transform 1 0 616 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768378
transform 1 0 752 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_512_6
timestamp 1730768378
transform 1 0 752 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768378
transform 1 0 888 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_513_6
timestamp 1730768378
transform 1 0 888 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768378
transform 1 0 1024 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_514_6
timestamp 1730768378
transform 1 0 1024 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768378
transform 1 0 1160 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_580_6
timestamp 1730768378
transform 1 0 1160 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768378
transform 1 0 1296 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_581_6
timestamp 1730768378
transform 1 0 1296 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768378
transform 1 0 1432 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_582_6
timestamp 1730768378
transform 1 0 1432 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768378
transform 1 0 1568 0 1 1448
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_583_6
timestamp 1730768378
transform 1 0 1568 0 1 1448
box 8 5 126 98
use welltap_svt  __well_tap__25
timestamp 1730768378
transform 1 0 1712 0 1 1472
box 8 4 12 24
use welltap_svt  __well_tap__25
timestamp 1730768378
transform 1 0 1712 0 1 1472
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768378
transform 1 0 216 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_55_6
timestamp 1730768378
transform 1 0 216 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768378
transform 1 0 352 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_56_6
timestamp 1730768378
transform 1 0 352 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768378
transform 1 0 488 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_57_6
timestamp 1730768378
transform 1 0 488 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768378
transform 1 0 624 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_58_6
timestamp 1730768378
transform 1 0 624 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768378
transform 1 0 760 0 -1 1660
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_59_6
timestamp 1730768378
transform 1 0 760 0 -1 1660
box 8 5 126 98
use welltap_svt  __well_tap__26
timestamp 1730768378
transform 1 0 104 0 -1 1636
box 8 4 12 24
use welltap_svt  __well_tap__26
timestamp 1730768378
transform 1 0 104 0 -1 1636
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768378
transform 1 0 1712 0 -1 1636
box 8 4 12 24
use welltap_svt  __well_tap__27
timestamp 1730768378
transform 1 0 1712 0 -1 1636
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768378
transform 1 0 128 0 1 1676
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768378
transform 1 0 104 0 1 1700
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_50_6
timestamp 1730768378
transform 1 0 128 0 1 1676
box 8 5 126 98
use welltap_svt  __well_tap__28
timestamp 1730768378
transform 1 0 104 0 1 1700
box 8 4 12 24
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768378
transform 1 0 264 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_51_6
timestamp 1730768378
transform 1 0 264 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768378
transform 1 0 400 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_52_6
timestamp 1730768378
transform 1 0 400 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768378
transform 1 0 536 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_53_6
timestamp 1730768378
transform 1 0 536 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768378
transform 1 0 672 0 1 1676
box 8 5 126 98
use _0_0std_0_0cells_0_0FAX1  fax_54_6
timestamp 1730768378
transform 1 0 672 0 1 1676
box 8 5 126 98
use welltap_svt  __well_tap__29
timestamp 1730768378
transform 1 0 1712 0 1 1700
box 8 4 12 24
use welltap_svt  __well_tap__29
timestamp 1730768378
transform 1 0 1712 0 1 1700
box 8 4 12 24
<< end >>
