VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.600000 BY 0.300000 ;
END CoreSite

LAYER li
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.056250 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.225000 ;
   PITCH 0.600000 0.600000 ;
END li

LAYER mcon
    TYPE CUT ;
    SPACING 0.225000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END mcon

LAYER met1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.150000 ;
   AREA 0.084375 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met1

LAYER v1
    TYPE CUT ;
    SPACING 0.075000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.075000 ;
END v1

LAYER met2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.150000 ;
   AREA 0.073125 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met2

LAYER v2
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v2

LAYER met3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met3

LAYER v3
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.450000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v3

LAYER met4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met4

LAYER v4
    TYPE CUT ;
    SPACING 0.450000 ;
    WIDTH 1.200000 ;
    ENCLOSURE ABOVE 0.150000 0.150000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END v4

LAYER met5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.650000 ;
   AREA 4.005000 ;
   WIDTH 1.650000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 1.650000 ;
   PITCH 3.300000 3.300000 ;
END met5

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA mcon_C DEFAULT
   LAYER li ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER mcon ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END mcon_C

VIA v1_C DEFAULT
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER met2 ;
     RECT -0.225000 -0.150000 0.225000 0.150000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_C

VIA v3_Ch
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Ch

VIA v3_Cv
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER met4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER met5 ;
     RECT -0.750000 -0.750000 0.750000 0.750000 ;
END v4_C

MACRO _0_0std_0_0cells_0_0AND2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0AND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.200000 BY 4.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 1.200000 3.600000 1.500000 3.900000 ;
        RECT 1.275000 3.375000 1.875000 3.600000 ;
        RECT 1.875000 3.375000 2.100000 3.600000 ;
        RECT 2.100000 3.375000 2.175000 3.600000 ;
        END
        ANTENNAGATEAREA 0.202500 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        RECT 0.675000 0.600000 1.275000 0.825000 ;
        RECT 1.275000 0.600000 1.500000 0.825000 ;
        RECT 1.500000 0.600000 1.575000 0.825000 ;
        END
        ANTENNAGATEAREA 0.202500 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 2.850000 3.000000 3.900000 3.225000 ;
        RECT 2.850000 2.850000 3.075000 3.000000 ;
        RECT 2.850000 2.625000 3.075000 2.850000 ;
        RECT 2.850000 1.725000 3.075000 2.625000 ;
        RECT 2.850000 1.500000 3.075000 1.725000 ;
        RECT 2.850000 1.425000 3.075000 1.500000 ;
        RECT 3.600000 3.225000 3.900000 3.300000 ;
        END
        ANTENNADIFFAREA 0.393750 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 1.275000 2.850000 1.500000 2.925000 ;
        RECT 1.275000 2.625000 1.500000 2.850000 ;
        RECT 1.275000 2.550000 1.500000 2.625000 ;
        RECT 2.325000 2.850000 2.550000 2.925000 ;
        RECT 2.325000 2.625000 2.550000 2.850000 ;
        RECT 2.325000 2.550000 2.550000 2.625000 ;
        LAYER mcon ;
        RECT 1.275000 2.625000 1.500000 2.850000 ;
        RECT 2.325000 2.625000 2.550000 2.850000 ;
        LAYER met1 ;
        RECT 1.200000 2.850000 2.625000 2.925000 ;
        RECT 1.200000 2.625000 1.275000 2.850000 ;
        RECT 1.200000 2.550000 2.625000 2.625000 ;
        RECT 1.275000 2.625000 1.500000 2.850000 ;
        RECT 1.500000 2.625000 2.325000 2.850000 ;
        RECT 2.325000 2.625000 2.550000 2.850000 ;
        RECT 2.550000 2.625000 2.625000 2.850000 ;
        END
        ANTENNADIFFAREA 0.450000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 2.325000 1.425000 2.550000 1.650000 ;
        RECT 2.325000 1.200000 2.550000 1.425000 ;
        RECT 2.325000 0.975000 2.400000 1.200000 ;
        RECT 2.325000 0.900000 2.700000 0.975000 ;
        RECT 2.325000 1.650000 2.550000 1.725000 ;
        RECT 2.400000 0.975000 2.625000 1.200000 ;
        RECT 2.625000 0.975000 2.700000 1.200000 ;
        LAYER mcon ;
        RECT 2.400000 0.975000 2.625000 1.200000 ;
        LAYER met1 ;
        RECT 2.325000 1.200000 2.700000 1.275000 ;
        RECT 2.325000 0.975000 2.400000 1.200000 ;
        RECT 2.325000 0.900000 2.700000 0.975000 ;
        RECT 2.400000 0.975000 2.625000 1.200000 ;
        RECT 2.625000 0.975000 2.700000 1.200000 ;
        END
        ANTENNADIFFAREA 0.258750 ;
    END GND
    OBS
        LAYER li ;
        RECT 1.275000 2.025000 1.500000 2.100000 ;
        RECT 1.275000 1.800000 1.500000 2.025000 ;
        RECT 1.275000 1.725000 1.500000 1.800000 ;
        RECT 1.275000 1.500000 1.500000 1.725000 ;
        RECT 1.275000 1.425000 1.500000 1.500000 ;
        RECT 1.800000 2.625000 2.025000 2.700000 ;
        RECT 1.800000 2.400000 2.025000 2.625000 ;
        RECT 1.800000 2.025000 2.025000 2.400000 ;
        RECT 1.800000 1.800000 2.025000 2.025000 ;
        RECT 1.800000 1.725000 2.025000 1.800000 ;
        RECT 3.375000 2.025000 3.600000 2.100000 ;
        RECT 3.375000 1.800000 3.600000 2.025000 ;
        RECT 3.375000 1.725000 3.600000 1.800000 ;
        LAYER met1 ;
        RECT 1.200000 2.025000 3.675000 2.100000 ;
        RECT 1.200000 1.800000 1.275000 2.025000 ;
        RECT 1.200000 1.725000 3.675000 1.800000 ;
        RECT 1.275000 1.800000 1.500000 2.025000 ;
        RECT 1.500000 1.800000 1.800000 2.025000 ;
        RECT 1.800000 1.800000 2.025000 2.025000 ;
        RECT 2.025000 1.800000 3.375000 2.025000 ;
        RECT 3.375000 1.800000 3.600000 2.025000 ;
        RECT 3.600000 1.800000 3.675000 2.025000 ;
    END
END _0_0std_0_0cells_0_0AND2X1

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 2.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.525000 1.725000 0.900000 1.800000 ;
        RECT 0.525000 1.500000 0.600000 1.725000 ;
        RECT 0.525000 1.425000 0.900000 1.500000 ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        RECT 0.825000 1.500000 0.900000 1.725000 ;
        LAYER mcon ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        LAYER met1 ;
        RECT 0.525000 1.725000 0.900000 1.800000 ;
        RECT 0.525000 1.500000 0.600000 1.725000 ;
        RECT 0.525000 1.425000 0.900000 1.500000 ;
        RECT 0.600000 1.500000 0.825000 1.725000 ;
        RECT 0.825000 1.500000 0.900000 1.725000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.525000 0.525000 0.900000 0.600000 ;
        RECT 0.525000 0.300000 0.600000 0.525000 ;
        RECT 0.525000 0.225000 0.900000 0.300000 ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        RECT 0.825000 0.300000 0.900000 0.525000 ;
        LAYER mcon ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        LAYER met1 ;
        RECT 0.525000 0.525000 0.900000 0.600000 ;
        RECT 0.525000 0.300000 0.600000 0.525000 ;
        RECT 0.525000 0.225000 0.900000 0.300000 ;
        RECT 0.600000 0.300000 0.825000 0.525000 ;
        RECT 0.825000 0.300000 0.900000 0.525000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 192.600000 BY 194.400000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 192.600000 BY 194.400000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

